$date
  Mon May 13 23:42:35 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_mef $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 1 # key_asc $end
$var reg 1 $ key_desc $end
$var reg 1 % enable_disp $end
$var reg 7 & segmentos[6:0] $end
$scope module uut $end
$var reg 1 ' clk $end
$var reg 1 ( reset $end
$var reg 1 ) key_asc $end
$var reg 1 * key_desc $end
$var reg 1 + enable_disp $end
$var reg 7 , segmentos[6:0] $end
$comment state is not handled $end
$comment secuencia is not handled $end
$var integer 32 - cuenta $end
$var reg 4 . bcd[3:0] $end
$scope module a $end
$var reg 1 / clk $end
$var reg 1 0 reset $end
$var reg 1 1 enable $end
$var reg 1 2 cout $end
$var integer 32 3 q $end
$upscope $end
$scope module b $end
$var reg 7 4 segmentos[6:0] $end
$var reg 4 5 bcd[3:0] $end
$var reg 1 6 enable $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
U#
U$
0%
b1001111 &
0'
0(
U)
U*
0+
b1001111 ,
b0 -
b0001 .
0/
00
11
U2
b0 3
b1001111 4
b0001 5
06
#10000000
1!
1'
1/
02
#20000000
0!
0'
b1 -
0/
b1 3
#30000000
1!
1'
1/
#40000000
0!
0'
b10 -
0/
b10 3
#50000000
1!
1'
1/
#60000000
0!
0'
b11 -
0/
b11 3
#70000000
1!
1'
1/
12
#80000000
0!
0'
b100 -
0/
b100 3
#90000000
1!
1'
1/
#100000000
0!
0'
b101 -
0/
b101 3
#110000000
1!
1'
1/
#120000000
0!
0'
b110 -
0/
b110 3
#130000000
1!
1'
1/
#140000000
0!
0'
b111 -
0/
b111 3
#150000000
1!
b0010010 &
1'
b0010010 ,
b0010 .
1/
02
b0010010 4
b0010 5
#160000000
0!
0'
b0 -
0/
b0 3
#170000000
1!
1'
1/
#180000000
0!
0'
b1 -
0/
b1 3
#190000000
1!
1'
1/
#200000000
0!
1#
0'
1)
b10 -
0/
b10 3
#210000000
1!
1'
1/
#220000000
0!
0'
b11 -
0/
b11 3
#230000000
1!
1'
1/
12
#240000000
0!
0#
0'
0)
b100 -
0/
b100 3
#250000000
1!
1'
1/
#260000000
0!
0'
b101 -
0/
b101 3
#270000000
1!
1'
1/
#280000000
0!
0'
b110 -
0/
b110 3
#290000000
1!
1'
1/
#300000000
0!
0'
b111 -
0/
b111 3
#310000000
1!
b0000110 &
1'
b0000110 ,
b0011 .
1/
02
b0000110 4
b0011 5
#320000000
0!
0'
b0 -
0/
b0 3
#330000000
1!
1'
1/
#340000000
0!
0'
b1 -
0/
b1 3
#350000000
1!
1'
1/
#360000000
0!
0'
b10 -
0/
b10 3
#370000000
1!
1'
1/
#380000000
0!
0'
b11 -
0/
b11 3
#390000000
1!
1'
1/
12
#400000000
0!
0'
b100 -
0/
b100 3
#410000000
1!
1'
1/
#420000000
0!
0'
b101 -
0/
b101 3
#430000000
1!
1'
1/
#440000000
0!
0'
b110 -
0/
b110 3
#450000000
1!
1'
1/
#460000000
0!
0'
b111 -
0/
b111 3
#470000000
1!
b0110001 &
1'
b0110001 ,
b1100 .
1/
02
b0110001 4
b1100 5
#480000000
0!
0'
b0 -
0/
b0 3
#490000000
1!
1'
1/
#500000000
0!
0'
b1 -
0/
b1 3
#510000000
1!
1'
1/
#520000000
0!
1$
0'
1*
b10 -
0/
b10 3
#530000000
1!
1'
1/
#540000000
0!
0'
b11 -
0/
b11 3
#550000000
1!
0$
1'
0*
1/
12
#560000000
0!
0'
b100 -
0/
b100 3
#570000000
1!
1'
1/
#580000000
0!
0'
b101 -
0/
b101 3
#590000000
1!
1'
1/
#600000000
0!
0'
b110 -
0/
b110 3
#610000000
1!
1'
1/
#620000000
0!
0'
b111 -
0/
b111 3
#630000000
1!
1'
1/
02
#640000000
0!
0'
b0 -
0/
b0 3
#650000000
1!
1'
1/
#660000000
0!
0'
b1 -
0/
b1 3
#670000000
1!
1'
1/
#680000000
0!
0'
b10 -
0/
b10 3
#690000000
1!
1'
1/
#700000000
0!
0'
b11 -
0/
b11 3
#710000000
1!
1'
1/
12
#720000000
0!
0'
b100 -
0/
b100 3
#730000000
1!
1'
1/
#740000000
0!
0'
b101 -
0/
b101 3
#750000000
1!
1'
1/
#760000000
0!
0'
b110 -
0/
b110 3
#770000000
1!
1'
1/
#780000000
0!
0'
b111 -
0/
b111 3
#790000000
1!
1'
1/
02
#800000000
0!
0'
b0 -
0/
b0 3
#810000000
1!
1'
1/
#820000000
0!
0'
b1 -
0/
b1 3
#830000000
1!
1'
1/
#840000000
0!
0'
b10 -
0/
b10 3
#850000000
1!
1'
1/
#860000000
0!
0'
b11 -
0/
b11 3
#870000000
1!
1'
1/
12
#880000000
0!
1#
0'
1)
b100 -
0/
b100 3
#890000000
1!
1'
1/
#900000000
0!
0'
b101 -
0/
b101 3
#910000000
1!
1'
1/
#920000000
0!
0#
0'
0)
b110 -
0/
b110 3
#930000000
1!
1'
1/
#940000000
0!
0'
b111 -
0/
b111 3
#950000000
1!
b1001111 &
1'
b1001111 ,
b0001 .
1/
02
b1001111 4
b0001 5
#960000000
0!
0'
b0 -
0/
b0 3
#970000000
1!
1'
1/
#980000000
0!
0'
b1 -
0/
b1 3
#990000000
1!
1'
1/
#1000000000
0!
0'
b10 -
0/
b10 3
#1010000000
1!
1'
1/
#1020000000
0!
0'
b11 -
0/
b11 3
#1030000000
1!
1'
1/
12
#1040000000
0!
0'
b100 -
0/
b100 3
#1050000000
1!
1'
1/
#1060000000
0!
0'
b101 -
0/
b101 3
#1070000000
1!
1'
1/
#1080000000
0!
0'
b110 -
0/
b110 3
#1090000000
1!
1'
1/
#1100000000
0!
0'
b111 -
0/
b111 3
#1110000000
1!
b0010010 &
1'
b0010010 ,
b0010 .
1/
02
b0010010 4
b0010 5
#1120000000
0!
0'
b0 -
0/
b0 3
#1130000000
1!
1'
1/
#1140000000
0!
0'
b1 -
0/
b1 3
#1150000000
1!
1'
1/
#1160000000
0!
0'
b10 -
0/
b10 3
#1170000000
1!
1'
1/
#1180000000
0!
0'
b11 -
0/
b11 3
#1190000000
1!
1'
1/
12
#1200000000
0!
1$
0'
1*
b100 -
0/
b100 3
#1210000000
1!
1'
1/
#1220000000
0!
0'
b101 -
0/
b101 3
#1230000000
1!
0$
1'
0*
1/
#1240000000
0!
0'
b110 -
0/
b110 3
#1250000000
1!
1'
1/
#1260000000
0!
0'
b111 -
0/
b111 3
#1270000000
1!
1'
1/
02
#1280000000
0!
0'
b0 -
0/
b0 3
#1290000000
1!
1'
1/
#1300000000
0!
0'
b1 -
0/
b1 3
#1310000000
1!
1'
1/
#1320000000
0!
0'
b10 -
0/
b10 3
#1330000000
1!
1'
1/
#1340000000
0!
0'
b11 -
0/
b11 3
#1350000000
1!
1'
1/
12
#1360000000
0!
0'
b100 -
0/
b100 3
#1370000000
1!
1'
1/
#1380000000
0!
0'
b101 -
0/
b101 3
#1390000000
1!
1'
1/
#1400000000
0!
0'
b110 -
0/
b110 3
#1410000000
1!
1'
1/
#1420000000
0!
0'
b111 -
0/
b111 3
#1430000000
1!
1'
1/
02
#1440000000
0!
0'
b0 -
0/
b0 3
#1450000000
1!
1'
1/
#1460000000
0!
0'
b1 -
0/
b1 3
#1470000000
1!
1'
1/
#1480000000
0!
0'
b10 -
0/
b10 3
#1490000000
1!
1'
1/
#1500000000
0!
0'
b11 -
0/
b11 3
#1510000000
1!
1'
1/
12
#1520000000
0!
0'
b100 -
0/
b100 3
#1530000000
1!
1'
1/
#1540000000
0!
0'
b101 -
0/
b101 3
#1550000000
1!
1'
1/
#1560000000
0!
1#
0'
1)
b110 -
0/
b110 3
#1570000000
1!
1'
1/
#1580000000
0!
0'
b111 -
0/
b111 3
#1590000000
1!
b0000110 &
1'
b0000110 ,
b0011 .
1/
02
b0000110 4
b0011 5
#1600000000
0!
0#
0'
0)
b0 -
0/
b0 3
#1610000000
1!
1'
1/
#1620000000
0!
0'
b1 -
0/
b1 3
#1630000000
1!
1'
1/
#1640000000
0!
0'
b10 -
0/
b10 3
#1650000000
1!
1'
1/
#1660000000
0!
0'
b11 -
0/
b11 3
#1670000000
1!
1'
1/
12
#1680000000
0!
0'
b100 -
0/
b100 3
#1690000000
1!
1'
1/
#1700000000
0!
0'
b101 -
0/
b101 3
#1710000000
1!
1'
1/
#1720000000
0!
0'
b110 -
0/
b110 3
#1730000000
1!
1'
1/
#1740000000
0!
0'
b111 -
0/
b111 3
#1750000000
1!
b0110001 &
1'
b0110001 ,
b1100 .
1/
02
b0110001 4
b1100 5
#1760000000
0!
0'
b0 -
0/
b0 3
#1770000000
1!
1'
1/
#1780000000
0!
0'
b1 -
0/
b1 3
#1790000000
1!
1'
1/
#1800000000
0!
0'
b10 -
0/
b10 3
#1810000000
1!
1'
1/
#1820000000
0!
0'
b11 -
0/
b11 3
#1830000000
1!
1'
1/
12
#1840000000
0!
0'
b100 -
0/
b100 3
#1850000000
1!
1'
1/
#1860000000
0!
0'
b101 -
0/
b101 3
#1870000000
1!
1'
1/
#1880000000
0!
1$
0'
1*
b110 -
0/
b110 3
#1890000000
1!
1'
1/
#1900000000
0!
0'
b111 -
0/
b111 3
#1910000000
1!
0$
1'
0*
1/
02
#1920000000
0!
0'
b0 -
0/
b0 3
#1930000000
1!
1'
1/
#1940000000
0!
0'
b1 -
0/
b1 3
#1950000000
1!
1'
1/
#1960000000
0!
0'
b10 -
0/
b10 3
#1970000000
1!
1'
1/
#1980000000
0!
0'
b11 -
0/
b11 3
#1990000000
1!
1'
1/
12
#2000000000
0!
0'
b100 -
0/
b100 3
#2010000000
1!
1'
1/
#2020000000
0!
0'
b101 -
0/
b101 3
#2030000000
1!
1'
1/
#2040000000
0!
0'
b110 -
0/
b110 3
#2050000000
1!
1'
1/
#2060000000
0!
0'
b111 -
0/
b111 3
#2070000000
1!
1'
1/
02
#2080000000
0!
0'
b0 -
0/
b0 3
#2090000000
1!
1'
1/
#2100000000
0!
0'
b1 -
0/
b1 3
#2110000000
1!
1'
1/
#2120000000
0!
0'
b10 -
0/
b10 3
#2130000000
1!
1'
1/
#2140000000
0!
0'
b11 -
0/
b11 3
#2150000000
1!
1'
1/
12
#2160000000
0!
0'
b100 -
0/
b100 3
#2170000000
1!
1'
1/
#2180000000
0!
0'
b101 -
0/
b101 3
#2190000000
1!
1'
1/
#2200000000
0!
0'
b110 -
0/
b110 3
#2210000000
1!
1'
1/
#2220000000
0!
0'
b111 -
0/
b111 3
#2230000000
1!
1'
1/
02
#2240000000
0!
1#
0'
1)
b0 -
0/
b0 3
#2250000000
1!
1'
1/
#2260000000
0!
0'
b1 -
0/
b1 3
#2270000000
1!
1'
1/
#2280000000
0!
0#
0'
0)
b10 -
0/
b10 3
#2290000000
1!
1'
1/
#2300000000
0!
0'
b11 -
0/
b11 3
#2310000000
1!
1'
1/
12
#2320000000
0!
0'
b100 -
0/
b100 3
#2330000000
1!
1'
1/
#2340000000
0!
0'
b101 -
0/
b101 3
#2350000000
1!
1'
1/
#2360000000
0!
0'
b110 -
0/
b110 3
#2370000000
1!
1'
1/
#2380000000
0!
0'
b111 -
0/
b111 3
#2390000000
1!
b1001111 &
1'
b1001111 ,
b0001 .
1/
02
b1001111 4
b0001 5
#2400000000
0!
0'
b0 -
0/
b0 3
#2410000000
1!
1'
1/
#2420000000
0!
0'
b1 -
0/
b1 3
#2430000000
1!
1'
1/
#2440000000
0!
0'
b10 -
0/
b10 3
#2450000000
1!
1'
1/
#2460000000
0!
0'
b11 -
0/
b11 3
#2470000000
1!
1'
1/
12
#2480000000
0!
0'
b100 -
0/
b100 3
#2490000000
1!
1'
1/
#2500000000
0!
0'
b101 -
0/
b101 3
#2510000000
1!
1'
1/
#2520000000
0!
0'
b110 -
0/
b110 3
#2530000000
1!
1'
1/
#2540000000
0!
0'
b111 -
0/
b111 3
#2550000000
1!
b0010010 &
1'
b0010010 ,
b0010 .
1/
02
b0010010 4
b0010 5
#2560000000
0!
1$
0'
1*
b0 -
0/
b0 3
#2570000000
1!
1'
1/
#2580000000
0!
0'
b1 -
0/
b1 3
#2590000000
1!
0$
1'
0*
1/
#2600000000
0!
0'
b10 -
0/
b10 3
#2610000000
1!
1'
1/
#2620000000
0!
0'
b11 -
0/
b11 3
#2630000000
1!
1'
1/
12
#2640000000
0!
0'
b100 -
0/
b100 3
#2650000000
1!
1'
1/
#2660000000
0!
0'
b101 -
0/
b101 3
#2670000000
1!
1'
1/
#2680000000
0!
0'
b110 -
0/
b110 3
#2690000000
1!
1'
1/
#2700000000
0!
0'
b111 -
0/
b111 3
#2710000000
1!
1'
1/
02
#2720000000
0!
0'
b0 -
0/
b0 3
#2730000000
1!
1'
1/
#2740000000
0!
0'
b1 -
0/
b1 3
#2750000000
1!
1'
1/
#2760000000
0!
0'
b10 -
0/
b10 3
#2770000000
1!
1'
1/
#2780000000
0!
0'
b11 -
0/
b11 3
#2790000000
1!
1'
1/
12
#2800000000
0!
0'
b100 -
0/
b100 3
#2810000000
1!
1'
1/
#2820000000
0!
0'
b101 -
0/
b101 3
#2830000000
1!
1'
1/
#2840000000
0!
0'
b110 -
0/
b110 3
#2850000000
1!
1'
1/
#2860000000
0!
0'
b111 -
0/
b111 3
#2870000000
1!
1'
1/
02
#2880000000
0!
0'
b0 -
0/
b0 3
#2890000000
1!
1'
1/
#2900000000
0!
0'
b1 -
0/
b1 3
#2910000000
1!
1'
1/
#2920000000
0!
1#
0'
1)
b10 -
0/
b10 3
#2930000000
1!
1'
1/
#2940000000
0!
0'
b11 -
0/
b11 3
#2950000000
1!
1'
1/
12
#2960000000
0!
0#
0'
0)
b100 -
0/
b100 3
#2970000000
1!
1'
1/
#2980000000
0!
0'
b101 -
0/
b101 3
#2990000000
1!
1'
1/
#3000000000
0!
0'
b110 -
0/
b110 3
#3010000000
1!
1'
1/
#3020000000
0!
0'
b111 -
0/
b111 3
#3030000000
1!
b0000110 &
1'
b0000110 ,
b0011 .
1/
02
b0000110 4
b0011 5
#3040000000
0!
0'
b0 -
0/
b0 3
#3050000000
1!
1'
1/
#3060000000
0!
0'
b1 -
0/
b1 3
#3070000000
1!
1'
1/
#3080000000
0!
0'
b10 -
0/
b10 3
#3090000000
1!
1'
1/
#3100000000
0!
0'
b11 -
0/
b11 3
#3110000000
1!
1'
1/
12
#3120000000
0!
0'
b100 -
0/
b100 3
#3130000000
1!
1'
1/
#3140000000
0!
0'
b101 -
0/
b101 3
#3150000000
1!
1'
1/
#3160000000
0!
0'
b110 -
0/
b110 3
#3170000000
1!
1'
1/
#3180000000
0!
0'
b111 -
0/
b111 3
#3190000000
1!
b0110001 &
1'
b0110001 ,
b1100 .
1/
02
b0110001 4
b1100 5
#3200000000
0!
0'
b0 -
0/
b0 3
#3210000000
1!
1'
1/
#3220000000
0!
0'
b1 -
0/
b1 3
#3230000000
1!
1'
1/
#3240000000
0!
1$
0'
1*
b10 -
0/
b10 3
#3250000000
1!
1'
1/
#3260000000
0!
0'
b11 -
0/
b11 3
#3270000000
1!
0$
1'
0*
1/
12
#3280000000
0!
0'
b100 -
0/
b100 3
#3290000000
1!
1'
1/
#3300000000
0!
0'
b101 -
0/
b101 3
#3310000000
1!
1'
1/
#3320000000
0!
0'
b110 -
0/
b110 3
#3330000000
1!
1'
1/
#3340000000
0!
0'
b111 -
0/
b111 3
#3350000000
1!
1'
1/
02
#3360000000
0!
0'
b0 -
0/
b0 3
#3370000000
1!
1'
1/
#3380000000
0!
0'
b1 -
0/
b1 3
#3390000000
1!
1'
1/
#3400000000
0!
0'
b10 -
0/
b10 3
#3410000000
1!
1'
1/
#3420000000
0!
0'
b11 -
0/
b11 3
#3430000000
1!
1'
1/
12
#3440000000
0!
0'
b100 -
0/
b100 3
#3450000000
1!
1'
1/
#3460000000
0!
0'
b101 -
0/
b101 3
#3470000000
1!
1'
1/
#3480000000
0!
0'
b110 -
0/
b110 3
#3490000000
1!
1'
1/
#3500000000
0!
0'
b111 -
0/
b111 3
#3510000000
1!
1'
1/
02
#3520000000
0!
0'
b0 -
0/
b0 3
#3530000000
1!
1'
1/
#3540000000
0!
0'
b1 -
0/
b1 3
#3550000000
1!
1'
1/
#3560000000
0!
0'
b10 -
0/
b10 3
#3570000000
1!
1'
1/
#3580000000
0!
0'
b11 -
0/
b11 3
#3590000000
1!
1'
1/
12
#3600000000
0!
1#
0'
1)
b100 -
0/
b100 3
#3610000000
1!
1'
1/
#3620000000
0!
0'
b101 -
0/
b101 3
#3630000000
1!
1'
1/
#3640000000
0!
0#
0'
0)
b110 -
0/
b110 3
#3650000000
1!
1'
1/
#3660000000
0!
0'
b111 -
0/
b111 3
#3670000000
1!
b1001111 &
1'
b1001111 ,
b0001 .
1/
02
b1001111 4
b0001 5
#3680000000
0!
0'
b0 -
0/
b0 3
#3690000000
1!
1'
1/
#3700000000
0!
0'
b1 -
0/
b1 3
#3710000000
1!
1'
1/
#3720000000
0!
0'
b10 -
0/
b10 3
#3730000000
1!
1'
1/
#3740000000
0!
0'
b11 -
0/
b11 3
#3750000000
1!
1'
1/
12
#3760000000
0!
0'
b100 -
0/
b100 3
#3770000000
1!
1'
1/
#3780000000
0!
0'
b101 -
0/
b101 3
#3790000000
1!
1'
1/
#3800000000
0!
0'
b110 -
0/
b110 3
#3810000000
1!
1'
1/
#3820000000
0!
0'
b111 -
0/
b111 3
#3830000000
1!
b0010010 &
1'
b0010010 ,
b0010 .
1/
02
b0010010 4
b0010 5
#3840000000
0!
0'
b0 -
0/
b0 3
#3850000000
1!
1'
1/
#3860000000
0!
0'
b1 -
0/
b1 3
#3870000000
1!
1'
1/
#3880000000
0!
0'
b10 -
0/
b10 3
#3890000000
1!
1'
1/
#3900000000
0!
0'
b11 -
0/
b11 3
#3910000000
1!
1'
1/
12
#3920000000
0!
1$
0'
1*
b100 -
0/
b100 3
#3930000000
1!
1'
1/
#3940000000
0!
0'
b101 -
0/
b101 3
#3950000000
1!
0$
1'
0*
1/
#3960000000
0!
0'
b110 -
0/
b110 3
#3970000000
1!
1'
1/
#3980000000
0!
0'
b111 -
0/
b111 3
#3990000000
1!
1'
1/
02
#4000000000
0!
0'
b0 -
0/
b0 3
#4010000000
1!
1'
1/
#4020000000
0!
0'
b1 -
0/
b1 3
#4030000000
1!
1'
1/
#4040000000
0!
0'
b10 -
0/
b10 3
#4050000000
1!
1'
1/
#4060000000
0!
0'
b11 -
0/
b11 3
#4070000000
1!
1'
1/
12
#4080000000
0!
0'
b100 -
0/
b100 3
#4090000000
1!
1'
1/
#4100000000
0!
0'
b101 -
0/
b101 3
#4110000000
1!
1'
1/
#4120000000
0!
0'
b110 -
0/
b110 3
#4130000000
1!
1'
1/
#4140000000
0!
0'
b111 -
0/
b111 3
#4150000000
1!
1'
1/
02
#4160000000
0!
0'
b0 -
0/
b0 3
#4170000000
1!
1'
1/
#4180000000
0!
0'
b1 -
0/
b1 3
#4190000000
1!
1'
1/
#4200000000
0!
0'
b10 -
0/
b10 3
#4210000000
1!
1'
1/
#4220000000
0!
0'
b11 -
0/
b11 3
#4230000000
1!
1'
1/
12
#4240000000
0!
0'
b100 -
0/
b100 3
#4250000000
1!
1'
1/
#4260000000
0!
0'
b101 -
0/
b101 3
#4270000000
1!
1'
1/
#4280000000
0!
1#
0'
1)
b110 -
0/
b110 3
#4290000000
1!
1'
1/
#4300000000
0!
0'
b111 -
0/
b111 3
#4310000000
1!
b0000110 &
1'
b0000110 ,
b0011 .
1/
02
b0000110 4
b0011 5
#4320000000
0!
0#
0'
0)
b0 -
0/
b0 3
#4330000000
1!
1'
1/
#4340000000
0!
0'
b1 -
0/
b1 3
#4350000000
1!
1'
1/
#4360000000
0!
0'
b10 -
0/
b10 3
#4370000000
1!
1'
1/
#4380000000
0!
0'
b11 -
0/
b11 3
#4390000000
1!
1'
1/
12
#4400000000
0!
0'
b100 -
0/
b100 3
#4410000000
1!
1'
1/
#4420000000
0!
0'
b101 -
0/
b101 3
#4430000000
1!
1'
1/
#4440000000
0!
0'
b110 -
0/
b110 3
#4450000000
1!
1'
1/
#4460000000
0!
0'
b111 -
0/
b111 3
#4470000000
1!
b0110001 &
1'
b0110001 ,
b1100 .
1/
02
b0110001 4
b1100 5
#4480000000
0!
0'
b0 -
0/
b0 3
#4490000000
1!
1'
1/
#4500000000
0!
0'
b1 -
0/
b1 3
#4510000000
1!
1'
1/
#4520000000
0!
0'
b10 -
0/
b10 3
#4530000000
1!
1'
1/
#4540000000
0!
0'
b11 -
0/
b11 3
#4550000000
1!
1'
1/
12
#4560000000
0!
0'
b100 -
0/
b100 3
#4570000000
1!
1'
1/
#4580000000
0!
0'
b101 -
0/
b101 3
#4590000000
1!
1'
1/
#4600000000
0!
1$
0'
1*
b110 -
0/
b110 3
#4610000000
1!
1'
1/
#4620000000
0!
0'
b111 -
0/
b111 3
#4630000000
1!
0$
1'
0*
1/
02
#4640000000
0!
0'
b0 -
0/
b0 3
#4650000000
1!
1'
1/
#4660000000
0!
0'
b1 -
0/
b1 3
#4670000000
1!
1'
1/
#4680000000
0!
0'
b10 -
0/
b10 3
#4690000000
1!
1'
1/
#4700000000
0!
0'
b11 -
0/
b11 3
#4710000000
1!
1'
1/
12
#4720000000
0!
0'
b100 -
0/
b100 3
#4730000000
1!
1'
1/
#4740000000
0!
0'
b101 -
0/
b101 3
#4750000000
1!
1'
1/
#4760000000
0!
0'
b110 -
0/
b110 3
#4770000000
1!
1'
1/
#4780000000
0!
0'
b111 -
0/
b111 3
#4790000000
1!
1'
1/
02
#4800000000
0!
0'
b0 -
0/
b0 3
#4810000000
1!
1'
1/
#4820000000
0!
0'
b1 -
0/
b1 3
#4830000000
1!
1'
1/
#4840000000
0!
0'
b10 -
0/
b10 3
#4850000000
1!
1'
1/
#4860000000
0!
0'
b11 -
0/
b11 3
#4870000000
1!
1'
1/
12
#4880000000
0!
0'
b100 -
0/
b100 3
#4890000000
1!
1'
1/
#4900000000
0!
0'
b101 -
0/
b101 3
#4910000000
1!
1'
1/
#4920000000
0!
0'
b110 -
0/
b110 3
#4930000000
1!
1'
1/
#4940000000
0!
0'
b111 -
0/
b111 3
#4950000000
1!
1'
1/
02
#4960000000
0!
1#
0'
1)
b0 -
0/
b0 3
#4970000000
1!
1'
1/
#4980000000
0!
0'
b1 -
0/
b1 3
#4990000000
1!
1'
1/
#5000000000
0!
0#
0'
0)
b10 -
0/
b10 3
#5010000000
1!
1'
1/
#5020000000
0!
0'
b11 -
0/
b11 3
#5030000000
1!
1'
1/
12
#5040000000
0!
0'
b100 -
0/
b100 3
#5050000000
1!
1'
1/
#5060000000
0!
0'
b101 -
0/
b101 3
#5070000000
1!
1'
1/
#5080000000
0!
0'
b110 -
0/
b110 3
#5090000000
1!
1'
1/
#5100000000
0!
0'
b111 -
0/
b111 3
#5110000000
1!
b1001111 &
1'
b1001111 ,
b0001 .
1/
02
b1001111 4
b0001 5
#5120000000
0!
0'
b0 -
0/
b0 3
#5130000000
1!
1'
1/
#5140000000
0!
0'
b1 -
0/
b1 3
#5150000000
1!
1'
1/
#5160000000
0!
0'
b10 -
0/
b10 3
#5170000000
1!
1'
1/
#5180000000
0!
0'
b11 -
0/
b11 3
#5190000000
1!
1'
1/
12
#5200000000
0!
0'
b100 -
0/
b100 3
#5210000000
1!
1'
1/
#5220000000
0!
0'
b101 -
0/
b101 3
#5230000000
1!
1'
1/
#5240000000
0!
0'
b110 -
0/
b110 3
#5250000000
1!
1'
1/
#5260000000
0!
0'
b111 -
0/
b111 3
#5270000000
1!
b0010010 &
1'
b0010010 ,
b0010 .
1/
02
b0010010 4
b0010 5
#5280000000
0!
1$
0'
1*
b0 -
0/
b0 3
#5290000000
1!
1'
1/
#5300000000
0!
0'
b1 -
0/
b1 3
#5310000000
1!
0$
1'
0*
1/
#5320000000
0!
0'
b10 -
0/
b10 3
#5330000000
1!
1'
1/
#5340000000
0!
0'
b11 -
0/
b11 3
#5350000000
1!
1'
1/
12
#5360000000
0!
0'
b100 -
0/
b100 3
#5370000000
1!
1'
1/
#5380000000
0!
0'
b101 -
0/
b101 3
#5390000000
1!
1'
1/
#5400000000
0!
0'
b110 -
0/
b110 3
#5410000000
1!
1'
1/
#5420000000
0!
0'
b111 -
0/
b111 3
#5430000000
1!
1'
1/
02
#5440000000
0!
0'
b0 -
0/
b0 3
#5450000000
1!
1'
1/
#5460000000
0!
0'
b1 -
0/
b1 3
#5470000000
1!
1'
1/
#5480000000
0!
0'
b10 -
0/
b10 3
#5490000000
1!
1'
1/
#5500000000
0!
0'
b11 -
0/
b11 3
#5510000000
1!
1'
1/
12
#5520000000
0!
0'
b100 -
0/
b100 3
#5530000000
1!
1'
1/
#5540000000
0!
0'
b101 -
0/
b101 3
#5550000000
1!
1'
1/
#5560000000
0!
0'
b110 -
0/
b110 3
#5570000000
1!
1'
1/
#5580000000
0!
0'
b111 -
0/
b111 3
#5590000000
1!
1'
1/
02
#5600000000
0!
0'
b0 -
0/
b0 3
#5610000000
1!
1'
1/
#5620000000
0!
0'
b1 -
0/
b1 3
#5630000000
1!
1'
1/
#5640000000
0!
1#
0'
1)
b10 -
0/
b10 3
#5650000000
1!
1'
1/
#5660000000
0!
0'
b11 -
0/
b11 3
#5670000000
1!
1'
1/
12
#5680000000
0!
0#
0'
0)
b100 -
0/
b100 3
#5690000000
1!
1'
1/
#5700000000
0!
0'
b101 -
0/
b101 3
#5710000000
1!
1'
1/
#5720000000
0!
0'
b110 -
0/
b110 3
#5730000000
1!
1'
1/
#5740000000
0!
0'
b111 -
0/
b111 3
#5750000000
1!
b0000110 &
1'
b0000110 ,
b0011 .
1/
02
b0000110 4
b0011 5
#5760000000
0!
0'
b0 -
0/
b0 3
#5770000000
1!
1'
1/
#5780000000
0!
0'
b1 -
0/
b1 3
#5790000000
1!
1'
1/
#5800000000
0!
0'
b10 -
0/
b10 3
#5810000000
1!
1'
1/
#5820000000
0!
0'
b11 -
0/
b11 3
#5830000000
1!
1'
1/
12
#5840000000
0!
0'
b100 -
0/
b100 3
#5850000000
1!
1'
1/
#5860000000
0!
0'
b101 -
0/
b101 3
#5870000000
1!
1'
1/
#5880000000
0!
0'
b110 -
0/
b110 3
#5890000000
1!
1'
1/
#5900000000
0!
0'
b111 -
0/
b111 3
#5910000000
1!
b0110001 &
1'
b0110001 ,
b1100 .
1/
02
b0110001 4
b1100 5
#5920000000
0!
0'
b0 -
0/
b0 3
#5930000000
1!
1'
1/
#5940000000
0!
0'
b1 -
0/
b1 3
#5950000000
1!
1'
1/
#5960000000
0!
1$
0'
1*
b10 -
0/
b10 3
#5970000000
1!
1'
1/
#5980000000
0!
0'
b11 -
0/
b11 3
#5990000000
1!
0$
1'
0*
1/
12
#6000000000
0!
0'
b100 -
0/
b100 3
#6010000000
1!
1'
1/
#6020000000
0!
0'
b101 -
0/
b101 3
#6030000000
1!
1'
1/
#6040000000
0!
0'
b110 -
0/
b110 3
#6050000000
1!
1'
1/
#6060000000
0!
0'
b111 -
0/
b111 3
#6070000000
1!
1'
1/
02
#6080000000
0!
0'
b0 -
0/
b0 3
#6090000000
1!
1'
1/
#6100000000
0!
0'
b1 -
0/
b1 3
#6110000000
1!
1'
1/
#6120000000
0!
0'
b10 -
0/
b10 3
#6130000000
1!
1'
1/
#6140000000
0!
0'
b11 -
0/
b11 3
#6150000000
1!
1'
1/
12
#6160000000
0!
0'
b100 -
0/
b100 3
#6170000000
1!
1'
1/
#6180000000
0!
0'
b101 -
0/
b101 3
#6190000000
1!
1'
1/
#6200000000
0!
0'
b110 -
0/
b110 3
#6210000000
1!
1'
1/
#6220000000
0!
0'
b111 -
0/
b111 3
#6230000000
1!
1'
1/
02
#6240000000
0!
0'
b0 -
0/
b0 3
#6250000000
1!
1'
1/
#6260000000
0!
0'
b1 -
0/
b1 3
#6270000000
1!
1'
1/
#6280000000
0!
0'
b10 -
0/
b10 3
#6290000000
1!
1'
1/
#6300000000
0!
0'
b11 -
0/
b11 3
#6310000000
1!
1'
1/
12
#6320000000
0!
1#
0'
1)
b100 -
0/
b100 3
#6330000000
1!
1'
1/
#6340000000
0!
0'
b101 -
0/
b101 3
#6350000000
1!
1'
1/
#6360000000
0!
0#
0'
0)
b110 -
0/
b110 3
#6370000000
1!
1'
1/
#6380000000
0!
0'
b111 -
0/
b111 3
#6390000000
1!
b1001111 &
1'
b1001111 ,
b0001 .
1/
02
b1001111 4
b0001 5
#6400000000
0!
0'
b0 -
0/
b0 3
#6410000000
1!
1'
1/
#6420000000
0!
0'
b1 -
0/
b1 3
#6430000000
1!
1'
1/
#6440000000
0!
0'
b10 -
0/
b10 3
#6450000000
1!
1'
1/
#6460000000
0!
0'
b11 -
0/
b11 3
#6470000000
1!
1'
1/
12
#6480000000
0!
0'
b100 -
0/
b100 3
#6490000000
1!
1'
1/
#6500000000
0!
0'
b101 -
0/
b101 3
#6510000000
1!
1'
1/
#6520000000
0!
0'
b110 -
0/
b110 3
#6530000000
1!
1'
1/
#6540000000
0!
0'
b111 -
0/
b111 3
#6550000000
1!
b0010010 &
1'
b0010010 ,
b0010 .
1/
02
b0010010 4
b0010 5
#6560000000
0!
0'
b0 -
0/
b0 3
#6570000000
1!
1'
1/
#6580000000
0!
0'
b1 -
0/
b1 3
#6590000000
1!
1'
1/
#6600000000
0!
0'
b10 -
0/
b10 3
#6610000000
1!
1'
1/
#6620000000
0!
0'
b11 -
0/
b11 3
#6630000000
1!
1'
1/
12
#6640000000
0!
1$
0'
1*
b100 -
0/
b100 3
#6650000000
1!
1'
1/
#6660000000
0!
0'
b101 -
0/
b101 3
#6670000000
1!
0$
1'
0*
1/
#6680000000
0!
0'
b110 -
0/
b110 3
#6690000000
1!
1'
1/
#6700000000
0!
0'
b111 -
0/
b111 3
#6710000000
1!
1'
1/
02
#6720000000
0!
0'
b0 -
0/
b0 3
#6730000000
1!
1'
1/
#6740000000
0!
0'
b1 -
0/
b1 3
#6750000000
1!
1'
1/
#6760000000
0!
0'
b10 -
0/
b10 3
#6770000000
1!
1'
1/
#6780000000
0!
0'
b11 -
0/
b11 3
#6790000000
1!
1'
1/
12
#6800000000
0!
0'
b100 -
0/
b100 3
#6810000000
1!
1'
1/
#6820000000
0!
0'
b101 -
0/
b101 3
#6830000000
1!
1'
1/
#6840000000
0!
0'
b110 -
0/
b110 3
#6850000000
1!
1'
1/
#6860000000
0!
0'
b111 -
0/
b111 3
#6870000000
1!
1'
1/
02
#6880000000
0!
0'
b0 -
0/
b0 3
#6890000000
1!
1'
1/
#6900000000
0!
0'
b1 -
0/
b1 3
#6910000000
1!
1'
1/
#6920000000
0!
0'
b10 -
0/
b10 3
#6930000000
1!
1'
1/
#6940000000
0!
0'
b11 -
0/
b11 3
#6950000000
1!
1'
1/
12
#6960000000
0!
0'
b100 -
0/
b100 3
#6970000000
1!
1'
1/
#6980000000
0!
0'
b101 -
0/
b101 3
#6990000000
1!
1'
1/
#7000000000
0!
1#
0'
1)
b110 -
0/
b110 3
#7010000000
1!
1'
1/
#7020000000
0!
0'
b111 -
0/
b111 3
#7030000000
1!
b0000110 &
1'
b0000110 ,
b0011 .
1/
02
b0000110 4
b0011 5
#7040000000
0!
0#
0'
0)
b0 -
0/
b0 3
#7050000000
1!
1'
1/
#7060000000
0!
0'
b1 -
0/
b1 3
#7070000000
1!
1'
1/
#7080000000
0!
0'
b10 -
0/
b10 3
#7090000000
1!
1'
1/
#7100000000
0!
0'
b11 -
0/
b11 3
#7110000000
1!
1'
1/
12
#7120000000
0!
0'
b100 -
0/
b100 3
#7130000000
1!
1'
1/
#7140000000
0!
0'
b101 -
0/
b101 3
#7150000000
1!
1'
1/
#7160000000
0!
0'
b110 -
0/
b110 3
#7170000000
1!
1'
1/
#7180000000
0!
0'
b111 -
0/
b111 3
#7190000000
1!
b0110001 &
1'
b0110001 ,
b1100 .
1/
02
b0110001 4
b1100 5
#7200000000
0!
0'
b0 -
0/
b0 3
#7210000000
1!
1'
1/
#7220000000
0!
0'
b1 -
0/
b1 3
#7230000000
1!
1'
1/
#7240000000
0!
0'
b10 -
0/
b10 3
#7250000000
1!
1'
1/
#7260000000
0!
0'
b11 -
0/
b11 3
#7270000000
1!
1'
1/
12
#7280000000
0!
0'
b100 -
0/
b100 3
#7290000000
1!
1'
1/
#7300000000
0!
0'
b101 -
0/
b101 3
#7310000000
1!
1'
1/
#7320000000
0!
1$
0'
1*
b110 -
0/
b110 3
#7330000000
1!
1'
1/
#7340000000
0!
0'
b111 -
0/
b111 3
#7350000000
1!
0$
1'
0*
1/
02
#7360000000
0!
0'
b0 -
0/
b0 3
#7370000000
1!
1'
1/
#7380000000
0!
0'
b1 -
0/
b1 3
#7390000000
1!
1'
1/
#7400000000
0!
0'
b10 -
0/
b10 3
#7410000000
1!
1'
1/
#7420000000
0!
0'
b11 -
0/
b11 3
#7430000000
1!
1'
1/
12
#7440000000
0!
0'
b100 -
0/
b100 3
#7450000000
1!
1'
1/
#7460000000
0!
0'
b101 -
0/
b101 3
#7470000000
1!
1'
1/
#7480000000
0!
0'
b110 -
0/
b110 3
#7490000000
1!
1'
1/
#7500000000
0!
0'
b111 -
0/
b111 3
#7510000000
1!
1'
1/
02
#7520000000
0!
0'
b0 -
0/
b0 3
#7530000000
1!
1'
1/
#7540000000
0!
0'
b1 -
0/
b1 3
#7550000000
1!
1'
1/
#7560000000
0!
0'
b10 -
0/
b10 3
#7570000000
1!
1'
1/
#7580000000
0!
0'
b11 -
0/
b11 3
#7590000000
1!
1'
1/
12
#7600000000
0!
0'
b100 -
0/
b100 3
#7610000000
1!
1'
1/
#7620000000
0!
0'
b101 -
0/
b101 3
#7630000000
1!
1'
1/
#7640000000
0!
0'
b110 -
0/
b110 3
#7650000000
1!
1'
1/
#7660000000
0!
0'
b111 -
0/
b111 3
#7670000000
1!
1'
1/
02
#7680000000
0!
1#
0'
1)
b0 -
0/
b0 3
#7690000000
1!
1'
1/
#7700000000
0!
0'
b1 -
0/
b1 3
#7710000000
1!
1'
1/
#7720000000
0!
0#
0'
0)
b10 -
0/
b10 3
#7730000000
1!
1'
1/
#7740000000
0!
0'
b11 -
0/
b11 3
#7750000000
1!
1'
1/
12
#7760000000
0!
0'
b100 -
0/
b100 3
#7770000000
1!
1'
1/
#7780000000
0!
0'
b101 -
0/
b101 3
#7790000000
1!
1'
1/
#7800000000
0!
0'
b110 -
0/
b110 3
#7810000000
1!
1'
1/
#7820000000
0!
0'
b111 -
0/
b111 3
#7830000000
1!
b1001111 &
1'
b1001111 ,
b0001 .
1/
02
b1001111 4
b0001 5
#7840000000
0!
0'
b0 -
0/
b0 3
#7850000000
1!
1'
1/
#7860000000
0!
0'
b1 -
0/
b1 3
#7870000000
1!
1'
1/
#7880000000
0!
0'
b10 -
0/
b10 3
#7890000000
1!
1'
1/
#7900000000
0!
0'
b11 -
0/
b11 3
#7910000000
1!
1'
1/
12
#7920000000
0!
0'
b100 -
0/
b100 3
#7930000000
1!
1'
1/
#7940000000
0!
0'
b101 -
0/
b101 3
#7950000000
1!
1'
1/
#7960000000
0!
0'
b110 -
0/
b110 3
#7970000000
1!
1'
1/
#7980000000
0!
0'
b111 -
0/
b111 3
#7990000000
1!
b0010010 &
1'
b0010010 ,
b0010 .
1/
02
b0010010 4
b0010 5
#8000000000
0!
1$
0'
1*
b0 -
0/
b0 3
#8010000000
1!
1'
1/
#8020000000
0!
0'
b1 -
0/
b1 3
#8030000000
1!
0$
1'
0*
1/
#8040000000
0!
0'
b10 -
0/
b10 3
#8050000000
1!
1'
1/
#8060000000
0!
0'
b11 -
0/
b11 3
#8070000000
1!
1'
1/
12
#8080000000
0!
0'
b100 -
0/
b100 3
#8090000000
1!
1'
1/
#8100000000
0!
0'
b101 -
0/
b101 3
#8110000000
1!
1'
1/
#8120000000
0!
0'
b110 -
0/
b110 3
#8130000000
1!
1'
1/
#8140000000
0!
0'
b111 -
0/
b111 3
#8150000000
1!
1'
1/
02
#8160000000
0!
0'
b0 -
0/
b0 3
#8170000000
1!
1'
1/
#8180000000
0!
0'
b1 -
0/
b1 3
#8190000000
1!
1'
1/
#8200000000
0!
0'
b10 -
0/
b10 3
#8210000000
1!
1'
1/
#8220000000
0!
0'
b11 -
0/
b11 3
#8230000000
1!
1'
1/
12
#8240000000
0!
0'
b100 -
0/
b100 3
#8250000000
1!
1'
1/
#8260000000
0!
0'
b101 -
0/
b101 3
#8270000000
1!
1'
1/
#8280000000
0!
0'
b110 -
0/
b110 3
#8290000000
1!
1'
1/
#8300000000
0!
0'
b111 -
0/
b111 3
#8310000000
1!
1'
1/
02
#8320000000
0!
0'
b0 -
0/
b0 3
#8330000000
1!
1'
1/
#8340000000
0!
0'
b1 -
0/
b1 3
#8350000000
1!
1'
1/
#8360000000
0!
1#
0'
1)
b10 -
0/
b10 3
#8370000000
1!
1'
1/
#8380000000
0!
0'
b11 -
0/
b11 3
#8390000000
1!
1'
1/
12
#8400000000
0!
0#
0'
0)
b100 -
0/
b100 3
#8410000000
1!
1'
1/
#8420000000
0!
0'
b101 -
0/
b101 3
#8430000000
1!
1'
1/
#8440000000
0!
0'
b110 -
0/
b110 3
#8450000000
1!
1'
1/
#8460000000
0!
0'
b111 -
0/
b111 3
#8470000000
1!
b0000110 &
1'
b0000110 ,
b0011 .
1/
02
b0000110 4
b0011 5
#8480000000
0!
0'
b0 -
0/
b0 3
#8490000000
1!
1'
1/
#8500000000
0!
0'
b1 -
0/
b1 3
#8510000000
1!
1'
1/
#8520000000
0!
0'
b10 -
0/
b10 3
#8530000000
1!
1'
1/
#8540000000
0!
0'
b11 -
0/
b11 3
#8550000000
1!
1'
1/
12
#8560000000
0!
0'
b100 -
0/
b100 3
#8570000000
1!
1'
1/
#8580000000
0!
0'
b101 -
0/
b101 3
#8590000000
1!
1'
1/
#8600000000
0!
0'
b110 -
0/
b110 3
#8610000000
1!
1'
1/
#8620000000
0!
0'
b111 -
0/
b111 3
#8630000000
1!
b0110001 &
1'
b0110001 ,
b1100 .
1/
02
b0110001 4
b1100 5
#8640000000
0!
0'
b0 -
0/
b0 3
#8650000000
1!
1'
1/
#8660000000
0!
0'
b1 -
0/
b1 3
#8670000000
1!
1'
1/
#8680000000
0!
1$
0'
1*
b10 -
0/
b10 3
#8690000000
1!
1'
1/
#8700000000
0!
0'
b11 -
0/
b11 3
#8710000000
1!
0$
1'
0*
1/
12
#8720000000
0!
0'
b100 -
0/
b100 3
#8730000000
1!
1'
1/
#8740000000
0!
0'
b101 -
0/
b101 3
#8750000000
1!
1'
1/
#8760000000
0!
0'
b110 -
0/
b110 3
#8770000000
1!
1'
1/
#8780000000
0!
0'
b111 -
0/
b111 3
#8790000000
1!
1'
1/
02
#8800000000
0!
0'
b0 -
0/
b0 3
#8810000000
1!
1'
1/
#8820000000
0!
0'
b1 -
0/
b1 3
#8830000000
1!
1'
1/
#8840000000
0!
0'
b10 -
0/
b10 3
#8850000000
1!
1'
1/
#8860000000
0!
0'
b11 -
0/
b11 3
#8870000000
1!
1'
1/
12
#8880000000
0!
0'
b100 -
0/
b100 3
#8890000000
1!
1'
1/
#8900000000
0!
0'
b101 -
0/
b101 3
#8910000000
1!
1'
1/
#8920000000
0!
0'
b110 -
0/
b110 3
#8930000000
1!
1'
1/
#8940000000
0!
0'
b111 -
0/
b111 3
#8950000000
1!
1'
1/
02
#8960000000
0!
0'
b0 -
0/
b0 3
#8970000000
1!
1'
1/
#8980000000
0!
0'
b1 -
0/
b1 3
#8990000000
1!
1'
1/
#9000000000
0!
0'
b10 -
0/
b10 3
#9010000000
1!
1'
1/
#9020000000
0!
0'
b11 -
0/
b11 3
#9030000000
1!
1'
1/
12
#9040000000
0!
1#
0'
1)
b100 -
0/
b100 3
#9050000000
1!
1'
1/
#9060000000
0!
0'
b101 -
0/
b101 3
#9070000000
1!
1'
1/
#9080000000
0!
0#
0'
0)
b110 -
0/
b110 3
#9090000000
1!
1'
1/
#9100000000
0!
0'
b111 -
0/
b111 3
#9110000000
1!
b1001111 &
1'
b1001111 ,
b0001 .
1/
02
b1001111 4
b0001 5
#9120000000
0!
0'
b0 -
0/
b0 3
#9130000000
1!
1'
1/
#9140000000
0!
0'
b1 -
0/
b1 3
#9150000000
1!
1'
1/
#9160000000
0!
0'
b10 -
0/
b10 3
#9170000000
1!
1'
1/
#9180000000
0!
0'
b11 -
0/
b11 3
#9190000000
1!
1'
1/
12
#9200000000
0!
0'
b100 -
0/
b100 3
#9210000000
1!
1'
1/
#9220000000
0!
0'
b101 -
0/
b101 3
#9230000000
1!
1'
1/
#9240000000
0!
0'
b110 -
0/
b110 3
#9250000000
1!
1'
1/
#9260000000
0!
0'
b111 -
0/
b111 3
#9270000000
1!
b0010010 &
1'
b0010010 ,
b0010 .
1/
02
b0010010 4
b0010 5
#9280000000
0!
0'
b0 -
0/
b0 3
#9290000000
1!
1'
1/
#9300000000
0!
0'
b1 -
0/
b1 3
#9310000000
1!
1'
1/
#9320000000
0!
0'
b10 -
0/
b10 3
#9330000000
1!
1'
1/
#9340000000
0!
0'
b11 -
0/
b11 3
#9350000000
1!
1'
1/
12
#9360000000
0!
1$
0'
1*
b100 -
0/
b100 3
#9370000000
1!
1'
1/
#9380000000
0!
0'
b101 -
0/
b101 3
#9390000000
1!
0$
1'
0*
1/
#9400000000
0!
0'
b110 -
0/
b110 3
#9410000000
1!
1'
1/
#9420000000
0!
0'
b111 -
0/
b111 3
#9430000000
1!
1'
1/
02
#9440000000
0!
0'
b0 -
0/
b0 3
#9450000000
1!
1'
1/
#9460000000
0!
0'
b1 -
0/
b1 3
#9470000000
1!
1'
1/
#9480000000
0!
0'
b10 -
0/
b10 3
#9490000000
1!
1'
1/
#9500000000
0!
0'
b11 -
0/
b11 3
#9510000000
1!
1'
1/
12
#9520000000
0!
0'
b100 -
0/
b100 3
#9530000000
1!
1'
1/
#9540000000
0!
0'
b101 -
0/
b101 3
#9550000000
1!
1'
1/
#9560000000
0!
0'
b110 -
0/
b110 3
#9570000000
1!
1'
1/
#9580000000
0!
0'
b111 -
0/
b111 3
#9590000000
1!
1'
1/
02
#9600000000
0!
0'
b0 -
0/
b0 3
#9610000000
1!
1'
1/
#9620000000
0!
0'
b1 -
0/
b1 3
#9630000000
1!
1'
1/
#9640000000
0!
0'
b10 -
0/
b10 3
#9650000000
1!
1'
1/
#9660000000
0!
0'
b11 -
0/
b11 3
#9670000000
1!
1'
1/
12
#9680000000
0!
0'
b100 -
0/
b100 3
#9690000000
1!
1'
1/
#9700000000
0!
0'
b101 -
0/
b101 3
#9710000000
1!
1'
1/
#9720000000
0!
1#
0'
1)
b110 -
0/
b110 3
#9730000000
1!
1'
1/
#9740000000
0!
0'
b111 -
0/
b111 3
#9750000000
1!
b0000110 &
1'
b0000110 ,
b0011 .
1/
02
b0000110 4
b0011 5
#9760000000
0!
0#
0'
0)
b0 -
0/
b0 3
#9770000000
1!
1'
1/
#9780000000
0!
0'
b1 -
0/
b1 3
#9790000000
1!
1'
1/
#9800000000
0!
0'
b10 -
0/
b10 3
#9810000000
1!
1'
1/
#9820000000
0!
0'
b11 -
0/
b11 3
#9830000000
1!
1'
1/
12
#9840000000
0!
0'
b100 -
0/
b100 3
#9850000000
1!
1'
1/
#9860000000
0!
0'
b101 -
0/
b101 3
#9870000000
1!
1'
1/
#9880000000
0!
0'
b110 -
0/
b110 3
#9890000000
1!
1'
1/
#9900000000
0!
0'
b111 -
0/
b111 3
#9910000000
1!
b0110001 &
1'
b0110001 ,
b1100 .
1/
02
b0110001 4
b1100 5
#9920000000
0!
0'
b0 -
0/
b0 3
#9930000000
1!
1'
1/
#9940000000
0!
0'
b1 -
0/
b1 3
#9950000000
1!
1'
1/
#9960000000
0!
0'
b10 -
0/
b10 3
#9970000000
1!
1'
1/
#9980000000
0!
0'
b11 -
0/
b11 3
#9990000000
1!
1'
1/
12
#10000000000
0!
0'
b100 -
0/
b100 3
