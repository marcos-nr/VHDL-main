$date
  Wed May 22 22:26:48 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module math_real $end
$upscope $end
$scope module tb_transmisor_uart $end
$var reg 1 ! clk $end
$var reg 1 " key $end
$var reg 1 # reset $end
$var reg 1 $ tx $end
$var reg 1 % done $end
$scope module uut $end
$var reg 1 & clk $end
$var reg 1 ' key $end
$var reg 1 ( reset $end
$var reg 1 ) tx $end
$var reg 1 * done $end
$var reg 1 + send $end
$var reg 1 , clk_tx $end
$var reg 1 - clk_11tx $end
$var reg 8 . cadena[7:0] $end
$scope module a $end
$var reg 1 / clk $end
$var reg 1 0 reset $end
$var reg 1 1 enable $end
$var reg 1 2 cout $end
$var integer 32 3 q $end
$upscope $end
$scope module b $end
$var reg 1 4 clk $end
$var reg 1 5 reset $end
$var reg 1 6 enable $end
$var reg 1 7 cout $end
$var integer 32 8 q $end
$upscope $end
$scope module c $end
$var reg 1 9 clk $end
$var reg 1 : reset $end
$var reg 1 ; enable $end
$var reg 1 < send $end
$var reg 8 = cadena[7:0] $end
$var reg 1 > tx $end
$var reg 1 ? done $end
$var reg 1 @ clkss $end
$var reg 1 A clkis $end
$var reg 1 B rst1s $end
$var reg 8 C ds[7:0] $end
$comment estado is not handled $end
$var integer 32 D cnt $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
U"
0#
1$
0%
0&
U'
0(
1)
0*
1+
U,
U-
bUUUUUUUU .
0/
00
11
U2
b0 3
04
05
16
U7
b0 8
U9
0:
1;
1<
bUUUUUUUU =
1>
0?
0@
0A
0B
bUUUUUUUU C
b1 D
#10000000
1!
1&
0,
0-
1/
02
b1 3
14
07
b1 8
09
#20000000
0!
0&
0/
04
#30000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#40000000
0!
0&
0/
04
#50000000
1!
1&
1/
b11 3
14
b11 8
#60000000
0!
1"
0&
1'
0/
04
#70000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#80000000
0!
0&
0/
04
#90000000
1!
1&
1/
b1 3
14
b101 8
#100000000
0!
0&
0/
04
#110000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#120000000
0!
0&
0/
04
#130000000
1!
1&
1/
b11 3
14
b111 8
#140000000
0!
0&
0/
04
#150000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#160000000
0!
0&
0/
04
#170000000
1!
1&
1/
b1 3
14
b1001 8
#180000000
0!
0&
0/
04
#190000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#200000000
0!
0&
0/
04
#210000000
1!
1&
1/
b11 3
14
b1011 8
#220000000
0!
0&
0/
04
#230000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#240000000
0!
0&
0/
04
#250000000
1!
1&
1/
b1 3
14
b1101 8
#260000000
0!
0&
0/
04
#270000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#280000000
0!
0&
0/
04
#290000000
1!
1&
1/
b11 3
14
b1111 8
#300000000
0!
0&
0/
04
#310000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#320000000
0!
0&
0/
04
#330000000
1!
1&
1/
b1 3
14
b10001 8
#340000000
0!
0&
0/
04
#350000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#360000000
0!
0&
0/
04
#370000000
1!
1&
1/
b11 3
14
b10011 8
#380000000
0!
0"
0&
0'
0/
04
#390000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#400000000
0!
0&
0/
04
#410000000
1!
1&
1/
b1 3
14
b10101 8
#420000000
0!
0&
0/
04
#430000000
1!
1&
1,
1-
1/
12
b10 3
14
17
b10110 8
19
#440000000
0!
0&
0/
04
#450000000
1!
1&
1/
b11 3
14
b10111 8
#460000000
0!
0&
0/
04
#470000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
#480000000
0!
0&
0/
04
#490000000
1!
1&
1/
b1 3
14
b11001 8
#500000000
0!
0&
0/
04
#510000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#520000000
0!
0&
0/
04
#530000000
1!
1&
1/
b11 3
14
b11011 8
#540000000
0!
0&
0/
04
#550000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#560000000
0!
0&
0/
04
#570000000
1!
1&
1/
b1 3
14
b11101 8
#580000000
0!
0&
0/
04
#590000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#600000000
0!
0&
0/
04
#610000000
1!
1&
1/
b11 3
14
b11111 8
#620000000
0!
0&
0/
04
#630000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#640000000
0!
0&
0/
04
#650000000
1!
1&
1/
b1 3
14
b100001 8
#660000000
0!
0&
0/
04
#670000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#680000000
0!
0&
0/
04
#690000000
1!
1&
1/
b11 3
14
b100011 8
#700000000
0!
0&
0/
04
#710000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#720000000
0!
0&
0/
04
#730000000
1!
1&
1/
b1 3
14
b100101 8
#740000000
0!
0&
0/
04
#750000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#760000000
0!
0&
0/
04
#770000000
1!
1&
1/
b11 3
14
b100111 8
#780000000
0!
0&
0/
04
#790000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#800000000
0!
0&
0/
04
#810000000
1!
1&
1/
b1 3
14
b101001 8
#820000000
0!
0&
0/
04
#830000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#840000000
0!
0&
0/
04
#850000000
1!
1&
1/
b11 3
14
b101011 8
#860000000
0!
0&
0/
04
#870000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#880000000
0!
0&
0/
04
#890000000
1!
1&
1/
b1 3
14
b1 8
#900000000
0!
0&
0/
04
#910000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#920000000
0!
0&
0/
04
#930000000
1!
1&
1/
b11 3
14
b11 8
#940000000
0!
0&
0/
04
#950000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#960000000
0!
0&
0/
04
#970000000
1!
1&
1/
b1 3
14
b101 8
#980000000
0!
0&
0/
04
#990000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#1000000000
0!
0&
0/
04
#1010000000
1!
1&
1/
b11 3
14
b111 8
#1020000000
0!
0&
0/
04
#1030000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#1040000000
0!
0&
0/
04
#1050000000
1!
1&
1/
b1 3
14
b1001 8
#1060000000
0!
0&
0/
04
#1070000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#1080000000
0!
0&
0/
04
#1090000000
1!
1&
1/
b11 3
14
b1011 8
#1100000000
0!
0&
0/
04
#1110000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#1120000000
0!
0&
0/
04
#1130000000
1!
1&
1/
b1 3
14
b1101 8
#1140000000
0!
0&
0/
04
#1150000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#1160000000
0!
0&
0/
04
#1170000000
1!
1&
1/
b11 3
14
b1111 8
#1180000000
0!
0&
0/
04
#1190000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#1200000000
0!
0&
0/
04
#1210000000
1!
1&
1/
b1 3
14
b10001 8
#1220000000
0!
0&
0/
04
#1230000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#1240000000
0!
0&
0/
04
#1250000000
1!
1&
1/
b11 3
14
b10011 8
#1260000000
0!
0&
0/
04
#1270000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#1280000000
0!
0&
0/
04
#1290000000
1!
1&
1/
b1 3
14
b10101 8
#1300000000
0!
0&
0/
04
#1310000000
1!
1&
1,
1-
1/
12
b10 3
14
17
b10110 8
19
#1320000000
0!
0&
0/
04
#1330000000
1!
1&
1/
b11 3
14
b10111 8
#1340000000
0!
0&
0/
04
#1350000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
#1360000000
0!
0&
0/
04
#1370000000
1!
1&
1/
b1 3
14
b11001 8
#1380000000
0!
0&
0/
04
#1390000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#1400000000
0!
0&
0/
04
#1410000000
1!
1&
1/
b11 3
14
b11011 8
#1420000000
0!
1"
0&
1'
0/
04
#1430000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#1440000000
0!
0&
0/
04
#1450000000
1!
1&
1/
b1 3
14
b11101 8
#1460000000
0!
0&
0/
04
#1470000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#1480000000
0!
0&
0/
04
#1490000000
1!
1&
1/
b11 3
14
b11111 8
#1500000000
0!
0&
0/
04
#1510000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#1520000000
0!
0&
0/
04
#1530000000
1!
1&
1/
b1 3
14
b100001 8
#1540000000
0!
0&
0/
04
#1550000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#1560000000
0!
0&
0/
04
#1570000000
1!
1&
1/
b11 3
14
b100011 8
#1580000000
0!
0&
0/
04
#1590000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#1600000000
0!
0&
0/
04
#1610000000
1!
1&
1/
b1 3
14
b100101 8
#1620000000
0!
0&
0/
04
#1630000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#1640000000
0!
0&
0/
04
#1650000000
1!
1&
1/
b11 3
14
b100111 8
#1660000000
0!
0&
0/
04
#1670000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#1680000000
0!
0&
0/
04
#1690000000
1!
1&
1/
b1 3
14
b101001 8
#1700000000
0!
0&
0/
04
#1710000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#1720000000
0!
0&
0/
04
#1730000000
1!
1&
1/
b11 3
14
b101011 8
#1740000000
0!
0"
0&
0'
0/
04
#1750000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#1760000000
0!
0&
0/
04
#1770000000
1!
1&
1/
b1 3
14
b1 8
#1780000000
0!
0&
0/
04
#1790000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#1800000000
0!
0&
0/
04
#1810000000
1!
1&
1/
b11 3
14
b11 8
#1820000000
0!
0&
0/
04
#1830000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#1840000000
0!
0&
0/
04
#1850000000
1!
1&
1/
b1 3
14
b101 8
#1860000000
0!
0&
0/
04
#1870000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#1880000000
0!
0&
0/
04
#1890000000
1!
1&
1/
b11 3
14
b111 8
#1900000000
0!
0&
0/
04
#1910000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#1920000000
0!
0&
0/
04
#1930000000
1!
1&
1/
b1 3
14
b1001 8
#1940000000
0!
0&
0/
04
#1950000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#1960000000
0!
0&
0/
04
#1970000000
1!
1&
1/
b11 3
14
b1011 8
#1980000000
0!
0&
0/
04
#1990000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#2000000000
0!
0&
0/
04
#2010000000
1!
1&
1/
b1 3
14
b1101 8
#2020000000
0!
0&
0/
04
#2030000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#2040000000
0!
0&
0/
04
#2050000000
1!
1&
1/
b11 3
14
b1111 8
#2060000000
0!
0&
0/
04
#2070000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#2080000000
0!
0&
0/
04
#2090000000
1!
1&
1/
b1 3
14
b10001 8
#2100000000
0!
0&
0/
04
#2110000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#2120000000
0!
0&
0/
04
#2130000000
1!
1&
1/
b11 3
14
b10011 8
#2140000000
0!
0&
0/
04
#2150000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#2160000000
0!
0&
0/
04
#2170000000
1!
1&
1/
b1 3
14
b10101 8
#2180000000
0!
0&
0/
04
#2190000000
1!
1&
1,
1-
1/
12
b10 3
14
17
b10110 8
19
#2200000000
0!
0&
0/
04
#2210000000
1!
1&
1/
b11 3
14
b10111 8
#2220000000
0!
0&
0/
04
#2230000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
#2240000000
0!
0&
0/
04
#2250000000
1!
1&
1/
b1 3
14
b11001 8
#2260000000
0!
0&
0/
04
#2270000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#2280000000
0!
0&
0/
04
#2290000000
1!
1&
1/
b11 3
14
b11011 8
#2300000000
0!
0&
0/
04
#2310000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#2320000000
0!
0&
0/
04
#2330000000
1!
1&
1/
b1 3
14
b11101 8
#2340000000
0!
0&
0/
04
#2350000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#2360000000
0!
0&
0/
04
#2370000000
1!
1&
1/
b11 3
14
b11111 8
#2380000000
0!
0&
0/
04
#2390000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#2400000000
0!
0&
0/
04
#2410000000
1!
1&
1/
b1 3
14
b100001 8
#2420000000
0!
0&
0/
04
#2430000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#2440000000
0!
0&
0/
04
#2450000000
1!
1&
1/
b11 3
14
b100011 8
#2460000000
0!
0&
0/
04
#2470000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#2480000000
0!
0&
0/
04
#2490000000
1!
1&
1/
b1 3
14
b100101 8
#2500000000
0!
0&
0/
04
#2510000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#2520000000
0!
0&
0/
04
#2530000000
1!
1&
1/
b11 3
14
b100111 8
#2540000000
0!
0&
0/
04
#2550000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#2560000000
0!
0&
0/
04
#2570000000
1!
1&
1/
b1 3
14
b101001 8
#2580000000
0!
0&
0/
04
#2590000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#2600000000
0!
0&
0/
04
#2610000000
1!
1&
1/
b11 3
14
b101011 8
#2620000000
0!
0&
0/
04
#2630000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#2640000000
0!
0&
0/
04
#2650000000
1!
1&
1/
b1 3
14
b1 8
#2660000000
0!
0&
0/
04
#2670000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#2680000000
0!
0&
0/
04
#2690000000
1!
1&
1/
b11 3
14
b11 8
#2700000000
0!
0&
0/
04
#2710000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#2720000000
0!
0&
0/
04
#2730000000
1!
1&
1/
b1 3
14
b101 8
#2740000000
0!
0&
0/
04
#2750000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#2760000000
0!
0&
0/
04
#2770000000
1!
1&
1/
b11 3
14
b111 8
#2780000000
0!
1"
0&
1'
0/
04
#2790000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#2800000000
0!
0&
0/
04
#2810000000
1!
1&
1/
b1 3
14
b1001 8
#2820000000
0!
0&
0/
04
#2830000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#2840000000
0!
0&
0/
04
#2850000000
1!
1&
1/
b11 3
14
b1011 8
#2860000000
0!
0&
0/
04
#2870000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#2880000000
0!
0&
0/
04
#2890000000
1!
1&
1/
b1 3
14
b1101 8
#2900000000
0!
0&
0/
04
#2910000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#2920000000
0!
0&
0/
04
#2930000000
1!
1&
1/
b11 3
14
b1111 8
#2940000000
0!
0&
0/
04
#2950000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#2960000000
0!
0&
0/
04
#2970000000
1!
1&
1/
b1 3
14
b10001 8
#2980000000
0!
0&
0/
04
#2990000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#3000000000
0!
0&
0/
04
#3010000000
1!
1&
1/
b11 3
14
b10011 8
#3020000000
0!
0&
0/
04
#3030000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#3040000000
0!
0&
0/
04
#3050000000
1!
1&
1/
b1 3
14
b10101 8
#3060000000
0!
0&
0/
04
#3070000000
1!
1&
1,
1-
b01110111 .
1/
12
b10 3
14
17
b10110 8
19
b01110111 =
#3080000000
0!
0&
0/
04
#3090000000
1!
1&
1/
b11 3
14
b10111 8
#3100000000
0!
0"
0&
0'
0/
04
#3110000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
b01110111 C
#3120000000
0!
0&
0/
04
#3130000000
1!
1&
1/
b1 3
14
b11001 8
#3140000000
0!
0&
0/
04
#3150000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#3160000000
0!
0&
0/
04
#3170000000
1!
1&
1/
b11 3
14
b11011 8
#3180000000
0!
0&
0/
04
#3190000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#3200000000
0!
0&
0/
04
#3210000000
1!
1&
1/
b1 3
14
b11101 8
#3220000000
0!
0&
0/
04
#3230000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#3240000000
0!
0&
0/
04
#3250000000
1!
1&
1/
b11 3
14
b11111 8
#3260000000
0!
0&
0/
04
#3270000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#3280000000
0!
0&
0/
04
#3290000000
1!
1&
1/
b1 3
14
b100001 8
#3300000000
0!
0&
0/
04
#3310000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#3320000000
0!
0&
0/
04
#3330000000
1!
1&
1/
b11 3
14
b100011 8
#3340000000
0!
0&
0/
04
#3350000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#3360000000
0!
0&
0/
04
#3370000000
1!
1&
1/
b1 3
14
b100101 8
#3380000000
0!
0&
0/
04
#3390000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#3400000000
0!
0&
0/
04
#3410000000
1!
1&
1/
b11 3
14
b100111 8
#3420000000
0!
0&
0/
04
#3430000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#3440000000
0!
0&
0/
04
#3450000000
1!
1&
1/
b1 3
14
b101001 8
#3460000000
0!
0&
0/
04
#3470000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#3480000000
0!
0&
0/
04
#3490000000
1!
1&
1/
b11 3
14
b101011 8
#3500000000
0!
0&
0/
04
#3510000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#3520000000
0!
0&
0/
04
#3530000000
1!
1&
1/
b1 3
14
b1 8
#3540000000
0!
0&
0/
04
#3550000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#3560000000
0!
0&
0/
04
#3570000000
1!
1&
1/
b11 3
14
b11 8
#3580000000
0!
0&
0/
04
#3590000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#3600000000
0!
0&
0/
04
#3610000000
1!
1&
1/
b1 3
14
b101 8
#3620000000
0!
0&
0/
04
#3630000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#3640000000
0!
0&
0/
04
#3650000000
1!
1&
1/
b11 3
14
b111 8
#3660000000
0!
0&
0/
04
#3670000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#3680000000
0!
0&
0/
04
#3690000000
1!
1&
1/
b1 3
14
b1001 8
#3700000000
0!
0&
0/
04
#3710000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#3720000000
0!
0&
0/
04
#3730000000
1!
1&
1/
b11 3
14
b1011 8
#3740000000
0!
0&
0/
04
#3750000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#3760000000
0!
0&
0/
04
#3770000000
1!
1&
1/
b1 3
14
b1101 8
#3780000000
0!
0&
0/
04
#3790000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#3800000000
0!
0&
0/
04
#3810000000
1!
1&
1/
b11 3
14
b1111 8
#3820000000
0!
0&
0/
04
#3830000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#3840000000
0!
0&
0/
04
#3850000000
1!
1&
1/
b1 3
14
b10001 8
#3860000000
0!
0&
0/
04
#3870000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#3880000000
0!
0&
0/
04
#3890000000
1!
1&
1/
b11 3
14
b10011 8
#3900000000
0!
0&
0/
04
#3910000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#3920000000
0!
0&
0/
04
#3930000000
1!
1&
1/
b1 3
14
b10101 8
#3940000000
0!
0&
0/
04
#3950000000
1!
1&
1,
1-
1/
12
b10 3
14
17
b10110 8
19
#3960000000
0!
0&
0/
04
#3970000000
1!
1&
1/
b11 3
14
b10111 8
#3980000000
0!
0&
0/
04
#3990000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
#4000000000
0!
0&
0/
04
#4010000000
1!
1&
1/
b1 3
14
b11001 8
#4020000000
0!
0&
0/
04
#4030000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#4040000000
0!
0&
0/
04
#4050000000
1!
1&
1/
b11 3
14
b11011 8
#4060000000
0!
0&
0/
04
#4070000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#4080000000
0!
0&
0/
04
#4090000000
1!
1&
1/
b1 3
14
b11101 8
#4100000000
0!
0&
0/
04
#4110000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#4120000000
0!
0&
0/
04
#4130000000
1!
1&
1/
b11 3
14
b11111 8
#4140000000
0!
1"
0&
1'
0/
04
#4150000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#4160000000
0!
0&
0/
04
#4170000000
1!
1&
1/
b1 3
14
b100001 8
#4180000000
0!
0&
0/
04
#4190000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#4200000000
0!
0&
0/
04
#4210000000
1!
1&
1/
b11 3
14
b100011 8
#4220000000
0!
0&
0/
04
#4230000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#4240000000
0!
0&
0/
04
#4250000000
1!
1&
1/
b1 3
14
b100101 8
#4260000000
0!
0&
0/
04
#4270000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#4280000000
0!
0&
0/
04
#4290000000
1!
1&
1/
b11 3
14
b100111 8
#4300000000
0!
0&
0/
04
#4310000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#4320000000
0!
0&
0/
04
#4330000000
1!
1&
1/
b1 3
14
b101001 8
#4340000000
0!
0&
0/
04
#4350000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#4360000000
0!
0&
0/
04
#4370000000
1!
1&
1/
b11 3
14
b101011 8
#4380000000
0!
0&
0/
04
#4390000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#4400000000
0!
0&
0/
04
#4410000000
1!
1&
1/
b1 3
14
b1 8
#4420000000
0!
0&
0/
04
#4430000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#4440000000
0!
0&
0/
04
#4450000000
1!
1&
1/
b11 3
14
b11 8
#4460000000
0!
0"
0&
0'
0/
04
#4470000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#4480000000
0!
0&
0/
04
#4490000000
1!
1&
1/
b1 3
14
b101 8
#4500000000
0!
0&
0/
04
#4510000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#4520000000
0!
0&
0/
04
#4530000000
1!
1&
1/
b11 3
14
b111 8
#4540000000
0!
0&
0/
04
#4550000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#4560000000
0!
0&
0/
04
#4570000000
1!
1&
1/
b1 3
14
b1001 8
#4580000000
0!
0&
0/
04
#4590000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#4600000000
0!
0&
0/
04
#4610000000
1!
1&
1/
b11 3
14
b1011 8
#4620000000
0!
0&
0/
04
#4630000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#4640000000
0!
0&
0/
04
#4650000000
1!
1&
1/
b1 3
14
b1101 8
#4660000000
0!
0&
0/
04
#4670000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#4680000000
0!
0&
0/
04
#4690000000
1!
1&
1/
b11 3
14
b1111 8
#4700000000
0!
0&
0/
04
#4710000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#4720000000
0!
0&
0/
04
#4730000000
1!
1&
1/
b1 3
14
b10001 8
#4740000000
0!
0&
0/
04
#4750000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#4760000000
0!
0&
0/
04
#4770000000
1!
1&
1/
b11 3
14
b10011 8
#4780000000
0!
0&
0/
04
#4790000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#4800000000
0!
0&
0/
04
#4810000000
1!
1&
1/
b1 3
14
b10101 8
#4820000000
0!
0&
0/
04
#4830000000
1!
1&
1,
1-
1/
12
b10 3
14
17
b10110 8
19
#4840000000
0!
0&
0/
04
#4850000000
1!
1&
1/
b11 3
14
b10111 8
#4860000000
0!
0&
0/
04
#4870000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
#4880000000
0!
0&
0/
04
#4890000000
1!
1&
1/
b1 3
14
b11001 8
#4900000000
0!
0&
0/
04
#4910000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#4920000000
0!
0&
0/
04
#4930000000
1!
1&
1/
b11 3
14
b11011 8
#4940000000
0!
0&
0/
04
#4950000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#4960000000
0!
0&
0/
04
#4970000000
1!
1&
1/
b1 3
14
b11101 8
#4980000000
0!
0&
0/
04
#4990000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#5000000000
0!
0&
0/
04
#5010000000
1!
1&
1/
b11 3
14
b11111 8
#5020000000
0!
0&
0/
04
#5030000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#5040000000
0!
0&
0/
04
#5050000000
1!
1&
1/
b1 3
14
b100001 8
#5060000000
0!
0&
0/
04
#5070000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#5080000000
0!
0&
0/
04
#5090000000
1!
1&
1/
b11 3
14
b100011 8
#5100000000
0!
0&
0/
04
#5110000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#5120000000
0!
0&
0/
04
#5130000000
1!
1&
1/
b1 3
14
b100101 8
#5140000000
0!
0&
0/
04
#5150000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#5160000000
0!
0&
0/
04
#5170000000
1!
1&
1/
b11 3
14
b100111 8
#5180000000
0!
0&
0/
04
#5190000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#5200000000
0!
0&
0/
04
#5210000000
1!
1&
1/
b1 3
14
b101001 8
#5220000000
0!
0&
0/
04
#5230000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#5240000000
0!
0&
0/
04
#5250000000
1!
1&
1/
b11 3
14
b101011 8
#5260000000
0!
0&
0/
04
#5270000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#5280000000
0!
0&
0/
04
#5290000000
1!
1&
1/
b1 3
14
b1 8
#5300000000
0!
0&
0/
04
#5310000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#5320000000
0!
0&
0/
04
#5330000000
1!
1&
1/
b11 3
14
b11 8
#5340000000
0!
0&
0/
04
#5350000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#5360000000
0!
0&
0/
04
#5370000000
1!
1&
1/
b1 3
14
b101 8
#5380000000
0!
0&
0/
04
#5390000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#5400000000
0!
0&
0/
04
#5410000000
1!
1&
1/
b11 3
14
b111 8
#5420000000
0!
0&
0/
04
#5430000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#5440000000
0!
0&
0/
04
#5450000000
1!
1&
1/
b1 3
14
b1001 8
#5460000000
0!
0&
0/
04
#5470000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#5480000000
0!
0&
0/
04
#5490000000
1!
1&
1/
b11 3
14
b1011 8
#5500000000
0!
1"
0&
1'
0/
04
#5510000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#5520000000
0!
0&
0/
04
#5530000000
1!
1&
1/
b1 3
14
b1101 8
#5540000000
0!
0&
0/
04
#5550000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#5560000000
0!
0&
0/
04
#5570000000
1!
1&
1/
b11 3
14
b1111 8
#5580000000
0!
0&
0/
04
#5590000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#5600000000
0!
0&
0/
04
#5610000000
1!
1&
1/
b1 3
14
b10001 8
#5620000000
0!
0&
0/
04
#5630000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#5640000000
0!
0&
0/
04
#5650000000
1!
1&
1/
b11 3
14
b10011 8
#5660000000
0!
0&
0/
04
#5670000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#5680000000
0!
0&
0/
04
#5690000000
1!
1&
1/
b1 3
14
b10101 8
#5700000000
0!
0&
0/
04
#5710000000
1!
1&
1,
1-
b01111000 .
1/
12
b10 3
14
17
b10110 8
19
b01111000 =
#5720000000
0!
0&
0/
04
#5730000000
1!
1&
1/
b11 3
14
b10111 8
#5740000000
0!
0&
0/
04
#5750000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
b01111000 C
#5760000000
0!
0&
0/
04
#5770000000
1!
1&
1/
b1 3
14
b11001 8
#5780000000
0!
0&
0/
04
#5790000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#5800000000
0!
0&
0/
04
#5810000000
1!
1&
1/
b11 3
14
b11011 8
#5820000000
0!
0"
0&
0'
0/
04
#5830000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#5840000000
0!
0&
0/
04
#5850000000
1!
1&
1/
b1 3
14
b11101 8
#5860000000
0!
0&
0/
04
#5870000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#5880000000
0!
0&
0/
04
#5890000000
1!
1&
1/
b11 3
14
b11111 8
#5900000000
0!
0&
0/
04
#5910000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#5920000000
0!
0&
0/
04
#5930000000
1!
1&
1/
b1 3
14
b100001 8
#5940000000
0!
0&
0/
04
#5950000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#5960000000
0!
0&
0/
04
#5970000000
1!
1&
1/
b11 3
14
b100011 8
#5980000000
0!
0&
0/
04
#5990000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#6000000000
0!
0&
0/
04
#6010000000
1!
1&
1/
b1 3
14
b100101 8
#6020000000
0!
0&
0/
04
#6030000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#6040000000
0!
0&
0/
04
#6050000000
1!
1&
1/
b11 3
14
b100111 8
#6060000000
0!
0&
0/
04
#6070000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#6080000000
0!
0&
0/
04
#6090000000
1!
1&
1/
b1 3
14
b101001 8
#6100000000
0!
0&
0/
04
#6110000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#6120000000
0!
0&
0/
04
#6130000000
1!
1&
1/
b11 3
14
b101011 8
#6140000000
0!
0&
0/
04
#6150000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#6160000000
0!
0&
0/
04
#6170000000
1!
1&
1/
b1 3
14
b1 8
#6180000000
0!
0&
0/
04
#6190000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#6200000000
0!
0&
0/
04
#6210000000
1!
1&
1/
b11 3
14
b11 8
#6220000000
0!
0&
0/
04
#6230000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#6240000000
0!
0&
0/
04
#6250000000
1!
1&
1/
b1 3
14
b101 8
#6260000000
0!
0&
0/
04
#6270000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#6280000000
0!
0&
0/
04
#6290000000
1!
1&
1/
b11 3
14
b111 8
#6300000000
0!
0&
0/
04
#6310000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#6320000000
0!
0&
0/
04
#6330000000
1!
1&
1/
b1 3
14
b1001 8
#6340000000
0!
0&
0/
04
#6350000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#6360000000
0!
0&
0/
04
#6370000000
1!
1&
1/
b11 3
14
b1011 8
#6380000000
0!
0&
0/
04
#6390000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#6400000000
0!
0&
0/
04
#6410000000
1!
1&
1/
b1 3
14
b1101 8
#6420000000
0!
0&
0/
04
#6430000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#6440000000
0!
0&
0/
04
#6450000000
1!
1&
1/
b11 3
14
b1111 8
#6460000000
0!
0&
0/
04
#6470000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#6480000000
0!
0&
0/
04
#6490000000
1!
1&
1/
b1 3
14
b10001 8
#6500000000
0!
0&
0/
04
#6510000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#6520000000
0!
0&
0/
04
#6530000000
1!
1&
1/
b11 3
14
b10011 8
#6540000000
0!
0&
0/
04
#6550000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#6560000000
0!
0&
0/
04
#6570000000
1!
1&
1/
b1 3
14
b10101 8
#6580000000
0!
0&
0/
04
#6590000000
1!
1&
1,
1-
1/
12
b10 3
14
17
b10110 8
19
#6600000000
0!
0&
0/
04
#6610000000
1!
1&
1/
b11 3
14
b10111 8
#6620000000
0!
0&
0/
04
#6630000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
#6640000000
0!
0&
0/
04
#6650000000
1!
1&
1/
b1 3
14
b11001 8
#6660000000
0!
0&
0/
04
#6670000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#6680000000
0!
0&
0/
04
#6690000000
1!
1&
1/
b11 3
14
b11011 8
#6700000000
0!
0&
0/
04
#6710000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#6720000000
0!
0&
0/
04
#6730000000
1!
1&
1/
b1 3
14
b11101 8
#6740000000
0!
0&
0/
04
#6750000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#6760000000
0!
0&
0/
04
#6770000000
1!
1&
1/
b11 3
14
b11111 8
#6780000000
0!
0&
0/
04
#6790000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#6800000000
0!
0&
0/
04
#6810000000
1!
1&
1/
b1 3
14
b100001 8
#6820000000
0!
0&
0/
04
#6830000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#6840000000
0!
0&
0/
04
#6850000000
1!
1&
1/
b11 3
14
b100011 8
#6860000000
0!
1"
0&
1'
0/
04
#6870000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#6880000000
0!
0&
0/
04
#6890000000
1!
1&
1/
b1 3
14
b100101 8
#6900000000
0!
0&
0/
04
#6910000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#6920000000
0!
0&
0/
04
#6930000000
1!
1&
1/
b11 3
14
b100111 8
#6940000000
0!
0&
0/
04
#6950000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#6960000000
0!
0&
0/
04
#6970000000
1!
1&
1/
b1 3
14
b101001 8
#6980000000
0!
0&
0/
04
#6990000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#7000000000
0!
0&
0/
04
#7010000000
1!
1&
1/
b11 3
14
b101011 8
#7020000000
0!
0&
0/
04
#7030000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#7040000000
0!
0&
0/
04
#7050000000
1!
1&
1/
b1 3
14
b1 8
#7060000000
0!
0&
0/
04
#7070000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#7080000000
0!
0&
0/
04
#7090000000
1!
1&
1/
b11 3
14
b11 8
#7100000000
0!
0&
0/
04
#7110000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#7120000000
0!
0&
0/
04
#7130000000
1!
1&
1/
b1 3
14
b101 8
#7140000000
0!
0&
0/
04
#7150000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#7160000000
0!
0&
0/
04
#7170000000
1!
1&
1/
b11 3
14
b111 8
#7180000000
0!
0"
0&
0'
0/
04
#7190000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#7200000000
0!
0&
0/
04
#7210000000
1!
1&
1/
b1 3
14
b1001 8
#7220000000
0!
0&
0/
04
#7230000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#7240000000
0!
0&
0/
04
#7250000000
1!
1&
1/
b11 3
14
b1011 8
#7260000000
0!
0&
0/
04
#7270000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#7280000000
0!
0&
0/
04
#7290000000
1!
1&
1/
b1 3
14
b1101 8
#7300000000
0!
0&
0/
04
#7310000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#7320000000
0!
0&
0/
04
#7330000000
1!
1&
1/
b11 3
14
b1111 8
#7340000000
0!
0&
0/
04
#7350000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#7360000000
0!
0&
0/
04
#7370000000
1!
1&
1/
b1 3
14
b10001 8
#7380000000
0!
0&
0/
04
#7390000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#7400000000
0!
0&
0/
04
#7410000000
1!
1&
1/
b11 3
14
b10011 8
#7420000000
0!
0&
0/
04
#7430000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#7440000000
0!
0&
0/
04
#7450000000
1!
1&
1/
b1 3
14
b10101 8
#7460000000
0!
0&
0/
04
#7470000000
1!
1&
1,
1-
1/
12
b10 3
14
17
b10110 8
19
#7480000000
0!
0&
0/
04
#7490000000
1!
1&
1/
b11 3
14
b10111 8
#7500000000
0!
0&
0/
04
#7510000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
#7520000000
0!
0&
0/
04
#7530000000
1!
1&
1/
b1 3
14
b11001 8
#7540000000
0!
0&
0/
04
#7550000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#7560000000
0!
0&
0/
04
#7570000000
1!
1&
1/
b11 3
14
b11011 8
#7580000000
0!
0&
0/
04
#7590000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#7600000000
0!
0&
0/
04
#7610000000
1!
1&
1/
b1 3
14
b11101 8
#7620000000
0!
0&
0/
04
#7630000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#7640000000
0!
0&
0/
04
#7650000000
1!
1&
1/
b11 3
14
b11111 8
#7660000000
0!
0&
0/
04
#7670000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#7680000000
0!
0&
0/
04
#7690000000
1!
1&
1/
b1 3
14
b100001 8
#7700000000
0!
0&
0/
04
#7710000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#7720000000
0!
0&
0/
04
#7730000000
1!
1&
1/
b11 3
14
b100011 8
#7740000000
0!
0&
0/
04
#7750000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#7760000000
0!
0&
0/
04
#7770000000
1!
1&
1/
b1 3
14
b100101 8
#7780000000
0!
0&
0/
04
#7790000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#7800000000
0!
0&
0/
04
#7810000000
1!
1&
1/
b11 3
14
b100111 8
#7820000000
0!
0&
0/
04
#7830000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#7840000000
0!
0&
0/
04
#7850000000
1!
1&
1/
b1 3
14
b101001 8
#7860000000
0!
0&
0/
04
#7870000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#7880000000
0!
0&
0/
04
#7890000000
1!
1&
1/
b11 3
14
b101011 8
#7900000000
0!
0&
0/
04
#7910000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#7920000000
0!
0&
0/
04
#7930000000
1!
1&
1/
b1 3
14
b1 8
#7940000000
0!
0&
0/
04
#7950000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#7960000000
0!
0&
0/
04
#7970000000
1!
1&
1/
b11 3
14
b11 8
#7980000000
0!
0&
0/
04
#7990000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#8000000000
0!
0&
0/
04
#8010000000
1!
1&
1/
b1 3
14
b101 8
#8020000000
0!
0&
0/
04
#8030000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#8040000000
0!
0&
0/
04
#8050000000
1!
1&
1/
b11 3
14
b111 8
#8060000000
0!
0&
0/
04
#8070000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#8080000000
0!
0&
0/
04
#8090000000
1!
1&
1/
b1 3
14
b1001 8
#8100000000
0!
0&
0/
04
#8110000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#8120000000
0!
0&
0/
04
#8130000000
1!
1&
1/
b11 3
14
b1011 8
#8140000000
0!
0&
0/
04
#8150000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#8160000000
0!
0&
0/
04
#8170000000
1!
1&
1/
b1 3
14
b1101 8
#8180000000
0!
0&
0/
04
#8190000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#8200000000
0!
0&
0/
04
#8210000000
1!
1&
1/
b11 3
14
b1111 8
#8220000000
0!
1"
0&
1'
0/
04
#8230000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#8240000000
0!
0&
0/
04
#8250000000
1!
1&
1/
b1 3
14
b10001 8
#8260000000
0!
0&
0/
04
#8270000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#8280000000
0!
0&
0/
04
#8290000000
1!
1&
1/
b11 3
14
b10011 8
#8300000000
0!
0&
0/
04
#8310000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#8320000000
0!
0&
0/
04
#8330000000
1!
1&
1/
b1 3
14
b10101 8
#8340000000
0!
0&
0/
04
#8350000000
1!
1&
1,
1-
b10000010 .
1/
12
b10 3
14
17
b10110 8
19
b10000010 =
#8360000000
0!
0&
0/
04
#8370000000
1!
1&
1/
b11 3
14
b10111 8
#8380000000
0!
0&
0/
04
#8390000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
b10000010 C
#8400000000
0!
0&
0/
04
#8410000000
1!
1&
1/
b1 3
14
b11001 8
#8420000000
0!
0&
0/
04
#8430000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#8440000000
0!
0&
0/
04
#8450000000
1!
1&
1/
b11 3
14
b11011 8
#8460000000
0!
0&
0/
04
#8470000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#8480000000
0!
0&
0/
04
#8490000000
1!
1&
1/
b1 3
14
b11101 8
#8500000000
0!
0&
0/
04
#8510000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#8520000000
0!
0&
0/
04
#8530000000
1!
1&
1/
b11 3
14
b11111 8
#8540000000
0!
0"
0&
0'
0/
04
#8550000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#8560000000
0!
0&
0/
04
#8570000000
1!
1&
1/
b1 3
14
b100001 8
#8580000000
0!
0&
0/
04
#8590000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#8600000000
0!
0&
0/
04
#8610000000
1!
1&
1/
b11 3
14
b100011 8
#8620000000
0!
0&
0/
04
#8630000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#8640000000
0!
0&
0/
04
#8650000000
1!
1&
1/
b1 3
14
b100101 8
#8660000000
0!
0&
0/
04
#8670000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#8680000000
0!
0&
0/
04
#8690000000
1!
1&
1/
b11 3
14
b100111 8
#8700000000
0!
0&
0/
04
#8710000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#8720000000
0!
0&
0/
04
#8730000000
1!
1&
1/
b1 3
14
b101001 8
#8740000000
0!
0&
0/
04
#8750000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#8760000000
0!
0&
0/
04
#8770000000
1!
1&
1/
b11 3
14
b101011 8
#8780000000
0!
0&
0/
04
#8790000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#8800000000
0!
0&
0/
04
#8810000000
1!
1&
1/
b1 3
14
b1 8
#8820000000
0!
0&
0/
04
#8830000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#8840000000
0!
0&
0/
04
#8850000000
1!
1&
1/
b11 3
14
b11 8
#8860000000
0!
0&
0/
04
#8870000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#8880000000
0!
0&
0/
04
#8890000000
1!
1&
1/
b1 3
14
b101 8
#8900000000
0!
0&
0/
04
#8910000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#8920000000
0!
0&
0/
04
#8930000000
1!
1&
1/
b11 3
14
b111 8
#8940000000
0!
0&
0/
04
#8950000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#8960000000
0!
0&
0/
04
#8970000000
1!
1&
1/
b1 3
14
b1001 8
#8980000000
0!
0&
0/
04
#8990000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#9000000000
0!
0&
0/
04
#9010000000
1!
1&
1/
b11 3
14
b1011 8
#9020000000
0!
0&
0/
04
#9030000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#9040000000
0!
0&
0/
04
#9050000000
1!
1&
1/
b1 3
14
b1101 8
#9060000000
0!
0&
0/
04
#9070000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#9080000000
0!
0&
0/
04
#9090000000
1!
1&
1/
b11 3
14
b1111 8
#9100000000
0!
0&
0/
04
#9110000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#9120000000
0!
0&
0/
04
#9130000000
1!
1&
1/
b1 3
14
b10001 8
#9140000000
0!
0&
0/
04
#9150000000
1!
1&
1,
1/
12
b10 3
14
b10010 8
19
#9160000000
0!
0&
0/
04
#9170000000
1!
1&
1/
b11 3
14
b10011 8
#9180000000
0!
0&
0/
04
#9190000000
1!
1&
0,
1/
02
b0 3
14
b10100 8
09
#9200000000
0!
0&
0/
04
#9210000000
1!
1&
1/
b1 3
14
b10101 8
#9220000000
0!
0&
0/
04
#9230000000
1!
1&
1,
1-
1/
12
b10 3
14
17
b10110 8
19
#9240000000
0!
0&
0/
04
#9250000000
1!
1&
1/
b11 3
14
b10111 8
#9260000000
0!
0&
0/
04
#9270000000
1!
1&
0,
1/
02
b0 3
14
b11000 8
09
#9280000000
0!
0&
0/
04
#9290000000
1!
1&
1/
b1 3
14
b11001 8
#9300000000
0!
0&
0/
04
#9310000000
1!
1&
1,
1/
12
b10 3
14
b11010 8
19
#9320000000
0!
0&
0/
04
#9330000000
1!
1&
1/
b11 3
14
b11011 8
#9340000000
0!
0&
0/
04
#9350000000
1!
1&
0,
1/
02
b0 3
14
b11100 8
09
#9360000000
0!
0&
0/
04
#9370000000
1!
1&
1/
b1 3
14
b11101 8
#9380000000
0!
0&
0/
04
#9390000000
1!
1&
1,
1/
12
b10 3
14
b11110 8
19
#9400000000
0!
0&
0/
04
#9410000000
1!
1&
1/
b11 3
14
b11111 8
#9420000000
0!
0&
0/
04
#9430000000
1!
1&
0,
1/
02
b0 3
14
b100000 8
09
#9440000000
0!
0&
0/
04
#9450000000
1!
1&
1/
b1 3
14
b100001 8
#9460000000
0!
0&
0/
04
#9470000000
1!
1&
1,
1/
12
b10 3
14
b100010 8
19
#9480000000
0!
0&
0/
04
#9490000000
1!
1&
1/
b11 3
14
b100011 8
#9500000000
0!
0&
0/
04
#9510000000
1!
1&
0,
1/
02
b0 3
14
b100100 8
09
#9520000000
0!
0&
0/
04
#9530000000
1!
1&
1/
b1 3
14
b100101 8
#9540000000
0!
0&
0/
04
#9550000000
1!
1&
1,
1/
12
b10 3
14
b100110 8
19
#9560000000
0!
0&
0/
04
#9570000000
1!
1&
1/
b11 3
14
b100111 8
#9580000000
0!
1"
0&
1'
0/
04
#9590000000
1!
1&
0,
1/
02
b0 3
14
b101000 8
09
#9600000000
0!
0&
0/
04
#9610000000
1!
1&
1/
b1 3
14
b101001 8
#9620000000
0!
0&
0/
04
#9630000000
1!
1&
1,
1/
12
b10 3
14
b101010 8
19
#9640000000
0!
0&
0/
04
#9650000000
1!
1&
1/
b11 3
14
b101011 8
#9660000000
0!
0&
0/
04
#9670000000
1!
1&
0,
0-
1/
02
b0 3
14
07
b0 8
09
#9680000000
0!
0&
0/
04
#9690000000
1!
1&
1/
b1 3
14
b1 8
#9700000000
0!
0&
0/
04
#9710000000
1!
1&
1,
1/
12
b10 3
14
b10 8
19
#9720000000
0!
0&
0/
04
#9730000000
1!
1&
1/
b11 3
14
b11 8
#9740000000
0!
0&
0/
04
#9750000000
1!
1&
0,
1/
02
b0 3
14
b100 8
09
#9760000000
0!
0&
0/
04
#9770000000
1!
1&
1/
b1 3
14
b101 8
#9780000000
0!
0&
0/
04
#9790000000
1!
1&
1,
1/
12
b10 3
14
b110 8
19
#9800000000
0!
0&
0/
04
#9810000000
1!
1&
1/
b11 3
14
b111 8
#9820000000
0!
0&
0/
04
#9830000000
1!
1&
0,
1/
02
b0 3
14
b1000 8
09
#9840000000
0!
0&
0/
04
#9850000000
1!
1&
1/
b1 3
14
b1001 8
#9860000000
0!
0&
0/
04
#9870000000
1!
1&
1,
1/
12
b10 3
14
b1010 8
19
#9880000000
0!
0&
0/
04
#9890000000
1!
1&
1/
b11 3
14
b1011 8
#9900000000
0!
0"
0&
0'
0/
04
#9910000000
1!
1&
0,
1/
02
b0 3
14
b1100 8
09
#9920000000
0!
0&
0/
04
#9930000000
1!
1&
1/
b1 3
14
b1101 8
#9940000000
0!
0&
0/
04
#9950000000
1!
1&
1,
1/
12
b10 3
14
b1110 8
19
#9960000000
0!
0&
0/
04
#9970000000
1!
1&
1/
b11 3
14
b1111 8
#9980000000
0!
0&
0/
04
#9990000000
1!
1&
0,
1/
02
b0 3
14
b10000 8
09
#10000000000
0!
0&
0/
04
