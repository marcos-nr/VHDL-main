$date
  Tue Apr 30 15:28:09 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp2_3 $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 4 # enable_disp[3:0] $end
$var reg 7 $ segmentos[6:0] $end
$scope module uut $end
$var reg 1 % clk $end
$var reg 1 & reset $end
$var reg 4 ' enable_disp[3:0] $end
$var reg 7 ( segmentos[6:0] $end
$comment state is not handled $end
$var reg 4 ) bcd[3:0] $end
$var integer 32 * cuenta $end
$var reg 1 + debounced_reset $end
$var reg 1 , enable_conta $end
$scope module a $end
$var reg 1 - clk $end
$var reg 1 . key $end
$var reg 1 / debounced_key $end
$var reg 1 0 key_stable $end
$var reg 1 1 last_key $end
$upscope $end
$scope module b $end
$var reg 1 2 clk $end
$var reg 1 3 reset $end
$var reg 1 4 enable $end
$var reg 1 5 cout $end
$var integer 32 6 q $end
$upscope $end
$scope module d $end
$var reg 7 7 segmentos[6:0] $end
$var reg 4 8 bcd[3:0] $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
U"
b1000 #
b0110000 $
0%
U&
b1000 '
b0110000 (
b0001 )
b0 *
U+
1,
0-
U.
U/
U0
U1
02
U3
14
U5
b0 6
b0110000 7
b0001 8
#10000000
1!
1%
1-
12
05
#20000000
0!
0%
b1 *
0-
02
b1 6
#30000000
1!
1%
1-
12
#40000000
0!
0%
b10 *
0-
02
b10 6
#50000000
1!
1%
1-
12
#60000000
0!
0%
b11 *
0-
02
b11 6
#70000000
1!
1%
1-
12
15
#80000000
0!
0%
b100 *
0-
02
b100 6
#90000000
1!
1%
1-
12
#100000000
0!
0%
b101 *
0-
02
b101 6
#110000000
1!
1%
1-
12
#120000000
0!
0%
b110 *
0-
02
b110 6
#130000000
1!
1%
1-
12
#140000000
0!
0%
b111 *
0-
02
b111 6
#150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#160000000
0!
0"
0%
0&
b0 *
0-
0.
02
b0 6
#170000000
1!
1%
0+
1-
0/
00
01
12
03
#180000000
0!
0%
b1 *
0-
02
b1 6
#190000000
1!
1%
1-
12
#200000000
0!
0%
b10 *
0-
02
b10 6
#210000000
1!
1%
1-
12
#220000000
0!
0%
b11 *
0-
02
b11 6
#230000000
1!
1%
1-
12
15
#240000000
0!
0%
b100 *
0-
02
b100 6
#250000000
1!
1%
1-
12
#260000000
0!
0%
b101 *
0-
02
b101 6
#270000000
1!
1%
1-
12
#280000000
0!
0%
b110 *
0-
02
b110 6
#290000000
1!
1%
1-
12
#300000000
0!
0%
b111 *
0-
02
b111 6
#310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#320000000
0!
0%
b0 *
0-
02
b0 6
#330000000
1!
1%
1-
12
#340000000
0!
0%
b1 *
0-
02
b1 6
#350000000
1!
1%
1-
12
#360000000
0!
0%
b10 *
0-
02
b10 6
#370000000
1!
1%
1-
12
#380000000
0!
0%
b11 *
0-
02
b11 6
#390000000
1!
1%
1-
12
15
#400000000
0!
0%
b100 *
0-
02
b100 6
#410000000
1!
1%
1-
12
#420000000
0!
0%
b101 *
0-
02
b101 6
#430000000
1!
1%
1-
12
#440000000
0!
0%
b110 *
0-
02
b110 6
#450000000
1!
1%
1-
12
#460000000
0!
0%
b111 *
0-
02
b111 6
#470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#480000000
0!
0%
b0 *
0-
02
b0 6
#490000000
1!
1%
1-
12
#500000000
0!
0%
b1 *
0-
02
b1 6
#510000000
1!
1%
1-
12
#520000000
0!
0%
b10 *
0-
02
b10 6
#530000000
1!
1%
1-
12
#540000000
0!
0%
b11 *
0-
02
b11 6
#550000000
1!
1%
1-
12
15
#560000000
0!
0%
b100 *
0-
02
b100 6
#570000000
1!
1%
1-
12
#580000000
0!
0%
b101 *
0-
02
b101 6
#590000000
1!
1%
1-
12
#600000000
0!
0%
b110 *
0-
02
b110 6
#610000000
1!
1%
1-
12
#620000000
0!
0%
b111 *
0-
02
b111 6
#630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#640000000
0!
0%
b0 *
0-
02
b0 6
#650000000
1!
1%
1-
12
#660000000
0!
0%
b1 *
0-
02
b1 6
#670000000
1!
1%
1-
12
#680000000
0!
0%
b10 *
0-
02
b10 6
#690000000
1!
1%
1-
12
#700000000
0!
0%
b11 *
0-
02
b11 6
#710000000
1!
1%
1-
12
15
#720000000
0!
0%
b100 *
0-
02
b100 6
#730000000
1!
1%
1-
12
#740000000
0!
0%
b101 *
0-
02
b101 6
#750000000
1!
1%
1-
12
#760000000
0!
0%
b110 *
0-
02
b110 6
#770000000
1!
1%
1-
12
#780000000
0!
0%
b111 *
0-
02
b111 6
#790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#800000000
0!
0%
b0 *
0-
02
b0 6
#810000000
1!
1%
1-
12
#820000000
0!
0%
b1 *
0-
02
b1 6
#830000000
1!
1%
1-
12
#840000000
0!
0%
b10 *
0-
02
b10 6
#850000000
1!
1%
1-
12
#860000000
0!
0%
b11 *
0-
02
b11 6
#870000000
1!
1%
1-
12
15
#880000000
0!
0%
b100 *
0-
02
b100 6
#890000000
1!
1%
1-
12
#900000000
0!
0%
b101 *
0-
02
b101 6
#910000000
1!
1%
1-
12
#920000000
0!
0%
b110 *
0-
02
b110 6
#930000000
1!
1%
1-
12
#940000000
0!
0%
b111 *
0-
02
b111 6
#950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#960000000
0!
0%
b0 *
0-
02
b0 6
#970000000
1!
1%
1-
12
#980000000
0!
0%
b1 *
0-
02
b1 6
#990000000
1!
1%
1-
12
#1000000000
0!
0%
b10 *
0-
02
b10 6
#1010000000
1!
1%
1-
12
#1020000000
0!
0%
b11 *
0-
02
b11 6
#1030000000
1!
1%
1-
12
15
#1040000000
0!
0%
b100 *
0-
02
b100 6
#1050000000
1!
1%
1-
12
#1060000000
0!
0%
b101 *
0-
02
b101 6
#1070000000
1!
1%
1-
12
#1080000000
0!
0%
b110 *
0-
02
b110 6
#1090000000
1!
1%
1-
12
#1100000000
0!
0%
b111 *
0-
02
b111 6
#1110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#1120000000
0!
0%
b0 *
0-
02
b0 6
#1130000000
1!
1%
1-
12
#1140000000
0!
0%
b1 *
0-
02
b1 6
#1150000000
1!
1%
1-
12
#1160000000
0!
0%
b10 *
0-
02
b10 6
#1170000000
1!
1%
1-
12
#1180000000
0!
0%
b11 *
0-
02
b11 6
#1190000000
1!
1%
1-
12
15
#1200000000
0!
0%
b100 *
0-
02
b100 6
#1210000000
1!
1%
1-
12
#1220000000
0!
0%
b101 *
0-
02
b101 6
#1230000000
1!
1%
1-
12
#1240000000
0!
0%
b110 *
0-
02
b110 6
#1250000000
1!
1%
1-
12
#1260000000
0!
0%
b111 *
0-
02
b111 6
#1270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#1280000000
0!
0%
b0 *
0-
02
b0 6
#1290000000
1!
1%
1-
12
#1300000000
0!
0%
b1 *
0-
02
b1 6
#1310000000
1!
1%
1-
12
#1320000000
0!
0%
b10 *
0-
02
b10 6
#1330000000
1!
1%
1-
12
#1340000000
0!
0%
b11 *
0-
02
b11 6
#1350000000
1!
1%
1-
12
15
#1360000000
0!
0%
b100 *
0-
02
b100 6
#1370000000
1!
1%
1-
12
#1380000000
0!
0%
b101 *
0-
02
b101 6
#1390000000
1!
1%
1-
12
#1400000000
0!
0%
b110 *
0-
02
b110 6
#1410000000
1!
1%
1-
12
#1420000000
0!
0%
b111 *
0-
02
b111 6
#1430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#1440000000
0!
0%
b0 *
0-
02
b0 6
#1450000000
1!
1%
1-
12
#1460000000
0!
0%
b1 *
0-
02
b1 6
#1470000000
1!
1%
1-
12
#1480000000
0!
0%
b10 *
0-
02
b10 6
#1490000000
1!
1%
1-
12
#1500000000
0!
0%
b11 *
0-
02
b11 6
#1510000000
1!
1%
1-
12
15
#1520000000
0!
0%
b100 *
0-
02
b100 6
#1530000000
1!
1%
1-
12
#1540000000
0!
0%
b101 *
0-
02
b101 6
#1550000000
1!
1%
1-
12
#1560000000
0!
0%
b110 *
0-
02
b110 6
#1570000000
1!
1%
1-
12
#1580000000
0!
0%
b111 *
0-
02
b111 6
#1590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#1600000000
0!
0%
b0 *
0-
02
b0 6
#1610000000
1!
1%
1-
12
#1620000000
0!
0%
b1 *
0-
02
b1 6
#1630000000
1!
1%
1-
12
#1640000000
0!
0%
b10 *
0-
02
b10 6
#1650000000
1!
1%
1-
12
#1660000000
0!
0%
b11 *
0-
02
b11 6
#1670000000
1!
1%
1-
12
15
#1680000000
0!
0%
b100 *
0-
02
b100 6
#1690000000
1!
1%
1-
12
#1700000000
0!
0%
b101 *
0-
02
b101 6
#1710000000
1!
1%
1-
12
#1720000000
0!
0%
b110 *
0-
02
b110 6
#1730000000
1!
1%
1-
12
#1740000000
0!
0%
b111 *
0-
02
b111 6
#1750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#1760000000
0!
0%
b0 *
0-
02
b0 6
#1770000000
1!
1%
1-
12
#1780000000
0!
0%
b1 *
0-
02
b1 6
#1790000000
1!
1%
1-
12
#1800000000
0!
0%
b10 *
0-
02
b10 6
#1810000000
1!
1%
1-
12
#1820000000
0!
0%
b11 *
0-
02
b11 6
#1830000000
1!
1%
1-
12
15
#1840000000
0!
0%
b100 *
0-
02
b100 6
#1850000000
1!
1%
1-
12
#1860000000
0!
0%
b101 *
0-
02
b101 6
#1870000000
1!
1%
1-
12
#1880000000
0!
0%
b110 *
0-
02
b110 6
#1890000000
1!
1%
1-
12
#1900000000
0!
0%
b111 *
0-
02
b111 6
#1910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#1920000000
0!
0%
b0 *
0-
02
b0 6
#1930000000
1!
1%
1-
12
#1940000000
0!
0%
b1 *
0-
02
b1 6
#1950000000
1!
1%
1-
12
#1960000000
0!
0%
b10 *
0-
02
b10 6
#1970000000
1!
1%
1-
12
#1980000000
0!
0%
b11 *
0-
02
b11 6
#1990000000
1!
1%
1-
12
15
#2000000000
0!
0%
b100 *
0-
02
b100 6
#2010000000
1!
1%
1-
12
#2020000000
0!
0%
b101 *
0-
02
b101 6
#2030000000
1!
1%
1-
12
#2040000000
0!
0%
b110 *
0-
02
b110 6
#2050000000
1!
1%
1-
12
#2060000000
0!
0%
b111 *
0-
02
b111 6
#2070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#2080000000
0!
0%
b0 *
0-
02
b0 6
#2090000000
1!
1%
1-
12
#2100000000
0!
0%
b1 *
0-
02
b1 6
#2110000000
1!
1%
1-
12
#2120000000
0!
0%
b10 *
0-
02
b10 6
#2130000000
1!
1%
1-
12
#2140000000
0!
0%
b11 *
0-
02
b11 6
#2150000000
1!
1%
1-
12
15
#2160000000
0!
0%
b100 *
0-
02
b100 6
#2170000000
1!
1%
1-
12
#2180000000
0!
0%
b101 *
0-
02
b101 6
#2190000000
1!
1%
1-
12
#2200000000
0!
0%
b110 *
0-
02
b110 6
#2210000000
1!
1%
1-
12
#2220000000
0!
0%
b111 *
0-
02
b111 6
#2230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#2240000000
0!
0%
b0 *
0-
02
b0 6
#2250000000
1!
1%
1-
12
#2260000000
0!
0%
b1 *
0-
02
b1 6
#2270000000
1!
1%
1-
12
#2280000000
0!
0%
b10 *
0-
02
b10 6
#2290000000
1!
1%
1-
12
#2300000000
0!
0%
b11 *
0-
02
b11 6
#2310000000
1!
1%
1-
12
15
#2320000000
0!
0%
b100 *
0-
02
b100 6
#2330000000
1!
1%
1-
12
#2340000000
0!
0%
b101 *
0-
02
b101 6
#2350000000
1!
1%
1-
12
#2360000000
0!
0%
b110 *
0-
02
b110 6
#2370000000
1!
1%
1-
12
#2380000000
0!
0%
b111 *
0-
02
b111 6
#2390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#2400000000
0!
0%
b0 *
0-
02
b0 6
#2410000000
1!
1%
1-
12
#2420000000
0!
0%
b1 *
0-
02
b1 6
#2430000000
1!
1%
1-
12
#2440000000
0!
0%
b10 *
0-
02
b10 6
#2450000000
1!
1%
1-
12
#2460000000
0!
0%
b11 *
0-
02
b11 6
#2470000000
1!
1%
1-
12
15
#2480000000
0!
0%
b100 *
0-
02
b100 6
#2490000000
1!
1%
1-
12
#2500000000
0!
0%
b101 *
0-
02
b101 6
#2510000000
1!
1%
1-
12
#2520000000
0!
0%
b110 *
0-
02
b110 6
#2530000000
1!
1%
1-
12
#2540000000
0!
0%
b111 *
0-
02
b111 6
#2550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#2560000000
0!
0%
b0 *
0-
02
b0 6
#2570000000
1!
1%
1-
12
#2580000000
0!
0%
b1 *
0-
02
b1 6
#2590000000
1!
1%
1-
12
#2600000000
0!
0%
b10 *
0-
02
b10 6
#2610000000
1!
1%
1-
12
#2620000000
0!
0%
b11 *
0-
02
b11 6
#2630000000
1!
1%
1-
12
15
#2640000000
0!
0%
b100 *
0-
02
b100 6
#2650000000
1!
1%
1-
12
#2660000000
0!
0%
b101 *
0-
02
b101 6
#2670000000
1!
1%
1-
12
#2680000000
0!
0%
b110 *
0-
02
b110 6
#2690000000
1!
1%
1-
12
#2700000000
0!
0%
b111 *
0-
02
b111 6
#2710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#2720000000
0!
0%
b0 *
0-
02
b0 6
#2730000000
1!
1%
1-
12
#2740000000
0!
0%
b1 *
0-
02
b1 6
#2750000000
1!
1%
1-
12
#2760000000
0!
0%
b10 *
0-
02
b10 6
#2770000000
1!
1%
1-
12
#2780000000
0!
0%
b11 *
0-
02
b11 6
#2790000000
1!
1%
1-
12
15
#2800000000
0!
0%
b100 *
0-
02
b100 6
#2810000000
1!
1%
1-
12
#2820000000
0!
0%
b101 *
0-
02
b101 6
#2830000000
1!
1%
1-
12
#2840000000
0!
0%
b110 *
0-
02
b110 6
#2850000000
1!
1%
1-
12
#2860000000
0!
0%
b111 *
0-
02
b111 6
#2870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#2880000000
0!
0%
b0 *
0-
02
b0 6
#2890000000
1!
1%
1-
12
#2900000000
0!
0%
b1 *
0-
02
b1 6
#2910000000
1!
1%
1-
12
#2920000000
0!
0%
b10 *
0-
02
b10 6
#2930000000
1!
1%
1-
12
#2940000000
0!
0%
b11 *
0-
02
b11 6
#2950000000
1!
1%
1-
12
15
#2960000000
0!
0%
b100 *
0-
02
b100 6
#2970000000
1!
1%
1-
12
#2980000000
0!
0%
b101 *
0-
02
b101 6
#2990000000
1!
1%
1-
12
#3000000000
0!
0%
b110 *
0-
02
b110 6
#3010000000
1!
1%
1-
12
#3020000000
0!
0%
b111 *
0-
02
b111 6
#3030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#3040000000
0!
0%
b0 *
0-
02
b0 6
#3050000000
1!
1%
1-
12
#3060000000
0!
0%
b1 *
0-
02
b1 6
#3070000000
1!
1%
1-
12
#3080000000
0!
0%
b10 *
0-
02
b10 6
#3090000000
1!
1%
1-
12
#3100000000
0!
0%
b11 *
0-
02
b11 6
#3110000000
1!
1%
1-
12
15
#3120000000
0!
0%
b100 *
0-
02
b100 6
#3130000000
1!
1%
1-
12
#3140000000
0!
0%
b101 *
0-
02
b101 6
#3150000000
1!
1%
1-
12
#3160000000
0!
0%
b110 *
0-
02
b110 6
#3170000000
1!
1%
1-
12
#3180000000
0!
0%
b111 *
0-
02
b111 6
#3190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#3200000000
0!
0%
b0 *
0-
02
b0 6
#3210000000
1!
1%
1-
12
#3220000000
0!
0%
b1 *
0-
02
b1 6
#3230000000
1!
1%
1-
12
#3240000000
0!
0%
b10 *
0-
02
b10 6
#3250000000
1!
1%
1-
12
#3260000000
0!
0%
b11 *
0-
02
b11 6
#3270000000
1!
1%
1-
12
15
#3280000000
0!
0%
b100 *
0-
02
b100 6
#3290000000
1!
1%
1-
12
#3300000000
0!
0%
b101 *
0-
02
b101 6
#3310000000
1!
1%
1-
12
#3320000000
0!
0%
b110 *
0-
02
b110 6
#3330000000
1!
1%
1-
12
#3340000000
0!
0%
b111 *
0-
02
b111 6
#3350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#3360000000
0!
0%
b0 *
0-
02
b0 6
#3370000000
1!
1%
1-
12
#3380000000
0!
0%
b1 *
0-
02
b1 6
#3390000000
1!
1%
1-
12
#3400000000
0!
0%
b10 *
0-
02
b10 6
#3410000000
1!
1%
1-
12
#3420000000
0!
0%
b11 *
0-
02
b11 6
#3430000000
1!
1%
1-
12
15
#3440000000
0!
0%
b100 *
0-
02
b100 6
#3450000000
1!
1%
1-
12
#3460000000
0!
0%
b101 *
0-
02
b101 6
#3470000000
1!
1%
1-
12
#3480000000
0!
0%
b110 *
0-
02
b110 6
#3490000000
1!
1%
1-
12
#3500000000
0!
0%
b111 *
0-
02
b111 6
#3510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#3520000000
0!
0%
b0 *
0-
02
b0 6
#3530000000
1!
1%
1-
12
#3540000000
0!
0%
b1 *
0-
02
b1 6
#3550000000
1!
1%
1-
12
#3560000000
0!
0%
b10 *
0-
02
b10 6
#3570000000
1!
1%
1-
12
#3580000000
0!
0%
b11 *
0-
02
b11 6
#3590000000
1!
1%
1-
12
15
#3600000000
0!
0%
b100 *
0-
02
b100 6
#3610000000
1!
1%
1-
12
#3620000000
0!
0%
b101 *
0-
02
b101 6
#3630000000
1!
1%
1-
12
#3640000000
0!
0%
b110 *
0-
02
b110 6
#3650000000
1!
1%
1-
12
#3660000000
0!
0%
b111 *
0-
02
b111 6
#3670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#3680000000
0!
0%
b0 *
0-
02
b0 6
#3690000000
1!
1%
1-
12
#3700000000
0!
0%
b1 *
0-
02
b1 6
#3710000000
1!
1%
1-
12
#3720000000
0!
0%
b10 *
0-
02
b10 6
#3730000000
1!
1%
1-
12
#3740000000
0!
0%
b11 *
0-
02
b11 6
#3750000000
1!
1%
1-
12
15
#3760000000
0!
0%
b100 *
0-
02
b100 6
#3770000000
1!
1%
1-
12
#3780000000
0!
0%
b101 *
0-
02
b101 6
#3790000000
1!
1%
1-
12
#3800000000
0!
0%
b110 *
0-
02
b110 6
#3810000000
1!
1%
1-
12
#3820000000
0!
0%
b111 *
0-
02
b111 6
#3830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#3840000000
0!
0%
b0 *
0-
02
b0 6
#3850000000
1!
1%
1-
12
#3860000000
0!
0%
b1 *
0-
02
b1 6
#3870000000
1!
1%
1-
12
#3880000000
0!
0%
b10 *
0-
02
b10 6
#3890000000
1!
1%
1-
12
#3900000000
0!
0%
b11 *
0-
02
b11 6
#3910000000
1!
1%
1-
12
15
#3920000000
0!
0%
b100 *
0-
02
b100 6
#3930000000
1!
1%
1-
12
#3940000000
0!
0%
b101 *
0-
02
b101 6
#3950000000
1!
1%
1-
12
#3960000000
0!
0%
b110 *
0-
02
b110 6
#3970000000
1!
1%
1-
12
#3980000000
0!
0%
b111 *
0-
02
b111 6
#3990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#4000000000
0!
0%
b0 *
0-
02
b0 6
#4010000000
1!
1%
1-
12
#4020000000
0!
0%
b1 *
0-
02
b1 6
#4030000000
1!
1%
1-
12
#4040000000
0!
0%
b10 *
0-
02
b10 6
#4050000000
1!
1%
1-
12
#4060000000
0!
0%
b11 *
0-
02
b11 6
#4070000000
1!
1%
1-
12
15
#4080000000
0!
0%
b100 *
0-
02
b100 6
#4090000000
1!
1%
1-
12
#4100000000
0!
0%
b101 *
0-
02
b101 6
#4110000000
1!
1%
1-
12
#4120000000
0!
0%
b110 *
0-
02
b110 6
#4130000000
1!
1%
1-
12
#4140000000
0!
0%
b111 *
0-
02
b111 6
#4150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#4160000000
0!
0%
b0 *
0-
02
b0 6
#4170000000
1!
1%
1-
12
#4180000000
0!
0%
b1 *
0-
02
b1 6
#4190000000
1!
1%
1-
12
#4200000000
0!
0%
b10 *
0-
02
b10 6
#4210000000
1!
1%
1-
12
#4220000000
0!
0%
b11 *
0-
02
b11 6
#4230000000
1!
1%
1-
12
15
#4240000000
0!
0%
b100 *
0-
02
b100 6
#4250000000
1!
1%
1-
12
#4260000000
0!
0%
b101 *
0-
02
b101 6
#4270000000
1!
1%
1-
12
#4280000000
0!
0%
b110 *
0-
02
b110 6
#4290000000
1!
1%
1-
12
#4300000000
0!
0%
b111 *
0-
02
b111 6
#4310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#4320000000
0!
0%
b0 *
0-
02
b0 6
#4330000000
1!
1%
1-
12
#4340000000
0!
0%
b1 *
0-
02
b1 6
#4350000000
1!
1%
1-
12
#4360000000
0!
0%
b10 *
0-
02
b10 6
#4370000000
1!
1%
1-
12
#4380000000
0!
0%
b11 *
0-
02
b11 6
#4390000000
1!
1%
1-
12
15
#4400000000
0!
0%
b100 *
0-
02
b100 6
#4410000000
1!
1%
1-
12
#4420000000
0!
0%
b101 *
0-
02
b101 6
#4430000000
1!
1%
1-
12
#4440000000
0!
0%
b110 *
0-
02
b110 6
#4450000000
1!
1%
1-
12
#4460000000
0!
0%
b111 *
0-
02
b111 6
#4470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#4480000000
0!
0%
b0 *
0-
02
b0 6
#4490000000
1!
1%
1-
12
#4500000000
0!
0%
b1 *
0-
02
b1 6
#4510000000
1!
1%
1-
12
#4520000000
0!
0%
b10 *
0-
02
b10 6
#4530000000
1!
1%
1-
12
#4540000000
0!
0%
b11 *
0-
02
b11 6
#4550000000
1!
1%
1-
12
15
#4560000000
0!
0%
b100 *
0-
02
b100 6
#4570000000
1!
1%
1-
12
#4580000000
0!
0%
b101 *
0-
02
b101 6
#4590000000
1!
1%
1-
12
#4600000000
0!
0%
b110 *
0-
02
b110 6
#4610000000
1!
1%
1-
12
#4620000000
0!
0%
b111 *
0-
02
b111 6
#4630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#4640000000
0!
0%
b0 *
0-
02
b0 6
#4650000000
1!
1%
1-
12
#4660000000
0!
0%
b1 *
0-
02
b1 6
#4670000000
1!
1%
1-
12
#4680000000
0!
0%
b10 *
0-
02
b10 6
#4690000000
1!
1%
1-
12
#4700000000
0!
0%
b11 *
0-
02
b11 6
#4710000000
1!
1%
1-
12
15
#4720000000
0!
0%
b100 *
0-
02
b100 6
#4730000000
1!
1%
1-
12
#4740000000
0!
0%
b101 *
0-
02
b101 6
#4750000000
1!
1%
1-
12
#4760000000
0!
0%
b110 *
0-
02
b110 6
#4770000000
1!
1%
1-
12
#4780000000
0!
0%
b111 *
0-
02
b111 6
#4790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#4800000000
0!
0%
b0 *
0-
02
b0 6
#4810000000
1!
1%
1-
12
#4820000000
0!
0%
b1 *
0-
02
b1 6
#4830000000
1!
1%
1-
12
#4840000000
0!
0%
b10 *
0-
02
b10 6
#4850000000
1!
1%
1-
12
#4860000000
0!
0%
b11 *
0-
02
b11 6
#4870000000
1!
1%
1-
12
15
#4880000000
0!
0%
b100 *
0-
02
b100 6
#4890000000
1!
1%
1-
12
#4900000000
0!
0%
b101 *
0-
02
b101 6
#4910000000
1!
1%
1-
12
#4920000000
0!
0%
b110 *
0-
02
b110 6
#4930000000
1!
1%
1-
12
#4940000000
0!
0%
b111 *
0-
02
b111 6
#4950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#4960000000
0!
0%
b0 *
0-
02
b0 6
#4970000000
1!
1%
1-
12
#4980000000
0!
0%
b1 *
0-
02
b1 6
#4990000000
1!
1%
1-
12
#5000000000
0!
0%
b10 *
0-
02
b10 6
#5010000000
1!
1%
1-
12
#5020000000
0!
0%
b11 *
0-
02
b11 6
#5030000000
1!
1%
1-
12
15
#5040000000
0!
0%
b100 *
0-
02
b100 6
#5050000000
1!
1%
1-
12
#5060000000
0!
0%
b101 *
0-
02
b101 6
#5070000000
1!
1%
1-
12
#5080000000
0!
0%
b110 *
0-
02
b110 6
#5090000000
1!
1%
1-
12
#5100000000
0!
0%
b111 *
0-
02
b111 6
#5110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#5120000000
0!
0%
b0 *
0-
02
b0 6
#5130000000
1!
1%
1-
12
#5140000000
0!
0%
b1 *
0-
02
b1 6
#5150000000
1!
1%
1-
12
#5160000000
0!
0%
b10 *
0-
02
b10 6
#5170000000
1!
1%
1-
12
#5180000000
0!
0%
b11 *
0-
02
b11 6
#5190000000
1!
1%
1-
12
15
#5200000000
0!
0%
b100 *
0-
02
b100 6
#5210000000
1!
1%
1-
12
#5220000000
0!
0%
b101 *
0-
02
b101 6
#5230000000
1!
1%
1-
12
#5240000000
0!
0%
b110 *
0-
02
b110 6
#5250000000
1!
1%
1-
12
#5260000000
0!
0%
b111 *
0-
02
b111 6
#5270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#5280000000
0!
0%
b0 *
0-
02
b0 6
#5290000000
1!
1%
1-
12
#5300000000
0!
0%
b1 *
0-
02
b1 6
#5310000000
1!
1%
1-
12
#5320000000
0!
0%
b10 *
0-
02
b10 6
#5330000000
1!
1%
1-
12
#5340000000
0!
0%
b11 *
0-
02
b11 6
#5350000000
1!
1%
1-
12
15
#5360000000
0!
0%
b100 *
0-
02
b100 6
#5370000000
1!
1%
1-
12
#5380000000
0!
0%
b101 *
0-
02
b101 6
#5390000000
1!
1%
1-
12
#5400000000
0!
0%
b110 *
0-
02
b110 6
#5410000000
1!
1%
1-
12
#5420000000
0!
0%
b111 *
0-
02
b111 6
#5430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#5440000000
0!
0%
b0 *
0-
02
b0 6
#5450000000
1!
1%
1-
12
#5460000000
0!
0%
b1 *
0-
02
b1 6
#5470000000
1!
1%
1-
12
#5480000000
0!
0%
b10 *
0-
02
b10 6
#5490000000
1!
1%
1-
12
#5500000000
0!
0%
b11 *
0-
02
b11 6
#5510000000
1!
1%
1-
12
15
#5520000000
0!
0%
b100 *
0-
02
b100 6
#5530000000
1!
1%
1-
12
#5540000000
0!
0%
b101 *
0-
02
b101 6
#5550000000
1!
1%
1-
12
#5560000000
0!
0%
b110 *
0-
02
b110 6
#5570000000
1!
1%
1-
12
#5580000000
0!
0%
b111 *
0-
02
b111 6
#5590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#5600000000
0!
0%
b0 *
0-
02
b0 6
#5610000000
1!
1%
1-
12
#5620000000
0!
0%
b1 *
0-
02
b1 6
#5630000000
1!
1%
1-
12
#5640000000
0!
0%
b10 *
0-
02
b10 6
#5650000000
1!
1%
1-
12
#5660000000
0!
0%
b11 *
0-
02
b11 6
#5670000000
1!
1%
1-
12
15
#5680000000
0!
0%
b100 *
0-
02
b100 6
#5690000000
1!
1%
1-
12
#5700000000
0!
0%
b101 *
0-
02
b101 6
#5710000000
1!
1%
1-
12
#5720000000
0!
0%
b110 *
0-
02
b110 6
#5730000000
1!
1%
1-
12
#5740000000
0!
0%
b111 *
0-
02
b111 6
#5750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#5760000000
0!
0%
b0 *
0-
02
b0 6
#5770000000
1!
1%
1-
12
#5780000000
0!
0%
b1 *
0-
02
b1 6
#5790000000
1!
1%
1-
12
#5800000000
0!
0%
b10 *
0-
02
b10 6
#5810000000
1!
1%
1-
12
#5820000000
0!
0%
b11 *
0-
02
b11 6
#5830000000
1!
1%
1-
12
15
#5840000000
0!
0%
b100 *
0-
02
b100 6
#5850000000
1!
1%
1-
12
#5860000000
0!
0%
b101 *
0-
02
b101 6
#5870000000
1!
1%
1-
12
#5880000000
0!
0%
b110 *
0-
02
b110 6
#5890000000
1!
1%
1-
12
#5900000000
0!
0%
b111 *
0-
02
b111 6
#5910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#5920000000
0!
0%
b0 *
0-
02
b0 6
#5930000000
1!
1%
1-
12
#5940000000
0!
0%
b1 *
0-
02
b1 6
#5950000000
1!
1%
1-
12
#5960000000
0!
0%
b10 *
0-
02
b10 6
#5970000000
1!
1%
1-
12
#5980000000
0!
0%
b11 *
0-
02
b11 6
#5990000000
1!
1%
1-
12
15
#6000000000
0!
0%
b100 *
0-
02
b100 6
#6010000000
1!
1%
1-
12
#6020000000
0!
0%
b101 *
0-
02
b101 6
#6030000000
1!
1%
1-
12
#6040000000
0!
0%
b110 *
0-
02
b110 6
#6050000000
1!
1%
1-
12
#6060000000
0!
0%
b111 *
0-
02
b111 6
#6070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#6080000000
0!
0%
b0 *
0-
02
b0 6
#6090000000
1!
1%
1-
12
#6100000000
0!
0%
b1 *
0-
02
b1 6
#6110000000
1!
1%
1-
12
#6120000000
0!
0%
b10 *
0-
02
b10 6
#6130000000
1!
1%
1-
12
#6140000000
0!
0%
b11 *
0-
02
b11 6
#6150000000
1!
1%
1-
12
15
#6160000000
0!
0%
b100 *
0-
02
b100 6
#6170000000
1!
1%
1-
12
#6180000000
0!
0%
b101 *
0-
02
b101 6
#6190000000
1!
1%
1-
12
#6200000000
0!
0%
b110 *
0-
02
b110 6
#6210000000
1!
1%
1-
12
#6220000000
0!
0%
b111 *
0-
02
b111 6
#6230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#6240000000
0!
0%
b0 *
0-
02
b0 6
#6250000000
1!
1%
1-
12
#6260000000
0!
0%
b1 *
0-
02
b1 6
#6270000000
1!
1%
1-
12
#6280000000
0!
0%
b10 *
0-
02
b10 6
#6290000000
1!
1%
1-
12
#6300000000
0!
0%
b11 *
0-
02
b11 6
#6310000000
1!
1%
1-
12
15
#6320000000
0!
0%
b100 *
0-
02
b100 6
#6330000000
1!
1%
1-
12
#6340000000
0!
0%
b101 *
0-
02
b101 6
#6350000000
1!
1%
1-
12
#6360000000
0!
0%
b110 *
0-
02
b110 6
#6370000000
1!
1%
1-
12
#6380000000
0!
0%
b111 *
0-
02
b111 6
#6390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#6400000000
0!
0%
b0 *
0-
02
b0 6
#6410000000
1!
1%
1-
12
#6420000000
0!
0%
b1 *
0-
02
b1 6
#6430000000
1!
1%
1-
12
#6440000000
0!
0%
b10 *
0-
02
b10 6
#6450000000
1!
1%
1-
12
#6460000000
0!
0%
b11 *
0-
02
b11 6
#6470000000
1!
1%
1-
12
15
#6480000000
0!
0%
b100 *
0-
02
b100 6
#6490000000
1!
1%
1-
12
#6500000000
0!
0%
b101 *
0-
02
b101 6
#6510000000
1!
1%
1-
12
#6520000000
0!
0%
b110 *
0-
02
b110 6
#6530000000
1!
1%
1-
12
#6540000000
0!
0%
b111 *
0-
02
b111 6
#6550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#6560000000
0!
0%
b0 *
0-
02
b0 6
#6570000000
1!
1%
1-
12
#6580000000
0!
0%
b1 *
0-
02
b1 6
#6590000000
1!
1%
1-
12
#6600000000
0!
0%
b10 *
0-
02
b10 6
#6610000000
1!
1%
1-
12
#6620000000
0!
0%
b11 *
0-
02
b11 6
#6630000000
1!
1%
1-
12
15
#6640000000
0!
0%
b100 *
0-
02
b100 6
#6650000000
1!
1%
1-
12
#6660000000
0!
0%
b101 *
0-
02
b101 6
#6670000000
1!
1%
1-
12
#6680000000
0!
0%
b110 *
0-
02
b110 6
#6690000000
1!
1%
1-
12
#6700000000
0!
0%
b111 *
0-
02
b111 6
#6710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#6720000000
0!
0%
b0 *
0-
02
b0 6
#6730000000
1!
1%
1-
12
#6740000000
0!
0%
b1 *
0-
02
b1 6
#6750000000
1!
1%
1-
12
#6760000000
0!
0%
b10 *
0-
02
b10 6
#6770000000
1!
1%
1-
12
#6780000000
0!
0%
b11 *
0-
02
b11 6
#6790000000
1!
1%
1-
12
15
#6800000000
0!
0%
b100 *
0-
02
b100 6
#6810000000
1!
1%
1-
12
#6820000000
0!
0%
b101 *
0-
02
b101 6
#6830000000
1!
1%
1-
12
#6840000000
0!
0%
b110 *
0-
02
b110 6
#6850000000
1!
1%
1-
12
#6860000000
0!
0%
b111 *
0-
02
b111 6
#6870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#6880000000
0!
0%
b0 *
0-
02
b0 6
#6890000000
1!
1%
1-
12
#6900000000
0!
0%
b1 *
0-
02
b1 6
#6910000000
1!
1%
1-
12
#6920000000
0!
0%
b10 *
0-
02
b10 6
#6930000000
1!
1%
1-
12
#6940000000
0!
0%
b11 *
0-
02
b11 6
#6950000000
1!
1%
1-
12
15
#6960000000
0!
0%
b100 *
0-
02
b100 6
#6970000000
1!
1%
1-
12
#6980000000
0!
0%
b101 *
0-
02
b101 6
#6990000000
1!
1%
1-
12
#7000000000
0!
0%
b110 *
0-
02
b110 6
#7010000000
1!
1%
1-
12
#7020000000
0!
0%
b111 *
0-
02
b111 6
#7030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#7040000000
0!
0%
b0 *
0-
02
b0 6
#7050000000
1!
1%
1-
12
#7060000000
0!
0%
b1 *
0-
02
b1 6
#7070000000
1!
1%
1-
12
#7080000000
0!
0%
b10 *
0-
02
b10 6
#7090000000
1!
1%
1-
12
#7100000000
0!
0%
b11 *
0-
02
b11 6
#7110000000
1!
1%
1-
12
15
#7120000000
0!
0%
b100 *
0-
02
b100 6
#7130000000
1!
1%
1-
12
#7140000000
0!
0%
b101 *
0-
02
b101 6
#7150000000
1!
1%
1-
12
#7160000000
0!
0%
b110 *
0-
02
b110 6
#7170000000
1!
1%
1-
12
#7180000000
0!
0%
b111 *
0-
02
b111 6
#7190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#7200000000
0!
0%
b0 *
0-
02
b0 6
#7210000000
1!
1%
1-
12
#7220000000
0!
0%
b1 *
0-
02
b1 6
#7230000000
1!
1%
1-
12
#7240000000
0!
0%
b10 *
0-
02
b10 6
#7250000000
1!
1%
1-
12
#7260000000
0!
0%
b11 *
0-
02
b11 6
#7270000000
1!
1%
1-
12
15
#7280000000
0!
0%
b100 *
0-
02
b100 6
#7290000000
1!
1%
1-
12
#7300000000
0!
0%
b101 *
0-
02
b101 6
#7310000000
1!
1%
1-
12
#7320000000
0!
0%
b110 *
0-
02
b110 6
#7330000000
1!
1%
1-
12
#7340000000
0!
0%
b111 *
0-
02
b111 6
#7350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#7360000000
0!
0%
b0 *
0-
02
b0 6
#7370000000
1!
1%
1-
12
#7380000000
0!
0%
b1 *
0-
02
b1 6
#7390000000
1!
1%
1-
12
#7400000000
0!
0%
b10 *
0-
02
b10 6
#7410000000
1!
1%
1-
12
#7420000000
0!
0%
b11 *
0-
02
b11 6
#7430000000
1!
1%
1-
12
15
#7440000000
0!
0%
b100 *
0-
02
b100 6
#7450000000
1!
1%
1-
12
#7460000000
0!
0%
b101 *
0-
02
b101 6
#7470000000
1!
1%
1-
12
#7480000000
0!
0%
b110 *
0-
02
b110 6
#7490000000
1!
1%
1-
12
#7500000000
0!
0%
b111 *
0-
02
b111 6
#7510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#7520000000
0!
0%
b0 *
0-
02
b0 6
#7530000000
1!
1%
1-
12
#7540000000
0!
0%
b1 *
0-
02
b1 6
#7550000000
1!
1%
1-
12
#7560000000
0!
0%
b10 *
0-
02
b10 6
#7570000000
1!
1%
1-
12
#7580000000
0!
0%
b11 *
0-
02
b11 6
#7590000000
1!
1%
1-
12
15
#7600000000
0!
0%
b100 *
0-
02
b100 6
#7610000000
1!
1%
1-
12
#7620000000
0!
0%
b101 *
0-
02
b101 6
#7630000000
1!
1%
1-
12
#7640000000
0!
0%
b110 *
0-
02
b110 6
#7650000000
1!
1%
1-
12
#7660000000
0!
0%
b111 *
0-
02
b111 6
#7670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#7680000000
0!
0%
b0 *
0-
02
b0 6
#7690000000
1!
1%
1-
12
#7700000000
0!
0%
b1 *
0-
02
b1 6
#7710000000
1!
1%
1-
12
#7720000000
0!
0%
b10 *
0-
02
b10 6
#7730000000
1!
1%
1-
12
#7740000000
0!
0%
b11 *
0-
02
b11 6
#7750000000
1!
1%
1-
12
15
#7760000000
0!
0%
b100 *
0-
02
b100 6
#7770000000
1!
1%
1-
12
#7780000000
0!
0%
b101 *
0-
02
b101 6
#7790000000
1!
1%
1-
12
#7800000000
0!
0%
b110 *
0-
02
b110 6
#7810000000
1!
1%
1-
12
#7820000000
0!
0%
b111 *
0-
02
b111 6
#7830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#7840000000
0!
0%
b0 *
0-
02
b0 6
#7850000000
1!
1%
1-
12
#7860000000
0!
0%
b1 *
0-
02
b1 6
#7870000000
1!
1%
1-
12
#7880000000
0!
0%
b10 *
0-
02
b10 6
#7890000000
1!
1%
1-
12
#7900000000
0!
0%
b11 *
0-
02
b11 6
#7910000000
1!
1%
1-
12
15
#7920000000
0!
0%
b100 *
0-
02
b100 6
#7930000000
1!
1%
1-
12
#7940000000
0!
0%
b101 *
0-
02
b101 6
#7950000000
1!
1%
1-
12
#7960000000
0!
0%
b110 *
0-
02
b110 6
#7970000000
1!
1%
1-
12
#7980000000
0!
0%
b111 *
0-
02
b111 6
#7990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#8000000000
0!
0%
b0 *
0-
02
b0 6
#8010000000
1!
1%
1-
12
#8020000000
0!
0%
b1 *
0-
02
b1 6
#8030000000
1!
1%
1-
12
#8040000000
0!
0%
b10 *
0-
02
b10 6
#8050000000
1!
1%
1-
12
#8060000000
0!
0%
b11 *
0-
02
b11 6
#8070000000
1!
1%
1-
12
15
#8080000000
0!
0%
b100 *
0-
02
b100 6
#8090000000
1!
1%
1-
12
#8100000000
0!
0%
b101 *
0-
02
b101 6
#8110000000
1!
1%
1-
12
#8120000000
0!
0%
b110 *
0-
02
b110 6
#8130000000
1!
1%
1-
12
#8140000000
0!
0%
b111 *
0-
02
b111 6
#8150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#8160000000
0!
0%
b0 *
0-
02
b0 6
#8170000000
1!
1%
1-
12
#8180000000
0!
0%
b1 *
0-
02
b1 6
#8190000000
1!
1%
1-
12
#8200000000
0!
0%
b10 *
0-
02
b10 6
#8210000000
1!
1%
1-
12
#8220000000
0!
0%
b11 *
0-
02
b11 6
#8230000000
1!
1%
1-
12
15
#8240000000
0!
0%
b100 *
0-
02
b100 6
#8250000000
1!
1%
1-
12
#8260000000
0!
0%
b101 *
0-
02
b101 6
#8270000000
1!
1%
1-
12
#8280000000
0!
0%
b110 *
0-
02
b110 6
#8290000000
1!
1%
1-
12
#8300000000
0!
0%
b111 *
0-
02
b111 6
#8310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#8320000000
0!
0%
b0 *
0-
02
b0 6
#8330000000
1!
1%
1-
12
#8340000000
0!
0%
b1 *
0-
02
b1 6
#8350000000
1!
1%
1-
12
#8360000000
0!
0%
b10 *
0-
02
b10 6
#8370000000
1!
1%
1-
12
#8380000000
0!
0%
b11 *
0-
02
b11 6
#8390000000
1!
1%
1-
12
15
#8400000000
0!
0%
b100 *
0-
02
b100 6
#8410000000
1!
1%
1-
12
#8420000000
0!
0%
b101 *
0-
02
b101 6
#8430000000
1!
1%
1-
12
#8440000000
0!
0%
b110 *
0-
02
b110 6
#8450000000
1!
1%
1-
12
#8460000000
0!
0%
b111 *
0-
02
b111 6
#8470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#8480000000
0!
0%
b0 *
0-
02
b0 6
#8490000000
1!
1%
1-
12
#8500000000
0!
0%
b1 *
0-
02
b1 6
#8510000000
1!
1%
1-
12
#8520000000
0!
0%
b10 *
0-
02
b10 6
#8530000000
1!
1%
1-
12
#8540000000
0!
0%
b11 *
0-
02
b11 6
#8550000000
1!
1%
1-
12
15
#8560000000
0!
0%
b100 *
0-
02
b100 6
#8570000000
1!
1%
1-
12
#8580000000
0!
0%
b101 *
0-
02
b101 6
#8590000000
1!
1%
1-
12
#8600000000
0!
0%
b110 *
0-
02
b110 6
#8610000000
1!
1%
1-
12
#8620000000
0!
0%
b111 *
0-
02
b111 6
#8630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#8640000000
0!
0%
b0 *
0-
02
b0 6
#8650000000
1!
1%
1-
12
#8660000000
0!
0%
b1 *
0-
02
b1 6
#8670000000
1!
1%
1-
12
#8680000000
0!
0%
b10 *
0-
02
b10 6
#8690000000
1!
1%
1-
12
#8700000000
0!
0%
b11 *
0-
02
b11 6
#8710000000
1!
1%
1-
12
15
#8720000000
0!
0%
b100 *
0-
02
b100 6
#8730000000
1!
1%
1-
12
#8740000000
0!
0%
b101 *
0-
02
b101 6
#8750000000
1!
1%
1-
12
#8760000000
0!
0%
b110 *
0-
02
b110 6
#8770000000
1!
1%
1-
12
#8780000000
0!
0%
b111 *
0-
02
b111 6
#8790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#8800000000
0!
0%
b0 *
0-
02
b0 6
#8810000000
1!
1%
1-
12
#8820000000
0!
0%
b1 *
0-
02
b1 6
#8830000000
1!
1%
1-
12
#8840000000
0!
0%
b10 *
0-
02
b10 6
#8850000000
1!
1%
1-
12
#8860000000
0!
0%
b11 *
0-
02
b11 6
#8870000000
1!
1%
1-
12
15
#8880000000
0!
0%
b100 *
0-
02
b100 6
#8890000000
1!
1%
1-
12
#8900000000
0!
0%
b101 *
0-
02
b101 6
#8910000000
1!
1%
1-
12
#8920000000
0!
0%
b110 *
0-
02
b110 6
#8930000000
1!
1%
1-
12
#8940000000
0!
0%
b111 *
0-
02
b111 6
#8950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#8960000000
0!
0%
b0 *
0-
02
b0 6
#8970000000
1!
1%
1-
12
#8980000000
0!
0%
b1 *
0-
02
b1 6
#8990000000
1!
1%
1-
12
#9000000000
0!
0%
b10 *
0-
02
b10 6
#9010000000
1!
1%
1-
12
#9020000000
0!
0%
b11 *
0-
02
b11 6
#9030000000
1!
1%
1-
12
15
#9040000000
0!
0%
b100 *
0-
02
b100 6
#9050000000
1!
1%
1-
12
#9060000000
0!
0%
b101 *
0-
02
b101 6
#9070000000
1!
1%
1-
12
#9080000000
0!
0%
b110 *
0-
02
b110 6
#9090000000
1!
1%
1-
12
#9100000000
0!
0%
b111 *
0-
02
b111 6
#9110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#9120000000
0!
0%
b0 *
0-
02
b0 6
#9130000000
1!
1%
1-
12
#9140000000
0!
0%
b1 *
0-
02
b1 6
#9150000000
1!
1%
1-
12
#9160000000
0!
0%
b10 *
0-
02
b10 6
#9170000000
1!
1%
1-
12
#9180000000
0!
0%
b11 *
0-
02
b11 6
#9190000000
1!
1%
1-
12
15
#9200000000
0!
0%
b100 *
0-
02
b100 6
#9210000000
1!
1%
1-
12
#9220000000
0!
0%
b101 *
0-
02
b101 6
#9230000000
1!
1%
1-
12
#9240000000
0!
0%
b110 *
0-
02
b110 6
#9250000000
1!
1%
1-
12
#9260000000
0!
0%
b111 *
0-
02
b111 6
#9270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#9280000000
0!
0%
b0 *
0-
02
b0 6
#9290000000
1!
1%
1-
12
#9300000000
0!
0%
b1 *
0-
02
b1 6
#9310000000
1!
1%
1-
12
#9320000000
0!
0%
b10 *
0-
02
b10 6
#9330000000
1!
1%
1-
12
#9340000000
0!
0%
b11 *
0-
02
b11 6
#9350000000
1!
1%
1-
12
15
#9360000000
0!
0%
b100 *
0-
02
b100 6
#9370000000
1!
1%
1-
12
#9380000000
0!
0%
b101 *
0-
02
b101 6
#9390000000
1!
1%
1-
12
#9400000000
0!
0%
b110 *
0-
02
b110 6
#9410000000
1!
1%
1-
12
#9420000000
0!
0%
b111 *
0-
02
b111 6
#9430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#9440000000
0!
0%
b0 *
0-
02
b0 6
#9450000000
1!
1%
1-
12
#9460000000
0!
0%
b1 *
0-
02
b1 6
#9470000000
1!
1%
1-
12
#9480000000
0!
0%
b10 *
0-
02
b10 6
#9490000000
1!
1%
1-
12
#9500000000
0!
0%
b11 *
0-
02
b11 6
#9510000000
1!
1%
1-
12
15
#9520000000
0!
0%
b100 *
0-
02
b100 6
#9530000000
1!
1%
1-
12
#9540000000
0!
0%
b101 *
0-
02
b101 6
#9550000000
1!
1%
1-
12
#9560000000
0!
0%
b110 *
0-
02
b110 6
#9570000000
1!
1%
1-
12
#9580000000
0!
0%
b111 *
0-
02
b111 6
#9590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#9600000000
0!
0%
b0 *
0-
02
b0 6
#9610000000
1!
1%
1-
12
#9620000000
0!
0%
b1 *
0-
02
b1 6
#9630000000
1!
1%
1-
12
#9640000000
0!
0%
b10 *
0-
02
b10 6
#9650000000
1!
1%
1-
12
#9660000000
0!
0%
b11 *
0-
02
b11 6
#9670000000
1!
1%
1-
12
15
#9680000000
0!
0%
b100 *
0-
02
b100 6
#9690000000
1!
1%
1-
12
#9700000000
0!
0%
b101 *
0-
02
b101 6
#9710000000
1!
1%
1-
12
#9720000000
0!
0%
b110 *
0-
02
b110 6
#9730000000
1!
1%
1-
12
#9740000000
0!
0%
b111 *
0-
02
b111 6
#9750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#9760000000
0!
0%
b0 *
0-
02
b0 6
#9770000000
1!
1%
1-
12
#9780000000
0!
0%
b1 *
0-
02
b1 6
#9790000000
1!
1%
1-
12
#9800000000
0!
0%
b10 *
0-
02
b10 6
#9810000000
1!
1%
1-
12
#9820000000
0!
0%
b11 *
0-
02
b11 6
#9830000000
1!
1%
1-
12
15
#9840000000
0!
0%
b100 *
0-
02
b100 6
#9850000000
1!
1%
1-
12
#9860000000
0!
0%
b101 *
0-
02
b101 6
#9870000000
1!
1%
1-
12
#9880000000
0!
0%
b110 *
0-
02
b110 6
#9890000000
1!
1%
1-
12
#9900000000
0!
0%
b111 *
0-
02
b111 6
#9910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#9920000000
0!
0%
b0 *
0-
02
b0 6
#9930000000
1!
1%
1-
12
#9940000000
0!
0%
b1 *
0-
02
b1 6
#9950000000
1!
1%
1-
12
#9960000000
0!
0%
b10 *
0-
02
b10 6
#9970000000
1!
1%
1-
12
#9980000000
0!
0%
b11 *
0-
02
b11 6
#9990000000
1!
1%
1-
12
15
#10000000000
0!
0%
b100 *
0-
02
b100 6
#10010000000
1!
1%
1-
12
#10020000000
0!
0%
b101 *
0-
02
b101 6
#10030000000
1!
1%
1-
12
#10040000000
0!
0%
b110 *
0-
02
b110 6
#10050000000
1!
1%
1-
12
#10060000000
0!
0%
b111 *
0-
02
b111 6
#10070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#10080000000
0!
0%
b0 *
0-
02
b0 6
#10090000000
1!
1%
1-
12
#10100000000
0!
0%
b1 *
0-
02
b1 6
#10110000000
1!
1%
1-
12
#10120000000
0!
0%
b10 *
0-
02
b10 6
#10130000000
1!
1%
1-
12
#10140000000
0!
0%
b11 *
0-
02
b11 6
#10150000000
1!
1%
1-
12
15
#10160000000
0!
0%
b100 *
0-
02
b100 6
#10170000000
1!
1%
1-
12
#10180000000
0!
0%
b101 *
0-
02
b101 6
#10190000000
1!
1%
1-
12
#10200000000
0!
0%
b110 *
0-
02
b110 6
#10210000000
1!
1%
1-
12
#10220000000
0!
0%
b111 *
0-
02
b111 6
#10230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#10240000000
0!
0%
b0 *
0-
02
b0 6
#10250000000
1!
1%
1-
12
#10260000000
0!
0%
b1 *
0-
02
b1 6
#10270000000
1!
1%
1-
12
#10280000000
0!
0%
b10 *
0-
02
b10 6
#10290000000
1!
1%
1-
12
#10300000000
0!
0%
b11 *
0-
02
b11 6
#10310000000
1!
1%
1-
12
15
#10320000000
0!
0%
b100 *
0-
02
b100 6
#10330000000
1!
1%
1-
12
#10340000000
0!
0%
b101 *
0-
02
b101 6
#10350000000
1!
1%
1-
12
#10360000000
0!
0%
b110 *
0-
02
b110 6
#10370000000
1!
1%
1-
12
#10380000000
0!
0%
b111 *
0-
02
b111 6
#10390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#10400000000
0!
0%
b0 *
0-
02
b0 6
#10410000000
1!
1%
1-
12
#10420000000
0!
0%
b1 *
0-
02
b1 6
#10430000000
1!
1%
1-
12
#10440000000
0!
0%
b10 *
0-
02
b10 6
#10450000000
1!
1%
1-
12
#10460000000
0!
0%
b11 *
0-
02
b11 6
#10470000000
1!
1%
1-
12
15
#10480000000
0!
0%
b100 *
0-
02
b100 6
#10490000000
1!
1%
1-
12
#10500000000
0!
0%
b101 *
0-
02
b101 6
#10510000000
1!
1%
1-
12
#10520000000
0!
0%
b110 *
0-
02
b110 6
#10530000000
1!
1%
1-
12
#10540000000
0!
0%
b111 *
0-
02
b111 6
#10550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#10560000000
0!
0%
b0 *
0-
02
b0 6
#10570000000
1!
1%
1-
12
#10580000000
0!
0%
b1 *
0-
02
b1 6
#10590000000
1!
1%
1-
12
#10600000000
0!
0%
b10 *
0-
02
b10 6
#10610000000
1!
1%
1-
12
#10620000000
0!
0%
b11 *
0-
02
b11 6
#10630000000
1!
1%
1-
12
15
#10640000000
0!
0%
b100 *
0-
02
b100 6
#10650000000
1!
1%
1-
12
#10660000000
0!
0%
b101 *
0-
02
b101 6
#10670000000
1!
1%
1-
12
#10680000000
0!
0%
b110 *
0-
02
b110 6
#10690000000
1!
1%
1-
12
#10700000000
0!
0%
b111 *
0-
02
b111 6
#10710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#10720000000
0!
0%
b0 *
0-
02
b0 6
#10730000000
1!
1%
1-
12
#10740000000
0!
0%
b1 *
0-
02
b1 6
#10750000000
1!
1%
1-
12
#10760000000
0!
0%
b10 *
0-
02
b10 6
#10770000000
1!
1%
1-
12
#10780000000
0!
0%
b11 *
0-
02
b11 6
#10790000000
1!
1%
1-
12
15
#10800000000
0!
0%
b100 *
0-
02
b100 6
#10810000000
1!
1%
1-
12
#10820000000
0!
0%
b101 *
0-
02
b101 6
#10830000000
1!
1%
1-
12
#10840000000
0!
0%
b110 *
0-
02
b110 6
#10850000000
1!
1%
1-
12
#10860000000
0!
0%
b111 *
0-
02
b111 6
#10870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#10880000000
0!
0%
b0 *
0-
02
b0 6
#10890000000
1!
1%
1-
12
#10900000000
0!
0%
b1 *
0-
02
b1 6
#10910000000
1!
1%
1-
12
#10920000000
0!
0%
b10 *
0-
02
b10 6
#10930000000
1!
1%
1-
12
#10940000000
0!
0%
b11 *
0-
02
b11 6
#10950000000
1!
1%
1-
12
15
#10960000000
0!
0%
b100 *
0-
02
b100 6
#10970000000
1!
1%
1-
12
#10980000000
0!
0%
b101 *
0-
02
b101 6
#10990000000
1!
1%
1-
12
#11000000000
0!
0%
b110 *
0-
02
b110 6
#11010000000
1!
1%
1-
12
#11020000000
0!
0%
b111 *
0-
02
b111 6
#11030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#11040000000
0!
0%
b0 *
0-
02
b0 6
#11050000000
1!
1%
1-
12
#11060000000
0!
0%
b1 *
0-
02
b1 6
#11070000000
1!
1%
1-
12
#11080000000
0!
0%
b10 *
0-
02
b10 6
#11090000000
1!
1%
1-
12
#11100000000
0!
0%
b11 *
0-
02
b11 6
#11110000000
1!
1%
1-
12
15
#11120000000
0!
0%
b100 *
0-
02
b100 6
#11130000000
1!
1%
1-
12
#11140000000
0!
0%
b101 *
0-
02
b101 6
#11150000000
1!
1%
1-
12
#11160000000
0!
0%
b110 *
0-
02
b110 6
#11170000000
1!
1%
1-
12
#11180000000
0!
0%
b111 *
0-
02
b111 6
#11190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#11200000000
0!
0%
b0 *
0-
02
b0 6
#11210000000
1!
1%
1-
12
#11220000000
0!
0%
b1 *
0-
02
b1 6
#11230000000
1!
1%
1-
12
#11240000000
0!
0%
b10 *
0-
02
b10 6
#11250000000
1!
1%
1-
12
#11260000000
0!
0%
b11 *
0-
02
b11 6
#11270000000
1!
1%
1-
12
15
#11280000000
0!
0%
b100 *
0-
02
b100 6
#11290000000
1!
1%
1-
12
#11300000000
0!
0%
b101 *
0-
02
b101 6
#11310000000
1!
1%
1-
12
#11320000000
0!
0%
b110 *
0-
02
b110 6
#11330000000
1!
1%
1-
12
#11340000000
0!
0%
b111 *
0-
02
b111 6
#11350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#11360000000
0!
0%
b0 *
0-
02
b0 6
#11370000000
1!
1%
1-
12
#11380000000
0!
0%
b1 *
0-
02
b1 6
#11390000000
1!
1%
1-
12
#11400000000
0!
0%
b10 *
0-
02
b10 6
#11410000000
1!
1%
1-
12
#11420000000
0!
0%
b11 *
0-
02
b11 6
#11430000000
1!
1%
1-
12
15
#11440000000
0!
0%
b100 *
0-
02
b100 6
#11450000000
1!
1%
1-
12
#11460000000
0!
0%
b101 *
0-
02
b101 6
#11470000000
1!
1%
1-
12
#11480000000
0!
0%
b110 *
0-
02
b110 6
#11490000000
1!
1%
1-
12
#11500000000
0!
0%
b111 *
0-
02
b111 6
#11510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#11520000000
0!
0%
b0 *
0-
02
b0 6
#11530000000
1!
1%
1-
12
#11540000000
0!
0%
b1 *
0-
02
b1 6
#11550000000
1!
1%
1-
12
#11560000000
0!
0%
b10 *
0-
02
b10 6
#11570000000
1!
1%
1-
12
#11580000000
0!
0%
b11 *
0-
02
b11 6
#11590000000
1!
1%
1-
12
15
#11600000000
0!
0%
b100 *
0-
02
b100 6
#11610000000
1!
1%
1-
12
#11620000000
0!
0%
b101 *
0-
02
b101 6
#11630000000
1!
1%
1-
12
#11640000000
0!
0%
b110 *
0-
02
b110 6
#11650000000
1!
1%
1-
12
#11660000000
0!
0%
b111 *
0-
02
b111 6
#11670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#11680000000
0!
0%
b0 *
0-
02
b0 6
#11690000000
1!
1%
1-
12
#11700000000
0!
0%
b1 *
0-
02
b1 6
#11710000000
1!
1%
1-
12
#11720000000
0!
0%
b10 *
0-
02
b10 6
#11730000000
1!
1%
1-
12
#11740000000
0!
0%
b11 *
0-
02
b11 6
#11750000000
1!
1%
1-
12
15
#11760000000
0!
0%
b100 *
0-
02
b100 6
#11770000000
1!
1%
1-
12
#11780000000
0!
0%
b101 *
0-
02
b101 6
#11790000000
1!
1%
1-
12
#11800000000
0!
0%
b110 *
0-
02
b110 6
#11810000000
1!
1%
1-
12
#11820000000
0!
0%
b111 *
0-
02
b111 6
#11830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#11840000000
0!
0%
b0 *
0-
02
b0 6
#11850000000
1!
1%
1-
12
#11860000000
0!
0%
b1 *
0-
02
b1 6
#11870000000
1!
1%
1-
12
#11880000000
0!
0%
b10 *
0-
02
b10 6
#11890000000
1!
1%
1-
12
#11900000000
0!
0%
b11 *
0-
02
b11 6
#11910000000
1!
1%
1-
12
15
#11920000000
0!
0%
b100 *
0-
02
b100 6
#11930000000
1!
1%
1-
12
#11940000000
0!
0%
b101 *
0-
02
b101 6
#11950000000
1!
1%
1-
12
#11960000000
0!
0%
b110 *
0-
02
b110 6
#11970000000
1!
1%
1-
12
#11980000000
0!
0%
b111 *
0-
02
b111 6
#11990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#12000000000
0!
0%
b0 *
0-
02
b0 6
#12010000000
1!
1%
1-
12
#12020000000
0!
0%
b1 *
0-
02
b1 6
#12030000000
1!
1%
1-
12
#12040000000
0!
0%
b10 *
0-
02
b10 6
#12050000000
1!
1%
1-
12
#12060000000
0!
0%
b11 *
0-
02
b11 6
#12070000000
1!
1%
1-
12
15
#12080000000
0!
0%
b100 *
0-
02
b100 6
#12090000000
1!
1%
1-
12
#12100000000
0!
0%
b101 *
0-
02
b101 6
#12110000000
1!
1%
1-
12
#12120000000
0!
0%
b110 *
0-
02
b110 6
#12130000000
1!
1%
1-
12
#12140000000
0!
0%
b111 *
0-
02
b111 6
#12150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#12160000000
0!
0%
b0 *
0-
02
b0 6
#12170000000
1!
1%
1-
12
#12180000000
0!
0%
b1 *
0-
02
b1 6
#12190000000
1!
1%
1-
12
#12200000000
0!
0%
b10 *
0-
02
b10 6
#12210000000
1!
1%
1-
12
#12220000000
0!
0%
b11 *
0-
02
b11 6
#12230000000
1!
1%
1-
12
15
#12240000000
0!
0%
b100 *
0-
02
b100 6
#12250000000
1!
1%
1-
12
#12260000000
0!
0%
b101 *
0-
02
b101 6
#12270000000
1!
1%
1-
12
#12280000000
0!
0%
b110 *
0-
02
b110 6
#12290000000
1!
1%
1-
12
#12300000000
0!
0%
b111 *
0-
02
b111 6
#12310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#12320000000
0!
0%
b0 *
0-
02
b0 6
#12330000000
1!
1%
1-
12
#12340000000
0!
0%
b1 *
0-
02
b1 6
#12350000000
1!
1%
1-
12
#12360000000
0!
0%
b10 *
0-
02
b10 6
#12370000000
1!
1%
1-
12
#12380000000
0!
0%
b11 *
0-
02
b11 6
#12390000000
1!
1%
1-
12
15
#12400000000
0!
0%
b100 *
0-
02
b100 6
#12410000000
1!
1%
1-
12
#12420000000
0!
0%
b101 *
0-
02
b101 6
#12430000000
1!
1%
1-
12
#12440000000
0!
0%
b110 *
0-
02
b110 6
#12450000000
1!
1%
1-
12
#12460000000
0!
0%
b111 *
0-
02
b111 6
#12470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#12480000000
0!
0%
b0 *
0-
02
b0 6
#12490000000
1!
1%
1-
12
#12500000000
0!
0%
b1 *
0-
02
b1 6
#12510000000
1!
1%
1-
12
#12520000000
0!
0%
b10 *
0-
02
b10 6
#12530000000
1!
1%
1-
12
#12540000000
0!
0%
b11 *
0-
02
b11 6
#12550000000
1!
1%
1-
12
15
#12560000000
0!
0%
b100 *
0-
02
b100 6
#12570000000
1!
1%
1-
12
#12580000000
0!
0%
b101 *
0-
02
b101 6
#12590000000
1!
1%
1-
12
#12600000000
0!
0%
b110 *
0-
02
b110 6
#12610000000
1!
1%
1-
12
#12620000000
0!
0%
b111 *
0-
02
b111 6
#12630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#12640000000
0!
0%
b0 *
0-
02
b0 6
#12650000000
1!
1%
1-
12
#12660000000
0!
0%
b1 *
0-
02
b1 6
#12670000000
1!
1%
1-
12
#12680000000
0!
0%
b10 *
0-
02
b10 6
#12690000000
1!
1%
1-
12
#12700000000
0!
0%
b11 *
0-
02
b11 6
#12710000000
1!
1%
1-
12
15
#12720000000
0!
0%
b100 *
0-
02
b100 6
#12730000000
1!
1%
1-
12
#12740000000
0!
0%
b101 *
0-
02
b101 6
#12750000000
1!
1%
1-
12
#12760000000
0!
0%
b110 *
0-
02
b110 6
#12770000000
1!
1%
1-
12
#12780000000
0!
0%
b111 *
0-
02
b111 6
#12790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#12800000000
0!
0%
b0 *
0-
02
b0 6
#12810000000
1!
1%
1-
12
#12820000000
0!
0%
b1 *
0-
02
b1 6
#12830000000
1!
1%
1-
12
#12840000000
0!
0%
b10 *
0-
02
b10 6
#12850000000
1!
1%
1-
12
#12860000000
0!
0%
b11 *
0-
02
b11 6
#12870000000
1!
1%
1-
12
15
#12880000000
0!
0%
b100 *
0-
02
b100 6
#12890000000
1!
1%
1-
12
#12900000000
0!
0%
b101 *
0-
02
b101 6
#12910000000
1!
1%
1-
12
#12920000000
0!
0%
b110 *
0-
02
b110 6
#12930000000
1!
1%
1-
12
#12940000000
0!
0%
b111 *
0-
02
b111 6
#12950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#12960000000
0!
0%
b0 *
0-
02
b0 6
#12970000000
1!
1%
1-
12
#12980000000
0!
0%
b1 *
0-
02
b1 6
#12990000000
1!
1%
1-
12
#13000000000
0!
0%
b10 *
0-
02
b10 6
#13010000000
1!
1%
1-
12
#13020000000
0!
0%
b11 *
0-
02
b11 6
#13030000000
1!
1%
1-
12
15
#13040000000
0!
0%
b100 *
0-
02
b100 6
#13050000000
1!
1%
1-
12
#13060000000
0!
0%
b101 *
0-
02
b101 6
#13070000000
1!
1%
1-
12
#13080000000
0!
0%
b110 *
0-
02
b110 6
#13090000000
1!
1%
1-
12
#13100000000
0!
0%
b111 *
0-
02
b111 6
#13110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#13120000000
0!
0%
b0 *
0-
02
b0 6
#13130000000
1!
1%
1-
12
#13140000000
0!
0%
b1 *
0-
02
b1 6
#13150000000
1!
1%
1-
12
#13160000000
0!
0%
b10 *
0-
02
b10 6
#13170000000
1!
1%
1-
12
#13180000000
0!
0%
b11 *
0-
02
b11 6
#13190000000
1!
1%
1-
12
15
#13200000000
0!
0%
b100 *
0-
02
b100 6
#13210000000
1!
1%
1-
12
#13220000000
0!
0%
b101 *
0-
02
b101 6
#13230000000
1!
1%
1-
12
#13240000000
0!
0%
b110 *
0-
02
b110 6
#13250000000
1!
1%
1-
12
#13260000000
0!
0%
b111 *
0-
02
b111 6
#13270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#13280000000
0!
0%
b0 *
0-
02
b0 6
#13290000000
1!
1%
1-
12
#13300000000
0!
0%
b1 *
0-
02
b1 6
#13310000000
1!
1%
1-
12
#13320000000
0!
0%
b10 *
0-
02
b10 6
#13330000000
1!
1%
1-
12
#13340000000
0!
0%
b11 *
0-
02
b11 6
#13350000000
1!
1%
1-
12
15
#13360000000
0!
0%
b100 *
0-
02
b100 6
#13370000000
1!
1%
1-
12
#13380000000
0!
0%
b101 *
0-
02
b101 6
#13390000000
1!
1%
1-
12
#13400000000
0!
0%
b110 *
0-
02
b110 6
#13410000000
1!
1%
1-
12
#13420000000
0!
0%
b111 *
0-
02
b111 6
#13430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#13440000000
0!
0%
b0 *
0-
02
b0 6
#13450000000
1!
1%
1-
12
#13460000000
0!
0%
b1 *
0-
02
b1 6
#13470000000
1!
1%
1-
12
#13480000000
0!
0%
b10 *
0-
02
b10 6
#13490000000
1!
1%
1-
12
#13500000000
0!
0%
b11 *
0-
02
b11 6
#13510000000
1!
1%
1-
12
15
#13520000000
0!
0%
b100 *
0-
02
b100 6
#13530000000
1!
1%
1-
12
#13540000000
0!
0%
b101 *
0-
02
b101 6
#13550000000
1!
1%
1-
12
#13560000000
0!
0%
b110 *
0-
02
b110 6
#13570000000
1!
1%
1-
12
#13580000000
0!
0%
b111 *
0-
02
b111 6
#13590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#13600000000
0!
0%
b0 *
0-
02
b0 6
#13610000000
1!
1%
1-
12
#13620000000
0!
0%
b1 *
0-
02
b1 6
#13630000000
1!
1%
1-
12
#13640000000
0!
0%
b10 *
0-
02
b10 6
#13650000000
1!
1%
1-
12
#13660000000
0!
0%
b11 *
0-
02
b11 6
#13670000000
1!
1%
1-
12
15
#13680000000
0!
0%
b100 *
0-
02
b100 6
#13690000000
1!
1%
1-
12
#13700000000
0!
0%
b101 *
0-
02
b101 6
#13710000000
1!
1%
1-
12
#13720000000
0!
0%
b110 *
0-
02
b110 6
#13730000000
1!
1%
1-
12
#13740000000
0!
0%
b111 *
0-
02
b111 6
#13750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#13760000000
0!
0%
b0 *
0-
02
b0 6
#13770000000
1!
1%
1-
12
#13780000000
0!
0%
b1 *
0-
02
b1 6
#13790000000
1!
1%
1-
12
#13800000000
0!
0%
b10 *
0-
02
b10 6
#13810000000
1!
1%
1-
12
#13820000000
0!
0%
b11 *
0-
02
b11 6
#13830000000
1!
1%
1-
12
15
#13840000000
0!
0%
b100 *
0-
02
b100 6
#13850000000
1!
1%
1-
12
#13860000000
0!
0%
b101 *
0-
02
b101 6
#13870000000
1!
1%
1-
12
#13880000000
0!
0%
b110 *
0-
02
b110 6
#13890000000
1!
1%
1-
12
#13900000000
0!
0%
b111 *
0-
02
b111 6
#13910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#13920000000
0!
0%
b0 *
0-
02
b0 6
#13930000000
1!
1%
1-
12
#13940000000
0!
0%
b1 *
0-
02
b1 6
#13950000000
1!
1%
1-
12
#13960000000
0!
0%
b10 *
0-
02
b10 6
#13970000000
1!
1%
1-
12
#13980000000
0!
0%
b11 *
0-
02
b11 6
#13990000000
1!
1%
1-
12
15
#14000000000
0!
0%
b100 *
0-
02
b100 6
#14010000000
1!
1%
1-
12
#14020000000
0!
0%
b101 *
0-
02
b101 6
#14030000000
1!
1%
1-
12
#14040000000
0!
0%
b110 *
0-
02
b110 6
#14050000000
1!
1%
1-
12
#14060000000
0!
0%
b111 *
0-
02
b111 6
#14070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#14080000000
0!
0%
b0 *
0-
02
b0 6
#14090000000
1!
1%
1-
12
#14100000000
0!
0%
b1 *
0-
02
b1 6
#14110000000
1!
1%
1-
12
#14120000000
0!
0%
b10 *
0-
02
b10 6
#14130000000
1!
1%
1-
12
#14140000000
0!
0%
b11 *
0-
02
b11 6
#14150000000
1!
1%
1-
12
15
#14160000000
0!
0%
b100 *
0-
02
b100 6
#14170000000
1!
1%
1-
12
#14180000000
0!
0%
b101 *
0-
02
b101 6
#14190000000
1!
1%
1-
12
#14200000000
0!
0%
b110 *
0-
02
b110 6
#14210000000
1!
1%
1-
12
#14220000000
0!
0%
b111 *
0-
02
b111 6
#14230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#14240000000
0!
0%
b0 *
0-
02
b0 6
#14250000000
1!
1%
1-
12
#14260000000
0!
0%
b1 *
0-
02
b1 6
#14270000000
1!
1%
1-
12
#14280000000
0!
0%
b10 *
0-
02
b10 6
#14290000000
1!
1%
1-
12
#14300000000
0!
0%
b11 *
0-
02
b11 6
#14310000000
1!
1%
1-
12
15
#14320000000
0!
0%
b100 *
0-
02
b100 6
#14330000000
1!
1%
1-
12
#14340000000
0!
0%
b101 *
0-
02
b101 6
#14350000000
1!
1%
1-
12
#14360000000
0!
0%
b110 *
0-
02
b110 6
#14370000000
1!
1%
1-
12
#14380000000
0!
0%
b111 *
0-
02
b111 6
#14390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#14400000000
0!
0%
b0 *
0-
02
b0 6
#14410000000
1!
1%
1-
12
#14420000000
0!
0%
b1 *
0-
02
b1 6
#14430000000
1!
1%
1-
12
#14440000000
0!
0%
b10 *
0-
02
b10 6
#14450000000
1!
1%
1-
12
#14460000000
0!
0%
b11 *
0-
02
b11 6
#14470000000
1!
1%
1-
12
15
#14480000000
0!
0%
b100 *
0-
02
b100 6
#14490000000
1!
1%
1-
12
#14500000000
0!
0%
b101 *
0-
02
b101 6
#14510000000
1!
1%
1-
12
#14520000000
0!
0%
b110 *
0-
02
b110 6
#14530000000
1!
1%
1-
12
#14540000000
0!
0%
b111 *
0-
02
b111 6
#14550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#14560000000
0!
0%
b0 *
0-
02
b0 6
#14570000000
1!
1%
1-
12
#14580000000
0!
0%
b1 *
0-
02
b1 6
#14590000000
1!
1%
1-
12
#14600000000
0!
0%
b10 *
0-
02
b10 6
#14610000000
1!
1%
1-
12
#14620000000
0!
0%
b11 *
0-
02
b11 6
#14630000000
1!
1%
1-
12
15
#14640000000
0!
0%
b100 *
0-
02
b100 6
#14650000000
1!
1%
1-
12
#14660000000
0!
0%
b101 *
0-
02
b101 6
#14670000000
1!
1%
1-
12
#14680000000
0!
0%
b110 *
0-
02
b110 6
#14690000000
1!
1%
1-
12
#14700000000
0!
0%
b111 *
0-
02
b111 6
#14710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#14720000000
0!
0%
b0 *
0-
02
b0 6
#14730000000
1!
1%
1-
12
#14740000000
0!
0%
b1 *
0-
02
b1 6
#14750000000
1!
1%
1-
12
#14760000000
0!
0%
b10 *
0-
02
b10 6
#14770000000
1!
1%
1-
12
#14780000000
0!
0%
b11 *
0-
02
b11 6
#14790000000
1!
1%
1-
12
15
#14800000000
0!
0%
b100 *
0-
02
b100 6
#14810000000
1!
1%
1-
12
#14820000000
0!
0%
b101 *
0-
02
b101 6
#14830000000
1!
1%
1-
12
#14840000000
0!
0%
b110 *
0-
02
b110 6
#14850000000
1!
1%
1-
12
#14860000000
0!
0%
b111 *
0-
02
b111 6
#14870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#14880000000
0!
0%
b0 *
0-
02
b0 6
#14890000000
1!
1%
1-
12
#14900000000
0!
0%
b1 *
0-
02
b1 6
#14910000000
1!
1%
1-
12
#14920000000
0!
0%
b10 *
0-
02
b10 6
#14930000000
1!
1%
1-
12
#14940000000
0!
0%
b11 *
0-
02
b11 6
#14950000000
1!
1%
1-
12
15
#14960000000
0!
0%
b100 *
0-
02
b100 6
#14970000000
1!
1%
1-
12
#14980000000
0!
0%
b101 *
0-
02
b101 6
#14990000000
1!
1%
1-
12
#15000000000
0!
0%
b110 *
0-
02
b110 6
#15010000000
1!
1%
1-
12
#15020000000
0!
0%
b111 *
0-
02
b111 6
#15030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#15040000000
0!
0%
b0 *
0-
02
b0 6
#15050000000
1!
1%
1-
12
#15060000000
0!
0%
b1 *
0-
02
b1 6
#15070000000
1!
1%
1-
12
#15080000000
0!
0%
b10 *
0-
02
b10 6
#15090000000
1!
1%
1-
12
#15100000000
0!
0%
b11 *
0-
02
b11 6
#15110000000
1!
1%
1-
12
15
#15120000000
0!
0%
b100 *
0-
02
b100 6
#15130000000
1!
1%
1-
12
#15140000000
0!
0%
b101 *
0-
02
b101 6
#15150000000
1!
1%
1-
12
#15160000000
0!
0%
b110 *
0-
02
b110 6
#15170000000
1!
1%
1-
12
#15180000000
0!
0%
b111 *
0-
02
b111 6
#15190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#15200000000
0!
0%
b0 *
0-
02
b0 6
#15210000000
1!
1%
1-
12
#15220000000
0!
0%
b1 *
0-
02
b1 6
#15230000000
1!
1%
1-
12
#15240000000
0!
0%
b10 *
0-
02
b10 6
#15250000000
1!
1%
1-
12
#15260000000
0!
0%
b11 *
0-
02
b11 6
#15270000000
1!
1%
1-
12
15
#15280000000
0!
0%
b100 *
0-
02
b100 6
#15290000000
1!
1%
1-
12
#15300000000
0!
0%
b101 *
0-
02
b101 6
#15310000000
1!
1%
1-
12
#15320000000
0!
0%
b110 *
0-
02
b110 6
#15330000000
1!
1%
1-
12
#15340000000
0!
0%
b111 *
0-
02
b111 6
#15350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#15360000000
0!
0%
b0 *
0-
02
b0 6
#15370000000
1!
1%
1-
12
#15380000000
0!
0%
b1 *
0-
02
b1 6
#15390000000
1!
1%
1-
12
#15400000000
0!
0%
b10 *
0-
02
b10 6
#15410000000
1!
1%
1-
12
#15420000000
0!
0%
b11 *
0-
02
b11 6
#15430000000
1!
1%
1-
12
15
#15440000000
0!
0%
b100 *
0-
02
b100 6
#15450000000
1!
1%
1-
12
#15460000000
0!
0%
b101 *
0-
02
b101 6
#15470000000
1!
1%
1-
12
#15480000000
0!
0%
b110 *
0-
02
b110 6
#15490000000
1!
1%
1-
12
#15500000000
0!
0%
b111 *
0-
02
b111 6
#15510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#15520000000
0!
0%
b0 *
0-
02
b0 6
#15530000000
1!
1%
1-
12
#15540000000
0!
0%
b1 *
0-
02
b1 6
#15550000000
1!
1%
1-
12
#15560000000
0!
0%
b10 *
0-
02
b10 6
#15570000000
1!
1%
1-
12
#15580000000
0!
0%
b11 *
0-
02
b11 6
#15590000000
1!
1%
1-
12
15
#15600000000
0!
0%
b100 *
0-
02
b100 6
#15610000000
1!
1%
1-
12
#15620000000
0!
0%
b101 *
0-
02
b101 6
#15630000000
1!
1%
1-
12
#15640000000
0!
0%
b110 *
0-
02
b110 6
#15650000000
1!
1%
1-
12
#15660000000
0!
0%
b111 *
0-
02
b111 6
#15670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#15680000000
0!
0%
b0 *
0-
02
b0 6
#15690000000
1!
1%
1-
12
#15700000000
0!
0%
b1 *
0-
02
b1 6
#15710000000
1!
1%
1-
12
#15720000000
0!
0%
b10 *
0-
02
b10 6
#15730000000
1!
1%
1-
12
#15740000000
0!
0%
b11 *
0-
02
b11 6
#15750000000
1!
1%
1-
12
15
#15760000000
0!
0%
b100 *
0-
02
b100 6
#15770000000
1!
1%
1-
12
#15780000000
0!
0%
b101 *
0-
02
b101 6
#15790000000
1!
1%
1-
12
#15800000000
0!
0%
b110 *
0-
02
b110 6
#15810000000
1!
1%
1-
12
#15820000000
0!
0%
b111 *
0-
02
b111 6
#15830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#15840000000
0!
0%
b0 *
0-
02
b0 6
#15850000000
1!
1%
1-
12
#15860000000
0!
0%
b1 *
0-
02
b1 6
#15870000000
1!
1%
1-
12
#15880000000
0!
0%
b10 *
0-
02
b10 6
#15890000000
1!
1%
1-
12
#15900000000
0!
0%
b11 *
0-
02
b11 6
#15910000000
1!
1%
1-
12
15
#15920000000
0!
0%
b100 *
0-
02
b100 6
#15930000000
1!
1%
1-
12
#15940000000
0!
0%
b101 *
0-
02
b101 6
#15950000000
1!
1%
1-
12
#15960000000
0!
0%
b110 *
0-
02
b110 6
#15970000000
1!
1%
1-
12
#15980000000
0!
0%
b111 *
0-
02
b111 6
#15990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#16000000000
0!
0%
b0 *
0-
02
b0 6
#16010000000
1!
1%
1-
12
#16020000000
0!
0%
b1 *
0-
02
b1 6
#16030000000
1!
1%
1-
12
#16040000000
0!
0%
b10 *
0-
02
b10 6
#16050000000
1!
1%
1-
12
#16060000000
0!
0%
b11 *
0-
02
b11 6
#16070000000
1!
1%
1-
12
15
#16080000000
0!
0%
b100 *
0-
02
b100 6
#16090000000
1!
1%
1-
12
#16100000000
0!
0%
b101 *
0-
02
b101 6
#16110000000
1!
1%
1-
12
#16120000000
0!
0%
b110 *
0-
02
b110 6
#16130000000
1!
1%
1-
12
#16140000000
0!
0%
b111 *
0-
02
b111 6
#16150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#16160000000
0!
0%
b0 *
0-
02
b0 6
#16170000000
1!
1%
1-
12
#16180000000
0!
0%
b1 *
0-
02
b1 6
#16190000000
1!
1%
1-
12
#16200000000
0!
0%
b10 *
0-
02
b10 6
#16210000000
1!
1%
1-
12
#16220000000
0!
0%
b11 *
0-
02
b11 6
#16230000000
1!
1%
1-
12
15
#16240000000
0!
0%
b100 *
0-
02
b100 6
#16250000000
1!
1%
1-
12
#16260000000
0!
0%
b101 *
0-
02
b101 6
#16270000000
1!
1%
1-
12
#16280000000
0!
0%
b110 *
0-
02
b110 6
#16290000000
1!
1%
1-
12
#16300000000
0!
0%
b111 *
0-
02
b111 6
#16310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#16320000000
0!
0%
b0 *
0-
02
b0 6
#16330000000
1!
1%
1-
12
#16340000000
0!
0%
b1 *
0-
02
b1 6
#16350000000
1!
1%
1-
12
#16360000000
0!
0%
b10 *
0-
02
b10 6
#16370000000
1!
1%
1-
12
#16380000000
0!
0%
b11 *
0-
02
b11 6
#16390000000
1!
1%
1-
12
15
#16400000000
0!
0%
b100 *
0-
02
b100 6
#16410000000
1!
1%
1-
12
#16420000000
0!
0%
b101 *
0-
02
b101 6
#16430000000
1!
1%
1-
12
#16440000000
0!
0%
b110 *
0-
02
b110 6
#16450000000
1!
1%
1-
12
#16460000000
0!
0%
b111 *
0-
02
b111 6
#16470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#16480000000
0!
0%
b0 *
0-
02
b0 6
#16490000000
1!
1%
1-
12
#16500000000
0!
0%
b1 *
0-
02
b1 6
#16510000000
1!
1%
1-
12
#16520000000
0!
0%
b10 *
0-
02
b10 6
#16530000000
1!
1%
1-
12
#16540000000
0!
0%
b11 *
0-
02
b11 6
#16550000000
1!
1%
1-
12
15
#16560000000
0!
0%
b100 *
0-
02
b100 6
#16570000000
1!
1%
1-
12
#16580000000
0!
0%
b101 *
0-
02
b101 6
#16590000000
1!
1%
1-
12
#16600000000
0!
0%
b110 *
0-
02
b110 6
#16610000000
1!
1%
1-
12
#16620000000
0!
0%
b111 *
0-
02
b111 6
#16630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#16640000000
0!
0%
b0 *
0-
02
b0 6
#16650000000
1!
1%
1-
12
#16660000000
0!
0%
b1 *
0-
02
b1 6
#16670000000
1!
1%
1-
12
#16680000000
0!
0%
b10 *
0-
02
b10 6
#16690000000
1!
1%
1-
12
#16700000000
0!
0%
b11 *
0-
02
b11 6
#16710000000
1!
1%
1-
12
15
#16720000000
0!
0%
b100 *
0-
02
b100 6
#16730000000
1!
1%
1-
12
#16740000000
0!
0%
b101 *
0-
02
b101 6
#16750000000
1!
1%
1-
12
#16760000000
0!
0%
b110 *
0-
02
b110 6
#16770000000
1!
1%
1-
12
#16780000000
0!
0%
b111 *
0-
02
b111 6
#16790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#16800000000
0!
0%
b0 *
0-
02
b0 6
#16810000000
1!
1%
1-
12
#16820000000
0!
0%
b1 *
0-
02
b1 6
#16830000000
1!
1%
1-
12
#16840000000
0!
0%
b10 *
0-
02
b10 6
#16850000000
1!
1%
1-
12
#16860000000
0!
0%
b11 *
0-
02
b11 6
#16870000000
1!
1%
1-
12
15
#16880000000
0!
0%
b100 *
0-
02
b100 6
#16890000000
1!
1%
1-
12
#16900000000
0!
0%
b101 *
0-
02
b101 6
#16910000000
1!
1%
1-
12
#16920000000
0!
0%
b110 *
0-
02
b110 6
#16930000000
1!
1%
1-
12
#16940000000
0!
0%
b111 *
0-
02
b111 6
#16950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#16960000000
0!
0%
b0 *
0-
02
b0 6
#16970000000
1!
1%
1-
12
#16980000000
0!
0%
b1 *
0-
02
b1 6
#16990000000
1!
1%
1-
12
#17000000000
0!
0%
b10 *
0-
02
b10 6
#17010000000
1!
1%
1-
12
#17020000000
0!
0%
b11 *
0-
02
b11 6
#17030000000
1!
1%
1-
12
15
#17040000000
0!
0%
b100 *
0-
02
b100 6
#17050000000
1!
1%
1-
12
#17060000000
0!
0%
b101 *
0-
02
b101 6
#17070000000
1!
1%
1-
12
#17080000000
0!
0%
b110 *
0-
02
b110 6
#17090000000
1!
1%
1-
12
#17100000000
0!
0%
b111 *
0-
02
b111 6
#17110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#17120000000
0!
0%
b0 *
0-
02
b0 6
#17130000000
1!
1%
1-
12
#17140000000
0!
0%
b1 *
0-
02
b1 6
#17150000000
1!
1%
1-
12
#17160000000
0!
0%
b10 *
0-
02
b10 6
#17170000000
1!
1%
1-
12
#17180000000
0!
0%
b11 *
0-
02
b11 6
#17190000000
1!
1%
1-
12
15
#17200000000
0!
0%
b100 *
0-
02
b100 6
#17210000000
1!
1%
1-
12
#17220000000
0!
0%
b101 *
0-
02
b101 6
#17230000000
1!
1%
1-
12
#17240000000
0!
0%
b110 *
0-
02
b110 6
#17250000000
1!
1%
1-
12
#17260000000
0!
0%
b111 *
0-
02
b111 6
#17270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#17280000000
0!
0%
b0 *
0-
02
b0 6
#17290000000
1!
1%
1-
12
#17300000000
0!
0%
b1 *
0-
02
b1 6
#17310000000
1!
1%
1-
12
#17320000000
0!
0%
b10 *
0-
02
b10 6
#17330000000
1!
1%
1-
12
#17340000000
0!
0%
b11 *
0-
02
b11 6
#17350000000
1!
1%
1-
12
15
#17360000000
0!
0%
b100 *
0-
02
b100 6
#17370000000
1!
1%
1-
12
#17380000000
0!
0%
b101 *
0-
02
b101 6
#17390000000
1!
1%
1-
12
#17400000000
0!
0%
b110 *
0-
02
b110 6
#17410000000
1!
1%
1-
12
#17420000000
0!
0%
b111 *
0-
02
b111 6
#17430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#17440000000
0!
0%
b0 *
0-
02
b0 6
#17450000000
1!
1%
1-
12
#17460000000
0!
0%
b1 *
0-
02
b1 6
#17470000000
1!
1%
1-
12
#17480000000
0!
0%
b10 *
0-
02
b10 6
#17490000000
1!
1%
1-
12
#17500000000
0!
0%
b11 *
0-
02
b11 6
#17510000000
1!
1%
1-
12
15
#17520000000
0!
0%
b100 *
0-
02
b100 6
#17530000000
1!
1%
1-
12
#17540000000
0!
0%
b101 *
0-
02
b101 6
#17550000000
1!
1%
1-
12
#17560000000
0!
0%
b110 *
0-
02
b110 6
#17570000000
1!
1%
1-
12
#17580000000
0!
0%
b111 *
0-
02
b111 6
#17590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#17600000000
0!
0%
b0 *
0-
02
b0 6
#17610000000
1!
1%
1-
12
#17620000000
0!
0%
b1 *
0-
02
b1 6
#17630000000
1!
1%
1-
12
#17640000000
0!
0%
b10 *
0-
02
b10 6
#17650000000
1!
1%
1-
12
#17660000000
0!
0%
b11 *
0-
02
b11 6
#17670000000
1!
1%
1-
12
15
#17680000000
0!
0%
b100 *
0-
02
b100 6
#17690000000
1!
1%
1-
12
#17700000000
0!
0%
b101 *
0-
02
b101 6
#17710000000
1!
1%
1-
12
#17720000000
0!
0%
b110 *
0-
02
b110 6
#17730000000
1!
1%
1-
12
#17740000000
0!
0%
b111 *
0-
02
b111 6
#17750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#17760000000
0!
0%
b0 *
0-
02
b0 6
#17770000000
1!
1%
1-
12
#17780000000
0!
0%
b1 *
0-
02
b1 6
#17790000000
1!
1%
1-
12
#17800000000
0!
0%
b10 *
0-
02
b10 6
#17810000000
1!
1%
1-
12
#17820000000
0!
0%
b11 *
0-
02
b11 6
#17830000000
1!
1%
1-
12
15
#17840000000
0!
0%
b100 *
0-
02
b100 6
#17850000000
1!
1%
1-
12
#17860000000
0!
0%
b101 *
0-
02
b101 6
#17870000000
1!
1%
1-
12
#17880000000
0!
0%
b110 *
0-
02
b110 6
#17890000000
1!
1%
1-
12
#17900000000
0!
0%
b111 *
0-
02
b111 6
#17910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#17920000000
0!
0%
b0 *
0-
02
b0 6
#17930000000
1!
1%
1-
12
#17940000000
0!
0%
b1 *
0-
02
b1 6
#17950000000
1!
1%
1-
12
#17960000000
0!
0%
b10 *
0-
02
b10 6
#17970000000
1!
1%
1-
12
#17980000000
0!
0%
b11 *
0-
02
b11 6
#17990000000
1!
1%
1-
12
15
#18000000000
0!
0%
b100 *
0-
02
b100 6
#18010000000
1!
1%
1-
12
#18020000000
0!
0%
b101 *
0-
02
b101 6
#18030000000
1!
1%
1-
12
#18040000000
0!
0%
b110 *
0-
02
b110 6
#18050000000
1!
1%
1-
12
#18060000000
0!
0%
b111 *
0-
02
b111 6
#18070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#18080000000
0!
0%
b0 *
0-
02
b0 6
#18090000000
1!
1%
1-
12
#18100000000
0!
0%
b1 *
0-
02
b1 6
#18110000000
1!
1%
1-
12
#18120000000
0!
0%
b10 *
0-
02
b10 6
#18130000000
1!
1%
1-
12
#18140000000
0!
0%
b11 *
0-
02
b11 6
#18150000000
1!
1%
1-
12
15
#18160000000
0!
0%
b100 *
0-
02
b100 6
#18170000000
1!
1%
1-
12
#18180000000
0!
0%
b101 *
0-
02
b101 6
#18190000000
1!
1%
1-
12
#18200000000
0!
0%
b110 *
0-
02
b110 6
#18210000000
1!
1%
1-
12
#18220000000
0!
0%
b111 *
0-
02
b111 6
#18230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#18240000000
0!
0%
b0 *
0-
02
b0 6
#18250000000
1!
1%
1-
12
#18260000000
0!
0%
b1 *
0-
02
b1 6
#18270000000
1!
1%
1-
12
#18280000000
0!
0%
b10 *
0-
02
b10 6
#18290000000
1!
1%
1-
12
#18300000000
0!
0%
b11 *
0-
02
b11 6
#18310000000
1!
1%
1-
12
15
#18320000000
0!
0%
b100 *
0-
02
b100 6
#18330000000
1!
1%
1-
12
#18340000000
0!
0%
b101 *
0-
02
b101 6
#18350000000
1!
1%
1-
12
#18360000000
0!
0%
b110 *
0-
02
b110 6
#18370000000
1!
1%
1-
12
#18380000000
0!
0%
b111 *
0-
02
b111 6
#18390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#18400000000
0!
0%
b0 *
0-
02
b0 6
#18410000000
1!
1%
1-
12
#18420000000
0!
0%
b1 *
0-
02
b1 6
#18430000000
1!
1%
1-
12
#18440000000
0!
0%
b10 *
0-
02
b10 6
#18450000000
1!
1%
1-
12
#18460000000
0!
0%
b11 *
0-
02
b11 6
#18470000000
1!
1%
1-
12
15
#18480000000
0!
0%
b100 *
0-
02
b100 6
#18490000000
1!
1%
1-
12
#18500000000
0!
0%
b101 *
0-
02
b101 6
#18510000000
1!
1%
1-
12
#18520000000
0!
0%
b110 *
0-
02
b110 6
#18530000000
1!
1%
1-
12
#18540000000
0!
0%
b111 *
0-
02
b111 6
#18550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#18560000000
0!
0%
b0 *
0-
02
b0 6
#18570000000
1!
1%
1-
12
#18580000000
0!
0%
b1 *
0-
02
b1 6
#18590000000
1!
1%
1-
12
#18600000000
0!
0%
b10 *
0-
02
b10 6
#18610000000
1!
1%
1-
12
#18620000000
0!
0%
b11 *
0-
02
b11 6
#18630000000
1!
1%
1-
12
15
#18640000000
0!
0%
b100 *
0-
02
b100 6
#18650000000
1!
1%
1-
12
#18660000000
0!
0%
b101 *
0-
02
b101 6
#18670000000
1!
1%
1-
12
#18680000000
0!
0%
b110 *
0-
02
b110 6
#18690000000
1!
1%
1-
12
#18700000000
0!
0%
b111 *
0-
02
b111 6
#18710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#18720000000
0!
0%
b0 *
0-
02
b0 6
#18730000000
1!
1%
1-
12
#18740000000
0!
0%
b1 *
0-
02
b1 6
#18750000000
1!
1%
1-
12
#18760000000
0!
0%
b10 *
0-
02
b10 6
#18770000000
1!
1%
1-
12
#18780000000
0!
0%
b11 *
0-
02
b11 6
#18790000000
1!
1%
1-
12
15
#18800000000
0!
0%
b100 *
0-
02
b100 6
#18810000000
1!
1%
1-
12
#18820000000
0!
0%
b101 *
0-
02
b101 6
#18830000000
1!
1%
1-
12
#18840000000
0!
0%
b110 *
0-
02
b110 6
#18850000000
1!
1%
1-
12
#18860000000
0!
0%
b111 *
0-
02
b111 6
#18870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#18880000000
0!
0%
b0 *
0-
02
b0 6
#18890000000
1!
1%
1-
12
#18900000000
0!
0%
b1 *
0-
02
b1 6
#18910000000
1!
1%
1-
12
#18920000000
0!
0%
b10 *
0-
02
b10 6
#18930000000
1!
1%
1-
12
#18940000000
0!
0%
b11 *
0-
02
b11 6
#18950000000
1!
1%
1-
12
15
#18960000000
0!
0%
b100 *
0-
02
b100 6
#18970000000
1!
1%
1-
12
#18980000000
0!
0%
b101 *
0-
02
b101 6
#18990000000
1!
1%
1-
12
#19000000000
0!
0%
b110 *
0-
02
b110 6
#19010000000
1!
1%
1-
12
#19020000000
0!
0%
b111 *
0-
02
b111 6
#19030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#19040000000
0!
0%
b0 *
0-
02
b0 6
#19050000000
1!
1%
1-
12
#19060000000
0!
0%
b1 *
0-
02
b1 6
#19070000000
1!
1%
1-
12
#19080000000
0!
0%
b10 *
0-
02
b10 6
#19090000000
1!
1%
1-
12
#19100000000
0!
0%
b11 *
0-
02
b11 6
#19110000000
1!
1%
1-
12
15
#19120000000
0!
0%
b100 *
0-
02
b100 6
#19130000000
1!
1%
1-
12
#19140000000
0!
0%
b101 *
0-
02
b101 6
#19150000000
1!
1%
1-
12
#19160000000
0!
0%
b110 *
0-
02
b110 6
#19170000000
1!
1%
1-
12
#19180000000
0!
0%
b111 *
0-
02
b111 6
#19190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#19200000000
0!
0%
b0 *
0-
02
b0 6
#19210000000
1!
1%
1-
12
#19220000000
0!
0%
b1 *
0-
02
b1 6
#19230000000
1!
1%
1-
12
#19240000000
0!
0%
b10 *
0-
02
b10 6
#19250000000
1!
1%
1-
12
#19260000000
0!
0%
b11 *
0-
02
b11 6
#19270000000
1!
1%
1-
12
15
#19280000000
0!
0%
b100 *
0-
02
b100 6
#19290000000
1!
1%
1-
12
#19300000000
0!
0%
b101 *
0-
02
b101 6
#19310000000
1!
1%
1-
12
#19320000000
0!
0%
b110 *
0-
02
b110 6
#19330000000
1!
1%
1-
12
#19340000000
0!
0%
b111 *
0-
02
b111 6
#19350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#19360000000
0!
0%
b0 *
0-
02
b0 6
#19370000000
1!
1%
1-
12
#19380000000
0!
0%
b1 *
0-
02
b1 6
#19390000000
1!
1%
1-
12
#19400000000
0!
0%
b10 *
0-
02
b10 6
#19410000000
1!
1%
1-
12
#19420000000
0!
0%
b11 *
0-
02
b11 6
#19430000000
1!
1%
1-
12
15
#19440000000
0!
0%
b100 *
0-
02
b100 6
#19450000000
1!
1%
1-
12
#19460000000
0!
0%
b101 *
0-
02
b101 6
#19470000000
1!
1%
1-
12
#19480000000
0!
0%
b110 *
0-
02
b110 6
#19490000000
1!
1%
1-
12
#19500000000
0!
0%
b111 *
0-
02
b111 6
#19510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#19520000000
0!
0%
b0 *
0-
02
b0 6
#19530000000
1!
1%
1-
12
#19540000000
0!
0%
b1 *
0-
02
b1 6
#19550000000
1!
1%
1-
12
#19560000000
0!
0%
b10 *
0-
02
b10 6
#19570000000
1!
1%
1-
12
#19580000000
0!
0%
b11 *
0-
02
b11 6
#19590000000
1!
1%
1-
12
15
#19600000000
0!
0%
b100 *
0-
02
b100 6
#19610000000
1!
1%
1-
12
#19620000000
0!
0%
b101 *
0-
02
b101 6
#19630000000
1!
1%
1-
12
#19640000000
0!
0%
b110 *
0-
02
b110 6
#19650000000
1!
1%
1-
12
#19660000000
0!
0%
b111 *
0-
02
b111 6
#19670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#19680000000
0!
0%
b0 *
0-
02
b0 6
#19690000000
1!
1%
1-
12
#19700000000
0!
0%
b1 *
0-
02
b1 6
#19710000000
1!
1%
1-
12
#19720000000
0!
0%
b10 *
0-
02
b10 6
#19730000000
1!
1%
1-
12
#19740000000
0!
0%
b11 *
0-
02
b11 6
#19750000000
1!
1%
1-
12
15
#19760000000
0!
0%
b100 *
0-
02
b100 6
#19770000000
1!
1%
1-
12
#19780000000
0!
0%
b101 *
0-
02
b101 6
#19790000000
1!
1%
1-
12
#19800000000
0!
0%
b110 *
0-
02
b110 6
#19810000000
1!
1%
1-
12
#19820000000
0!
0%
b111 *
0-
02
b111 6
#19830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#19840000000
0!
0%
b0 *
0-
02
b0 6
#19850000000
1!
1%
1-
12
#19860000000
0!
0%
b1 *
0-
02
b1 6
#19870000000
1!
1%
1-
12
#19880000000
0!
0%
b10 *
0-
02
b10 6
#19890000000
1!
1%
1-
12
#19900000000
0!
0%
b11 *
0-
02
b11 6
#19910000000
1!
1%
1-
12
15
#19920000000
0!
0%
b100 *
0-
02
b100 6
#19930000000
1!
1%
1-
12
#19940000000
0!
0%
b101 *
0-
02
b101 6
#19950000000
1!
1%
1-
12
#19960000000
0!
0%
b110 *
0-
02
b110 6
#19970000000
1!
1%
1-
12
#19980000000
0!
0%
b111 *
0-
02
b111 6
#19990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#20000000000
0!
0%
b0 *
0-
02
b0 6
#20010000000
1!
1%
1-
12
#20020000000
0!
0%
b1 *
0-
02
b1 6
#20030000000
1!
1%
1-
12
#20040000000
0!
0%
b10 *
0-
02
b10 6
#20050000000
1!
1%
1-
12
#20060000000
0!
0%
b11 *
0-
02
b11 6
#20070000000
1!
1%
1-
12
15
#20080000000
0!
0%
b100 *
0-
02
b100 6
#20090000000
1!
1%
1-
12
#20100000000
0!
0%
b101 *
0-
02
b101 6
#20110000000
1!
1%
1-
12
#20120000000
0!
0%
b110 *
0-
02
b110 6
#20130000000
1!
1%
1-
12
#20140000000
0!
0%
b111 *
0-
02
b111 6
#20150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#20160000000
0!
0%
b0 *
0-
02
b0 6
#20170000000
1!
1%
1-
12
#20180000000
0!
0%
b1 *
0-
02
b1 6
#20190000000
1!
1%
1-
12
#20200000000
0!
0%
b10 *
0-
02
b10 6
#20210000000
1!
1%
1-
12
#20220000000
0!
0%
b11 *
0-
02
b11 6
#20230000000
1!
1%
1-
12
15
#20240000000
0!
0%
b100 *
0-
02
b100 6
#20250000000
1!
1%
1-
12
#20260000000
0!
0%
b101 *
0-
02
b101 6
#20270000000
1!
1%
1-
12
#20280000000
0!
0%
b110 *
0-
02
b110 6
#20290000000
1!
1%
1-
12
#20300000000
0!
0%
b111 *
0-
02
b111 6
#20310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#20320000000
0!
0%
b0 *
0-
02
b0 6
#20330000000
1!
1%
1-
12
#20340000000
0!
0%
b1 *
0-
02
b1 6
#20350000000
1!
1%
1-
12
#20360000000
0!
0%
b10 *
0-
02
b10 6
#20370000000
1!
1%
1-
12
#20380000000
0!
0%
b11 *
0-
02
b11 6
#20390000000
1!
1%
1-
12
15
#20400000000
0!
0%
b100 *
0-
02
b100 6
#20410000000
1!
1%
1-
12
#20420000000
0!
0%
b101 *
0-
02
b101 6
#20430000000
1!
1%
1-
12
#20440000000
0!
0%
b110 *
0-
02
b110 6
#20450000000
1!
1%
1-
12
#20460000000
0!
0%
b111 *
0-
02
b111 6
#20470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#20480000000
0!
0%
b0 *
0-
02
b0 6
#20490000000
1!
1%
1-
12
#20500000000
0!
0%
b1 *
0-
02
b1 6
#20510000000
1!
1%
1-
12
#20520000000
0!
0%
b10 *
0-
02
b10 6
#20530000000
1!
1%
1-
12
#20540000000
0!
0%
b11 *
0-
02
b11 6
#20550000000
1!
1%
1-
12
15
#20560000000
0!
0%
b100 *
0-
02
b100 6
#20570000000
1!
1%
1-
12
#20580000000
0!
0%
b101 *
0-
02
b101 6
#20590000000
1!
1%
1-
12
#20600000000
0!
0%
b110 *
0-
02
b110 6
#20610000000
1!
1%
1-
12
#20620000000
0!
0%
b111 *
0-
02
b111 6
#20630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#20640000000
0!
0%
b0 *
0-
02
b0 6
#20650000000
1!
1%
1-
12
#20660000000
0!
0%
b1 *
0-
02
b1 6
#20670000000
1!
1%
1-
12
#20680000000
0!
0%
b10 *
0-
02
b10 6
#20690000000
1!
1%
1-
12
#20700000000
0!
0%
b11 *
0-
02
b11 6
#20710000000
1!
1%
1-
12
15
#20720000000
0!
0%
b100 *
0-
02
b100 6
#20730000000
1!
1%
1-
12
#20740000000
0!
0%
b101 *
0-
02
b101 6
#20750000000
1!
1%
1-
12
#20760000000
0!
0%
b110 *
0-
02
b110 6
#20770000000
1!
1%
1-
12
#20780000000
0!
0%
b111 *
0-
02
b111 6
#20790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#20800000000
0!
0%
b0 *
0-
02
b0 6
#20810000000
1!
1%
1-
12
#20820000000
0!
0%
b1 *
0-
02
b1 6
#20830000000
1!
1%
1-
12
#20840000000
0!
0%
b10 *
0-
02
b10 6
#20850000000
1!
1%
1-
12
#20860000000
0!
0%
b11 *
0-
02
b11 6
#20870000000
1!
1%
1-
12
15
#20880000000
0!
0%
b100 *
0-
02
b100 6
#20890000000
1!
1%
1-
12
#20900000000
0!
0%
b101 *
0-
02
b101 6
#20910000000
1!
1%
1-
12
#20920000000
0!
0%
b110 *
0-
02
b110 6
#20930000000
1!
1%
1-
12
#20940000000
0!
0%
b111 *
0-
02
b111 6
#20950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#20960000000
0!
0%
b0 *
0-
02
b0 6
#20970000000
1!
1%
1-
12
#20980000000
0!
0%
b1 *
0-
02
b1 6
#20990000000
1!
1%
1-
12
#21000000000
0!
0%
b10 *
0-
02
b10 6
#21010000000
1!
1%
1-
12
#21020000000
0!
0%
b11 *
0-
02
b11 6
#21030000000
1!
1%
1-
12
15
#21040000000
0!
0%
b100 *
0-
02
b100 6
#21050000000
1!
1%
1-
12
#21060000000
0!
0%
b101 *
0-
02
b101 6
#21070000000
1!
1%
1-
12
#21080000000
0!
0%
b110 *
0-
02
b110 6
#21090000000
1!
1%
1-
12
#21100000000
0!
0%
b111 *
0-
02
b111 6
#21110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#21120000000
0!
0%
b0 *
0-
02
b0 6
#21130000000
1!
1%
1-
12
#21140000000
0!
0%
b1 *
0-
02
b1 6
#21150000000
1!
1%
1-
12
#21160000000
0!
0%
b10 *
0-
02
b10 6
#21170000000
1!
1%
1-
12
#21180000000
0!
0%
b11 *
0-
02
b11 6
#21190000000
1!
1%
1-
12
15
#21200000000
0!
0%
b100 *
0-
02
b100 6
#21210000000
1!
1%
1-
12
#21220000000
0!
0%
b101 *
0-
02
b101 6
#21230000000
1!
1%
1-
12
#21240000000
0!
0%
b110 *
0-
02
b110 6
#21250000000
1!
1%
1-
12
#21260000000
0!
0%
b111 *
0-
02
b111 6
#21270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#21280000000
0!
0%
b0 *
0-
02
b0 6
#21290000000
1!
1%
1-
12
#21300000000
0!
0%
b1 *
0-
02
b1 6
#21310000000
1!
1%
1-
12
#21320000000
0!
0%
b10 *
0-
02
b10 6
#21330000000
1!
1%
1-
12
#21340000000
0!
0%
b11 *
0-
02
b11 6
#21350000000
1!
1%
1-
12
15
#21360000000
0!
0%
b100 *
0-
02
b100 6
#21370000000
1!
1%
1-
12
#21380000000
0!
0%
b101 *
0-
02
b101 6
#21390000000
1!
1%
1-
12
#21400000000
0!
0%
b110 *
0-
02
b110 6
#21410000000
1!
1%
1-
12
#21420000000
0!
0%
b111 *
0-
02
b111 6
#21430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#21440000000
0!
0%
b0 *
0-
02
b0 6
#21450000000
1!
1%
1-
12
#21460000000
0!
0%
b1 *
0-
02
b1 6
#21470000000
1!
1%
1-
12
#21480000000
0!
0%
b10 *
0-
02
b10 6
#21490000000
1!
1%
1-
12
#21500000000
0!
0%
b11 *
0-
02
b11 6
#21510000000
1!
1%
1-
12
15
#21520000000
0!
0%
b100 *
0-
02
b100 6
#21530000000
1!
1%
1-
12
#21540000000
0!
0%
b101 *
0-
02
b101 6
#21550000000
1!
1%
1-
12
#21560000000
0!
0%
b110 *
0-
02
b110 6
#21570000000
1!
1%
1-
12
#21580000000
0!
0%
b111 *
0-
02
b111 6
#21590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#21600000000
0!
0%
b0 *
0-
02
b0 6
#21610000000
1!
1%
1-
12
#21620000000
0!
0%
b1 *
0-
02
b1 6
#21630000000
1!
1%
1-
12
#21640000000
0!
0%
b10 *
0-
02
b10 6
#21650000000
1!
1%
1-
12
#21660000000
0!
0%
b11 *
0-
02
b11 6
#21670000000
1!
1%
1-
12
15
#21680000000
0!
0%
b100 *
0-
02
b100 6
#21690000000
1!
1%
1-
12
#21700000000
0!
0%
b101 *
0-
02
b101 6
#21710000000
1!
1%
1-
12
#21720000000
0!
0%
b110 *
0-
02
b110 6
#21730000000
1!
1%
1-
12
#21740000000
0!
0%
b111 *
0-
02
b111 6
#21750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#21760000000
0!
0%
b0 *
0-
02
b0 6
#21770000000
1!
1%
1-
12
#21780000000
0!
0%
b1 *
0-
02
b1 6
#21790000000
1!
1%
1-
12
#21800000000
0!
0%
b10 *
0-
02
b10 6
#21810000000
1!
1%
1-
12
#21820000000
0!
0%
b11 *
0-
02
b11 6
#21830000000
1!
1%
1-
12
15
#21840000000
0!
0%
b100 *
0-
02
b100 6
#21850000000
1!
1%
1-
12
#21860000000
0!
0%
b101 *
0-
02
b101 6
#21870000000
1!
1%
1-
12
#21880000000
0!
0%
b110 *
0-
02
b110 6
#21890000000
1!
1%
1-
12
#21900000000
0!
0%
b111 *
0-
02
b111 6
#21910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#21920000000
0!
0%
b0 *
0-
02
b0 6
#21930000000
1!
1%
1-
12
#21940000000
0!
0%
b1 *
0-
02
b1 6
#21950000000
1!
1%
1-
12
#21960000000
0!
0%
b10 *
0-
02
b10 6
#21970000000
1!
1%
1-
12
#21980000000
0!
0%
b11 *
0-
02
b11 6
#21990000000
1!
1%
1-
12
15
#22000000000
0!
0%
b100 *
0-
02
b100 6
#22010000000
1!
1%
1-
12
#22020000000
0!
0%
b101 *
0-
02
b101 6
#22030000000
1!
1%
1-
12
#22040000000
0!
0%
b110 *
0-
02
b110 6
#22050000000
1!
1%
1-
12
#22060000000
0!
0%
b111 *
0-
02
b111 6
#22070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#22080000000
0!
0%
b0 *
0-
02
b0 6
#22090000000
1!
1%
1-
12
#22100000000
0!
0%
b1 *
0-
02
b1 6
#22110000000
1!
1%
1-
12
#22120000000
0!
0%
b10 *
0-
02
b10 6
#22130000000
1!
1%
1-
12
#22140000000
0!
0%
b11 *
0-
02
b11 6
#22150000000
1!
1%
1-
12
15
#22160000000
0!
0%
b100 *
0-
02
b100 6
#22170000000
1!
1%
1-
12
#22180000000
0!
0%
b101 *
0-
02
b101 6
#22190000000
1!
1%
1-
12
#22200000000
0!
0%
b110 *
0-
02
b110 6
#22210000000
1!
1%
1-
12
#22220000000
0!
0%
b111 *
0-
02
b111 6
#22230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#22240000000
0!
0%
b0 *
0-
02
b0 6
#22250000000
1!
1%
1-
12
#22260000000
0!
0%
b1 *
0-
02
b1 6
#22270000000
1!
1%
1-
12
#22280000000
0!
0%
b10 *
0-
02
b10 6
#22290000000
1!
1%
1-
12
#22300000000
0!
0%
b11 *
0-
02
b11 6
#22310000000
1!
1%
1-
12
15
#22320000000
0!
0%
b100 *
0-
02
b100 6
#22330000000
1!
1%
1-
12
#22340000000
0!
0%
b101 *
0-
02
b101 6
#22350000000
1!
1%
1-
12
#22360000000
0!
0%
b110 *
0-
02
b110 6
#22370000000
1!
1%
1-
12
#22380000000
0!
0%
b111 *
0-
02
b111 6
#22390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#22400000000
0!
0%
b0 *
0-
02
b0 6
#22410000000
1!
1%
1-
12
#22420000000
0!
0%
b1 *
0-
02
b1 6
#22430000000
1!
1%
1-
12
#22440000000
0!
0%
b10 *
0-
02
b10 6
#22450000000
1!
1%
1-
12
#22460000000
0!
0%
b11 *
0-
02
b11 6
#22470000000
1!
1%
1-
12
15
#22480000000
0!
0%
b100 *
0-
02
b100 6
#22490000000
1!
1%
1-
12
#22500000000
0!
0%
b101 *
0-
02
b101 6
#22510000000
1!
1%
1-
12
#22520000000
0!
0%
b110 *
0-
02
b110 6
#22530000000
1!
1%
1-
12
#22540000000
0!
0%
b111 *
0-
02
b111 6
#22550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#22560000000
0!
0%
b0 *
0-
02
b0 6
#22570000000
1!
1%
1-
12
#22580000000
0!
0%
b1 *
0-
02
b1 6
#22590000000
1!
1%
1-
12
#22600000000
0!
0%
b10 *
0-
02
b10 6
#22610000000
1!
1%
1-
12
#22620000000
0!
0%
b11 *
0-
02
b11 6
#22630000000
1!
1%
1-
12
15
#22640000000
0!
0%
b100 *
0-
02
b100 6
#22650000000
1!
1%
1-
12
#22660000000
0!
0%
b101 *
0-
02
b101 6
#22670000000
1!
1%
1-
12
#22680000000
0!
0%
b110 *
0-
02
b110 6
#22690000000
1!
1%
1-
12
#22700000000
0!
0%
b111 *
0-
02
b111 6
#22710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#22720000000
0!
0%
b0 *
0-
02
b0 6
#22730000000
1!
1%
1-
12
#22740000000
0!
0%
b1 *
0-
02
b1 6
#22750000000
1!
1%
1-
12
#22760000000
0!
0%
b10 *
0-
02
b10 6
#22770000000
1!
1%
1-
12
#22780000000
0!
0%
b11 *
0-
02
b11 6
#22790000000
1!
1%
1-
12
15
#22800000000
0!
0%
b100 *
0-
02
b100 6
#22810000000
1!
1%
1-
12
#22820000000
0!
0%
b101 *
0-
02
b101 6
#22830000000
1!
1%
1-
12
#22840000000
0!
0%
b110 *
0-
02
b110 6
#22850000000
1!
1%
1-
12
#22860000000
0!
0%
b111 *
0-
02
b111 6
#22870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#22880000000
0!
0%
b0 *
0-
02
b0 6
#22890000000
1!
1%
1-
12
#22900000000
0!
0%
b1 *
0-
02
b1 6
#22910000000
1!
1%
1-
12
#22920000000
0!
0%
b10 *
0-
02
b10 6
#22930000000
1!
1%
1-
12
#22940000000
0!
0%
b11 *
0-
02
b11 6
#22950000000
1!
1%
1-
12
15
#22960000000
0!
0%
b100 *
0-
02
b100 6
#22970000000
1!
1%
1-
12
#22980000000
0!
0%
b101 *
0-
02
b101 6
#22990000000
1!
1%
1-
12
#23000000000
0!
0%
b110 *
0-
02
b110 6
#23010000000
1!
1%
1-
12
#23020000000
0!
0%
b111 *
0-
02
b111 6
#23030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#23040000000
0!
0%
b0 *
0-
02
b0 6
#23050000000
1!
1%
1-
12
#23060000000
0!
0%
b1 *
0-
02
b1 6
#23070000000
1!
1%
1-
12
#23080000000
0!
0%
b10 *
0-
02
b10 6
#23090000000
1!
1%
1-
12
#23100000000
0!
0%
b11 *
0-
02
b11 6
#23110000000
1!
1%
1-
12
15
#23120000000
0!
0%
b100 *
0-
02
b100 6
#23130000000
1!
1%
1-
12
#23140000000
0!
0%
b101 *
0-
02
b101 6
#23150000000
1!
1%
1-
12
#23160000000
0!
0%
b110 *
0-
02
b110 6
#23170000000
1!
1%
1-
12
#23180000000
0!
0%
b111 *
0-
02
b111 6
#23190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#23200000000
0!
0%
b0 *
0-
02
b0 6
#23210000000
1!
1%
1-
12
#23220000000
0!
0%
b1 *
0-
02
b1 6
#23230000000
1!
1%
1-
12
#23240000000
0!
0%
b10 *
0-
02
b10 6
#23250000000
1!
1%
1-
12
#23260000000
0!
0%
b11 *
0-
02
b11 6
#23270000000
1!
1%
1-
12
15
#23280000000
0!
0%
b100 *
0-
02
b100 6
#23290000000
1!
1%
1-
12
#23300000000
0!
0%
b101 *
0-
02
b101 6
#23310000000
1!
1%
1-
12
#23320000000
0!
0%
b110 *
0-
02
b110 6
#23330000000
1!
1%
1-
12
#23340000000
0!
0%
b111 *
0-
02
b111 6
#23350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#23360000000
0!
0%
b0 *
0-
02
b0 6
#23370000000
1!
1%
1-
12
#23380000000
0!
0%
b1 *
0-
02
b1 6
#23390000000
1!
1%
1-
12
#23400000000
0!
0%
b10 *
0-
02
b10 6
#23410000000
1!
1%
1-
12
#23420000000
0!
0%
b11 *
0-
02
b11 6
#23430000000
1!
1%
1-
12
15
#23440000000
0!
0%
b100 *
0-
02
b100 6
#23450000000
1!
1%
1-
12
#23460000000
0!
0%
b101 *
0-
02
b101 6
#23470000000
1!
1%
1-
12
#23480000000
0!
0%
b110 *
0-
02
b110 6
#23490000000
1!
1%
1-
12
#23500000000
0!
0%
b111 *
0-
02
b111 6
#23510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#23520000000
0!
0%
b0 *
0-
02
b0 6
#23530000000
1!
1%
1-
12
#23540000000
0!
0%
b1 *
0-
02
b1 6
#23550000000
1!
1%
1-
12
#23560000000
0!
0%
b10 *
0-
02
b10 6
#23570000000
1!
1%
1-
12
#23580000000
0!
0%
b11 *
0-
02
b11 6
#23590000000
1!
1%
1-
12
15
#23600000000
0!
0%
b100 *
0-
02
b100 6
#23610000000
1!
1%
1-
12
#23620000000
0!
0%
b101 *
0-
02
b101 6
#23630000000
1!
1%
1-
12
#23640000000
0!
0%
b110 *
0-
02
b110 6
#23650000000
1!
1%
1-
12
#23660000000
0!
0%
b111 *
0-
02
b111 6
#23670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#23680000000
0!
0%
b0 *
0-
02
b0 6
#23690000000
1!
1%
1-
12
#23700000000
0!
0%
b1 *
0-
02
b1 6
#23710000000
1!
1%
1-
12
#23720000000
0!
0%
b10 *
0-
02
b10 6
#23730000000
1!
1%
1-
12
#23740000000
0!
0%
b11 *
0-
02
b11 6
#23750000000
1!
1%
1-
12
15
#23760000000
0!
0%
b100 *
0-
02
b100 6
#23770000000
1!
1%
1-
12
#23780000000
0!
0%
b101 *
0-
02
b101 6
#23790000000
1!
1%
1-
12
#23800000000
0!
0%
b110 *
0-
02
b110 6
#23810000000
1!
1%
1-
12
#23820000000
0!
0%
b111 *
0-
02
b111 6
#23830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#23840000000
0!
0%
b0 *
0-
02
b0 6
#23850000000
1!
1%
1-
12
#23860000000
0!
0%
b1 *
0-
02
b1 6
#23870000000
1!
1%
1-
12
#23880000000
0!
0%
b10 *
0-
02
b10 6
#23890000000
1!
1%
1-
12
#23900000000
0!
0%
b11 *
0-
02
b11 6
#23910000000
1!
1%
1-
12
15
#23920000000
0!
0%
b100 *
0-
02
b100 6
#23930000000
1!
1%
1-
12
#23940000000
0!
0%
b101 *
0-
02
b101 6
#23950000000
1!
1%
1-
12
#23960000000
0!
0%
b110 *
0-
02
b110 6
#23970000000
1!
1%
1-
12
#23980000000
0!
0%
b111 *
0-
02
b111 6
#23990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#24000000000
0!
0%
b0 *
0-
02
b0 6
#24010000000
1!
1%
1-
12
#24020000000
0!
0%
b1 *
0-
02
b1 6
#24030000000
1!
1%
1-
12
#24040000000
0!
0%
b10 *
0-
02
b10 6
#24050000000
1!
1%
1-
12
#24060000000
0!
0%
b11 *
0-
02
b11 6
#24070000000
1!
1%
1-
12
15
#24080000000
0!
0%
b100 *
0-
02
b100 6
#24090000000
1!
1%
1-
12
#24100000000
0!
0%
b101 *
0-
02
b101 6
#24110000000
1!
1%
1-
12
#24120000000
0!
0%
b110 *
0-
02
b110 6
#24130000000
1!
1%
1-
12
#24140000000
0!
0%
b111 *
0-
02
b111 6
#24150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#24160000000
0!
0%
b0 *
0-
02
b0 6
#24170000000
1!
1%
1-
12
#24180000000
0!
0%
b1 *
0-
02
b1 6
#24190000000
1!
1%
1-
12
#24200000000
0!
0%
b10 *
0-
02
b10 6
#24210000000
1!
1%
1-
12
#24220000000
0!
0%
b11 *
0-
02
b11 6
#24230000000
1!
1%
1-
12
15
#24240000000
0!
0%
b100 *
0-
02
b100 6
#24250000000
1!
1%
1-
12
#24260000000
0!
0%
b101 *
0-
02
b101 6
#24270000000
1!
1%
1-
12
#24280000000
0!
0%
b110 *
0-
02
b110 6
#24290000000
1!
1%
1-
12
#24300000000
0!
0%
b111 *
0-
02
b111 6
#24310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#24320000000
0!
0%
b0 *
0-
02
b0 6
#24330000000
1!
1%
1-
12
#24340000000
0!
0%
b1 *
0-
02
b1 6
#24350000000
1!
1%
1-
12
#24360000000
0!
0%
b10 *
0-
02
b10 6
#24370000000
1!
1%
1-
12
#24380000000
0!
0%
b11 *
0-
02
b11 6
#24390000000
1!
1%
1-
12
15
#24400000000
0!
0%
b100 *
0-
02
b100 6
#24410000000
1!
1%
1-
12
#24420000000
0!
0%
b101 *
0-
02
b101 6
#24430000000
1!
1%
1-
12
#24440000000
0!
0%
b110 *
0-
02
b110 6
#24450000000
1!
1%
1-
12
#24460000000
0!
0%
b111 *
0-
02
b111 6
#24470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#24480000000
0!
0%
b0 *
0-
02
b0 6
#24490000000
1!
1%
1-
12
#24500000000
0!
0%
b1 *
0-
02
b1 6
#24510000000
1!
1%
1-
12
#24520000000
0!
0%
b10 *
0-
02
b10 6
#24530000000
1!
1%
1-
12
#24540000000
0!
0%
b11 *
0-
02
b11 6
#24550000000
1!
1%
1-
12
15
#24560000000
0!
0%
b100 *
0-
02
b100 6
#24570000000
1!
1%
1-
12
#24580000000
0!
0%
b101 *
0-
02
b101 6
#24590000000
1!
1%
1-
12
#24600000000
0!
0%
b110 *
0-
02
b110 6
#24610000000
1!
1%
1-
12
#24620000000
0!
0%
b111 *
0-
02
b111 6
#24630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#24640000000
0!
0%
b0 *
0-
02
b0 6
#24650000000
1!
1%
1-
12
#24660000000
0!
0%
b1 *
0-
02
b1 6
#24670000000
1!
1%
1-
12
#24680000000
0!
0%
b10 *
0-
02
b10 6
#24690000000
1!
1%
1-
12
#24700000000
0!
0%
b11 *
0-
02
b11 6
#24710000000
1!
1%
1-
12
15
#24720000000
0!
0%
b100 *
0-
02
b100 6
#24730000000
1!
1%
1-
12
#24740000000
0!
0%
b101 *
0-
02
b101 6
#24750000000
1!
1%
1-
12
#24760000000
0!
0%
b110 *
0-
02
b110 6
#24770000000
1!
1%
1-
12
#24780000000
0!
0%
b111 *
0-
02
b111 6
#24790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#24800000000
0!
0%
b0 *
0-
02
b0 6
#24810000000
1!
1%
1-
12
#24820000000
0!
0%
b1 *
0-
02
b1 6
#24830000000
1!
1%
1-
12
#24840000000
0!
0%
b10 *
0-
02
b10 6
#24850000000
1!
1%
1-
12
#24860000000
0!
0%
b11 *
0-
02
b11 6
#24870000000
1!
1%
1-
12
15
#24880000000
0!
0%
b100 *
0-
02
b100 6
#24890000000
1!
1%
1-
12
#24900000000
0!
0%
b101 *
0-
02
b101 6
#24910000000
1!
1%
1-
12
#24920000000
0!
0%
b110 *
0-
02
b110 6
#24930000000
1!
1%
1-
12
#24940000000
0!
0%
b111 *
0-
02
b111 6
#24950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#24960000000
0!
0%
b0 *
0-
02
b0 6
#24970000000
1!
1%
1-
12
#24980000000
0!
0%
b1 *
0-
02
b1 6
#24990000000
1!
1%
1-
12
#25000000000
0!
0%
b10 *
0-
02
b10 6
#25010000000
1!
1%
1-
12
#25020000000
0!
0%
b11 *
0-
02
b11 6
#25030000000
1!
1%
1-
12
15
#25040000000
0!
0%
b100 *
0-
02
b100 6
#25050000000
1!
1%
1-
12
#25060000000
0!
0%
b101 *
0-
02
b101 6
#25070000000
1!
1%
1-
12
#25080000000
0!
0%
b110 *
0-
02
b110 6
#25090000000
1!
1%
1-
12
#25100000000
0!
0%
b111 *
0-
02
b111 6
#25110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#25120000000
0!
0%
b0 *
0-
02
b0 6
#25130000000
1!
1%
1-
12
#25140000000
0!
0%
b1 *
0-
02
b1 6
#25150000000
1!
1%
1-
12
#25160000000
0!
0%
b10 *
0-
02
b10 6
#25170000000
1!
1%
1-
12
#25180000000
0!
0%
b11 *
0-
02
b11 6
#25190000000
1!
1%
1-
12
15
#25200000000
0!
0%
b100 *
0-
02
b100 6
#25210000000
1!
1%
1-
12
#25220000000
0!
0%
b101 *
0-
02
b101 6
#25230000000
1!
1%
1-
12
#25240000000
0!
0%
b110 *
0-
02
b110 6
#25250000000
1!
1%
1-
12
#25260000000
0!
0%
b111 *
0-
02
b111 6
#25270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#25280000000
0!
0%
b0 *
0-
02
b0 6
#25290000000
1!
1%
1-
12
#25300000000
0!
0%
b1 *
0-
02
b1 6
#25310000000
1!
1%
1-
12
#25320000000
0!
0%
b10 *
0-
02
b10 6
#25330000000
1!
1%
1-
12
#25340000000
0!
0%
b11 *
0-
02
b11 6
#25350000000
1!
1%
1-
12
15
#25360000000
0!
0%
b100 *
0-
02
b100 6
#25370000000
1!
1%
1-
12
#25380000000
0!
0%
b101 *
0-
02
b101 6
#25390000000
1!
1%
1-
12
#25400000000
0!
0%
b110 *
0-
02
b110 6
#25410000000
1!
1%
1-
12
#25420000000
0!
0%
b111 *
0-
02
b111 6
#25430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#25440000000
0!
0%
b0 *
0-
02
b0 6
#25450000000
1!
1%
1-
12
#25460000000
0!
0%
b1 *
0-
02
b1 6
#25470000000
1!
1%
1-
12
#25480000000
0!
0%
b10 *
0-
02
b10 6
#25490000000
1!
1%
1-
12
#25500000000
0!
0%
b11 *
0-
02
b11 6
#25510000000
1!
1%
1-
12
15
#25520000000
0!
0%
b100 *
0-
02
b100 6
#25530000000
1!
1%
1-
12
#25540000000
0!
0%
b101 *
0-
02
b101 6
#25550000000
1!
1%
1-
12
#25560000000
0!
0%
b110 *
0-
02
b110 6
#25570000000
1!
1%
1-
12
#25580000000
0!
0%
b111 *
0-
02
b111 6
#25590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#25600000000
0!
0%
b0 *
0-
02
b0 6
#25610000000
1!
1%
1-
12
#25620000000
0!
0%
b1 *
0-
02
b1 6
#25630000000
1!
1%
1-
12
#25640000000
0!
0%
b10 *
0-
02
b10 6
#25650000000
1!
1%
1-
12
#25660000000
0!
0%
b11 *
0-
02
b11 6
#25670000000
1!
1%
1-
12
15
#25680000000
0!
0%
b100 *
0-
02
b100 6
#25690000000
1!
1%
1-
12
#25700000000
0!
0%
b101 *
0-
02
b101 6
#25710000000
1!
1%
1-
12
#25720000000
0!
0%
b110 *
0-
02
b110 6
#25730000000
1!
1%
1-
12
#25740000000
0!
0%
b111 *
0-
02
b111 6
#25750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#25760000000
0!
0%
b0 *
0-
02
b0 6
#25770000000
1!
1%
1-
12
#25780000000
0!
0%
b1 *
0-
02
b1 6
#25790000000
1!
1%
1-
12
#25800000000
0!
0%
b10 *
0-
02
b10 6
#25810000000
1!
1%
1-
12
#25820000000
0!
0%
b11 *
0-
02
b11 6
#25830000000
1!
1%
1-
12
15
#25840000000
0!
0%
b100 *
0-
02
b100 6
#25850000000
1!
1%
1-
12
#25860000000
0!
0%
b101 *
0-
02
b101 6
#25870000000
1!
1%
1-
12
#25880000000
0!
0%
b110 *
0-
02
b110 6
#25890000000
1!
1%
1-
12
#25900000000
0!
0%
b111 *
0-
02
b111 6
#25910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#25920000000
0!
0%
b0 *
0-
02
b0 6
#25930000000
1!
1%
1-
12
#25940000000
0!
0%
b1 *
0-
02
b1 6
#25950000000
1!
1%
1-
12
#25960000000
0!
0%
b10 *
0-
02
b10 6
#25970000000
1!
1%
1-
12
#25980000000
0!
0%
b11 *
0-
02
b11 6
#25990000000
1!
1%
1-
12
15
#26000000000
0!
0%
b100 *
0-
02
b100 6
#26010000000
1!
1%
1-
12
#26020000000
0!
0%
b101 *
0-
02
b101 6
#26030000000
1!
1%
1-
12
#26040000000
0!
0%
b110 *
0-
02
b110 6
#26050000000
1!
1%
1-
12
#26060000000
0!
0%
b111 *
0-
02
b111 6
#26070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#26080000000
0!
0%
b0 *
0-
02
b0 6
#26090000000
1!
1%
1-
12
#26100000000
0!
0%
b1 *
0-
02
b1 6
#26110000000
1!
1%
1-
12
#26120000000
0!
0%
b10 *
0-
02
b10 6
#26130000000
1!
1%
1-
12
#26140000000
0!
0%
b11 *
0-
02
b11 6
#26150000000
1!
1%
1-
12
15
#26160000000
0!
0%
b100 *
0-
02
b100 6
#26170000000
1!
1%
1-
12
#26180000000
0!
0%
b101 *
0-
02
b101 6
#26190000000
1!
1%
1-
12
#26200000000
0!
0%
b110 *
0-
02
b110 6
#26210000000
1!
1%
1-
12
#26220000000
0!
0%
b111 *
0-
02
b111 6
#26230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#26240000000
0!
0%
b0 *
0-
02
b0 6
#26250000000
1!
1%
1-
12
#26260000000
0!
0%
b1 *
0-
02
b1 6
#26270000000
1!
1%
1-
12
#26280000000
0!
0%
b10 *
0-
02
b10 6
#26290000000
1!
1%
1-
12
#26300000000
0!
0%
b11 *
0-
02
b11 6
#26310000000
1!
1%
1-
12
15
#26320000000
0!
0%
b100 *
0-
02
b100 6
#26330000000
1!
1%
1-
12
#26340000000
0!
0%
b101 *
0-
02
b101 6
#26350000000
1!
1%
1-
12
#26360000000
0!
0%
b110 *
0-
02
b110 6
#26370000000
1!
1%
1-
12
#26380000000
0!
0%
b111 *
0-
02
b111 6
#26390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#26400000000
0!
0%
b0 *
0-
02
b0 6
#26410000000
1!
1%
1-
12
#26420000000
0!
0%
b1 *
0-
02
b1 6
#26430000000
1!
1%
1-
12
#26440000000
0!
0%
b10 *
0-
02
b10 6
#26450000000
1!
1%
1-
12
#26460000000
0!
0%
b11 *
0-
02
b11 6
#26470000000
1!
1%
1-
12
15
#26480000000
0!
0%
b100 *
0-
02
b100 6
#26490000000
1!
1%
1-
12
#26500000000
0!
0%
b101 *
0-
02
b101 6
#26510000000
1!
1%
1-
12
#26520000000
0!
0%
b110 *
0-
02
b110 6
#26530000000
1!
1%
1-
12
#26540000000
0!
0%
b111 *
0-
02
b111 6
#26550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#26560000000
0!
0%
b0 *
0-
02
b0 6
#26570000000
1!
1%
1-
12
#26580000000
0!
0%
b1 *
0-
02
b1 6
#26590000000
1!
1%
1-
12
#26600000000
0!
0%
b10 *
0-
02
b10 6
#26610000000
1!
1%
1-
12
#26620000000
0!
0%
b11 *
0-
02
b11 6
#26630000000
1!
1%
1-
12
15
#26640000000
0!
0%
b100 *
0-
02
b100 6
#26650000000
1!
1%
1-
12
#26660000000
0!
0%
b101 *
0-
02
b101 6
#26670000000
1!
1%
1-
12
#26680000000
0!
0%
b110 *
0-
02
b110 6
#26690000000
1!
1%
1-
12
#26700000000
0!
0%
b111 *
0-
02
b111 6
#26710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#26720000000
0!
0%
b0 *
0-
02
b0 6
#26730000000
1!
1%
1-
12
#26740000000
0!
0%
b1 *
0-
02
b1 6
#26750000000
1!
1%
1-
12
#26760000000
0!
0%
b10 *
0-
02
b10 6
#26770000000
1!
1%
1-
12
#26780000000
0!
0%
b11 *
0-
02
b11 6
#26790000000
1!
1%
1-
12
15
#26800000000
0!
0%
b100 *
0-
02
b100 6
#26810000000
1!
1%
1-
12
#26820000000
0!
0%
b101 *
0-
02
b101 6
#26830000000
1!
1%
1-
12
#26840000000
0!
0%
b110 *
0-
02
b110 6
#26850000000
1!
1%
1-
12
#26860000000
0!
0%
b111 *
0-
02
b111 6
#26870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#26880000000
0!
0%
b0 *
0-
02
b0 6
#26890000000
1!
1%
1-
12
#26900000000
0!
0%
b1 *
0-
02
b1 6
#26910000000
1!
1%
1-
12
#26920000000
0!
0%
b10 *
0-
02
b10 6
#26930000000
1!
1%
1-
12
#26940000000
0!
0%
b11 *
0-
02
b11 6
#26950000000
1!
1%
1-
12
15
#26960000000
0!
0%
b100 *
0-
02
b100 6
#26970000000
1!
1%
1-
12
#26980000000
0!
0%
b101 *
0-
02
b101 6
#26990000000
1!
1%
1-
12
#27000000000
0!
0%
b110 *
0-
02
b110 6
#27010000000
1!
1%
1-
12
#27020000000
0!
0%
b111 *
0-
02
b111 6
#27030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#27040000000
0!
0%
b0 *
0-
02
b0 6
#27050000000
1!
1%
1-
12
#27060000000
0!
0%
b1 *
0-
02
b1 6
#27070000000
1!
1%
1-
12
#27080000000
0!
0%
b10 *
0-
02
b10 6
#27090000000
1!
1%
1-
12
#27100000000
0!
0%
b11 *
0-
02
b11 6
#27110000000
1!
1%
1-
12
15
#27120000000
0!
0%
b100 *
0-
02
b100 6
#27130000000
1!
1%
1-
12
#27140000000
0!
0%
b101 *
0-
02
b101 6
#27150000000
1!
1%
1-
12
#27160000000
0!
0%
b110 *
0-
02
b110 6
#27170000000
1!
1%
1-
12
#27180000000
0!
0%
b111 *
0-
02
b111 6
#27190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#27200000000
0!
0%
b0 *
0-
02
b0 6
#27210000000
1!
1%
1-
12
#27220000000
0!
0%
b1 *
0-
02
b1 6
#27230000000
1!
1%
1-
12
#27240000000
0!
0%
b10 *
0-
02
b10 6
#27250000000
1!
1%
1-
12
#27260000000
0!
0%
b11 *
0-
02
b11 6
#27270000000
1!
1%
1-
12
15
#27280000000
0!
0%
b100 *
0-
02
b100 6
#27290000000
1!
1%
1-
12
#27300000000
0!
0%
b101 *
0-
02
b101 6
#27310000000
1!
1%
1-
12
#27320000000
0!
0%
b110 *
0-
02
b110 6
#27330000000
1!
1%
1-
12
#27340000000
0!
0%
b111 *
0-
02
b111 6
#27350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#27360000000
0!
0%
b0 *
0-
02
b0 6
#27370000000
1!
1%
1-
12
#27380000000
0!
0%
b1 *
0-
02
b1 6
#27390000000
1!
1%
1-
12
#27400000000
0!
0%
b10 *
0-
02
b10 6
#27410000000
1!
1%
1-
12
#27420000000
0!
0%
b11 *
0-
02
b11 6
#27430000000
1!
1%
1-
12
15
#27440000000
0!
0%
b100 *
0-
02
b100 6
#27450000000
1!
1%
1-
12
#27460000000
0!
0%
b101 *
0-
02
b101 6
#27470000000
1!
1%
1-
12
#27480000000
0!
0%
b110 *
0-
02
b110 6
#27490000000
1!
1%
1-
12
#27500000000
0!
0%
b111 *
0-
02
b111 6
#27510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#27520000000
0!
0%
b0 *
0-
02
b0 6
#27530000000
1!
1%
1-
12
#27540000000
0!
0%
b1 *
0-
02
b1 6
#27550000000
1!
1%
1-
12
#27560000000
0!
0%
b10 *
0-
02
b10 6
#27570000000
1!
1%
1-
12
#27580000000
0!
0%
b11 *
0-
02
b11 6
#27590000000
1!
1%
1-
12
15
#27600000000
0!
0%
b100 *
0-
02
b100 6
#27610000000
1!
1%
1-
12
#27620000000
0!
0%
b101 *
0-
02
b101 6
#27630000000
1!
1%
1-
12
#27640000000
0!
0%
b110 *
0-
02
b110 6
#27650000000
1!
1%
1-
12
#27660000000
0!
0%
b111 *
0-
02
b111 6
#27670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#27680000000
0!
0%
b0 *
0-
02
b0 6
#27690000000
1!
1%
1-
12
#27700000000
0!
0%
b1 *
0-
02
b1 6
#27710000000
1!
1%
1-
12
#27720000000
0!
0%
b10 *
0-
02
b10 6
#27730000000
1!
1%
1-
12
#27740000000
0!
0%
b11 *
0-
02
b11 6
#27750000000
1!
1%
1-
12
15
#27760000000
0!
0%
b100 *
0-
02
b100 6
#27770000000
1!
1%
1-
12
#27780000000
0!
0%
b101 *
0-
02
b101 6
#27790000000
1!
1%
1-
12
#27800000000
0!
0%
b110 *
0-
02
b110 6
#27810000000
1!
1%
1-
12
#27820000000
0!
0%
b111 *
0-
02
b111 6
#27830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#27840000000
0!
0%
b0 *
0-
02
b0 6
#27850000000
1!
1%
1-
12
#27860000000
0!
0%
b1 *
0-
02
b1 6
#27870000000
1!
1%
1-
12
#27880000000
0!
0%
b10 *
0-
02
b10 6
#27890000000
1!
1%
1-
12
#27900000000
0!
0%
b11 *
0-
02
b11 6
#27910000000
1!
1%
1-
12
15
#27920000000
0!
0%
b100 *
0-
02
b100 6
#27930000000
1!
1%
1-
12
#27940000000
0!
0%
b101 *
0-
02
b101 6
#27950000000
1!
1%
1-
12
#27960000000
0!
0%
b110 *
0-
02
b110 6
#27970000000
1!
1%
1-
12
#27980000000
0!
0%
b111 *
0-
02
b111 6
#27990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#28000000000
0!
0%
b0 *
0-
02
b0 6
#28010000000
1!
1%
1-
12
#28020000000
0!
0%
b1 *
0-
02
b1 6
#28030000000
1!
1%
1-
12
#28040000000
0!
0%
b10 *
0-
02
b10 6
#28050000000
1!
1%
1-
12
#28060000000
0!
0%
b11 *
0-
02
b11 6
#28070000000
1!
1%
1-
12
15
#28080000000
0!
0%
b100 *
0-
02
b100 6
#28090000000
1!
1%
1-
12
#28100000000
0!
0%
b101 *
0-
02
b101 6
#28110000000
1!
1%
1-
12
#28120000000
0!
0%
b110 *
0-
02
b110 6
#28130000000
1!
1%
1-
12
#28140000000
0!
0%
b111 *
0-
02
b111 6
#28150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#28160000000
0!
0%
b0 *
0-
02
b0 6
#28170000000
1!
1%
1-
12
#28180000000
0!
0%
b1 *
0-
02
b1 6
#28190000000
1!
1%
1-
12
#28200000000
0!
0%
b10 *
0-
02
b10 6
#28210000000
1!
1%
1-
12
#28220000000
0!
0%
b11 *
0-
02
b11 6
#28230000000
1!
1%
1-
12
15
#28240000000
0!
0%
b100 *
0-
02
b100 6
#28250000000
1!
1%
1-
12
#28260000000
0!
0%
b101 *
0-
02
b101 6
#28270000000
1!
1%
1-
12
#28280000000
0!
0%
b110 *
0-
02
b110 6
#28290000000
1!
1%
1-
12
#28300000000
0!
0%
b111 *
0-
02
b111 6
#28310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#28320000000
0!
0%
b0 *
0-
02
b0 6
#28330000000
1!
1%
1-
12
#28340000000
0!
0%
b1 *
0-
02
b1 6
#28350000000
1!
1%
1-
12
#28360000000
0!
0%
b10 *
0-
02
b10 6
#28370000000
1!
1%
1-
12
#28380000000
0!
0%
b11 *
0-
02
b11 6
#28390000000
1!
1%
1-
12
15
#28400000000
0!
0%
b100 *
0-
02
b100 6
#28410000000
1!
1%
1-
12
#28420000000
0!
0%
b101 *
0-
02
b101 6
#28430000000
1!
1%
1-
12
#28440000000
0!
0%
b110 *
0-
02
b110 6
#28450000000
1!
1%
1-
12
#28460000000
0!
0%
b111 *
0-
02
b111 6
#28470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#28480000000
0!
0%
b0 *
0-
02
b0 6
#28490000000
1!
1%
1-
12
#28500000000
0!
0%
b1 *
0-
02
b1 6
#28510000000
1!
1%
1-
12
#28520000000
0!
0%
b10 *
0-
02
b10 6
#28530000000
1!
1%
1-
12
#28540000000
0!
0%
b11 *
0-
02
b11 6
#28550000000
1!
1%
1-
12
15
#28560000000
0!
0%
b100 *
0-
02
b100 6
#28570000000
1!
1%
1-
12
#28580000000
0!
0%
b101 *
0-
02
b101 6
#28590000000
1!
1%
1-
12
#28600000000
0!
0%
b110 *
0-
02
b110 6
#28610000000
1!
1%
1-
12
#28620000000
0!
0%
b111 *
0-
02
b111 6
#28630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#28640000000
0!
0%
b0 *
0-
02
b0 6
#28650000000
1!
1%
1-
12
#28660000000
0!
0%
b1 *
0-
02
b1 6
#28670000000
1!
1%
1-
12
#28680000000
0!
0%
b10 *
0-
02
b10 6
#28690000000
1!
1%
1-
12
#28700000000
0!
0%
b11 *
0-
02
b11 6
#28710000000
1!
1%
1-
12
15
#28720000000
0!
0%
b100 *
0-
02
b100 6
#28730000000
1!
1%
1-
12
#28740000000
0!
0%
b101 *
0-
02
b101 6
#28750000000
1!
1%
1-
12
#28760000000
0!
0%
b110 *
0-
02
b110 6
#28770000000
1!
1%
1-
12
#28780000000
0!
0%
b111 *
0-
02
b111 6
#28790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#28800000000
0!
0%
b0 *
0-
02
b0 6
#28810000000
1!
1%
1-
12
#28820000000
0!
0%
b1 *
0-
02
b1 6
#28830000000
1!
1%
1-
12
#28840000000
0!
0%
b10 *
0-
02
b10 6
#28850000000
1!
1%
1-
12
#28860000000
0!
0%
b11 *
0-
02
b11 6
#28870000000
1!
1%
1-
12
15
#28880000000
0!
0%
b100 *
0-
02
b100 6
#28890000000
1!
1%
1-
12
#28900000000
0!
0%
b101 *
0-
02
b101 6
#28910000000
1!
1%
1-
12
#28920000000
0!
0%
b110 *
0-
02
b110 6
#28930000000
1!
1%
1-
12
#28940000000
0!
0%
b111 *
0-
02
b111 6
#28950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#28960000000
0!
0%
b0 *
0-
02
b0 6
#28970000000
1!
1%
1-
12
#28980000000
0!
0%
b1 *
0-
02
b1 6
#28990000000
1!
1%
1-
12
#29000000000
0!
0%
b10 *
0-
02
b10 6
#29010000000
1!
1%
1-
12
#29020000000
0!
0%
b11 *
0-
02
b11 6
#29030000000
1!
1%
1-
12
15
#29040000000
0!
0%
b100 *
0-
02
b100 6
#29050000000
1!
1%
1-
12
#29060000000
0!
0%
b101 *
0-
02
b101 6
#29070000000
1!
1%
1-
12
#29080000000
0!
0%
b110 *
0-
02
b110 6
#29090000000
1!
1%
1-
12
#29100000000
0!
0%
b111 *
0-
02
b111 6
#29110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#29120000000
0!
0%
b0 *
0-
02
b0 6
#29130000000
1!
1%
1-
12
#29140000000
0!
0%
b1 *
0-
02
b1 6
#29150000000
1!
1%
1-
12
#29160000000
0!
0%
b10 *
0-
02
b10 6
#29170000000
1!
1%
1-
12
#29180000000
0!
0%
b11 *
0-
02
b11 6
#29190000000
1!
1%
1-
12
15
#29200000000
0!
0%
b100 *
0-
02
b100 6
#29210000000
1!
1%
1-
12
#29220000000
0!
0%
b101 *
0-
02
b101 6
#29230000000
1!
1%
1-
12
#29240000000
0!
0%
b110 *
0-
02
b110 6
#29250000000
1!
1%
1-
12
#29260000000
0!
0%
b111 *
0-
02
b111 6
#29270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#29280000000
0!
0%
b0 *
0-
02
b0 6
#29290000000
1!
1%
1-
12
#29300000000
0!
0%
b1 *
0-
02
b1 6
#29310000000
1!
1%
1-
12
#29320000000
0!
0%
b10 *
0-
02
b10 6
#29330000000
1!
1%
1-
12
#29340000000
0!
0%
b11 *
0-
02
b11 6
#29350000000
1!
1%
1-
12
15
#29360000000
0!
0%
b100 *
0-
02
b100 6
#29370000000
1!
1%
1-
12
#29380000000
0!
0%
b101 *
0-
02
b101 6
#29390000000
1!
1%
1-
12
#29400000000
0!
0%
b110 *
0-
02
b110 6
#29410000000
1!
1%
1-
12
#29420000000
0!
0%
b111 *
0-
02
b111 6
#29430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#29440000000
0!
0%
b0 *
0-
02
b0 6
#29450000000
1!
1%
1-
12
#29460000000
0!
0%
b1 *
0-
02
b1 6
#29470000000
1!
1%
1-
12
#29480000000
0!
0%
b10 *
0-
02
b10 6
#29490000000
1!
1%
1-
12
#29500000000
0!
0%
b11 *
0-
02
b11 6
#29510000000
1!
1%
1-
12
15
#29520000000
0!
0%
b100 *
0-
02
b100 6
#29530000000
1!
1%
1-
12
#29540000000
0!
0%
b101 *
0-
02
b101 6
#29550000000
1!
1%
1-
12
#29560000000
0!
0%
b110 *
0-
02
b110 6
#29570000000
1!
1%
1-
12
#29580000000
0!
0%
b111 *
0-
02
b111 6
#29590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#29600000000
0!
0%
b0 *
0-
02
b0 6
#29610000000
1!
1%
1-
12
#29620000000
0!
0%
b1 *
0-
02
b1 6
#29630000000
1!
1%
1-
12
#29640000000
0!
0%
b10 *
0-
02
b10 6
#29650000000
1!
1%
1-
12
#29660000000
0!
0%
b11 *
0-
02
b11 6
#29670000000
1!
1%
1-
12
15
#29680000000
0!
0%
b100 *
0-
02
b100 6
#29690000000
1!
1%
1-
12
#29700000000
0!
0%
b101 *
0-
02
b101 6
#29710000000
1!
1%
1-
12
#29720000000
0!
0%
b110 *
0-
02
b110 6
#29730000000
1!
1%
1-
12
#29740000000
0!
0%
b111 *
0-
02
b111 6
#29750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#29760000000
0!
0%
b0 *
0-
02
b0 6
#29770000000
1!
1%
1-
12
#29780000000
0!
0%
b1 *
0-
02
b1 6
#29790000000
1!
1%
1-
12
#29800000000
0!
0%
b10 *
0-
02
b10 6
#29810000000
1!
1%
1-
12
#29820000000
0!
0%
b11 *
0-
02
b11 6
#29830000000
1!
1%
1-
12
15
#29840000000
0!
0%
b100 *
0-
02
b100 6
#29850000000
1!
1%
1-
12
#29860000000
0!
0%
b101 *
0-
02
b101 6
#29870000000
1!
1%
1-
12
#29880000000
0!
0%
b110 *
0-
02
b110 6
#29890000000
1!
1%
1-
12
#29900000000
0!
0%
b111 *
0-
02
b111 6
#29910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#29920000000
0!
0%
b0 *
0-
02
b0 6
#29930000000
1!
1%
1-
12
#29940000000
0!
0%
b1 *
0-
02
b1 6
#29950000000
1!
1%
1-
12
#29960000000
0!
0%
b10 *
0-
02
b10 6
#29970000000
1!
1%
1-
12
#29980000000
0!
0%
b11 *
0-
02
b11 6
#29990000000
1!
1%
1-
12
15
#30000000000
0!
0%
b100 *
0-
02
b100 6
#30010000000
1!
1%
1-
12
#30020000000
0!
0%
b101 *
0-
02
b101 6
#30030000000
1!
1%
1-
12
#30040000000
0!
0%
b110 *
0-
02
b110 6
#30050000000
1!
1%
1-
12
#30060000000
0!
0%
b111 *
0-
02
b111 6
#30070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#30080000000
0!
0%
b0 *
0-
02
b0 6
#30090000000
1!
1%
1-
12
#30100000000
0!
0%
b1 *
0-
02
b1 6
#30110000000
1!
1%
1-
12
#30120000000
0!
0%
b10 *
0-
02
b10 6
#30130000000
1!
1%
1-
12
#30140000000
0!
0%
b11 *
0-
02
b11 6
#30150000000
1!
1%
1-
12
15
#30160000000
0!
0%
b100 *
0-
02
b100 6
#30170000000
1!
1%
1-
12
#30180000000
0!
0%
b101 *
0-
02
b101 6
#30190000000
1!
1%
1-
12
#30200000000
0!
0%
b110 *
0-
02
b110 6
#30210000000
1!
1%
1-
12
#30220000000
0!
0%
b111 *
0-
02
b111 6
#30230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#30240000000
0!
0%
b0 *
0-
02
b0 6
#30250000000
1!
1%
1-
12
#30260000000
0!
0%
b1 *
0-
02
b1 6
#30270000000
1!
1%
1-
12
#30280000000
0!
0%
b10 *
0-
02
b10 6
#30290000000
1!
1%
1-
12
#30300000000
0!
0%
b11 *
0-
02
b11 6
#30310000000
1!
1%
1-
12
15
#30320000000
0!
0%
b100 *
0-
02
b100 6
#30330000000
1!
1%
1-
12
#30340000000
0!
0%
b101 *
0-
02
b101 6
#30350000000
1!
1%
1-
12
#30360000000
0!
0%
b110 *
0-
02
b110 6
#30370000000
1!
1%
1-
12
#30380000000
0!
0%
b111 *
0-
02
b111 6
#30390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#30400000000
0!
0%
b0 *
0-
02
b0 6
#30410000000
1!
1%
1-
12
#30420000000
0!
0%
b1 *
0-
02
b1 6
#30430000000
1!
1%
1-
12
#30440000000
0!
0%
b10 *
0-
02
b10 6
#30450000000
1!
1%
1-
12
#30460000000
0!
0%
b11 *
0-
02
b11 6
#30470000000
1!
1%
1-
12
15
#30480000000
0!
0%
b100 *
0-
02
b100 6
#30490000000
1!
1%
1-
12
#30500000000
0!
0%
b101 *
0-
02
b101 6
#30510000000
1!
1%
1-
12
#30520000000
0!
0%
b110 *
0-
02
b110 6
#30530000000
1!
1%
1-
12
#30540000000
0!
0%
b111 *
0-
02
b111 6
#30550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#30560000000
0!
0%
b0 *
0-
02
b0 6
#30570000000
1!
1%
1-
12
#30580000000
0!
0%
b1 *
0-
02
b1 6
#30590000000
1!
1%
1-
12
#30600000000
0!
0%
b10 *
0-
02
b10 6
#30610000000
1!
1%
1-
12
#30620000000
0!
0%
b11 *
0-
02
b11 6
#30630000000
1!
1%
1-
12
15
#30640000000
0!
0%
b100 *
0-
02
b100 6
#30650000000
1!
1%
1-
12
#30660000000
0!
0%
b101 *
0-
02
b101 6
#30670000000
1!
1%
1-
12
#30680000000
0!
0%
b110 *
0-
02
b110 6
#30690000000
1!
1%
1-
12
#30700000000
0!
0%
b111 *
0-
02
b111 6
#30710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#30720000000
0!
0%
b0 *
0-
02
b0 6
#30730000000
1!
1%
1-
12
#30740000000
0!
0%
b1 *
0-
02
b1 6
#30750000000
1!
1%
1-
12
#30760000000
0!
0%
b10 *
0-
02
b10 6
#30770000000
1!
1%
1-
12
#30780000000
0!
0%
b11 *
0-
02
b11 6
#30790000000
1!
1%
1-
12
15
#30800000000
0!
0%
b100 *
0-
02
b100 6
#30810000000
1!
1%
1-
12
#30820000000
0!
0%
b101 *
0-
02
b101 6
#30830000000
1!
1%
1-
12
#30840000000
0!
0%
b110 *
0-
02
b110 6
#30850000000
1!
1%
1-
12
#30860000000
0!
0%
b111 *
0-
02
b111 6
#30870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#30880000000
0!
0%
b0 *
0-
02
b0 6
#30890000000
1!
1%
1-
12
#30900000000
0!
0%
b1 *
0-
02
b1 6
#30910000000
1!
1%
1-
12
#30920000000
0!
0%
b10 *
0-
02
b10 6
#30930000000
1!
1%
1-
12
#30940000000
0!
0%
b11 *
0-
02
b11 6
#30950000000
1!
1%
1-
12
15
#30960000000
0!
0%
b100 *
0-
02
b100 6
#30970000000
1!
1%
1-
12
#30980000000
0!
0%
b101 *
0-
02
b101 6
#30990000000
1!
1%
1-
12
#31000000000
0!
0%
b110 *
0-
02
b110 6
#31010000000
1!
1%
1-
12
#31020000000
0!
0%
b111 *
0-
02
b111 6
#31030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#31040000000
0!
0%
b0 *
0-
02
b0 6
#31050000000
1!
1%
1-
12
#31060000000
0!
0%
b1 *
0-
02
b1 6
#31070000000
1!
1%
1-
12
#31080000000
0!
0%
b10 *
0-
02
b10 6
#31090000000
1!
1%
1-
12
#31100000000
0!
0%
b11 *
0-
02
b11 6
#31110000000
1!
1%
1-
12
15
#31120000000
0!
0%
b100 *
0-
02
b100 6
#31130000000
1!
1%
1-
12
#31140000000
0!
0%
b101 *
0-
02
b101 6
#31150000000
1!
1%
1-
12
#31160000000
0!
0%
b110 *
0-
02
b110 6
#31170000000
1!
1%
1-
12
#31180000000
0!
0%
b111 *
0-
02
b111 6
#31190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#31200000000
0!
0%
b0 *
0-
02
b0 6
#31210000000
1!
1%
1-
12
#31220000000
0!
0%
b1 *
0-
02
b1 6
#31230000000
1!
1%
1-
12
#31240000000
0!
0%
b10 *
0-
02
b10 6
#31250000000
1!
1%
1-
12
#31260000000
0!
0%
b11 *
0-
02
b11 6
#31270000000
1!
1%
1-
12
15
#31280000000
0!
0%
b100 *
0-
02
b100 6
#31290000000
1!
1%
1-
12
#31300000000
0!
0%
b101 *
0-
02
b101 6
#31310000000
1!
1%
1-
12
#31320000000
0!
0%
b110 *
0-
02
b110 6
#31330000000
1!
1%
1-
12
#31340000000
0!
0%
b111 *
0-
02
b111 6
#31350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#31360000000
0!
0%
b0 *
0-
02
b0 6
#31370000000
1!
1%
1-
12
#31380000000
0!
0%
b1 *
0-
02
b1 6
#31390000000
1!
1%
1-
12
#31400000000
0!
0%
b10 *
0-
02
b10 6
#31410000000
1!
1%
1-
12
#31420000000
0!
0%
b11 *
0-
02
b11 6
#31430000000
1!
1%
1-
12
15
#31440000000
0!
0%
b100 *
0-
02
b100 6
#31450000000
1!
1%
1-
12
#31460000000
0!
0%
b101 *
0-
02
b101 6
#31470000000
1!
1%
1-
12
#31480000000
0!
0%
b110 *
0-
02
b110 6
#31490000000
1!
1%
1-
12
#31500000000
0!
0%
b111 *
0-
02
b111 6
#31510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#31520000000
0!
0%
b0 *
0-
02
b0 6
#31530000000
1!
1%
1-
12
#31540000000
0!
0%
b1 *
0-
02
b1 6
#31550000000
1!
1%
1-
12
#31560000000
0!
0%
b10 *
0-
02
b10 6
#31570000000
1!
1%
1-
12
#31580000000
0!
0%
b11 *
0-
02
b11 6
#31590000000
1!
1%
1-
12
15
#31600000000
0!
0%
b100 *
0-
02
b100 6
#31610000000
1!
1%
1-
12
#31620000000
0!
0%
b101 *
0-
02
b101 6
#31630000000
1!
1%
1-
12
#31640000000
0!
0%
b110 *
0-
02
b110 6
#31650000000
1!
1%
1-
12
#31660000000
0!
0%
b111 *
0-
02
b111 6
#31670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#31680000000
0!
0%
b0 *
0-
02
b0 6
#31690000000
1!
1%
1-
12
#31700000000
0!
0%
b1 *
0-
02
b1 6
#31710000000
1!
1%
1-
12
#31720000000
0!
0%
b10 *
0-
02
b10 6
#31730000000
1!
1%
1-
12
#31740000000
0!
0%
b11 *
0-
02
b11 6
#31750000000
1!
1%
1-
12
15
#31760000000
0!
0%
b100 *
0-
02
b100 6
#31770000000
1!
1%
1-
12
#31780000000
0!
0%
b101 *
0-
02
b101 6
#31790000000
1!
1%
1-
12
#31800000000
0!
0%
b110 *
0-
02
b110 6
#31810000000
1!
1%
1-
12
#31820000000
0!
0%
b111 *
0-
02
b111 6
#31830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#31840000000
0!
0%
b0 *
0-
02
b0 6
#31850000000
1!
1%
1-
12
#31860000000
0!
0%
b1 *
0-
02
b1 6
#31870000000
1!
1%
1-
12
#31880000000
0!
0%
b10 *
0-
02
b10 6
#31890000000
1!
1%
1-
12
#31900000000
0!
0%
b11 *
0-
02
b11 6
#31910000000
1!
1%
1-
12
15
#31920000000
0!
0%
b100 *
0-
02
b100 6
#31930000000
1!
1%
1-
12
#31940000000
0!
0%
b101 *
0-
02
b101 6
#31950000000
1!
1%
1-
12
#31960000000
0!
0%
b110 *
0-
02
b110 6
#31970000000
1!
1%
1-
12
#31980000000
0!
0%
b111 *
0-
02
b111 6
#31990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#32000000000
0!
0%
b0 *
0-
02
b0 6
#32010000000
1!
1%
1-
12
#32020000000
0!
0%
b1 *
0-
02
b1 6
#32030000000
1!
1%
1-
12
#32040000000
0!
0%
b10 *
0-
02
b10 6
#32050000000
1!
1%
1-
12
#32060000000
0!
0%
b11 *
0-
02
b11 6
#32070000000
1!
1%
1-
12
15
#32080000000
0!
0%
b100 *
0-
02
b100 6
#32090000000
1!
1%
1-
12
#32100000000
0!
0%
b101 *
0-
02
b101 6
#32110000000
1!
1%
1-
12
#32120000000
0!
0%
b110 *
0-
02
b110 6
#32130000000
1!
1%
1-
12
#32140000000
0!
0%
b111 *
0-
02
b111 6
#32150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#32160000000
0!
0%
b0 *
0-
02
b0 6
#32170000000
1!
1%
1-
12
#32180000000
0!
0%
b1 *
0-
02
b1 6
#32190000000
1!
1%
1-
12
#32200000000
0!
0%
b10 *
0-
02
b10 6
#32210000000
1!
1%
1-
12
#32220000000
0!
0%
b11 *
0-
02
b11 6
#32230000000
1!
1%
1-
12
15
#32240000000
0!
0%
b100 *
0-
02
b100 6
#32250000000
1!
1%
1-
12
#32260000000
0!
0%
b101 *
0-
02
b101 6
#32270000000
1!
1%
1-
12
#32280000000
0!
0%
b110 *
0-
02
b110 6
#32290000000
1!
1%
1-
12
#32300000000
0!
0%
b111 *
0-
02
b111 6
#32310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#32320000000
0!
0%
b0 *
0-
02
b0 6
#32330000000
1!
1%
1-
12
#32340000000
0!
0%
b1 *
0-
02
b1 6
#32350000000
1!
1%
1-
12
#32360000000
0!
0%
b10 *
0-
02
b10 6
#32370000000
1!
1%
1-
12
#32380000000
0!
0%
b11 *
0-
02
b11 6
#32390000000
1!
1%
1-
12
15
#32400000000
0!
0%
b100 *
0-
02
b100 6
#32410000000
1!
1%
1-
12
#32420000000
0!
0%
b101 *
0-
02
b101 6
#32430000000
1!
1%
1-
12
#32440000000
0!
0%
b110 *
0-
02
b110 6
#32450000000
1!
1%
1-
12
#32460000000
0!
0%
b111 *
0-
02
b111 6
#32470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#32480000000
0!
0%
b0 *
0-
02
b0 6
#32490000000
1!
1%
1-
12
#32500000000
0!
0%
b1 *
0-
02
b1 6
#32510000000
1!
1%
1-
12
#32520000000
0!
0%
b10 *
0-
02
b10 6
#32530000000
1!
1%
1-
12
#32540000000
0!
0%
b11 *
0-
02
b11 6
#32550000000
1!
1%
1-
12
15
#32560000000
0!
0%
b100 *
0-
02
b100 6
#32570000000
1!
1%
1-
12
#32580000000
0!
0%
b101 *
0-
02
b101 6
#32590000000
1!
1%
1-
12
#32600000000
0!
0%
b110 *
0-
02
b110 6
#32610000000
1!
1%
1-
12
#32620000000
0!
0%
b111 *
0-
02
b111 6
#32630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#32640000000
0!
0%
b0 *
0-
02
b0 6
#32650000000
1!
1%
1-
12
#32660000000
0!
0%
b1 *
0-
02
b1 6
#32670000000
1!
1%
1-
12
#32680000000
0!
0%
b10 *
0-
02
b10 6
#32690000000
1!
1%
1-
12
#32700000000
0!
0%
b11 *
0-
02
b11 6
#32710000000
1!
1%
1-
12
15
#32720000000
0!
0%
b100 *
0-
02
b100 6
#32730000000
1!
1%
1-
12
#32740000000
0!
0%
b101 *
0-
02
b101 6
#32750000000
1!
1%
1-
12
#32760000000
0!
0%
b110 *
0-
02
b110 6
#32770000000
1!
1%
1-
12
#32780000000
0!
0%
b111 *
0-
02
b111 6
#32790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#32800000000
0!
0%
b0 *
0-
02
b0 6
#32810000000
1!
1%
1-
12
#32820000000
0!
0%
b1 *
0-
02
b1 6
#32830000000
1!
1%
1-
12
#32840000000
0!
0%
b10 *
0-
02
b10 6
#32850000000
1!
1%
1-
12
#32860000000
0!
0%
b11 *
0-
02
b11 6
#32870000000
1!
1%
1-
12
15
#32880000000
0!
0%
b100 *
0-
02
b100 6
#32890000000
1!
1%
1-
12
#32900000000
0!
0%
b101 *
0-
02
b101 6
#32910000000
1!
1%
1-
12
#32920000000
0!
0%
b110 *
0-
02
b110 6
#32930000000
1!
1%
1-
12
#32940000000
0!
0%
b111 *
0-
02
b111 6
#32950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#32960000000
0!
0%
b0 *
0-
02
b0 6
#32970000000
1!
1%
1-
12
#32980000000
0!
0%
b1 *
0-
02
b1 6
#32990000000
1!
1%
1-
12
#33000000000
0!
0%
b10 *
0-
02
b10 6
#33010000000
1!
1%
1-
12
#33020000000
0!
0%
b11 *
0-
02
b11 6
#33030000000
1!
1%
1-
12
15
#33040000000
0!
0%
b100 *
0-
02
b100 6
#33050000000
1!
1%
1-
12
#33060000000
0!
0%
b101 *
0-
02
b101 6
#33070000000
1!
1%
1-
12
#33080000000
0!
0%
b110 *
0-
02
b110 6
#33090000000
1!
1%
1-
12
#33100000000
0!
0%
b111 *
0-
02
b111 6
#33110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#33120000000
0!
0%
b0 *
0-
02
b0 6
#33130000000
1!
1%
1-
12
#33140000000
0!
0%
b1 *
0-
02
b1 6
#33150000000
1!
1%
1-
12
#33160000000
0!
0%
b10 *
0-
02
b10 6
#33170000000
1!
1%
1-
12
#33180000000
0!
0%
b11 *
0-
02
b11 6
#33190000000
1!
1%
1-
12
15
#33200000000
0!
0%
b100 *
0-
02
b100 6
#33210000000
1!
1%
1-
12
#33220000000
0!
0%
b101 *
0-
02
b101 6
#33230000000
1!
1%
1-
12
#33240000000
0!
0%
b110 *
0-
02
b110 6
#33250000000
1!
1%
1-
12
#33260000000
0!
0%
b111 *
0-
02
b111 6
#33270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#33280000000
0!
0%
b0 *
0-
02
b0 6
#33290000000
1!
1%
1-
12
#33300000000
0!
0%
b1 *
0-
02
b1 6
#33310000000
1!
1%
1-
12
#33320000000
0!
0%
b10 *
0-
02
b10 6
#33330000000
1!
1%
1-
12
#33340000000
0!
0%
b11 *
0-
02
b11 6
#33350000000
1!
1%
1-
12
15
#33360000000
0!
0%
b100 *
0-
02
b100 6
#33370000000
1!
1%
1-
12
#33380000000
0!
0%
b101 *
0-
02
b101 6
#33390000000
1!
1%
1-
12
#33400000000
0!
0%
b110 *
0-
02
b110 6
#33410000000
1!
1%
1-
12
#33420000000
0!
0%
b111 *
0-
02
b111 6
#33430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#33440000000
0!
0%
b0 *
0-
02
b0 6
#33450000000
1!
1%
1-
12
#33460000000
0!
0%
b1 *
0-
02
b1 6
#33470000000
1!
1%
1-
12
#33480000000
0!
0%
b10 *
0-
02
b10 6
#33490000000
1!
1%
1-
12
#33500000000
0!
0%
b11 *
0-
02
b11 6
#33510000000
1!
1%
1-
12
15
#33520000000
0!
0%
b100 *
0-
02
b100 6
#33530000000
1!
1%
1-
12
#33540000000
0!
0%
b101 *
0-
02
b101 6
#33550000000
1!
1%
1-
12
#33560000000
0!
0%
b110 *
0-
02
b110 6
#33570000000
1!
1%
1-
12
#33580000000
0!
0%
b111 *
0-
02
b111 6
#33590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#33600000000
0!
0%
b0 *
0-
02
b0 6
#33610000000
1!
1%
1-
12
#33620000000
0!
0%
b1 *
0-
02
b1 6
#33630000000
1!
1%
1-
12
#33640000000
0!
0%
b10 *
0-
02
b10 6
#33650000000
1!
1%
1-
12
#33660000000
0!
0%
b11 *
0-
02
b11 6
#33670000000
1!
1%
1-
12
15
#33680000000
0!
0%
b100 *
0-
02
b100 6
#33690000000
1!
1%
1-
12
#33700000000
0!
0%
b101 *
0-
02
b101 6
#33710000000
1!
1%
1-
12
#33720000000
0!
0%
b110 *
0-
02
b110 6
#33730000000
1!
1%
1-
12
#33740000000
0!
0%
b111 *
0-
02
b111 6
#33750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#33760000000
0!
0%
b0 *
0-
02
b0 6
#33770000000
1!
1%
1-
12
#33780000000
0!
0%
b1 *
0-
02
b1 6
#33790000000
1!
1%
1-
12
#33800000000
0!
0%
b10 *
0-
02
b10 6
#33810000000
1!
1%
1-
12
#33820000000
0!
0%
b11 *
0-
02
b11 6
#33830000000
1!
1%
1-
12
15
#33840000000
0!
0%
b100 *
0-
02
b100 6
#33850000000
1!
1%
1-
12
#33860000000
0!
0%
b101 *
0-
02
b101 6
#33870000000
1!
1%
1-
12
#33880000000
0!
0%
b110 *
0-
02
b110 6
#33890000000
1!
1%
1-
12
#33900000000
0!
0%
b111 *
0-
02
b111 6
#33910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#33920000000
0!
0%
b0 *
0-
02
b0 6
#33930000000
1!
1%
1-
12
#33940000000
0!
0%
b1 *
0-
02
b1 6
#33950000000
1!
1%
1-
12
#33960000000
0!
0%
b10 *
0-
02
b10 6
#33970000000
1!
1%
1-
12
#33980000000
0!
0%
b11 *
0-
02
b11 6
#33990000000
1!
1%
1-
12
15
#34000000000
0!
0%
b100 *
0-
02
b100 6
#34010000000
1!
1%
1-
12
#34020000000
0!
0%
b101 *
0-
02
b101 6
#34030000000
1!
1%
1-
12
#34040000000
0!
0%
b110 *
0-
02
b110 6
#34050000000
1!
1%
1-
12
#34060000000
0!
0%
b111 *
0-
02
b111 6
#34070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#34080000000
0!
0%
b0 *
0-
02
b0 6
#34090000000
1!
1%
1-
12
#34100000000
0!
0%
b1 *
0-
02
b1 6
#34110000000
1!
1%
1-
12
#34120000000
0!
0%
b10 *
0-
02
b10 6
#34130000000
1!
1%
1-
12
#34140000000
0!
0%
b11 *
0-
02
b11 6
#34150000000
1!
1%
1-
12
15
#34160000000
0!
0%
b100 *
0-
02
b100 6
#34170000000
1!
1%
1-
12
#34180000000
0!
0%
b101 *
0-
02
b101 6
#34190000000
1!
1%
1-
12
#34200000000
0!
0%
b110 *
0-
02
b110 6
#34210000000
1!
1%
1-
12
#34220000000
0!
0%
b111 *
0-
02
b111 6
#34230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#34240000000
0!
0%
b0 *
0-
02
b0 6
#34250000000
1!
1%
1-
12
#34260000000
0!
0%
b1 *
0-
02
b1 6
#34270000000
1!
1%
1-
12
#34280000000
0!
0%
b10 *
0-
02
b10 6
#34290000000
1!
1%
1-
12
#34300000000
0!
0%
b11 *
0-
02
b11 6
#34310000000
1!
1%
1-
12
15
#34320000000
0!
0%
b100 *
0-
02
b100 6
#34330000000
1!
1%
1-
12
#34340000000
0!
0%
b101 *
0-
02
b101 6
#34350000000
1!
1%
1-
12
#34360000000
0!
0%
b110 *
0-
02
b110 6
#34370000000
1!
1%
1-
12
#34380000000
0!
0%
b111 *
0-
02
b111 6
#34390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#34400000000
0!
0%
b0 *
0-
02
b0 6
#34410000000
1!
1%
1-
12
#34420000000
0!
0%
b1 *
0-
02
b1 6
#34430000000
1!
1%
1-
12
#34440000000
0!
0%
b10 *
0-
02
b10 6
#34450000000
1!
1%
1-
12
#34460000000
0!
0%
b11 *
0-
02
b11 6
#34470000000
1!
1%
1-
12
15
#34480000000
0!
0%
b100 *
0-
02
b100 6
#34490000000
1!
1%
1-
12
#34500000000
0!
0%
b101 *
0-
02
b101 6
#34510000000
1!
1%
1-
12
#34520000000
0!
0%
b110 *
0-
02
b110 6
#34530000000
1!
1%
1-
12
#34540000000
0!
0%
b111 *
0-
02
b111 6
#34550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#34560000000
0!
0%
b0 *
0-
02
b0 6
#34570000000
1!
1%
1-
12
#34580000000
0!
0%
b1 *
0-
02
b1 6
#34590000000
1!
1%
1-
12
#34600000000
0!
0%
b10 *
0-
02
b10 6
#34610000000
1!
1%
1-
12
#34620000000
0!
0%
b11 *
0-
02
b11 6
#34630000000
1!
1%
1-
12
15
#34640000000
0!
0%
b100 *
0-
02
b100 6
#34650000000
1!
1%
1-
12
#34660000000
0!
0%
b101 *
0-
02
b101 6
#34670000000
1!
1%
1-
12
#34680000000
0!
0%
b110 *
0-
02
b110 6
#34690000000
1!
1%
1-
12
#34700000000
0!
0%
b111 *
0-
02
b111 6
#34710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#34720000000
0!
0%
b0 *
0-
02
b0 6
#34730000000
1!
1%
1-
12
#34740000000
0!
0%
b1 *
0-
02
b1 6
#34750000000
1!
1%
1-
12
#34760000000
0!
0%
b10 *
0-
02
b10 6
#34770000000
1!
1%
1-
12
#34780000000
0!
0%
b11 *
0-
02
b11 6
#34790000000
1!
1%
1-
12
15
#34800000000
0!
0%
b100 *
0-
02
b100 6
#34810000000
1!
1%
1-
12
#34820000000
0!
0%
b101 *
0-
02
b101 6
#34830000000
1!
1%
1-
12
#34840000000
0!
0%
b110 *
0-
02
b110 6
#34850000000
1!
1%
1-
12
#34860000000
0!
0%
b111 *
0-
02
b111 6
#34870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#34880000000
0!
0%
b0 *
0-
02
b0 6
#34890000000
1!
1%
1-
12
#34900000000
0!
0%
b1 *
0-
02
b1 6
#34910000000
1!
1%
1-
12
#34920000000
0!
0%
b10 *
0-
02
b10 6
#34930000000
1!
1%
1-
12
#34940000000
0!
0%
b11 *
0-
02
b11 6
#34950000000
1!
1%
1-
12
15
#34960000000
0!
0%
b100 *
0-
02
b100 6
#34970000000
1!
1%
1-
12
#34980000000
0!
0%
b101 *
0-
02
b101 6
#34990000000
1!
1%
1-
12
#35000000000
0!
0%
b110 *
0-
02
b110 6
#35010000000
1!
1%
1-
12
#35020000000
0!
0%
b111 *
0-
02
b111 6
#35030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#35040000000
0!
0%
b0 *
0-
02
b0 6
#35050000000
1!
1%
1-
12
#35060000000
0!
0%
b1 *
0-
02
b1 6
#35070000000
1!
1%
1-
12
#35080000000
0!
0%
b10 *
0-
02
b10 6
#35090000000
1!
1%
1-
12
#35100000000
0!
0%
b11 *
0-
02
b11 6
#35110000000
1!
1%
1-
12
15
#35120000000
0!
0%
b100 *
0-
02
b100 6
#35130000000
1!
1%
1-
12
#35140000000
0!
0%
b101 *
0-
02
b101 6
#35150000000
1!
1%
1-
12
#35160000000
0!
0%
b110 *
0-
02
b110 6
#35170000000
1!
1%
1-
12
#35180000000
0!
0%
b111 *
0-
02
b111 6
#35190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#35200000000
0!
0%
b0 *
0-
02
b0 6
#35210000000
1!
1%
1-
12
#35220000000
0!
0%
b1 *
0-
02
b1 6
#35230000000
1!
1%
1-
12
#35240000000
0!
0%
b10 *
0-
02
b10 6
#35250000000
1!
1%
1-
12
#35260000000
0!
0%
b11 *
0-
02
b11 6
#35270000000
1!
1%
1-
12
15
#35280000000
0!
0%
b100 *
0-
02
b100 6
#35290000000
1!
1%
1-
12
#35300000000
0!
0%
b101 *
0-
02
b101 6
#35310000000
1!
1%
1-
12
#35320000000
0!
0%
b110 *
0-
02
b110 6
#35330000000
1!
1%
1-
12
#35340000000
0!
0%
b111 *
0-
02
b111 6
#35350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#35360000000
0!
0%
b0 *
0-
02
b0 6
#35370000000
1!
1%
1-
12
#35380000000
0!
0%
b1 *
0-
02
b1 6
#35390000000
1!
1%
1-
12
#35400000000
0!
0%
b10 *
0-
02
b10 6
#35410000000
1!
1%
1-
12
#35420000000
0!
0%
b11 *
0-
02
b11 6
#35430000000
1!
1%
1-
12
15
#35440000000
0!
0%
b100 *
0-
02
b100 6
#35450000000
1!
1%
1-
12
#35460000000
0!
0%
b101 *
0-
02
b101 6
#35470000000
1!
1%
1-
12
#35480000000
0!
0%
b110 *
0-
02
b110 6
#35490000000
1!
1%
1-
12
#35500000000
0!
0%
b111 *
0-
02
b111 6
#35510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#35520000000
0!
0%
b0 *
0-
02
b0 6
#35530000000
1!
1%
1-
12
#35540000000
0!
0%
b1 *
0-
02
b1 6
#35550000000
1!
1%
1-
12
#35560000000
0!
0%
b10 *
0-
02
b10 6
#35570000000
1!
1%
1-
12
#35580000000
0!
0%
b11 *
0-
02
b11 6
#35590000000
1!
1%
1-
12
15
#35600000000
0!
0%
b100 *
0-
02
b100 6
#35610000000
1!
1%
1-
12
#35620000000
0!
0%
b101 *
0-
02
b101 6
#35630000000
1!
1%
1-
12
#35640000000
0!
0%
b110 *
0-
02
b110 6
#35650000000
1!
1%
1-
12
#35660000000
0!
0%
b111 *
0-
02
b111 6
#35670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#35680000000
0!
0%
b0 *
0-
02
b0 6
#35690000000
1!
1%
1-
12
#35700000000
0!
0%
b1 *
0-
02
b1 6
#35710000000
1!
1%
1-
12
#35720000000
0!
0%
b10 *
0-
02
b10 6
#35730000000
1!
1%
1-
12
#35740000000
0!
0%
b11 *
0-
02
b11 6
#35750000000
1!
1%
1-
12
15
#35760000000
0!
0%
b100 *
0-
02
b100 6
#35770000000
1!
1%
1-
12
#35780000000
0!
0%
b101 *
0-
02
b101 6
#35790000000
1!
1%
1-
12
#35800000000
0!
0%
b110 *
0-
02
b110 6
#35810000000
1!
1%
1-
12
#35820000000
0!
0%
b111 *
0-
02
b111 6
#35830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#35840000000
0!
0%
b0 *
0-
02
b0 6
#35850000000
1!
1%
1-
12
#35860000000
0!
0%
b1 *
0-
02
b1 6
#35870000000
1!
1%
1-
12
#35880000000
0!
0%
b10 *
0-
02
b10 6
#35890000000
1!
1%
1-
12
#35900000000
0!
0%
b11 *
0-
02
b11 6
#35910000000
1!
1%
1-
12
15
#35920000000
0!
0%
b100 *
0-
02
b100 6
#35930000000
1!
1%
1-
12
#35940000000
0!
0%
b101 *
0-
02
b101 6
#35950000000
1!
1%
1-
12
#35960000000
0!
0%
b110 *
0-
02
b110 6
#35970000000
1!
1%
1-
12
#35980000000
0!
0%
b111 *
0-
02
b111 6
#35990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#36000000000
0!
0%
b0 *
0-
02
b0 6
#36010000000
1!
1%
1-
12
#36020000000
0!
0%
b1 *
0-
02
b1 6
#36030000000
1!
1%
1-
12
#36040000000
0!
0%
b10 *
0-
02
b10 6
#36050000000
1!
1%
1-
12
#36060000000
0!
0%
b11 *
0-
02
b11 6
#36070000000
1!
1%
1-
12
15
#36080000000
0!
0%
b100 *
0-
02
b100 6
#36090000000
1!
1%
1-
12
#36100000000
0!
0%
b101 *
0-
02
b101 6
#36110000000
1!
1%
1-
12
#36120000000
0!
0%
b110 *
0-
02
b110 6
#36130000000
1!
1%
1-
12
#36140000000
0!
0%
b111 *
0-
02
b111 6
#36150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#36160000000
0!
0%
b0 *
0-
02
b0 6
#36170000000
1!
1%
1-
12
#36180000000
0!
0%
b1 *
0-
02
b1 6
#36190000000
1!
1%
1-
12
#36200000000
0!
0%
b10 *
0-
02
b10 6
#36210000000
1!
1%
1-
12
#36220000000
0!
0%
b11 *
0-
02
b11 6
#36230000000
1!
1%
1-
12
15
#36240000000
0!
0%
b100 *
0-
02
b100 6
#36250000000
1!
1%
1-
12
#36260000000
0!
0%
b101 *
0-
02
b101 6
#36270000000
1!
1%
1-
12
#36280000000
0!
0%
b110 *
0-
02
b110 6
#36290000000
1!
1%
1-
12
#36300000000
0!
0%
b111 *
0-
02
b111 6
#36310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#36320000000
0!
0%
b0 *
0-
02
b0 6
#36330000000
1!
1%
1-
12
#36340000000
0!
0%
b1 *
0-
02
b1 6
#36350000000
1!
1%
1-
12
#36360000000
0!
0%
b10 *
0-
02
b10 6
#36370000000
1!
1%
1-
12
#36380000000
0!
0%
b11 *
0-
02
b11 6
#36390000000
1!
1%
1-
12
15
#36400000000
0!
0%
b100 *
0-
02
b100 6
#36410000000
1!
1%
1-
12
#36420000000
0!
0%
b101 *
0-
02
b101 6
#36430000000
1!
1%
1-
12
#36440000000
0!
0%
b110 *
0-
02
b110 6
#36450000000
1!
1%
1-
12
#36460000000
0!
0%
b111 *
0-
02
b111 6
#36470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#36480000000
0!
0%
b0 *
0-
02
b0 6
#36490000000
1!
1%
1-
12
#36500000000
0!
0%
b1 *
0-
02
b1 6
#36510000000
1!
1%
1-
12
#36520000000
0!
0%
b10 *
0-
02
b10 6
#36530000000
1!
1%
1-
12
#36540000000
0!
0%
b11 *
0-
02
b11 6
#36550000000
1!
1%
1-
12
15
#36560000000
0!
0%
b100 *
0-
02
b100 6
#36570000000
1!
1%
1-
12
#36580000000
0!
0%
b101 *
0-
02
b101 6
#36590000000
1!
1%
1-
12
#36600000000
0!
0%
b110 *
0-
02
b110 6
#36610000000
1!
1%
1-
12
#36620000000
0!
0%
b111 *
0-
02
b111 6
#36630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#36640000000
0!
0%
b0 *
0-
02
b0 6
#36650000000
1!
1%
1-
12
#36660000000
0!
0%
b1 *
0-
02
b1 6
#36670000000
1!
1%
1-
12
#36680000000
0!
0%
b10 *
0-
02
b10 6
#36690000000
1!
1%
1-
12
#36700000000
0!
0%
b11 *
0-
02
b11 6
#36710000000
1!
1%
1-
12
15
#36720000000
0!
0%
b100 *
0-
02
b100 6
#36730000000
1!
1%
1-
12
#36740000000
0!
0%
b101 *
0-
02
b101 6
#36750000000
1!
1%
1-
12
#36760000000
0!
0%
b110 *
0-
02
b110 6
#36770000000
1!
1%
1-
12
#36780000000
0!
0%
b111 *
0-
02
b111 6
#36790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#36800000000
0!
0%
b0 *
0-
02
b0 6
#36810000000
1!
1%
1-
12
#36820000000
0!
0%
b1 *
0-
02
b1 6
#36830000000
1!
1%
1-
12
#36840000000
0!
0%
b10 *
0-
02
b10 6
#36850000000
1!
1%
1-
12
#36860000000
0!
0%
b11 *
0-
02
b11 6
#36870000000
1!
1%
1-
12
15
#36880000000
0!
0%
b100 *
0-
02
b100 6
#36890000000
1!
1%
1-
12
#36900000000
0!
0%
b101 *
0-
02
b101 6
#36910000000
1!
1%
1-
12
#36920000000
0!
0%
b110 *
0-
02
b110 6
#36930000000
1!
1%
1-
12
#36940000000
0!
0%
b111 *
0-
02
b111 6
#36950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#36960000000
0!
0%
b0 *
0-
02
b0 6
#36970000000
1!
1%
1-
12
#36980000000
0!
0%
b1 *
0-
02
b1 6
#36990000000
1!
1%
1-
12
#37000000000
0!
0%
b10 *
0-
02
b10 6
#37010000000
1!
1%
1-
12
#37020000000
0!
0%
b11 *
0-
02
b11 6
#37030000000
1!
1%
1-
12
15
#37040000000
0!
0%
b100 *
0-
02
b100 6
#37050000000
1!
1%
1-
12
#37060000000
0!
0%
b101 *
0-
02
b101 6
#37070000000
1!
1%
1-
12
#37080000000
0!
0%
b110 *
0-
02
b110 6
#37090000000
1!
1%
1-
12
#37100000000
0!
0%
b111 *
0-
02
b111 6
#37110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#37120000000
0!
0%
b0 *
0-
02
b0 6
#37130000000
1!
1%
1-
12
#37140000000
0!
0%
b1 *
0-
02
b1 6
#37150000000
1!
1%
1-
12
#37160000000
0!
0%
b10 *
0-
02
b10 6
#37170000000
1!
1%
1-
12
#37180000000
0!
0%
b11 *
0-
02
b11 6
#37190000000
1!
1%
1-
12
15
#37200000000
0!
0%
b100 *
0-
02
b100 6
#37210000000
1!
1%
1-
12
#37220000000
0!
0%
b101 *
0-
02
b101 6
#37230000000
1!
1%
1-
12
#37240000000
0!
0%
b110 *
0-
02
b110 6
#37250000000
1!
1%
1-
12
#37260000000
0!
0%
b111 *
0-
02
b111 6
#37270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#37280000000
0!
0%
b0 *
0-
02
b0 6
#37290000000
1!
1%
1-
12
#37300000000
0!
0%
b1 *
0-
02
b1 6
#37310000000
1!
1%
1-
12
#37320000000
0!
0%
b10 *
0-
02
b10 6
#37330000000
1!
1%
1-
12
#37340000000
0!
0%
b11 *
0-
02
b11 6
#37350000000
1!
1%
1-
12
15
#37360000000
0!
0%
b100 *
0-
02
b100 6
#37370000000
1!
1%
1-
12
#37380000000
0!
0%
b101 *
0-
02
b101 6
#37390000000
1!
1%
1-
12
#37400000000
0!
0%
b110 *
0-
02
b110 6
#37410000000
1!
1%
1-
12
#37420000000
0!
0%
b111 *
0-
02
b111 6
#37430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#37440000000
0!
0%
b0 *
0-
02
b0 6
#37450000000
1!
1%
1-
12
#37460000000
0!
0%
b1 *
0-
02
b1 6
#37470000000
1!
1%
1-
12
#37480000000
0!
0%
b10 *
0-
02
b10 6
#37490000000
1!
1%
1-
12
#37500000000
0!
0%
b11 *
0-
02
b11 6
#37510000000
1!
1%
1-
12
15
#37520000000
0!
0%
b100 *
0-
02
b100 6
#37530000000
1!
1%
1-
12
#37540000000
0!
0%
b101 *
0-
02
b101 6
#37550000000
1!
1%
1-
12
#37560000000
0!
0%
b110 *
0-
02
b110 6
#37570000000
1!
1%
1-
12
#37580000000
0!
0%
b111 *
0-
02
b111 6
#37590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#37600000000
0!
0%
b0 *
0-
02
b0 6
#37610000000
1!
1%
1-
12
#37620000000
0!
0%
b1 *
0-
02
b1 6
#37630000000
1!
1%
1-
12
#37640000000
0!
0%
b10 *
0-
02
b10 6
#37650000000
1!
1%
1-
12
#37660000000
0!
0%
b11 *
0-
02
b11 6
#37670000000
1!
1%
1-
12
15
#37680000000
0!
0%
b100 *
0-
02
b100 6
#37690000000
1!
1%
1-
12
#37700000000
0!
0%
b101 *
0-
02
b101 6
#37710000000
1!
1%
1-
12
#37720000000
0!
0%
b110 *
0-
02
b110 6
#37730000000
1!
1%
1-
12
#37740000000
0!
0%
b111 *
0-
02
b111 6
#37750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#37760000000
0!
0%
b0 *
0-
02
b0 6
#37770000000
1!
1%
1-
12
#37780000000
0!
0%
b1 *
0-
02
b1 6
#37790000000
1!
1%
1-
12
#37800000000
0!
0%
b10 *
0-
02
b10 6
#37810000000
1!
1%
1-
12
#37820000000
0!
0%
b11 *
0-
02
b11 6
#37830000000
1!
1%
1-
12
15
#37840000000
0!
0%
b100 *
0-
02
b100 6
#37850000000
1!
1%
1-
12
#37860000000
0!
0%
b101 *
0-
02
b101 6
#37870000000
1!
1%
1-
12
#37880000000
0!
0%
b110 *
0-
02
b110 6
#37890000000
1!
1%
1-
12
#37900000000
0!
0%
b111 *
0-
02
b111 6
#37910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#37920000000
0!
0%
b0 *
0-
02
b0 6
#37930000000
1!
1%
1-
12
#37940000000
0!
0%
b1 *
0-
02
b1 6
#37950000000
1!
1%
1-
12
#37960000000
0!
0%
b10 *
0-
02
b10 6
#37970000000
1!
1%
1-
12
#37980000000
0!
0%
b11 *
0-
02
b11 6
#37990000000
1!
1%
1-
12
15
#38000000000
0!
0%
b100 *
0-
02
b100 6
#38010000000
1!
1%
1-
12
#38020000000
0!
0%
b101 *
0-
02
b101 6
#38030000000
1!
1%
1-
12
#38040000000
0!
0%
b110 *
0-
02
b110 6
#38050000000
1!
1%
1-
12
#38060000000
0!
0%
b111 *
0-
02
b111 6
#38070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#38080000000
0!
0%
b0 *
0-
02
b0 6
#38090000000
1!
1%
1-
12
#38100000000
0!
0%
b1 *
0-
02
b1 6
#38110000000
1!
1%
1-
12
#38120000000
0!
0%
b10 *
0-
02
b10 6
#38130000000
1!
1%
1-
12
#38140000000
0!
0%
b11 *
0-
02
b11 6
#38150000000
1!
1%
1-
12
15
#38160000000
0!
0%
b100 *
0-
02
b100 6
#38170000000
1!
1%
1-
12
#38180000000
0!
0%
b101 *
0-
02
b101 6
#38190000000
1!
1%
1-
12
#38200000000
0!
0%
b110 *
0-
02
b110 6
#38210000000
1!
1%
1-
12
#38220000000
0!
0%
b111 *
0-
02
b111 6
#38230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#38240000000
0!
0%
b0 *
0-
02
b0 6
#38250000000
1!
1%
1-
12
#38260000000
0!
0%
b1 *
0-
02
b1 6
#38270000000
1!
1%
1-
12
#38280000000
0!
0%
b10 *
0-
02
b10 6
#38290000000
1!
1%
1-
12
#38300000000
0!
0%
b11 *
0-
02
b11 6
#38310000000
1!
1%
1-
12
15
#38320000000
0!
0%
b100 *
0-
02
b100 6
#38330000000
1!
1%
1-
12
#38340000000
0!
0%
b101 *
0-
02
b101 6
#38350000000
1!
1%
1-
12
#38360000000
0!
0%
b110 *
0-
02
b110 6
#38370000000
1!
1%
1-
12
#38380000000
0!
0%
b111 *
0-
02
b111 6
#38390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#38400000000
0!
0%
b0 *
0-
02
b0 6
#38410000000
1!
1%
1-
12
#38420000000
0!
0%
b1 *
0-
02
b1 6
#38430000000
1!
1%
1-
12
#38440000000
0!
0%
b10 *
0-
02
b10 6
#38450000000
1!
1%
1-
12
#38460000000
0!
0%
b11 *
0-
02
b11 6
#38470000000
1!
1%
1-
12
15
#38480000000
0!
0%
b100 *
0-
02
b100 6
#38490000000
1!
1%
1-
12
#38500000000
0!
0%
b101 *
0-
02
b101 6
#38510000000
1!
1%
1-
12
#38520000000
0!
0%
b110 *
0-
02
b110 6
#38530000000
1!
1%
1-
12
#38540000000
0!
0%
b111 *
0-
02
b111 6
#38550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#38560000000
0!
0%
b0 *
0-
02
b0 6
#38570000000
1!
1%
1-
12
#38580000000
0!
0%
b1 *
0-
02
b1 6
#38590000000
1!
1%
1-
12
#38600000000
0!
0%
b10 *
0-
02
b10 6
#38610000000
1!
1%
1-
12
#38620000000
0!
0%
b11 *
0-
02
b11 6
#38630000000
1!
1%
1-
12
15
#38640000000
0!
0%
b100 *
0-
02
b100 6
#38650000000
1!
1%
1-
12
#38660000000
0!
0%
b101 *
0-
02
b101 6
#38670000000
1!
1%
1-
12
#38680000000
0!
0%
b110 *
0-
02
b110 6
#38690000000
1!
1%
1-
12
#38700000000
0!
0%
b111 *
0-
02
b111 6
#38710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#38720000000
0!
0%
b0 *
0-
02
b0 6
#38730000000
1!
1%
1-
12
#38740000000
0!
0%
b1 *
0-
02
b1 6
#38750000000
1!
1%
1-
12
#38760000000
0!
0%
b10 *
0-
02
b10 6
#38770000000
1!
1%
1-
12
#38780000000
0!
0%
b11 *
0-
02
b11 6
#38790000000
1!
1%
1-
12
15
#38800000000
0!
0%
b100 *
0-
02
b100 6
#38810000000
1!
1%
1-
12
#38820000000
0!
0%
b101 *
0-
02
b101 6
#38830000000
1!
1%
1-
12
#38840000000
0!
0%
b110 *
0-
02
b110 6
#38850000000
1!
1%
1-
12
#38860000000
0!
0%
b111 *
0-
02
b111 6
#38870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#38880000000
0!
0%
b0 *
0-
02
b0 6
#38890000000
1!
1%
1-
12
#38900000000
0!
0%
b1 *
0-
02
b1 6
#38910000000
1!
1%
1-
12
#38920000000
0!
0%
b10 *
0-
02
b10 6
#38930000000
1!
1%
1-
12
#38940000000
0!
0%
b11 *
0-
02
b11 6
#38950000000
1!
1%
1-
12
15
#38960000000
0!
0%
b100 *
0-
02
b100 6
#38970000000
1!
1%
1-
12
#38980000000
0!
0%
b101 *
0-
02
b101 6
#38990000000
1!
1%
1-
12
#39000000000
0!
0%
b110 *
0-
02
b110 6
#39010000000
1!
1%
1-
12
#39020000000
0!
0%
b111 *
0-
02
b111 6
#39030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#39040000000
0!
0%
b0 *
0-
02
b0 6
#39050000000
1!
1%
1-
12
#39060000000
0!
0%
b1 *
0-
02
b1 6
#39070000000
1!
1%
1-
12
#39080000000
0!
0%
b10 *
0-
02
b10 6
#39090000000
1!
1%
1-
12
#39100000000
0!
0%
b11 *
0-
02
b11 6
#39110000000
1!
1%
1-
12
15
#39120000000
0!
0%
b100 *
0-
02
b100 6
#39130000000
1!
1%
1-
12
#39140000000
0!
0%
b101 *
0-
02
b101 6
#39150000000
1!
1%
1-
12
#39160000000
0!
0%
b110 *
0-
02
b110 6
#39170000000
1!
1%
1-
12
#39180000000
0!
0%
b111 *
0-
02
b111 6
#39190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#39200000000
0!
0%
b0 *
0-
02
b0 6
#39210000000
1!
1%
1-
12
#39220000000
0!
0%
b1 *
0-
02
b1 6
#39230000000
1!
1%
1-
12
#39240000000
0!
0%
b10 *
0-
02
b10 6
#39250000000
1!
1%
1-
12
#39260000000
0!
0%
b11 *
0-
02
b11 6
#39270000000
1!
1%
1-
12
15
#39280000000
0!
0%
b100 *
0-
02
b100 6
#39290000000
1!
1%
1-
12
#39300000000
0!
0%
b101 *
0-
02
b101 6
#39310000000
1!
1%
1-
12
#39320000000
0!
0%
b110 *
0-
02
b110 6
#39330000000
1!
1%
1-
12
#39340000000
0!
0%
b111 *
0-
02
b111 6
#39350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#39360000000
0!
0%
b0 *
0-
02
b0 6
#39370000000
1!
1%
1-
12
#39380000000
0!
0%
b1 *
0-
02
b1 6
#39390000000
1!
1%
1-
12
#39400000000
0!
0%
b10 *
0-
02
b10 6
#39410000000
1!
1%
1-
12
#39420000000
0!
0%
b11 *
0-
02
b11 6
#39430000000
1!
1%
1-
12
15
#39440000000
0!
0%
b100 *
0-
02
b100 6
#39450000000
1!
1%
1-
12
#39460000000
0!
0%
b101 *
0-
02
b101 6
#39470000000
1!
1%
1-
12
#39480000000
0!
0%
b110 *
0-
02
b110 6
#39490000000
1!
1%
1-
12
#39500000000
0!
0%
b111 *
0-
02
b111 6
#39510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#39520000000
0!
0%
b0 *
0-
02
b0 6
#39530000000
1!
1%
1-
12
#39540000000
0!
0%
b1 *
0-
02
b1 6
#39550000000
1!
1%
1-
12
#39560000000
0!
0%
b10 *
0-
02
b10 6
#39570000000
1!
1%
1-
12
#39580000000
0!
0%
b11 *
0-
02
b11 6
#39590000000
1!
1%
1-
12
15
#39600000000
0!
0%
b100 *
0-
02
b100 6
#39610000000
1!
1%
1-
12
#39620000000
0!
0%
b101 *
0-
02
b101 6
#39630000000
1!
1%
1-
12
#39640000000
0!
0%
b110 *
0-
02
b110 6
#39650000000
1!
1%
1-
12
#39660000000
0!
0%
b111 *
0-
02
b111 6
#39670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#39680000000
0!
0%
b0 *
0-
02
b0 6
#39690000000
1!
1%
1-
12
#39700000000
0!
0%
b1 *
0-
02
b1 6
#39710000000
1!
1%
1-
12
#39720000000
0!
0%
b10 *
0-
02
b10 6
#39730000000
1!
1%
1-
12
#39740000000
0!
0%
b11 *
0-
02
b11 6
#39750000000
1!
1%
1-
12
15
#39760000000
0!
0%
b100 *
0-
02
b100 6
#39770000000
1!
1%
1-
12
#39780000000
0!
0%
b101 *
0-
02
b101 6
#39790000000
1!
1%
1-
12
#39800000000
0!
0%
b110 *
0-
02
b110 6
#39810000000
1!
1%
1-
12
#39820000000
0!
0%
b111 *
0-
02
b111 6
#39830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#39840000000
0!
0%
b0 *
0-
02
b0 6
#39850000000
1!
1%
1-
12
#39860000000
0!
0%
b1 *
0-
02
b1 6
#39870000000
1!
1%
1-
12
#39880000000
0!
0%
b10 *
0-
02
b10 6
#39890000000
1!
1%
1-
12
#39900000000
0!
0%
b11 *
0-
02
b11 6
#39910000000
1!
1%
1-
12
15
#39920000000
0!
0%
b100 *
0-
02
b100 6
#39930000000
1!
1%
1-
12
#39940000000
0!
0%
b101 *
0-
02
b101 6
#39950000000
1!
1%
1-
12
#39960000000
0!
0%
b110 *
0-
02
b110 6
#39970000000
1!
1%
1-
12
#39980000000
0!
0%
b111 *
0-
02
b111 6
#39990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#40000000000
0!
0%
b0 *
0-
02
b0 6
#40010000000
1!
1%
1-
12
#40020000000
0!
0%
b1 *
0-
02
b1 6
#40030000000
1!
1%
1-
12
#40040000000
0!
0%
b10 *
0-
02
b10 6
#40050000000
1!
1%
1-
12
#40060000000
0!
0%
b11 *
0-
02
b11 6
#40070000000
1!
1%
1-
12
15
#40080000000
0!
0%
b100 *
0-
02
b100 6
#40090000000
1!
1%
1-
12
#40100000000
0!
0%
b101 *
0-
02
b101 6
#40110000000
1!
1%
1-
12
#40120000000
0!
0%
b110 *
0-
02
b110 6
#40130000000
1!
1%
1-
12
#40140000000
0!
0%
b111 *
0-
02
b111 6
#40150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#40160000000
0!
0%
b0 *
0-
02
b0 6
#40170000000
1!
1%
1-
12
#40180000000
0!
0%
b1 *
0-
02
b1 6
#40190000000
1!
1%
1-
12
#40200000000
0!
0%
b10 *
0-
02
b10 6
#40210000000
1!
1%
1-
12
#40220000000
0!
0%
b11 *
0-
02
b11 6
#40230000000
1!
1%
1-
12
15
#40240000000
0!
0%
b100 *
0-
02
b100 6
#40250000000
1!
1%
1-
12
#40260000000
0!
0%
b101 *
0-
02
b101 6
#40270000000
1!
1%
1-
12
#40280000000
0!
0%
b110 *
0-
02
b110 6
#40290000000
1!
1%
1-
12
#40300000000
0!
0%
b111 *
0-
02
b111 6
#40310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#40320000000
0!
0%
b0 *
0-
02
b0 6
#40330000000
1!
1%
1-
12
#40340000000
0!
0%
b1 *
0-
02
b1 6
#40350000000
1!
1%
1-
12
#40360000000
0!
0%
b10 *
0-
02
b10 6
#40370000000
1!
1%
1-
12
#40380000000
0!
0%
b11 *
0-
02
b11 6
#40390000000
1!
1%
1-
12
15
#40400000000
0!
0%
b100 *
0-
02
b100 6
#40410000000
1!
1%
1-
12
#40420000000
0!
0%
b101 *
0-
02
b101 6
#40430000000
1!
1%
1-
12
#40440000000
0!
0%
b110 *
0-
02
b110 6
#40450000000
1!
1%
1-
12
#40460000000
0!
0%
b111 *
0-
02
b111 6
#40470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#40480000000
0!
0%
b0 *
0-
02
b0 6
#40490000000
1!
1%
1-
12
#40500000000
0!
0%
b1 *
0-
02
b1 6
#40510000000
1!
1%
1-
12
#40520000000
0!
0%
b10 *
0-
02
b10 6
#40530000000
1!
1%
1-
12
#40540000000
0!
0%
b11 *
0-
02
b11 6
#40550000000
1!
1%
1-
12
15
#40560000000
0!
0%
b100 *
0-
02
b100 6
#40570000000
1!
1%
1-
12
#40580000000
0!
0%
b101 *
0-
02
b101 6
#40590000000
1!
1%
1-
12
#40600000000
0!
0%
b110 *
0-
02
b110 6
#40610000000
1!
1%
1-
12
#40620000000
0!
0%
b111 *
0-
02
b111 6
#40630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#40640000000
0!
0%
b0 *
0-
02
b0 6
#40650000000
1!
1%
1-
12
#40660000000
0!
0%
b1 *
0-
02
b1 6
#40670000000
1!
1%
1-
12
#40680000000
0!
0%
b10 *
0-
02
b10 6
#40690000000
1!
1%
1-
12
#40700000000
0!
0%
b11 *
0-
02
b11 6
#40710000000
1!
1%
1-
12
15
#40720000000
0!
0%
b100 *
0-
02
b100 6
#40730000000
1!
1%
1-
12
#40740000000
0!
0%
b101 *
0-
02
b101 6
#40750000000
1!
1%
1-
12
#40760000000
0!
0%
b110 *
0-
02
b110 6
#40770000000
1!
1%
1-
12
#40780000000
0!
0%
b111 *
0-
02
b111 6
#40790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#40800000000
0!
0%
b0 *
0-
02
b0 6
#40810000000
1!
1%
1-
12
#40820000000
0!
0%
b1 *
0-
02
b1 6
#40830000000
1!
1%
1-
12
#40840000000
0!
0%
b10 *
0-
02
b10 6
#40850000000
1!
1%
1-
12
#40860000000
0!
0%
b11 *
0-
02
b11 6
#40870000000
1!
1%
1-
12
15
#40880000000
0!
0%
b100 *
0-
02
b100 6
#40890000000
1!
1%
1-
12
#40900000000
0!
0%
b101 *
0-
02
b101 6
#40910000000
1!
1%
1-
12
#40920000000
0!
0%
b110 *
0-
02
b110 6
#40930000000
1!
1%
1-
12
#40940000000
0!
0%
b111 *
0-
02
b111 6
#40950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#40960000000
0!
0%
b0 *
0-
02
b0 6
#40970000000
1!
1%
1-
12
#40980000000
0!
0%
b1 *
0-
02
b1 6
#40990000000
1!
1%
1-
12
#41000000000
0!
0%
b10 *
0-
02
b10 6
#41010000000
1!
1%
1-
12
#41020000000
0!
0%
b11 *
0-
02
b11 6
#41030000000
1!
1%
1-
12
15
#41040000000
0!
0%
b100 *
0-
02
b100 6
#41050000000
1!
1%
1-
12
#41060000000
0!
0%
b101 *
0-
02
b101 6
#41070000000
1!
1%
1-
12
#41080000000
0!
0%
b110 *
0-
02
b110 6
#41090000000
1!
1%
1-
12
#41100000000
0!
0%
b111 *
0-
02
b111 6
#41110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#41120000000
0!
0%
b0 *
0-
02
b0 6
#41130000000
1!
1%
1-
12
#41140000000
0!
0%
b1 *
0-
02
b1 6
#41150000000
1!
1%
1-
12
#41160000000
0!
0%
b10 *
0-
02
b10 6
#41170000000
1!
1%
1-
12
#41180000000
0!
0%
b11 *
0-
02
b11 6
#41190000000
1!
1%
1-
12
15
#41200000000
0!
0%
b100 *
0-
02
b100 6
#41210000000
1!
1%
1-
12
#41220000000
0!
0%
b101 *
0-
02
b101 6
#41230000000
1!
1%
1-
12
#41240000000
0!
0%
b110 *
0-
02
b110 6
#41250000000
1!
1%
1-
12
#41260000000
0!
0%
b111 *
0-
02
b111 6
#41270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#41280000000
0!
0%
b0 *
0-
02
b0 6
#41290000000
1!
1%
1-
12
#41300000000
0!
0%
b1 *
0-
02
b1 6
#41310000000
1!
1%
1-
12
#41320000000
0!
0%
b10 *
0-
02
b10 6
#41330000000
1!
1%
1-
12
#41340000000
0!
0%
b11 *
0-
02
b11 6
#41350000000
1!
1%
1-
12
15
#41360000000
0!
0%
b100 *
0-
02
b100 6
#41370000000
1!
1%
1-
12
#41380000000
0!
0%
b101 *
0-
02
b101 6
#41390000000
1!
1%
1-
12
#41400000000
0!
0%
b110 *
0-
02
b110 6
#41410000000
1!
1%
1-
12
#41420000000
0!
0%
b111 *
0-
02
b111 6
#41430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#41440000000
0!
0%
b0 *
0-
02
b0 6
#41450000000
1!
1%
1-
12
#41460000000
0!
0%
b1 *
0-
02
b1 6
#41470000000
1!
1%
1-
12
#41480000000
0!
0%
b10 *
0-
02
b10 6
#41490000000
1!
1%
1-
12
#41500000000
0!
0%
b11 *
0-
02
b11 6
#41510000000
1!
1%
1-
12
15
#41520000000
0!
0%
b100 *
0-
02
b100 6
#41530000000
1!
1%
1-
12
#41540000000
0!
0%
b101 *
0-
02
b101 6
#41550000000
1!
1%
1-
12
#41560000000
0!
0%
b110 *
0-
02
b110 6
#41570000000
1!
1%
1-
12
#41580000000
0!
0%
b111 *
0-
02
b111 6
#41590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#41600000000
0!
0%
b0 *
0-
02
b0 6
#41610000000
1!
1%
1-
12
#41620000000
0!
0%
b1 *
0-
02
b1 6
#41630000000
1!
1%
1-
12
#41640000000
0!
0%
b10 *
0-
02
b10 6
#41650000000
1!
1%
1-
12
#41660000000
0!
0%
b11 *
0-
02
b11 6
#41670000000
1!
1%
1-
12
15
#41680000000
0!
0%
b100 *
0-
02
b100 6
#41690000000
1!
1%
1-
12
#41700000000
0!
0%
b101 *
0-
02
b101 6
#41710000000
1!
1%
1-
12
#41720000000
0!
0%
b110 *
0-
02
b110 6
#41730000000
1!
1%
1-
12
#41740000000
0!
0%
b111 *
0-
02
b111 6
#41750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#41760000000
0!
0%
b0 *
0-
02
b0 6
#41770000000
1!
1%
1-
12
#41780000000
0!
0%
b1 *
0-
02
b1 6
#41790000000
1!
1%
1-
12
#41800000000
0!
0%
b10 *
0-
02
b10 6
#41810000000
1!
1%
1-
12
#41820000000
0!
0%
b11 *
0-
02
b11 6
#41830000000
1!
1%
1-
12
15
#41840000000
0!
0%
b100 *
0-
02
b100 6
#41850000000
1!
1%
1-
12
#41860000000
0!
0%
b101 *
0-
02
b101 6
#41870000000
1!
1%
1-
12
#41880000000
0!
0%
b110 *
0-
02
b110 6
#41890000000
1!
1%
1-
12
#41900000000
0!
0%
b111 *
0-
02
b111 6
#41910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#41920000000
0!
0%
b0 *
0-
02
b0 6
#41930000000
1!
1%
1-
12
#41940000000
0!
0%
b1 *
0-
02
b1 6
#41950000000
1!
1%
1-
12
#41960000000
0!
0%
b10 *
0-
02
b10 6
#41970000000
1!
1%
1-
12
#41980000000
0!
0%
b11 *
0-
02
b11 6
#41990000000
1!
1%
1-
12
15
#42000000000
0!
0%
b100 *
0-
02
b100 6
#42010000000
1!
1%
1-
12
#42020000000
0!
0%
b101 *
0-
02
b101 6
#42030000000
1!
1%
1-
12
#42040000000
0!
0%
b110 *
0-
02
b110 6
#42050000000
1!
1%
1-
12
#42060000000
0!
0%
b111 *
0-
02
b111 6
#42070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#42080000000
0!
0%
b0 *
0-
02
b0 6
#42090000000
1!
1%
1-
12
#42100000000
0!
0%
b1 *
0-
02
b1 6
#42110000000
1!
1%
1-
12
#42120000000
0!
0%
b10 *
0-
02
b10 6
#42130000000
1!
1%
1-
12
#42140000000
0!
0%
b11 *
0-
02
b11 6
#42150000000
1!
1%
1-
12
15
#42160000000
0!
0%
b100 *
0-
02
b100 6
#42170000000
1!
1%
1-
12
#42180000000
0!
0%
b101 *
0-
02
b101 6
#42190000000
1!
1%
1-
12
#42200000000
0!
0%
b110 *
0-
02
b110 6
#42210000000
1!
1%
1-
12
#42220000000
0!
0%
b111 *
0-
02
b111 6
#42230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#42240000000
0!
0%
b0 *
0-
02
b0 6
#42250000000
1!
1%
1-
12
#42260000000
0!
0%
b1 *
0-
02
b1 6
#42270000000
1!
1%
1-
12
#42280000000
0!
0%
b10 *
0-
02
b10 6
#42290000000
1!
1%
1-
12
#42300000000
0!
0%
b11 *
0-
02
b11 6
#42310000000
1!
1%
1-
12
15
#42320000000
0!
0%
b100 *
0-
02
b100 6
#42330000000
1!
1%
1-
12
#42340000000
0!
0%
b101 *
0-
02
b101 6
#42350000000
1!
1%
1-
12
#42360000000
0!
0%
b110 *
0-
02
b110 6
#42370000000
1!
1%
1-
12
#42380000000
0!
0%
b111 *
0-
02
b111 6
#42390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#42400000000
0!
0%
b0 *
0-
02
b0 6
#42410000000
1!
1%
1-
12
#42420000000
0!
0%
b1 *
0-
02
b1 6
#42430000000
1!
1%
1-
12
#42440000000
0!
0%
b10 *
0-
02
b10 6
#42450000000
1!
1%
1-
12
#42460000000
0!
0%
b11 *
0-
02
b11 6
#42470000000
1!
1%
1-
12
15
#42480000000
0!
0%
b100 *
0-
02
b100 6
#42490000000
1!
1%
1-
12
#42500000000
0!
0%
b101 *
0-
02
b101 6
#42510000000
1!
1%
1-
12
#42520000000
0!
0%
b110 *
0-
02
b110 6
#42530000000
1!
1%
1-
12
#42540000000
0!
0%
b111 *
0-
02
b111 6
#42550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#42560000000
0!
0%
b0 *
0-
02
b0 6
#42570000000
1!
1%
1-
12
#42580000000
0!
0%
b1 *
0-
02
b1 6
#42590000000
1!
1%
1-
12
#42600000000
0!
0%
b10 *
0-
02
b10 6
#42610000000
1!
1%
1-
12
#42620000000
0!
0%
b11 *
0-
02
b11 6
#42630000000
1!
1%
1-
12
15
#42640000000
0!
0%
b100 *
0-
02
b100 6
#42650000000
1!
1%
1-
12
#42660000000
0!
0%
b101 *
0-
02
b101 6
#42670000000
1!
1%
1-
12
#42680000000
0!
0%
b110 *
0-
02
b110 6
#42690000000
1!
1%
1-
12
#42700000000
0!
0%
b111 *
0-
02
b111 6
#42710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#42720000000
0!
0%
b0 *
0-
02
b0 6
#42730000000
1!
1%
1-
12
#42740000000
0!
0%
b1 *
0-
02
b1 6
#42750000000
1!
1%
1-
12
#42760000000
0!
0%
b10 *
0-
02
b10 6
#42770000000
1!
1%
1-
12
#42780000000
0!
0%
b11 *
0-
02
b11 6
#42790000000
1!
1%
1-
12
15
#42800000000
0!
0%
b100 *
0-
02
b100 6
#42810000000
1!
1%
1-
12
#42820000000
0!
0%
b101 *
0-
02
b101 6
#42830000000
1!
1%
1-
12
#42840000000
0!
0%
b110 *
0-
02
b110 6
#42850000000
1!
1%
1-
12
#42860000000
0!
0%
b111 *
0-
02
b111 6
#42870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#42880000000
0!
0%
b0 *
0-
02
b0 6
#42890000000
1!
1%
1-
12
#42900000000
0!
0%
b1 *
0-
02
b1 6
#42910000000
1!
1%
1-
12
#42920000000
0!
0%
b10 *
0-
02
b10 6
#42930000000
1!
1%
1-
12
#42940000000
0!
0%
b11 *
0-
02
b11 6
#42950000000
1!
1%
1-
12
15
#42960000000
0!
0%
b100 *
0-
02
b100 6
#42970000000
1!
1%
1-
12
#42980000000
0!
0%
b101 *
0-
02
b101 6
#42990000000
1!
1%
1-
12
#43000000000
0!
0%
b110 *
0-
02
b110 6
#43010000000
1!
1%
1-
12
#43020000000
0!
0%
b111 *
0-
02
b111 6
#43030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#43040000000
0!
0%
b0 *
0-
02
b0 6
#43050000000
1!
1%
1-
12
#43060000000
0!
0%
b1 *
0-
02
b1 6
#43070000000
1!
1%
1-
12
#43080000000
0!
0%
b10 *
0-
02
b10 6
#43090000000
1!
1%
1-
12
#43100000000
0!
0%
b11 *
0-
02
b11 6
#43110000000
1!
1%
1-
12
15
#43120000000
0!
0%
b100 *
0-
02
b100 6
#43130000000
1!
1%
1-
12
#43140000000
0!
0%
b101 *
0-
02
b101 6
#43150000000
1!
1%
1-
12
#43160000000
0!
0%
b110 *
0-
02
b110 6
#43170000000
1!
1%
1-
12
#43180000000
0!
0%
b111 *
0-
02
b111 6
#43190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#43200000000
0!
0%
b0 *
0-
02
b0 6
#43210000000
1!
1%
1-
12
#43220000000
0!
0%
b1 *
0-
02
b1 6
#43230000000
1!
1%
1-
12
#43240000000
0!
0%
b10 *
0-
02
b10 6
#43250000000
1!
1%
1-
12
#43260000000
0!
0%
b11 *
0-
02
b11 6
#43270000000
1!
1%
1-
12
15
#43280000000
0!
0%
b100 *
0-
02
b100 6
#43290000000
1!
1%
1-
12
#43300000000
0!
0%
b101 *
0-
02
b101 6
#43310000000
1!
1%
1-
12
#43320000000
0!
0%
b110 *
0-
02
b110 6
#43330000000
1!
1%
1-
12
#43340000000
0!
0%
b111 *
0-
02
b111 6
#43350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#43360000000
0!
0%
b0 *
0-
02
b0 6
#43370000000
1!
1%
1-
12
#43380000000
0!
0%
b1 *
0-
02
b1 6
#43390000000
1!
1%
1-
12
#43400000000
0!
0%
b10 *
0-
02
b10 6
#43410000000
1!
1%
1-
12
#43420000000
0!
0%
b11 *
0-
02
b11 6
#43430000000
1!
1%
1-
12
15
#43440000000
0!
0%
b100 *
0-
02
b100 6
#43450000000
1!
1%
1-
12
#43460000000
0!
0%
b101 *
0-
02
b101 6
#43470000000
1!
1%
1-
12
#43480000000
0!
0%
b110 *
0-
02
b110 6
#43490000000
1!
1%
1-
12
#43500000000
0!
0%
b111 *
0-
02
b111 6
#43510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#43520000000
0!
0%
b0 *
0-
02
b0 6
#43530000000
1!
1%
1-
12
#43540000000
0!
0%
b1 *
0-
02
b1 6
#43550000000
1!
1%
1-
12
#43560000000
0!
0%
b10 *
0-
02
b10 6
#43570000000
1!
1%
1-
12
#43580000000
0!
0%
b11 *
0-
02
b11 6
#43590000000
1!
1%
1-
12
15
#43600000000
0!
0%
b100 *
0-
02
b100 6
#43610000000
1!
1%
1-
12
#43620000000
0!
0%
b101 *
0-
02
b101 6
#43630000000
1!
1%
1-
12
#43640000000
0!
0%
b110 *
0-
02
b110 6
#43650000000
1!
1%
1-
12
#43660000000
0!
0%
b111 *
0-
02
b111 6
#43670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#43680000000
0!
0%
b0 *
0-
02
b0 6
#43690000000
1!
1%
1-
12
#43700000000
0!
0%
b1 *
0-
02
b1 6
#43710000000
1!
1%
1-
12
#43720000000
0!
0%
b10 *
0-
02
b10 6
#43730000000
1!
1%
1-
12
#43740000000
0!
0%
b11 *
0-
02
b11 6
#43750000000
1!
1%
1-
12
15
#43760000000
0!
0%
b100 *
0-
02
b100 6
#43770000000
1!
1%
1-
12
#43780000000
0!
0%
b101 *
0-
02
b101 6
#43790000000
1!
1%
1-
12
#43800000000
0!
0%
b110 *
0-
02
b110 6
#43810000000
1!
1%
1-
12
#43820000000
0!
0%
b111 *
0-
02
b111 6
#43830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#43840000000
0!
0%
b0 *
0-
02
b0 6
#43850000000
1!
1%
1-
12
#43860000000
0!
0%
b1 *
0-
02
b1 6
#43870000000
1!
1%
1-
12
#43880000000
0!
0%
b10 *
0-
02
b10 6
#43890000000
1!
1%
1-
12
#43900000000
0!
0%
b11 *
0-
02
b11 6
#43910000000
1!
1%
1-
12
15
#43920000000
0!
0%
b100 *
0-
02
b100 6
#43930000000
1!
1%
1-
12
#43940000000
0!
0%
b101 *
0-
02
b101 6
#43950000000
1!
1%
1-
12
#43960000000
0!
0%
b110 *
0-
02
b110 6
#43970000000
1!
1%
1-
12
#43980000000
0!
0%
b111 *
0-
02
b111 6
#43990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#44000000000
0!
0%
b0 *
0-
02
b0 6
#44010000000
1!
1%
1-
12
#44020000000
0!
0%
b1 *
0-
02
b1 6
#44030000000
1!
1%
1-
12
#44040000000
0!
0%
b10 *
0-
02
b10 6
#44050000000
1!
1%
1-
12
#44060000000
0!
0%
b11 *
0-
02
b11 6
#44070000000
1!
1%
1-
12
15
#44080000000
0!
0%
b100 *
0-
02
b100 6
#44090000000
1!
1%
1-
12
#44100000000
0!
0%
b101 *
0-
02
b101 6
#44110000000
1!
1%
1-
12
#44120000000
0!
0%
b110 *
0-
02
b110 6
#44130000000
1!
1%
1-
12
#44140000000
0!
0%
b111 *
0-
02
b111 6
#44150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#44160000000
0!
0%
b0 *
0-
02
b0 6
#44170000000
1!
1%
1-
12
#44180000000
0!
0%
b1 *
0-
02
b1 6
#44190000000
1!
1%
1-
12
#44200000000
0!
0%
b10 *
0-
02
b10 6
#44210000000
1!
1%
1-
12
#44220000000
0!
0%
b11 *
0-
02
b11 6
#44230000000
1!
1%
1-
12
15
#44240000000
0!
0%
b100 *
0-
02
b100 6
#44250000000
1!
1%
1-
12
#44260000000
0!
0%
b101 *
0-
02
b101 6
#44270000000
1!
1%
1-
12
#44280000000
0!
0%
b110 *
0-
02
b110 6
#44290000000
1!
1%
1-
12
#44300000000
0!
0%
b111 *
0-
02
b111 6
#44310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#44320000000
0!
0%
b0 *
0-
02
b0 6
#44330000000
1!
1%
1-
12
#44340000000
0!
0%
b1 *
0-
02
b1 6
#44350000000
1!
1%
1-
12
#44360000000
0!
0%
b10 *
0-
02
b10 6
#44370000000
1!
1%
1-
12
#44380000000
0!
0%
b11 *
0-
02
b11 6
#44390000000
1!
1%
1-
12
15
#44400000000
0!
0%
b100 *
0-
02
b100 6
#44410000000
1!
1%
1-
12
#44420000000
0!
0%
b101 *
0-
02
b101 6
#44430000000
1!
1%
1-
12
#44440000000
0!
0%
b110 *
0-
02
b110 6
#44450000000
1!
1%
1-
12
#44460000000
0!
0%
b111 *
0-
02
b111 6
#44470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#44480000000
0!
0%
b0 *
0-
02
b0 6
#44490000000
1!
1%
1-
12
#44500000000
0!
0%
b1 *
0-
02
b1 6
#44510000000
1!
1%
1-
12
#44520000000
0!
0%
b10 *
0-
02
b10 6
#44530000000
1!
1%
1-
12
#44540000000
0!
0%
b11 *
0-
02
b11 6
#44550000000
1!
1%
1-
12
15
#44560000000
0!
0%
b100 *
0-
02
b100 6
#44570000000
1!
1%
1-
12
#44580000000
0!
0%
b101 *
0-
02
b101 6
#44590000000
1!
1%
1-
12
#44600000000
0!
0%
b110 *
0-
02
b110 6
#44610000000
1!
1%
1-
12
#44620000000
0!
0%
b111 *
0-
02
b111 6
#44630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#44640000000
0!
0%
b0 *
0-
02
b0 6
#44650000000
1!
1%
1-
12
#44660000000
0!
0%
b1 *
0-
02
b1 6
#44670000000
1!
1%
1-
12
#44680000000
0!
0%
b10 *
0-
02
b10 6
#44690000000
1!
1%
1-
12
#44700000000
0!
0%
b11 *
0-
02
b11 6
#44710000000
1!
1%
1-
12
15
#44720000000
0!
0%
b100 *
0-
02
b100 6
#44730000000
1!
1%
1-
12
#44740000000
0!
0%
b101 *
0-
02
b101 6
#44750000000
1!
1%
1-
12
#44760000000
0!
0%
b110 *
0-
02
b110 6
#44770000000
1!
1%
1-
12
#44780000000
0!
0%
b111 *
0-
02
b111 6
#44790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#44800000000
0!
0%
b0 *
0-
02
b0 6
#44810000000
1!
1%
1-
12
#44820000000
0!
0%
b1 *
0-
02
b1 6
#44830000000
1!
1%
1-
12
#44840000000
0!
0%
b10 *
0-
02
b10 6
#44850000000
1!
1%
1-
12
#44860000000
0!
0%
b11 *
0-
02
b11 6
#44870000000
1!
1%
1-
12
15
#44880000000
0!
0%
b100 *
0-
02
b100 6
#44890000000
1!
1%
1-
12
#44900000000
0!
0%
b101 *
0-
02
b101 6
#44910000000
1!
1%
1-
12
#44920000000
0!
0%
b110 *
0-
02
b110 6
#44930000000
1!
1%
1-
12
#44940000000
0!
0%
b111 *
0-
02
b111 6
#44950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#44960000000
0!
0%
b0 *
0-
02
b0 6
#44970000000
1!
1%
1-
12
#44980000000
0!
0%
b1 *
0-
02
b1 6
#44990000000
1!
1%
1-
12
#45000000000
0!
0%
b10 *
0-
02
b10 6
#45010000000
1!
1%
1-
12
#45020000000
0!
0%
b11 *
0-
02
b11 6
#45030000000
1!
1%
1-
12
15
#45040000000
0!
0%
b100 *
0-
02
b100 6
#45050000000
1!
1%
1-
12
#45060000000
0!
0%
b101 *
0-
02
b101 6
#45070000000
1!
1%
1-
12
#45080000000
0!
0%
b110 *
0-
02
b110 6
#45090000000
1!
1%
1-
12
#45100000000
0!
0%
b111 *
0-
02
b111 6
#45110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#45120000000
0!
0%
b0 *
0-
02
b0 6
#45130000000
1!
1%
1-
12
#45140000000
0!
0%
b1 *
0-
02
b1 6
#45150000000
1!
1%
1-
12
#45160000000
0!
0%
b10 *
0-
02
b10 6
#45170000000
1!
1%
1-
12
#45180000000
0!
0%
b11 *
0-
02
b11 6
#45190000000
1!
1%
1-
12
15
#45200000000
0!
0%
b100 *
0-
02
b100 6
#45210000000
1!
1%
1-
12
#45220000000
0!
0%
b101 *
0-
02
b101 6
#45230000000
1!
1%
1-
12
#45240000000
0!
0%
b110 *
0-
02
b110 6
#45250000000
1!
1%
1-
12
#45260000000
0!
0%
b111 *
0-
02
b111 6
#45270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#45280000000
0!
0%
b0 *
0-
02
b0 6
#45290000000
1!
1%
1-
12
#45300000000
0!
0%
b1 *
0-
02
b1 6
#45310000000
1!
1%
1-
12
#45320000000
0!
0%
b10 *
0-
02
b10 6
#45330000000
1!
1%
1-
12
#45340000000
0!
0%
b11 *
0-
02
b11 6
#45350000000
1!
1%
1-
12
15
#45360000000
0!
0%
b100 *
0-
02
b100 6
#45370000000
1!
1%
1-
12
#45380000000
0!
0%
b101 *
0-
02
b101 6
#45390000000
1!
1%
1-
12
#45400000000
0!
0%
b110 *
0-
02
b110 6
#45410000000
1!
1%
1-
12
#45420000000
0!
0%
b111 *
0-
02
b111 6
#45430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#45440000000
0!
0%
b0 *
0-
02
b0 6
#45450000000
1!
1%
1-
12
#45460000000
0!
0%
b1 *
0-
02
b1 6
#45470000000
1!
1%
1-
12
#45480000000
0!
0%
b10 *
0-
02
b10 6
#45490000000
1!
1%
1-
12
#45500000000
0!
0%
b11 *
0-
02
b11 6
#45510000000
1!
1%
1-
12
15
#45520000000
0!
0%
b100 *
0-
02
b100 6
#45530000000
1!
1%
1-
12
#45540000000
0!
0%
b101 *
0-
02
b101 6
#45550000000
1!
1%
1-
12
#45560000000
0!
0%
b110 *
0-
02
b110 6
#45570000000
1!
1%
1-
12
#45580000000
0!
0%
b111 *
0-
02
b111 6
#45590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#45600000000
0!
0%
b0 *
0-
02
b0 6
#45610000000
1!
1%
1-
12
#45620000000
0!
0%
b1 *
0-
02
b1 6
#45630000000
1!
1%
1-
12
#45640000000
0!
0%
b10 *
0-
02
b10 6
#45650000000
1!
1%
1-
12
#45660000000
0!
0%
b11 *
0-
02
b11 6
#45670000000
1!
1%
1-
12
15
#45680000000
0!
0%
b100 *
0-
02
b100 6
#45690000000
1!
1%
1-
12
#45700000000
0!
0%
b101 *
0-
02
b101 6
#45710000000
1!
1%
1-
12
#45720000000
0!
0%
b110 *
0-
02
b110 6
#45730000000
1!
1%
1-
12
#45740000000
0!
0%
b111 *
0-
02
b111 6
#45750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#45760000000
0!
0%
b0 *
0-
02
b0 6
#45770000000
1!
1%
1-
12
#45780000000
0!
0%
b1 *
0-
02
b1 6
#45790000000
1!
1%
1-
12
#45800000000
0!
0%
b10 *
0-
02
b10 6
#45810000000
1!
1%
1-
12
#45820000000
0!
0%
b11 *
0-
02
b11 6
#45830000000
1!
1%
1-
12
15
#45840000000
0!
0%
b100 *
0-
02
b100 6
#45850000000
1!
1%
1-
12
#45860000000
0!
0%
b101 *
0-
02
b101 6
#45870000000
1!
1%
1-
12
#45880000000
0!
0%
b110 *
0-
02
b110 6
#45890000000
1!
1%
1-
12
#45900000000
0!
0%
b111 *
0-
02
b111 6
#45910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#45920000000
0!
0%
b0 *
0-
02
b0 6
#45930000000
1!
1%
1-
12
#45940000000
0!
0%
b1 *
0-
02
b1 6
#45950000000
1!
1%
1-
12
#45960000000
0!
0%
b10 *
0-
02
b10 6
#45970000000
1!
1%
1-
12
#45980000000
0!
0%
b11 *
0-
02
b11 6
#45990000000
1!
1%
1-
12
15
#46000000000
0!
0%
b100 *
0-
02
b100 6
#46010000000
1!
1%
1-
12
#46020000000
0!
0%
b101 *
0-
02
b101 6
#46030000000
1!
1%
1-
12
#46040000000
0!
0%
b110 *
0-
02
b110 6
#46050000000
1!
1%
1-
12
#46060000000
0!
0%
b111 *
0-
02
b111 6
#46070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#46080000000
0!
0%
b0 *
0-
02
b0 6
#46090000000
1!
1%
1-
12
#46100000000
0!
0%
b1 *
0-
02
b1 6
#46110000000
1!
1%
1-
12
#46120000000
0!
0%
b10 *
0-
02
b10 6
#46130000000
1!
1%
1-
12
#46140000000
0!
0%
b11 *
0-
02
b11 6
#46150000000
1!
1%
1-
12
15
#46160000000
0!
0%
b100 *
0-
02
b100 6
#46170000000
1!
1%
1-
12
#46180000000
0!
0%
b101 *
0-
02
b101 6
#46190000000
1!
1%
1-
12
#46200000000
0!
0%
b110 *
0-
02
b110 6
#46210000000
1!
1%
1-
12
#46220000000
0!
0%
b111 *
0-
02
b111 6
#46230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#46240000000
0!
0%
b0 *
0-
02
b0 6
#46250000000
1!
1%
1-
12
#46260000000
0!
0%
b1 *
0-
02
b1 6
#46270000000
1!
1%
1-
12
#46280000000
0!
0%
b10 *
0-
02
b10 6
#46290000000
1!
1%
1-
12
#46300000000
0!
0%
b11 *
0-
02
b11 6
#46310000000
1!
1%
1-
12
15
#46320000000
0!
0%
b100 *
0-
02
b100 6
#46330000000
1!
1%
1-
12
#46340000000
0!
0%
b101 *
0-
02
b101 6
#46350000000
1!
1%
1-
12
#46360000000
0!
0%
b110 *
0-
02
b110 6
#46370000000
1!
1%
1-
12
#46380000000
0!
0%
b111 *
0-
02
b111 6
#46390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#46400000000
0!
0%
b0 *
0-
02
b0 6
#46410000000
1!
1%
1-
12
#46420000000
0!
0%
b1 *
0-
02
b1 6
#46430000000
1!
1%
1-
12
#46440000000
0!
0%
b10 *
0-
02
b10 6
#46450000000
1!
1%
1-
12
#46460000000
0!
0%
b11 *
0-
02
b11 6
#46470000000
1!
1%
1-
12
15
#46480000000
0!
0%
b100 *
0-
02
b100 6
#46490000000
1!
1%
1-
12
#46500000000
0!
0%
b101 *
0-
02
b101 6
#46510000000
1!
1%
1-
12
#46520000000
0!
0%
b110 *
0-
02
b110 6
#46530000000
1!
1%
1-
12
#46540000000
0!
0%
b111 *
0-
02
b111 6
#46550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#46560000000
0!
0%
b0 *
0-
02
b0 6
#46570000000
1!
1%
1-
12
#46580000000
0!
0%
b1 *
0-
02
b1 6
#46590000000
1!
1%
1-
12
#46600000000
0!
0%
b10 *
0-
02
b10 6
#46610000000
1!
1%
1-
12
#46620000000
0!
0%
b11 *
0-
02
b11 6
#46630000000
1!
1%
1-
12
15
#46640000000
0!
0%
b100 *
0-
02
b100 6
#46650000000
1!
1%
1-
12
#46660000000
0!
0%
b101 *
0-
02
b101 6
#46670000000
1!
1%
1-
12
#46680000000
0!
0%
b110 *
0-
02
b110 6
#46690000000
1!
1%
1-
12
#46700000000
0!
0%
b111 *
0-
02
b111 6
#46710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#46720000000
0!
0%
b0 *
0-
02
b0 6
#46730000000
1!
1%
1-
12
#46740000000
0!
0%
b1 *
0-
02
b1 6
#46750000000
1!
1%
1-
12
#46760000000
0!
0%
b10 *
0-
02
b10 6
#46770000000
1!
1%
1-
12
#46780000000
0!
0%
b11 *
0-
02
b11 6
#46790000000
1!
1%
1-
12
15
#46800000000
0!
0%
b100 *
0-
02
b100 6
#46810000000
1!
1%
1-
12
#46820000000
0!
0%
b101 *
0-
02
b101 6
#46830000000
1!
1%
1-
12
#46840000000
0!
0%
b110 *
0-
02
b110 6
#46850000000
1!
1%
1-
12
#46860000000
0!
0%
b111 *
0-
02
b111 6
#46870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#46880000000
0!
0%
b0 *
0-
02
b0 6
#46890000000
1!
1%
1-
12
#46900000000
0!
0%
b1 *
0-
02
b1 6
#46910000000
1!
1%
1-
12
#46920000000
0!
0%
b10 *
0-
02
b10 6
#46930000000
1!
1%
1-
12
#46940000000
0!
0%
b11 *
0-
02
b11 6
#46950000000
1!
1%
1-
12
15
#46960000000
0!
0%
b100 *
0-
02
b100 6
#46970000000
1!
1%
1-
12
#46980000000
0!
0%
b101 *
0-
02
b101 6
#46990000000
1!
1%
1-
12
#47000000000
0!
0%
b110 *
0-
02
b110 6
#47010000000
1!
1%
1-
12
#47020000000
0!
0%
b111 *
0-
02
b111 6
#47030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#47040000000
0!
0%
b0 *
0-
02
b0 6
#47050000000
1!
1%
1-
12
#47060000000
0!
0%
b1 *
0-
02
b1 6
#47070000000
1!
1%
1-
12
#47080000000
0!
0%
b10 *
0-
02
b10 6
#47090000000
1!
1%
1-
12
#47100000000
0!
0%
b11 *
0-
02
b11 6
#47110000000
1!
1%
1-
12
15
#47120000000
0!
0%
b100 *
0-
02
b100 6
#47130000000
1!
1%
1-
12
#47140000000
0!
0%
b101 *
0-
02
b101 6
#47150000000
1!
1%
1-
12
#47160000000
0!
0%
b110 *
0-
02
b110 6
#47170000000
1!
1%
1-
12
#47180000000
0!
0%
b111 *
0-
02
b111 6
#47190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#47200000000
0!
0%
b0 *
0-
02
b0 6
#47210000000
1!
1%
1-
12
#47220000000
0!
0%
b1 *
0-
02
b1 6
#47230000000
1!
1%
1-
12
#47240000000
0!
0%
b10 *
0-
02
b10 6
#47250000000
1!
1%
1-
12
#47260000000
0!
0%
b11 *
0-
02
b11 6
#47270000000
1!
1%
1-
12
15
#47280000000
0!
0%
b100 *
0-
02
b100 6
#47290000000
1!
1%
1-
12
#47300000000
0!
0%
b101 *
0-
02
b101 6
#47310000000
1!
1%
1-
12
#47320000000
0!
0%
b110 *
0-
02
b110 6
#47330000000
1!
1%
1-
12
#47340000000
0!
0%
b111 *
0-
02
b111 6
#47350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#47360000000
0!
0%
b0 *
0-
02
b0 6
#47370000000
1!
1%
1-
12
#47380000000
0!
0%
b1 *
0-
02
b1 6
#47390000000
1!
1%
1-
12
#47400000000
0!
0%
b10 *
0-
02
b10 6
#47410000000
1!
1%
1-
12
#47420000000
0!
0%
b11 *
0-
02
b11 6
#47430000000
1!
1%
1-
12
15
#47440000000
0!
0%
b100 *
0-
02
b100 6
#47450000000
1!
1%
1-
12
#47460000000
0!
0%
b101 *
0-
02
b101 6
#47470000000
1!
1%
1-
12
#47480000000
0!
0%
b110 *
0-
02
b110 6
#47490000000
1!
1%
1-
12
#47500000000
0!
0%
b111 *
0-
02
b111 6
#47510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#47520000000
0!
0%
b0 *
0-
02
b0 6
#47530000000
1!
1%
1-
12
#47540000000
0!
0%
b1 *
0-
02
b1 6
#47550000000
1!
1%
1-
12
#47560000000
0!
0%
b10 *
0-
02
b10 6
#47570000000
1!
1%
1-
12
#47580000000
0!
0%
b11 *
0-
02
b11 6
#47590000000
1!
1%
1-
12
15
#47600000000
0!
0%
b100 *
0-
02
b100 6
#47610000000
1!
1%
1-
12
#47620000000
0!
0%
b101 *
0-
02
b101 6
#47630000000
1!
1%
1-
12
#47640000000
0!
0%
b110 *
0-
02
b110 6
#47650000000
1!
1%
1-
12
#47660000000
0!
0%
b111 *
0-
02
b111 6
#47670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#47680000000
0!
0%
b0 *
0-
02
b0 6
#47690000000
1!
1%
1-
12
#47700000000
0!
0%
b1 *
0-
02
b1 6
#47710000000
1!
1%
1-
12
#47720000000
0!
0%
b10 *
0-
02
b10 6
#47730000000
1!
1%
1-
12
#47740000000
0!
0%
b11 *
0-
02
b11 6
#47750000000
1!
1%
1-
12
15
#47760000000
0!
0%
b100 *
0-
02
b100 6
#47770000000
1!
1%
1-
12
#47780000000
0!
0%
b101 *
0-
02
b101 6
#47790000000
1!
1%
1-
12
#47800000000
0!
0%
b110 *
0-
02
b110 6
#47810000000
1!
1%
1-
12
#47820000000
0!
0%
b111 *
0-
02
b111 6
#47830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#47840000000
0!
0%
b0 *
0-
02
b0 6
#47850000000
1!
1%
1-
12
#47860000000
0!
0%
b1 *
0-
02
b1 6
#47870000000
1!
1%
1-
12
#47880000000
0!
0%
b10 *
0-
02
b10 6
#47890000000
1!
1%
1-
12
#47900000000
0!
0%
b11 *
0-
02
b11 6
#47910000000
1!
1%
1-
12
15
#47920000000
0!
0%
b100 *
0-
02
b100 6
#47930000000
1!
1%
1-
12
#47940000000
0!
0%
b101 *
0-
02
b101 6
#47950000000
1!
1%
1-
12
#47960000000
0!
0%
b110 *
0-
02
b110 6
#47970000000
1!
1%
1-
12
#47980000000
0!
0%
b111 *
0-
02
b111 6
#47990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#48000000000
0!
0%
b0 *
0-
02
b0 6
#48010000000
1!
1%
1-
12
#48020000000
0!
0%
b1 *
0-
02
b1 6
#48030000000
1!
1%
1-
12
#48040000000
0!
0%
b10 *
0-
02
b10 6
#48050000000
1!
1%
1-
12
#48060000000
0!
0%
b11 *
0-
02
b11 6
#48070000000
1!
1%
1-
12
15
#48080000000
0!
0%
b100 *
0-
02
b100 6
#48090000000
1!
1%
1-
12
#48100000000
0!
0%
b101 *
0-
02
b101 6
#48110000000
1!
1%
1-
12
#48120000000
0!
0%
b110 *
0-
02
b110 6
#48130000000
1!
1%
1-
12
#48140000000
0!
0%
b111 *
0-
02
b111 6
#48150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#48160000000
0!
0%
b0 *
0-
02
b0 6
#48170000000
1!
1%
1-
12
#48180000000
0!
0%
b1 *
0-
02
b1 6
#48190000000
1!
1%
1-
12
#48200000000
0!
0%
b10 *
0-
02
b10 6
#48210000000
1!
1%
1-
12
#48220000000
0!
0%
b11 *
0-
02
b11 6
#48230000000
1!
1%
1-
12
15
#48240000000
0!
0%
b100 *
0-
02
b100 6
#48250000000
1!
1%
1-
12
#48260000000
0!
0%
b101 *
0-
02
b101 6
#48270000000
1!
1%
1-
12
#48280000000
0!
0%
b110 *
0-
02
b110 6
#48290000000
1!
1%
1-
12
#48300000000
0!
0%
b111 *
0-
02
b111 6
#48310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#48320000000
0!
0%
b0 *
0-
02
b0 6
#48330000000
1!
1%
1-
12
#48340000000
0!
0%
b1 *
0-
02
b1 6
#48350000000
1!
1%
1-
12
#48360000000
0!
0%
b10 *
0-
02
b10 6
#48370000000
1!
1%
1-
12
#48380000000
0!
0%
b11 *
0-
02
b11 6
#48390000000
1!
1%
1-
12
15
#48400000000
0!
0%
b100 *
0-
02
b100 6
#48410000000
1!
1%
1-
12
#48420000000
0!
0%
b101 *
0-
02
b101 6
#48430000000
1!
1%
1-
12
#48440000000
0!
0%
b110 *
0-
02
b110 6
#48450000000
1!
1%
1-
12
#48460000000
0!
0%
b111 *
0-
02
b111 6
#48470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#48480000000
0!
0%
b0 *
0-
02
b0 6
#48490000000
1!
1%
1-
12
#48500000000
0!
0%
b1 *
0-
02
b1 6
#48510000000
1!
1%
1-
12
#48520000000
0!
0%
b10 *
0-
02
b10 6
#48530000000
1!
1%
1-
12
#48540000000
0!
0%
b11 *
0-
02
b11 6
#48550000000
1!
1%
1-
12
15
#48560000000
0!
0%
b100 *
0-
02
b100 6
#48570000000
1!
1%
1-
12
#48580000000
0!
0%
b101 *
0-
02
b101 6
#48590000000
1!
1%
1-
12
#48600000000
0!
0%
b110 *
0-
02
b110 6
#48610000000
1!
1%
1-
12
#48620000000
0!
0%
b111 *
0-
02
b111 6
#48630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#48640000000
0!
0%
b0 *
0-
02
b0 6
#48650000000
1!
1%
1-
12
#48660000000
0!
0%
b1 *
0-
02
b1 6
#48670000000
1!
1%
1-
12
#48680000000
0!
0%
b10 *
0-
02
b10 6
#48690000000
1!
1%
1-
12
#48700000000
0!
0%
b11 *
0-
02
b11 6
#48710000000
1!
1%
1-
12
15
#48720000000
0!
0%
b100 *
0-
02
b100 6
#48730000000
1!
1%
1-
12
#48740000000
0!
0%
b101 *
0-
02
b101 6
#48750000000
1!
1%
1-
12
#48760000000
0!
0%
b110 *
0-
02
b110 6
#48770000000
1!
1%
1-
12
#48780000000
0!
0%
b111 *
0-
02
b111 6
#48790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#48800000000
0!
0%
b0 *
0-
02
b0 6
#48810000000
1!
1%
1-
12
#48820000000
0!
0%
b1 *
0-
02
b1 6
#48830000000
1!
1%
1-
12
#48840000000
0!
0%
b10 *
0-
02
b10 6
#48850000000
1!
1%
1-
12
#48860000000
0!
0%
b11 *
0-
02
b11 6
#48870000000
1!
1%
1-
12
15
#48880000000
0!
0%
b100 *
0-
02
b100 6
#48890000000
1!
1%
1-
12
#48900000000
0!
0%
b101 *
0-
02
b101 6
#48910000000
1!
1%
1-
12
#48920000000
0!
0%
b110 *
0-
02
b110 6
#48930000000
1!
1%
1-
12
#48940000000
0!
0%
b111 *
0-
02
b111 6
#48950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#48960000000
0!
0%
b0 *
0-
02
b0 6
#48970000000
1!
1%
1-
12
#48980000000
0!
0%
b1 *
0-
02
b1 6
#48990000000
1!
1%
1-
12
#49000000000
0!
0%
b10 *
0-
02
b10 6
#49010000000
1!
1%
1-
12
#49020000000
0!
0%
b11 *
0-
02
b11 6
#49030000000
1!
1%
1-
12
15
#49040000000
0!
0%
b100 *
0-
02
b100 6
#49050000000
1!
1%
1-
12
#49060000000
0!
0%
b101 *
0-
02
b101 6
#49070000000
1!
1%
1-
12
#49080000000
0!
0%
b110 *
0-
02
b110 6
#49090000000
1!
1%
1-
12
#49100000000
0!
0%
b111 *
0-
02
b111 6
#49110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#49120000000
0!
0%
b0 *
0-
02
b0 6
#49130000000
1!
1%
1-
12
#49140000000
0!
0%
b1 *
0-
02
b1 6
#49150000000
1!
1%
1-
12
#49160000000
0!
0%
b10 *
0-
02
b10 6
#49170000000
1!
1%
1-
12
#49180000000
0!
0%
b11 *
0-
02
b11 6
#49190000000
1!
1%
1-
12
15
#49200000000
0!
0%
b100 *
0-
02
b100 6
#49210000000
1!
1%
1-
12
#49220000000
0!
0%
b101 *
0-
02
b101 6
#49230000000
1!
1%
1-
12
#49240000000
0!
0%
b110 *
0-
02
b110 6
#49250000000
1!
1%
1-
12
#49260000000
0!
0%
b111 *
0-
02
b111 6
#49270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#49280000000
0!
0%
b0 *
0-
02
b0 6
#49290000000
1!
1%
1-
12
#49300000000
0!
0%
b1 *
0-
02
b1 6
#49310000000
1!
1%
1-
12
#49320000000
0!
0%
b10 *
0-
02
b10 6
#49330000000
1!
1%
1-
12
#49340000000
0!
0%
b11 *
0-
02
b11 6
#49350000000
1!
1%
1-
12
15
#49360000000
0!
0%
b100 *
0-
02
b100 6
#49370000000
1!
1%
1-
12
#49380000000
0!
0%
b101 *
0-
02
b101 6
#49390000000
1!
1%
1-
12
#49400000000
0!
0%
b110 *
0-
02
b110 6
#49410000000
1!
1%
1-
12
#49420000000
0!
0%
b111 *
0-
02
b111 6
#49430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#49440000000
0!
0%
b0 *
0-
02
b0 6
#49450000000
1!
1%
1-
12
#49460000000
0!
0%
b1 *
0-
02
b1 6
#49470000000
1!
1%
1-
12
#49480000000
0!
0%
b10 *
0-
02
b10 6
#49490000000
1!
1%
1-
12
#49500000000
0!
0%
b11 *
0-
02
b11 6
#49510000000
1!
1%
1-
12
15
#49520000000
0!
0%
b100 *
0-
02
b100 6
#49530000000
1!
1%
1-
12
#49540000000
0!
0%
b101 *
0-
02
b101 6
#49550000000
1!
1%
1-
12
#49560000000
0!
0%
b110 *
0-
02
b110 6
#49570000000
1!
1%
1-
12
#49580000000
0!
0%
b111 *
0-
02
b111 6
#49590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#49600000000
0!
0%
b0 *
0-
02
b0 6
#49610000000
1!
1%
1-
12
#49620000000
0!
0%
b1 *
0-
02
b1 6
#49630000000
1!
1%
1-
12
#49640000000
0!
0%
b10 *
0-
02
b10 6
#49650000000
1!
1%
1-
12
#49660000000
0!
0%
b11 *
0-
02
b11 6
#49670000000
1!
1%
1-
12
15
#49680000000
0!
0%
b100 *
0-
02
b100 6
#49690000000
1!
1%
1-
12
#49700000000
0!
0%
b101 *
0-
02
b101 6
#49710000000
1!
1%
1-
12
#49720000000
0!
0%
b110 *
0-
02
b110 6
#49730000000
1!
1%
1-
12
#49740000000
0!
0%
b111 *
0-
02
b111 6
#49750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#49760000000
0!
0%
b0 *
0-
02
b0 6
#49770000000
1!
1%
1-
12
#49780000000
0!
0%
b1 *
0-
02
b1 6
#49790000000
1!
1%
1-
12
#49800000000
0!
0%
b10 *
0-
02
b10 6
#49810000000
1!
1%
1-
12
#49820000000
0!
0%
b11 *
0-
02
b11 6
#49830000000
1!
1%
1-
12
15
#49840000000
0!
0%
b100 *
0-
02
b100 6
#49850000000
1!
1%
1-
12
#49860000000
0!
0%
b101 *
0-
02
b101 6
#49870000000
1!
1%
1-
12
#49880000000
0!
0%
b110 *
0-
02
b110 6
#49890000000
1!
1%
1-
12
#49900000000
0!
0%
b111 *
0-
02
b111 6
#49910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#49920000000
0!
0%
b0 *
0-
02
b0 6
#49930000000
1!
1%
1-
12
#49940000000
0!
0%
b1 *
0-
02
b1 6
#49950000000
1!
1%
1-
12
#49960000000
0!
0%
b10 *
0-
02
b10 6
#49970000000
1!
1%
1-
12
#49980000000
0!
0%
b11 *
0-
02
b11 6
#49990000000
1!
1%
1-
12
15
#50000000000
0!
0%
b100 *
0-
02
b100 6
#50010000000
1!
1%
1-
12
#50020000000
0!
0%
b101 *
0-
02
b101 6
#50030000000
1!
1%
1-
12
#50040000000
0!
0%
b110 *
0-
02
b110 6
#50050000000
1!
1%
1-
12
#50060000000
0!
0%
b111 *
0-
02
b111 6
#50070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#50080000000
0!
0%
b0 *
0-
02
b0 6
#50090000000
1!
1%
1-
12
#50100000000
0!
0%
b1 *
0-
02
b1 6
#50110000000
1!
1%
1-
12
#50120000000
0!
0%
b10 *
0-
02
b10 6
#50130000000
1!
1%
1-
12
#50140000000
0!
0%
b11 *
0-
02
b11 6
#50150000000
1!
1%
1-
12
15
#50160000000
0!
0%
b100 *
0-
02
b100 6
#50170000000
1!
1%
1-
12
#50180000000
0!
0%
b101 *
0-
02
b101 6
#50190000000
1!
1%
1-
12
#50200000000
0!
0%
b110 *
0-
02
b110 6
#50210000000
1!
1%
1-
12
#50220000000
0!
0%
b111 *
0-
02
b111 6
#50230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#50240000000
0!
0%
b0 *
0-
02
b0 6
#50250000000
1!
1%
1-
12
#50260000000
0!
0%
b1 *
0-
02
b1 6
#50270000000
1!
1%
1-
12
#50280000000
0!
0%
b10 *
0-
02
b10 6
#50290000000
1!
1%
1-
12
#50300000000
0!
0%
b11 *
0-
02
b11 6
#50310000000
1!
1%
1-
12
15
#50320000000
0!
0%
b100 *
0-
02
b100 6
#50330000000
1!
1%
1-
12
#50340000000
0!
0%
b101 *
0-
02
b101 6
#50350000000
1!
1%
1-
12
#50360000000
0!
0%
b110 *
0-
02
b110 6
#50370000000
1!
1%
1-
12
#50380000000
0!
0%
b111 *
0-
02
b111 6
#50390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#50400000000
0!
0%
b0 *
0-
02
b0 6
#50410000000
1!
1%
1-
12
#50420000000
0!
0%
b1 *
0-
02
b1 6
#50430000000
1!
1%
1-
12
#50440000000
0!
0%
b10 *
0-
02
b10 6
#50450000000
1!
1%
1-
12
#50460000000
0!
0%
b11 *
0-
02
b11 6
#50470000000
1!
1%
1-
12
15
#50480000000
0!
0%
b100 *
0-
02
b100 6
#50490000000
1!
1%
1-
12
#50500000000
0!
0%
b101 *
0-
02
b101 6
#50510000000
1!
1%
1-
12
#50520000000
0!
0%
b110 *
0-
02
b110 6
#50530000000
1!
1%
1-
12
#50540000000
0!
0%
b111 *
0-
02
b111 6
#50550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#50560000000
0!
0%
b0 *
0-
02
b0 6
#50570000000
1!
1%
1-
12
#50580000000
0!
0%
b1 *
0-
02
b1 6
#50590000000
1!
1%
1-
12
#50600000000
0!
0%
b10 *
0-
02
b10 6
#50610000000
1!
1%
1-
12
#50620000000
0!
0%
b11 *
0-
02
b11 6
#50630000000
1!
1%
1-
12
15
#50640000000
0!
0%
b100 *
0-
02
b100 6
#50650000000
1!
1%
1-
12
#50660000000
0!
0%
b101 *
0-
02
b101 6
#50670000000
1!
1%
1-
12
#50680000000
0!
0%
b110 *
0-
02
b110 6
#50690000000
1!
1%
1-
12
#50700000000
0!
0%
b111 *
0-
02
b111 6
#50710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#50720000000
0!
0%
b0 *
0-
02
b0 6
#50730000000
1!
1%
1-
12
#50740000000
0!
0%
b1 *
0-
02
b1 6
#50750000000
1!
1%
1-
12
#50760000000
0!
0%
b10 *
0-
02
b10 6
#50770000000
1!
1%
1-
12
#50780000000
0!
0%
b11 *
0-
02
b11 6
#50790000000
1!
1%
1-
12
15
#50800000000
0!
0%
b100 *
0-
02
b100 6
#50810000000
1!
1%
1-
12
#50820000000
0!
0%
b101 *
0-
02
b101 6
#50830000000
1!
1%
1-
12
#50840000000
0!
0%
b110 *
0-
02
b110 6
#50850000000
1!
1%
1-
12
#50860000000
0!
0%
b111 *
0-
02
b111 6
#50870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#50880000000
0!
0%
b0 *
0-
02
b0 6
#50890000000
1!
1%
1-
12
#50900000000
0!
0%
b1 *
0-
02
b1 6
#50910000000
1!
1%
1-
12
#50920000000
0!
0%
b10 *
0-
02
b10 6
#50930000000
1!
1%
1-
12
#50940000000
0!
0%
b11 *
0-
02
b11 6
#50950000000
1!
1%
1-
12
15
#50960000000
0!
0%
b100 *
0-
02
b100 6
#50970000000
1!
1%
1-
12
#50980000000
0!
0%
b101 *
0-
02
b101 6
#50990000000
1!
1%
1-
12
#51000000000
0!
0%
b110 *
0-
02
b110 6
#51010000000
1!
1%
1-
12
#51020000000
0!
0%
b111 *
0-
02
b111 6
#51030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#51040000000
0!
0%
b0 *
0-
02
b0 6
#51050000000
1!
1%
1-
12
#51060000000
0!
0%
b1 *
0-
02
b1 6
#51070000000
1!
1%
1-
12
#51080000000
0!
0%
b10 *
0-
02
b10 6
#51090000000
1!
1%
1-
12
#51100000000
0!
0%
b11 *
0-
02
b11 6
#51110000000
1!
1%
1-
12
15
#51120000000
0!
0%
b100 *
0-
02
b100 6
#51130000000
1!
1%
1-
12
#51140000000
0!
0%
b101 *
0-
02
b101 6
#51150000000
1!
1%
1-
12
#51160000000
0!
0%
b110 *
0-
02
b110 6
#51170000000
1!
1%
1-
12
#51180000000
0!
0%
b111 *
0-
02
b111 6
#51190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#51200000000
0!
0%
b0 *
0-
02
b0 6
#51210000000
1!
1%
1-
12
#51220000000
0!
0%
b1 *
0-
02
b1 6
#51230000000
1!
1%
1-
12
#51240000000
0!
0%
b10 *
0-
02
b10 6
#51250000000
1!
1%
1-
12
#51260000000
0!
0%
b11 *
0-
02
b11 6
#51270000000
1!
1%
1-
12
15
#51280000000
0!
0%
b100 *
0-
02
b100 6
#51290000000
1!
1%
1-
12
#51300000000
0!
0%
b101 *
0-
02
b101 6
#51310000000
1!
1%
1-
12
#51320000000
0!
0%
b110 *
0-
02
b110 6
#51330000000
1!
1%
1-
12
#51340000000
0!
0%
b111 *
0-
02
b111 6
#51350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#51360000000
0!
0%
b0 *
0-
02
b0 6
#51370000000
1!
1%
1-
12
#51380000000
0!
0%
b1 *
0-
02
b1 6
#51390000000
1!
1%
1-
12
#51400000000
0!
0%
b10 *
0-
02
b10 6
#51410000000
1!
1%
1-
12
#51420000000
0!
0%
b11 *
0-
02
b11 6
#51430000000
1!
1%
1-
12
15
#51440000000
0!
0%
b100 *
0-
02
b100 6
#51450000000
1!
1%
1-
12
#51460000000
0!
0%
b101 *
0-
02
b101 6
#51470000000
1!
1%
1-
12
#51480000000
0!
0%
b110 *
0-
02
b110 6
#51490000000
1!
1%
1-
12
#51500000000
0!
0%
b111 *
0-
02
b111 6
#51510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#51520000000
0!
0%
b0 *
0-
02
b0 6
#51530000000
1!
1%
1-
12
#51540000000
0!
0%
b1 *
0-
02
b1 6
#51550000000
1!
1%
1-
12
#51560000000
0!
0%
b10 *
0-
02
b10 6
#51570000000
1!
1%
1-
12
#51580000000
0!
0%
b11 *
0-
02
b11 6
#51590000000
1!
1%
1-
12
15
#51600000000
0!
0%
b100 *
0-
02
b100 6
#51610000000
1!
1%
1-
12
#51620000000
0!
0%
b101 *
0-
02
b101 6
#51630000000
1!
1%
1-
12
#51640000000
0!
0%
b110 *
0-
02
b110 6
#51650000000
1!
1%
1-
12
#51660000000
0!
0%
b111 *
0-
02
b111 6
#51670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#51680000000
0!
0%
b0 *
0-
02
b0 6
#51690000000
1!
1%
1-
12
#51700000000
0!
0%
b1 *
0-
02
b1 6
#51710000000
1!
1%
1-
12
#51720000000
0!
0%
b10 *
0-
02
b10 6
#51730000000
1!
1%
1-
12
#51740000000
0!
0%
b11 *
0-
02
b11 6
#51750000000
1!
1%
1-
12
15
#51760000000
0!
0%
b100 *
0-
02
b100 6
#51770000000
1!
1%
1-
12
#51780000000
0!
0%
b101 *
0-
02
b101 6
#51790000000
1!
1%
1-
12
#51800000000
0!
0%
b110 *
0-
02
b110 6
#51810000000
1!
1%
1-
12
#51820000000
0!
0%
b111 *
0-
02
b111 6
#51830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#51840000000
0!
0%
b0 *
0-
02
b0 6
#51850000000
1!
1%
1-
12
#51860000000
0!
0%
b1 *
0-
02
b1 6
#51870000000
1!
1%
1-
12
#51880000000
0!
0%
b10 *
0-
02
b10 6
#51890000000
1!
1%
1-
12
#51900000000
0!
0%
b11 *
0-
02
b11 6
#51910000000
1!
1%
1-
12
15
#51920000000
0!
0%
b100 *
0-
02
b100 6
#51930000000
1!
1%
1-
12
#51940000000
0!
0%
b101 *
0-
02
b101 6
#51950000000
1!
1%
1-
12
#51960000000
0!
0%
b110 *
0-
02
b110 6
#51970000000
1!
1%
1-
12
#51980000000
0!
0%
b111 *
0-
02
b111 6
#51990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#52000000000
0!
0%
b0 *
0-
02
b0 6
#52010000000
1!
1%
1-
12
#52020000000
0!
0%
b1 *
0-
02
b1 6
#52030000000
1!
1%
1-
12
#52040000000
0!
0%
b10 *
0-
02
b10 6
#52050000000
1!
1%
1-
12
#52060000000
0!
0%
b11 *
0-
02
b11 6
#52070000000
1!
1%
1-
12
15
#52080000000
0!
0%
b100 *
0-
02
b100 6
#52090000000
1!
1%
1-
12
#52100000000
0!
0%
b101 *
0-
02
b101 6
#52110000000
1!
1%
1-
12
#52120000000
0!
0%
b110 *
0-
02
b110 6
#52130000000
1!
1%
1-
12
#52140000000
0!
0%
b111 *
0-
02
b111 6
#52150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#52160000000
0!
0%
b0 *
0-
02
b0 6
#52170000000
1!
1%
1-
12
#52180000000
0!
0%
b1 *
0-
02
b1 6
#52190000000
1!
1%
1-
12
#52200000000
0!
0%
b10 *
0-
02
b10 6
#52210000000
1!
1%
1-
12
#52220000000
0!
0%
b11 *
0-
02
b11 6
#52230000000
1!
1%
1-
12
15
#52240000000
0!
0%
b100 *
0-
02
b100 6
#52250000000
1!
1%
1-
12
#52260000000
0!
0%
b101 *
0-
02
b101 6
#52270000000
1!
1%
1-
12
#52280000000
0!
0%
b110 *
0-
02
b110 6
#52290000000
1!
1%
1-
12
#52300000000
0!
0%
b111 *
0-
02
b111 6
#52310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#52320000000
0!
0%
b0 *
0-
02
b0 6
#52330000000
1!
1%
1-
12
#52340000000
0!
0%
b1 *
0-
02
b1 6
#52350000000
1!
1%
1-
12
#52360000000
0!
0%
b10 *
0-
02
b10 6
#52370000000
1!
1%
1-
12
#52380000000
0!
0%
b11 *
0-
02
b11 6
#52390000000
1!
1%
1-
12
15
#52400000000
0!
0%
b100 *
0-
02
b100 6
#52410000000
1!
1%
1-
12
#52420000000
0!
0%
b101 *
0-
02
b101 6
#52430000000
1!
1%
1-
12
#52440000000
0!
0%
b110 *
0-
02
b110 6
#52450000000
1!
1%
1-
12
#52460000000
0!
0%
b111 *
0-
02
b111 6
#52470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#52480000000
0!
0%
b0 *
0-
02
b0 6
#52490000000
1!
1%
1-
12
#52500000000
0!
0%
b1 *
0-
02
b1 6
#52510000000
1!
1%
1-
12
#52520000000
0!
0%
b10 *
0-
02
b10 6
#52530000000
1!
1%
1-
12
#52540000000
0!
0%
b11 *
0-
02
b11 6
#52550000000
1!
1%
1-
12
15
#52560000000
0!
0%
b100 *
0-
02
b100 6
#52570000000
1!
1%
1-
12
#52580000000
0!
0%
b101 *
0-
02
b101 6
#52590000000
1!
1%
1-
12
#52600000000
0!
0%
b110 *
0-
02
b110 6
#52610000000
1!
1%
1-
12
#52620000000
0!
0%
b111 *
0-
02
b111 6
#52630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#52640000000
0!
0%
b0 *
0-
02
b0 6
#52650000000
1!
1%
1-
12
#52660000000
0!
0%
b1 *
0-
02
b1 6
#52670000000
1!
1%
1-
12
#52680000000
0!
0%
b10 *
0-
02
b10 6
#52690000000
1!
1%
1-
12
#52700000000
0!
0%
b11 *
0-
02
b11 6
#52710000000
1!
1%
1-
12
15
#52720000000
0!
0%
b100 *
0-
02
b100 6
#52730000000
1!
1%
1-
12
#52740000000
0!
0%
b101 *
0-
02
b101 6
#52750000000
1!
1%
1-
12
#52760000000
0!
0%
b110 *
0-
02
b110 6
#52770000000
1!
1%
1-
12
#52780000000
0!
0%
b111 *
0-
02
b111 6
#52790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#52800000000
0!
0%
b0 *
0-
02
b0 6
#52810000000
1!
1%
1-
12
#52820000000
0!
0%
b1 *
0-
02
b1 6
#52830000000
1!
1%
1-
12
#52840000000
0!
0%
b10 *
0-
02
b10 6
#52850000000
1!
1%
1-
12
#52860000000
0!
0%
b11 *
0-
02
b11 6
#52870000000
1!
1%
1-
12
15
#52880000000
0!
0%
b100 *
0-
02
b100 6
#52890000000
1!
1%
1-
12
#52900000000
0!
0%
b101 *
0-
02
b101 6
#52910000000
1!
1%
1-
12
#52920000000
0!
0%
b110 *
0-
02
b110 6
#52930000000
1!
1%
1-
12
#52940000000
0!
0%
b111 *
0-
02
b111 6
#52950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#52960000000
0!
0%
b0 *
0-
02
b0 6
#52970000000
1!
1%
1-
12
#52980000000
0!
0%
b1 *
0-
02
b1 6
#52990000000
1!
1%
1-
12
#53000000000
0!
0%
b10 *
0-
02
b10 6
#53010000000
1!
1%
1-
12
#53020000000
0!
0%
b11 *
0-
02
b11 6
#53030000000
1!
1%
1-
12
15
#53040000000
0!
0%
b100 *
0-
02
b100 6
#53050000000
1!
1%
1-
12
#53060000000
0!
0%
b101 *
0-
02
b101 6
#53070000000
1!
1%
1-
12
#53080000000
0!
0%
b110 *
0-
02
b110 6
#53090000000
1!
1%
1-
12
#53100000000
0!
0%
b111 *
0-
02
b111 6
#53110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#53120000000
0!
0%
b0 *
0-
02
b0 6
#53130000000
1!
1%
1-
12
#53140000000
0!
0%
b1 *
0-
02
b1 6
#53150000000
1!
1%
1-
12
#53160000000
0!
0%
b10 *
0-
02
b10 6
#53170000000
1!
1%
1-
12
#53180000000
0!
0%
b11 *
0-
02
b11 6
#53190000000
1!
1%
1-
12
15
#53200000000
0!
0%
b100 *
0-
02
b100 6
#53210000000
1!
1%
1-
12
#53220000000
0!
0%
b101 *
0-
02
b101 6
#53230000000
1!
1%
1-
12
#53240000000
0!
0%
b110 *
0-
02
b110 6
#53250000000
1!
1%
1-
12
#53260000000
0!
0%
b111 *
0-
02
b111 6
#53270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#53280000000
0!
0%
b0 *
0-
02
b0 6
#53290000000
1!
1%
1-
12
#53300000000
0!
0%
b1 *
0-
02
b1 6
#53310000000
1!
1%
1-
12
#53320000000
0!
0%
b10 *
0-
02
b10 6
#53330000000
1!
1%
1-
12
#53340000000
0!
0%
b11 *
0-
02
b11 6
#53350000000
1!
1%
1-
12
15
#53360000000
0!
0%
b100 *
0-
02
b100 6
#53370000000
1!
1%
1-
12
#53380000000
0!
0%
b101 *
0-
02
b101 6
#53390000000
1!
1%
1-
12
#53400000000
0!
0%
b110 *
0-
02
b110 6
#53410000000
1!
1%
1-
12
#53420000000
0!
0%
b111 *
0-
02
b111 6
#53430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#53440000000
0!
0%
b0 *
0-
02
b0 6
#53450000000
1!
1%
1-
12
#53460000000
0!
0%
b1 *
0-
02
b1 6
#53470000000
1!
1%
1-
12
#53480000000
0!
0%
b10 *
0-
02
b10 6
#53490000000
1!
1%
1-
12
#53500000000
0!
0%
b11 *
0-
02
b11 6
#53510000000
1!
1%
1-
12
15
#53520000000
0!
0%
b100 *
0-
02
b100 6
#53530000000
1!
1%
1-
12
#53540000000
0!
0%
b101 *
0-
02
b101 6
#53550000000
1!
1%
1-
12
#53560000000
0!
0%
b110 *
0-
02
b110 6
#53570000000
1!
1%
1-
12
#53580000000
0!
0%
b111 *
0-
02
b111 6
#53590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#53600000000
0!
0%
b0 *
0-
02
b0 6
#53610000000
1!
1%
1-
12
#53620000000
0!
0%
b1 *
0-
02
b1 6
#53630000000
1!
1%
1-
12
#53640000000
0!
0%
b10 *
0-
02
b10 6
#53650000000
1!
1%
1-
12
#53660000000
0!
0%
b11 *
0-
02
b11 6
#53670000000
1!
1%
1-
12
15
#53680000000
0!
0%
b100 *
0-
02
b100 6
#53690000000
1!
1%
1-
12
#53700000000
0!
0%
b101 *
0-
02
b101 6
#53710000000
1!
1%
1-
12
#53720000000
0!
0%
b110 *
0-
02
b110 6
#53730000000
1!
1%
1-
12
#53740000000
0!
0%
b111 *
0-
02
b111 6
#53750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#53760000000
0!
0%
b0 *
0-
02
b0 6
#53770000000
1!
1%
1-
12
#53780000000
0!
0%
b1 *
0-
02
b1 6
#53790000000
1!
1%
1-
12
#53800000000
0!
0%
b10 *
0-
02
b10 6
#53810000000
1!
1%
1-
12
#53820000000
0!
0%
b11 *
0-
02
b11 6
#53830000000
1!
1%
1-
12
15
#53840000000
0!
0%
b100 *
0-
02
b100 6
#53850000000
1!
1%
1-
12
#53860000000
0!
0%
b101 *
0-
02
b101 6
#53870000000
1!
1%
1-
12
#53880000000
0!
0%
b110 *
0-
02
b110 6
#53890000000
1!
1%
1-
12
#53900000000
0!
0%
b111 *
0-
02
b111 6
#53910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#53920000000
0!
0%
b0 *
0-
02
b0 6
#53930000000
1!
1%
1-
12
#53940000000
0!
0%
b1 *
0-
02
b1 6
#53950000000
1!
1%
1-
12
#53960000000
0!
0%
b10 *
0-
02
b10 6
#53970000000
1!
1%
1-
12
#53980000000
0!
0%
b11 *
0-
02
b11 6
#53990000000
1!
1%
1-
12
15
#54000000000
0!
0%
b100 *
0-
02
b100 6
#54010000000
1!
1%
1-
12
#54020000000
0!
0%
b101 *
0-
02
b101 6
#54030000000
1!
1%
1-
12
#54040000000
0!
0%
b110 *
0-
02
b110 6
#54050000000
1!
1%
1-
12
#54060000000
0!
0%
b111 *
0-
02
b111 6
#54070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#54080000000
0!
0%
b0 *
0-
02
b0 6
#54090000000
1!
1%
1-
12
#54100000000
0!
0%
b1 *
0-
02
b1 6
#54110000000
1!
1%
1-
12
#54120000000
0!
0%
b10 *
0-
02
b10 6
#54130000000
1!
1%
1-
12
#54140000000
0!
0%
b11 *
0-
02
b11 6
#54150000000
1!
1%
1-
12
15
#54160000000
0!
0%
b100 *
0-
02
b100 6
#54170000000
1!
1%
1-
12
#54180000000
0!
0%
b101 *
0-
02
b101 6
#54190000000
1!
1%
1-
12
#54200000000
0!
0%
b110 *
0-
02
b110 6
#54210000000
1!
1%
1-
12
#54220000000
0!
0%
b111 *
0-
02
b111 6
#54230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#54240000000
0!
0%
b0 *
0-
02
b0 6
#54250000000
1!
1%
1-
12
#54260000000
0!
0%
b1 *
0-
02
b1 6
#54270000000
1!
1%
1-
12
#54280000000
0!
0%
b10 *
0-
02
b10 6
#54290000000
1!
1%
1-
12
#54300000000
0!
0%
b11 *
0-
02
b11 6
#54310000000
1!
1%
1-
12
15
#54320000000
0!
0%
b100 *
0-
02
b100 6
#54330000000
1!
1%
1-
12
#54340000000
0!
0%
b101 *
0-
02
b101 6
#54350000000
1!
1%
1-
12
#54360000000
0!
0%
b110 *
0-
02
b110 6
#54370000000
1!
1%
1-
12
#54380000000
0!
0%
b111 *
0-
02
b111 6
#54390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#54400000000
0!
0%
b0 *
0-
02
b0 6
#54410000000
1!
1%
1-
12
#54420000000
0!
0%
b1 *
0-
02
b1 6
#54430000000
1!
1%
1-
12
#54440000000
0!
0%
b10 *
0-
02
b10 6
#54450000000
1!
1%
1-
12
#54460000000
0!
0%
b11 *
0-
02
b11 6
#54470000000
1!
1%
1-
12
15
#54480000000
0!
0%
b100 *
0-
02
b100 6
#54490000000
1!
1%
1-
12
#54500000000
0!
0%
b101 *
0-
02
b101 6
#54510000000
1!
1%
1-
12
#54520000000
0!
0%
b110 *
0-
02
b110 6
#54530000000
1!
1%
1-
12
#54540000000
0!
0%
b111 *
0-
02
b111 6
#54550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#54560000000
0!
0%
b0 *
0-
02
b0 6
#54570000000
1!
1%
1-
12
#54580000000
0!
0%
b1 *
0-
02
b1 6
#54590000000
1!
1%
1-
12
#54600000000
0!
0%
b10 *
0-
02
b10 6
#54610000000
1!
1%
1-
12
#54620000000
0!
0%
b11 *
0-
02
b11 6
#54630000000
1!
1%
1-
12
15
#54640000000
0!
0%
b100 *
0-
02
b100 6
#54650000000
1!
1%
1-
12
#54660000000
0!
0%
b101 *
0-
02
b101 6
#54670000000
1!
1%
1-
12
#54680000000
0!
0%
b110 *
0-
02
b110 6
#54690000000
1!
1%
1-
12
#54700000000
0!
0%
b111 *
0-
02
b111 6
#54710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#54720000000
0!
0%
b0 *
0-
02
b0 6
#54730000000
1!
1%
1-
12
#54740000000
0!
0%
b1 *
0-
02
b1 6
#54750000000
1!
1%
1-
12
#54760000000
0!
0%
b10 *
0-
02
b10 6
#54770000000
1!
1%
1-
12
#54780000000
0!
0%
b11 *
0-
02
b11 6
#54790000000
1!
1%
1-
12
15
#54800000000
0!
0%
b100 *
0-
02
b100 6
#54810000000
1!
1%
1-
12
#54820000000
0!
0%
b101 *
0-
02
b101 6
#54830000000
1!
1%
1-
12
#54840000000
0!
0%
b110 *
0-
02
b110 6
#54850000000
1!
1%
1-
12
#54860000000
0!
0%
b111 *
0-
02
b111 6
#54870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#54880000000
0!
0%
b0 *
0-
02
b0 6
#54890000000
1!
1%
1-
12
#54900000000
0!
0%
b1 *
0-
02
b1 6
#54910000000
1!
1%
1-
12
#54920000000
0!
0%
b10 *
0-
02
b10 6
#54930000000
1!
1%
1-
12
#54940000000
0!
0%
b11 *
0-
02
b11 6
#54950000000
1!
1%
1-
12
15
#54960000000
0!
0%
b100 *
0-
02
b100 6
#54970000000
1!
1%
1-
12
#54980000000
0!
0%
b101 *
0-
02
b101 6
#54990000000
1!
1%
1-
12
#55000000000
0!
0%
b110 *
0-
02
b110 6
#55010000000
1!
1%
1-
12
#55020000000
0!
0%
b111 *
0-
02
b111 6
#55030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#55040000000
0!
0%
b0 *
0-
02
b0 6
#55050000000
1!
1%
1-
12
#55060000000
0!
0%
b1 *
0-
02
b1 6
#55070000000
1!
1%
1-
12
#55080000000
0!
0%
b10 *
0-
02
b10 6
#55090000000
1!
1%
1-
12
#55100000000
0!
0%
b11 *
0-
02
b11 6
#55110000000
1!
1%
1-
12
15
#55120000000
0!
0%
b100 *
0-
02
b100 6
#55130000000
1!
1%
1-
12
#55140000000
0!
0%
b101 *
0-
02
b101 6
#55150000000
1!
1%
1-
12
#55160000000
0!
0%
b110 *
0-
02
b110 6
#55170000000
1!
1%
1-
12
#55180000000
0!
0%
b111 *
0-
02
b111 6
#55190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#55200000000
0!
0%
b0 *
0-
02
b0 6
#55210000000
1!
1%
1-
12
#55220000000
0!
0%
b1 *
0-
02
b1 6
#55230000000
1!
1%
1-
12
#55240000000
0!
0%
b10 *
0-
02
b10 6
#55250000000
1!
1%
1-
12
#55260000000
0!
0%
b11 *
0-
02
b11 6
#55270000000
1!
1%
1-
12
15
#55280000000
0!
0%
b100 *
0-
02
b100 6
#55290000000
1!
1%
1-
12
#55300000000
0!
0%
b101 *
0-
02
b101 6
#55310000000
1!
1%
1-
12
#55320000000
0!
0%
b110 *
0-
02
b110 6
#55330000000
1!
1%
1-
12
#55340000000
0!
0%
b111 *
0-
02
b111 6
#55350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#55360000000
0!
0%
b0 *
0-
02
b0 6
#55370000000
1!
1%
1-
12
#55380000000
0!
0%
b1 *
0-
02
b1 6
#55390000000
1!
1%
1-
12
#55400000000
0!
0%
b10 *
0-
02
b10 6
#55410000000
1!
1%
1-
12
#55420000000
0!
0%
b11 *
0-
02
b11 6
#55430000000
1!
1%
1-
12
15
#55440000000
0!
0%
b100 *
0-
02
b100 6
#55450000000
1!
1%
1-
12
#55460000000
0!
0%
b101 *
0-
02
b101 6
#55470000000
1!
1%
1-
12
#55480000000
0!
0%
b110 *
0-
02
b110 6
#55490000000
1!
1%
1-
12
#55500000000
0!
0%
b111 *
0-
02
b111 6
#55510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#55520000000
0!
0%
b0 *
0-
02
b0 6
#55530000000
1!
1%
1-
12
#55540000000
0!
0%
b1 *
0-
02
b1 6
#55550000000
1!
1%
1-
12
#55560000000
0!
0%
b10 *
0-
02
b10 6
#55570000000
1!
1%
1-
12
#55580000000
0!
0%
b11 *
0-
02
b11 6
#55590000000
1!
1%
1-
12
15
#55600000000
0!
0%
b100 *
0-
02
b100 6
#55610000000
1!
1%
1-
12
#55620000000
0!
0%
b101 *
0-
02
b101 6
#55630000000
1!
1%
1-
12
#55640000000
0!
0%
b110 *
0-
02
b110 6
#55650000000
1!
1%
1-
12
#55660000000
0!
0%
b111 *
0-
02
b111 6
#55670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#55680000000
0!
0%
b0 *
0-
02
b0 6
#55690000000
1!
1%
1-
12
#55700000000
0!
0%
b1 *
0-
02
b1 6
#55710000000
1!
1%
1-
12
#55720000000
0!
0%
b10 *
0-
02
b10 6
#55730000000
1!
1%
1-
12
#55740000000
0!
0%
b11 *
0-
02
b11 6
#55750000000
1!
1%
1-
12
15
#55760000000
0!
0%
b100 *
0-
02
b100 6
#55770000000
1!
1%
1-
12
#55780000000
0!
0%
b101 *
0-
02
b101 6
#55790000000
1!
1%
1-
12
#55800000000
0!
0%
b110 *
0-
02
b110 6
#55810000000
1!
1%
1-
12
#55820000000
0!
0%
b111 *
0-
02
b111 6
#55830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#55840000000
0!
0%
b0 *
0-
02
b0 6
#55850000000
1!
1%
1-
12
#55860000000
0!
0%
b1 *
0-
02
b1 6
#55870000000
1!
1%
1-
12
#55880000000
0!
0%
b10 *
0-
02
b10 6
#55890000000
1!
1%
1-
12
#55900000000
0!
0%
b11 *
0-
02
b11 6
#55910000000
1!
1%
1-
12
15
#55920000000
0!
0%
b100 *
0-
02
b100 6
#55930000000
1!
1%
1-
12
#55940000000
0!
0%
b101 *
0-
02
b101 6
#55950000000
1!
1%
1-
12
#55960000000
0!
0%
b110 *
0-
02
b110 6
#55970000000
1!
1%
1-
12
#55980000000
0!
0%
b111 *
0-
02
b111 6
#55990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#56000000000
0!
0%
b0 *
0-
02
b0 6
#56010000000
1!
1%
1-
12
#56020000000
0!
0%
b1 *
0-
02
b1 6
#56030000000
1!
1%
1-
12
#56040000000
0!
0%
b10 *
0-
02
b10 6
#56050000000
1!
1%
1-
12
#56060000000
0!
0%
b11 *
0-
02
b11 6
#56070000000
1!
1%
1-
12
15
#56080000000
0!
0%
b100 *
0-
02
b100 6
#56090000000
1!
1%
1-
12
#56100000000
0!
0%
b101 *
0-
02
b101 6
#56110000000
1!
1%
1-
12
#56120000000
0!
0%
b110 *
0-
02
b110 6
#56130000000
1!
1%
1-
12
#56140000000
0!
0%
b111 *
0-
02
b111 6
#56150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#56160000000
0!
0%
b0 *
0-
02
b0 6
#56170000000
1!
1%
1-
12
#56180000000
0!
0%
b1 *
0-
02
b1 6
#56190000000
1!
1%
1-
12
#56200000000
0!
0%
b10 *
0-
02
b10 6
#56210000000
1!
1%
1-
12
#56220000000
0!
0%
b11 *
0-
02
b11 6
#56230000000
1!
1%
1-
12
15
#56240000000
0!
0%
b100 *
0-
02
b100 6
#56250000000
1!
1%
1-
12
#56260000000
0!
0%
b101 *
0-
02
b101 6
#56270000000
1!
1%
1-
12
#56280000000
0!
0%
b110 *
0-
02
b110 6
#56290000000
1!
1%
1-
12
#56300000000
0!
0%
b111 *
0-
02
b111 6
#56310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#56320000000
0!
0%
b0 *
0-
02
b0 6
#56330000000
1!
1%
1-
12
#56340000000
0!
0%
b1 *
0-
02
b1 6
#56350000000
1!
1%
1-
12
#56360000000
0!
0%
b10 *
0-
02
b10 6
#56370000000
1!
1%
1-
12
#56380000000
0!
0%
b11 *
0-
02
b11 6
#56390000000
1!
1%
1-
12
15
#56400000000
0!
0%
b100 *
0-
02
b100 6
#56410000000
1!
1%
1-
12
#56420000000
0!
0%
b101 *
0-
02
b101 6
#56430000000
1!
1%
1-
12
#56440000000
0!
0%
b110 *
0-
02
b110 6
#56450000000
1!
1%
1-
12
#56460000000
0!
0%
b111 *
0-
02
b111 6
#56470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#56480000000
0!
0%
b0 *
0-
02
b0 6
#56490000000
1!
1%
1-
12
#56500000000
0!
0%
b1 *
0-
02
b1 6
#56510000000
1!
1%
1-
12
#56520000000
0!
0%
b10 *
0-
02
b10 6
#56530000000
1!
1%
1-
12
#56540000000
0!
0%
b11 *
0-
02
b11 6
#56550000000
1!
1%
1-
12
15
#56560000000
0!
0%
b100 *
0-
02
b100 6
#56570000000
1!
1%
1-
12
#56580000000
0!
0%
b101 *
0-
02
b101 6
#56590000000
1!
1%
1-
12
#56600000000
0!
0%
b110 *
0-
02
b110 6
#56610000000
1!
1%
1-
12
#56620000000
0!
0%
b111 *
0-
02
b111 6
#56630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#56640000000
0!
0%
b0 *
0-
02
b0 6
#56650000000
1!
1%
1-
12
#56660000000
0!
0%
b1 *
0-
02
b1 6
#56670000000
1!
1%
1-
12
#56680000000
0!
0%
b10 *
0-
02
b10 6
#56690000000
1!
1%
1-
12
#56700000000
0!
0%
b11 *
0-
02
b11 6
#56710000000
1!
1%
1-
12
15
#56720000000
0!
0%
b100 *
0-
02
b100 6
#56730000000
1!
1%
1-
12
#56740000000
0!
0%
b101 *
0-
02
b101 6
#56750000000
1!
1%
1-
12
#56760000000
0!
0%
b110 *
0-
02
b110 6
#56770000000
1!
1%
1-
12
#56780000000
0!
0%
b111 *
0-
02
b111 6
#56790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#56800000000
0!
0%
b0 *
0-
02
b0 6
#56810000000
1!
1%
1-
12
#56820000000
0!
0%
b1 *
0-
02
b1 6
#56830000000
1!
1%
1-
12
#56840000000
0!
0%
b10 *
0-
02
b10 6
#56850000000
1!
1%
1-
12
#56860000000
0!
0%
b11 *
0-
02
b11 6
#56870000000
1!
1%
1-
12
15
#56880000000
0!
0%
b100 *
0-
02
b100 6
#56890000000
1!
1%
1-
12
#56900000000
0!
0%
b101 *
0-
02
b101 6
#56910000000
1!
1%
1-
12
#56920000000
0!
0%
b110 *
0-
02
b110 6
#56930000000
1!
1%
1-
12
#56940000000
0!
0%
b111 *
0-
02
b111 6
#56950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#56960000000
0!
0%
b0 *
0-
02
b0 6
#56970000000
1!
1%
1-
12
#56980000000
0!
0%
b1 *
0-
02
b1 6
#56990000000
1!
1%
1-
12
#57000000000
0!
0%
b10 *
0-
02
b10 6
#57010000000
1!
1%
1-
12
#57020000000
0!
0%
b11 *
0-
02
b11 6
#57030000000
1!
1%
1-
12
15
#57040000000
0!
0%
b100 *
0-
02
b100 6
#57050000000
1!
1%
1-
12
#57060000000
0!
0%
b101 *
0-
02
b101 6
#57070000000
1!
1%
1-
12
#57080000000
0!
0%
b110 *
0-
02
b110 6
#57090000000
1!
1%
1-
12
#57100000000
0!
0%
b111 *
0-
02
b111 6
#57110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#57120000000
0!
0%
b0 *
0-
02
b0 6
#57130000000
1!
1%
1-
12
#57140000000
0!
0%
b1 *
0-
02
b1 6
#57150000000
1!
1%
1-
12
#57160000000
0!
0%
b10 *
0-
02
b10 6
#57170000000
1!
1%
1-
12
#57180000000
0!
0%
b11 *
0-
02
b11 6
#57190000000
1!
1%
1-
12
15
#57200000000
0!
0%
b100 *
0-
02
b100 6
#57210000000
1!
1%
1-
12
#57220000000
0!
0%
b101 *
0-
02
b101 6
#57230000000
1!
1%
1-
12
#57240000000
0!
0%
b110 *
0-
02
b110 6
#57250000000
1!
1%
1-
12
#57260000000
0!
0%
b111 *
0-
02
b111 6
#57270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#57280000000
0!
0%
b0 *
0-
02
b0 6
#57290000000
1!
1%
1-
12
#57300000000
0!
0%
b1 *
0-
02
b1 6
#57310000000
1!
1%
1-
12
#57320000000
0!
0%
b10 *
0-
02
b10 6
#57330000000
1!
1%
1-
12
#57340000000
0!
0%
b11 *
0-
02
b11 6
#57350000000
1!
1%
1-
12
15
#57360000000
0!
0%
b100 *
0-
02
b100 6
#57370000000
1!
1%
1-
12
#57380000000
0!
0%
b101 *
0-
02
b101 6
#57390000000
1!
1%
1-
12
#57400000000
0!
0%
b110 *
0-
02
b110 6
#57410000000
1!
1%
1-
12
#57420000000
0!
0%
b111 *
0-
02
b111 6
#57430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#57440000000
0!
0%
b0 *
0-
02
b0 6
#57450000000
1!
1%
1-
12
#57460000000
0!
0%
b1 *
0-
02
b1 6
#57470000000
1!
1%
1-
12
#57480000000
0!
0%
b10 *
0-
02
b10 6
#57490000000
1!
1%
1-
12
#57500000000
0!
0%
b11 *
0-
02
b11 6
#57510000000
1!
1%
1-
12
15
#57520000000
0!
0%
b100 *
0-
02
b100 6
#57530000000
1!
1%
1-
12
#57540000000
0!
0%
b101 *
0-
02
b101 6
#57550000000
1!
1%
1-
12
#57560000000
0!
0%
b110 *
0-
02
b110 6
#57570000000
1!
1%
1-
12
#57580000000
0!
0%
b111 *
0-
02
b111 6
#57590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#57600000000
0!
0%
b0 *
0-
02
b0 6
#57610000000
1!
1%
1-
12
#57620000000
0!
0%
b1 *
0-
02
b1 6
#57630000000
1!
1%
1-
12
#57640000000
0!
0%
b10 *
0-
02
b10 6
#57650000000
1!
1%
1-
12
#57660000000
0!
0%
b11 *
0-
02
b11 6
#57670000000
1!
1%
1-
12
15
#57680000000
0!
0%
b100 *
0-
02
b100 6
#57690000000
1!
1%
1-
12
#57700000000
0!
0%
b101 *
0-
02
b101 6
#57710000000
1!
1%
1-
12
#57720000000
0!
0%
b110 *
0-
02
b110 6
#57730000000
1!
1%
1-
12
#57740000000
0!
0%
b111 *
0-
02
b111 6
#57750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#57760000000
0!
0%
b0 *
0-
02
b0 6
#57770000000
1!
1%
1-
12
#57780000000
0!
0%
b1 *
0-
02
b1 6
#57790000000
1!
1%
1-
12
#57800000000
0!
0%
b10 *
0-
02
b10 6
#57810000000
1!
1%
1-
12
#57820000000
0!
0%
b11 *
0-
02
b11 6
#57830000000
1!
1%
1-
12
15
#57840000000
0!
0%
b100 *
0-
02
b100 6
#57850000000
1!
1%
1-
12
#57860000000
0!
0%
b101 *
0-
02
b101 6
#57870000000
1!
1%
1-
12
#57880000000
0!
0%
b110 *
0-
02
b110 6
#57890000000
1!
1%
1-
12
#57900000000
0!
0%
b111 *
0-
02
b111 6
#57910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#57920000000
0!
0%
b0 *
0-
02
b0 6
#57930000000
1!
1%
1-
12
#57940000000
0!
0%
b1 *
0-
02
b1 6
#57950000000
1!
1%
1-
12
#57960000000
0!
0%
b10 *
0-
02
b10 6
#57970000000
1!
1%
1-
12
#57980000000
0!
0%
b11 *
0-
02
b11 6
#57990000000
1!
1%
1-
12
15
#58000000000
0!
0%
b100 *
0-
02
b100 6
#58010000000
1!
1%
1-
12
#58020000000
0!
0%
b101 *
0-
02
b101 6
#58030000000
1!
1%
1-
12
#58040000000
0!
0%
b110 *
0-
02
b110 6
#58050000000
1!
1%
1-
12
#58060000000
0!
0%
b111 *
0-
02
b111 6
#58070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#58080000000
0!
0%
b0 *
0-
02
b0 6
#58090000000
1!
1%
1-
12
#58100000000
0!
0%
b1 *
0-
02
b1 6
#58110000000
1!
1%
1-
12
#58120000000
0!
0%
b10 *
0-
02
b10 6
#58130000000
1!
1%
1-
12
#58140000000
0!
0%
b11 *
0-
02
b11 6
#58150000000
1!
1%
1-
12
15
#58160000000
0!
0%
b100 *
0-
02
b100 6
#58170000000
1!
1%
1-
12
#58180000000
0!
0%
b101 *
0-
02
b101 6
#58190000000
1!
1%
1-
12
#58200000000
0!
0%
b110 *
0-
02
b110 6
#58210000000
1!
1%
1-
12
#58220000000
0!
0%
b111 *
0-
02
b111 6
#58230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#58240000000
0!
0%
b0 *
0-
02
b0 6
#58250000000
1!
1%
1-
12
#58260000000
0!
0%
b1 *
0-
02
b1 6
#58270000000
1!
1%
1-
12
#58280000000
0!
0%
b10 *
0-
02
b10 6
#58290000000
1!
1%
1-
12
#58300000000
0!
0%
b11 *
0-
02
b11 6
#58310000000
1!
1%
1-
12
15
#58320000000
0!
0%
b100 *
0-
02
b100 6
#58330000000
1!
1%
1-
12
#58340000000
0!
0%
b101 *
0-
02
b101 6
#58350000000
1!
1%
1-
12
#58360000000
0!
0%
b110 *
0-
02
b110 6
#58370000000
1!
1%
1-
12
#58380000000
0!
0%
b111 *
0-
02
b111 6
#58390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#58400000000
0!
0%
b0 *
0-
02
b0 6
#58410000000
1!
1%
1-
12
#58420000000
0!
0%
b1 *
0-
02
b1 6
#58430000000
1!
1%
1-
12
#58440000000
0!
0%
b10 *
0-
02
b10 6
#58450000000
1!
1%
1-
12
#58460000000
0!
0%
b11 *
0-
02
b11 6
#58470000000
1!
1%
1-
12
15
#58480000000
0!
0%
b100 *
0-
02
b100 6
#58490000000
1!
1%
1-
12
#58500000000
0!
0%
b101 *
0-
02
b101 6
#58510000000
1!
1%
1-
12
#58520000000
0!
0%
b110 *
0-
02
b110 6
#58530000000
1!
1%
1-
12
#58540000000
0!
0%
b111 *
0-
02
b111 6
#58550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#58560000000
0!
0%
b0 *
0-
02
b0 6
#58570000000
1!
1%
1-
12
#58580000000
0!
0%
b1 *
0-
02
b1 6
#58590000000
1!
1%
1-
12
#58600000000
0!
0%
b10 *
0-
02
b10 6
#58610000000
1!
1%
1-
12
#58620000000
0!
0%
b11 *
0-
02
b11 6
#58630000000
1!
1%
1-
12
15
#58640000000
0!
0%
b100 *
0-
02
b100 6
#58650000000
1!
1%
1-
12
#58660000000
0!
0%
b101 *
0-
02
b101 6
#58670000000
1!
1%
1-
12
#58680000000
0!
0%
b110 *
0-
02
b110 6
#58690000000
1!
1%
1-
12
#58700000000
0!
0%
b111 *
0-
02
b111 6
#58710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#58720000000
0!
0%
b0 *
0-
02
b0 6
#58730000000
1!
1%
1-
12
#58740000000
0!
0%
b1 *
0-
02
b1 6
#58750000000
1!
1%
1-
12
#58760000000
0!
0%
b10 *
0-
02
b10 6
#58770000000
1!
1%
1-
12
#58780000000
0!
0%
b11 *
0-
02
b11 6
#58790000000
1!
1%
1-
12
15
#58800000000
0!
0%
b100 *
0-
02
b100 6
#58810000000
1!
1%
1-
12
#58820000000
0!
0%
b101 *
0-
02
b101 6
#58830000000
1!
1%
1-
12
#58840000000
0!
0%
b110 *
0-
02
b110 6
#58850000000
1!
1%
1-
12
#58860000000
0!
0%
b111 *
0-
02
b111 6
#58870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#58880000000
0!
0%
b0 *
0-
02
b0 6
#58890000000
1!
1%
1-
12
#58900000000
0!
0%
b1 *
0-
02
b1 6
#58910000000
1!
1%
1-
12
#58920000000
0!
0%
b10 *
0-
02
b10 6
#58930000000
1!
1%
1-
12
#58940000000
0!
0%
b11 *
0-
02
b11 6
#58950000000
1!
1%
1-
12
15
#58960000000
0!
0%
b100 *
0-
02
b100 6
#58970000000
1!
1%
1-
12
#58980000000
0!
0%
b101 *
0-
02
b101 6
#58990000000
1!
1%
1-
12
#59000000000
0!
0%
b110 *
0-
02
b110 6
#59010000000
1!
1%
1-
12
#59020000000
0!
0%
b111 *
0-
02
b111 6
#59030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#59040000000
0!
0%
b0 *
0-
02
b0 6
#59050000000
1!
1%
1-
12
#59060000000
0!
0%
b1 *
0-
02
b1 6
#59070000000
1!
1%
1-
12
#59080000000
0!
0%
b10 *
0-
02
b10 6
#59090000000
1!
1%
1-
12
#59100000000
0!
0%
b11 *
0-
02
b11 6
#59110000000
1!
1%
1-
12
15
#59120000000
0!
0%
b100 *
0-
02
b100 6
#59130000000
1!
1%
1-
12
#59140000000
0!
0%
b101 *
0-
02
b101 6
#59150000000
1!
1%
1-
12
#59160000000
0!
0%
b110 *
0-
02
b110 6
#59170000000
1!
1%
1-
12
#59180000000
0!
0%
b111 *
0-
02
b111 6
#59190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#59200000000
0!
0%
b0 *
0-
02
b0 6
#59210000000
1!
1%
1-
12
#59220000000
0!
0%
b1 *
0-
02
b1 6
#59230000000
1!
1%
1-
12
#59240000000
0!
0%
b10 *
0-
02
b10 6
#59250000000
1!
1%
1-
12
#59260000000
0!
0%
b11 *
0-
02
b11 6
#59270000000
1!
1%
1-
12
15
#59280000000
0!
0%
b100 *
0-
02
b100 6
#59290000000
1!
1%
1-
12
#59300000000
0!
0%
b101 *
0-
02
b101 6
#59310000000
1!
1%
1-
12
#59320000000
0!
0%
b110 *
0-
02
b110 6
#59330000000
1!
1%
1-
12
#59340000000
0!
0%
b111 *
0-
02
b111 6
#59350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#59360000000
0!
0%
b0 *
0-
02
b0 6
#59370000000
1!
1%
1-
12
#59380000000
0!
0%
b1 *
0-
02
b1 6
#59390000000
1!
1%
1-
12
#59400000000
0!
0%
b10 *
0-
02
b10 6
#59410000000
1!
1%
1-
12
#59420000000
0!
0%
b11 *
0-
02
b11 6
#59430000000
1!
1%
1-
12
15
#59440000000
0!
0%
b100 *
0-
02
b100 6
#59450000000
1!
1%
1-
12
#59460000000
0!
0%
b101 *
0-
02
b101 6
#59470000000
1!
1%
1-
12
#59480000000
0!
0%
b110 *
0-
02
b110 6
#59490000000
1!
1%
1-
12
#59500000000
0!
0%
b111 *
0-
02
b111 6
#59510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#59520000000
0!
0%
b0 *
0-
02
b0 6
#59530000000
1!
1%
1-
12
#59540000000
0!
0%
b1 *
0-
02
b1 6
#59550000000
1!
1%
1-
12
#59560000000
0!
0%
b10 *
0-
02
b10 6
#59570000000
1!
1%
1-
12
#59580000000
0!
0%
b11 *
0-
02
b11 6
#59590000000
1!
1%
1-
12
15
#59600000000
0!
0%
b100 *
0-
02
b100 6
#59610000000
1!
1%
1-
12
#59620000000
0!
0%
b101 *
0-
02
b101 6
#59630000000
1!
1%
1-
12
#59640000000
0!
0%
b110 *
0-
02
b110 6
#59650000000
1!
1%
1-
12
#59660000000
0!
0%
b111 *
0-
02
b111 6
#59670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#59680000000
0!
0%
b0 *
0-
02
b0 6
#59690000000
1!
1%
1-
12
#59700000000
0!
0%
b1 *
0-
02
b1 6
#59710000000
1!
1%
1-
12
#59720000000
0!
0%
b10 *
0-
02
b10 6
#59730000000
1!
1%
1-
12
#59740000000
0!
0%
b11 *
0-
02
b11 6
#59750000000
1!
1%
1-
12
15
#59760000000
0!
0%
b100 *
0-
02
b100 6
#59770000000
1!
1%
1-
12
#59780000000
0!
0%
b101 *
0-
02
b101 6
#59790000000
1!
1%
1-
12
#59800000000
0!
0%
b110 *
0-
02
b110 6
#59810000000
1!
1%
1-
12
#59820000000
0!
0%
b111 *
0-
02
b111 6
#59830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#59840000000
0!
0%
b0 *
0-
02
b0 6
#59850000000
1!
1%
1-
12
#59860000000
0!
0%
b1 *
0-
02
b1 6
#59870000000
1!
1%
1-
12
#59880000000
0!
0%
b10 *
0-
02
b10 6
#59890000000
1!
1%
1-
12
#59900000000
0!
0%
b11 *
0-
02
b11 6
#59910000000
1!
1%
1-
12
15
#59920000000
0!
0%
b100 *
0-
02
b100 6
#59930000000
1!
1%
1-
12
#59940000000
0!
0%
b101 *
0-
02
b101 6
#59950000000
1!
1%
1-
12
#59960000000
0!
0%
b110 *
0-
02
b110 6
#59970000000
1!
1%
1-
12
#59980000000
0!
0%
b111 *
0-
02
b111 6
#59990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#60000000000
0!
0%
b0 *
0-
02
b0 6
#60010000000
1!
1%
1-
12
#60020000000
0!
0%
b1 *
0-
02
b1 6
#60030000000
1!
1%
1-
12
#60040000000
0!
0%
b10 *
0-
02
b10 6
#60050000000
1!
1%
1-
12
#60060000000
0!
0%
b11 *
0-
02
b11 6
#60070000000
1!
1%
1-
12
15
#60080000000
0!
0%
b100 *
0-
02
b100 6
#60090000000
1!
1%
1-
12
#60100000000
0!
0%
b101 *
0-
02
b101 6
#60110000000
1!
1%
1-
12
#60120000000
0!
0%
b110 *
0-
02
b110 6
#60130000000
1!
1%
1-
12
#60140000000
0!
0%
b111 *
0-
02
b111 6
#60150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#60160000000
0!
0%
b0 *
0-
02
b0 6
#60170000000
1!
1%
1-
12
#60180000000
0!
0%
b1 *
0-
02
b1 6
#60190000000
1!
1%
1-
12
#60200000000
0!
0%
b10 *
0-
02
b10 6
#60210000000
1!
1%
1-
12
#60220000000
0!
0%
b11 *
0-
02
b11 6
#60230000000
1!
1%
1-
12
15
#60240000000
0!
0%
b100 *
0-
02
b100 6
#60250000000
1!
1%
1-
12
#60260000000
0!
0%
b101 *
0-
02
b101 6
#60270000000
1!
1%
1-
12
#60280000000
0!
0%
b110 *
0-
02
b110 6
#60290000000
1!
1%
1-
12
#60300000000
0!
0%
b111 *
0-
02
b111 6
#60310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#60320000000
0!
0%
b0 *
0-
02
b0 6
#60330000000
1!
1%
1-
12
#60340000000
0!
0%
b1 *
0-
02
b1 6
#60350000000
1!
1%
1-
12
#60360000000
0!
0%
b10 *
0-
02
b10 6
#60370000000
1!
1%
1-
12
#60380000000
0!
0%
b11 *
0-
02
b11 6
#60390000000
1!
1%
1-
12
15
#60400000000
0!
0%
b100 *
0-
02
b100 6
#60410000000
1!
1%
1-
12
#60420000000
0!
0%
b101 *
0-
02
b101 6
#60430000000
1!
1%
1-
12
#60440000000
0!
0%
b110 *
0-
02
b110 6
#60450000000
1!
1%
1-
12
#60460000000
0!
0%
b111 *
0-
02
b111 6
#60470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#60480000000
0!
0%
b0 *
0-
02
b0 6
#60490000000
1!
1%
1-
12
#60500000000
0!
0%
b1 *
0-
02
b1 6
#60510000000
1!
1%
1-
12
#60520000000
0!
0%
b10 *
0-
02
b10 6
#60530000000
1!
1%
1-
12
#60540000000
0!
0%
b11 *
0-
02
b11 6
#60550000000
1!
1%
1-
12
15
#60560000000
0!
0%
b100 *
0-
02
b100 6
#60570000000
1!
1%
1-
12
#60580000000
0!
0%
b101 *
0-
02
b101 6
#60590000000
1!
1%
1-
12
#60600000000
0!
0%
b110 *
0-
02
b110 6
#60610000000
1!
1%
1-
12
#60620000000
0!
0%
b111 *
0-
02
b111 6
#60630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#60640000000
0!
0%
b0 *
0-
02
b0 6
#60650000000
1!
1%
1-
12
#60660000000
0!
0%
b1 *
0-
02
b1 6
#60670000000
1!
1%
1-
12
#60680000000
0!
0%
b10 *
0-
02
b10 6
#60690000000
1!
1%
1-
12
#60700000000
0!
0%
b11 *
0-
02
b11 6
#60710000000
1!
1%
1-
12
15
#60720000000
0!
0%
b100 *
0-
02
b100 6
#60730000000
1!
1%
1-
12
#60740000000
0!
0%
b101 *
0-
02
b101 6
#60750000000
1!
1%
1-
12
#60760000000
0!
0%
b110 *
0-
02
b110 6
#60770000000
1!
1%
1-
12
#60780000000
0!
0%
b111 *
0-
02
b111 6
#60790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#60800000000
0!
0%
b0 *
0-
02
b0 6
#60810000000
1!
1%
1-
12
#60820000000
0!
0%
b1 *
0-
02
b1 6
#60830000000
1!
1%
1-
12
#60840000000
0!
0%
b10 *
0-
02
b10 6
#60850000000
1!
1%
1-
12
#60860000000
0!
0%
b11 *
0-
02
b11 6
#60870000000
1!
1%
1-
12
15
#60880000000
0!
0%
b100 *
0-
02
b100 6
#60890000000
1!
1%
1-
12
#60900000000
0!
0%
b101 *
0-
02
b101 6
#60910000000
1!
1%
1-
12
#60920000000
0!
0%
b110 *
0-
02
b110 6
#60930000000
1!
1%
1-
12
#60940000000
0!
0%
b111 *
0-
02
b111 6
#60950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#60960000000
0!
0%
b0 *
0-
02
b0 6
#60970000000
1!
1%
1-
12
#60980000000
0!
0%
b1 *
0-
02
b1 6
#60990000000
1!
1%
1-
12
#61000000000
0!
0%
b10 *
0-
02
b10 6
#61010000000
1!
1%
1-
12
#61020000000
0!
0%
b11 *
0-
02
b11 6
#61030000000
1!
1%
1-
12
15
#61040000000
0!
0%
b100 *
0-
02
b100 6
#61050000000
1!
1%
1-
12
#61060000000
0!
0%
b101 *
0-
02
b101 6
#61070000000
1!
1%
1-
12
#61080000000
0!
0%
b110 *
0-
02
b110 6
#61090000000
1!
1%
1-
12
#61100000000
0!
0%
b111 *
0-
02
b111 6
#61110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#61120000000
0!
0%
b0 *
0-
02
b0 6
#61130000000
1!
1%
1-
12
#61140000000
0!
0%
b1 *
0-
02
b1 6
#61150000000
1!
1%
1-
12
#61160000000
0!
0%
b10 *
0-
02
b10 6
#61170000000
1!
1%
1-
12
#61180000000
0!
0%
b11 *
0-
02
b11 6
#61190000000
1!
1%
1-
12
15
#61200000000
0!
0%
b100 *
0-
02
b100 6
#61210000000
1!
1%
1-
12
#61220000000
0!
0%
b101 *
0-
02
b101 6
#61230000000
1!
1%
1-
12
#61240000000
0!
0%
b110 *
0-
02
b110 6
#61250000000
1!
1%
1-
12
#61260000000
0!
0%
b111 *
0-
02
b111 6
#61270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#61280000000
0!
0%
b0 *
0-
02
b0 6
#61290000000
1!
1%
1-
12
#61300000000
0!
0%
b1 *
0-
02
b1 6
#61310000000
1!
1%
1-
12
#61320000000
0!
0%
b10 *
0-
02
b10 6
#61330000000
1!
1%
1-
12
#61340000000
0!
0%
b11 *
0-
02
b11 6
#61350000000
1!
1%
1-
12
15
#61360000000
0!
0%
b100 *
0-
02
b100 6
#61370000000
1!
1%
1-
12
#61380000000
0!
0%
b101 *
0-
02
b101 6
#61390000000
1!
1%
1-
12
#61400000000
0!
0%
b110 *
0-
02
b110 6
#61410000000
1!
1%
1-
12
#61420000000
0!
0%
b111 *
0-
02
b111 6
#61430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#61440000000
0!
0%
b0 *
0-
02
b0 6
#61450000000
1!
1%
1-
12
#61460000000
0!
0%
b1 *
0-
02
b1 6
#61470000000
1!
1%
1-
12
#61480000000
0!
0%
b10 *
0-
02
b10 6
#61490000000
1!
1%
1-
12
#61500000000
0!
0%
b11 *
0-
02
b11 6
#61510000000
1!
1%
1-
12
15
#61520000000
0!
0%
b100 *
0-
02
b100 6
#61530000000
1!
1%
1-
12
#61540000000
0!
0%
b101 *
0-
02
b101 6
#61550000000
1!
1%
1-
12
#61560000000
0!
0%
b110 *
0-
02
b110 6
#61570000000
1!
1%
1-
12
#61580000000
0!
0%
b111 *
0-
02
b111 6
#61590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#61600000000
0!
0%
b0 *
0-
02
b0 6
#61610000000
1!
1%
1-
12
#61620000000
0!
0%
b1 *
0-
02
b1 6
#61630000000
1!
1%
1-
12
#61640000000
0!
0%
b10 *
0-
02
b10 6
#61650000000
1!
1%
1-
12
#61660000000
0!
0%
b11 *
0-
02
b11 6
#61670000000
1!
1%
1-
12
15
#61680000000
0!
0%
b100 *
0-
02
b100 6
#61690000000
1!
1%
1-
12
#61700000000
0!
0%
b101 *
0-
02
b101 6
#61710000000
1!
1%
1-
12
#61720000000
0!
0%
b110 *
0-
02
b110 6
#61730000000
1!
1%
1-
12
#61740000000
0!
0%
b111 *
0-
02
b111 6
#61750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#61760000000
0!
0%
b0 *
0-
02
b0 6
#61770000000
1!
1%
1-
12
#61780000000
0!
0%
b1 *
0-
02
b1 6
#61790000000
1!
1%
1-
12
#61800000000
0!
0%
b10 *
0-
02
b10 6
#61810000000
1!
1%
1-
12
#61820000000
0!
0%
b11 *
0-
02
b11 6
#61830000000
1!
1%
1-
12
15
#61840000000
0!
0%
b100 *
0-
02
b100 6
#61850000000
1!
1%
1-
12
#61860000000
0!
0%
b101 *
0-
02
b101 6
#61870000000
1!
1%
1-
12
#61880000000
0!
0%
b110 *
0-
02
b110 6
#61890000000
1!
1%
1-
12
#61900000000
0!
0%
b111 *
0-
02
b111 6
#61910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#61920000000
0!
0%
b0 *
0-
02
b0 6
#61930000000
1!
1%
1-
12
#61940000000
0!
0%
b1 *
0-
02
b1 6
#61950000000
1!
1%
1-
12
#61960000000
0!
0%
b10 *
0-
02
b10 6
#61970000000
1!
1%
1-
12
#61980000000
0!
0%
b11 *
0-
02
b11 6
#61990000000
1!
1%
1-
12
15
#62000000000
0!
0%
b100 *
0-
02
b100 6
#62010000000
1!
1%
1-
12
#62020000000
0!
0%
b101 *
0-
02
b101 6
#62030000000
1!
1%
1-
12
#62040000000
0!
0%
b110 *
0-
02
b110 6
#62050000000
1!
1%
1-
12
#62060000000
0!
0%
b111 *
0-
02
b111 6
#62070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#62080000000
0!
0%
b0 *
0-
02
b0 6
#62090000000
1!
1%
1-
12
#62100000000
0!
0%
b1 *
0-
02
b1 6
#62110000000
1!
1%
1-
12
#62120000000
0!
0%
b10 *
0-
02
b10 6
#62130000000
1!
1%
1-
12
#62140000000
0!
0%
b11 *
0-
02
b11 6
#62150000000
1!
1%
1-
12
15
#62160000000
0!
0%
b100 *
0-
02
b100 6
#62170000000
1!
1%
1-
12
#62180000000
0!
0%
b101 *
0-
02
b101 6
#62190000000
1!
1%
1-
12
#62200000000
0!
0%
b110 *
0-
02
b110 6
#62210000000
1!
1%
1-
12
#62220000000
0!
0%
b111 *
0-
02
b111 6
#62230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#62240000000
0!
0%
b0 *
0-
02
b0 6
#62250000000
1!
1%
1-
12
#62260000000
0!
0%
b1 *
0-
02
b1 6
#62270000000
1!
1%
1-
12
#62280000000
0!
0%
b10 *
0-
02
b10 6
#62290000000
1!
1%
1-
12
#62300000000
0!
0%
b11 *
0-
02
b11 6
#62310000000
1!
1%
1-
12
15
#62320000000
0!
0%
b100 *
0-
02
b100 6
#62330000000
1!
1%
1-
12
#62340000000
0!
0%
b101 *
0-
02
b101 6
#62350000000
1!
1%
1-
12
#62360000000
0!
0%
b110 *
0-
02
b110 6
#62370000000
1!
1%
1-
12
#62380000000
0!
0%
b111 *
0-
02
b111 6
#62390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#62400000000
0!
0%
b0 *
0-
02
b0 6
#62410000000
1!
1%
1-
12
#62420000000
0!
0%
b1 *
0-
02
b1 6
#62430000000
1!
1%
1-
12
#62440000000
0!
0%
b10 *
0-
02
b10 6
#62450000000
1!
1%
1-
12
#62460000000
0!
0%
b11 *
0-
02
b11 6
#62470000000
1!
1%
1-
12
15
#62480000000
0!
0%
b100 *
0-
02
b100 6
#62490000000
1!
1%
1-
12
#62500000000
0!
0%
b101 *
0-
02
b101 6
#62510000000
1!
1%
1-
12
#62520000000
0!
0%
b110 *
0-
02
b110 6
#62530000000
1!
1%
1-
12
#62540000000
0!
0%
b111 *
0-
02
b111 6
#62550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#62560000000
0!
0%
b0 *
0-
02
b0 6
#62570000000
1!
1%
1-
12
#62580000000
0!
0%
b1 *
0-
02
b1 6
#62590000000
1!
1%
1-
12
#62600000000
0!
0%
b10 *
0-
02
b10 6
#62610000000
1!
1%
1-
12
#62620000000
0!
0%
b11 *
0-
02
b11 6
#62630000000
1!
1%
1-
12
15
#62640000000
0!
0%
b100 *
0-
02
b100 6
#62650000000
1!
1%
1-
12
#62660000000
0!
0%
b101 *
0-
02
b101 6
#62670000000
1!
1%
1-
12
#62680000000
0!
0%
b110 *
0-
02
b110 6
#62690000000
1!
1%
1-
12
#62700000000
0!
0%
b111 *
0-
02
b111 6
#62710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#62720000000
0!
0%
b0 *
0-
02
b0 6
#62730000000
1!
1%
1-
12
#62740000000
0!
0%
b1 *
0-
02
b1 6
#62750000000
1!
1%
1-
12
#62760000000
0!
0%
b10 *
0-
02
b10 6
#62770000000
1!
1%
1-
12
#62780000000
0!
0%
b11 *
0-
02
b11 6
#62790000000
1!
1%
1-
12
15
#62800000000
0!
0%
b100 *
0-
02
b100 6
#62810000000
1!
1%
1-
12
#62820000000
0!
0%
b101 *
0-
02
b101 6
#62830000000
1!
1%
1-
12
#62840000000
0!
0%
b110 *
0-
02
b110 6
#62850000000
1!
1%
1-
12
#62860000000
0!
0%
b111 *
0-
02
b111 6
#62870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#62880000000
0!
0%
b0 *
0-
02
b0 6
#62890000000
1!
1%
1-
12
#62900000000
0!
0%
b1 *
0-
02
b1 6
#62910000000
1!
1%
1-
12
#62920000000
0!
0%
b10 *
0-
02
b10 6
#62930000000
1!
1%
1-
12
#62940000000
0!
0%
b11 *
0-
02
b11 6
#62950000000
1!
1%
1-
12
15
#62960000000
0!
0%
b100 *
0-
02
b100 6
#62970000000
1!
1%
1-
12
#62980000000
0!
0%
b101 *
0-
02
b101 6
#62990000000
1!
1%
1-
12
#63000000000
0!
0%
b110 *
0-
02
b110 6
#63010000000
1!
1%
1-
12
#63020000000
0!
0%
b111 *
0-
02
b111 6
#63030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#63040000000
0!
0%
b0 *
0-
02
b0 6
#63050000000
1!
1%
1-
12
#63060000000
0!
0%
b1 *
0-
02
b1 6
#63070000000
1!
1%
1-
12
#63080000000
0!
0%
b10 *
0-
02
b10 6
#63090000000
1!
1%
1-
12
#63100000000
0!
0%
b11 *
0-
02
b11 6
#63110000000
1!
1%
1-
12
15
#63120000000
0!
0%
b100 *
0-
02
b100 6
#63130000000
1!
1%
1-
12
#63140000000
0!
0%
b101 *
0-
02
b101 6
#63150000000
1!
1%
1-
12
#63160000000
0!
0%
b110 *
0-
02
b110 6
#63170000000
1!
1%
1-
12
#63180000000
0!
0%
b111 *
0-
02
b111 6
#63190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#63200000000
0!
0%
b0 *
0-
02
b0 6
#63210000000
1!
1%
1-
12
#63220000000
0!
0%
b1 *
0-
02
b1 6
#63230000000
1!
1%
1-
12
#63240000000
0!
0%
b10 *
0-
02
b10 6
#63250000000
1!
1%
1-
12
#63260000000
0!
0%
b11 *
0-
02
b11 6
#63270000000
1!
1%
1-
12
15
#63280000000
0!
0%
b100 *
0-
02
b100 6
#63290000000
1!
1%
1-
12
#63300000000
0!
0%
b101 *
0-
02
b101 6
#63310000000
1!
1%
1-
12
#63320000000
0!
0%
b110 *
0-
02
b110 6
#63330000000
1!
1%
1-
12
#63340000000
0!
0%
b111 *
0-
02
b111 6
#63350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#63360000000
0!
0%
b0 *
0-
02
b0 6
#63370000000
1!
1%
1-
12
#63380000000
0!
0%
b1 *
0-
02
b1 6
#63390000000
1!
1%
1-
12
#63400000000
0!
0%
b10 *
0-
02
b10 6
#63410000000
1!
1%
1-
12
#63420000000
0!
0%
b11 *
0-
02
b11 6
#63430000000
1!
1%
1-
12
15
#63440000000
0!
0%
b100 *
0-
02
b100 6
#63450000000
1!
1%
1-
12
#63460000000
0!
0%
b101 *
0-
02
b101 6
#63470000000
1!
1%
1-
12
#63480000000
0!
0%
b110 *
0-
02
b110 6
#63490000000
1!
1%
1-
12
#63500000000
0!
0%
b111 *
0-
02
b111 6
#63510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#63520000000
0!
0%
b0 *
0-
02
b0 6
#63530000000
1!
1%
1-
12
#63540000000
0!
0%
b1 *
0-
02
b1 6
#63550000000
1!
1%
1-
12
#63560000000
0!
0%
b10 *
0-
02
b10 6
#63570000000
1!
1%
1-
12
#63580000000
0!
0%
b11 *
0-
02
b11 6
#63590000000
1!
1%
1-
12
15
#63600000000
0!
0%
b100 *
0-
02
b100 6
#63610000000
1!
1%
1-
12
#63620000000
0!
0%
b101 *
0-
02
b101 6
#63630000000
1!
1%
1-
12
#63640000000
0!
0%
b110 *
0-
02
b110 6
#63650000000
1!
1%
1-
12
#63660000000
0!
0%
b111 *
0-
02
b111 6
#63670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#63680000000
0!
0%
b0 *
0-
02
b0 6
#63690000000
1!
1%
1-
12
#63700000000
0!
0%
b1 *
0-
02
b1 6
#63710000000
1!
1%
1-
12
#63720000000
0!
0%
b10 *
0-
02
b10 6
#63730000000
1!
1%
1-
12
#63740000000
0!
0%
b11 *
0-
02
b11 6
#63750000000
1!
1%
1-
12
15
#63760000000
0!
0%
b100 *
0-
02
b100 6
#63770000000
1!
1%
1-
12
#63780000000
0!
0%
b101 *
0-
02
b101 6
#63790000000
1!
1%
1-
12
#63800000000
0!
0%
b110 *
0-
02
b110 6
#63810000000
1!
1%
1-
12
#63820000000
0!
0%
b111 *
0-
02
b111 6
#63830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#63840000000
0!
0%
b0 *
0-
02
b0 6
#63850000000
1!
1%
1-
12
#63860000000
0!
0%
b1 *
0-
02
b1 6
#63870000000
1!
1%
1-
12
#63880000000
0!
0%
b10 *
0-
02
b10 6
#63890000000
1!
1%
1-
12
#63900000000
0!
0%
b11 *
0-
02
b11 6
#63910000000
1!
1%
1-
12
15
#63920000000
0!
0%
b100 *
0-
02
b100 6
#63930000000
1!
1%
1-
12
#63940000000
0!
0%
b101 *
0-
02
b101 6
#63950000000
1!
1%
1-
12
#63960000000
0!
0%
b110 *
0-
02
b110 6
#63970000000
1!
1%
1-
12
#63980000000
0!
0%
b111 *
0-
02
b111 6
#63990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#64000000000
0!
0%
b0 *
0-
02
b0 6
#64010000000
1!
1%
1-
12
#64020000000
0!
0%
b1 *
0-
02
b1 6
#64030000000
1!
1%
1-
12
#64040000000
0!
0%
b10 *
0-
02
b10 6
#64050000000
1!
1%
1-
12
#64060000000
0!
0%
b11 *
0-
02
b11 6
#64070000000
1!
1%
1-
12
15
#64080000000
0!
0%
b100 *
0-
02
b100 6
#64090000000
1!
1%
1-
12
#64100000000
0!
0%
b101 *
0-
02
b101 6
#64110000000
1!
1%
1-
12
#64120000000
0!
0%
b110 *
0-
02
b110 6
#64130000000
1!
1%
1-
12
#64140000000
0!
0%
b111 *
0-
02
b111 6
#64150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#64160000000
0!
0%
b0 *
0-
02
b0 6
#64170000000
1!
1%
1-
12
#64180000000
0!
0%
b1 *
0-
02
b1 6
#64190000000
1!
1%
1-
12
#64200000000
0!
0%
b10 *
0-
02
b10 6
#64210000000
1!
1%
1-
12
#64220000000
0!
0%
b11 *
0-
02
b11 6
#64230000000
1!
1%
1-
12
15
#64240000000
0!
0%
b100 *
0-
02
b100 6
#64250000000
1!
1%
1-
12
#64260000000
0!
0%
b101 *
0-
02
b101 6
#64270000000
1!
1%
1-
12
#64280000000
0!
0%
b110 *
0-
02
b110 6
#64290000000
1!
1%
1-
12
#64300000000
0!
0%
b111 *
0-
02
b111 6
#64310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#64320000000
0!
0%
b0 *
0-
02
b0 6
#64330000000
1!
1%
1-
12
#64340000000
0!
0%
b1 *
0-
02
b1 6
#64350000000
1!
1%
1-
12
#64360000000
0!
0%
b10 *
0-
02
b10 6
#64370000000
1!
1%
1-
12
#64380000000
0!
0%
b11 *
0-
02
b11 6
#64390000000
1!
1%
1-
12
15
#64400000000
0!
0%
b100 *
0-
02
b100 6
#64410000000
1!
1%
1-
12
#64420000000
0!
0%
b101 *
0-
02
b101 6
#64430000000
1!
1%
1-
12
#64440000000
0!
0%
b110 *
0-
02
b110 6
#64450000000
1!
1%
1-
12
#64460000000
0!
0%
b111 *
0-
02
b111 6
#64470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#64480000000
0!
0%
b0 *
0-
02
b0 6
#64490000000
1!
1%
1-
12
#64500000000
0!
0%
b1 *
0-
02
b1 6
#64510000000
1!
1%
1-
12
#64520000000
0!
0%
b10 *
0-
02
b10 6
#64530000000
1!
1%
1-
12
#64540000000
0!
0%
b11 *
0-
02
b11 6
#64550000000
1!
1%
1-
12
15
#64560000000
0!
0%
b100 *
0-
02
b100 6
#64570000000
1!
1%
1-
12
#64580000000
0!
0%
b101 *
0-
02
b101 6
#64590000000
1!
1%
1-
12
#64600000000
0!
0%
b110 *
0-
02
b110 6
#64610000000
1!
1%
1-
12
#64620000000
0!
0%
b111 *
0-
02
b111 6
#64630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#64640000000
0!
0%
b0 *
0-
02
b0 6
#64650000000
1!
1%
1-
12
#64660000000
0!
0%
b1 *
0-
02
b1 6
#64670000000
1!
1%
1-
12
#64680000000
0!
0%
b10 *
0-
02
b10 6
#64690000000
1!
1%
1-
12
#64700000000
0!
0%
b11 *
0-
02
b11 6
#64710000000
1!
1%
1-
12
15
#64720000000
0!
0%
b100 *
0-
02
b100 6
#64730000000
1!
1%
1-
12
#64740000000
0!
0%
b101 *
0-
02
b101 6
#64750000000
1!
1%
1-
12
#64760000000
0!
0%
b110 *
0-
02
b110 6
#64770000000
1!
1%
1-
12
#64780000000
0!
0%
b111 *
0-
02
b111 6
#64790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#64800000000
0!
0%
b0 *
0-
02
b0 6
#64810000000
1!
1%
1-
12
#64820000000
0!
0%
b1 *
0-
02
b1 6
#64830000000
1!
1%
1-
12
#64840000000
0!
0%
b10 *
0-
02
b10 6
#64850000000
1!
1%
1-
12
#64860000000
0!
0%
b11 *
0-
02
b11 6
#64870000000
1!
1%
1-
12
15
#64880000000
0!
0%
b100 *
0-
02
b100 6
#64890000000
1!
1%
1-
12
#64900000000
0!
0%
b101 *
0-
02
b101 6
#64910000000
1!
1%
1-
12
#64920000000
0!
0%
b110 *
0-
02
b110 6
#64930000000
1!
1%
1-
12
#64940000000
0!
0%
b111 *
0-
02
b111 6
#64950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#64960000000
0!
0%
b0 *
0-
02
b0 6
#64970000000
1!
1%
1-
12
#64980000000
0!
0%
b1 *
0-
02
b1 6
#64990000000
1!
1%
1-
12
#65000000000
0!
0%
b10 *
0-
02
b10 6
#65010000000
1!
1%
1-
12
#65020000000
0!
0%
b11 *
0-
02
b11 6
#65030000000
1!
1%
1-
12
15
#65040000000
0!
0%
b100 *
0-
02
b100 6
#65050000000
1!
1%
1-
12
#65060000000
0!
0%
b101 *
0-
02
b101 6
#65070000000
1!
1%
1-
12
#65080000000
0!
0%
b110 *
0-
02
b110 6
#65090000000
1!
1%
1-
12
#65100000000
0!
0%
b111 *
0-
02
b111 6
#65110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#65120000000
0!
0%
b0 *
0-
02
b0 6
#65130000000
1!
1%
1-
12
#65140000000
0!
0%
b1 *
0-
02
b1 6
#65150000000
1!
1%
1-
12
#65160000000
0!
0%
b10 *
0-
02
b10 6
#65170000000
1!
1%
1-
12
#65180000000
0!
0%
b11 *
0-
02
b11 6
#65190000000
1!
1%
1-
12
15
#65200000000
0!
0%
b100 *
0-
02
b100 6
#65210000000
1!
1%
1-
12
#65220000000
0!
0%
b101 *
0-
02
b101 6
#65230000000
1!
1%
1-
12
#65240000000
0!
0%
b110 *
0-
02
b110 6
#65250000000
1!
1%
1-
12
#65260000000
0!
0%
b111 *
0-
02
b111 6
#65270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#65280000000
0!
0%
b0 *
0-
02
b0 6
#65290000000
1!
1%
1-
12
#65300000000
0!
0%
b1 *
0-
02
b1 6
#65310000000
1!
1%
1-
12
#65320000000
0!
0%
b10 *
0-
02
b10 6
#65330000000
1!
1%
1-
12
#65340000000
0!
0%
b11 *
0-
02
b11 6
#65350000000
1!
1%
1-
12
15
#65360000000
0!
0%
b100 *
0-
02
b100 6
#65370000000
1!
1%
1-
12
#65380000000
0!
0%
b101 *
0-
02
b101 6
#65390000000
1!
1%
1-
12
#65400000000
0!
0%
b110 *
0-
02
b110 6
#65410000000
1!
1%
1-
12
#65420000000
0!
0%
b111 *
0-
02
b111 6
#65430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#65440000000
0!
0%
b0 *
0-
02
b0 6
#65450000000
1!
1%
1-
12
#65460000000
0!
0%
b1 *
0-
02
b1 6
#65470000000
1!
1%
1-
12
#65480000000
0!
0%
b10 *
0-
02
b10 6
#65490000000
1!
1%
1-
12
#65500000000
0!
0%
b11 *
0-
02
b11 6
#65510000000
1!
1%
1-
12
15
#65520000000
0!
0%
b100 *
0-
02
b100 6
#65530000000
1!
1%
1-
12
#65540000000
0!
0%
b101 *
0-
02
b101 6
#65550000000
1!
1%
1-
12
#65560000000
0!
0%
b110 *
0-
02
b110 6
#65570000000
1!
1%
1-
12
#65580000000
0!
0%
b111 *
0-
02
b111 6
#65590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#65600000000
0!
0%
b0 *
0-
02
b0 6
#65610000000
1!
1%
1-
12
#65620000000
0!
0%
b1 *
0-
02
b1 6
#65630000000
1!
1%
1-
12
#65640000000
0!
0%
b10 *
0-
02
b10 6
#65650000000
1!
1%
1-
12
#65660000000
0!
0%
b11 *
0-
02
b11 6
#65670000000
1!
1%
1-
12
15
#65680000000
0!
0%
b100 *
0-
02
b100 6
#65690000000
1!
1%
1-
12
#65700000000
0!
0%
b101 *
0-
02
b101 6
#65710000000
1!
1%
1-
12
#65720000000
0!
0%
b110 *
0-
02
b110 6
#65730000000
1!
1%
1-
12
#65740000000
0!
0%
b111 *
0-
02
b111 6
#65750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#65760000000
0!
0%
b0 *
0-
02
b0 6
#65770000000
1!
1%
1-
12
#65780000000
0!
0%
b1 *
0-
02
b1 6
#65790000000
1!
1%
1-
12
#65800000000
0!
0%
b10 *
0-
02
b10 6
#65810000000
1!
1%
1-
12
#65820000000
0!
0%
b11 *
0-
02
b11 6
#65830000000
1!
1%
1-
12
15
#65840000000
0!
0%
b100 *
0-
02
b100 6
#65850000000
1!
1%
1-
12
#65860000000
0!
0%
b101 *
0-
02
b101 6
#65870000000
1!
1%
1-
12
#65880000000
0!
0%
b110 *
0-
02
b110 6
#65890000000
1!
1%
1-
12
#65900000000
0!
0%
b111 *
0-
02
b111 6
#65910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#65920000000
0!
0%
b0 *
0-
02
b0 6
#65930000000
1!
1%
1-
12
#65940000000
0!
0%
b1 *
0-
02
b1 6
#65950000000
1!
1%
1-
12
#65960000000
0!
0%
b10 *
0-
02
b10 6
#65970000000
1!
1%
1-
12
#65980000000
0!
0%
b11 *
0-
02
b11 6
#65990000000
1!
1%
1-
12
15
#66000000000
0!
0%
b100 *
0-
02
b100 6
#66010000000
1!
1%
1-
12
#66020000000
0!
0%
b101 *
0-
02
b101 6
#66030000000
1!
1%
1-
12
#66040000000
0!
0%
b110 *
0-
02
b110 6
#66050000000
1!
1%
1-
12
#66060000000
0!
0%
b111 *
0-
02
b111 6
#66070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#66080000000
0!
0%
b0 *
0-
02
b0 6
#66090000000
1!
1%
1-
12
#66100000000
0!
0%
b1 *
0-
02
b1 6
#66110000000
1!
1%
1-
12
#66120000000
0!
0%
b10 *
0-
02
b10 6
#66130000000
1!
1%
1-
12
#66140000000
0!
0%
b11 *
0-
02
b11 6
#66150000000
1!
1%
1-
12
15
#66160000000
0!
0%
b100 *
0-
02
b100 6
#66170000000
1!
1%
1-
12
#66180000000
0!
0%
b101 *
0-
02
b101 6
#66190000000
1!
1%
1-
12
#66200000000
0!
0%
b110 *
0-
02
b110 6
#66210000000
1!
1%
1-
12
#66220000000
0!
0%
b111 *
0-
02
b111 6
#66230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#66240000000
0!
0%
b0 *
0-
02
b0 6
#66250000000
1!
1%
1-
12
#66260000000
0!
0%
b1 *
0-
02
b1 6
#66270000000
1!
1%
1-
12
#66280000000
0!
0%
b10 *
0-
02
b10 6
#66290000000
1!
1%
1-
12
#66300000000
0!
0%
b11 *
0-
02
b11 6
#66310000000
1!
1%
1-
12
15
#66320000000
0!
0%
b100 *
0-
02
b100 6
#66330000000
1!
1%
1-
12
#66340000000
0!
0%
b101 *
0-
02
b101 6
#66350000000
1!
1%
1-
12
#66360000000
0!
0%
b110 *
0-
02
b110 6
#66370000000
1!
1%
1-
12
#66380000000
0!
0%
b111 *
0-
02
b111 6
#66390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#66400000000
0!
0%
b0 *
0-
02
b0 6
#66410000000
1!
1%
1-
12
#66420000000
0!
0%
b1 *
0-
02
b1 6
#66430000000
1!
1%
1-
12
#66440000000
0!
0%
b10 *
0-
02
b10 6
#66450000000
1!
1%
1-
12
#66460000000
0!
0%
b11 *
0-
02
b11 6
#66470000000
1!
1%
1-
12
15
#66480000000
0!
0%
b100 *
0-
02
b100 6
#66490000000
1!
1%
1-
12
#66500000000
0!
0%
b101 *
0-
02
b101 6
#66510000000
1!
1%
1-
12
#66520000000
0!
0%
b110 *
0-
02
b110 6
#66530000000
1!
1%
1-
12
#66540000000
0!
0%
b111 *
0-
02
b111 6
#66550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#66560000000
0!
0%
b0 *
0-
02
b0 6
#66570000000
1!
1%
1-
12
#66580000000
0!
0%
b1 *
0-
02
b1 6
#66590000000
1!
1%
1-
12
#66600000000
0!
0%
b10 *
0-
02
b10 6
#66610000000
1!
1%
1-
12
#66620000000
0!
0%
b11 *
0-
02
b11 6
#66630000000
1!
1%
1-
12
15
#66640000000
0!
0%
b100 *
0-
02
b100 6
#66650000000
1!
1%
1-
12
#66660000000
0!
0%
b101 *
0-
02
b101 6
#66670000000
1!
1%
1-
12
#66680000000
0!
0%
b110 *
0-
02
b110 6
#66690000000
1!
1%
1-
12
#66700000000
0!
0%
b111 *
0-
02
b111 6
#66710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#66720000000
0!
0%
b0 *
0-
02
b0 6
#66730000000
1!
1%
1-
12
#66740000000
0!
0%
b1 *
0-
02
b1 6
#66750000000
1!
1%
1-
12
#66760000000
0!
0%
b10 *
0-
02
b10 6
#66770000000
1!
1%
1-
12
#66780000000
0!
0%
b11 *
0-
02
b11 6
#66790000000
1!
1%
1-
12
15
#66800000000
0!
0%
b100 *
0-
02
b100 6
#66810000000
1!
1%
1-
12
#66820000000
0!
0%
b101 *
0-
02
b101 6
#66830000000
1!
1%
1-
12
#66840000000
0!
0%
b110 *
0-
02
b110 6
#66850000000
1!
1%
1-
12
#66860000000
0!
0%
b111 *
0-
02
b111 6
#66870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#66880000000
0!
0%
b0 *
0-
02
b0 6
#66890000000
1!
1%
1-
12
#66900000000
0!
0%
b1 *
0-
02
b1 6
#66910000000
1!
1%
1-
12
#66920000000
0!
0%
b10 *
0-
02
b10 6
#66930000000
1!
1%
1-
12
#66940000000
0!
0%
b11 *
0-
02
b11 6
#66950000000
1!
1%
1-
12
15
#66960000000
0!
0%
b100 *
0-
02
b100 6
#66970000000
1!
1%
1-
12
#66980000000
0!
0%
b101 *
0-
02
b101 6
#66990000000
1!
1%
1-
12
#67000000000
0!
0%
b110 *
0-
02
b110 6
#67010000000
1!
1%
1-
12
#67020000000
0!
0%
b111 *
0-
02
b111 6
#67030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#67040000000
0!
0%
b0 *
0-
02
b0 6
#67050000000
1!
1%
1-
12
#67060000000
0!
0%
b1 *
0-
02
b1 6
#67070000000
1!
1%
1-
12
#67080000000
0!
0%
b10 *
0-
02
b10 6
#67090000000
1!
1%
1-
12
#67100000000
0!
0%
b11 *
0-
02
b11 6
#67110000000
1!
1%
1-
12
15
#67120000000
0!
0%
b100 *
0-
02
b100 6
#67130000000
1!
1%
1-
12
#67140000000
0!
0%
b101 *
0-
02
b101 6
#67150000000
1!
1%
1-
12
#67160000000
0!
0%
b110 *
0-
02
b110 6
#67170000000
1!
1%
1-
12
#67180000000
0!
0%
b111 *
0-
02
b111 6
#67190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#67200000000
0!
0%
b0 *
0-
02
b0 6
#67210000000
1!
1%
1-
12
#67220000000
0!
0%
b1 *
0-
02
b1 6
#67230000000
1!
1%
1-
12
#67240000000
0!
0%
b10 *
0-
02
b10 6
#67250000000
1!
1%
1-
12
#67260000000
0!
0%
b11 *
0-
02
b11 6
#67270000000
1!
1%
1-
12
15
#67280000000
0!
0%
b100 *
0-
02
b100 6
#67290000000
1!
1%
1-
12
#67300000000
0!
0%
b101 *
0-
02
b101 6
#67310000000
1!
1%
1-
12
#67320000000
0!
0%
b110 *
0-
02
b110 6
#67330000000
1!
1%
1-
12
#67340000000
0!
0%
b111 *
0-
02
b111 6
#67350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#67360000000
0!
0%
b0 *
0-
02
b0 6
#67370000000
1!
1%
1-
12
#67380000000
0!
0%
b1 *
0-
02
b1 6
#67390000000
1!
1%
1-
12
#67400000000
0!
0%
b10 *
0-
02
b10 6
#67410000000
1!
1%
1-
12
#67420000000
0!
0%
b11 *
0-
02
b11 6
#67430000000
1!
1%
1-
12
15
#67440000000
0!
0%
b100 *
0-
02
b100 6
#67450000000
1!
1%
1-
12
#67460000000
0!
0%
b101 *
0-
02
b101 6
#67470000000
1!
1%
1-
12
#67480000000
0!
0%
b110 *
0-
02
b110 6
#67490000000
1!
1%
1-
12
#67500000000
0!
0%
b111 *
0-
02
b111 6
#67510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#67520000000
0!
0%
b0 *
0-
02
b0 6
#67530000000
1!
1%
1-
12
#67540000000
0!
0%
b1 *
0-
02
b1 6
#67550000000
1!
1%
1-
12
#67560000000
0!
0%
b10 *
0-
02
b10 6
#67570000000
1!
1%
1-
12
#67580000000
0!
0%
b11 *
0-
02
b11 6
#67590000000
1!
1%
1-
12
15
#67600000000
0!
0%
b100 *
0-
02
b100 6
#67610000000
1!
1%
1-
12
#67620000000
0!
0%
b101 *
0-
02
b101 6
#67630000000
1!
1%
1-
12
#67640000000
0!
0%
b110 *
0-
02
b110 6
#67650000000
1!
1%
1-
12
#67660000000
0!
0%
b111 *
0-
02
b111 6
#67670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#67680000000
0!
0%
b0 *
0-
02
b0 6
#67690000000
1!
1%
1-
12
#67700000000
0!
0%
b1 *
0-
02
b1 6
#67710000000
1!
1%
1-
12
#67720000000
0!
0%
b10 *
0-
02
b10 6
#67730000000
1!
1%
1-
12
#67740000000
0!
0%
b11 *
0-
02
b11 6
#67750000000
1!
1%
1-
12
15
#67760000000
0!
0%
b100 *
0-
02
b100 6
#67770000000
1!
1%
1-
12
#67780000000
0!
0%
b101 *
0-
02
b101 6
#67790000000
1!
1%
1-
12
#67800000000
0!
0%
b110 *
0-
02
b110 6
#67810000000
1!
1%
1-
12
#67820000000
0!
0%
b111 *
0-
02
b111 6
#67830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#67840000000
0!
0%
b0 *
0-
02
b0 6
#67850000000
1!
1%
1-
12
#67860000000
0!
0%
b1 *
0-
02
b1 6
#67870000000
1!
1%
1-
12
#67880000000
0!
0%
b10 *
0-
02
b10 6
#67890000000
1!
1%
1-
12
#67900000000
0!
0%
b11 *
0-
02
b11 6
#67910000000
1!
1%
1-
12
15
#67920000000
0!
0%
b100 *
0-
02
b100 6
#67930000000
1!
1%
1-
12
#67940000000
0!
0%
b101 *
0-
02
b101 6
#67950000000
1!
1%
1-
12
#67960000000
0!
0%
b110 *
0-
02
b110 6
#67970000000
1!
1%
1-
12
#67980000000
0!
0%
b111 *
0-
02
b111 6
#67990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#68000000000
0!
0%
b0 *
0-
02
b0 6
#68010000000
1!
1%
1-
12
#68020000000
0!
0%
b1 *
0-
02
b1 6
#68030000000
1!
1%
1-
12
#68040000000
0!
0%
b10 *
0-
02
b10 6
#68050000000
1!
1%
1-
12
#68060000000
0!
0%
b11 *
0-
02
b11 6
#68070000000
1!
1%
1-
12
15
#68080000000
0!
0%
b100 *
0-
02
b100 6
#68090000000
1!
1%
1-
12
#68100000000
0!
0%
b101 *
0-
02
b101 6
#68110000000
1!
1%
1-
12
#68120000000
0!
0%
b110 *
0-
02
b110 6
#68130000000
1!
1%
1-
12
#68140000000
0!
0%
b111 *
0-
02
b111 6
#68150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#68160000000
0!
0%
b0 *
0-
02
b0 6
#68170000000
1!
1%
1-
12
#68180000000
0!
0%
b1 *
0-
02
b1 6
#68190000000
1!
1%
1-
12
#68200000000
0!
0%
b10 *
0-
02
b10 6
#68210000000
1!
1%
1-
12
#68220000000
0!
0%
b11 *
0-
02
b11 6
#68230000000
1!
1%
1-
12
15
#68240000000
0!
0%
b100 *
0-
02
b100 6
#68250000000
1!
1%
1-
12
#68260000000
0!
0%
b101 *
0-
02
b101 6
#68270000000
1!
1%
1-
12
#68280000000
0!
0%
b110 *
0-
02
b110 6
#68290000000
1!
1%
1-
12
#68300000000
0!
0%
b111 *
0-
02
b111 6
#68310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#68320000000
0!
0%
b0 *
0-
02
b0 6
#68330000000
1!
1%
1-
12
#68340000000
0!
0%
b1 *
0-
02
b1 6
#68350000000
1!
1%
1-
12
#68360000000
0!
0%
b10 *
0-
02
b10 6
#68370000000
1!
1%
1-
12
#68380000000
0!
0%
b11 *
0-
02
b11 6
#68390000000
1!
1%
1-
12
15
#68400000000
0!
0%
b100 *
0-
02
b100 6
#68410000000
1!
1%
1-
12
#68420000000
0!
0%
b101 *
0-
02
b101 6
#68430000000
1!
1%
1-
12
#68440000000
0!
0%
b110 *
0-
02
b110 6
#68450000000
1!
1%
1-
12
#68460000000
0!
0%
b111 *
0-
02
b111 6
#68470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#68480000000
0!
0%
b0 *
0-
02
b0 6
#68490000000
1!
1%
1-
12
#68500000000
0!
0%
b1 *
0-
02
b1 6
#68510000000
1!
1%
1-
12
#68520000000
0!
0%
b10 *
0-
02
b10 6
#68530000000
1!
1%
1-
12
#68540000000
0!
0%
b11 *
0-
02
b11 6
#68550000000
1!
1%
1-
12
15
#68560000000
0!
0%
b100 *
0-
02
b100 6
#68570000000
1!
1%
1-
12
#68580000000
0!
0%
b101 *
0-
02
b101 6
#68590000000
1!
1%
1-
12
#68600000000
0!
0%
b110 *
0-
02
b110 6
#68610000000
1!
1%
1-
12
#68620000000
0!
0%
b111 *
0-
02
b111 6
#68630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#68640000000
0!
0%
b0 *
0-
02
b0 6
#68650000000
1!
1%
1-
12
#68660000000
0!
0%
b1 *
0-
02
b1 6
#68670000000
1!
1%
1-
12
#68680000000
0!
0%
b10 *
0-
02
b10 6
#68690000000
1!
1%
1-
12
#68700000000
0!
0%
b11 *
0-
02
b11 6
#68710000000
1!
1%
1-
12
15
#68720000000
0!
0%
b100 *
0-
02
b100 6
#68730000000
1!
1%
1-
12
#68740000000
0!
0%
b101 *
0-
02
b101 6
#68750000000
1!
1%
1-
12
#68760000000
0!
0%
b110 *
0-
02
b110 6
#68770000000
1!
1%
1-
12
#68780000000
0!
0%
b111 *
0-
02
b111 6
#68790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#68800000000
0!
0%
b0 *
0-
02
b0 6
#68810000000
1!
1%
1-
12
#68820000000
0!
0%
b1 *
0-
02
b1 6
#68830000000
1!
1%
1-
12
#68840000000
0!
0%
b10 *
0-
02
b10 6
#68850000000
1!
1%
1-
12
#68860000000
0!
0%
b11 *
0-
02
b11 6
#68870000000
1!
1%
1-
12
15
#68880000000
0!
0%
b100 *
0-
02
b100 6
#68890000000
1!
1%
1-
12
#68900000000
0!
0%
b101 *
0-
02
b101 6
#68910000000
1!
1%
1-
12
#68920000000
0!
0%
b110 *
0-
02
b110 6
#68930000000
1!
1%
1-
12
#68940000000
0!
0%
b111 *
0-
02
b111 6
#68950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#68960000000
0!
0%
b0 *
0-
02
b0 6
#68970000000
1!
1%
1-
12
#68980000000
0!
0%
b1 *
0-
02
b1 6
#68990000000
1!
1%
1-
12
#69000000000
0!
0%
b10 *
0-
02
b10 6
#69010000000
1!
1%
1-
12
#69020000000
0!
0%
b11 *
0-
02
b11 6
#69030000000
1!
1%
1-
12
15
#69040000000
0!
0%
b100 *
0-
02
b100 6
#69050000000
1!
1%
1-
12
#69060000000
0!
0%
b101 *
0-
02
b101 6
#69070000000
1!
1%
1-
12
#69080000000
0!
0%
b110 *
0-
02
b110 6
#69090000000
1!
1%
1-
12
#69100000000
0!
0%
b111 *
0-
02
b111 6
#69110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#69120000000
0!
0%
b0 *
0-
02
b0 6
#69130000000
1!
1%
1-
12
#69140000000
0!
0%
b1 *
0-
02
b1 6
#69150000000
1!
1%
1-
12
#69160000000
0!
0%
b10 *
0-
02
b10 6
#69170000000
1!
1%
1-
12
#69180000000
0!
0%
b11 *
0-
02
b11 6
#69190000000
1!
1%
1-
12
15
#69200000000
0!
0%
b100 *
0-
02
b100 6
#69210000000
1!
1%
1-
12
#69220000000
0!
0%
b101 *
0-
02
b101 6
#69230000000
1!
1%
1-
12
#69240000000
0!
0%
b110 *
0-
02
b110 6
#69250000000
1!
1%
1-
12
#69260000000
0!
0%
b111 *
0-
02
b111 6
#69270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#69280000000
0!
0%
b0 *
0-
02
b0 6
#69290000000
1!
1%
1-
12
#69300000000
0!
0%
b1 *
0-
02
b1 6
#69310000000
1!
1%
1-
12
#69320000000
0!
0%
b10 *
0-
02
b10 6
#69330000000
1!
1%
1-
12
#69340000000
0!
0%
b11 *
0-
02
b11 6
#69350000000
1!
1%
1-
12
15
#69360000000
0!
0%
b100 *
0-
02
b100 6
#69370000000
1!
1%
1-
12
#69380000000
0!
0%
b101 *
0-
02
b101 6
#69390000000
1!
1%
1-
12
#69400000000
0!
0%
b110 *
0-
02
b110 6
#69410000000
1!
1%
1-
12
#69420000000
0!
0%
b111 *
0-
02
b111 6
#69430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#69440000000
0!
0%
b0 *
0-
02
b0 6
#69450000000
1!
1%
1-
12
#69460000000
0!
0%
b1 *
0-
02
b1 6
#69470000000
1!
1%
1-
12
#69480000000
0!
0%
b10 *
0-
02
b10 6
#69490000000
1!
1%
1-
12
#69500000000
0!
0%
b11 *
0-
02
b11 6
#69510000000
1!
1%
1-
12
15
#69520000000
0!
0%
b100 *
0-
02
b100 6
#69530000000
1!
1%
1-
12
#69540000000
0!
0%
b101 *
0-
02
b101 6
#69550000000
1!
1%
1-
12
#69560000000
0!
0%
b110 *
0-
02
b110 6
#69570000000
1!
1%
1-
12
#69580000000
0!
0%
b111 *
0-
02
b111 6
#69590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#69600000000
0!
0%
b0 *
0-
02
b0 6
#69610000000
1!
1%
1-
12
#69620000000
0!
0%
b1 *
0-
02
b1 6
#69630000000
1!
1%
1-
12
#69640000000
0!
0%
b10 *
0-
02
b10 6
#69650000000
1!
1%
1-
12
#69660000000
0!
0%
b11 *
0-
02
b11 6
#69670000000
1!
1%
1-
12
15
#69680000000
0!
0%
b100 *
0-
02
b100 6
#69690000000
1!
1%
1-
12
#69700000000
0!
0%
b101 *
0-
02
b101 6
#69710000000
1!
1%
1-
12
#69720000000
0!
0%
b110 *
0-
02
b110 6
#69730000000
1!
1%
1-
12
#69740000000
0!
0%
b111 *
0-
02
b111 6
#69750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#69760000000
0!
0%
b0 *
0-
02
b0 6
#69770000000
1!
1%
1-
12
#69780000000
0!
0%
b1 *
0-
02
b1 6
#69790000000
1!
1%
1-
12
#69800000000
0!
0%
b10 *
0-
02
b10 6
#69810000000
1!
1%
1-
12
#69820000000
0!
0%
b11 *
0-
02
b11 6
#69830000000
1!
1%
1-
12
15
#69840000000
0!
0%
b100 *
0-
02
b100 6
#69850000000
1!
1%
1-
12
#69860000000
0!
0%
b101 *
0-
02
b101 6
#69870000000
1!
1%
1-
12
#69880000000
0!
0%
b110 *
0-
02
b110 6
#69890000000
1!
1%
1-
12
#69900000000
0!
0%
b111 *
0-
02
b111 6
#69910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#69920000000
0!
0%
b0 *
0-
02
b0 6
#69930000000
1!
1%
1-
12
#69940000000
0!
0%
b1 *
0-
02
b1 6
#69950000000
1!
1%
1-
12
#69960000000
0!
0%
b10 *
0-
02
b10 6
#69970000000
1!
1%
1-
12
#69980000000
0!
0%
b11 *
0-
02
b11 6
#69990000000
1!
1%
1-
12
15
#70000000000
0!
0%
b100 *
0-
02
b100 6
#70010000000
1!
1%
1-
12
#70020000000
0!
0%
b101 *
0-
02
b101 6
#70030000000
1!
1%
1-
12
#70040000000
0!
0%
b110 *
0-
02
b110 6
#70050000000
1!
1%
1-
12
#70060000000
0!
0%
b111 *
0-
02
b111 6
#70070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#70080000000
0!
0%
b0 *
0-
02
b0 6
#70090000000
1!
1%
1-
12
#70100000000
0!
0%
b1 *
0-
02
b1 6
#70110000000
1!
1%
1-
12
#70120000000
0!
0%
b10 *
0-
02
b10 6
#70130000000
1!
1%
1-
12
#70140000000
0!
0%
b11 *
0-
02
b11 6
#70150000000
1!
1%
1-
12
15
#70160000000
0!
0%
b100 *
0-
02
b100 6
#70170000000
1!
1%
1-
12
#70180000000
0!
0%
b101 *
0-
02
b101 6
#70190000000
1!
1%
1-
12
#70200000000
0!
0%
b110 *
0-
02
b110 6
#70210000000
1!
1%
1-
12
#70220000000
0!
0%
b111 *
0-
02
b111 6
#70230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#70240000000
0!
0%
b0 *
0-
02
b0 6
#70250000000
1!
1%
1-
12
#70260000000
0!
0%
b1 *
0-
02
b1 6
#70270000000
1!
1%
1-
12
#70280000000
0!
0%
b10 *
0-
02
b10 6
#70290000000
1!
1%
1-
12
#70300000000
0!
0%
b11 *
0-
02
b11 6
#70310000000
1!
1%
1-
12
15
#70320000000
0!
0%
b100 *
0-
02
b100 6
#70330000000
1!
1%
1-
12
#70340000000
0!
0%
b101 *
0-
02
b101 6
#70350000000
1!
1%
1-
12
#70360000000
0!
0%
b110 *
0-
02
b110 6
#70370000000
1!
1%
1-
12
#70380000000
0!
0%
b111 *
0-
02
b111 6
#70390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#70400000000
0!
0%
b0 *
0-
02
b0 6
#70410000000
1!
1%
1-
12
#70420000000
0!
0%
b1 *
0-
02
b1 6
#70430000000
1!
1%
1-
12
#70440000000
0!
0%
b10 *
0-
02
b10 6
#70450000000
1!
1%
1-
12
#70460000000
0!
0%
b11 *
0-
02
b11 6
#70470000000
1!
1%
1-
12
15
#70480000000
0!
0%
b100 *
0-
02
b100 6
#70490000000
1!
1%
1-
12
#70500000000
0!
0%
b101 *
0-
02
b101 6
#70510000000
1!
1%
1-
12
#70520000000
0!
0%
b110 *
0-
02
b110 6
#70530000000
1!
1%
1-
12
#70540000000
0!
0%
b111 *
0-
02
b111 6
#70550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#70560000000
0!
0%
b0 *
0-
02
b0 6
#70570000000
1!
1%
1-
12
#70580000000
0!
0%
b1 *
0-
02
b1 6
#70590000000
1!
1%
1-
12
#70600000000
0!
0%
b10 *
0-
02
b10 6
#70610000000
1!
1%
1-
12
#70620000000
0!
0%
b11 *
0-
02
b11 6
#70630000000
1!
1%
1-
12
15
#70640000000
0!
0%
b100 *
0-
02
b100 6
#70650000000
1!
1%
1-
12
#70660000000
0!
0%
b101 *
0-
02
b101 6
#70670000000
1!
1%
1-
12
#70680000000
0!
0%
b110 *
0-
02
b110 6
#70690000000
1!
1%
1-
12
#70700000000
0!
0%
b111 *
0-
02
b111 6
#70710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#70720000000
0!
0%
b0 *
0-
02
b0 6
#70730000000
1!
1%
1-
12
#70740000000
0!
0%
b1 *
0-
02
b1 6
#70750000000
1!
1%
1-
12
#70760000000
0!
0%
b10 *
0-
02
b10 6
#70770000000
1!
1%
1-
12
#70780000000
0!
0%
b11 *
0-
02
b11 6
#70790000000
1!
1%
1-
12
15
#70800000000
0!
0%
b100 *
0-
02
b100 6
#70810000000
1!
1%
1-
12
#70820000000
0!
0%
b101 *
0-
02
b101 6
#70830000000
1!
1%
1-
12
#70840000000
0!
0%
b110 *
0-
02
b110 6
#70850000000
1!
1%
1-
12
#70860000000
0!
0%
b111 *
0-
02
b111 6
#70870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#70880000000
0!
0%
b0 *
0-
02
b0 6
#70890000000
1!
1%
1-
12
#70900000000
0!
0%
b1 *
0-
02
b1 6
#70910000000
1!
1%
1-
12
#70920000000
0!
0%
b10 *
0-
02
b10 6
#70930000000
1!
1%
1-
12
#70940000000
0!
0%
b11 *
0-
02
b11 6
#70950000000
1!
1%
1-
12
15
#70960000000
0!
0%
b100 *
0-
02
b100 6
#70970000000
1!
1%
1-
12
#70980000000
0!
0%
b101 *
0-
02
b101 6
#70990000000
1!
1%
1-
12
#71000000000
0!
0%
b110 *
0-
02
b110 6
#71010000000
1!
1%
1-
12
#71020000000
0!
0%
b111 *
0-
02
b111 6
#71030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#71040000000
0!
0%
b0 *
0-
02
b0 6
#71050000000
1!
1%
1-
12
#71060000000
0!
0%
b1 *
0-
02
b1 6
#71070000000
1!
1%
1-
12
#71080000000
0!
0%
b10 *
0-
02
b10 6
#71090000000
1!
1%
1-
12
#71100000000
0!
0%
b11 *
0-
02
b11 6
#71110000000
1!
1%
1-
12
15
#71120000000
0!
0%
b100 *
0-
02
b100 6
#71130000000
1!
1%
1-
12
#71140000000
0!
0%
b101 *
0-
02
b101 6
#71150000000
1!
1%
1-
12
#71160000000
0!
0%
b110 *
0-
02
b110 6
#71170000000
1!
1%
1-
12
#71180000000
0!
0%
b111 *
0-
02
b111 6
#71190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#71200000000
0!
0%
b0 *
0-
02
b0 6
#71210000000
1!
1%
1-
12
#71220000000
0!
0%
b1 *
0-
02
b1 6
#71230000000
1!
1%
1-
12
#71240000000
0!
0%
b10 *
0-
02
b10 6
#71250000000
1!
1%
1-
12
#71260000000
0!
0%
b11 *
0-
02
b11 6
#71270000000
1!
1%
1-
12
15
#71280000000
0!
0%
b100 *
0-
02
b100 6
#71290000000
1!
1%
1-
12
#71300000000
0!
0%
b101 *
0-
02
b101 6
#71310000000
1!
1%
1-
12
#71320000000
0!
0%
b110 *
0-
02
b110 6
#71330000000
1!
1%
1-
12
#71340000000
0!
0%
b111 *
0-
02
b111 6
#71350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#71360000000
0!
0%
b0 *
0-
02
b0 6
#71370000000
1!
1%
1-
12
#71380000000
0!
0%
b1 *
0-
02
b1 6
#71390000000
1!
1%
1-
12
#71400000000
0!
0%
b10 *
0-
02
b10 6
#71410000000
1!
1%
1-
12
#71420000000
0!
0%
b11 *
0-
02
b11 6
#71430000000
1!
1%
1-
12
15
#71440000000
0!
0%
b100 *
0-
02
b100 6
#71450000000
1!
1%
1-
12
#71460000000
0!
0%
b101 *
0-
02
b101 6
#71470000000
1!
1%
1-
12
#71480000000
0!
0%
b110 *
0-
02
b110 6
#71490000000
1!
1%
1-
12
#71500000000
0!
0%
b111 *
0-
02
b111 6
#71510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#71520000000
0!
0%
b0 *
0-
02
b0 6
#71530000000
1!
1%
1-
12
#71540000000
0!
0%
b1 *
0-
02
b1 6
#71550000000
1!
1%
1-
12
#71560000000
0!
0%
b10 *
0-
02
b10 6
#71570000000
1!
1%
1-
12
#71580000000
0!
0%
b11 *
0-
02
b11 6
#71590000000
1!
1%
1-
12
15
#71600000000
0!
0%
b100 *
0-
02
b100 6
#71610000000
1!
1%
1-
12
#71620000000
0!
0%
b101 *
0-
02
b101 6
#71630000000
1!
1%
1-
12
#71640000000
0!
0%
b110 *
0-
02
b110 6
#71650000000
1!
1%
1-
12
#71660000000
0!
0%
b111 *
0-
02
b111 6
#71670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#71680000000
0!
0%
b0 *
0-
02
b0 6
#71690000000
1!
1%
1-
12
#71700000000
0!
0%
b1 *
0-
02
b1 6
#71710000000
1!
1%
1-
12
#71720000000
0!
0%
b10 *
0-
02
b10 6
#71730000000
1!
1%
1-
12
#71740000000
0!
0%
b11 *
0-
02
b11 6
#71750000000
1!
1%
1-
12
15
#71760000000
0!
0%
b100 *
0-
02
b100 6
#71770000000
1!
1%
1-
12
#71780000000
0!
0%
b101 *
0-
02
b101 6
#71790000000
1!
1%
1-
12
#71800000000
0!
0%
b110 *
0-
02
b110 6
#71810000000
1!
1%
1-
12
#71820000000
0!
0%
b111 *
0-
02
b111 6
#71830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#71840000000
0!
0%
b0 *
0-
02
b0 6
#71850000000
1!
1%
1-
12
#71860000000
0!
0%
b1 *
0-
02
b1 6
#71870000000
1!
1%
1-
12
#71880000000
0!
0%
b10 *
0-
02
b10 6
#71890000000
1!
1%
1-
12
#71900000000
0!
0%
b11 *
0-
02
b11 6
#71910000000
1!
1%
1-
12
15
#71920000000
0!
0%
b100 *
0-
02
b100 6
#71930000000
1!
1%
1-
12
#71940000000
0!
0%
b101 *
0-
02
b101 6
#71950000000
1!
1%
1-
12
#71960000000
0!
0%
b110 *
0-
02
b110 6
#71970000000
1!
1%
1-
12
#71980000000
0!
0%
b111 *
0-
02
b111 6
#71990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#72000000000
0!
0%
b0 *
0-
02
b0 6
#72010000000
1!
1%
1-
12
#72020000000
0!
0%
b1 *
0-
02
b1 6
#72030000000
1!
1%
1-
12
#72040000000
0!
0%
b10 *
0-
02
b10 6
#72050000000
1!
1%
1-
12
#72060000000
0!
0%
b11 *
0-
02
b11 6
#72070000000
1!
1%
1-
12
15
#72080000000
0!
0%
b100 *
0-
02
b100 6
#72090000000
1!
1%
1-
12
#72100000000
0!
0%
b101 *
0-
02
b101 6
#72110000000
1!
1%
1-
12
#72120000000
0!
0%
b110 *
0-
02
b110 6
#72130000000
1!
1%
1-
12
#72140000000
0!
0%
b111 *
0-
02
b111 6
#72150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#72160000000
0!
0%
b0 *
0-
02
b0 6
#72170000000
1!
1%
1-
12
#72180000000
0!
0%
b1 *
0-
02
b1 6
#72190000000
1!
1%
1-
12
#72200000000
0!
0%
b10 *
0-
02
b10 6
#72210000000
1!
1%
1-
12
#72220000000
0!
0%
b11 *
0-
02
b11 6
#72230000000
1!
1%
1-
12
15
#72240000000
0!
0%
b100 *
0-
02
b100 6
#72250000000
1!
1%
1-
12
#72260000000
0!
0%
b101 *
0-
02
b101 6
#72270000000
1!
1%
1-
12
#72280000000
0!
0%
b110 *
0-
02
b110 6
#72290000000
1!
1%
1-
12
#72300000000
0!
0%
b111 *
0-
02
b111 6
#72310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#72320000000
0!
0%
b0 *
0-
02
b0 6
#72330000000
1!
1%
1-
12
#72340000000
0!
0%
b1 *
0-
02
b1 6
#72350000000
1!
1%
1-
12
#72360000000
0!
0%
b10 *
0-
02
b10 6
#72370000000
1!
1%
1-
12
#72380000000
0!
0%
b11 *
0-
02
b11 6
#72390000000
1!
1%
1-
12
15
#72400000000
0!
0%
b100 *
0-
02
b100 6
#72410000000
1!
1%
1-
12
#72420000000
0!
0%
b101 *
0-
02
b101 6
#72430000000
1!
1%
1-
12
#72440000000
0!
0%
b110 *
0-
02
b110 6
#72450000000
1!
1%
1-
12
#72460000000
0!
0%
b111 *
0-
02
b111 6
#72470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#72480000000
0!
0%
b0 *
0-
02
b0 6
#72490000000
1!
1%
1-
12
#72500000000
0!
0%
b1 *
0-
02
b1 6
#72510000000
1!
1%
1-
12
#72520000000
0!
0%
b10 *
0-
02
b10 6
#72530000000
1!
1%
1-
12
#72540000000
0!
0%
b11 *
0-
02
b11 6
#72550000000
1!
1%
1-
12
15
#72560000000
0!
0%
b100 *
0-
02
b100 6
#72570000000
1!
1%
1-
12
#72580000000
0!
0%
b101 *
0-
02
b101 6
#72590000000
1!
1%
1-
12
#72600000000
0!
0%
b110 *
0-
02
b110 6
#72610000000
1!
1%
1-
12
#72620000000
0!
0%
b111 *
0-
02
b111 6
#72630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#72640000000
0!
0%
b0 *
0-
02
b0 6
#72650000000
1!
1%
1-
12
#72660000000
0!
0%
b1 *
0-
02
b1 6
#72670000000
1!
1%
1-
12
#72680000000
0!
0%
b10 *
0-
02
b10 6
#72690000000
1!
1%
1-
12
#72700000000
0!
0%
b11 *
0-
02
b11 6
#72710000000
1!
1%
1-
12
15
#72720000000
0!
0%
b100 *
0-
02
b100 6
#72730000000
1!
1%
1-
12
#72740000000
0!
0%
b101 *
0-
02
b101 6
#72750000000
1!
1%
1-
12
#72760000000
0!
0%
b110 *
0-
02
b110 6
#72770000000
1!
1%
1-
12
#72780000000
0!
0%
b111 *
0-
02
b111 6
#72790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#72800000000
0!
0%
b0 *
0-
02
b0 6
#72810000000
1!
1%
1-
12
#72820000000
0!
0%
b1 *
0-
02
b1 6
#72830000000
1!
1%
1-
12
#72840000000
0!
0%
b10 *
0-
02
b10 6
#72850000000
1!
1%
1-
12
#72860000000
0!
0%
b11 *
0-
02
b11 6
#72870000000
1!
1%
1-
12
15
#72880000000
0!
0%
b100 *
0-
02
b100 6
#72890000000
1!
1%
1-
12
#72900000000
0!
0%
b101 *
0-
02
b101 6
#72910000000
1!
1%
1-
12
#72920000000
0!
0%
b110 *
0-
02
b110 6
#72930000000
1!
1%
1-
12
#72940000000
0!
0%
b111 *
0-
02
b111 6
#72950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#72960000000
0!
0%
b0 *
0-
02
b0 6
#72970000000
1!
1%
1-
12
#72980000000
0!
0%
b1 *
0-
02
b1 6
#72990000000
1!
1%
1-
12
#73000000000
0!
0%
b10 *
0-
02
b10 6
#73010000000
1!
1%
1-
12
#73020000000
0!
0%
b11 *
0-
02
b11 6
#73030000000
1!
1%
1-
12
15
#73040000000
0!
0%
b100 *
0-
02
b100 6
#73050000000
1!
1%
1-
12
#73060000000
0!
0%
b101 *
0-
02
b101 6
#73070000000
1!
1%
1-
12
#73080000000
0!
0%
b110 *
0-
02
b110 6
#73090000000
1!
1%
1-
12
#73100000000
0!
0%
b111 *
0-
02
b111 6
#73110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#73120000000
0!
0%
b0 *
0-
02
b0 6
#73130000000
1!
1%
1-
12
#73140000000
0!
0%
b1 *
0-
02
b1 6
#73150000000
1!
1%
1-
12
#73160000000
0!
0%
b10 *
0-
02
b10 6
#73170000000
1!
1%
1-
12
#73180000000
0!
0%
b11 *
0-
02
b11 6
#73190000000
1!
1%
1-
12
15
#73200000000
0!
0%
b100 *
0-
02
b100 6
#73210000000
1!
1%
1-
12
#73220000000
0!
0%
b101 *
0-
02
b101 6
#73230000000
1!
1%
1-
12
#73240000000
0!
0%
b110 *
0-
02
b110 6
#73250000000
1!
1%
1-
12
#73260000000
0!
0%
b111 *
0-
02
b111 6
#73270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#73280000000
0!
0%
b0 *
0-
02
b0 6
#73290000000
1!
1%
1-
12
#73300000000
0!
0%
b1 *
0-
02
b1 6
#73310000000
1!
1%
1-
12
#73320000000
0!
0%
b10 *
0-
02
b10 6
#73330000000
1!
1%
1-
12
#73340000000
0!
0%
b11 *
0-
02
b11 6
#73350000000
1!
1%
1-
12
15
#73360000000
0!
0%
b100 *
0-
02
b100 6
#73370000000
1!
1%
1-
12
#73380000000
0!
0%
b101 *
0-
02
b101 6
#73390000000
1!
1%
1-
12
#73400000000
0!
0%
b110 *
0-
02
b110 6
#73410000000
1!
1%
1-
12
#73420000000
0!
0%
b111 *
0-
02
b111 6
#73430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#73440000000
0!
0%
b0 *
0-
02
b0 6
#73450000000
1!
1%
1-
12
#73460000000
0!
0%
b1 *
0-
02
b1 6
#73470000000
1!
1%
1-
12
#73480000000
0!
0%
b10 *
0-
02
b10 6
#73490000000
1!
1%
1-
12
#73500000000
0!
0%
b11 *
0-
02
b11 6
#73510000000
1!
1%
1-
12
15
#73520000000
0!
0%
b100 *
0-
02
b100 6
#73530000000
1!
1%
1-
12
#73540000000
0!
0%
b101 *
0-
02
b101 6
#73550000000
1!
1%
1-
12
#73560000000
0!
0%
b110 *
0-
02
b110 6
#73570000000
1!
1%
1-
12
#73580000000
0!
0%
b111 *
0-
02
b111 6
#73590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#73600000000
0!
0%
b0 *
0-
02
b0 6
#73610000000
1!
1%
1-
12
#73620000000
0!
0%
b1 *
0-
02
b1 6
#73630000000
1!
1%
1-
12
#73640000000
0!
0%
b10 *
0-
02
b10 6
#73650000000
1!
1%
1-
12
#73660000000
0!
0%
b11 *
0-
02
b11 6
#73670000000
1!
1%
1-
12
15
#73680000000
0!
0%
b100 *
0-
02
b100 6
#73690000000
1!
1%
1-
12
#73700000000
0!
0%
b101 *
0-
02
b101 6
#73710000000
1!
1%
1-
12
#73720000000
0!
0%
b110 *
0-
02
b110 6
#73730000000
1!
1%
1-
12
#73740000000
0!
0%
b111 *
0-
02
b111 6
#73750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#73760000000
0!
0%
b0 *
0-
02
b0 6
#73770000000
1!
1%
1-
12
#73780000000
0!
0%
b1 *
0-
02
b1 6
#73790000000
1!
1%
1-
12
#73800000000
0!
0%
b10 *
0-
02
b10 6
#73810000000
1!
1%
1-
12
#73820000000
0!
0%
b11 *
0-
02
b11 6
#73830000000
1!
1%
1-
12
15
#73840000000
0!
0%
b100 *
0-
02
b100 6
#73850000000
1!
1%
1-
12
#73860000000
0!
0%
b101 *
0-
02
b101 6
#73870000000
1!
1%
1-
12
#73880000000
0!
0%
b110 *
0-
02
b110 6
#73890000000
1!
1%
1-
12
#73900000000
0!
0%
b111 *
0-
02
b111 6
#73910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#73920000000
0!
0%
b0 *
0-
02
b0 6
#73930000000
1!
1%
1-
12
#73940000000
0!
0%
b1 *
0-
02
b1 6
#73950000000
1!
1%
1-
12
#73960000000
0!
0%
b10 *
0-
02
b10 6
#73970000000
1!
1%
1-
12
#73980000000
0!
0%
b11 *
0-
02
b11 6
#73990000000
1!
1%
1-
12
15
#74000000000
0!
0%
b100 *
0-
02
b100 6
#74010000000
1!
1%
1-
12
#74020000000
0!
0%
b101 *
0-
02
b101 6
#74030000000
1!
1%
1-
12
#74040000000
0!
0%
b110 *
0-
02
b110 6
#74050000000
1!
1%
1-
12
#74060000000
0!
0%
b111 *
0-
02
b111 6
#74070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#74080000000
0!
0%
b0 *
0-
02
b0 6
#74090000000
1!
1%
1-
12
#74100000000
0!
0%
b1 *
0-
02
b1 6
#74110000000
1!
1%
1-
12
#74120000000
0!
0%
b10 *
0-
02
b10 6
#74130000000
1!
1%
1-
12
#74140000000
0!
0%
b11 *
0-
02
b11 6
#74150000000
1!
1%
1-
12
15
#74160000000
0!
0%
b100 *
0-
02
b100 6
#74170000000
1!
1%
1-
12
#74180000000
0!
0%
b101 *
0-
02
b101 6
#74190000000
1!
1%
1-
12
#74200000000
0!
0%
b110 *
0-
02
b110 6
#74210000000
1!
1%
1-
12
#74220000000
0!
0%
b111 *
0-
02
b111 6
#74230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#74240000000
0!
0%
b0 *
0-
02
b0 6
#74250000000
1!
1%
1-
12
#74260000000
0!
0%
b1 *
0-
02
b1 6
#74270000000
1!
1%
1-
12
#74280000000
0!
0%
b10 *
0-
02
b10 6
#74290000000
1!
1%
1-
12
#74300000000
0!
0%
b11 *
0-
02
b11 6
#74310000000
1!
1%
1-
12
15
#74320000000
0!
0%
b100 *
0-
02
b100 6
#74330000000
1!
1%
1-
12
#74340000000
0!
0%
b101 *
0-
02
b101 6
#74350000000
1!
1%
1-
12
#74360000000
0!
0%
b110 *
0-
02
b110 6
#74370000000
1!
1%
1-
12
#74380000000
0!
0%
b111 *
0-
02
b111 6
#74390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#74400000000
0!
0%
b0 *
0-
02
b0 6
#74410000000
1!
1%
1-
12
#74420000000
0!
0%
b1 *
0-
02
b1 6
#74430000000
1!
1%
1-
12
#74440000000
0!
0%
b10 *
0-
02
b10 6
#74450000000
1!
1%
1-
12
#74460000000
0!
0%
b11 *
0-
02
b11 6
#74470000000
1!
1%
1-
12
15
#74480000000
0!
0%
b100 *
0-
02
b100 6
#74490000000
1!
1%
1-
12
#74500000000
0!
0%
b101 *
0-
02
b101 6
#74510000000
1!
1%
1-
12
#74520000000
0!
0%
b110 *
0-
02
b110 6
#74530000000
1!
1%
1-
12
#74540000000
0!
0%
b111 *
0-
02
b111 6
#74550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#74560000000
0!
0%
b0 *
0-
02
b0 6
#74570000000
1!
1%
1-
12
#74580000000
0!
0%
b1 *
0-
02
b1 6
#74590000000
1!
1%
1-
12
#74600000000
0!
0%
b10 *
0-
02
b10 6
#74610000000
1!
1%
1-
12
#74620000000
0!
0%
b11 *
0-
02
b11 6
#74630000000
1!
1%
1-
12
15
#74640000000
0!
0%
b100 *
0-
02
b100 6
#74650000000
1!
1%
1-
12
#74660000000
0!
0%
b101 *
0-
02
b101 6
#74670000000
1!
1%
1-
12
#74680000000
0!
0%
b110 *
0-
02
b110 6
#74690000000
1!
1%
1-
12
#74700000000
0!
0%
b111 *
0-
02
b111 6
#74710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#74720000000
0!
0%
b0 *
0-
02
b0 6
#74730000000
1!
1%
1-
12
#74740000000
0!
0%
b1 *
0-
02
b1 6
#74750000000
1!
1%
1-
12
#74760000000
0!
0%
b10 *
0-
02
b10 6
#74770000000
1!
1%
1-
12
#74780000000
0!
0%
b11 *
0-
02
b11 6
#74790000000
1!
1%
1-
12
15
#74800000000
0!
0%
b100 *
0-
02
b100 6
#74810000000
1!
1%
1-
12
#74820000000
0!
0%
b101 *
0-
02
b101 6
#74830000000
1!
1%
1-
12
#74840000000
0!
0%
b110 *
0-
02
b110 6
#74850000000
1!
1%
1-
12
#74860000000
0!
0%
b111 *
0-
02
b111 6
#74870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#74880000000
0!
0%
b0 *
0-
02
b0 6
#74890000000
1!
1%
1-
12
#74900000000
0!
0%
b1 *
0-
02
b1 6
#74910000000
1!
1%
1-
12
#74920000000
0!
0%
b10 *
0-
02
b10 6
#74930000000
1!
1%
1-
12
#74940000000
0!
0%
b11 *
0-
02
b11 6
#74950000000
1!
1%
1-
12
15
#74960000000
0!
0%
b100 *
0-
02
b100 6
#74970000000
1!
1%
1-
12
#74980000000
0!
0%
b101 *
0-
02
b101 6
#74990000000
1!
1%
1-
12
#75000000000
0!
0%
b110 *
0-
02
b110 6
#75010000000
1!
1%
1-
12
#75020000000
0!
0%
b111 *
0-
02
b111 6
#75030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#75040000000
0!
0%
b0 *
0-
02
b0 6
#75050000000
1!
1%
1-
12
#75060000000
0!
0%
b1 *
0-
02
b1 6
#75070000000
1!
1%
1-
12
#75080000000
0!
0%
b10 *
0-
02
b10 6
#75090000000
1!
1%
1-
12
#75100000000
0!
0%
b11 *
0-
02
b11 6
#75110000000
1!
1%
1-
12
15
#75120000000
0!
0%
b100 *
0-
02
b100 6
#75130000000
1!
1%
1-
12
#75140000000
0!
0%
b101 *
0-
02
b101 6
#75150000000
1!
1%
1-
12
#75160000000
0!
0%
b110 *
0-
02
b110 6
#75170000000
1!
1%
1-
12
#75180000000
0!
0%
b111 *
0-
02
b111 6
#75190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#75200000000
0!
0%
b0 *
0-
02
b0 6
#75210000000
1!
1%
1-
12
#75220000000
0!
0%
b1 *
0-
02
b1 6
#75230000000
1!
1%
1-
12
#75240000000
0!
0%
b10 *
0-
02
b10 6
#75250000000
1!
1%
1-
12
#75260000000
0!
0%
b11 *
0-
02
b11 6
#75270000000
1!
1%
1-
12
15
#75280000000
0!
0%
b100 *
0-
02
b100 6
#75290000000
1!
1%
1-
12
#75300000000
0!
0%
b101 *
0-
02
b101 6
#75310000000
1!
1%
1-
12
#75320000000
0!
0%
b110 *
0-
02
b110 6
#75330000000
1!
1%
1-
12
#75340000000
0!
0%
b111 *
0-
02
b111 6
#75350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#75360000000
0!
0%
b0 *
0-
02
b0 6
#75370000000
1!
1%
1-
12
#75380000000
0!
0%
b1 *
0-
02
b1 6
#75390000000
1!
1%
1-
12
#75400000000
0!
0%
b10 *
0-
02
b10 6
#75410000000
1!
1%
1-
12
#75420000000
0!
0%
b11 *
0-
02
b11 6
#75430000000
1!
1%
1-
12
15
#75440000000
0!
0%
b100 *
0-
02
b100 6
#75450000000
1!
1%
1-
12
#75460000000
0!
0%
b101 *
0-
02
b101 6
#75470000000
1!
1%
1-
12
#75480000000
0!
0%
b110 *
0-
02
b110 6
#75490000000
1!
1%
1-
12
#75500000000
0!
0%
b111 *
0-
02
b111 6
#75510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#75520000000
0!
0%
b0 *
0-
02
b0 6
#75530000000
1!
1%
1-
12
#75540000000
0!
0%
b1 *
0-
02
b1 6
#75550000000
1!
1%
1-
12
#75560000000
0!
0%
b10 *
0-
02
b10 6
#75570000000
1!
1%
1-
12
#75580000000
0!
0%
b11 *
0-
02
b11 6
#75590000000
1!
1%
1-
12
15
#75600000000
0!
0%
b100 *
0-
02
b100 6
#75610000000
1!
1%
1-
12
#75620000000
0!
0%
b101 *
0-
02
b101 6
#75630000000
1!
1%
1-
12
#75640000000
0!
0%
b110 *
0-
02
b110 6
#75650000000
1!
1%
1-
12
#75660000000
0!
0%
b111 *
0-
02
b111 6
#75670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#75680000000
0!
0%
b0 *
0-
02
b0 6
#75690000000
1!
1%
1-
12
#75700000000
0!
0%
b1 *
0-
02
b1 6
#75710000000
1!
1%
1-
12
#75720000000
0!
0%
b10 *
0-
02
b10 6
#75730000000
1!
1%
1-
12
#75740000000
0!
0%
b11 *
0-
02
b11 6
#75750000000
1!
1%
1-
12
15
#75760000000
0!
0%
b100 *
0-
02
b100 6
#75770000000
1!
1%
1-
12
#75780000000
0!
0%
b101 *
0-
02
b101 6
#75790000000
1!
1%
1-
12
#75800000000
0!
0%
b110 *
0-
02
b110 6
#75810000000
1!
1%
1-
12
#75820000000
0!
0%
b111 *
0-
02
b111 6
#75830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#75840000000
0!
0%
b0 *
0-
02
b0 6
#75850000000
1!
1%
1-
12
#75860000000
0!
0%
b1 *
0-
02
b1 6
#75870000000
1!
1%
1-
12
#75880000000
0!
0%
b10 *
0-
02
b10 6
#75890000000
1!
1%
1-
12
#75900000000
0!
0%
b11 *
0-
02
b11 6
#75910000000
1!
1%
1-
12
15
#75920000000
0!
0%
b100 *
0-
02
b100 6
#75930000000
1!
1%
1-
12
#75940000000
0!
0%
b101 *
0-
02
b101 6
#75950000000
1!
1%
1-
12
#75960000000
0!
0%
b110 *
0-
02
b110 6
#75970000000
1!
1%
1-
12
#75980000000
0!
0%
b111 *
0-
02
b111 6
#75990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#76000000000
0!
0%
b0 *
0-
02
b0 6
#76010000000
1!
1%
1-
12
#76020000000
0!
0%
b1 *
0-
02
b1 6
#76030000000
1!
1%
1-
12
#76040000000
0!
0%
b10 *
0-
02
b10 6
#76050000000
1!
1%
1-
12
#76060000000
0!
0%
b11 *
0-
02
b11 6
#76070000000
1!
1%
1-
12
15
#76080000000
0!
0%
b100 *
0-
02
b100 6
#76090000000
1!
1%
1-
12
#76100000000
0!
0%
b101 *
0-
02
b101 6
#76110000000
1!
1%
1-
12
#76120000000
0!
0%
b110 *
0-
02
b110 6
#76130000000
1!
1%
1-
12
#76140000000
0!
0%
b111 *
0-
02
b111 6
#76150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#76160000000
0!
0%
b0 *
0-
02
b0 6
#76170000000
1!
1%
1-
12
#76180000000
0!
0%
b1 *
0-
02
b1 6
#76190000000
1!
1%
1-
12
#76200000000
0!
0%
b10 *
0-
02
b10 6
#76210000000
1!
1%
1-
12
#76220000000
0!
0%
b11 *
0-
02
b11 6
#76230000000
1!
1%
1-
12
15
#76240000000
0!
0%
b100 *
0-
02
b100 6
#76250000000
1!
1%
1-
12
#76260000000
0!
0%
b101 *
0-
02
b101 6
#76270000000
1!
1%
1-
12
#76280000000
0!
0%
b110 *
0-
02
b110 6
#76290000000
1!
1%
1-
12
#76300000000
0!
0%
b111 *
0-
02
b111 6
#76310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#76320000000
0!
0%
b0 *
0-
02
b0 6
#76330000000
1!
1%
1-
12
#76340000000
0!
0%
b1 *
0-
02
b1 6
#76350000000
1!
1%
1-
12
#76360000000
0!
0%
b10 *
0-
02
b10 6
#76370000000
1!
1%
1-
12
#76380000000
0!
0%
b11 *
0-
02
b11 6
#76390000000
1!
1%
1-
12
15
#76400000000
0!
0%
b100 *
0-
02
b100 6
#76410000000
1!
1%
1-
12
#76420000000
0!
0%
b101 *
0-
02
b101 6
#76430000000
1!
1%
1-
12
#76440000000
0!
0%
b110 *
0-
02
b110 6
#76450000000
1!
1%
1-
12
#76460000000
0!
0%
b111 *
0-
02
b111 6
#76470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#76480000000
0!
0%
b0 *
0-
02
b0 6
#76490000000
1!
1%
1-
12
#76500000000
0!
0%
b1 *
0-
02
b1 6
#76510000000
1!
1%
1-
12
#76520000000
0!
0%
b10 *
0-
02
b10 6
#76530000000
1!
1%
1-
12
#76540000000
0!
0%
b11 *
0-
02
b11 6
#76550000000
1!
1%
1-
12
15
#76560000000
0!
0%
b100 *
0-
02
b100 6
#76570000000
1!
1%
1-
12
#76580000000
0!
0%
b101 *
0-
02
b101 6
#76590000000
1!
1%
1-
12
#76600000000
0!
0%
b110 *
0-
02
b110 6
#76610000000
1!
1%
1-
12
#76620000000
0!
0%
b111 *
0-
02
b111 6
#76630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#76640000000
0!
0%
b0 *
0-
02
b0 6
#76650000000
1!
1%
1-
12
#76660000000
0!
0%
b1 *
0-
02
b1 6
#76670000000
1!
1%
1-
12
#76680000000
0!
0%
b10 *
0-
02
b10 6
#76690000000
1!
1%
1-
12
#76700000000
0!
0%
b11 *
0-
02
b11 6
#76710000000
1!
1%
1-
12
15
#76720000000
0!
0%
b100 *
0-
02
b100 6
#76730000000
1!
1%
1-
12
#76740000000
0!
0%
b101 *
0-
02
b101 6
#76750000000
1!
1%
1-
12
#76760000000
0!
0%
b110 *
0-
02
b110 6
#76770000000
1!
1%
1-
12
#76780000000
0!
0%
b111 *
0-
02
b111 6
#76790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#76800000000
0!
0%
b0 *
0-
02
b0 6
#76810000000
1!
1%
1-
12
#76820000000
0!
0%
b1 *
0-
02
b1 6
#76830000000
1!
1%
1-
12
#76840000000
0!
0%
b10 *
0-
02
b10 6
#76850000000
1!
1%
1-
12
#76860000000
0!
0%
b11 *
0-
02
b11 6
#76870000000
1!
1%
1-
12
15
#76880000000
0!
0%
b100 *
0-
02
b100 6
#76890000000
1!
1%
1-
12
#76900000000
0!
0%
b101 *
0-
02
b101 6
#76910000000
1!
1%
1-
12
#76920000000
0!
0%
b110 *
0-
02
b110 6
#76930000000
1!
1%
1-
12
#76940000000
0!
0%
b111 *
0-
02
b111 6
#76950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#76960000000
0!
0%
b0 *
0-
02
b0 6
#76970000000
1!
1%
1-
12
#76980000000
0!
0%
b1 *
0-
02
b1 6
#76990000000
1!
1%
1-
12
#77000000000
0!
0%
b10 *
0-
02
b10 6
#77010000000
1!
1%
1-
12
#77020000000
0!
0%
b11 *
0-
02
b11 6
#77030000000
1!
1%
1-
12
15
#77040000000
0!
0%
b100 *
0-
02
b100 6
#77050000000
1!
1%
1-
12
#77060000000
0!
0%
b101 *
0-
02
b101 6
#77070000000
1!
1%
1-
12
#77080000000
0!
0%
b110 *
0-
02
b110 6
#77090000000
1!
1%
1-
12
#77100000000
0!
0%
b111 *
0-
02
b111 6
#77110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#77120000000
0!
0%
b0 *
0-
02
b0 6
#77130000000
1!
1%
1-
12
#77140000000
0!
0%
b1 *
0-
02
b1 6
#77150000000
1!
1%
1-
12
#77160000000
0!
0%
b10 *
0-
02
b10 6
#77170000000
1!
1%
1-
12
#77180000000
0!
0%
b11 *
0-
02
b11 6
#77190000000
1!
1%
1-
12
15
#77200000000
0!
0%
b100 *
0-
02
b100 6
#77210000000
1!
1%
1-
12
#77220000000
0!
0%
b101 *
0-
02
b101 6
#77230000000
1!
1%
1-
12
#77240000000
0!
0%
b110 *
0-
02
b110 6
#77250000000
1!
1%
1-
12
#77260000000
0!
0%
b111 *
0-
02
b111 6
#77270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#77280000000
0!
0%
b0 *
0-
02
b0 6
#77290000000
1!
1%
1-
12
#77300000000
0!
0%
b1 *
0-
02
b1 6
#77310000000
1!
1%
1-
12
#77320000000
0!
0%
b10 *
0-
02
b10 6
#77330000000
1!
1%
1-
12
#77340000000
0!
0%
b11 *
0-
02
b11 6
#77350000000
1!
1%
1-
12
15
#77360000000
0!
0%
b100 *
0-
02
b100 6
#77370000000
1!
1%
1-
12
#77380000000
0!
0%
b101 *
0-
02
b101 6
#77390000000
1!
1%
1-
12
#77400000000
0!
0%
b110 *
0-
02
b110 6
#77410000000
1!
1%
1-
12
#77420000000
0!
0%
b111 *
0-
02
b111 6
#77430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#77440000000
0!
0%
b0 *
0-
02
b0 6
#77450000000
1!
1%
1-
12
#77460000000
0!
0%
b1 *
0-
02
b1 6
#77470000000
1!
1%
1-
12
#77480000000
0!
0%
b10 *
0-
02
b10 6
#77490000000
1!
1%
1-
12
#77500000000
0!
0%
b11 *
0-
02
b11 6
#77510000000
1!
1%
1-
12
15
#77520000000
0!
0%
b100 *
0-
02
b100 6
#77530000000
1!
1%
1-
12
#77540000000
0!
0%
b101 *
0-
02
b101 6
#77550000000
1!
1%
1-
12
#77560000000
0!
0%
b110 *
0-
02
b110 6
#77570000000
1!
1%
1-
12
#77580000000
0!
0%
b111 *
0-
02
b111 6
#77590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#77600000000
0!
0%
b0 *
0-
02
b0 6
#77610000000
1!
1%
1-
12
#77620000000
0!
0%
b1 *
0-
02
b1 6
#77630000000
1!
1%
1-
12
#77640000000
0!
0%
b10 *
0-
02
b10 6
#77650000000
1!
1%
1-
12
#77660000000
0!
0%
b11 *
0-
02
b11 6
#77670000000
1!
1%
1-
12
15
#77680000000
0!
0%
b100 *
0-
02
b100 6
#77690000000
1!
1%
1-
12
#77700000000
0!
0%
b101 *
0-
02
b101 6
#77710000000
1!
1%
1-
12
#77720000000
0!
0%
b110 *
0-
02
b110 6
#77730000000
1!
1%
1-
12
#77740000000
0!
0%
b111 *
0-
02
b111 6
#77750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#77760000000
0!
0%
b0 *
0-
02
b0 6
#77770000000
1!
1%
1-
12
#77780000000
0!
0%
b1 *
0-
02
b1 6
#77790000000
1!
1%
1-
12
#77800000000
0!
0%
b10 *
0-
02
b10 6
#77810000000
1!
1%
1-
12
#77820000000
0!
0%
b11 *
0-
02
b11 6
#77830000000
1!
1%
1-
12
15
#77840000000
0!
0%
b100 *
0-
02
b100 6
#77850000000
1!
1%
1-
12
#77860000000
0!
0%
b101 *
0-
02
b101 6
#77870000000
1!
1%
1-
12
#77880000000
0!
0%
b110 *
0-
02
b110 6
#77890000000
1!
1%
1-
12
#77900000000
0!
0%
b111 *
0-
02
b111 6
#77910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#77920000000
0!
0%
b0 *
0-
02
b0 6
#77930000000
1!
1%
1-
12
#77940000000
0!
0%
b1 *
0-
02
b1 6
#77950000000
1!
1%
1-
12
#77960000000
0!
0%
b10 *
0-
02
b10 6
#77970000000
1!
1%
1-
12
#77980000000
0!
0%
b11 *
0-
02
b11 6
#77990000000
1!
1%
1-
12
15
#78000000000
0!
0%
b100 *
0-
02
b100 6
#78010000000
1!
1%
1-
12
#78020000000
0!
0%
b101 *
0-
02
b101 6
#78030000000
1!
1%
1-
12
#78040000000
0!
0%
b110 *
0-
02
b110 6
#78050000000
1!
1%
1-
12
#78060000000
0!
0%
b111 *
0-
02
b111 6
#78070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#78080000000
0!
0%
b0 *
0-
02
b0 6
#78090000000
1!
1%
1-
12
#78100000000
0!
0%
b1 *
0-
02
b1 6
#78110000000
1!
1%
1-
12
#78120000000
0!
0%
b10 *
0-
02
b10 6
#78130000000
1!
1%
1-
12
#78140000000
0!
0%
b11 *
0-
02
b11 6
#78150000000
1!
1%
1-
12
15
#78160000000
0!
0%
b100 *
0-
02
b100 6
#78170000000
1!
1%
1-
12
#78180000000
0!
0%
b101 *
0-
02
b101 6
#78190000000
1!
1%
1-
12
#78200000000
0!
0%
b110 *
0-
02
b110 6
#78210000000
1!
1%
1-
12
#78220000000
0!
0%
b111 *
0-
02
b111 6
#78230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#78240000000
0!
0%
b0 *
0-
02
b0 6
#78250000000
1!
1%
1-
12
#78260000000
0!
0%
b1 *
0-
02
b1 6
#78270000000
1!
1%
1-
12
#78280000000
0!
0%
b10 *
0-
02
b10 6
#78290000000
1!
1%
1-
12
#78300000000
0!
0%
b11 *
0-
02
b11 6
#78310000000
1!
1%
1-
12
15
#78320000000
0!
0%
b100 *
0-
02
b100 6
#78330000000
1!
1%
1-
12
#78340000000
0!
0%
b101 *
0-
02
b101 6
#78350000000
1!
1%
1-
12
#78360000000
0!
0%
b110 *
0-
02
b110 6
#78370000000
1!
1%
1-
12
#78380000000
0!
0%
b111 *
0-
02
b111 6
#78390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#78400000000
0!
0%
b0 *
0-
02
b0 6
#78410000000
1!
1%
1-
12
#78420000000
0!
0%
b1 *
0-
02
b1 6
#78430000000
1!
1%
1-
12
#78440000000
0!
0%
b10 *
0-
02
b10 6
#78450000000
1!
1%
1-
12
#78460000000
0!
0%
b11 *
0-
02
b11 6
#78470000000
1!
1%
1-
12
15
#78480000000
0!
0%
b100 *
0-
02
b100 6
#78490000000
1!
1%
1-
12
#78500000000
0!
0%
b101 *
0-
02
b101 6
#78510000000
1!
1%
1-
12
#78520000000
0!
0%
b110 *
0-
02
b110 6
#78530000000
1!
1%
1-
12
#78540000000
0!
0%
b111 *
0-
02
b111 6
#78550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#78560000000
0!
0%
b0 *
0-
02
b0 6
#78570000000
1!
1%
1-
12
#78580000000
0!
0%
b1 *
0-
02
b1 6
#78590000000
1!
1%
1-
12
#78600000000
0!
0%
b10 *
0-
02
b10 6
#78610000000
1!
1%
1-
12
#78620000000
0!
0%
b11 *
0-
02
b11 6
#78630000000
1!
1%
1-
12
15
#78640000000
0!
0%
b100 *
0-
02
b100 6
#78650000000
1!
1%
1-
12
#78660000000
0!
0%
b101 *
0-
02
b101 6
#78670000000
1!
1%
1-
12
#78680000000
0!
0%
b110 *
0-
02
b110 6
#78690000000
1!
1%
1-
12
#78700000000
0!
0%
b111 *
0-
02
b111 6
#78710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#78720000000
0!
0%
b0 *
0-
02
b0 6
#78730000000
1!
1%
1-
12
#78740000000
0!
0%
b1 *
0-
02
b1 6
#78750000000
1!
1%
1-
12
#78760000000
0!
0%
b10 *
0-
02
b10 6
#78770000000
1!
1%
1-
12
#78780000000
0!
0%
b11 *
0-
02
b11 6
#78790000000
1!
1%
1-
12
15
#78800000000
0!
0%
b100 *
0-
02
b100 6
#78810000000
1!
1%
1-
12
#78820000000
0!
0%
b101 *
0-
02
b101 6
#78830000000
1!
1%
1-
12
#78840000000
0!
0%
b110 *
0-
02
b110 6
#78850000000
1!
1%
1-
12
#78860000000
0!
0%
b111 *
0-
02
b111 6
#78870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#78880000000
0!
0%
b0 *
0-
02
b0 6
#78890000000
1!
1%
1-
12
#78900000000
0!
0%
b1 *
0-
02
b1 6
#78910000000
1!
1%
1-
12
#78920000000
0!
0%
b10 *
0-
02
b10 6
#78930000000
1!
1%
1-
12
#78940000000
0!
0%
b11 *
0-
02
b11 6
#78950000000
1!
1%
1-
12
15
#78960000000
0!
0%
b100 *
0-
02
b100 6
#78970000000
1!
1%
1-
12
#78980000000
0!
0%
b101 *
0-
02
b101 6
#78990000000
1!
1%
1-
12
#79000000000
0!
0%
b110 *
0-
02
b110 6
#79010000000
1!
1%
1-
12
#79020000000
0!
0%
b111 *
0-
02
b111 6
#79030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#79040000000
0!
0%
b0 *
0-
02
b0 6
#79050000000
1!
1%
1-
12
#79060000000
0!
0%
b1 *
0-
02
b1 6
#79070000000
1!
1%
1-
12
#79080000000
0!
0%
b10 *
0-
02
b10 6
#79090000000
1!
1%
1-
12
#79100000000
0!
0%
b11 *
0-
02
b11 6
#79110000000
1!
1%
1-
12
15
#79120000000
0!
0%
b100 *
0-
02
b100 6
#79130000000
1!
1%
1-
12
#79140000000
0!
0%
b101 *
0-
02
b101 6
#79150000000
1!
1%
1-
12
#79160000000
0!
0%
b110 *
0-
02
b110 6
#79170000000
1!
1%
1-
12
#79180000000
0!
0%
b111 *
0-
02
b111 6
#79190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#79200000000
0!
0%
b0 *
0-
02
b0 6
#79210000000
1!
1%
1-
12
#79220000000
0!
0%
b1 *
0-
02
b1 6
#79230000000
1!
1%
1-
12
#79240000000
0!
0%
b10 *
0-
02
b10 6
#79250000000
1!
1%
1-
12
#79260000000
0!
0%
b11 *
0-
02
b11 6
#79270000000
1!
1%
1-
12
15
#79280000000
0!
0%
b100 *
0-
02
b100 6
#79290000000
1!
1%
1-
12
#79300000000
0!
0%
b101 *
0-
02
b101 6
#79310000000
1!
1%
1-
12
#79320000000
0!
0%
b110 *
0-
02
b110 6
#79330000000
1!
1%
1-
12
#79340000000
0!
0%
b111 *
0-
02
b111 6
#79350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#79360000000
0!
0%
b0 *
0-
02
b0 6
#79370000000
1!
1%
1-
12
#79380000000
0!
0%
b1 *
0-
02
b1 6
#79390000000
1!
1%
1-
12
#79400000000
0!
0%
b10 *
0-
02
b10 6
#79410000000
1!
1%
1-
12
#79420000000
0!
0%
b11 *
0-
02
b11 6
#79430000000
1!
1%
1-
12
15
#79440000000
0!
0%
b100 *
0-
02
b100 6
#79450000000
1!
1%
1-
12
#79460000000
0!
0%
b101 *
0-
02
b101 6
#79470000000
1!
1%
1-
12
#79480000000
0!
0%
b110 *
0-
02
b110 6
#79490000000
1!
1%
1-
12
#79500000000
0!
0%
b111 *
0-
02
b111 6
#79510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#79520000000
0!
0%
b0 *
0-
02
b0 6
#79530000000
1!
1%
1-
12
#79540000000
0!
0%
b1 *
0-
02
b1 6
#79550000000
1!
1%
1-
12
#79560000000
0!
0%
b10 *
0-
02
b10 6
#79570000000
1!
1%
1-
12
#79580000000
0!
0%
b11 *
0-
02
b11 6
#79590000000
1!
1%
1-
12
15
#79600000000
0!
0%
b100 *
0-
02
b100 6
#79610000000
1!
1%
1-
12
#79620000000
0!
0%
b101 *
0-
02
b101 6
#79630000000
1!
1%
1-
12
#79640000000
0!
0%
b110 *
0-
02
b110 6
#79650000000
1!
1%
1-
12
#79660000000
0!
0%
b111 *
0-
02
b111 6
#79670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#79680000000
0!
0%
b0 *
0-
02
b0 6
#79690000000
1!
1%
1-
12
#79700000000
0!
0%
b1 *
0-
02
b1 6
#79710000000
1!
1%
1-
12
#79720000000
0!
0%
b10 *
0-
02
b10 6
#79730000000
1!
1%
1-
12
#79740000000
0!
0%
b11 *
0-
02
b11 6
#79750000000
1!
1%
1-
12
15
#79760000000
0!
0%
b100 *
0-
02
b100 6
#79770000000
1!
1%
1-
12
#79780000000
0!
0%
b101 *
0-
02
b101 6
#79790000000
1!
1%
1-
12
#79800000000
0!
0%
b110 *
0-
02
b110 6
#79810000000
1!
1%
1-
12
#79820000000
0!
0%
b111 *
0-
02
b111 6
#79830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#79840000000
0!
0%
b0 *
0-
02
b0 6
#79850000000
1!
1%
1-
12
#79860000000
0!
0%
b1 *
0-
02
b1 6
#79870000000
1!
1%
1-
12
#79880000000
0!
0%
b10 *
0-
02
b10 6
#79890000000
1!
1%
1-
12
#79900000000
0!
0%
b11 *
0-
02
b11 6
#79910000000
1!
1%
1-
12
15
#79920000000
0!
0%
b100 *
0-
02
b100 6
#79930000000
1!
1%
1-
12
#79940000000
0!
0%
b101 *
0-
02
b101 6
#79950000000
1!
1%
1-
12
#79960000000
0!
0%
b110 *
0-
02
b110 6
#79970000000
1!
1%
1-
12
#79980000000
0!
0%
b111 *
0-
02
b111 6
#79990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#80000000000
0!
0%
b0 *
0-
02
b0 6
#80010000000
1!
1%
1-
12
#80020000000
0!
0%
b1 *
0-
02
b1 6
#80030000000
1!
1%
1-
12
#80040000000
0!
0%
b10 *
0-
02
b10 6
#80050000000
1!
1%
1-
12
#80060000000
0!
0%
b11 *
0-
02
b11 6
#80070000000
1!
1%
1-
12
15
#80080000000
0!
0%
b100 *
0-
02
b100 6
#80090000000
1!
1%
1-
12
#80100000000
0!
0%
b101 *
0-
02
b101 6
#80110000000
1!
1%
1-
12
#80120000000
0!
0%
b110 *
0-
02
b110 6
#80130000000
1!
1%
1-
12
#80140000000
0!
0%
b111 *
0-
02
b111 6
#80150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#80160000000
0!
0%
b0 *
0-
02
b0 6
#80170000000
1!
1%
1-
12
#80180000000
0!
0%
b1 *
0-
02
b1 6
#80190000000
1!
1%
1-
12
#80200000000
0!
0%
b10 *
0-
02
b10 6
#80210000000
1!
1%
1-
12
#80220000000
0!
0%
b11 *
0-
02
b11 6
#80230000000
1!
1%
1-
12
15
#80240000000
0!
0%
b100 *
0-
02
b100 6
#80250000000
1!
1%
1-
12
#80260000000
0!
0%
b101 *
0-
02
b101 6
#80270000000
1!
1%
1-
12
#80280000000
0!
0%
b110 *
0-
02
b110 6
#80290000000
1!
1%
1-
12
#80300000000
0!
0%
b111 *
0-
02
b111 6
#80310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#80320000000
0!
0%
b0 *
0-
02
b0 6
#80330000000
1!
1%
1-
12
#80340000000
0!
0%
b1 *
0-
02
b1 6
#80350000000
1!
1%
1-
12
#80360000000
0!
0%
b10 *
0-
02
b10 6
#80370000000
1!
1%
1-
12
#80380000000
0!
0%
b11 *
0-
02
b11 6
#80390000000
1!
1%
1-
12
15
#80400000000
0!
0%
b100 *
0-
02
b100 6
#80410000000
1!
1%
1-
12
#80420000000
0!
0%
b101 *
0-
02
b101 6
#80430000000
1!
1%
1-
12
#80440000000
0!
0%
b110 *
0-
02
b110 6
#80450000000
1!
1%
1-
12
#80460000000
0!
0%
b111 *
0-
02
b111 6
#80470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#80480000000
0!
0%
b0 *
0-
02
b0 6
#80490000000
1!
1%
1-
12
#80500000000
0!
0%
b1 *
0-
02
b1 6
#80510000000
1!
1%
1-
12
#80520000000
0!
0%
b10 *
0-
02
b10 6
#80530000000
1!
1%
1-
12
#80540000000
0!
0%
b11 *
0-
02
b11 6
#80550000000
1!
1%
1-
12
15
#80560000000
0!
0%
b100 *
0-
02
b100 6
#80570000000
1!
1%
1-
12
#80580000000
0!
0%
b101 *
0-
02
b101 6
#80590000000
1!
1%
1-
12
#80600000000
0!
0%
b110 *
0-
02
b110 6
#80610000000
1!
1%
1-
12
#80620000000
0!
0%
b111 *
0-
02
b111 6
#80630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#80640000000
0!
0%
b0 *
0-
02
b0 6
#80650000000
1!
1%
1-
12
#80660000000
0!
0%
b1 *
0-
02
b1 6
#80670000000
1!
1%
1-
12
#80680000000
0!
0%
b10 *
0-
02
b10 6
#80690000000
1!
1%
1-
12
#80700000000
0!
0%
b11 *
0-
02
b11 6
#80710000000
1!
1%
1-
12
15
#80720000000
0!
0%
b100 *
0-
02
b100 6
#80730000000
1!
1%
1-
12
#80740000000
0!
0%
b101 *
0-
02
b101 6
#80750000000
1!
1%
1-
12
#80760000000
0!
0%
b110 *
0-
02
b110 6
#80770000000
1!
1%
1-
12
#80780000000
0!
0%
b111 *
0-
02
b111 6
#80790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#80800000000
0!
0%
b0 *
0-
02
b0 6
#80810000000
1!
1%
1-
12
#80820000000
0!
0%
b1 *
0-
02
b1 6
#80830000000
1!
1%
1-
12
#80840000000
0!
0%
b10 *
0-
02
b10 6
#80850000000
1!
1%
1-
12
#80860000000
0!
0%
b11 *
0-
02
b11 6
#80870000000
1!
1%
1-
12
15
#80880000000
0!
0%
b100 *
0-
02
b100 6
#80890000000
1!
1%
1-
12
#80900000000
0!
0%
b101 *
0-
02
b101 6
#80910000000
1!
1%
1-
12
#80920000000
0!
0%
b110 *
0-
02
b110 6
#80930000000
1!
1%
1-
12
#80940000000
0!
0%
b111 *
0-
02
b111 6
#80950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#80960000000
0!
0%
b0 *
0-
02
b0 6
#80970000000
1!
1%
1-
12
#80980000000
0!
0%
b1 *
0-
02
b1 6
#80990000000
1!
1%
1-
12
#81000000000
0!
0%
b10 *
0-
02
b10 6
#81010000000
1!
1%
1-
12
#81020000000
0!
0%
b11 *
0-
02
b11 6
#81030000000
1!
1%
1-
12
15
#81040000000
0!
0%
b100 *
0-
02
b100 6
#81050000000
1!
1%
1-
12
#81060000000
0!
0%
b101 *
0-
02
b101 6
#81070000000
1!
1%
1-
12
#81080000000
0!
0%
b110 *
0-
02
b110 6
#81090000000
1!
1%
1-
12
#81100000000
0!
0%
b111 *
0-
02
b111 6
#81110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#81120000000
0!
0%
b0 *
0-
02
b0 6
#81130000000
1!
1%
1-
12
#81140000000
0!
0%
b1 *
0-
02
b1 6
#81150000000
1!
1%
1-
12
#81160000000
0!
0%
b10 *
0-
02
b10 6
#81170000000
1!
1%
1-
12
#81180000000
0!
0%
b11 *
0-
02
b11 6
#81190000000
1!
1%
1-
12
15
#81200000000
0!
0%
b100 *
0-
02
b100 6
#81210000000
1!
1%
1-
12
#81220000000
0!
0%
b101 *
0-
02
b101 6
#81230000000
1!
1%
1-
12
#81240000000
0!
0%
b110 *
0-
02
b110 6
#81250000000
1!
1%
1-
12
#81260000000
0!
0%
b111 *
0-
02
b111 6
#81270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#81280000000
0!
0%
b0 *
0-
02
b0 6
#81290000000
1!
1%
1-
12
#81300000000
0!
0%
b1 *
0-
02
b1 6
#81310000000
1!
1%
1-
12
#81320000000
0!
0%
b10 *
0-
02
b10 6
#81330000000
1!
1%
1-
12
#81340000000
0!
0%
b11 *
0-
02
b11 6
#81350000000
1!
1%
1-
12
15
#81360000000
0!
0%
b100 *
0-
02
b100 6
#81370000000
1!
1%
1-
12
#81380000000
0!
0%
b101 *
0-
02
b101 6
#81390000000
1!
1%
1-
12
#81400000000
0!
0%
b110 *
0-
02
b110 6
#81410000000
1!
1%
1-
12
#81420000000
0!
0%
b111 *
0-
02
b111 6
#81430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#81440000000
0!
0%
b0 *
0-
02
b0 6
#81450000000
1!
1%
1-
12
#81460000000
0!
0%
b1 *
0-
02
b1 6
#81470000000
1!
1%
1-
12
#81480000000
0!
0%
b10 *
0-
02
b10 6
#81490000000
1!
1%
1-
12
#81500000000
0!
0%
b11 *
0-
02
b11 6
#81510000000
1!
1%
1-
12
15
#81520000000
0!
0%
b100 *
0-
02
b100 6
#81530000000
1!
1%
1-
12
#81540000000
0!
0%
b101 *
0-
02
b101 6
#81550000000
1!
1%
1-
12
#81560000000
0!
0%
b110 *
0-
02
b110 6
#81570000000
1!
1%
1-
12
#81580000000
0!
0%
b111 *
0-
02
b111 6
#81590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#81600000000
0!
0%
b0 *
0-
02
b0 6
#81610000000
1!
1%
1-
12
#81620000000
0!
0%
b1 *
0-
02
b1 6
#81630000000
1!
1%
1-
12
#81640000000
0!
0%
b10 *
0-
02
b10 6
#81650000000
1!
1%
1-
12
#81660000000
0!
0%
b11 *
0-
02
b11 6
#81670000000
1!
1%
1-
12
15
#81680000000
0!
0%
b100 *
0-
02
b100 6
#81690000000
1!
1%
1-
12
#81700000000
0!
0%
b101 *
0-
02
b101 6
#81710000000
1!
1%
1-
12
#81720000000
0!
0%
b110 *
0-
02
b110 6
#81730000000
1!
1%
1-
12
#81740000000
0!
0%
b111 *
0-
02
b111 6
#81750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#81760000000
0!
0%
b0 *
0-
02
b0 6
#81770000000
1!
1%
1-
12
#81780000000
0!
0%
b1 *
0-
02
b1 6
#81790000000
1!
1%
1-
12
#81800000000
0!
0%
b10 *
0-
02
b10 6
#81810000000
1!
1%
1-
12
#81820000000
0!
0%
b11 *
0-
02
b11 6
#81830000000
1!
1%
1-
12
15
#81840000000
0!
0%
b100 *
0-
02
b100 6
#81850000000
1!
1%
1-
12
#81860000000
0!
0%
b101 *
0-
02
b101 6
#81870000000
1!
1%
1-
12
#81880000000
0!
0%
b110 *
0-
02
b110 6
#81890000000
1!
1%
1-
12
#81900000000
0!
0%
b111 *
0-
02
b111 6
#81910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#81920000000
0!
0%
b0 *
0-
02
b0 6
#81930000000
1!
1%
1-
12
#81940000000
0!
0%
b1 *
0-
02
b1 6
#81950000000
1!
1%
1-
12
#81960000000
0!
0%
b10 *
0-
02
b10 6
#81970000000
1!
1%
1-
12
#81980000000
0!
0%
b11 *
0-
02
b11 6
#81990000000
1!
1%
1-
12
15
#82000000000
0!
0%
b100 *
0-
02
b100 6
#82010000000
1!
1%
1-
12
#82020000000
0!
0%
b101 *
0-
02
b101 6
#82030000000
1!
1%
1-
12
#82040000000
0!
0%
b110 *
0-
02
b110 6
#82050000000
1!
1%
1-
12
#82060000000
0!
0%
b111 *
0-
02
b111 6
#82070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#82080000000
0!
0%
b0 *
0-
02
b0 6
#82090000000
1!
1%
1-
12
#82100000000
0!
0%
b1 *
0-
02
b1 6
#82110000000
1!
1%
1-
12
#82120000000
0!
0%
b10 *
0-
02
b10 6
#82130000000
1!
1%
1-
12
#82140000000
0!
0%
b11 *
0-
02
b11 6
#82150000000
1!
1%
1-
12
15
#82160000000
0!
0%
b100 *
0-
02
b100 6
#82170000000
1!
1%
1-
12
#82180000000
0!
0%
b101 *
0-
02
b101 6
#82190000000
1!
1%
1-
12
#82200000000
0!
0%
b110 *
0-
02
b110 6
#82210000000
1!
1%
1-
12
#82220000000
0!
0%
b111 *
0-
02
b111 6
#82230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#82240000000
0!
0%
b0 *
0-
02
b0 6
#82250000000
1!
1%
1-
12
#82260000000
0!
0%
b1 *
0-
02
b1 6
#82270000000
1!
1%
1-
12
#82280000000
0!
0%
b10 *
0-
02
b10 6
#82290000000
1!
1%
1-
12
#82300000000
0!
0%
b11 *
0-
02
b11 6
#82310000000
1!
1%
1-
12
15
#82320000000
0!
0%
b100 *
0-
02
b100 6
#82330000000
1!
1%
1-
12
#82340000000
0!
0%
b101 *
0-
02
b101 6
#82350000000
1!
1%
1-
12
#82360000000
0!
0%
b110 *
0-
02
b110 6
#82370000000
1!
1%
1-
12
#82380000000
0!
0%
b111 *
0-
02
b111 6
#82390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#82400000000
0!
0%
b0 *
0-
02
b0 6
#82410000000
1!
1%
1-
12
#82420000000
0!
0%
b1 *
0-
02
b1 6
#82430000000
1!
1%
1-
12
#82440000000
0!
0%
b10 *
0-
02
b10 6
#82450000000
1!
1%
1-
12
#82460000000
0!
0%
b11 *
0-
02
b11 6
#82470000000
1!
1%
1-
12
15
#82480000000
0!
0%
b100 *
0-
02
b100 6
#82490000000
1!
1%
1-
12
#82500000000
0!
0%
b101 *
0-
02
b101 6
#82510000000
1!
1%
1-
12
#82520000000
0!
0%
b110 *
0-
02
b110 6
#82530000000
1!
1%
1-
12
#82540000000
0!
0%
b111 *
0-
02
b111 6
#82550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#82560000000
0!
0%
b0 *
0-
02
b0 6
#82570000000
1!
1%
1-
12
#82580000000
0!
0%
b1 *
0-
02
b1 6
#82590000000
1!
1%
1-
12
#82600000000
0!
0%
b10 *
0-
02
b10 6
#82610000000
1!
1%
1-
12
#82620000000
0!
0%
b11 *
0-
02
b11 6
#82630000000
1!
1%
1-
12
15
#82640000000
0!
0%
b100 *
0-
02
b100 6
#82650000000
1!
1%
1-
12
#82660000000
0!
0%
b101 *
0-
02
b101 6
#82670000000
1!
1%
1-
12
#82680000000
0!
0%
b110 *
0-
02
b110 6
#82690000000
1!
1%
1-
12
#82700000000
0!
0%
b111 *
0-
02
b111 6
#82710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#82720000000
0!
0%
b0 *
0-
02
b0 6
#82730000000
1!
1%
1-
12
#82740000000
0!
0%
b1 *
0-
02
b1 6
#82750000000
1!
1%
1-
12
#82760000000
0!
0%
b10 *
0-
02
b10 6
#82770000000
1!
1%
1-
12
#82780000000
0!
0%
b11 *
0-
02
b11 6
#82790000000
1!
1%
1-
12
15
#82800000000
0!
0%
b100 *
0-
02
b100 6
#82810000000
1!
1%
1-
12
#82820000000
0!
0%
b101 *
0-
02
b101 6
#82830000000
1!
1%
1-
12
#82840000000
0!
0%
b110 *
0-
02
b110 6
#82850000000
1!
1%
1-
12
#82860000000
0!
0%
b111 *
0-
02
b111 6
#82870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#82880000000
0!
0%
b0 *
0-
02
b0 6
#82890000000
1!
1%
1-
12
#82900000000
0!
0%
b1 *
0-
02
b1 6
#82910000000
1!
1%
1-
12
#82920000000
0!
0%
b10 *
0-
02
b10 6
#82930000000
1!
1%
1-
12
#82940000000
0!
0%
b11 *
0-
02
b11 6
#82950000000
1!
1%
1-
12
15
#82960000000
0!
0%
b100 *
0-
02
b100 6
#82970000000
1!
1%
1-
12
#82980000000
0!
0%
b101 *
0-
02
b101 6
#82990000000
1!
1%
1-
12
#83000000000
0!
0%
b110 *
0-
02
b110 6
#83010000000
1!
1%
1-
12
#83020000000
0!
0%
b111 *
0-
02
b111 6
#83030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#83040000000
0!
0%
b0 *
0-
02
b0 6
#83050000000
1!
1%
1-
12
#83060000000
0!
0%
b1 *
0-
02
b1 6
#83070000000
1!
1%
1-
12
#83080000000
0!
0%
b10 *
0-
02
b10 6
#83090000000
1!
1%
1-
12
#83100000000
0!
0%
b11 *
0-
02
b11 6
#83110000000
1!
1%
1-
12
15
#83120000000
0!
0%
b100 *
0-
02
b100 6
#83130000000
1!
1%
1-
12
#83140000000
0!
0%
b101 *
0-
02
b101 6
#83150000000
1!
1%
1-
12
#83160000000
0!
0%
b110 *
0-
02
b110 6
#83170000000
1!
1%
1-
12
#83180000000
0!
0%
b111 *
0-
02
b111 6
#83190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#83200000000
0!
0%
b0 *
0-
02
b0 6
#83210000000
1!
1%
1-
12
#83220000000
0!
0%
b1 *
0-
02
b1 6
#83230000000
1!
1%
1-
12
#83240000000
0!
0%
b10 *
0-
02
b10 6
#83250000000
1!
1%
1-
12
#83260000000
0!
0%
b11 *
0-
02
b11 6
#83270000000
1!
1%
1-
12
15
#83280000000
0!
0%
b100 *
0-
02
b100 6
#83290000000
1!
1%
1-
12
#83300000000
0!
0%
b101 *
0-
02
b101 6
#83310000000
1!
1%
1-
12
#83320000000
0!
0%
b110 *
0-
02
b110 6
#83330000000
1!
1%
1-
12
#83340000000
0!
0%
b111 *
0-
02
b111 6
#83350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#83360000000
0!
0%
b0 *
0-
02
b0 6
#83370000000
1!
1%
1-
12
#83380000000
0!
0%
b1 *
0-
02
b1 6
#83390000000
1!
1%
1-
12
#83400000000
0!
0%
b10 *
0-
02
b10 6
#83410000000
1!
1%
1-
12
#83420000000
0!
0%
b11 *
0-
02
b11 6
#83430000000
1!
1%
1-
12
15
#83440000000
0!
0%
b100 *
0-
02
b100 6
#83450000000
1!
1%
1-
12
#83460000000
0!
0%
b101 *
0-
02
b101 6
#83470000000
1!
1%
1-
12
#83480000000
0!
0%
b110 *
0-
02
b110 6
#83490000000
1!
1%
1-
12
#83500000000
0!
0%
b111 *
0-
02
b111 6
#83510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#83520000000
0!
0%
b0 *
0-
02
b0 6
#83530000000
1!
1%
1-
12
#83540000000
0!
0%
b1 *
0-
02
b1 6
#83550000000
1!
1%
1-
12
#83560000000
0!
0%
b10 *
0-
02
b10 6
#83570000000
1!
1%
1-
12
#83580000000
0!
0%
b11 *
0-
02
b11 6
#83590000000
1!
1%
1-
12
15
#83600000000
0!
0%
b100 *
0-
02
b100 6
#83610000000
1!
1%
1-
12
#83620000000
0!
0%
b101 *
0-
02
b101 6
#83630000000
1!
1%
1-
12
#83640000000
0!
0%
b110 *
0-
02
b110 6
#83650000000
1!
1%
1-
12
#83660000000
0!
0%
b111 *
0-
02
b111 6
#83670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#83680000000
0!
0%
b0 *
0-
02
b0 6
#83690000000
1!
1%
1-
12
#83700000000
0!
0%
b1 *
0-
02
b1 6
#83710000000
1!
1%
1-
12
#83720000000
0!
0%
b10 *
0-
02
b10 6
#83730000000
1!
1%
1-
12
#83740000000
0!
0%
b11 *
0-
02
b11 6
#83750000000
1!
1%
1-
12
15
#83760000000
0!
0%
b100 *
0-
02
b100 6
#83770000000
1!
1%
1-
12
#83780000000
0!
0%
b101 *
0-
02
b101 6
#83790000000
1!
1%
1-
12
#83800000000
0!
0%
b110 *
0-
02
b110 6
#83810000000
1!
1%
1-
12
#83820000000
0!
0%
b111 *
0-
02
b111 6
#83830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#83840000000
0!
0%
b0 *
0-
02
b0 6
#83850000000
1!
1%
1-
12
#83860000000
0!
0%
b1 *
0-
02
b1 6
#83870000000
1!
1%
1-
12
#83880000000
0!
0%
b10 *
0-
02
b10 6
#83890000000
1!
1%
1-
12
#83900000000
0!
0%
b11 *
0-
02
b11 6
#83910000000
1!
1%
1-
12
15
#83920000000
0!
0%
b100 *
0-
02
b100 6
#83930000000
1!
1%
1-
12
#83940000000
0!
0%
b101 *
0-
02
b101 6
#83950000000
1!
1%
1-
12
#83960000000
0!
0%
b110 *
0-
02
b110 6
#83970000000
1!
1%
1-
12
#83980000000
0!
0%
b111 *
0-
02
b111 6
#83990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#84000000000
0!
0%
b0 *
0-
02
b0 6
#84010000000
1!
1%
1-
12
#84020000000
0!
0%
b1 *
0-
02
b1 6
#84030000000
1!
1%
1-
12
#84040000000
0!
0%
b10 *
0-
02
b10 6
#84050000000
1!
1%
1-
12
#84060000000
0!
0%
b11 *
0-
02
b11 6
#84070000000
1!
1%
1-
12
15
#84080000000
0!
0%
b100 *
0-
02
b100 6
#84090000000
1!
1%
1-
12
#84100000000
0!
0%
b101 *
0-
02
b101 6
#84110000000
1!
1%
1-
12
#84120000000
0!
0%
b110 *
0-
02
b110 6
#84130000000
1!
1%
1-
12
#84140000000
0!
0%
b111 *
0-
02
b111 6
#84150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#84160000000
0!
0%
b0 *
0-
02
b0 6
#84170000000
1!
1%
1-
12
#84180000000
0!
0%
b1 *
0-
02
b1 6
#84190000000
1!
1%
1-
12
#84200000000
0!
0%
b10 *
0-
02
b10 6
#84210000000
1!
1%
1-
12
#84220000000
0!
0%
b11 *
0-
02
b11 6
#84230000000
1!
1%
1-
12
15
#84240000000
0!
0%
b100 *
0-
02
b100 6
#84250000000
1!
1%
1-
12
#84260000000
0!
0%
b101 *
0-
02
b101 6
#84270000000
1!
1%
1-
12
#84280000000
0!
0%
b110 *
0-
02
b110 6
#84290000000
1!
1%
1-
12
#84300000000
0!
0%
b111 *
0-
02
b111 6
#84310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#84320000000
0!
0%
b0 *
0-
02
b0 6
#84330000000
1!
1%
1-
12
#84340000000
0!
0%
b1 *
0-
02
b1 6
#84350000000
1!
1%
1-
12
#84360000000
0!
0%
b10 *
0-
02
b10 6
#84370000000
1!
1%
1-
12
#84380000000
0!
0%
b11 *
0-
02
b11 6
#84390000000
1!
1%
1-
12
15
#84400000000
0!
0%
b100 *
0-
02
b100 6
#84410000000
1!
1%
1-
12
#84420000000
0!
0%
b101 *
0-
02
b101 6
#84430000000
1!
1%
1-
12
#84440000000
0!
0%
b110 *
0-
02
b110 6
#84450000000
1!
1%
1-
12
#84460000000
0!
0%
b111 *
0-
02
b111 6
#84470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#84480000000
0!
0%
b0 *
0-
02
b0 6
#84490000000
1!
1%
1-
12
#84500000000
0!
0%
b1 *
0-
02
b1 6
#84510000000
1!
1%
1-
12
#84520000000
0!
0%
b10 *
0-
02
b10 6
#84530000000
1!
1%
1-
12
#84540000000
0!
0%
b11 *
0-
02
b11 6
#84550000000
1!
1%
1-
12
15
#84560000000
0!
0%
b100 *
0-
02
b100 6
#84570000000
1!
1%
1-
12
#84580000000
0!
0%
b101 *
0-
02
b101 6
#84590000000
1!
1%
1-
12
#84600000000
0!
0%
b110 *
0-
02
b110 6
#84610000000
1!
1%
1-
12
#84620000000
0!
0%
b111 *
0-
02
b111 6
#84630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#84640000000
0!
0%
b0 *
0-
02
b0 6
#84650000000
1!
1%
1-
12
#84660000000
0!
0%
b1 *
0-
02
b1 6
#84670000000
1!
1%
1-
12
#84680000000
0!
0%
b10 *
0-
02
b10 6
#84690000000
1!
1%
1-
12
#84700000000
0!
0%
b11 *
0-
02
b11 6
#84710000000
1!
1%
1-
12
15
#84720000000
0!
0%
b100 *
0-
02
b100 6
#84730000000
1!
1%
1-
12
#84740000000
0!
0%
b101 *
0-
02
b101 6
#84750000000
1!
1%
1-
12
#84760000000
0!
0%
b110 *
0-
02
b110 6
#84770000000
1!
1%
1-
12
#84780000000
0!
0%
b111 *
0-
02
b111 6
#84790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#84800000000
0!
0%
b0 *
0-
02
b0 6
#84810000000
1!
1%
1-
12
#84820000000
0!
0%
b1 *
0-
02
b1 6
#84830000000
1!
1%
1-
12
#84840000000
0!
0%
b10 *
0-
02
b10 6
#84850000000
1!
1%
1-
12
#84860000000
0!
0%
b11 *
0-
02
b11 6
#84870000000
1!
1%
1-
12
15
#84880000000
0!
0%
b100 *
0-
02
b100 6
#84890000000
1!
1%
1-
12
#84900000000
0!
0%
b101 *
0-
02
b101 6
#84910000000
1!
1%
1-
12
#84920000000
0!
0%
b110 *
0-
02
b110 6
#84930000000
1!
1%
1-
12
#84940000000
0!
0%
b111 *
0-
02
b111 6
#84950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#84960000000
0!
0%
b0 *
0-
02
b0 6
#84970000000
1!
1%
1-
12
#84980000000
0!
0%
b1 *
0-
02
b1 6
#84990000000
1!
1%
1-
12
#85000000000
0!
0%
b10 *
0-
02
b10 6
#85010000000
1!
1%
1-
12
#85020000000
0!
0%
b11 *
0-
02
b11 6
#85030000000
1!
1%
1-
12
15
#85040000000
0!
0%
b100 *
0-
02
b100 6
#85050000000
1!
1%
1-
12
#85060000000
0!
0%
b101 *
0-
02
b101 6
#85070000000
1!
1%
1-
12
#85080000000
0!
0%
b110 *
0-
02
b110 6
#85090000000
1!
1%
1-
12
#85100000000
0!
0%
b111 *
0-
02
b111 6
#85110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#85120000000
0!
0%
b0 *
0-
02
b0 6
#85130000000
1!
1%
1-
12
#85140000000
0!
0%
b1 *
0-
02
b1 6
#85150000000
1!
1%
1-
12
#85160000000
0!
0%
b10 *
0-
02
b10 6
#85170000000
1!
1%
1-
12
#85180000000
0!
0%
b11 *
0-
02
b11 6
#85190000000
1!
1%
1-
12
15
#85200000000
0!
0%
b100 *
0-
02
b100 6
#85210000000
1!
1%
1-
12
#85220000000
0!
0%
b101 *
0-
02
b101 6
#85230000000
1!
1%
1-
12
#85240000000
0!
0%
b110 *
0-
02
b110 6
#85250000000
1!
1%
1-
12
#85260000000
0!
0%
b111 *
0-
02
b111 6
#85270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#85280000000
0!
0%
b0 *
0-
02
b0 6
#85290000000
1!
1%
1-
12
#85300000000
0!
0%
b1 *
0-
02
b1 6
#85310000000
1!
1%
1-
12
#85320000000
0!
0%
b10 *
0-
02
b10 6
#85330000000
1!
1%
1-
12
#85340000000
0!
0%
b11 *
0-
02
b11 6
#85350000000
1!
1%
1-
12
15
#85360000000
0!
0%
b100 *
0-
02
b100 6
#85370000000
1!
1%
1-
12
#85380000000
0!
0%
b101 *
0-
02
b101 6
#85390000000
1!
1%
1-
12
#85400000000
0!
0%
b110 *
0-
02
b110 6
#85410000000
1!
1%
1-
12
#85420000000
0!
0%
b111 *
0-
02
b111 6
#85430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#85440000000
0!
0%
b0 *
0-
02
b0 6
#85450000000
1!
1%
1-
12
#85460000000
0!
0%
b1 *
0-
02
b1 6
#85470000000
1!
1%
1-
12
#85480000000
0!
0%
b10 *
0-
02
b10 6
#85490000000
1!
1%
1-
12
#85500000000
0!
0%
b11 *
0-
02
b11 6
#85510000000
1!
1%
1-
12
15
#85520000000
0!
0%
b100 *
0-
02
b100 6
#85530000000
1!
1%
1-
12
#85540000000
0!
0%
b101 *
0-
02
b101 6
#85550000000
1!
1%
1-
12
#85560000000
0!
0%
b110 *
0-
02
b110 6
#85570000000
1!
1%
1-
12
#85580000000
0!
0%
b111 *
0-
02
b111 6
#85590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#85600000000
0!
0%
b0 *
0-
02
b0 6
#85610000000
1!
1%
1-
12
#85620000000
0!
0%
b1 *
0-
02
b1 6
#85630000000
1!
1%
1-
12
#85640000000
0!
0%
b10 *
0-
02
b10 6
#85650000000
1!
1%
1-
12
#85660000000
0!
0%
b11 *
0-
02
b11 6
#85670000000
1!
1%
1-
12
15
#85680000000
0!
0%
b100 *
0-
02
b100 6
#85690000000
1!
1%
1-
12
#85700000000
0!
0%
b101 *
0-
02
b101 6
#85710000000
1!
1%
1-
12
#85720000000
0!
0%
b110 *
0-
02
b110 6
#85730000000
1!
1%
1-
12
#85740000000
0!
0%
b111 *
0-
02
b111 6
#85750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#85760000000
0!
0%
b0 *
0-
02
b0 6
#85770000000
1!
1%
1-
12
#85780000000
0!
0%
b1 *
0-
02
b1 6
#85790000000
1!
1%
1-
12
#85800000000
0!
0%
b10 *
0-
02
b10 6
#85810000000
1!
1%
1-
12
#85820000000
0!
0%
b11 *
0-
02
b11 6
#85830000000
1!
1%
1-
12
15
#85840000000
0!
0%
b100 *
0-
02
b100 6
#85850000000
1!
1%
1-
12
#85860000000
0!
0%
b101 *
0-
02
b101 6
#85870000000
1!
1%
1-
12
#85880000000
0!
0%
b110 *
0-
02
b110 6
#85890000000
1!
1%
1-
12
#85900000000
0!
0%
b111 *
0-
02
b111 6
#85910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#85920000000
0!
0%
b0 *
0-
02
b0 6
#85930000000
1!
1%
1-
12
#85940000000
0!
0%
b1 *
0-
02
b1 6
#85950000000
1!
1%
1-
12
#85960000000
0!
0%
b10 *
0-
02
b10 6
#85970000000
1!
1%
1-
12
#85980000000
0!
0%
b11 *
0-
02
b11 6
#85990000000
1!
1%
1-
12
15
#86000000000
0!
0%
b100 *
0-
02
b100 6
#86010000000
1!
1%
1-
12
#86020000000
0!
0%
b101 *
0-
02
b101 6
#86030000000
1!
1%
1-
12
#86040000000
0!
0%
b110 *
0-
02
b110 6
#86050000000
1!
1%
1-
12
#86060000000
0!
0%
b111 *
0-
02
b111 6
#86070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#86080000000
0!
0%
b0 *
0-
02
b0 6
#86090000000
1!
1%
1-
12
#86100000000
0!
0%
b1 *
0-
02
b1 6
#86110000000
1!
1%
1-
12
#86120000000
0!
0%
b10 *
0-
02
b10 6
#86130000000
1!
1%
1-
12
#86140000000
0!
0%
b11 *
0-
02
b11 6
#86150000000
1!
1%
1-
12
15
#86160000000
0!
0%
b100 *
0-
02
b100 6
#86170000000
1!
1%
1-
12
#86180000000
0!
0%
b101 *
0-
02
b101 6
#86190000000
1!
1%
1-
12
#86200000000
0!
0%
b110 *
0-
02
b110 6
#86210000000
1!
1%
1-
12
#86220000000
0!
0%
b111 *
0-
02
b111 6
#86230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#86240000000
0!
0%
b0 *
0-
02
b0 6
#86250000000
1!
1%
1-
12
#86260000000
0!
0%
b1 *
0-
02
b1 6
#86270000000
1!
1%
1-
12
#86280000000
0!
0%
b10 *
0-
02
b10 6
#86290000000
1!
1%
1-
12
#86300000000
0!
0%
b11 *
0-
02
b11 6
#86310000000
1!
1%
1-
12
15
#86320000000
0!
0%
b100 *
0-
02
b100 6
#86330000000
1!
1%
1-
12
#86340000000
0!
0%
b101 *
0-
02
b101 6
#86350000000
1!
1%
1-
12
#86360000000
0!
0%
b110 *
0-
02
b110 6
#86370000000
1!
1%
1-
12
#86380000000
0!
0%
b111 *
0-
02
b111 6
#86390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#86400000000
0!
0%
b0 *
0-
02
b0 6
#86410000000
1!
1%
1-
12
#86420000000
0!
0%
b1 *
0-
02
b1 6
#86430000000
1!
1%
1-
12
#86440000000
0!
0%
b10 *
0-
02
b10 6
#86450000000
1!
1%
1-
12
#86460000000
0!
0%
b11 *
0-
02
b11 6
#86470000000
1!
1%
1-
12
15
#86480000000
0!
0%
b100 *
0-
02
b100 6
#86490000000
1!
1%
1-
12
#86500000000
0!
0%
b101 *
0-
02
b101 6
#86510000000
1!
1%
1-
12
#86520000000
0!
0%
b110 *
0-
02
b110 6
#86530000000
1!
1%
1-
12
#86540000000
0!
0%
b111 *
0-
02
b111 6
#86550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#86560000000
0!
0%
b0 *
0-
02
b0 6
#86570000000
1!
1%
1-
12
#86580000000
0!
0%
b1 *
0-
02
b1 6
#86590000000
1!
1%
1-
12
#86600000000
0!
0%
b10 *
0-
02
b10 6
#86610000000
1!
1%
1-
12
#86620000000
0!
0%
b11 *
0-
02
b11 6
#86630000000
1!
1%
1-
12
15
#86640000000
0!
0%
b100 *
0-
02
b100 6
#86650000000
1!
1%
1-
12
#86660000000
0!
0%
b101 *
0-
02
b101 6
#86670000000
1!
1%
1-
12
#86680000000
0!
0%
b110 *
0-
02
b110 6
#86690000000
1!
1%
1-
12
#86700000000
0!
0%
b111 *
0-
02
b111 6
#86710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#86720000000
0!
0%
b0 *
0-
02
b0 6
#86730000000
1!
1%
1-
12
#86740000000
0!
0%
b1 *
0-
02
b1 6
#86750000000
1!
1%
1-
12
#86760000000
0!
0%
b10 *
0-
02
b10 6
#86770000000
1!
1%
1-
12
#86780000000
0!
0%
b11 *
0-
02
b11 6
#86790000000
1!
1%
1-
12
15
#86800000000
0!
0%
b100 *
0-
02
b100 6
#86810000000
1!
1%
1-
12
#86820000000
0!
0%
b101 *
0-
02
b101 6
#86830000000
1!
1%
1-
12
#86840000000
0!
0%
b110 *
0-
02
b110 6
#86850000000
1!
1%
1-
12
#86860000000
0!
0%
b111 *
0-
02
b111 6
#86870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#86880000000
0!
0%
b0 *
0-
02
b0 6
#86890000000
1!
1%
1-
12
#86900000000
0!
0%
b1 *
0-
02
b1 6
#86910000000
1!
1%
1-
12
#86920000000
0!
0%
b10 *
0-
02
b10 6
#86930000000
1!
1%
1-
12
#86940000000
0!
0%
b11 *
0-
02
b11 6
#86950000000
1!
1%
1-
12
15
#86960000000
0!
0%
b100 *
0-
02
b100 6
#86970000000
1!
1%
1-
12
#86980000000
0!
0%
b101 *
0-
02
b101 6
#86990000000
1!
1%
1-
12
#87000000000
0!
0%
b110 *
0-
02
b110 6
#87010000000
1!
1%
1-
12
#87020000000
0!
0%
b111 *
0-
02
b111 6
#87030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#87040000000
0!
0%
b0 *
0-
02
b0 6
#87050000000
1!
1%
1-
12
#87060000000
0!
0%
b1 *
0-
02
b1 6
#87070000000
1!
1%
1-
12
#87080000000
0!
0%
b10 *
0-
02
b10 6
#87090000000
1!
1%
1-
12
#87100000000
0!
0%
b11 *
0-
02
b11 6
#87110000000
1!
1%
1-
12
15
#87120000000
0!
0%
b100 *
0-
02
b100 6
#87130000000
1!
1%
1-
12
#87140000000
0!
0%
b101 *
0-
02
b101 6
#87150000000
1!
1%
1-
12
#87160000000
0!
0%
b110 *
0-
02
b110 6
#87170000000
1!
1%
1-
12
#87180000000
0!
0%
b111 *
0-
02
b111 6
#87190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#87200000000
0!
0%
b0 *
0-
02
b0 6
#87210000000
1!
1%
1-
12
#87220000000
0!
0%
b1 *
0-
02
b1 6
#87230000000
1!
1%
1-
12
#87240000000
0!
0%
b10 *
0-
02
b10 6
#87250000000
1!
1%
1-
12
#87260000000
0!
0%
b11 *
0-
02
b11 6
#87270000000
1!
1%
1-
12
15
#87280000000
0!
0%
b100 *
0-
02
b100 6
#87290000000
1!
1%
1-
12
#87300000000
0!
0%
b101 *
0-
02
b101 6
#87310000000
1!
1%
1-
12
#87320000000
0!
0%
b110 *
0-
02
b110 6
#87330000000
1!
1%
1-
12
#87340000000
0!
0%
b111 *
0-
02
b111 6
#87350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#87360000000
0!
0%
b0 *
0-
02
b0 6
#87370000000
1!
1%
1-
12
#87380000000
0!
0%
b1 *
0-
02
b1 6
#87390000000
1!
1%
1-
12
#87400000000
0!
0%
b10 *
0-
02
b10 6
#87410000000
1!
1%
1-
12
#87420000000
0!
0%
b11 *
0-
02
b11 6
#87430000000
1!
1%
1-
12
15
#87440000000
0!
0%
b100 *
0-
02
b100 6
#87450000000
1!
1%
1-
12
#87460000000
0!
0%
b101 *
0-
02
b101 6
#87470000000
1!
1%
1-
12
#87480000000
0!
0%
b110 *
0-
02
b110 6
#87490000000
1!
1%
1-
12
#87500000000
0!
0%
b111 *
0-
02
b111 6
#87510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#87520000000
0!
0%
b0 *
0-
02
b0 6
#87530000000
1!
1%
1-
12
#87540000000
0!
0%
b1 *
0-
02
b1 6
#87550000000
1!
1%
1-
12
#87560000000
0!
0%
b10 *
0-
02
b10 6
#87570000000
1!
1%
1-
12
#87580000000
0!
0%
b11 *
0-
02
b11 6
#87590000000
1!
1%
1-
12
15
#87600000000
0!
0%
b100 *
0-
02
b100 6
#87610000000
1!
1%
1-
12
#87620000000
0!
0%
b101 *
0-
02
b101 6
#87630000000
1!
1%
1-
12
#87640000000
0!
0%
b110 *
0-
02
b110 6
#87650000000
1!
1%
1-
12
#87660000000
0!
0%
b111 *
0-
02
b111 6
#87670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#87680000000
0!
0%
b0 *
0-
02
b0 6
#87690000000
1!
1%
1-
12
#87700000000
0!
0%
b1 *
0-
02
b1 6
#87710000000
1!
1%
1-
12
#87720000000
0!
0%
b10 *
0-
02
b10 6
#87730000000
1!
1%
1-
12
#87740000000
0!
0%
b11 *
0-
02
b11 6
#87750000000
1!
1%
1-
12
15
#87760000000
0!
0%
b100 *
0-
02
b100 6
#87770000000
1!
1%
1-
12
#87780000000
0!
0%
b101 *
0-
02
b101 6
#87790000000
1!
1%
1-
12
#87800000000
0!
0%
b110 *
0-
02
b110 6
#87810000000
1!
1%
1-
12
#87820000000
0!
0%
b111 *
0-
02
b111 6
#87830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#87840000000
0!
0%
b0 *
0-
02
b0 6
#87850000000
1!
1%
1-
12
#87860000000
0!
0%
b1 *
0-
02
b1 6
#87870000000
1!
1%
1-
12
#87880000000
0!
0%
b10 *
0-
02
b10 6
#87890000000
1!
1%
1-
12
#87900000000
0!
0%
b11 *
0-
02
b11 6
#87910000000
1!
1%
1-
12
15
#87920000000
0!
0%
b100 *
0-
02
b100 6
#87930000000
1!
1%
1-
12
#87940000000
0!
0%
b101 *
0-
02
b101 6
#87950000000
1!
1%
1-
12
#87960000000
0!
0%
b110 *
0-
02
b110 6
#87970000000
1!
1%
1-
12
#87980000000
0!
0%
b111 *
0-
02
b111 6
#87990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#88000000000
0!
0%
b0 *
0-
02
b0 6
#88010000000
1!
1%
1-
12
#88020000000
0!
0%
b1 *
0-
02
b1 6
#88030000000
1!
1%
1-
12
#88040000000
0!
0%
b10 *
0-
02
b10 6
#88050000000
1!
1%
1-
12
#88060000000
0!
0%
b11 *
0-
02
b11 6
#88070000000
1!
1%
1-
12
15
#88080000000
0!
0%
b100 *
0-
02
b100 6
#88090000000
1!
1%
1-
12
#88100000000
0!
0%
b101 *
0-
02
b101 6
#88110000000
1!
1%
1-
12
#88120000000
0!
0%
b110 *
0-
02
b110 6
#88130000000
1!
1%
1-
12
#88140000000
0!
0%
b111 *
0-
02
b111 6
#88150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#88160000000
0!
0%
b0 *
0-
02
b0 6
#88170000000
1!
1%
1-
12
#88180000000
0!
0%
b1 *
0-
02
b1 6
#88190000000
1!
1%
1-
12
#88200000000
0!
0%
b10 *
0-
02
b10 6
#88210000000
1!
1%
1-
12
#88220000000
0!
0%
b11 *
0-
02
b11 6
#88230000000
1!
1%
1-
12
15
#88240000000
0!
0%
b100 *
0-
02
b100 6
#88250000000
1!
1%
1-
12
#88260000000
0!
0%
b101 *
0-
02
b101 6
#88270000000
1!
1%
1-
12
#88280000000
0!
0%
b110 *
0-
02
b110 6
#88290000000
1!
1%
1-
12
#88300000000
0!
0%
b111 *
0-
02
b111 6
#88310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#88320000000
0!
0%
b0 *
0-
02
b0 6
#88330000000
1!
1%
1-
12
#88340000000
0!
0%
b1 *
0-
02
b1 6
#88350000000
1!
1%
1-
12
#88360000000
0!
0%
b10 *
0-
02
b10 6
#88370000000
1!
1%
1-
12
#88380000000
0!
0%
b11 *
0-
02
b11 6
#88390000000
1!
1%
1-
12
15
#88400000000
0!
0%
b100 *
0-
02
b100 6
#88410000000
1!
1%
1-
12
#88420000000
0!
0%
b101 *
0-
02
b101 6
#88430000000
1!
1%
1-
12
#88440000000
0!
0%
b110 *
0-
02
b110 6
#88450000000
1!
1%
1-
12
#88460000000
0!
0%
b111 *
0-
02
b111 6
#88470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#88480000000
0!
0%
b0 *
0-
02
b0 6
#88490000000
1!
1%
1-
12
#88500000000
0!
0%
b1 *
0-
02
b1 6
#88510000000
1!
1%
1-
12
#88520000000
0!
0%
b10 *
0-
02
b10 6
#88530000000
1!
1%
1-
12
#88540000000
0!
0%
b11 *
0-
02
b11 6
#88550000000
1!
1%
1-
12
15
#88560000000
0!
0%
b100 *
0-
02
b100 6
#88570000000
1!
1%
1-
12
#88580000000
0!
0%
b101 *
0-
02
b101 6
#88590000000
1!
1%
1-
12
#88600000000
0!
0%
b110 *
0-
02
b110 6
#88610000000
1!
1%
1-
12
#88620000000
0!
0%
b111 *
0-
02
b111 6
#88630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#88640000000
0!
0%
b0 *
0-
02
b0 6
#88650000000
1!
1%
1-
12
#88660000000
0!
0%
b1 *
0-
02
b1 6
#88670000000
1!
1%
1-
12
#88680000000
0!
0%
b10 *
0-
02
b10 6
#88690000000
1!
1%
1-
12
#88700000000
0!
0%
b11 *
0-
02
b11 6
#88710000000
1!
1%
1-
12
15
#88720000000
0!
0%
b100 *
0-
02
b100 6
#88730000000
1!
1%
1-
12
#88740000000
0!
0%
b101 *
0-
02
b101 6
#88750000000
1!
1%
1-
12
#88760000000
0!
0%
b110 *
0-
02
b110 6
#88770000000
1!
1%
1-
12
#88780000000
0!
0%
b111 *
0-
02
b111 6
#88790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#88800000000
0!
0%
b0 *
0-
02
b0 6
#88810000000
1!
1%
1-
12
#88820000000
0!
0%
b1 *
0-
02
b1 6
#88830000000
1!
1%
1-
12
#88840000000
0!
0%
b10 *
0-
02
b10 6
#88850000000
1!
1%
1-
12
#88860000000
0!
0%
b11 *
0-
02
b11 6
#88870000000
1!
1%
1-
12
15
#88880000000
0!
0%
b100 *
0-
02
b100 6
#88890000000
1!
1%
1-
12
#88900000000
0!
0%
b101 *
0-
02
b101 6
#88910000000
1!
1%
1-
12
#88920000000
0!
0%
b110 *
0-
02
b110 6
#88930000000
1!
1%
1-
12
#88940000000
0!
0%
b111 *
0-
02
b111 6
#88950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#88960000000
0!
0%
b0 *
0-
02
b0 6
#88970000000
1!
1%
1-
12
#88980000000
0!
0%
b1 *
0-
02
b1 6
#88990000000
1!
1%
1-
12
#89000000000
0!
0%
b10 *
0-
02
b10 6
#89010000000
1!
1%
1-
12
#89020000000
0!
0%
b11 *
0-
02
b11 6
#89030000000
1!
1%
1-
12
15
#89040000000
0!
0%
b100 *
0-
02
b100 6
#89050000000
1!
1%
1-
12
#89060000000
0!
0%
b101 *
0-
02
b101 6
#89070000000
1!
1%
1-
12
#89080000000
0!
0%
b110 *
0-
02
b110 6
#89090000000
1!
1%
1-
12
#89100000000
0!
0%
b111 *
0-
02
b111 6
#89110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#89120000000
0!
0%
b0 *
0-
02
b0 6
#89130000000
1!
1%
1-
12
#89140000000
0!
0%
b1 *
0-
02
b1 6
#89150000000
1!
1%
1-
12
#89160000000
0!
0%
b10 *
0-
02
b10 6
#89170000000
1!
1%
1-
12
#89180000000
0!
0%
b11 *
0-
02
b11 6
#89190000000
1!
1%
1-
12
15
#89200000000
0!
0%
b100 *
0-
02
b100 6
#89210000000
1!
1%
1-
12
#89220000000
0!
0%
b101 *
0-
02
b101 6
#89230000000
1!
1%
1-
12
#89240000000
0!
0%
b110 *
0-
02
b110 6
#89250000000
1!
1%
1-
12
#89260000000
0!
0%
b111 *
0-
02
b111 6
#89270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#89280000000
0!
0%
b0 *
0-
02
b0 6
#89290000000
1!
1%
1-
12
#89300000000
0!
0%
b1 *
0-
02
b1 6
#89310000000
1!
1%
1-
12
#89320000000
0!
0%
b10 *
0-
02
b10 6
#89330000000
1!
1%
1-
12
#89340000000
0!
0%
b11 *
0-
02
b11 6
#89350000000
1!
1%
1-
12
15
#89360000000
0!
0%
b100 *
0-
02
b100 6
#89370000000
1!
1%
1-
12
#89380000000
0!
0%
b101 *
0-
02
b101 6
#89390000000
1!
1%
1-
12
#89400000000
0!
0%
b110 *
0-
02
b110 6
#89410000000
1!
1%
1-
12
#89420000000
0!
0%
b111 *
0-
02
b111 6
#89430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#89440000000
0!
0%
b0 *
0-
02
b0 6
#89450000000
1!
1%
1-
12
#89460000000
0!
0%
b1 *
0-
02
b1 6
#89470000000
1!
1%
1-
12
#89480000000
0!
0%
b10 *
0-
02
b10 6
#89490000000
1!
1%
1-
12
#89500000000
0!
0%
b11 *
0-
02
b11 6
#89510000000
1!
1%
1-
12
15
#89520000000
0!
0%
b100 *
0-
02
b100 6
#89530000000
1!
1%
1-
12
#89540000000
0!
0%
b101 *
0-
02
b101 6
#89550000000
1!
1%
1-
12
#89560000000
0!
0%
b110 *
0-
02
b110 6
#89570000000
1!
1%
1-
12
#89580000000
0!
0%
b111 *
0-
02
b111 6
#89590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#89600000000
0!
0%
b0 *
0-
02
b0 6
#89610000000
1!
1%
1-
12
#89620000000
0!
0%
b1 *
0-
02
b1 6
#89630000000
1!
1%
1-
12
#89640000000
0!
0%
b10 *
0-
02
b10 6
#89650000000
1!
1%
1-
12
#89660000000
0!
0%
b11 *
0-
02
b11 6
#89670000000
1!
1%
1-
12
15
#89680000000
0!
0%
b100 *
0-
02
b100 6
#89690000000
1!
1%
1-
12
#89700000000
0!
0%
b101 *
0-
02
b101 6
#89710000000
1!
1%
1-
12
#89720000000
0!
0%
b110 *
0-
02
b110 6
#89730000000
1!
1%
1-
12
#89740000000
0!
0%
b111 *
0-
02
b111 6
#89750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#89760000000
0!
0%
b0 *
0-
02
b0 6
#89770000000
1!
1%
1-
12
#89780000000
0!
0%
b1 *
0-
02
b1 6
#89790000000
1!
1%
1-
12
#89800000000
0!
0%
b10 *
0-
02
b10 6
#89810000000
1!
1%
1-
12
#89820000000
0!
0%
b11 *
0-
02
b11 6
#89830000000
1!
1%
1-
12
15
#89840000000
0!
0%
b100 *
0-
02
b100 6
#89850000000
1!
1%
1-
12
#89860000000
0!
0%
b101 *
0-
02
b101 6
#89870000000
1!
1%
1-
12
#89880000000
0!
0%
b110 *
0-
02
b110 6
#89890000000
1!
1%
1-
12
#89900000000
0!
0%
b111 *
0-
02
b111 6
#89910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#89920000000
0!
0%
b0 *
0-
02
b0 6
#89930000000
1!
1%
1-
12
#89940000000
0!
0%
b1 *
0-
02
b1 6
#89950000000
1!
1%
1-
12
#89960000000
0!
0%
b10 *
0-
02
b10 6
#89970000000
1!
1%
1-
12
#89980000000
0!
0%
b11 *
0-
02
b11 6
#89990000000
1!
1%
1-
12
15
#90000000000
0!
0%
b100 *
0-
02
b100 6
#90010000000
1!
1%
1-
12
#90020000000
0!
0%
b101 *
0-
02
b101 6
#90030000000
1!
1%
1-
12
#90040000000
0!
0%
b110 *
0-
02
b110 6
#90050000000
1!
1%
1-
12
#90060000000
0!
0%
b111 *
0-
02
b111 6
#90070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#90080000000
0!
0%
b0 *
0-
02
b0 6
#90090000000
1!
1%
1-
12
#90100000000
0!
0%
b1 *
0-
02
b1 6
#90110000000
1!
1%
1-
12
#90120000000
0!
0%
b10 *
0-
02
b10 6
#90130000000
1!
1%
1-
12
#90140000000
0!
0%
b11 *
0-
02
b11 6
#90150000000
1!
1%
1-
12
15
#90160000000
0!
0%
b100 *
0-
02
b100 6
#90170000000
1!
1%
1-
12
#90180000000
0!
0%
b101 *
0-
02
b101 6
#90190000000
1!
1%
1-
12
#90200000000
0!
0%
b110 *
0-
02
b110 6
#90210000000
1!
1%
1-
12
#90220000000
0!
0%
b111 *
0-
02
b111 6
#90230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#90240000000
0!
0%
b0 *
0-
02
b0 6
#90250000000
1!
1%
1-
12
#90260000000
0!
0%
b1 *
0-
02
b1 6
#90270000000
1!
1%
1-
12
#90280000000
0!
0%
b10 *
0-
02
b10 6
#90290000000
1!
1%
1-
12
#90300000000
0!
0%
b11 *
0-
02
b11 6
#90310000000
1!
1%
1-
12
15
#90320000000
0!
0%
b100 *
0-
02
b100 6
#90330000000
1!
1%
1-
12
#90340000000
0!
0%
b101 *
0-
02
b101 6
#90350000000
1!
1%
1-
12
#90360000000
0!
0%
b110 *
0-
02
b110 6
#90370000000
1!
1%
1-
12
#90380000000
0!
0%
b111 *
0-
02
b111 6
#90390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#90400000000
0!
0%
b0 *
0-
02
b0 6
#90410000000
1!
1%
1-
12
#90420000000
0!
0%
b1 *
0-
02
b1 6
#90430000000
1!
1%
1-
12
#90440000000
0!
0%
b10 *
0-
02
b10 6
#90450000000
1!
1%
1-
12
#90460000000
0!
0%
b11 *
0-
02
b11 6
#90470000000
1!
1%
1-
12
15
#90480000000
0!
0%
b100 *
0-
02
b100 6
#90490000000
1!
1%
1-
12
#90500000000
0!
0%
b101 *
0-
02
b101 6
#90510000000
1!
1%
1-
12
#90520000000
0!
0%
b110 *
0-
02
b110 6
#90530000000
1!
1%
1-
12
#90540000000
0!
0%
b111 *
0-
02
b111 6
#90550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#90560000000
0!
0%
b0 *
0-
02
b0 6
#90570000000
1!
1%
1-
12
#90580000000
0!
0%
b1 *
0-
02
b1 6
#90590000000
1!
1%
1-
12
#90600000000
0!
0%
b10 *
0-
02
b10 6
#90610000000
1!
1%
1-
12
#90620000000
0!
0%
b11 *
0-
02
b11 6
#90630000000
1!
1%
1-
12
15
#90640000000
0!
0%
b100 *
0-
02
b100 6
#90650000000
1!
1%
1-
12
#90660000000
0!
0%
b101 *
0-
02
b101 6
#90670000000
1!
1%
1-
12
#90680000000
0!
0%
b110 *
0-
02
b110 6
#90690000000
1!
1%
1-
12
#90700000000
0!
0%
b111 *
0-
02
b111 6
#90710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#90720000000
0!
0%
b0 *
0-
02
b0 6
#90730000000
1!
1%
1-
12
#90740000000
0!
0%
b1 *
0-
02
b1 6
#90750000000
1!
1%
1-
12
#90760000000
0!
0%
b10 *
0-
02
b10 6
#90770000000
1!
1%
1-
12
#90780000000
0!
0%
b11 *
0-
02
b11 6
#90790000000
1!
1%
1-
12
15
#90800000000
0!
0%
b100 *
0-
02
b100 6
#90810000000
1!
1%
1-
12
#90820000000
0!
0%
b101 *
0-
02
b101 6
#90830000000
1!
1%
1-
12
#90840000000
0!
0%
b110 *
0-
02
b110 6
#90850000000
1!
1%
1-
12
#90860000000
0!
0%
b111 *
0-
02
b111 6
#90870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#90880000000
0!
0%
b0 *
0-
02
b0 6
#90890000000
1!
1%
1-
12
#90900000000
0!
0%
b1 *
0-
02
b1 6
#90910000000
1!
1%
1-
12
#90920000000
0!
0%
b10 *
0-
02
b10 6
#90930000000
1!
1%
1-
12
#90940000000
0!
0%
b11 *
0-
02
b11 6
#90950000000
1!
1%
1-
12
15
#90960000000
0!
0%
b100 *
0-
02
b100 6
#90970000000
1!
1%
1-
12
#90980000000
0!
0%
b101 *
0-
02
b101 6
#90990000000
1!
1%
1-
12
#91000000000
0!
0%
b110 *
0-
02
b110 6
#91010000000
1!
1%
1-
12
#91020000000
0!
0%
b111 *
0-
02
b111 6
#91030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#91040000000
0!
0%
b0 *
0-
02
b0 6
#91050000000
1!
1%
1-
12
#91060000000
0!
0%
b1 *
0-
02
b1 6
#91070000000
1!
1%
1-
12
#91080000000
0!
0%
b10 *
0-
02
b10 6
#91090000000
1!
1%
1-
12
#91100000000
0!
0%
b11 *
0-
02
b11 6
#91110000000
1!
1%
1-
12
15
#91120000000
0!
0%
b100 *
0-
02
b100 6
#91130000000
1!
1%
1-
12
#91140000000
0!
0%
b101 *
0-
02
b101 6
#91150000000
1!
1%
1-
12
#91160000000
0!
0%
b110 *
0-
02
b110 6
#91170000000
1!
1%
1-
12
#91180000000
0!
0%
b111 *
0-
02
b111 6
#91190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#91200000000
0!
0%
b0 *
0-
02
b0 6
#91210000000
1!
1%
1-
12
#91220000000
0!
0%
b1 *
0-
02
b1 6
#91230000000
1!
1%
1-
12
#91240000000
0!
0%
b10 *
0-
02
b10 6
#91250000000
1!
1%
1-
12
#91260000000
0!
0%
b11 *
0-
02
b11 6
#91270000000
1!
1%
1-
12
15
#91280000000
0!
0%
b100 *
0-
02
b100 6
#91290000000
1!
1%
1-
12
#91300000000
0!
0%
b101 *
0-
02
b101 6
#91310000000
1!
1%
1-
12
#91320000000
0!
0%
b110 *
0-
02
b110 6
#91330000000
1!
1%
1-
12
#91340000000
0!
0%
b111 *
0-
02
b111 6
#91350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#91360000000
0!
0%
b0 *
0-
02
b0 6
#91370000000
1!
1%
1-
12
#91380000000
0!
0%
b1 *
0-
02
b1 6
#91390000000
1!
1%
1-
12
#91400000000
0!
0%
b10 *
0-
02
b10 6
#91410000000
1!
1%
1-
12
#91420000000
0!
0%
b11 *
0-
02
b11 6
#91430000000
1!
1%
1-
12
15
#91440000000
0!
0%
b100 *
0-
02
b100 6
#91450000000
1!
1%
1-
12
#91460000000
0!
0%
b101 *
0-
02
b101 6
#91470000000
1!
1%
1-
12
#91480000000
0!
0%
b110 *
0-
02
b110 6
#91490000000
1!
1%
1-
12
#91500000000
0!
0%
b111 *
0-
02
b111 6
#91510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#91520000000
0!
0%
b0 *
0-
02
b0 6
#91530000000
1!
1%
1-
12
#91540000000
0!
0%
b1 *
0-
02
b1 6
#91550000000
1!
1%
1-
12
#91560000000
0!
0%
b10 *
0-
02
b10 6
#91570000000
1!
1%
1-
12
#91580000000
0!
0%
b11 *
0-
02
b11 6
#91590000000
1!
1%
1-
12
15
#91600000000
0!
0%
b100 *
0-
02
b100 6
#91610000000
1!
1%
1-
12
#91620000000
0!
0%
b101 *
0-
02
b101 6
#91630000000
1!
1%
1-
12
#91640000000
0!
0%
b110 *
0-
02
b110 6
#91650000000
1!
1%
1-
12
#91660000000
0!
0%
b111 *
0-
02
b111 6
#91670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#91680000000
0!
0%
b0 *
0-
02
b0 6
#91690000000
1!
1%
1-
12
#91700000000
0!
0%
b1 *
0-
02
b1 6
#91710000000
1!
1%
1-
12
#91720000000
0!
0%
b10 *
0-
02
b10 6
#91730000000
1!
1%
1-
12
#91740000000
0!
0%
b11 *
0-
02
b11 6
#91750000000
1!
1%
1-
12
15
#91760000000
0!
0%
b100 *
0-
02
b100 6
#91770000000
1!
1%
1-
12
#91780000000
0!
0%
b101 *
0-
02
b101 6
#91790000000
1!
1%
1-
12
#91800000000
0!
0%
b110 *
0-
02
b110 6
#91810000000
1!
1%
1-
12
#91820000000
0!
0%
b111 *
0-
02
b111 6
#91830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#91840000000
0!
0%
b0 *
0-
02
b0 6
#91850000000
1!
1%
1-
12
#91860000000
0!
0%
b1 *
0-
02
b1 6
#91870000000
1!
1%
1-
12
#91880000000
0!
0%
b10 *
0-
02
b10 6
#91890000000
1!
1%
1-
12
#91900000000
0!
0%
b11 *
0-
02
b11 6
#91910000000
1!
1%
1-
12
15
#91920000000
0!
0%
b100 *
0-
02
b100 6
#91930000000
1!
1%
1-
12
#91940000000
0!
0%
b101 *
0-
02
b101 6
#91950000000
1!
1%
1-
12
#91960000000
0!
0%
b110 *
0-
02
b110 6
#91970000000
1!
1%
1-
12
#91980000000
0!
0%
b111 *
0-
02
b111 6
#91990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#92000000000
0!
0%
b0 *
0-
02
b0 6
#92010000000
1!
1%
1-
12
#92020000000
0!
0%
b1 *
0-
02
b1 6
#92030000000
1!
1%
1-
12
#92040000000
0!
0%
b10 *
0-
02
b10 6
#92050000000
1!
1%
1-
12
#92060000000
0!
0%
b11 *
0-
02
b11 6
#92070000000
1!
1%
1-
12
15
#92080000000
0!
0%
b100 *
0-
02
b100 6
#92090000000
1!
1%
1-
12
#92100000000
0!
0%
b101 *
0-
02
b101 6
#92110000000
1!
1%
1-
12
#92120000000
0!
0%
b110 *
0-
02
b110 6
#92130000000
1!
1%
1-
12
#92140000000
0!
0%
b111 *
0-
02
b111 6
#92150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#92160000000
0!
0%
b0 *
0-
02
b0 6
#92170000000
1!
1%
1-
12
#92180000000
0!
0%
b1 *
0-
02
b1 6
#92190000000
1!
1%
1-
12
#92200000000
0!
0%
b10 *
0-
02
b10 6
#92210000000
1!
1%
1-
12
#92220000000
0!
0%
b11 *
0-
02
b11 6
#92230000000
1!
1%
1-
12
15
#92240000000
0!
0%
b100 *
0-
02
b100 6
#92250000000
1!
1%
1-
12
#92260000000
0!
0%
b101 *
0-
02
b101 6
#92270000000
1!
1%
1-
12
#92280000000
0!
0%
b110 *
0-
02
b110 6
#92290000000
1!
1%
1-
12
#92300000000
0!
0%
b111 *
0-
02
b111 6
#92310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#92320000000
0!
0%
b0 *
0-
02
b0 6
#92330000000
1!
1%
1-
12
#92340000000
0!
0%
b1 *
0-
02
b1 6
#92350000000
1!
1%
1-
12
#92360000000
0!
0%
b10 *
0-
02
b10 6
#92370000000
1!
1%
1-
12
#92380000000
0!
0%
b11 *
0-
02
b11 6
#92390000000
1!
1%
1-
12
15
#92400000000
0!
0%
b100 *
0-
02
b100 6
#92410000000
1!
1%
1-
12
#92420000000
0!
0%
b101 *
0-
02
b101 6
#92430000000
1!
1%
1-
12
#92440000000
0!
0%
b110 *
0-
02
b110 6
#92450000000
1!
1%
1-
12
#92460000000
0!
0%
b111 *
0-
02
b111 6
#92470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#92480000000
0!
0%
b0 *
0-
02
b0 6
#92490000000
1!
1%
1-
12
#92500000000
0!
0%
b1 *
0-
02
b1 6
#92510000000
1!
1%
1-
12
#92520000000
0!
0%
b10 *
0-
02
b10 6
#92530000000
1!
1%
1-
12
#92540000000
0!
0%
b11 *
0-
02
b11 6
#92550000000
1!
1%
1-
12
15
#92560000000
0!
0%
b100 *
0-
02
b100 6
#92570000000
1!
1%
1-
12
#92580000000
0!
0%
b101 *
0-
02
b101 6
#92590000000
1!
1%
1-
12
#92600000000
0!
0%
b110 *
0-
02
b110 6
#92610000000
1!
1%
1-
12
#92620000000
0!
0%
b111 *
0-
02
b111 6
#92630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#92640000000
0!
0%
b0 *
0-
02
b0 6
#92650000000
1!
1%
1-
12
#92660000000
0!
0%
b1 *
0-
02
b1 6
#92670000000
1!
1%
1-
12
#92680000000
0!
0%
b10 *
0-
02
b10 6
#92690000000
1!
1%
1-
12
#92700000000
0!
0%
b11 *
0-
02
b11 6
#92710000000
1!
1%
1-
12
15
#92720000000
0!
0%
b100 *
0-
02
b100 6
#92730000000
1!
1%
1-
12
#92740000000
0!
0%
b101 *
0-
02
b101 6
#92750000000
1!
1%
1-
12
#92760000000
0!
0%
b110 *
0-
02
b110 6
#92770000000
1!
1%
1-
12
#92780000000
0!
0%
b111 *
0-
02
b111 6
#92790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#92800000000
0!
0%
b0 *
0-
02
b0 6
#92810000000
1!
1%
1-
12
#92820000000
0!
0%
b1 *
0-
02
b1 6
#92830000000
1!
1%
1-
12
#92840000000
0!
0%
b10 *
0-
02
b10 6
#92850000000
1!
1%
1-
12
#92860000000
0!
0%
b11 *
0-
02
b11 6
#92870000000
1!
1%
1-
12
15
#92880000000
0!
0%
b100 *
0-
02
b100 6
#92890000000
1!
1%
1-
12
#92900000000
0!
0%
b101 *
0-
02
b101 6
#92910000000
1!
1%
1-
12
#92920000000
0!
0%
b110 *
0-
02
b110 6
#92930000000
1!
1%
1-
12
#92940000000
0!
0%
b111 *
0-
02
b111 6
#92950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#92960000000
0!
0%
b0 *
0-
02
b0 6
#92970000000
1!
1%
1-
12
#92980000000
0!
0%
b1 *
0-
02
b1 6
#92990000000
1!
1%
1-
12
#93000000000
0!
0%
b10 *
0-
02
b10 6
#93010000000
1!
1%
1-
12
#93020000000
0!
0%
b11 *
0-
02
b11 6
#93030000000
1!
1%
1-
12
15
#93040000000
0!
0%
b100 *
0-
02
b100 6
#93050000000
1!
1%
1-
12
#93060000000
0!
0%
b101 *
0-
02
b101 6
#93070000000
1!
1%
1-
12
#93080000000
0!
0%
b110 *
0-
02
b110 6
#93090000000
1!
1%
1-
12
#93100000000
0!
0%
b111 *
0-
02
b111 6
#93110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#93120000000
0!
0%
b0 *
0-
02
b0 6
#93130000000
1!
1%
1-
12
#93140000000
0!
0%
b1 *
0-
02
b1 6
#93150000000
1!
1%
1-
12
#93160000000
0!
0%
b10 *
0-
02
b10 6
#93170000000
1!
1%
1-
12
#93180000000
0!
0%
b11 *
0-
02
b11 6
#93190000000
1!
1%
1-
12
15
#93200000000
0!
0%
b100 *
0-
02
b100 6
#93210000000
1!
1%
1-
12
#93220000000
0!
0%
b101 *
0-
02
b101 6
#93230000000
1!
1%
1-
12
#93240000000
0!
0%
b110 *
0-
02
b110 6
#93250000000
1!
1%
1-
12
#93260000000
0!
0%
b111 *
0-
02
b111 6
#93270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#93280000000
0!
0%
b0 *
0-
02
b0 6
#93290000000
1!
1%
1-
12
#93300000000
0!
0%
b1 *
0-
02
b1 6
#93310000000
1!
1%
1-
12
#93320000000
0!
0%
b10 *
0-
02
b10 6
#93330000000
1!
1%
1-
12
#93340000000
0!
0%
b11 *
0-
02
b11 6
#93350000000
1!
1%
1-
12
15
#93360000000
0!
0%
b100 *
0-
02
b100 6
#93370000000
1!
1%
1-
12
#93380000000
0!
0%
b101 *
0-
02
b101 6
#93390000000
1!
1%
1-
12
#93400000000
0!
0%
b110 *
0-
02
b110 6
#93410000000
1!
1%
1-
12
#93420000000
0!
0%
b111 *
0-
02
b111 6
#93430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#93440000000
0!
0%
b0 *
0-
02
b0 6
#93450000000
1!
1%
1-
12
#93460000000
0!
0%
b1 *
0-
02
b1 6
#93470000000
1!
1%
1-
12
#93480000000
0!
0%
b10 *
0-
02
b10 6
#93490000000
1!
1%
1-
12
#93500000000
0!
0%
b11 *
0-
02
b11 6
#93510000000
1!
1%
1-
12
15
#93520000000
0!
0%
b100 *
0-
02
b100 6
#93530000000
1!
1%
1-
12
#93540000000
0!
0%
b101 *
0-
02
b101 6
#93550000000
1!
1%
1-
12
#93560000000
0!
0%
b110 *
0-
02
b110 6
#93570000000
1!
1%
1-
12
#93580000000
0!
0%
b111 *
0-
02
b111 6
#93590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#93600000000
0!
0%
b0 *
0-
02
b0 6
#93610000000
1!
1%
1-
12
#93620000000
0!
0%
b1 *
0-
02
b1 6
#93630000000
1!
1%
1-
12
#93640000000
0!
0%
b10 *
0-
02
b10 6
#93650000000
1!
1%
1-
12
#93660000000
0!
0%
b11 *
0-
02
b11 6
#93670000000
1!
1%
1-
12
15
#93680000000
0!
0%
b100 *
0-
02
b100 6
#93690000000
1!
1%
1-
12
#93700000000
0!
0%
b101 *
0-
02
b101 6
#93710000000
1!
1%
1-
12
#93720000000
0!
0%
b110 *
0-
02
b110 6
#93730000000
1!
1%
1-
12
#93740000000
0!
0%
b111 *
0-
02
b111 6
#93750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#93760000000
0!
0%
b0 *
0-
02
b0 6
#93770000000
1!
1%
1-
12
#93780000000
0!
0%
b1 *
0-
02
b1 6
#93790000000
1!
1%
1-
12
#93800000000
0!
0%
b10 *
0-
02
b10 6
#93810000000
1!
1%
1-
12
#93820000000
0!
0%
b11 *
0-
02
b11 6
#93830000000
1!
1%
1-
12
15
#93840000000
0!
0%
b100 *
0-
02
b100 6
#93850000000
1!
1%
1-
12
#93860000000
0!
0%
b101 *
0-
02
b101 6
#93870000000
1!
1%
1-
12
#93880000000
0!
0%
b110 *
0-
02
b110 6
#93890000000
1!
1%
1-
12
#93900000000
0!
0%
b111 *
0-
02
b111 6
#93910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#93920000000
0!
0%
b0 *
0-
02
b0 6
#93930000000
1!
1%
1-
12
#93940000000
0!
0%
b1 *
0-
02
b1 6
#93950000000
1!
1%
1-
12
#93960000000
0!
0%
b10 *
0-
02
b10 6
#93970000000
1!
1%
1-
12
#93980000000
0!
0%
b11 *
0-
02
b11 6
#93990000000
1!
1%
1-
12
15
#94000000000
0!
0%
b100 *
0-
02
b100 6
#94010000000
1!
1%
1-
12
#94020000000
0!
0%
b101 *
0-
02
b101 6
#94030000000
1!
1%
1-
12
#94040000000
0!
0%
b110 *
0-
02
b110 6
#94050000000
1!
1%
1-
12
#94060000000
0!
0%
b111 *
0-
02
b111 6
#94070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#94080000000
0!
0%
b0 *
0-
02
b0 6
#94090000000
1!
1%
1-
12
#94100000000
0!
0%
b1 *
0-
02
b1 6
#94110000000
1!
1%
1-
12
#94120000000
0!
0%
b10 *
0-
02
b10 6
#94130000000
1!
1%
1-
12
#94140000000
0!
0%
b11 *
0-
02
b11 6
#94150000000
1!
1%
1-
12
15
#94160000000
0!
0%
b100 *
0-
02
b100 6
#94170000000
1!
1%
1-
12
#94180000000
0!
0%
b101 *
0-
02
b101 6
#94190000000
1!
1%
1-
12
#94200000000
0!
0%
b110 *
0-
02
b110 6
#94210000000
1!
1%
1-
12
#94220000000
0!
0%
b111 *
0-
02
b111 6
#94230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#94240000000
0!
0%
b0 *
0-
02
b0 6
#94250000000
1!
1%
1-
12
#94260000000
0!
0%
b1 *
0-
02
b1 6
#94270000000
1!
1%
1-
12
#94280000000
0!
0%
b10 *
0-
02
b10 6
#94290000000
1!
1%
1-
12
#94300000000
0!
0%
b11 *
0-
02
b11 6
#94310000000
1!
1%
1-
12
15
#94320000000
0!
0%
b100 *
0-
02
b100 6
#94330000000
1!
1%
1-
12
#94340000000
0!
0%
b101 *
0-
02
b101 6
#94350000000
1!
1%
1-
12
#94360000000
0!
0%
b110 *
0-
02
b110 6
#94370000000
1!
1%
1-
12
#94380000000
0!
0%
b111 *
0-
02
b111 6
#94390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#94400000000
0!
0%
b0 *
0-
02
b0 6
#94410000000
1!
1%
1-
12
#94420000000
0!
0%
b1 *
0-
02
b1 6
#94430000000
1!
1%
1-
12
#94440000000
0!
0%
b10 *
0-
02
b10 6
#94450000000
1!
1%
1-
12
#94460000000
0!
0%
b11 *
0-
02
b11 6
#94470000000
1!
1%
1-
12
15
#94480000000
0!
0%
b100 *
0-
02
b100 6
#94490000000
1!
1%
1-
12
#94500000000
0!
0%
b101 *
0-
02
b101 6
#94510000000
1!
1%
1-
12
#94520000000
0!
0%
b110 *
0-
02
b110 6
#94530000000
1!
1%
1-
12
#94540000000
0!
0%
b111 *
0-
02
b111 6
#94550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#94560000000
0!
0%
b0 *
0-
02
b0 6
#94570000000
1!
1%
1-
12
#94580000000
0!
0%
b1 *
0-
02
b1 6
#94590000000
1!
1%
1-
12
#94600000000
0!
0%
b10 *
0-
02
b10 6
#94610000000
1!
1%
1-
12
#94620000000
0!
0%
b11 *
0-
02
b11 6
#94630000000
1!
1%
1-
12
15
#94640000000
0!
0%
b100 *
0-
02
b100 6
#94650000000
1!
1%
1-
12
#94660000000
0!
0%
b101 *
0-
02
b101 6
#94670000000
1!
1%
1-
12
#94680000000
0!
0%
b110 *
0-
02
b110 6
#94690000000
1!
1%
1-
12
#94700000000
0!
0%
b111 *
0-
02
b111 6
#94710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#94720000000
0!
0%
b0 *
0-
02
b0 6
#94730000000
1!
1%
1-
12
#94740000000
0!
0%
b1 *
0-
02
b1 6
#94750000000
1!
1%
1-
12
#94760000000
0!
0%
b10 *
0-
02
b10 6
#94770000000
1!
1%
1-
12
#94780000000
0!
0%
b11 *
0-
02
b11 6
#94790000000
1!
1%
1-
12
15
#94800000000
0!
0%
b100 *
0-
02
b100 6
#94810000000
1!
1%
1-
12
#94820000000
0!
0%
b101 *
0-
02
b101 6
#94830000000
1!
1%
1-
12
#94840000000
0!
0%
b110 *
0-
02
b110 6
#94850000000
1!
1%
1-
12
#94860000000
0!
0%
b111 *
0-
02
b111 6
#94870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#94880000000
0!
0%
b0 *
0-
02
b0 6
#94890000000
1!
1%
1-
12
#94900000000
0!
0%
b1 *
0-
02
b1 6
#94910000000
1!
1%
1-
12
#94920000000
0!
0%
b10 *
0-
02
b10 6
#94930000000
1!
1%
1-
12
#94940000000
0!
0%
b11 *
0-
02
b11 6
#94950000000
1!
1%
1-
12
15
#94960000000
0!
0%
b100 *
0-
02
b100 6
#94970000000
1!
1%
1-
12
#94980000000
0!
0%
b101 *
0-
02
b101 6
#94990000000
1!
1%
1-
12
#95000000000
0!
0%
b110 *
0-
02
b110 6
#95010000000
1!
1%
1-
12
#95020000000
0!
0%
b111 *
0-
02
b111 6
#95030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#95040000000
0!
0%
b0 *
0-
02
b0 6
#95050000000
1!
1%
1-
12
#95060000000
0!
0%
b1 *
0-
02
b1 6
#95070000000
1!
1%
1-
12
#95080000000
0!
0%
b10 *
0-
02
b10 6
#95090000000
1!
1%
1-
12
#95100000000
0!
0%
b11 *
0-
02
b11 6
#95110000000
1!
1%
1-
12
15
#95120000000
0!
0%
b100 *
0-
02
b100 6
#95130000000
1!
1%
1-
12
#95140000000
0!
0%
b101 *
0-
02
b101 6
#95150000000
1!
1%
1-
12
#95160000000
0!
0%
b110 *
0-
02
b110 6
#95170000000
1!
1%
1-
12
#95180000000
0!
0%
b111 *
0-
02
b111 6
#95190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#95200000000
0!
0%
b0 *
0-
02
b0 6
#95210000000
1!
1%
1-
12
#95220000000
0!
0%
b1 *
0-
02
b1 6
#95230000000
1!
1%
1-
12
#95240000000
0!
0%
b10 *
0-
02
b10 6
#95250000000
1!
1%
1-
12
#95260000000
0!
0%
b11 *
0-
02
b11 6
#95270000000
1!
1%
1-
12
15
#95280000000
0!
0%
b100 *
0-
02
b100 6
#95290000000
1!
1%
1-
12
#95300000000
0!
0%
b101 *
0-
02
b101 6
#95310000000
1!
1%
1-
12
#95320000000
0!
0%
b110 *
0-
02
b110 6
#95330000000
1!
1%
1-
12
#95340000000
0!
0%
b111 *
0-
02
b111 6
#95350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#95360000000
0!
0%
b0 *
0-
02
b0 6
#95370000000
1!
1%
1-
12
#95380000000
0!
0%
b1 *
0-
02
b1 6
#95390000000
1!
1%
1-
12
#95400000000
0!
0%
b10 *
0-
02
b10 6
#95410000000
1!
1%
1-
12
#95420000000
0!
0%
b11 *
0-
02
b11 6
#95430000000
1!
1%
1-
12
15
#95440000000
0!
0%
b100 *
0-
02
b100 6
#95450000000
1!
1%
1-
12
#95460000000
0!
0%
b101 *
0-
02
b101 6
#95470000000
1!
1%
1-
12
#95480000000
0!
0%
b110 *
0-
02
b110 6
#95490000000
1!
1%
1-
12
#95500000000
0!
0%
b111 *
0-
02
b111 6
#95510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#95520000000
0!
0%
b0 *
0-
02
b0 6
#95530000000
1!
1%
1-
12
#95540000000
0!
0%
b1 *
0-
02
b1 6
#95550000000
1!
1%
1-
12
#95560000000
0!
0%
b10 *
0-
02
b10 6
#95570000000
1!
1%
1-
12
#95580000000
0!
0%
b11 *
0-
02
b11 6
#95590000000
1!
1%
1-
12
15
#95600000000
0!
0%
b100 *
0-
02
b100 6
#95610000000
1!
1%
1-
12
#95620000000
0!
0%
b101 *
0-
02
b101 6
#95630000000
1!
1%
1-
12
#95640000000
0!
0%
b110 *
0-
02
b110 6
#95650000000
1!
1%
1-
12
#95660000000
0!
0%
b111 *
0-
02
b111 6
#95670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#95680000000
0!
0%
b0 *
0-
02
b0 6
#95690000000
1!
1%
1-
12
#95700000000
0!
0%
b1 *
0-
02
b1 6
#95710000000
1!
1%
1-
12
#95720000000
0!
0%
b10 *
0-
02
b10 6
#95730000000
1!
1%
1-
12
#95740000000
0!
0%
b11 *
0-
02
b11 6
#95750000000
1!
1%
1-
12
15
#95760000000
0!
0%
b100 *
0-
02
b100 6
#95770000000
1!
1%
1-
12
#95780000000
0!
0%
b101 *
0-
02
b101 6
#95790000000
1!
1%
1-
12
#95800000000
0!
0%
b110 *
0-
02
b110 6
#95810000000
1!
1%
1-
12
#95820000000
0!
0%
b111 *
0-
02
b111 6
#95830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#95840000000
0!
0%
b0 *
0-
02
b0 6
#95850000000
1!
1%
1-
12
#95860000000
0!
0%
b1 *
0-
02
b1 6
#95870000000
1!
1%
1-
12
#95880000000
0!
0%
b10 *
0-
02
b10 6
#95890000000
1!
1%
1-
12
#95900000000
0!
0%
b11 *
0-
02
b11 6
#95910000000
1!
1%
1-
12
15
#95920000000
0!
0%
b100 *
0-
02
b100 6
#95930000000
1!
1%
1-
12
#95940000000
0!
0%
b101 *
0-
02
b101 6
#95950000000
1!
1%
1-
12
#95960000000
0!
0%
b110 *
0-
02
b110 6
#95970000000
1!
1%
1-
12
#95980000000
0!
0%
b111 *
0-
02
b111 6
#95990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#96000000000
0!
0%
b0 *
0-
02
b0 6
#96010000000
1!
1%
1-
12
#96020000000
0!
0%
b1 *
0-
02
b1 6
#96030000000
1!
1%
1-
12
#96040000000
0!
0%
b10 *
0-
02
b10 6
#96050000000
1!
1%
1-
12
#96060000000
0!
0%
b11 *
0-
02
b11 6
#96070000000
1!
1%
1-
12
15
#96080000000
0!
0%
b100 *
0-
02
b100 6
#96090000000
1!
1%
1-
12
#96100000000
0!
0%
b101 *
0-
02
b101 6
#96110000000
1!
1%
1-
12
#96120000000
0!
0%
b110 *
0-
02
b110 6
#96130000000
1!
1%
1-
12
#96140000000
0!
0%
b111 *
0-
02
b111 6
#96150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#96160000000
0!
0%
b0 *
0-
02
b0 6
#96170000000
1!
1%
1-
12
#96180000000
0!
0%
b1 *
0-
02
b1 6
#96190000000
1!
1%
1-
12
#96200000000
0!
0%
b10 *
0-
02
b10 6
#96210000000
1!
1%
1-
12
#96220000000
0!
0%
b11 *
0-
02
b11 6
#96230000000
1!
1%
1-
12
15
#96240000000
0!
0%
b100 *
0-
02
b100 6
#96250000000
1!
1%
1-
12
#96260000000
0!
0%
b101 *
0-
02
b101 6
#96270000000
1!
1%
1-
12
#96280000000
0!
0%
b110 *
0-
02
b110 6
#96290000000
1!
1%
1-
12
#96300000000
0!
0%
b111 *
0-
02
b111 6
#96310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#96320000000
0!
0%
b0 *
0-
02
b0 6
#96330000000
1!
1%
1-
12
#96340000000
0!
0%
b1 *
0-
02
b1 6
#96350000000
1!
1%
1-
12
#96360000000
0!
0%
b10 *
0-
02
b10 6
#96370000000
1!
1%
1-
12
#96380000000
0!
0%
b11 *
0-
02
b11 6
#96390000000
1!
1%
1-
12
15
#96400000000
0!
0%
b100 *
0-
02
b100 6
#96410000000
1!
1%
1-
12
#96420000000
0!
0%
b101 *
0-
02
b101 6
#96430000000
1!
1%
1-
12
#96440000000
0!
0%
b110 *
0-
02
b110 6
#96450000000
1!
1%
1-
12
#96460000000
0!
0%
b111 *
0-
02
b111 6
#96470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#96480000000
0!
0%
b0 *
0-
02
b0 6
#96490000000
1!
1%
1-
12
#96500000000
0!
0%
b1 *
0-
02
b1 6
#96510000000
1!
1%
1-
12
#96520000000
0!
0%
b10 *
0-
02
b10 6
#96530000000
1!
1%
1-
12
#96540000000
0!
0%
b11 *
0-
02
b11 6
#96550000000
1!
1%
1-
12
15
#96560000000
0!
0%
b100 *
0-
02
b100 6
#96570000000
1!
1%
1-
12
#96580000000
0!
0%
b101 *
0-
02
b101 6
#96590000000
1!
1%
1-
12
#96600000000
0!
0%
b110 *
0-
02
b110 6
#96610000000
1!
1%
1-
12
#96620000000
0!
0%
b111 *
0-
02
b111 6
#96630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#96640000000
0!
0%
b0 *
0-
02
b0 6
#96650000000
1!
1%
1-
12
#96660000000
0!
0%
b1 *
0-
02
b1 6
#96670000000
1!
1%
1-
12
#96680000000
0!
0%
b10 *
0-
02
b10 6
#96690000000
1!
1%
1-
12
#96700000000
0!
0%
b11 *
0-
02
b11 6
#96710000000
1!
1%
1-
12
15
#96720000000
0!
0%
b100 *
0-
02
b100 6
#96730000000
1!
1%
1-
12
#96740000000
0!
0%
b101 *
0-
02
b101 6
#96750000000
1!
1%
1-
12
#96760000000
0!
0%
b110 *
0-
02
b110 6
#96770000000
1!
1%
1-
12
#96780000000
0!
0%
b111 *
0-
02
b111 6
#96790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#96800000000
0!
0%
b0 *
0-
02
b0 6
#96810000000
1!
1%
1-
12
#96820000000
0!
0%
b1 *
0-
02
b1 6
#96830000000
1!
1%
1-
12
#96840000000
0!
0%
b10 *
0-
02
b10 6
#96850000000
1!
1%
1-
12
#96860000000
0!
0%
b11 *
0-
02
b11 6
#96870000000
1!
1%
1-
12
15
#96880000000
0!
0%
b100 *
0-
02
b100 6
#96890000000
1!
1%
1-
12
#96900000000
0!
0%
b101 *
0-
02
b101 6
#96910000000
1!
1%
1-
12
#96920000000
0!
0%
b110 *
0-
02
b110 6
#96930000000
1!
1%
1-
12
#96940000000
0!
0%
b111 *
0-
02
b111 6
#96950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#96960000000
0!
0%
b0 *
0-
02
b0 6
#96970000000
1!
1%
1-
12
#96980000000
0!
0%
b1 *
0-
02
b1 6
#96990000000
1!
1%
1-
12
#97000000000
0!
0%
b10 *
0-
02
b10 6
#97010000000
1!
1%
1-
12
#97020000000
0!
0%
b11 *
0-
02
b11 6
#97030000000
1!
1%
1-
12
15
#97040000000
0!
0%
b100 *
0-
02
b100 6
#97050000000
1!
1%
1-
12
#97060000000
0!
0%
b101 *
0-
02
b101 6
#97070000000
1!
1%
1-
12
#97080000000
0!
0%
b110 *
0-
02
b110 6
#97090000000
1!
1%
1-
12
#97100000000
0!
0%
b111 *
0-
02
b111 6
#97110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#97120000000
0!
0%
b0 *
0-
02
b0 6
#97130000000
1!
1%
1-
12
#97140000000
0!
0%
b1 *
0-
02
b1 6
#97150000000
1!
1%
1-
12
#97160000000
0!
0%
b10 *
0-
02
b10 6
#97170000000
1!
1%
1-
12
#97180000000
0!
0%
b11 *
0-
02
b11 6
#97190000000
1!
1%
1-
12
15
#97200000000
0!
0%
b100 *
0-
02
b100 6
#97210000000
1!
1%
1-
12
#97220000000
0!
0%
b101 *
0-
02
b101 6
#97230000000
1!
1%
1-
12
#97240000000
0!
0%
b110 *
0-
02
b110 6
#97250000000
1!
1%
1-
12
#97260000000
0!
0%
b111 *
0-
02
b111 6
#97270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#97280000000
0!
0%
b0 *
0-
02
b0 6
#97290000000
1!
1%
1-
12
#97300000000
0!
0%
b1 *
0-
02
b1 6
#97310000000
1!
1%
1-
12
#97320000000
0!
0%
b10 *
0-
02
b10 6
#97330000000
1!
1%
1-
12
#97340000000
0!
0%
b11 *
0-
02
b11 6
#97350000000
1!
1%
1-
12
15
#97360000000
0!
0%
b100 *
0-
02
b100 6
#97370000000
1!
1%
1-
12
#97380000000
0!
0%
b101 *
0-
02
b101 6
#97390000000
1!
1%
1-
12
#97400000000
0!
0%
b110 *
0-
02
b110 6
#97410000000
1!
1%
1-
12
#97420000000
0!
0%
b111 *
0-
02
b111 6
#97430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#97440000000
0!
0%
b0 *
0-
02
b0 6
#97450000000
1!
1%
1-
12
#97460000000
0!
0%
b1 *
0-
02
b1 6
#97470000000
1!
1%
1-
12
#97480000000
0!
0%
b10 *
0-
02
b10 6
#97490000000
1!
1%
1-
12
#97500000000
0!
0%
b11 *
0-
02
b11 6
#97510000000
1!
1%
1-
12
15
#97520000000
0!
0%
b100 *
0-
02
b100 6
#97530000000
1!
1%
1-
12
#97540000000
0!
0%
b101 *
0-
02
b101 6
#97550000000
1!
1%
1-
12
#97560000000
0!
0%
b110 *
0-
02
b110 6
#97570000000
1!
1%
1-
12
#97580000000
0!
0%
b111 *
0-
02
b111 6
#97590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#97600000000
0!
0%
b0 *
0-
02
b0 6
#97610000000
1!
1%
1-
12
#97620000000
0!
0%
b1 *
0-
02
b1 6
#97630000000
1!
1%
1-
12
#97640000000
0!
0%
b10 *
0-
02
b10 6
#97650000000
1!
1%
1-
12
#97660000000
0!
0%
b11 *
0-
02
b11 6
#97670000000
1!
1%
1-
12
15
#97680000000
0!
0%
b100 *
0-
02
b100 6
#97690000000
1!
1%
1-
12
#97700000000
0!
0%
b101 *
0-
02
b101 6
#97710000000
1!
1%
1-
12
#97720000000
0!
0%
b110 *
0-
02
b110 6
#97730000000
1!
1%
1-
12
#97740000000
0!
0%
b111 *
0-
02
b111 6
#97750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#97760000000
0!
0%
b0 *
0-
02
b0 6
#97770000000
1!
1%
1-
12
#97780000000
0!
0%
b1 *
0-
02
b1 6
#97790000000
1!
1%
1-
12
#97800000000
0!
0%
b10 *
0-
02
b10 6
#97810000000
1!
1%
1-
12
#97820000000
0!
0%
b11 *
0-
02
b11 6
#97830000000
1!
1%
1-
12
15
#97840000000
0!
0%
b100 *
0-
02
b100 6
#97850000000
1!
1%
1-
12
#97860000000
0!
0%
b101 *
0-
02
b101 6
#97870000000
1!
1%
1-
12
#97880000000
0!
0%
b110 *
0-
02
b110 6
#97890000000
1!
1%
1-
12
#97900000000
0!
0%
b111 *
0-
02
b111 6
#97910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#97920000000
0!
0%
b0 *
0-
02
b0 6
#97930000000
1!
1%
1-
12
#97940000000
0!
0%
b1 *
0-
02
b1 6
#97950000000
1!
1%
1-
12
#97960000000
0!
0%
b10 *
0-
02
b10 6
#97970000000
1!
1%
1-
12
#97980000000
0!
0%
b11 *
0-
02
b11 6
#97990000000
1!
1%
1-
12
15
#98000000000
0!
0%
b100 *
0-
02
b100 6
#98010000000
1!
1%
1-
12
#98020000000
0!
0%
b101 *
0-
02
b101 6
#98030000000
1!
1%
1-
12
#98040000000
0!
0%
b110 *
0-
02
b110 6
#98050000000
1!
1%
1-
12
#98060000000
0!
0%
b111 *
0-
02
b111 6
#98070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#98080000000
0!
0%
b0 *
0-
02
b0 6
#98090000000
1!
1%
1-
12
#98100000000
0!
0%
b1 *
0-
02
b1 6
#98110000000
1!
1%
1-
12
#98120000000
0!
0%
b10 *
0-
02
b10 6
#98130000000
1!
1%
1-
12
#98140000000
0!
0%
b11 *
0-
02
b11 6
#98150000000
1!
1%
1-
12
15
#98160000000
0!
0%
b100 *
0-
02
b100 6
#98170000000
1!
1%
1-
12
#98180000000
0!
0%
b101 *
0-
02
b101 6
#98190000000
1!
1%
1-
12
#98200000000
0!
0%
b110 *
0-
02
b110 6
#98210000000
1!
1%
1-
12
#98220000000
0!
0%
b111 *
0-
02
b111 6
#98230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#98240000000
0!
0%
b0 *
0-
02
b0 6
#98250000000
1!
1%
1-
12
#98260000000
0!
0%
b1 *
0-
02
b1 6
#98270000000
1!
1%
1-
12
#98280000000
0!
0%
b10 *
0-
02
b10 6
#98290000000
1!
1%
1-
12
#98300000000
0!
0%
b11 *
0-
02
b11 6
#98310000000
1!
1%
1-
12
15
#98320000000
0!
0%
b100 *
0-
02
b100 6
#98330000000
1!
1%
1-
12
#98340000000
0!
0%
b101 *
0-
02
b101 6
#98350000000
1!
1%
1-
12
#98360000000
0!
0%
b110 *
0-
02
b110 6
#98370000000
1!
1%
1-
12
#98380000000
0!
0%
b111 *
0-
02
b111 6
#98390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#98400000000
0!
0%
b0 *
0-
02
b0 6
#98410000000
1!
1%
1-
12
#98420000000
0!
0%
b1 *
0-
02
b1 6
#98430000000
1!
1%
1-
12
#98440000000
0!
0%
b10 *
0-
02
b10 6
#98450000000
1!
1%
1-
12
#98460000000
0!
0%
b11 *
0-
02
b11 6
#98470000000
1!
1%
1-
12
15
#98480000000
0!
0%
b100 *
0-
02
b100 6
#98490000000
1!
1%
1-
12
#98500000000
0!
0%
b101 *
0-
02
b101 6
#98510000000
1!
1%
1-
12
#98520000000
0!
0%
b110 *
0-
02
b110 6
#98530000000
1!
1%
1-
12
#98540000000
0!
0%
b111 *
0-
02
b111 6
#98550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#98560000000
0!
0%
b0 *
0-
02
b0 6
#98570000000
1!
1%
1-
12
#98580000000
0!
0%
b1 *
0-
02
b1 6
#98590000000
1!
1%
1-
12
#98600000000
0!
0%
b10 *
0-
02
b10 6
#98610000000
1!
1%
1-
12
#98620000000
0!
0%
b11 *
0-
02
b11 6
#98630000000
1!
1%
1-
12
15
#98640000000
0!
0%
b100 *
0-
02
b100 6
#98650000000
1!
1%
1-
12
#98660000000
0!
0%
b101 *
0-
02
b101 6
#98670000000
1!
1%
1-
12
#98680000000
0!
0%
b110 *
0-
02
b110 6
#98690000000
1!
1%
1-
12
#98700000000
0!
0%
b111 *
0-
02
b111 6
#98710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#98720000000
0!
0%
b0 *
0-
02
b0 6
#98730000000
1!
1%
1-
12
#98740000000
0!
0%
b1 *
0-
02
b1 6
#98750000000
1!
1%
1-
12
#98760000000
0!
0%
b10 *
0-
02
b10 6
#98770000000
1!
1%
1-
12
#98780000000
0!
0%
b11 *
0-
02
b11 6
#98790000000
1!
1%
1-
12
15
#98800000000
0!
0%
b100 *
0-
02
b100 6
#98810000000
1!
1%
1-
12
#98820000000
0!
0%
b101 *
0-
02
b101 6
#98830000000
1!
1%
1-
12
#98840000000
0!
0%
b110 *
0-
02
b110 6
#98850000000
1!
1%
1-
12
#98860000000
0!
0%
b111 *
0-
02
b111 6
#98870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#98880000000
0!
0%
b0 *
0-
02
b0 6
#98890000000
1!
1%
1-
12
#98900000000
0!
0%
b1 *
0-
02
b1 6
#98910000000
1!
1%
1-
12
#98920000000
0!
0%
b10 *
0-
02
b10 6
#98930000000
1!
1%
1-
12
#98940000000
0!
0%
b11 *
0-
02
b11 6
#98950000000
1!
1%
1-
12
15
#98960000000
0!
0%
b100 *
0-
02
b100 6
#98970000000
1!
1%
1-
12
#98980000000
0!
0%
b101 *
0-
02
b101 6
#98990000000
1!
1%
1-
12
#99000000000
0!
0%
b110 *
0-
02
b110 6
#99010000000
1!
1%
1-
12
#99020000000
0!
0%
b111 *
0-
02
b111 6
#99030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#99040000000
0!
0%
b0 *
0-
02
b0 6
#99050000000
1!
1%
1-
12
#99060000000
0!
0%
b1 *
0-
02
b1 6
#99070000000
1!
1%
1-
12
#99080000000
0!
0%
b10 *
0-
02
b10 6
#99090000000
1!
1%
1-
12
#99100000000
0!
0%
b11 *
0-
02
b11 6
#99110000000
1!
1%
1-
12
15
#99120000000
0!
0%
b100 *
0-
02
b100 6
#99130000000
1!
1%
1-
12
#99140000000
0!
0%
b101 *
0-
02
b101 6
#99150000000
1!
1%
1-
12
#99160000000
0!
0%
b110 *
0-
02
b110 6
#99170000000
1!
1%
1-
12
#99180000000
0!
0%
b111 *
0-
02
b111 6
#99190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#99200000000
0!
0%
b0 *
0-
02
b0 6
#99210000000
1!
1%
1-
12
#99220000000
0!
0%
b1 *
0-
02
b1 6
#99230000000
1!
1%
1-
12
#99240000000
0!
0%
b10 *
0-
02
b10 6
#99250000000
1!
1%
1-
12
#99260000000
0!
0%
b11 *
0-
02
b11 6
#99270000000
1!
1%
1-
12
15
#99280000000
0!
0%
b100 *
0-
02
b100 6
#99290000000
1!
1%
1-
12
#99300000000
0!
0%
b101 *
0-
02
b101 6
#99310000000
1!
1%
1-
12
#99320000000
0!
0%
b110 *
0-
02
b110 6
#99330000000
1!
1%
1-
12
#99340000000
0!
0%
b111 *
0-
02
b111 6
#99350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#99360000000
0!
0%
b0 *
0-
02
b0 6
#99370000000
1!
1%
1-
12
#99380000000
0!
0%
b1 *
0-
02
b1 6
#99390000000
1!
1%
1-
12
#99400000000
0!
0%
b10 *
0-
02
b10 6
#99410000000
1!
1%
1-
12
#99420000000
0!
0%
b11 *
0-
02
b11 6
#99430000000
1!
1%
1-
12
15
#99440000000
0!
0%
b100 *
0-
02
b100 6
#99450000000
1!
1%
1-
12
#99460000000
0!
0%
b101 *
0-
02
b101 6
#99470000000
1!
1%
1-
12
#99480000000
0!
0%
b110 *
0-
02
b110 6
#99490000000
1!
1%
1-
12
#99500000000
0!
0%
b111 *
0-
02
b111 6
#99510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#99520000000
0!
0%
b0 *
0-
02
b0 6
#99530000000
1!
1%
1-
12
#99540000000
0!
0%
b1 *
0-
02
b1 6
#99550000000
1!
1%
1-
12
#99560000000
0!
0%
b10 *
0-
02
b10 6
#99570000000
1!
1%
1-
12
#99580000000
0!
0%
b11 *
0-
02
b11 6
#99590000000
1!
1%
1-
12
15
#99600000000
0!
0%
b100 *
0-
02
b100 6
#99610000000
1!
1%
1-
12
#99620000000
0!
0%
b101 *
0-
02
b101 6
#99630000000
1!
1%
1-
12
#99640000000
0!
0%
b110 *
0-
02
b110 6
#99650000000
1!
1%
1-
12
#99660000000
0!
0%
b111 *
0-
02
b111 6
#99670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#99680000000
0!
0%
b0 *
0-
02
b0 6
#99690000000
1!
1%
1-
12
#99700000000
0!
0%
b1 *
0-
02
b1 6
#99710000000
1!
1%
1-
12
#99720000000
0!
0%
b10 *
0-
02
b10 6
#99730000000
1!
1%
1-
12
#99740000000
0!
0%
b11 *
0-
02
b11 6
#99750000000
1!
1%
1-
12
15
#99760000000
0!
0%
b100 *
0-
02
b100 6
#99770000000
1!
1%
1-
12
#99780000000
0!
0%
b101 *
0-
02
b101 6
#99790000000
1!
1%
1-
12
#99800000000
0!
0%
b110 *
0-
02
b110 6
#99810000000
1!
1%
1-
12
#99820000000
0!
0%
b111 *
0-
02
b111 6
#99830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#99840000000
0!
0%
b0 *
0-
02
b0 6
#99850000000
1!
1%
1-
12
#99860000000
0!
0%
b1 *
0-
02
b1 6
#99870000000
1!
1%
1-
12
#99880000000
0!
0%
b10 *
0-
02
b10 6
#99890000000
1!
1%
1-
12
#99900000000
0!
0%
b11 *
0-
02
b11 6
#99910000000
1!
1%
1-
12
15
#99920000000
0!
0%
b100 *
0-
02
b100 6
#99930000000
1!
1%
1-
12
#99940000000
0!
0%
b101 *
0-
02
b101 6
#99950000000
1!
1%
1-
12
#99960000000
0!
0%
b110 *
0-
02
b110 6
#99970000000
1!
1%
1-
12
#99980000000
0!
0%
b111 *
0-
02
b111 6
#99990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#100000000000
0!
0%
b0 *
0-
02
b0 6
#100010000000
1!
1%
1-
12
#100020000000
0!
0%
b1 *
0-
02
b1 6
#100030000000
1!
1%
1-
12
#100040000000
0!
0%
b10 *
0-
02
b10 6
#100050000000
1!
1%
1-
12
#100060000000
0!
0%
b11 *
0-
02
b11 6
#100070000000
1!
1%
1-
12
15
#100080000000
0!
0%
b100 *
0-
02
b100 6
#100090000000
1!
1%
1-
12
#100100000000
0!
0%
b101 *
0-
02
b101 6
#100110000000
1!
1%
1-
12
#100120000000
0!
0%
b110 *
0-
02
b110 6
#100130000000
1!
1%
1-
12
#100140000000
0!
0%
b111 *
0-
02
b111 6
#100150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#100160000000
0!
0%
b0 *
0-
02
b0 6
#100170000000
1!
1%
1-
12
#100180000000
0!
0%
b1 *
0-
02
b1 6
#100190000000
1!
1%
1-
12
#100200000000
0!
0%
b10 *
0-
02
b10 6
#100210000000
1!
1%
1-
12
#100220000000
0!
0%
b11 *
0-
02
b11 6
#100230000000
1!
1%
1-
12
15
#100240000000
0!
0%
b100 *
0-
02
b100 6
#100250000000
1!
1%
1-
12
#100260000000
0!
0%
b101 *
0-
02
b101 6
#100270000000
1!
1%
1-
12
#100280000000
0!
0%
b110 *
0-
02
b110 6
#100290000000
1!
1%
1-
12
#100300000000
0!
0%
b111 *
0-
02
b111 6
#100310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#100320000000
0!
0%
b0 *
0-
02
b0 6
#100330000000
1!
1%
1-
12
#100340000000
0!
0%
b1 *
0-
02
b1 6
#100350000000
1!
1%
1-
12
#100360000000
0!
0%
b10 *
0-
02
b10 6
#100370000000
1!
1%
1-
12
#100380000000
0!
0%
b11 *
0-
02
b11 6
#100390000000
1!
1%
1-
12
15
#100400000000
0!
0%
b100 *
0-
02
b100 6
#100410000000
1!
1%
1-
12
#100420000000
0!
0%
b101 *
0-
02
b101 6
#100430000000
1!
1%
1-
12
#100440000000
0!
0%
b110 *
0-
02
b110 6
#100450000000
1!
1%
1-
12
#100460000000
0!
0%
b111 *
0-
02
b111 6
#100470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#100480000000
0!
0%
b0 *
0-
02
b0 6
#100490000000
1!
1%
1-
12
#100500000000
0!
0%
b1 *
0-
02
b1 6
#100510000000
1!
1%
1-
12
#100520000000
0!
0%
b10 *
0-
02
b10 6
#100530000000
1!
1%
1-
12
#100540000000
0!
0%
b11 *
0-
02
b11 6
#100550000000
1!
1%
1-
12
15
#100560000000
0!
0%
b100 *
0-
02
b100 6
#100570000000
1!
1%
1-
12
#100580000000
0!
0%
b101 *
0-
02
b101 6
#100590000000
1!
1%
1-
12
#100600000000
0!
0%
b110 *
0-
02
b110 6
#100610000000
1!
1%
1-
12
#100620000000
0!
0%
b111 *
0-
02
b111 6
#100630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#100640000000
0!
0%
b0 *
0-
02
b0 6
#100650000000
1!
1%
1-
12
#100660000000
0!
0%
b1 *
0-
02
b1 6
#100670000000
1!
1%
1-
12
#100680000000
0!
0%
b10 *
0-
02
b10 6
#100690000000
1!
1%
1-
12
#100700000000
0!
0%
b11 *
0-
02
b11 6
#100710000000
1!
1%
1-
12
15
#100720000000
0!
0%
b100 *
0-
02
b100 6
#100730000000
1!
1%
1-
12
#100740000000
0!
0%
b101 *
0-
02
b101 6
#100750000000
1!
1%
1-
12
#100760000000
0!
0%
b110 *
0-
02
b110 6
#100770000000
1!
1%
1-
12
#100780000000
0!
0%
b111 *
0-
02
b111 6
#100790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#100800000000
0!
0%
b0 *
0-
02
b0 6
#100810000000
1!
1%
1-
12
#100820000000
0!
0%
b1 *
0-
02
b1 6
#100830000000
1!
1%
1-
12
#100840000000
0!
0%
b10 *
0-
02
b10 6
#100850000000
1!
1%
1-
12
#100860000000
0!
0%
b11 *
0-
02
b11 6
#100870000000
1!
1%
1-
12
15
#100880000000
0!
0%
b100 *
0-
02
b100 6
#100890000000
1!
1%
1-
12
#100900000000
0!
0%
b101 *
0-
02
b101 6
#100910000000
1!
1%
1-
12
#100920000000
0!
0%
b110 *
0-
02
b110 6
#100930000000
1!
1%
1-
12
#100940000000
0!
0%
b111 *
0-
02
b111 6
#100950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#100960000000
0!
0%
b0 *
0-
02
b0 6
#100970000000
1!
1%
1-
12
#100980000000
0!
0%
b1 *
0-
02
b1 6
#100990000000
1!
1%
1-
12
#101000000000
0!
0%
b10 *
0-
02
b10 6
#101010000000
1!
1%
1-
12
#101020000000
0!
0%
b11 *
0-
02
b11 6
#101030000000
1!
1%
1-
12
15
#101040000000
0!
0%
b100 *
0-
02
b100 6
#101050000000
1!
1%
1-
12
#101060000000
0!
0%
b101 *
0-
02
b101 6
#101070000000
1!
1%
1-
12
#101080000000
0!
0%
b110 *
0-
02
b110 6
#101090000000
1!
1%
1-
12
#101100000000
0!
0%
b111 *
0-
02
b111 6
#101110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#101120000000
0!
0%
b0 *
0-
02
b0 6
#101130000000
1!
1%
1-
12
#101140000000
0!
0%
b1 *
0-
02
b1 6
#101150000000
1!
1%
1-
12
#101160000000
0!
0%
b10 *
0-
02
b10 6
#101170000000
1!
1%
1-
12
#101180000000
0!
0%
b11 *
0-
02
b11 6
#101190000000
1!
1%
1-
12
15
#101200000000
0!
0%
b100 *
0-
02
b100 6
#101210000000
1!
1%
1-
12
#101220000000
0!
0%
b101 *
0-
02
b101 6
#101230000000
1!
1%
1-
12
#101240000000
0!
0%
b110 *
0-
02
b110 6
#101250000000
1!
1%
1-
12
#101260000000
0!
0%
b111 *
0-
02
b111 6
#101270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#101280000000
0!
0%
b0 *
0-
02
b0 6
#101290000000
1!
1%
1-
12
#101300000000
0!
0%
b1 *
0-
02
b1 6
#101310000000
1!
1%
1-
12
#101320000000
0!
0%
b10 *
0-
02
b10 6
#101330000000
1!
1%
1-
12
#101340000000
0!
0%
b11 *
0-
02
b11 6
#101350000000
1!
1%
1-
12
15
#101360000000
0!
0%
b100 *
0-
02
b100 6
#101370000000
1!
1%
1-
12
#101380000000
0!
0%
b101 *
0-
02
b101 6
#101390000000
1!
1%
1-
12
#101400000000
0!
0%
b110 *
0-
02
b110 6
#101410000000
1!
1%
1-
12
#101420000000
0!
0%
b111 *
0-
02
b111 6
#101430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#101440000000
0!
0%
b0 *
0-
02
b0 6
#101450000000
1!
1%
1-
12
#101460000000
0!
0%
b1 *
0-
02
b1 6
#101470000000
1!
1%
1-
12
#101480000000
0!
0%
b10 *
0-
02
b10 6
#101490000000
1!
1%
1-
12
#101500000000
0!
0%
b11 *
0-
02
b11 6
#101510000000
1!
1%
1-
12
15
#101520000000
0!
0%
b100 *
0-
02
b100 6
#101530000000
1!
1%
1-
12
#101540000000
0!
0%
b101 *
0-
02
b101 6
#101550000000
1!
1%
1-
12
#101560000000
0!
0%
b110 *
0-
02
b110 6
#101570000000
1!
1%
1-
12
#101580000000
0!
0%
b111 *
0-
02
b111 6
#101590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#101600000000
0!
0%
b0 *
0-
02
b0 6
#101610000000
1!
1%
1-
12
#101620000000
0!
0%
b1 *
0-
02
b1 6
#101630000000
1!
1%
1-
12
#101640000000
0!
0%
b10 *
0-
02
b10 6
#101650000000
1!
1%
1-
12
#101660000000
0!
0%
b11 *
0-
02
b11 6
#101670000000
1!
1%
1-
12
15
#101680000000
0!
0%
b100 *
0-
02
b100 6
#101690000000
1!
1%
1-
12
#101700000000
0!
0%
b101 *
0-
02
b101 6
#101710000000
1!
1%
1-
12
#101720000000
0!
0%
b110 *
0-
02
b110 6
#101730000000
1!
1%
1-
12
#101740000000
0!
0%
b111 *
0-
02
b111 6
#101750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#101760000000
0!
0%
b0 *
0-
02
b0 6
#101770000000
1!
1%
1-
12
#101780000000
0!
0%
b1 *
0-
02
b1 6
#101790000000
1!
1%
1-
12
#101800000000
0!
0%
b10 *
0-
02
b10 6
#101810000000
1!
1%
1-
12
#101820000000
0!
0%
b11 *
0-
02
b11 6
#101830000000
1!
1%
1-
12
15
#101840000000
0!
0%
b100 *
0-
02
b100 6
#101850000000
1!
1%
1-
12
#101860000000
0!
0%
b101 *
0-
02
b101 6
#101870000000
1!
1%
1-
12
#101880000000
0!
0%
b110 *
0-
02
b110 6
#101890000000
1!
1%
1-
12
#101900000000
0!
0%
b111 *
0-
02
b111 6
#101910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#101920000000
0!
0%
b0 *
0-
02
b0 6
#101930000000
1!
1%
1-
12
#101940000000
0!
0%
b1 *
0-
02
b1 6
#101950000000
1!
1%
1-
12
#101960000000
0!
0%
b10 *
0-
02
b10 6
#101970000000
1!
1%
1-
12
#101980000000
0!
0%
b11 *
0-
02
b11 6
#101990000000
1!
1%
1-
12
15
#102000000000
0!
0%
b100 *
0-
02
b100 6
#102010000000
1!
1%
1-
12
#102020000000
0!
0%
b101 *
0-
02
b101 6
#102030000000
1!
1%
1-
12
#102040000000
0!
0%
b110 *
0-
02
b110 6
#102050000000
1!
1%
1-
12
#102060000000
0!
0%
b111 *
0-
02
b111 6
#102070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#102080000000
0!
0%
b0 *
0-
02
b0 6
#102090000000
1!
1%
1-
12
#102100000000
0!
0%
b1 *
0-
02
b1 6
#102110000000
1!
1%
1-
12
#102120000000
0!
0%
b10 *
0-
02
b10 6
#102130000000
1!
1%
1-
12
#102140000000
0!
0%
b11 *
0-
02
b11 6
#102150000000
1!
1%
1-
12
15
#102160000000
0!
0%
b100 *
0-
02
b100 6
#102170000000
1!
1%
1-
12
#102180000000
0!
0%
b101 *
0-
02
b101 6
#102190000000
1!
1%
1-
12
#102200000000
0!
0%
b110 *
0-
02
b110 6
#102210000000
1!
1%
1-
12
#102220000000
0!
0%
b111 *
0-
02
b111 6
#102230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#102240000000
0!
0%
b0 *
0-
02
b0 6
#102250000000
1!
1%
1-
12
#102260000000
0!
0%
b1 *
0-
02
b1 6
#102270000000
1!
1%
1-
12
#102280000000
0!
0%
b10 *
0-
02
b10 6
#102290000000
1!
1%
1-
12
#102300000000
0!
0%
b11 *
0-
02
b11 6
#102310000000
1!
1%
1-
12
15
#102320000000
0!
0%
b100 *
0-
02
b100 6
#102330000000
1!
1%
1-
12
#102340000000
0!
0%
b101 *
0-
02
b101 6
#102350000000
1!
1%
1-
12
#102360000000
0!
0%
b110 *
0-
02
b110 6
#102370000000
1!
1%
1-
12
#102380000000
0!
0%
b111 *
0-
02
b111 6
#102390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#102400000000
0!
0%
b0 *
0-
02
b0 6
#102410000000
1!
1%
1-
12
#102420000000
0!
0%
b1 *
0-
02
b1 6
#102430000000
1!
1%
1-
12
#102440000000
0!
0%
b10 *
0-
02
b10 6
#102450000000
1!
1%
1-
12
#102460000000
0!
0%
b11 *
0-
02
b11 6
#102470000000
1!
1%
1-
12
15
#102480000000
0!
0%
b100 *
0-
02
b100 6
#102490000000
1!
1%
1-
12
#102500000000
0!
0%
b101 *
0-
02
b101 6
#102510000000
1!
1%
1-
12
#102520000000
0!
0%
b110 *
0-
02
b110 6
#102530000000
1!
1%
1-
12
#102540000000
0!
0%
b111 *
0-
02
b111 6
#102550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#102560000000
0!
0%
b0 *
0-
02
b0 6
#102570000000
1!
1%
1-
12
#102580000000
0!
0%
b1 *
0-
02
b1 6
#102590000000
1!
1%
1-
12
#102600000000
0!
0%
b10 *
0-
02
b10 6
#102610000000
1!
1%
1-
12
#102620000000
0!
0%
b11 *
0-
02
b11 6
#102630000000
1!
1%
1-
12
15
#102640000000
0!
0%
b100 *
0-
02
b100 6
#102650000000
1!
1%
1-
12
#102660000000
0!
0%
b101 *
0-
02
b101 6
#102670000000
1!
1%
1-
12
#102680000000
0!
0%
b110 *
0-
02
b110 6
#102690000000
1!
1%
1-
12
#102700000000
0!
0%
b111 *
0-
02
b111 6
#102710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#102720000000
0!
0%
b0 *
0-
02
b0 6
#102730000000
1!
1%
1-
12
#102740000000
0!
0%
b1 *
0-
02
b1 6
#102750000000
1!
1%
1-
12
#102760000000
0!
0%
b10 *
0-
02
b10 6
#102770000000
1!
1%
1-
12
#102780000000
0!
0%
b11 *
0-
02
b11 6
#102790000000
1!
1%
1-
12
15
#102800000000
0!
0%
b100 *
0-
02
b100 6
#102810000000
1!
1%
1-
12
#102820000000
0!
0%
b101 *
0-
02
b101 6
#102830000000
1!
1%
1-
12
#102840000000
0!
0%
b110 *
0-
02
b110 6
#102850000000
1!
1%
1-
12
#102860000000
0!
0%
b111 *
0-
02
b111 6
#102870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#102880000000
0!
0%
b0 *
0-
02
b0 6
#102890000000
1!
1%
1-
12
#102900000000
0!
0%
b1 *
0-
02
b1 6
#102910000000
1!
1%
1-
12
#102920000000
0!
0%
b10 *
0-
02
b10 6
#102930000000
1!
1%
1-
12
#102940000000
0!
0%
b11 *
0-
02
b11 6
#102950000000
1!
1%
1-
12
15
#102960000000
0!
0%
b100 *
0-
02
b100 6
#102970000000
1!
1%
1-
12
#102980000000
0!
0%
b101 *
0-
02
b101 6
#102990000000
1!
1%
1-
12
#103000000000
0!
0%
b110 *
0-
02
b110 6
#103010000000
1!
1%
1-
12
#103020000000
0!
0%
b111 *
0-
02
b111 6
#103030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#103040000000
0!
0%
b0 *
0-
02
b0 6
#103050000000
1!
1%
1-
12
#103060000000
0!
0%
b1 *
0-
02
b1 6
#103070000000
1!
1%
1-
12
#103080000000
0!
0%
b10 *
0-
02
b10 6
#103090000000
1!
1%
1-
12
#103100000000
0!
0%
b11 *
0-
02
b11 6
#103110000000
1!
1%
1-
12
15
#103120000000
0!
0%
b100 *
0-
02
b100 6
#103130000000
1!
1%
1-
12
#103140000000
0!
0%
b101 *
0-
02
b101 6
#103150000000
1!
1%
1-
12
#103160000000
0!
0%
b110 *
0-
02
b110 6
#103170000000
1!
1%
1-
12
#103180000000
0!
0%
b111 *
0-
02
b111 6
#103190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#103200000000
0!
0%
b0 *
0-
02
b0 6
#103210000000
1!
1%
1-
12
#103220000000
0!
0%
b1 *
0-
02
b1 6
#103230000000
1!
1%
1-
12
#103240000000
0!
0%
b10 *
0-
02
b10 6
#103250000000
1!
1%
1-
12
#103260000000
0!
0%
b11 *
0-
02
b11 6
#103270000000
1!
1%
1-
12
15
#103280000000
0!
0%
b100 *
0-
02
b100 6
#103290000000
1!
1%
1-
12
#103300000000
0!
0%
b101 *
0-
02
b101 6
#103310000000
1!
1%
1-
12
#103320000000
0!
0%
b110 *
0-
02
b110 6
#103330000000
1!
1%
1-
12
#103340000000
0!
0%
b111 *
0-
02
b111 6
#103350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#103360000000
0!
0%
b0 *
0-
02
b0 6
#103370000000
1!
1%
1-
12
#103380000000
0!
0%
b1 *
0-
02
b1 6
#103390000000
1!
1%
1-
12
#103400000000
0!
0%
b10 *
0-
02
b10 6
#103410000000
1!
1%
1-
12
#103420000000
0!
0%
b11 *
0-
02
b11 6
#103430000000
1!
1%
1-
12
15
#103440000000
0!
0%
b100 *
0-
02
b100 6
#103450000000
1!
1%
1-
12
#103460000000
0!
0%
b101 *
0-
02
b101 6
#103470000000
1!
1%
1-
12
#103480000000
0!
0%
b110 *
0-
02
b110 6
#103490000000
1!
1%
1-
12
#103500000000
0!
0%
b111 *
0-
02
b111 6
#103510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#103520000000
0!
0%
b0 *
0-
02
b0 6
#103530000000
1!
1%
1-
12
#103540000000
0!
0%
b1 *
0-
02
b1 6
#103550000000
1!
1%
1-
12
#103560000000
0!
0%
b10 *
0-
02
b10 6
#103570000000
1!
1%
1-
12
#103580000000
0!
0%
b11 *
0-
02
b11 6
#103590000000
1!
1%
1-
12
15
#103600000000
0!
0%
b100 *
0-
02
b100 6
#103610000000
1!
1%
1-
12
#103620000000
0!
0%
b101 *
0-
02
b101 6
#103630000000
1!
1%
1-
12
#103640000000
0!
0%
b110 *
0-
02
b110 6
#103650000000
1!
1%
1-
12
#103660000000
0!
0%
b111 *
0-
02
b111 6
#103670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#103680000000
0!
0%
b0 *
0-
02
b0 6
#103690000000
1!
1%
1-
12
#103700000000
0!
0%
b1 *
0-
02
b1 6
#103710000000
1!
1%
1-
12
#103720000000
0!
0%
b10 *
0-
02
b10 6
#103730000000
1!
1%
1-
12
#103740000000
0!
0%
b11 *
0-
02
b11 6
#103750000000
1!
1%
1-
12
15
#103760000000
0!
0%
b100 *
0-
02
b100 6
#103770000000
1!
1%
1-
12
#103780000000
0!
0%
b101 *
0-
02
b101 6
#103790000000
1!
1%
1-
12
#103800000000
0!
0%
b110 *
0-
02
b110 6
#103810000000
1!
1%
1-
12
#103820000000
0!
0%
b111 *
0-
02
b111 6
#103830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#103840000000
0!
0%
b0 *
0-
02
b0 6
#103850000000
1!
1%
1-
12
#103860000000
0!
0%
b1 *
0-
02
b1 6
#103870000000
1!
1%
1-
12
#103880000000
0!
0%
b10 *
0-
02
b10 6
#103890000000
1!
1%
1-
12
#103900000000
0!
0%
b11 *
0-
02
b11 6
#103910000000
1!
1%
1-
12
15
#103920000000
0!
0%
b100 *
0-
02
b100 6
#103930000000
1!
1%
1-
12
#103940000000
0!
0%
b101 *
0-
02
b101 6
#103950000000
1!
1%
1-
12
#103960000000
0!
0%
b110 *
0-
02
b110 6
#103970000000
1!
1%
1-
12
#103980000000
0!
0%
b111 *
0-
02
b111 6
#103990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#104000000000
0!
0%
b0 *
0-
02
b0 6
#104010000000
1!
1%
1-
12
#104020000000
0!
0%
b1 *
0-
02
b1 6
#104030000000
1!
1%
1-
12
#104040000000
0!
0%
b10 *
0-
02
b10 6
#104050000000
1!
1%
1-
12
#104060000000
0!
0%
b11 *
0-
02
b11 6
#104070000000
1!
1%
1-
12
15
#104080000000
0!
0%
b100 *
0-
02
b100 6
#104090000000
1!
1%
1-
12
#104100000000
0!
0%
b101 *
0-
02
b101 6
#104110000000
1!
1%
1-
12
#104120000000
0!
0%
b110 *
0-
02
b110 6
#104130000000
1!
1%
1-
12
#104140000000
0!
0%
b111 *
0-
02
b111 6
#104150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#104160000000
0!
0%
b0 *
0-
02
b0 6
#104170000000
1!
1%
1-
12
#104180000000
0!
0%
b1 *
0-
02
b1 6
#104190000000
1!
1%
1-
12
#104200000000
0!
0%
b10 *
0-
02
b10 6
#104210000000
1!
1%
1-
12
#104220000000
0!
0%
b11 *
0-
02
b11 6
#104230000000
1!
1%
1-
12
15
#104240000000
0!
0%
b100 *
0-
02
b100 6
#104250000000
1!
1%
1-
12
#104260000000
0!
0%
b101 *
0-
02
b101 6
#104270000000
1!
1%
1-
12
#104280000000
0!
0%
b110 *
0-
02
b110 6
#104290000000
1!
1%
1-
12
#104300000000
0!
0%
b111 *
0-
02
b111 6
#104310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#104320000000
0!
0%
b0 *
0-
02
b0 6
#104330000000
1!
1%
1-
12
#104340000000
0!
0%
b1 *
0-
02
b1 6
#104350000000
1!
1%
1-
12
#104360000000
0!
0%
b10 *
0-
02
b10 6
#104370000000
1!
1%
1-
12
#104380000000
0!
0%
b11 *
0-
02
b11 6
#104390000000
1!
1%
1-
12
15
#104400000000
0!
0%
b100 *
0-
02
b100 6
#104410000000
1!
1%
1-
12
#104420000000
0!
0%
b101 *
0-
02
b101 6
#104430000000
1!
1%
1-
12
#104440000000
0!
0%
b110 *
0-
02
b110 6
#104450000000
1!
1%
1-
12
#104460000000
0!
0%
b111 *
0-
02
b111 6
#104470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#104480000000
0!
0%
b0 *
0-
02
b0 6
#104490000000
1!
1%
1-
12
#104500000000
0!
0%
b1 *
0-
02
b1 6
#104510000000
1!
1%
1-
12
#104520000000
0!
0%
b10 *
0-
02
b10 6
#104530000000
1!
1%
1-
12
#104540000000
0!
0%
b11 *
0-
02
b11 6
#104550000000
1!
1%
1-
12
15
#104560000000
0!
0%
b100 *
0-
02
b100 6
#104570000000
1!
1%
1-
12
#104580000000
0!
0%
b101 *
0-
02
b101 6
#104590000000
1!
1%
1-
12
#104600000000
0!
0%
b110 *
0-
02
b110 6
#104610000000
1!
1%
1-
12
#104620000000
0!
0%
b111 *
0-
02
b111 6
#104630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#104640000000
0!
0%
b0 *
0-
02
b0 6
#104650000000
1!
1%
1-
12
#104660000000
0!
0%
b1 *
0-
02
b1 6
#104670000000
1!
1%
1-
12
#104680000000
0!
0%
b10 *
0-
02
b10 6
#104690000000
1!
1%
1-
12
#104700000000
0!
0%
b11 *
0-
02
b11 6
#104710000000
1!
1%
1-
12
15
#104720000000
0!
0%
b100 *
0-
02
b100 6
#104730000000
1!
1%
1-
12
#104740000000
0!
0%
b101 *
0-
02
b101 6
#104750000000
1!
1%
1-
12
#104760000000
0!
0%
b110 *
0-
02
b110 6
#104770000000
1!
1%
1-
12
#104780000000
0!
0%
b111 *
0-
02
b111 6
#104790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#104800000000
0!
0%
b0 *
0-
02
b0 6
#104810000000
1!
1%
1-
12
#104820000000
0!
0%
b1 *
0-
02
b1 6
#104830000000
1!
1%
1-
12
#104840000000
0!
0%
b10 *
0-
02
b10 6
#104850000000
1!
1%
1-
12
#104860000000
0!
0%
b11 *
0-
02
b11 6
#104870000000
1!
1%
1-
12
15
#104880000000
0!
0%
b100 *
0-
02
b100 6
#104890000000
1!
1%
1-
12
#104900000000
0!
0%
b101 *
0-
02
b101 6
#104910000000
1!
1%
1-
12
#104920000000
0!
0%
b110 *
0-
02
b110 6
#104930000000
1!
1%
1-
12
#104940000000
0!
0%
b111 *
0-
02
b111 6
#104950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#104960000000
0!
0%
b0 *
0-
02
b0 6
#104970000000
1!
1%
1-
12
#104980000000
0!
0%
b1 *
0-
02
b1 6
#104990000000
1!
1%
1-
12
#105000000000
0!
0%
b10 *
0-
02
b10 6
#105010000000
1!
1%
1-
12
#105020000000
0!
0%
b11 *
0-
02
b11 6
#105030000000
1!
1%
1-
12
15
#105040000000
0!
0%
b100 *
0-
02
b100 6
#105050000000
1!
1%
1-
12
#105060000000
0!
0%
b101 *
0-
02
b101 6
#105070000000
1!
1%
1-
12
#105080000000
0!
0%
b110 *
0-
02
b110 6
#105090000000
1!
1%
1-
12
#105100000000
0!
0%
b111 *
0-
02
b111 6
#105110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#105120000000
0!
0%
b0 *
0-
02
b0 6
#105130000000
1!
1%
1-
12
#105140000000
0!
0%
b1 *
0-
02
b1 6
#105150000000
1!
1%
1-
12
#105160000000
0!
0%
b10 *
0-
02
b10 6
#105170000000
1!
1%
1-
12
#105180000000
0!
0%
b11 *
0-
02
b11 6
#105190000000
1!
1%
1-
12
15
#105200000000
0!
0%
b100 *
0-
02
b100 6
#105210000000
1!
1%
1-
12
#105220000000
0!
0%
b101 *
0-
02
b101 6
#105230000000
1!
1%
1-
12
#105240000000
0!
0%
b110 *
0-
02
b110 6
#105250000000
1!
1%
1-
12
#105260000000
0!
0%
b111 *
0-
02
b111 6
#105270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#105280000000
0!
0%
b0 *
0-
02
b0 6
#105290000000
1!
1%
1-
12
#105300000000
0!
0%
b1 *
0-
02
b1 6
#105310000000
1!
1%
1-
12
#105320000000
0!
0%
b10 *
0-
02
b10 6
#105330000000
1!
1%
1-
12
#105340000000
0!
0%
b11 *
0-
02
b11 6
#105350000000
1!
1%
1-
12
15
#105360000000
0!
0%
b100 *
0-
02
b100 6
#105370000000
1!
1%
1-
12
#105380000000
0!
0%
b101 *
0-
02
b101 6
#105390000000
1!
1%
1-
12
#105400000000
0!
0%
b110 *
0-
02
b110 6
#105410000000
1!
1%
1-
12
#105420000000
0!
0%
b111 *
0-
02
b111 6
#105430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#105440000000
0!
0%
b0 *
0-
02
b0 6
#105450000000
1!
1%
1-
12
#105460000000
0!
0%
b1 *
0-
02
b1 6
#105470000000
1!
1%
1-
12
#105480000000
0!
0%
b10 *
0-
02
b10 6
#105490000000
1!
1%
1-
12
#105500000000
0!
0%
b11 *
0-
02
b11 6
#105510000000
1!
1%
1-
12
15
#105520000000
0!
0%
b100 *
0-
02
b100 6
#105530000000
1!
1%
1-
12
#105540000000
0!
0%
b101 *
0-
02
b101 6
#105550000000
1!
1%
1-
12
#105560000000
0!
0%
b110 *
0-
02
b110 6
#105570000000
1!
1%
1-
12
#105580000000
0!
0%
b111 *
0-
02
b111 6
#105590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#105600000000
0!
0%
b0 *
0-
02
b0 6
#105610000000
1!
1%
1-
12
#105620000000
0!
0%
b1 *
0-
02
b1 6
#105630000000
1!
1%
1-
12
#105640000000
0!
0%
b10 *
0-
02
b10 6
#105650000000
1!
1%
1-
12
#105660000000
0!
0%
b11 *
0-
02
b11 6
#105670000000
1!
1%
1-
12
15
#105680000000
0!
0%
b100 *
0-
02
b100 6
#105690000000
1!
1%
1-
12
#105700000000
0!
0%
b101 *
0-
02
b101 6
#105710000000
1!
1%
1-
12
#105720000000
0!
0%
b110 *
0-
02
b110 6
#105730000000
1!
1%
1-
12
#105740000000
0!
0%
b111 *
0-
02
b111 6
#105750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#105760000000
0!
0%
b0 *
0-
02
b0 6
#105770000000
1!
1%
1-
12
#105780000000
0!
0%
b1 *
0-
02
b1 6
#105790000000
1!
1%
1-
12
#105800000000
0!
0%
b10 *
0-
02
b10 6
#105810000000
1!
1%
1-
12
#105820000000
0!
0%
b11 *
0-
02
b11 6
#105830000000
1!
1%
1-
12
15
#105840000000
0!
0%
b100 *
0-
02
b100 6
#105850000000
1!
1%
1-
12
#105860000000
0!
0%
b101 *
0-
02
b101 6
#105870000000
1!
1%
1-
12
#105880000000
0!
0%
b110 *
0-
02
b110 6
#105890000000
1!
1%
1-
12
#105900000000
0!
0%
b111 *
0-
02
b111 6
#105910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#105920000000
0!
0%
b0 *
0-
02
b0 6
#105930000000
1!
1%
1-
12
#105940000000
0!
0%
b1 *
0-
02
b1 6
#105950000000
1!
1%
1-
12
#105960000000
0!
0%
b10 *
0-
02
b10 6
#105970000000
1!
1%
1-
12
#105980000000
0!
0%
b11 *
0-
02
b11 6
#105990000000
1!
1%
1-
12
15
#106000000000
0!
0%
b100 *
0-
02
b100 6
#106010000000
1!
1%
1-
12
#106020000000
0!
0%
b101 *
0-
02
b101 6
#106030000000
1!
1%
1-
12
#106040000000
0!
0%
b110 *
0-
02
b110 6
#106050000000
1!
1%
1-
12
#106060000000
0!
0%
b111 *
0-
02
b111 6
#106070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#106080000000
0!
0%
b0 *
0-
02
b0 6
#106090000000
1!
1%
1-
12
#106100000000
0!
0%
b1 *
0-
02
b1 6
#106110000000
1!
1%
1-
12
#106120000000
0!
0%
b10 *
0-
02
b10 6
#106130000000
1!
1%
1-
12
#106140000000
0!
0%
b11 *
0-
02
b11 6
#106150000000
1!
1%
1-
12
15
#106160000000
0!
0%
b100 *
0-
02
b100 6
#106170000000
1!
1%
1-
12
#106180000000
0!
0%
b101 *
0-
02
b101 6
#106190000000
1!
1%
1-
12
#106200000000
0!
0%
b110 *
0-
02
b110 6
#106210000000
1!
1%
1-
12
#106220000000
0!
0%
b111 *
0-
02
b111 6
#106230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#106240000000
0!
0%
b0 *
0-
02
b0 6
#106250000000
1!
1%
1-
12
#106260000000
0!
0%
b1 *
0-
02
b1 6
#106270000000
1!
1%
1-
12
#106280000000
0!
0%
b10 *
0-
02
b10 6
#106290000000
1!
1%
1-
12
#106300000000
0!
0%
b11 *
0-
02
b11 6
#106310000000
1!
1%
1-
12
15
#106320000000
0!
0%
b100 *
0-
02
b100 6
#106330000000
1!
1%
1-
12
#106340000000
0!
0%
b101 *
0-
02
b101 6
#106350000000
1!
1%
1-
12
#106360000000
0!
0%
b110 *
0-
02
b110 6
#106370000000
1!
1%
1-
12
#106380000000
0!
0%
b111 *
0-
02
b111 6
#106390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#106400000000
0!
0%
b0 *
0-
02
b0 6
#106410000000
1!
1%
1-
12
#106420000000
0!
0%
b1 *
0-
02
b1 6
#106430000000
1!
1%
1-
12
#106440000000
0!
0%
b10 *
0-
02
b10 6
#106450000000
1!
1%
1-
12
#106460000000
0!
0%
b11 *
0-
02
b11 6
#106470000000
1!
1%
1-
12
15
#106480000000
0!
0%
b100 *
0-
02
b100 6
#106490000000
1!
1%
1-
12
#106500000000
0!
0%
b101 *
0-
02
b101 6
#106510000000
1!
1%
1-
12
#106520000000
0!
0%
b110 *
0-
02
b110 6
#106530000000
1!
1%
1-
12
#106540000000
0!
0%
b111 *
0-
02
b111 6
#106550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#106560000000
0!
0%
b0 *
0-
02
b0 6
#106570000000
1!
1%
1-
12
#106580000000
0!
0%
b1 *
0-
02
b1 6
#106590000000
1!
1%
1-
12
#106600000000
0!
0%
b10 *
0-
02
b10 6
#106610000000
1!
1%
1-
12
#106620000000
0!
0%
b11 *
0-
02
b11 6
#106630000000
1!
1%
1-
12
15
#106640000000
0!
0%
b100 *
0-
02
b100 6
#106650000000
1!
1%
1-
12
#106660000000
0!
0%
b101 *
0-
02
b101 6
#106670000000
1!
1%
1-
12
#106680000000
0!
0%
b110 *
0-
02
b110 6
#106690000000
1!
1%
1-
12
#106700000000
0!
0%
b111 *
0-
02
b111 6
#106710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#106720000000
0!
0%
b0 *
0-
02
b0 6
#106730000000
1!
1%
1-
12
#106740000000
0!
0%
b1 *
0-
02
b1 6
#106750000000
1!
1%
1-
12
#106760000000
0!
0%
b10 *
0-
02
b10 6
#106770000000
1!
1%
1-
12
#106780000000
0!
0%
b11 *
0-
02
b11 6
#106790000000
1!
1%
1-
12
15
#106800000000
0!
0%
b100 *
0-
02
b100 6
#106810000000
1!
1%
1-
12
#106820000000
0!
0%
b101 *
0-
02
b101 6
#106830000000
1!
1%
1-
12
#106840000000
0!
0%
b110 *
0-
02
b110 6
#106850000000
1!
1%
1-
12
#106860000000
0!
0%
b111 *
0-
02
b111 6
#106870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#106880000000
0!
0%
b0 *
0-
02
b0 6
#106890000000
1!
1%
1-
12
#106900000000
0!
0%
b1 *
0-
02
b1 6
#106910000000
1!
1%
1-
12
#106920000000
0!
0%
b10 *
0-
02
b10 6
#106930000000
1!
1%
1-
12
#106940000000
0!
0%
b11 *
0-
02
b11 6
#106950000000
1!
1%
1-
12
15
#106960000000
0!
0%
b100 *
0-
02
b100 6
#106970000000
1!
1%
1-
12
#106980000000
0!
0%
b101 *
0-
02
b101 6
#106990000000
1!
1%
1-
12
#107000000000
0!
0%
b110 *
0-
02
b110 6
#107010000000
1!
1%
1-
12
#107020000000
0!
0%
b111 *
0-
02
b111 6
#107030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#107040000000
0!
0%
b0 *
0-
02
b0 6
#107050000000
1!
1%
1-
12
#107060000000
0!
0%
b1 *
0-
02
b1 6
#107070000000
1!
1%
1-
12
#107080000000
0!
0%
b10 *
0-
02
b10 6
#107090000000
1!
1%
1-
12
#107100000000
0!
0%
b11 *
0-
02
b11 6
#107110000000
1!
1%
1-
12
15
#107120000000
0!
0%
b100 *
0-
02
b100 6
#107130000000
1!
1%
1-
12
#107140000000
0!
0%
b101 *
0-
02
b101 6
#107150000000
1!
1%
1-
12
#107160000000
0!
0%
b110 *
0-
02
b110 6
#107170000000
1!
1%
1-
12
#107180000000
0!
0%
b111 *
0-
02
b111 6
#107190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#107200000000
0!
0%
b0 *
0-
02
b0 6
#107210000000
1!
1%
1-
12
#107220000000
0!
0%
b1 *
0-
02
b1 6
#107230000000
1!
1%
1-
12
#107240000000
0!
0%
b10 *
0-
02
b10 6
#107250000000
1!
1%
1-
12
#107260000000
0!
0%
b11 *
0-
02
b11 6
#107270000000
1!
1%
1-
12
15
#107280000000
0!
0%
b100 *
0-
02
b100 6
#107290000000
1!
1%
1-
12
#107300000000
0!
0%
b101 *
0-
02
b101 6
#107310000000
1!
1%
1-
12
#107320000000
0!
0%
b110 *
0-
02
b110 6
#107330000000
1!
1%
1-
12
#107340000000
0!
0%
b111 *
0-
02
b111 6
#107350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#107360000000
0!
0%
b0 *
0-
02
b0 6
#107370000000
1!
1%
1-
12
#107380000000
0!
0%
b1 *
0-
02
b1 6
#107390000000
1!
1%
1-
12
#107400000000
0!
0%
b10 *
0-
02
b10 6
#107410000000
1!
1%
1-
12
#107420000000
0!
0%
b11 *
0-
02
b11 6
#107430000000
1!
1%
1-
12
15
#107440000000
0!
0%
b100 *
0-
02
b100 6
#107450000000
1!
1%
1-
12
#107460000000
0!
0%
b101 *
0-
02
b101 6
#107470000000
1!
1%
1-
12
#107480000000
0!
0%
b110 *
0-
02
b110 6
#107490000000
1!
1%
1-
12
#107500000000
0!
0%
b111 *
0-
02
b111 6
#107510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#107520000000
0!
0%
b0 *
0-
02
b0 6
#107530000000
1!
1%
1-
12
#107540000000
0!
0%
b1 *
0-
02
b1 6
#107550000000
1!
1%
1-
12
#107560000000
0!
0%
b10 *
0-
02
b10 6
#107570000000
1!
1%
1-
12
#107580000000
0!
0%
b11 *
0-
02
b11 6
#107590000000
1!
1%
1-
12
15
#107600000000
0!
0%
b100 *
0-
02
b100 6
#107610000000
1!
1%
1-
12
#107620000000
0!
0%
b101 *
0-
02
b101 6
#107630000000
1!
1%
1-
12
#107640000000
0!
0%
b110 *
0-
02
b110 6
#107650000000
1!
1%
1-
12
#107660000000
0!
0%
b111 *
0-
02
b111 6
#107670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#107680000000
0!
0%
b0 *
0-
02
b0 6
#107690000000
1!
1%
1-
12
#107700000000
0!
0%
b1 *
0-
02
b1 6
#107710000000
1!
1%
1-
12
#107720000000
0!
0%
b10 *
0-
02
b10 6
#107730000000
1!
1%
1-
12
#107740000000
0!
0%
b11 *
0-
02
b11 6
#107750000000
1!
1%
1-
12
15
#107760000000
0!
0%
b100 *
0-
02
b100 6
#107770000000
1!
1%
1-
12
#107780000000
0!
0%
b101 *
0-
02
b101 6
#107790000000
1!
1%
1-
12
#107800000000
0!
0%
b110 *
0-
02
b110 6
#107810000000
1!
1%
1-
12
#107820000000
0!
0%
b111 *
0-
02
b111 6
#107830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#107840000000
0!
0%
b0 *
0-
02
b0 6
#107850000000
1!
1%
1-
12
#107860000000
0!
0%
b1 *
0-
02
b1 6
#107870000000
1!
1%
1-
12
#107880000000
0!
0%
b10 *
0-
02
b10 6
#107890000000
1!
1%
1-
12
#107900000000
0!
0%
b11 *
0-
02
b11 6
#107910000000
1!
1%
1-
12
15
#107920000000
0!
0%
b100 *
0-
02
b100 6
#107930000000
1!
1%
1-
12
#107940000000
0!
0%
b101 *
0-
02
b101 6
#107950000000
1!
1%
1-
12
#107960000000
0!
0%
b110 *
0-
02
b110 6
#107970000000
1!
1%
1-
12
#107980000000
0!
0%
b111 *
0-
02
b111 6
#107990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#108000000000
0!
0%
b0 *
0-
02
b0 6
#108010000000
1!
1%
1-
12
#108020000000
0!
0%
b1 *
0-
02
b1 6
#108030000000
1!
1%
1-
12
#108040000000
0!
0%
b10 *
0-
02
b10 6
#108050000000
1!
1%
1-
12
#108060000000
0!
0%
b11 *
0-
02
b11 6
#108070000000
1!
1%
1-
12
15
#108080000000
0!
0%
b100 *
0-
02
b100 6
#108090000000
1!
1%
1-
12
#108100000000
0!
0%
b101 *
0-
02
b101 6
#108110000000
1!
1%
1-
12
#108120000000
0!
0%
b110 *
0-
02
b110 6
#108130000000
1!
1%
1-
12
#108140000000
0!
0%
b111 *
0-
02
b111 6
#108150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#108160000000
0!
0%
b0 *
0-
02
b0 6
#108170000000
1!
1%
1-
12
#108180000000
0!
0%
b1 *
0-
02
b1 6
#108190000000
1!
1%
1-
12
#108200000000
0!
0%
b10 *
0-
02
b10 6
#108210000000
1!
1%
1-
12
#108220000000
0!
0%
b11 *
0-
02
b11 6
#108230000000
1!
1%
1-
12
15
#108240000000
0!
0%
b100 *
0-
02
b100 6
#108250000000
1!
1%
1-
12
#108260000000
0!
0%
b101 *
0-
02
b101 6
#108270000000
1!
1%
1-
12
#108280000000
0!
0%
b110 *
0-
02
b110 6
#108290000000
1!
1%
1-
12
#108300000000
0!
0%
b111 *
0-
02
b111 6
#108310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#108320000000
0!
0%
b0 *
0-
02
b0 6
#108330000000
1!
1%
1-
12
#108340000000
0!
0%
b1 *
0-
02
b1 6
#108350000000
1!
1%
1-
12
#108360000000
0!
0%
b10 *
0-
02
b10 6
#108370000000
1!
1%
1-
12
#108380000000
0!
0%
b11 *
0-
02
b11 6
#108390000000
1!
1%
1-
12
15
#108400000000
0!
0%
b100 *
0-
02
b100 6
#108410000000
1!
1%
1-
12
#108420000000
0!
0%
b101 *
0-
02
b101 6
#108430000000
1!
1%
1-
12
#108440000000
0!
0%
b110 *
0-
02
b110 6
#108450000000
1!
1%
1-
12
#108460000000
0!
0%
b111 *
0-
02
b111 6
#108470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#108480000000
0!
0%
b0 *
0-
02
b0 6
#108490000000
1!
1%
1-
12
#108500000000
0!
0%
b1 *
0-
02
b1 6
#108510000000
1!
1%
1-
12
#108520000000
0!
0%
b10 *
0-
02
b10 6
#108530000000
1!
1%
1-
12
#108540000000
0!
0%
b11 *
0-
02
b11 6
#108550000000
1!
1%
1-
12
15
#108560000000
0!
0%
b100 *
0-
02
b100 6
#108570000000
1!
1%
1-
12
#108580000000
0!
0%
b101 *
0-
02
b101 6
#108590000000
1!
1%
1-
12
#108600000000
0!
0%
b110 *
0-
02
b110 6
#108610000000
1!
1%
1-
12
#108620000000
0!
0%
b111 *
0-
02
b111 6
#108630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#108640000000
0!
0%
b0 *
0-
02
b0 6
#108650000000
1!
1%
1-
12
#108660000000
0!
0%
b1 *
0-
02
b1 6
#108670000000
1!
1%
1-
12
#108680000000
0!
0%
b10 *
0-
02
b10 6
#108690000000
1!
1%
1-
12
#108700000000
0!
0%
b11 *
0-
02
b11 6
#108710000000
1!
1%
1-
12
15
#108720000000
0!
0%
b100 *
0-
02
b100 6
#108730000000
1!
1%
1-
12
#108740000000
0!
0%
b101 *
0-
02
b101 6
#108750000000
1!
1%
1-
12
#108760000000
0!
0%
b110 *
0-
02
b110 6
#108770000000
1!
1%
1-
12
#108780000000
0!
0%
b111 *
0-
02
b111 6
#108790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#108800000000
0!
0%
b0 *
0-
02
b0 6
#108810000000
1!
1%
1-
12
#108820000000
0!
0%
b1 *
0-
02
b1 6
#108830000000
1!
1%
1-
12
#108840000000
0!
0%
b10 *
0-
02
b10 6
#108850000000
1!
1%
1-
12
#108860000000
0!
0%
b11 *
0-
02
b11 6
#108870000000
1!
1%
1-
12
15
#108880000000
0!
0%
b100 *
0-
02
b100 6
#108890000000
1!
1%
1-
12
#108900000000
0!
0%
b101 *
0-
02
b101 6
#108910000000
1!
1%
1-
12
#108920000000
0!
0%
b110 *
0-
02
b110 6
#108930000000
1!
1%
1-
12
#108940000000
0!
0%
b111 *
0-
02
b111 6
#108950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#108960000000
0!
0%
b0 *
0-
02
b0 6
#108970000000
1!
1%
1-
12
#108980000000
0!
0%
b1 *
0-
02
b1 6
#108990000000
1!
1%
1-
12
#109000000000
0!
0%
b10 *
0-
02
b10 6
#109010000000
1!
1%
1-
12
#109020000000
0!
0%
b11 *
0-
02
b11 6
#109030000000
1!
1%
1-
12
15
#109040000000
0!
0%
b100 *
0-
02
b100 6
#109050000000
1!
1%
1-
12
#109060000000
0!
0%
b101 *
0-
02
b101 6
#109070000000
1!
1%
1-
12
#109080000000
0!
0%
b110 *
0-
02
b110 6
#109090000000
1!
1%
1-
12
#109100000000
0!
0%
b111 *
0-
02
b111 6
#109110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#109120000000
0!
0%
b0 *
0-
02
b0 6
#109130000000
1!
1%
1-
12
#109140000000
0!
0%
b1 *
0-
02
b1 6
#109150000000
1!
1%
1-
12
#109160000000
0!
0%
b10 *
0-
02
b10 6
#109170000000
1!
1%
1-
12
#109180000000
0!
0%
b11 *
0-
02
b11 6
#109190000000
1!
1%
1-
12
15
#109200000000
0!
0%
b100 *
0-
02
b100 6
#109210000000
1!
1%
1-
12
#109220000000
0!
0%
b101 *
0-
02
b101 6
#109230000000
1!
1%
1-
12
#109240000000
0!
0%
b110 *
0-
02
b110 6
#109250000000
1!
1%
1-
12
#109260000000
0!
0%
b111 *
0-
02
b111 6
#109270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#109280000000
0!
0%
b0 *
0-
02
b0 6
#109290000000
1!
1%
1-
12
#109300000000
0!
0%
b1 *
0-
02
b1 6
#109310000000
1!
1%
1-
12
#109320000000
0!
0%
b10 *
0-
02
b10 6
#109330000000
1!
1%
1-
12
#109340000000
0!
0%
b11 *
0-
02
b11 6
#109350000000
1!
1%
1-
12
15
#109360000000
0!
0%
b100 *
0-
02
b100 6
#109370000000
1!
1%
1-
12
#109380000000
0!
0%
b101 *
0-
02
b101 6
#109390000000
1!
1%
1-
12
#109400000000
0!
0%
b110 *
0-
02
b110 6
#109410000000
1!
1%
1-
12
#109420000000
0!
0%
b111 *
0-
02
b111 6
#109430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#109440000000
0!
0%
b0 *
0-
02
b0 6
#109450000000
1!
1%
1-
12
#109460000000
0!
0%
b1 *
0-
02
b1 6
#109470000000
1!
1%
1-
12
#109480000000
0!
0%
b10 *
0-
02
b10 6
#109490000000
1!
1%
1-
12
#109500000000
0!
0%
b11 *
0-
02
b11 6
#109510000000
1!
1%
1-
12
15
#109520000000
0!
0%
b100 *
0-
02
b100 6
#109530000000
1!
1%
1-
12
#109540000000
0!
0%
b101 *
0-
02
b101 6
#109550000000
1!
1%
1-
12
#109560000000
0!
0%
b110 *
0-
02
b110 6
#109570000000
1!
1%
1-
12
#109580000000
0!
0%
b111 *
0-
02
b111 6
#109590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#109600000000
0!
0%
b0 *
0-
02
b0 6
#109610000000
1!
1%
1-
12
#109620000000
0!
0%
b1 *
0-
02
b1 6
#109630000000
1!
1%
1-
12
#109640000000
0!
0%
b10 *
0-
02
b10 6
#109650000000
1!
1%
1-
12
#109660000000
0!
0%
b11 *
0-
02
b11 6
#109670000000
1!
1%
1-
12
15
#109680000000
0!
0%
b100 *
0-
02
b100 6
#109690000000
1!
1%
1-
12
#109700000000
0!
0%
b101 *
0-
02
b101 6
#109710000000
1!
1%
1-
12
#109720000000
0!
0%
b110 *
0-
02
b110 6
#109730000000
1!
1%
1-
12
#109740000000
0!
0%
b111 *
0-
02
b111 6
#109750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#109760000000
0!
0%
b0 *
0-
02
b0 6
#109770000000
1!
1%
1-
12
#109780000000
0!
0%
b1 *
0-
02
b1 6
#109790000000
1!
1%
1-
12
#109800000000
0!
0%
b10 *
0-
02
b10 6
#109810000000
1!
1%
1-
12
#109820000000
0!
0%
b11 *
0-
02
b11 6
#109830000000
1!
1%
1-
12
15
#109840000000
0!
0%
b100 *
0-
02
b100 6
#109850000000
1!
1%
1-
12
#109860000000
0!
0%
b101 *
0-
02
b101 6
#109870000000
1!
1%
1-
12
#109880000000
0!
0%
b110 *
0-
02
b110 6
#109890000000
1!
1%
1-
12
#109900000000
0!
0%
b111 *
0-
02
b111 6
#109910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#109920000000
0!
0%
b0 *
0-
02
b0 6
#109930000000
1!
1%
1-
12
#109940000000
0!
0%
b1 *
0-
02
b1 6
#109950000000
1!
1%
1-
12
#109960000000
0!
0%
b10 *
0-
02
b10 6
#109970000000
1!
1%
1-
12
#109980000000
0!
0%
b11 *
0-
02
b11 6
#109990000000
1!
1%
1-
12
15
#110000000000
0!
0%
b100 *
0-
02
b100 6
#110010000000
1!
1%
1-
12
#110020000000
0!
0%
b101 *
0-
02
b101 6
#110030000000
1!
1%
1-
12
#110040000000
0!
0%
b110 *
0-
02
b110 6
#110050000000
1!
1%
1-
12
#110060000000
0!
0%
b111 *
0-
02
b111 6
#110070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#110080000000
0!
0%
b0 *
0-
02
b0 6
#110090000000
1!
1%
1-
12
#110100000000
0!
0%
b1 *
0-
02
b1 6
#110110000000
1!
1%
1-
12
#110120000000
0!
0%
b10 *
0-
02
b10 6
#110130000000
1!
1%
1-
12
#110140000000
0!
0%
b11 *
0-
02
b11 6
#110150000000
1!
1%
1-
12
15
#110160000000
0!
0%
b100 *
0-
02
b100 6
#110170000000
1!
1%
1-
12
#110180000000
0!
0%
b101 *
0-
02
b101 6
#110190000000
1!
1%
1-
12
#110200000000
0!
0%
b110 *
0-
02
b110 6
#110210000000
1!
1%
1-
12
#110220000000
0!
0%
b111 *
0-
02
b111 6
#110230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#110240000000
0!
0%
b0 *
0-
02
b0 6
#110250000000
1!
1%
1-
12
#110260000000
0!
0%
b1 *
0-
02
b1 6
#110270000000
1!
1%
1-
12
#110280000000
0!
0%
b10 *
0-
02
b10 6
#110290000000
1!
1%
1-
12
#110300000000
0!
0%
b11 *
0-
02
b11 6
#110310000000
1!
1%
1-
12
15
#110320000000
0!
0%
b100 *
0-
02
b100 6
#110330000000
1!
1%
1-
12
#110340000000
0!
0%
b101 *
0-
02
b101 6
#110350000000
1!
1%
1-
12
#110360000000
0!
0%
b110 *
0-
02
b110 6
#110370000000
1!
1%
1-
12
#110380000000
0!
0%
b111 *
0-
02
b111 6
#110390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#110400000000
0!
0%
b0 *
0-
02
b0 6
#110410000000
1!
1%
1-
12
#110420000000
0!
0%
b1 *
0-
02
b1 6
#110430000000
1!
1%
1-
12
#110440000000
0!
0%
b10 *
0-
02
b10 6
#110450000000
1!
1%
1-
12
#110460000000
0!
0%
b11 *
0-
02
b11 6
#110470000000
1!
1%
1-
12
15
#110480000000
0!
0%
b100 *
0-
02
b100 6
#110490000000
1!
1%
1-
12
#110500000000
0!
0%
b101 *
0-
02
b101 6
#110510000000
1!
1%
1-
12
#110520000000
0!
0%
b110 *
0-
02
b110 6
#110530000000
1!
1%
1-
12
#110540000000
0!
0%
b111 *
0-
02
b111 6
#110550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#110560000000
0!
0%
b0 *
0-
02
b0 6
#110570000000
1!
1%
1-
12
#110580000000
0!
0%
b1 *
0-
02
b1 6
#110590000000
1!
1%
1-
12
#110600000000
0!
0%
b10 *
0-
02
b10 6
#110610000000
1!
1%
1-
12
#110620000000
0!
0%
b11 *
0-
02
b11 6
#110630000000
1!
1%
1-
12
15
#110640000000
0!
0%
b100 *
0-
02
b100 6
#110650000000
1!
1%
1-
12
#110660000000
0!
0%
b101 *
0-
02
b101 6
#110670000000
1!
1%
1-
12
#110680000000
0!
0%
b110 *
0-
02
b110 6
#110690000000
1!
1%
1-
12
#110700000000
0!
0%
b111 *
0-
02
b111 6
#110710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#110720000000
0!
0%
b0 *
0-
02
b0 6
#110730000000
1!
1%
1-
12
#110740000000
0!
0%
b1 *
0-
02
b1 6
#110750000000
1!
1%
1-
12
#110760000000
0!
0%
b10 *
0-
02
b10 6
#110770000000
1!
1%
1-
12
#110780000000
0!
0%
b11 *
0-
02
b11 6
#110790000000
1!
1%
1-
12
15
#110800000000
0!
0%
b100 *
0-
02
b100 6
#110810000000
1!
1%
1-
12
#110820000000
0!
0%
b101 *
0-
02
b101 6
#110830000000
1!
1%
1-
12
#110840000000
0!
0%
b110 *
0-
02
b110 6
#110850000000
1!
1%
1-
12
#110860000000
0!
0%
b111 *
0-
02
b111 6
#110870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#110880000000
0!
0%
b0 *
0-
02
b0 6
#110890000000
1!
1%
1-
12
#110900000000
0!
0%
b1 *
0-
02
b1 6
#110910000000
1!
1%
1-
12
#110920000000
0!
0%
b10 *
0-
02
b10 6
#110930000000
1!
1%
1-
12
#110940000000
0!
0%
b11 *
0-
02
b11 6
#110950000000
1!
1%
1-
12
15
#110960000000
0!
0%
b100 *
0-
02
b100 6
#110970000000
1!
1%
1-
12
#110980000000
0!
0%
b101 *
0-
02
b101 6
#110990000000
1!
1%
1-
12
#111000000000
0!
0%
b110 *
0-
02
b110 6
#111010000000
1!
1%
1-
12
#111020000000
0!
0%
b111 *
0-
02
b111 6
#111030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#111040000000
0!
0%
b0 *
0-
02
b0 6
#111050000000
1!
1%
1-
12
#111060000000
0!
0%
b1 *
0-
02
b1 6
#111070000000
1!
1%
1-
12
#111080000000
0!
0%
b10 *
0-
02
b10 6
#111090000000
1!
1%
1-
12
#111100000000
0!
0%
b11 *
0-
02
b11 6
#111110000000
1!
1%
1-
12
15
#111120000000
0!
0%
b100 *
0-
02
b100 6
#111130000000
1!
1%
1-
12
#111140000000
0!
0%
b101 *
0-
02
b101 6
#111150000000
1!
1%
1-
12
#111160000000
0!
0%
b110 *
0-
02
b110 6
#111170000000
1!
1%
1-
12
#111180000000
0!
0%
b111 *
0-
02
b111 6
#111190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#111200000000
0!
0%
b0 *
0-
02
b0 6
#111210000000
1!
1%
1-
12
#111220000000
0!
0%
b1 *
0-
02
b1 6
#111230000000
1!
1%
1-
12
#111240000000
0!
0%
b10 *
0-
02
b10 6
#111250000000
1!
1%
1-
12
#111260000000
0!
0%
b11 *
0-
02
b11 6
#111270000000
1!
1%
1-
12
15
#111280000000
0!
0%
b100 *
0-
02
b100 6
#111290000000
1!
1%
1-
12
#111300000000
0!
0%
b101 *
0-
02
b101 6
#111310000000
1!
1%
1-
12
#111320000000
0!
0%
b110 *
0-
02
b110 6
#111330000000
1!
1%
1-
12
#111340000000
0!
0%
b111 *
0-
02
b111 6
#111350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#111360000000
0!
0%
b0 *
0-
02
b0 6
#111370000000
1!
1%
1-
12
#111380000000
0!
0%
b1 *
0-
02
b1 6
#111390000000
1!
1%
1-
12
#111400000000
0!
0%
b10 *
0-
02
b10 6
#111410000000
1!
1%
1-
12
#111420000000
0!
0%
b11 *
0-
02
b11 6
#111430000000
1!
1%
1-
12
15
#111440000000
0!
0%
b100 *
0-
02
b100 6
#111450000000
1!
1%
1-
12
#111460000000
0!
0%
b101 *
0-
02
b101 6
#111470000000
1!
1%
1-
12
#111480000000
0!
0%
b110 *
0-
02
b110 6
#111490000000
1!
1%
1-
12
#111500000000
0!
0%
b111 *
0-
02
b111 6
#111510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#111520000000
0!
0%
b0 *
0-
02
b0 6
#111530000000
1!
1%
1-
12
#111540000000
0!
0%
b1 *
0-
02
b1 6
#111550000000
1!
1%
1-
12
#111560000000
0!
0%
b10 *
0-
02
b10 6
#111570000000
1!
1%
1-
12
#111580000000
0!
0%
b11 *
0-
02
b11 6
#111590000000
1!
1%
1-
12
15
#111600000000
0!
0%
b100 *
0-
02
b100 6
#111610000000
1!
1%
1-
12
#111620000000
0!
0%
b101 *
0-
02
b101 6
#111630000000
1!
1%
1-
12
#111640000000
0!
0%
b110 *
0-
02
b110 6
#111650000000
1!
1%
1-
12
#111660000000
0!
0%
b111 *
0-
02
b111 6
#111670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#111680000000
0!
0%
b0 *
0-
02
b0 6
#111690000000
1!
1%
1-
12
#111700000000
0!
0%
b1 *
0-
02
b1 6
#111710000000
1!
1%
1-
12
#111720000000
0!
0%
b10 *
0-
02
b10 6
#111730000000
1!
1%
1-
12
#111740000000
0!
0%
b11 *
0-
02
b11 6
#111750000000
1!
1%
1-
12
15
#111760000000
0!
0%
b100 *
0-
02
b100 6
#111770000000
1!
1%
1-
12
#111780000000
0!
0%
b101 *
0-
02
b101 6
#111790000000
1!
1%
1-
12
#111800000000
0!
0%
b110 *
0-
02
b110 6
#111810000000
1!
1%
1-
12
#111820000000
0!
0%
b111 *
0-
02
b111 6
#111830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#111840000000
0!
0%
b0 *
0-
02
b0 6
#111850000000
1!
1%
1-
12
#111860000000
0!
0%
b1 *
0-
02
b1 6
#111870000000
1!
1%
1-
12
#111880000000
0!
0%
b10 *
0-
02
b10 6
#111890000000
1!
1%
1-
12
#111900000000
0!
0%
b11 *
0-
02
b11 6
#111910000000
1!
1%
1-
12
15
#111920000000
0!
0%
b100 *
0-
02
b100 6
#111930000000
1!
1%
1-
12
#111940000000
0!
0%
b101 *
0-
02
b101 6
#111950000000
1!
1%
1-
12
#111960000000
0!
0%
b110 *
0-
02
b110 6
#111970000000
1!
1%
1-
12
#111980000000
0!
0%
b111 *
0-
02
b111 6
#111990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#112000000000
0!
0%
b0 *
0-
02
b0 6
#112010000000
1!
1%
1-
12
#112020000000
0!
0%
b1 *
0-
02
b1 6
#112030000000
1!
1%
1-
12
#112040000000
0!
0%
b10 *
0-
02
b10 6
#112050000000
1!
1%
1-
12
#112060000000
0!
0%
b11 *
0-
02
b11 6
#112070000000
1!
1%
1-
12
15
#112080000000
0!
0%
b100 *
0-
02
b100 6
#112090000000
1!
1%
1-
12
#112100000000
0!
0%
b101 *
0-
02
b101 6
#112110000000
1!
1%
1-
12
#112120000000
0!
0%
b110 *
0-
02
b110 6
#112130000000
1!
1%
1-
12
#112140000000
0!
0%
b111 *
0-
02
b111 6
#112150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#112160000000
0!
0%
b0 *
0-
02
b0 6
#112170000000
1!
1%
1-
12
#112180000000
0!
0%
b1 *
0-
02
b1 6
#112190000000
1!
1%
1-
12
#112200000000
0!
0%
b10 *
0-
02
b10 6
#112210000000
1!
1%
1-
12
#112220000000
0!
0%
b11 *
0-
02
b11 6
#112230000000
1!
1%
1-
12
15
#112240000000
0!
0%
b100 *
0-
02
b100 6
#112250000000
1!
1%
1-
12
#112260000000
0!
0%
b101 *
0-
02
b101 6
#112270000000
1!
1%
1-
12
#112280000000
0!
0%
b110 *
0-
02
b110 6
#112290000000
1!
1%
1-
12
#112300000000
0!
0%
b111 *
0-
02
b111 6
#112310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#112320000000
0!
0%
b0 *
0-
02
b0 6
#112330000000
1!
1%
1-
12
#112340000000
0!
0%
b1 *
0-
02
b1 6
#112350000000
1!
1%
1-
12
#112360000000
0!
0%
b10 *
0-
02
b10 6
#112370000000
1!
1%
1-
12
#112380000000
0!
0%
b11 *
0-
02
b11 6
#112390000000
1!
1%
1-
12
15
#112400000000
0!
0%
b100 *
0-
02
b100 6
#112410000000
1!
1%
1-
12
#112420000000
0!
0%
b101 *
0-
02
b101 6
#112430000000
1!
1%
1-
12
#112440000000
0!
0%
b110 *
0-
02
b110 6
#112450000000
1!
1%
1-
12
#112460000000
0!
0%
b111 *
0-
02
b111 6
#112470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#112480000000
0!
0%
b0 *
0-
02
b0 6
#112490000000
1!
1%
1-
12
#112500000000
0!
0%
b1 *
0-
02
b1 6
#112510000000
1!
1%
1-
12
#112520000000
0!
0%
b10 *
0-
02
b10 6
#112530000000
1!
1%
1-
12
#112540000000
0!
0%
b11 *
0-
02
b11 6
#112550000000
1!
1%
1-
12
15
#112560000000
0!
0%
b100 *
0-
02
b100 6
#112570000000
1!
1%
1-
12
#112580000000
0!
0%
b101 *
0-
02
b101 6
#112590000000
1!
1%
1-
12
#112600000000
0!
0%
b110 *
0-
02
b110 6
#112610000000
1!
1%
1-
12
#112620000000
0!
0%
b111 *
0-
02
b111 6
#112630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#112640000000
0!
0%
b0 *
0-
02
b0 6
#112650000000
1!
1%
1-
12
#112660000000
0!
0%
b1 *
0-
02
b1 6
#112670000000
1!
1%
1-
12
#112680000000
0!
0%
b10 *
0-
02
b10 6
#112690000000
1!
1%
1-
12
#112700000000
0!
0%
b11 *
0-
02
b11 6
#112710000000
1!
1%
1-
12
15
#112720000000
0!
0%
b100 *
0-
02
b100 6
#112730000000
1!
1%
1-
12
#112740000000
0!
0%
b101 *
0-
02
b101 6
#112750000000
1!
1%
1-
12
#112760000000
0!
0%
b110 *
0-
02
b110 6
#112770000000
1!
1%
1-
12
#112780000000
0!
0%
b111 *
0-
02
b111 6
#112790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#112800000000
0!
0%
b0 *
0-
02
b0 6
#112810000000
1!
1%
1-
12
#112820000000
0!
0%
b1 *
0-
02
b1 6
#112830000000
1!
1%
1-
12
#112840000000
0!
0%
b10 *
0-
02
b10 6
#112850000000
1!
1%
1-
12
#112860000000
0!
0%
b11 *
0-
02
b11 6
#112870000000
1!
1%
1-
12
15
#112880000000
0!
0%
b100 *
0-
02
b100 6
#112890000000
1!
1%
1-
12
#112900000000
0!
0%
b101 *
0-
02
b101 6
#112910000000
1!
1%
1-
12
#112920000000
0!
0%
b110 *
0-
02
b110 6
#112930000000
1!
1%
1-
12
#112940000000
0!
0%
b111 *
0-
02
b111 6
#112950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#112960000000
0!
0%
b0 *
0-
02
b0 6
#112970000000
1!
1%
1-
12
#112980000000
0!
0%
b1 *
0-
02
b1 6
#112990000000
1!
1%
1-
12
#113000000000
0!
0%
b10 *
0-
02
b10 6
#113010000000
1!
1%
1-
12
#113020000000
0!
0%
b11 *
0-
02
b11 6
#113030000000
1!
1%
1-
12
15
#113040000000
0!
0%
b100 *
0-
02
b100 6
#113050000000
1!
1%
1-
12
#113060000000
0!
0%
b101 *
0-
02
b101 6
#113070000000
1!
1%
1-
12
#113080000000
0!
0%
b110 *
0-
02
b110 6
#113090000000
1!
1%
1-
12
#113100000000
0!
0%
b111 *
0-
02
b111 6
#113110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#113120000000
0!
0%
b0 *
0-
02
b0 6
#113130000000
1!
1%
1-
12
#113140000000
0!
0%
b1 *
0-
02
b1 6
#113150000000
1!
1%
1-
12
#113160000000
0!
0%
b10 *
0-
02
b10 6
#113170000000
1!
1%
1-
12
#113180000000
0!
0%
b11 *
0-
02
b11 6
#113190000000
1!
1%
1-
12
15
#113200000000
0!
0%
b100 *
0-
02
b100 6
#113210000000
1!
1%
1-
12
#113220000000
0!
0%
b101 *
0-
02
b101 6
#113230000000
1!
1%
1-
12
#113240000000
0!
0%
b110 *
0-
02
b110 6
#113250000000
1!
1%
1-
12
#113260000000
0!
0%
b111 *
0-
02
b111 6
#113270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#113280000000
0!
0%
b0 *
0-
02
b0 6
#113290000000
1!
1%
1-
12
#113300000000
0!
0%
b1 *
0-
02
b1 6
#113310000000
1!
1%
1-
12
#113320000000
0!
0%
b10 *
0-
02
b10 6
#113330000000
1!
1%
1-
12
#113340000000
0!
0%
b11 *
0-
02
b11 6
#113350000000
1!
1%
1-
12
15
#113360000000
0!
0%
b100 *
0-
02
b100 6
#113370000000
1!
1%
1-
12
#113380000000
0!
0%
b101 *
0-
02
b101 6
#113390000000
1!
1%
1-
12
#113400000000
0!
0%
b110 *
0-
02
b110 6
#113410000000
1!
1%
1-
12
#113420000000
0!
0%
b111 *
0-
02
b111 6
#113430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#113440000000
0!
0%
b0 *
0-
02
b0 6
#113450000000
1!
1%
1-
12
#113460000000
0!
0%
b1 *
0-
02
b1 6
#113470000000
1!
1%
1-
12
#113480000000
0!
0%
b10 *
0-
02
b10 6
#113490000000
1!
1%
1-
12
#113500000000
0!
0%
b11 *
0-
02
b11 6
#113510000000
1!
1%
1-
12
15
#113520000000
0!
0%
b100 *
0-
02
b100 6
#113530000000
1!
1%
1-
12
#113540000000
0!
0%
b101 *
0-
02
b101 6
#113550000000
1!
1%
1-
12
#113560000000
0!
0%
b110 *
0-
02
b110 6
#113570000000
1!
1%
1-
12
#113580000000
0!
0%
b111 *
0-
02
b111 6
#113590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#113600000000
0!
0%
b0 *
0-
02
b0 6
#113610000000
1!
1%
1-
12
#113620000000
0!
0%
b1 *
0-
02
b1 6
#113630000000
1!
1%
1-
12
#113640000000
0!
0%
b10 *
0-
02
b10 6
#113650000000
1!
1%
1-
12
#113660000000
0!
0%
b11 *
0-
02
b11 6
#113670000000
1!
1%
1-
12
15
#113680000000
0!
0%
b100 *
0-
02
b100 6
#113690000000
1!
1%
1-
12
#113700000000
0!
0%
b101 *
0-
02
b101 6
#113710000000
1!
1%
1-
12
#113720000000
0!
0%
b110 *
0-
02
b110 6
#113730000000
1!
1%
1-
12
#113740000000
0!
0%
b111 *
0-
02
b111 6
#113750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#113760000000
0!
0%
b0 *
0-
02
b0 6
#113770000000
1!
1%
1-
12
#113780000000
0!
0%
b1 *
0-
02
b1 6
#113790000000
1!
1%
1-
12
#113800000000
0!
0%
b10 *
0-
02
b10 6
#113810000000
1!
1%
1-
12
#113820000000
0!
0%
b11 *
0-
02
b11 6
#113830000000
1!
1%
1-
12
15
#113840000000
0!
0%
b100 *
0-
02
b100 6
#113850000000
1!
1%
1-
12
#113860000000
0!
0%
b101 *
0-
02
b101 6
#113870000000
1!
1%
1-
12
#113880000000
0!
0%
b110 *
0-
02
b110 6
#113890000000
1!
1%
1-
12
#113900000000
0!
0%
b111 *
0-
02
b111 6
#113910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#113920000000
0!
0%
b0 *
0-
02
b0 6
#113930000000
1!
1%
1-
12
#113940000000
0!
0%
b1 *
0-
02
b1 6
#113950000000
1!
1%
1-
12
#113960000000
0!
0%
b10 *
0-
02
b10 6
#113970000000
1!
1%
1-
12
#113980000000
0!
0%
b11 *
0-
02
b11 6
#113990000000
1!
1%
1-
12
15
#114000000000
0!
0%
b100 *
0-
02
b100 6
#114010000000
1!
1%
1-
12
#114020000000
0!
0%
b101 *
0-
02
b101 6
#114030000000
1!
1%
1-
12
#114040000000
0!
0%
b110 *
0-
02
b110 6
#114050000000
1!
1%
1-
12
#114060000000
0!
0%
b111 *
0-
02
b111 6
#114070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#114080000000
0!
0%
b0 *
0-
02
b0 6
#114090000000
1!
1%
1-
12
#114100000000
0!
0%
b1 *
0-
02
b1 6
#114110000000
1!
1%
1-
12
#114120000000
0!
0%
b10 *
0-
02
b10 6
#114130000000
1!
1%
1-
12
#114140000000
0!
0%
b11 *
0-
02
b11 6
#114150000000
1!
1%
1-
12
15
#114160000000
0!
0%
b100 *
0-
02
b100 6
#114170000000
1!
1%
1-
12
#114180000000
0!
0%
b101 *
0-
02
b101 6
#114190000000
1!
1%
1-
12
#114200000000
0!
0%
b110 *
0-
02
b110 6
#114210000000
1!
1%
1-
12
#114220000000
0!
0%
b111 *
0-
02
b111 6
#114230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#114240000000
0!
0%
b0 *
0-
02
b0 6
#114250000000
1!
1%
1-
12
#114260000000
0!
0%
b1 *
0-
02
b1 6
#114270000000
1!
1%
1-
12
#114280000000
0!
0%
b10 *
0-
02
b10 6
#114290000000
1!
1%
1-
12
#114300000000
0!
0%
b11 *
0-
02
b11 6
#114310000000
1!
1%
1-
12
15
#114320000000
0!
0%
b100 *
0-
02
b100 6
#114330000000
1!
1%
1-
12
#114340000000
0!
0%
b101 *
0-
02
b101 6
#114350000000
1!
1%
1-
12
#114360000000
0!
0%
b110 *
0-
02
b110 6
#114370000000
1!
1%
1-
12
#114380000000
0!
0%
b111 *
0-
02
b111 6
#114390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#114400000000
0!
0%
b0 *
0-
02
b0 6
#114410000000
1!
1%
1-
12
#114420000000
0!
0%
b1 *
0-
02
b1 6
#114430000000
1!
1%
1-
12
#114440000000
0!
0%
b10 *
0-
02
b10 6
#114450000000
1!
1%
1-
12
#114460000000
0!
0%
b11 *
0-
02
b11 6
#114470000000
1!
1%
1-
12
15
#114480000000
0!
0%
b100 *
0-
02
b100 6
#114490000000
1!
1%
1-
12
#114500000000
0!
0%
b101 *
0-
02
b101 6
#114510000000
1!
1%
1-
12
#114520000000
0!
0%
b110 *
0-
02
b110 6
#114530000000
1!
1%
1-
12
#114540000000
0!
0%
b111 *
0-
02
b111 6
#114550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#114560000000
0!
0%
b0 *
0-
02
b0 6
#114570000000
1!
1%
1-
12
#114580000000
0!
0%
b1 *
0-
02
b1 6
#114590000000
1!
1%
1-
12
#114600000000
0!
0%
b10 *
0-
02
b10 6
#114610000000
1!
1%
1-
12
#114620000000
0!
0%
b11 *
0-
02
b11 6
#114630000000
1!
1%
1-
12
15
#114640000000
0!
0%
b100 *
0-
02
b100 6
#114650000000
1!
1%
1-
12
#114660000000
0!
0%
b101 *
0-
02
b101 6
#114670000000
1!
1%
1-
12
#114680000000
0!
0%
b110 *
0-
02
b110 6
#114690000000
1!
1%
1-
12
#114700000000
0!
0%
b111 *
0-
02
b111 6
#114710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#114720000000
0!
0%
b0 *
0-
02
b0 6
#114730000000
1!
1%
1-
12
#114740000000
0!
0%
b1 *
0-
02
b1 6
#114750000000
1!
1%
1-
12
#114760000000
0!
0%
b10 *
0-
02
b10 6
#114770000000
1!
1%
1-
12
#114780000000
0!
0%
b11 *
0-
02
b11 6
#114790000000
1!
1%
1-
12
15
#114800000000
0!
0%
b100 *
0-
02
b100 6
#114810000000
1!
1%
1-
12
#114820000000
0!
0%
b101 *
0-
02
b101 6
#114830000000
1!
1%
1-
12
#114840000000
0!
0%
b110 *
0-
02
b110 6
#114850000000
1!
1%
1-
12
#114860000000
0!
0%
b111 *
0-
02
b111 6
#114870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#114880000000
0!
0%
b0 *
0-
02
b0 6
#114890000000
1!
1%
1-
12
#114900000000
0!
0%
b1 *
0-
02
b1 6
#114910000000
1!
1%
1-
12
#114920000000
0!
0%
b10 *
0-
02
b10 6
#114930000000
1!
1%
1-
12
#114940000000
0!
0%
b11 *
0-
02
b11 6
#114950000000
1!
1%
1-
12
15
#114960000000
0!
0%
b100 *
0-
02
b100 6
#114970000000
1!
1%
1-
12
#114980000000
0!
0%
b101 *
0-
02
b101 6
#114990000000
1!
1%
1-
12
#115000000000
0!
0%
b110 *
0-
02
b110 6
#115010000000
1!
1%
1-
12
#115020000000
0!
0%
b111 *
0-
02
b111 6
#115030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#115040000000
0!
0%
b0 *
0-
02
b0 6
#115050000000
1!
1%
1-
12
#115060000000
0!
0%
b1 *
0-
02
b1 6
#115070000000
1!
1%
1-
12
#115080000000
0!
0%
b10 *
0-
02
b10 6
#115090000000
1!
1%
1-
12
#115100000000
0!
0%
b11 *
0-
02
b11 6
#115110000000
1!
1%
1-
12
15
#115120000000
0!
0%
b100 *
0-
02
b100 6
#115130000000
1!
1%
1-
12
#115140000000
0!
0%
b101 *
0-
02
b101 6
#115150000000
1!
1%
1-
12
#115160000000
0!
0%
b110 *
0-
02
b110 6
#115170000000
1!
1%
1-
12
#115180000000
0!
0%
b111 *
0-
02
b111 6
#115190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#115200000000
0!
0%
b0 *
0-
02
b0 6
#115210000000
1!
1%
1-
12
#115220000000
0!
0%
b1 *
0-
02
b1 6
#115230000000
1!
1%
1-
12
#115240000000
0!
0%
b10 *
0-
02
b10 6
#115250000000
1!
1%
1-
12
#115260000000
0!
0%
b11 *
0-
02
b11 6
#115270000000
1!
1%
1-
12
15
#115280000000
0!
0%
b100 *
0-
02
b100 6
#115290000000
1!
1%
1-
12
#115300000000
0!
0%
b101 *
0-
02
b101 6
#115310000000
1!
1%
1-
12
#115320000000
0!
0%
b110 *
0-
02
b110 6
#115330000000
1!
1%
1-
12
#115340000000
0!
0%
b111 *
0-
02
b111 6
#115350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#115360000000
0!
0%
b0 *
0-
02
b0 6
#115370000000
1!
1%
1-
12
#115380000000
0!
0%
b1 *
0-
02
b1 6
#115390000000
1!
1%
1-
12
#115400000000
0!
0%
b10 *
0-
02
b10 6
#115410000000
1!
1%
1-
12
#115420000000
0!
0%
b11 *
0-
02
b11 6
#115430000000
1!
1%
1-
12
15
#115440000000
0!
0%
b100 *
0-
02
b100 6
#115450000000
1!
1%
1-
12
#115460000000
0!
0%
b101 *
0-
02
b101 6
#115470000000
1!
1%
1-
12
#115480000000
0!
0%
b110 *
0-
02
b110 6
#115490000000
1!
1%
1-
12
#115500000000
0!
0%
b111 *
0-
02
b111 6
#115510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#115520000000
0!
0%
b0 *
0-
02
b0 6
#115530000000
1!
1%
1-
12
#115540000000
0!
0%
b1 *
0-
02
b1 6
#115550000000
1!
1%
1-
12
#115560000000
0!
0%
b10 *
0-
02
b10 6
#115570000000
1!
1%
1-
12
#115580000000
0!
0%
b11 *
0-
02
b11 6
#115590000000
1!
1%
1-
12
15
#115600000000
0!
0%
b100 *
0-
02
b100 6
#115610000000
1!
1%
1-
12
#115620000000
0!
0%
b101 *
0-
02
b101 6
#115630000000
1!
1%
1-
12
#115640000000
0!
0%
b110 *
0-
02
b110 6
#115650000000
1!
1%
1-
12
#115660000000
0!
0%
b111 *
0-
02
b111 6
#115670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#115680000000
0!
0%
b0 *
0-
02
b0 6
#115690000000
1!
1%
1-
12
#115700000000
0!
0%
b1 *
0-
02
b1 6
#115710000000
1!
1%
1-
12
#115720000000
0!
0%
b10 *
0-
02
b10 6
#115730000000
1!
1%
1-
12
#115740000000
0!
0%
b11 *
0-
02
b11 6
#115750000000
1!
1%
1-
12
15
#115760000000
0!
0%
b100 *
0-
02
b100 6
#115770000000
1!
1%
1-
12
#115780000000
0!
0%
b101 *
0-
02
b101 6
#115790000000
1!
1%
1-
12
#115800000000
0!
0%
b110 *
0-
02
b110 6
#115810000000
1!
1%
1-
12
#115820000000
0!
0%
b111 *
0-
02
b111 6
#115830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#115840000000
0!
0%
b0 *
0-
02
b0 6
#115850000000
1!
1%
1-
12
#115860000000
0!
0%
b1 *
0-
02
b1 6
#115870000000
1!
1%
1-
12
#115880000000
0!
0%
b10 *
0-
02
b10 6
#115890000000
1!
1%
1-
12
#115900000000
0!
0%
b11 *
0-
02
b11 6
#115910000000
1!
1%
1-
12
15
#115920000000
0!
0%
b100 *
0-
02
b100 6
#115930000000
1!
1%
1-
12
#115940000000
0!
0%
b101 *
0-
02
b101 6
#115950000000
1!
1%
1-
12
#115960000000
0!
0%
b110 *
0-
02
b110 6
#115970000000
1!
1%
1-
12
#115980000000
0!
0%
b111 *
0-
02
b111 6
#115990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#116000000000
0!
0%
b0 *
0-
02
b0 6
#116010000000
1!
1%
1-
12
#116020000000
0!
0%
b1 *
0-
02
b1 6
#116030000000
1!
1%
1-
12
#116040000000
0!
0%
b10 *
0-
02
b10 6
#116050000000
1!
1%
1-
12
#116060000000
0!
0%
b11 *
0-
02
b11 6
#116070000000
1!
1%
1-
12
15
#116080000000
0!
0%
b100 *
0-
02
b100 6
#116090000000
1!
1%
1-
12
#116100000000
0!
0%
b101 *
0-
02
b101 6
#116110000000
1!
1%
1-
12
#116120000000
0!
0%
b110 *
0-
02
b110 6
#116130000000
1!
1%
1-
12
#116140000000
0!
0%
b111 *
0-
02
b111 6
#116150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#116160000000
0!
0%
b0 *
0-
02
b0 6
#116170000000
1!
1%
1-
12
#116180000000
0!
0%
b1 *
0-
02
b1 6
#116190000000
1!
1%
1-
12
#116200000000
0!
0%
b10 *
0-
02
b10 6
#116210000000
1!
1%
1-
12
#116220000000
0!
0%
b11 *
0-
02
b11 6
#116230000000
1!
1%
1-
12
15
#116240000000
0!
0%
b100 *
0-
02
b100 6
#116250000000
1!
1%
1-
12
#116260000000
0!
0%
b101 *
0-
02
b101 6
#116270000000
1!
1%
1-
12
#116280000000
0!
0%
b110 *
0-
02
b110 6
#116290000000
1!
1%
1-
12
#116300000000
0!
0%
b111 *
0-
02
b111 6
#116310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#116320000000
0!
0%
b0 *
0-
02
b0 6
#116330000000
1!
1%
1-
12
#116340000000
0!
0%
b1 *
0-
02
b1 6
#116350000000
1!
1%
1-
12
#116360000000
0!
0%
b10 *
0-
02
b10 6
#116370000000
1!
1%
1-
12
#116380000000
0!
0%
b11 *
0-
02
b11 6
#116390000000
1!
1%
1-
12
15
#116400000000
0!
0%
b100 *
0-
02
b100 6
#116410000000
1!
1%
1-
12
#116420000000
0!
0%
b101 *
0-
02
b101 6
#116430000000
1!
1%
1-
12
#116440000000
0!
0%
b110 *
0-
02
b110 6
#116450000000
1!
1%
1-
12
#116460000000
0!
0%
b111 *
0-
02
b111 6
#116470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#116480000000
0!
0%
b0 *
0-
02
b0 6
#116490000000
1!
1%
1-
12
#116500000000
0!
0%
b1 *
0-
02
b1 6
#116510000000
1!
1%
1-
12
#116520000000
0!
0%
b10 *
0-
02
b10 6
#116530000000
1!
1%
1-
12
#116540000000
0!
0%
b11 *
0-
02
b11 6
#116550000000
1!
1%
1-
12
15
#116560000000
0!
0%
b100 *
0-
02
b100 6
#116570000000
1!
1%
1-
12
#116580000000
0!
0%
b101 *
0-
02
b101 6
#116590000000
1!
1%
1-
12
#116600000000
0!
0%
b110 *
0-
02
b110 6
#116610000000
1!
1%
1-
12
#116620000000
0!
0%
b111 *
0-
02
b111 6
#116630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#116640000000
0!
0%
b0 *
0-
02
b0 6
#116650000000
1!
1%
1-
12
#116660000000
0!
0%
b1 *
0-
02
b1 6
#116670000000
1!
1%
1-
12
#116680000000
0!
0%
b10 *
0-
02
b10 6
#116690000000
1!
1%
1-
12
#116700000000
0!
0%
b11 *
0-
02
b11 6
#116710000000
1!
1%
1-
12
15
#116720000000
0!
0%
b100 *
0-
02
b100 6
#116730000000
1!
1%
1-
12
#116740000000
0!
0%
b101 *
0-
02
b101 6
#116750000000
1!
1%
1-
12
#116760000000
0!
0%
b110 *
0-
02
b110 6
#116770000000
1!
1%
1-
12
#116780000000
0!
0%
b111 *
0-
02
b111 6
#116790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#116800000000
0!
0%
b0 *
0-
02
b0 6
#116810000000
1!
1%
1-
12
#116820000000
0!
0%
b1 *
0-
02
b1 6
#116830000000
1!
1%
1-
12
#116840000000
0!
0%
b10 *
0-
02
b10 6
#116850000000
1!
1%
1-
12
#116860000000
0!
0%
b11 *
0-
02
b11 6
#116870000000
1!
1%
1-
12
15
#116880000000
0!
0%
b100 *
0-
02
b100 6
#116890000000
1!
1%
1-
12
#116900000000
0!
0%
b101 *
0-
02
b101 6
#116910000000
1!
1%
1-
12
#116920000000
0!
0%
b110 *
0-
02
b110 6
#116930000000
1!
1%
1-
12
#116940000000
0!
0%
b111 *
0-
02
b111 6
#116950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#116960000000
0!
0%
b0 *
0-
02
b0 6
#116970000000
1!
1%
1-
12
#116980000000
0!
0%
b1 *
0-
02
b1 6
#116990000000
1!
1%
1-
12
#117000000000
0!
0%
b10 *
0-
02
b10 6
#117010000000
1!
1%
1-
12
#117020000000
0!
0%
b11 *
0-
02
b11 6
#117030000000
1!
1%
1-
12
15
#117040000000
0!
0%
b100 *
0-
02
b100 6
#117050000000
1!
1%
1-
12
#117060000000
0!
0%
b101 *
0-
02
b101 6
#117070000000
1!
1%
1-
12
#117080000000
0!
0%
b110 *
0-
02
b110 6
#117090000000
1!
1%
1-
12
#117100000000
0!
0%
b111 *
0-
02
b111 6
#117110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#117120000000
0!
0%
b0 *
0-
02
b0 6
#117130000000
1!
1%
1-
12
#117140000000
0!
0%
b1 *
0-
02
b1 6
#117150000000
1!
1%
1-
12
#117160000000
0!
0%
b10 *
0-
02
b10 6
#117170000000
1!
1%
1-
12
#117180000000
0!
0%
b11 *
0-
02
b11 6
#117190000000
1!
1%
1-
12
15
#117200000000
0!
0%
b100 *
0-
02
b100 6
#117210000000
1!
1%
1-
12
#117220000000
0!
0%
b101 *
0-
02
b101 6
#117230000000
1!
1%
1-
12
#117240000000
0!
0%
b110 *
0-
02
b110 6
#117250000000
1!
1%
1-
12
#117260000000
0!
0%
b111 *
0-
02
b111 6
#117270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#117280000000
0!
0%
b0 *
0-
02
b0 6
#117290000000
1!
1%
1-
12
#117300000000
0!
0%
b1 *
0-
02
b1 6
#117310000000
1!
1%
1-
12
#117320000000
0!
0%
b10 *
0-
02
b10 6
#117330000000
1!
1%
1-
12
#117340000000
0!
0%
b11 *
0-
02
b11 6
#117350000000
1!
1%
1-
12
15
#117360000000
0!
0%
b100 *
0-
02
b100 6
#117370000000
1!
1%
1-
12
#117380000000
0!
0%
b101 *
0-
02
b101 6
#117390000000
1!
1%
1-
12
#117400000000
0!
0%
b110 *
0-
02
b110 6
#117410000000
1!
1%
1-
12
#117420000000
0!
0%
b111 *
0-
02
b111 6
#117430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#117440000000
0!
0%
b0 *
0-
02
b0 6
#117450000000
1!
1%
1-
12
#117460000000
0!
0%
b1 *
0-
02
b1 6
#117470000000
1!
1%
1-
12
#117480000000
0!
0%
b10 *
0-
02
b10 6
#117490000000
1!
1%
1-
12
#117500000000
0!
0%
b11 *
0-
02
b11 6
#117510000000
1!
1%
1-
12
15
#117520000000
0!
0%
b100 *
0-
02
b100 6
#117530000000
1!
1%
1-
12
#117540000000
0!
0%
b101 *
0-
02
b101 6
#117550000000
1!
1%
1-
12
#117560000000
0!
0%
b110 *
0-
02
b110 6
#117570000000
1!
1%
1-
12
#117580000000
0!
0%
b111 *
0-
02
b111 6
#117590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#117600000000
0!
0%
b0 *
0-
02
b0 6
#117610000000
1!
1%
1-
12
#117620000000
0!
0%
b1 *
0-
02
b1 6
#117630000000
1!
1%
1-
12
#117640000000
0!
0%
b10 *
0-
02
b10 6
#117650000000
1!
1%
1-
12
#117660000000
0!
0%
b11 *
0-
02
b11 6
#117670000000
1!
1%
1-
12
15
#117680000000
0!
0%
b100 *
0-
02
b100 6
#117690000000
1!
1%
1-
12
#117700000000
0!
0%
b101 *
0-
02
b101 6
#117710000000
1!
1%
1-
12
#117720000000
0!
0%
b110 *
0-
02
b110 6
#117730000000
1!
1%
1-
12
#117740000000
0!
0%
b111 *
0-
02
b111 6
#117750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#117760000000
0!
0%
b0 *
0-
02
b0 6
#117770000000
1!
1%
1-
12
#117780000000
0!
0%
b1 *
0-
02
b1 6
#117790000000
1!
1%
1-
12
#117800000000
0!
0%
b10 *
0-
02
b10 6
#117810000000
1!
1%
1-
12
#117820000000
0!
0%
b11 *
0-
02
b11 6
#117830000000
1!
1%
1-
12
15
#117840000000
0!
0%
b100 *
0-
02
b100 6
#117850000000
1!
1%
1-
12
#117860000000
0!
0%
b101 *
0-
02
b101 6
#117870000000
1!
1%
1-
12
#117880000000
0!
0%
b110 *
0-
02
b110 6
#117890000000
1!
1%
1-
12
#117900000000
0!
0%
b111 *
0-
02
b111 6
#117910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#117920000000
0!
0%
b0 *
0-
02
b0 6
#117930000000
1!
1%
1-
12
#117940000000
0!
0%
b1 *
0-
02
b1 6
#117950000000
1!
1%
1-
12
#117960000000
0!
0%
b10 *
0-
02
b10 6
#117970000000
1!
1%
1-
12
#117980000000
0!
0%
b11 *
0-
02
b11 6
#117990000000
1!
1%
1-
12
15
#118000000000
0!
0%
b100 *
0-
02
b100 6
#118010000000
1!
1%
1-
12
#118020000000
0!
0%
b101 *
0-
02
b101 6
#118030000000
1!
1%
1-
12
#118040000000
0!
0%
b110 *
0-
02
b110 6
#118050000000
1!
1%
1-
12
#118060000000
0!
0%
b111 *
0-
02
b111 6
#118070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#118080000000
0!
0%
b0 *
0-
02
b0 6
#118090000000
1!
1%
1-
12
#118100000000
0!
0%
b1 *
0-
02
b1 6
#118110000000
1!
1%
1-
12
#118120000000
0!
0%
b10 *
0-
02
b10 6
#118130000000
1!
1%
1-
12
#118140000000
0!
0%
b11 *
0-
02
b11 6
#118150000000
1!
1%
1-
12
15
#118160000000
0!
0%
b100 *
0-
02
b100 6
#118170000000
1!
1%
1-
12
#118180000000
0!
0%
b101 *
0-
02
b101 6
#118190000000
1!
1%
1-
12
#118200000000
0!
0%
b110 *
0-
02
b110 6
#118210000000
1!
1%
1-
12
#118220000000
0!
0%
b111 *
0-
02
b111 6
#118230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#118240000000
0!
0%
b0 *
0-
02
b0 6
#118250000000
1!
1%
1-
12
#118260000000
0!
0%
b1 *
0-
02
b1 6
#118270000000
1!
1%
1-
12
#118280000000
0!
0%
b10 *
0-
02
b10 6
#118290000000
1!
1%
1-
12
#118300000000
0!
0%
b11 *
0-
02
b11 6
#118310000000
1!
1%
1-
12
15
#118320000000
0!
0%
b100 *
0-
02
b100 6
#118330000000
1!
1%
1-
12
#118340000000
0!
0%
b101 *
0-
02
b101 6
#118350000000
1!
1%
1-
12
#118360000000
0!
0%
b110 *
0-
02
b110 6
#118370000000
1!
1%
1-
12
#118380000000
0!
0%
b111 *
0-
02
b111 6
#118390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#118400000000
0!
0%
b0 *
0-
02
b0 6
#118410000000
1!
1%
1-
12
#118420000000
0!
0%
b1 *
0-
02
b1 6
#118430000000
1!
1%
1-
12
#118440000000
0!
0%
b10 *
0-
02
b10 6
#118450000000
1!
1%
1-
12
#118460000000
0!
0%
b11 *
0-
02
b11 6
#118470000000
1!
1%
1-
12
15
#118480000000
0!
0%
b100 *
0-
02
b100 6
#118490000000
1!
1%
1-
12
#118500000000
0!
0%
b101 *
0-
02
b101 6
#118510000000
1!
1%
1-
12
#118520000000
0!
0%
b110 *
0-
02
b110 6
#118530000000
1!
1%
1-
12
#118540000000
0!
0%
b111 *
0-
02
b111 6
#118550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#118560000000
0!
0%
b0 *
0-
02
b0 6
#118570000000
1!
1%
1-
12
#118580000000
0!
0%
b1 *
0-
02
b1 6
#118590000000
1!
1%
1-
12
#118600000000
0!
0%
b10 *
0-
02
b10 6
#118610000000
1!
1%
1-
12
#118620000000
0!
0%
b11 *
0-
02
b11 6
#118630000000
1!
1%
1-
12
15
#118640000000
0!
0%
b100 *
0-
02
b100 6
#118650000000
1!
1%
1-
12
#118660000000
0!
0%
b101 *
0-
02
b101 6
#118670000000
1!
1%
1-
12
#118680000000
0!
0%
b110 *
0-
02
b110 6
#118690000000
1!
1%
1-
12
#118700000000
0!
0%
b111 *
0-
02
b111 6
#118710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#118720000000
0!
0%
b0 *
0-
02
b0 6
#118730000000
1!
1%
1-
12
#118740000000
0!
0%
b1 *
0-
02
b1 6
#118750000000
1!
1%
1-
12
#118760000000
0!
0%
b10 *
0-
02
b10 6
#118770000000
1!
1%
1-
12
#118780000000
0!
0%
b11 *
0-
02
b11 6
#118790000000
1!
1%
1-
12
15
#118800000000
0!
0%
b100 *
0-
02
b100 6
#118810000000
1!
1%
1-
12
#118820000000
0!
0%
b101 *
0-
02
b101 6
#118830000000
1!
1%
1-
12
#118840000000
0!
0%
b110 *
0-
02
b110 6
#118850000000
1!
1%
1-
12
#118860000000
0!
0%
b111 *
0-
02
b111 6
#118870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#118880000000
0!
0%
b0 *
0-
02
b0 6
#118890000000
1!
1%
1-
12
#118900000000
0!
0%
b1 *
0-
02
b1 6
#118910000000
1!
1%
1-
12
#118920000000
0!
0%
b10 *
0-
02
b10 6
#118930000000
1!
1%
1-
12
#118940000000
0!
0%
b11 *
0-
02
b11 6
#118950000000
1!
1%
1-
12
15
#118960000000
0!
0%
b100 *
0-
02
b100 6
#118970000000
1!
1%
1-
12
#118980000000
0!
0%
b101 *
0-
02
b101 6
#118990000000
1!
1%
1-
12
#119000000000
0!
0%
b110 *
0-
02
b110 6
#119010000000
1!
1%
1-
12
#119020000000
0!
0%
b111 *
0-
02
b111 6
#119030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#119040000000
0!
0%
b0 *
0-
02
b0 6
#119050000000
1!
1%
1-
12
#119060000000
0!
0%
b1 *
0-
02
b1 6
#119070000000
1!
1%
1-
12
#119080000000
0!
0%
b10 *
0-
02
b10 6
#119090000000
1!
1%
1-
12
#119100000000
0!
0%
b11 *
0-
02
b11 6
#119110000000
1!
1%
1-
12
15
#119120000000
0!
0%
b100 *
0-
02
b100 6
#119130000000
1!
1%
1-
12
#119140000000
0!
0%
b101 *
0-
02
b101 6
#119150000000
1!
1%
1-
12
#119160000000
0!
0%
b110 *
0-
02
b110 6
#119170000000
1!
1%
1-
12
#119180000000
0!
0%
b111 *
0-
02
b111 6
#119190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#119200000000
0!
0%
b0 *
0-
02
b0 6
#119210000000
1!
1%
1-
12
#119220000000
0!
0%
b1 *
0-
02
b1 6
#119230000000
1!
1%
1-
12
#119240000000
0!
0%
b10 *
0-
02
b10 6
#119250000000
1!
1%
1-
12
#119260000000
0!
0%
b11 *
0-
02
b11 6
#119270000000
1!
1%
1-
12
15
#119280000000
0!
0%
b100 *
0-
02
b100 6
#119290000000
1!
1%
1-
12
#119300000000
0!
0%
b101 *
0-
02
b101 6
#119310000000
1!
1%
1-
12
#119320000000
0!
0%
b110 *
0-
02
b110 6
#119330000000
1!
1%
1-
12
#119340000000
0!
0%
b111 *
0-
02
b111 6
#119350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#119360000000
0!
0%
b0 *
0-
02
b0 6
#119370000000
1!
1%
1-
12
#119380000000
0!
0%
b1 *
0-
02
b1 6
#119390000000
1!
1%
1-
12
#119400000000
0!
0%
b10 *
0-
02
b10 6
#119410000000
1!
1%
1-
12
#119420000000
0!
0%
b11 *
0-
02
b11 6
#119430000000
1!
1%
1-
12
15
#119440000000
0!
0%
b100 *
0-
02
b100 6
#119450000000
1!
1%
1-
12
#119460000000
0!
0%
b101 *
0-
02
b101 6
#119470000000
1!
1%
1-
12
#119480000000
0!
0%
b110 *
0-
02
b110 6
#119490000000
1!
1%
1-
12
#119500000000
0!
0%
b111 *
0-
02
b111 6
#119510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#119520000000
0!
0%
b0 *
0-
02
b0 6
#119530000000
1!
1%
1-
12
#119540000000
0!
0%
b1 *
0-
02
b1 6
#119550000000
1!
1%
1-
12
#119560000000
0!
0%
b10 *
0-
02
b10 6
#119570000000
1!
1%
1-
12
#119580000000
0!
0%
b11 *
0-
02
b11 6
#119590000000
1!
1%
1-
12
15
#119600000000
0!
0%
b100 *
0-
02
b100 6
#119610000000
1!
1%
1-
12
#119620000000
0!
0%
b101 *
0-
02
b101 6
#119630000000
1!
1%
1-
12
#119640000000
0!
0%
b110 *
0-
02
b110 6
#119650000000
1!
1%
1-
12
#119660000000
0!
0%
b111 *
0-
02
b111 6
#119670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#119680000000
0!
0%
b0 *
0-
02
b0 6
#119690000000
1!
1%
1-
12
#119700000000
0!
0%
b1 *
0-
02
b1 6
#119710000000
1!
1%
1-
12
#119720000000
0!
0%
b10 *
0-
02
b10 6
#119730000000
1!
1%
1-
12
#119740000000
0!
0%
b11 *
0-
02
b11 6
#119750000000
1!
1%
1-
12
15
#119760000000
0!
0%
b100 *
0-
02
b100 6
#119770000000
1!
1%
1-
12
#119780000000
0!
0%
b101 *
0-
02
b101 6
#119790000000
1!
1%
1-
12
#119800000000
0!
0%
b110 *
0-
02
b110 6
#119810000000
1!
1%
1-
12
#119820000000
0!
0%
b111 *
0-
02
b111 6
#119830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#119840000000
0!
0%
b0 *
0-
02
b0 6
#119850000000
1!
1%
1-
12
#119860000000
0!
0%
b1 *
0-
02
b1 6
#119870000000
1!
1%
1-
12
#119880000000
0!
0%
b10 *
0-
02
b10 6
#119890000000
1!
1%
1-
12
#119900000000
0!
0%
b11 *
0-
02
b11 6
#119910000000
1!
1%
1-
12
15
#119920000000
0!
0%
b100 *
0-
02
b100 6
#119930000000
1!
1%
1-
12
#119940000000
0!
0%
b101 *
0-
02
b101 6
#119950000000
1!
1%
1-
12
#119960000000
0!
0%
b110 *
0-
02
b110 6
#119970000000
1!
1%
1-
12
#119980000000
0!
0%
b111 *
0-
02
b111 6
#119990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#120000000000
0!
0%
b0 *
0-
02
b0 6
#120010000000
1!
1%
1-
12
#120020000000
0!
0%
b1 *
0-
02
b1 6
#120030000000
1!
1%
1-
12
#120040000000
0!
0%
b10 *
0-
02
b10 6
#120050000000
1!
1%
1-
12
#120060000000
0!
0%
b11 *
0-
02
b11 6
#120070000000
1!
1%
1-
12
15
#120080000000
0!
0%
b100 *
0-
02
b100 6
#120090000000
1!
1%
1-
12
#120100000000
0!
0%
b101 *
0-
02
b101 6
#120110000000
1!
1%
1-
12
#120120000000
0!
0%
b110 *
0-
02
b110 6
#120130000000
1!
1%
1-
12
#120140000000
0!
0%
b111 *
0-
02
b111 6
#120150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#120160000000
0!
0%
b0 *
0-
02
b0 6
#120170000000
1!
1%
1-
12
#120180000000
0!
0%
b1 *
0-
02
b1 6
#120190000000
1!
1%
1-
12
#120200000000
0!
0%
b10 *
0-
02
b10 6
#120210000000
1!
1%
1-
12
#120220000000
0!
0%
b11 *
0-
02
b11 6
#120230000000
1!
1%
1-
12
15
#120240000000
0!
0%
b100 *
0-
02
b100 6
#120250000000
1!
1%
1-
12
#120260000000
0!
0%
b101 *
0-
02
b101 6
#120270000000
1!
1%
1-
12
#120280000000
0!
0%
b110 *
0-
02
b110 6
#120290000000
1!
1%
1-
12
#120300000000
0!
0%
b111 *
0-
02
b111 6
#120310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#120320000000
0!
0%
b0 *
0-
02
b0 6
#120330000000
1!
1%
1-
12
#120340000000
0!
0%
b1 *
0-
02
b1 6
#120350000000
1!
1%
1-
12
#120360000000
0!
0%
b10 *
0-
02
b10 6
#120370000000
1!
1%
1-
12
#120380000000
0!
0%
b11 *
0-
02
b11 6
#120390000000
1!
1%
1-
12
15
#120400000000
0!
0%
b100 *
0-
02
b100 6
#120410000000
1!
1%
1-
12
#120420000000
0!
0%
b101 *
0-
02
b101 6
#120430000000
1!
1%
1-
12
#120440000000
0!
0%
b110 *
0-
02
b110 6
#120450000000
1!
1%
1-
12
#120460000000
0!
0%
b111 *
0-
02
b111 6
#120470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#120480000000
0!
0%
b0 *
0-
02
b0 6
#120490000000
1!
1%
1-
12
#120500000000
0!
0%
b1 *
0-
02
b1 6
#120510000000
1!
1%
1-
12
#120520000000
0!
0%
b10 *
0-
02
b10 6
#120530000000
1!
1%
1-
12
#120540000000
0!
0%
b11 *
0-
02
b11 6
#120550000000
1!
1%
1-
12
15
#120560000000
0!
0%
b100 *
0-
02
b100 6
#120570000000
1!
1%
1-
12
#120580000000
0!
0%
b101 *
0-
02
b101 6
#120590000000
1!
1%
1-
12
#120600000000
0!
0%
b110 *
0-
02
b110 6
#120610000000
1!
1%
1-
12
#120620000000
0!
0%
b111 *
0-
02
b111 6
#120630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#120640000000
0!
0%
b0 *
0-
02
b0 6
#120650000000
1!
1%
1-
12
#120660000000
0!
0%
b1 *
0-
02
b1 6
#120670000000
1!
1%
1-
12
#120680000000
0!
0%
b10 *
0-
02
b10 6
#120690000000
1!
1%
1-
12
#120700000000
0!
0%
b11 *
0-
02
b11 6
#120710000000
1!
1%
1-
12
15
#120720000000
0!
0%
b100 *
0-
02
b100 6
#120730000000
1!
1%
1-
12
#120740000000
0!
0%
b101 *
0-
02
b101 6
#120750000000
1!
1%
1-
12
#120760000000
0!
0%
b110 *
0-
02
b110 6
#120770000000
1!
1%
1-
12
#120780000000
0!
0%
b111 *
0-
02
b111 6
#120790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#120800000000
0!
0%
b0 *
0-
02
b0 6
#120810000000
1!
1%
1-
12
#120820000000
0!
0%
b1 *
0-
02
b1 6
#120830000000
1!
1%
1-
12
#120840000000
0!
0%
b10 *
0-
02
b10 6
#120850000000
1!
1%
1-
12
#120860000000
0!
0%
b11 *
0-
02
b11 6
#120870000000
1!
1%
1-
12
15
#120880000000
0!
0%
b100 *
0-
02
b100 6
#120890000000
1!
1%
1-
12
#120900000000
0!
0%
b101 *
0-
02
b101 6
#120910000000
1!
1%
1-
12
#120920000000
0!
0%
b110 *
0-
02
b110 6
#120930000000
1!
1%
1-
12
#120940000000
0!
0%
b111 *
0-
02
b111 6
#120950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#120960000000
0!
0%
b0 *
0-
02
b0 6
#120970000000
1!
1%
1-
12
#120980000000
0!
0%
b1 *
0-
02
b1 6
#120990000000
1!
1%
1-
12
#121000000000
0!
0%
b10 *
0-
02
b10 6
#121010000000
1!
1%
1-
12
#121020000000
0!
0%
b11 *
0-
02
b11 6
#121030000000
1!
1%
1-
12
15
#121040000000
0!
0%
b100 *
0-
02
b100 6
#121050000000
1!
1%
1-
12
#121060000000
0!
0%
b101 *
0-
02
b101 6
#121070000000
1!
1%
1-
12
#121080000000
0!
0%
b110 *
0-
02
b110 6
#121090000000
1!
1%
1-
12
#121100000000
0!
0%
b111 *
0-
02
b111 6
#121110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#121120000000
0!
0%
b0 *
0-
02
b0 6
#121130000000
1!
1%
1-
12
#121140000000
0!
0%
b1 *
0-
02
b1 6
#121150000000
1!
1%
1-
12
#121160000000
0!
0%
b10 *
0-
02
b10 6
#121170000000
1!
1%
1-
12
#121180000000
0!
0%
b11 *
0-
02
b11 6
#121190000000
1!
1%
1-
12
15
#121200000000
0!
0%
b100 *
0-
02
b100 6
#121210000000
1!
1%
1-
12
#121220000000
0!
0%
b101 *
0-
02
b101 6
#121230000000
1!
1%
1-
12
#121240000000
0!
0%
b110 *
0-
02
b110 6
#121250000000
1!
1%
1-
12
#121260000000
0!
0%
b111 *
0-
02
b111 6
#121270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#121280000000
0!
0%
b0 *
0-
02
b0 6
#121290000000
1!
1%
1-
12
#121300000000
0!
0%
b1 *
0-
02
b1 6
#121310000000
1!
1%
1-
12
#121320000000
0!
0%
b10 *
0-
02
b10 6
#121330000000
1!
1%
1-
12
#121340000000
0!
0%
b11 *
0-
02
b11 6
#121350000000
1!
1%
1-
12
15
#121360000000
0!
0%
b100 *
0-
02
b100 6
#121370000000
1!
1%
1-
12
#121380000000
0!
0%
b101 *
0-
02
b101 6
#121390000000
1!
1%
1-
12
#121400000000
0!
0%
b110 *
0-
02
b110 6
#121410000000
1!
1%
1-
12
#121420000000
0!
0%
b111 *
0-
02
b111 6
#121430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#121440000000
0!
0%
b0 *
0-
02
b0 6
#121450000000
1!
1%
1-
12
#121460000000
0!
0%
b1 *
0-
02
b1 6
#121470000000
1!
1%
1-
12
#121480000000
0!
0%
b10 *
0-
02
b10 6
#121490000000
1!
1%
1-
12
#121500000000
0!
0%
b11 *
0-
02
b11 6
#121510000000
1!
1%
1-
12
15
#121520000000
0!
0%
b100 *
0-
02
b100 6
#121530000000
1!
1%
1-
12
#121540000000
0!
0%
b101 *
0-
02
b101 6
#121550000000
1!
1%
1-
12
#121560000000
0!
0%
b110 *
0-
02
b110 6
#121570000000
1!
1%
1-
12
#121580000000
0!
0%
b111 *
0-
02
b111 6
#121590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#121600000000
0!
0%
b0 *
0-
02
b0 6
#121610000000
1!
1%
1-
12
#121620000000
0!
0%
b1 *
0-
02
b1 6
#121630000000
1!
1%
1-
12
#121640000000
0!
0%
b10 *
0-
02
b10 6
#121650000000
1!
1%
1-
12
#121660000000
0!
0%
b11 *
0-
02
b11 6
#121670000000
1!
1%
1-
12
15
#121680000000
0!
0%
b100 *
0-
02
b100 6
#121690000000
1!
1%
1-
12
#121700000000
0!
0%
b101 *
0-
02
b101 6
#121710000000
1!
1%
1-
12
#121720000000
0!
0%
b110 *
0-
02
b110 6
#121730000000
1!
1%
1-
12
#121740000000
0!
0%
b111 *
0-
02
b111 6
#121750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#121760000000
0!
0%
b0 *
0-
02
b0 6
#121770000000
1!
1%
1-
12
#121780000000
0!
0%
b1 *
0-
02
b1 6
#121790000000
1!
1%
1-
12
#121800000000
0!
0%
b10 *
0-
02
b10 6
#121810000000
1!
1%
1-
12
#121820000000
0!
0%
b11 *
0-
02
b11 6
#121830000000
1!
1%
1-
12
15
#121840000000
0!
0%
b100 *
0-
02
b100 6
#121850000000
1!
1%
1-
12
#121860000000
0!
0%
b101 *
0-
02
b101 6
#121870000000
1!
1%
1-
12
#121880000000
0!
0%
b110 *
0-
02
b110 6
#121890000000
1!
1%
1-
12
#121900000000
0!
0%
b111 *
0-
02
b111 6
#121910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#121920000000
0!
0%
b0 *
0-
02
b0 6
#121930000000
1!
1%
1-
12
#121940000000
0!
0%
b1 *
0-
02
b1 6
#121950000000
1!
1%
1-
12
#121960000000
0!
0%
b10 *
0-
02
b10 6
#121970000000
1!
1%
1-
12
#121980000000
0!
0%
b11 *
0-
02
b11 6
#121990000000
1!
1%
1-
12
15
#122000000000
0!
0%
b100 *
0-
02
b100 6
#122010000000
1!
1%
1-
12
#122020000000
0!
0%
b101 *
0-
02
b101 6
#122030000000
1!
1%
1-
12
#122040000000
0!
0%
b110 *
0-
02
b110 6
#122050000000
1!
1%
1-
12
#122060000000
0!
0%
b111 *
0-
02
b111 6
#122070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#122080000000
0!
0%
b0 *
0-
02
b0 6
#122090000000
1!
1%
1-
12
#122100000000
0!
0%
b1 *
0-
02
b1 6
#122110000000
1!
1%
1-
12
#122120000000
0!
0%
b10 *
0-
02
b10 6
#122130000000
1!
1%
1-
12
#122140000000
0!
0%
b11 *
0-
02
b11 6
#122150000000
1!
1%
1-
12
15
#122160000000
0!
0%
b100 *
0-
02
b100 6
#122170000000
1!
1%
1-
12
#122180000000
0!
0%
b101 *
0-
02
b101 6
#122190000000
1!
1%
1-
12
#122200000000
0!
0%
b110 *
0-
02
b110 6
#122210000000
1!
1%
1-
12
#122220000000
0!
0%
b111 *
0-
02
b111 6
#122230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#122240000000
0!
0%
b0 *
0-
02
b0 6
#122250000000
1!
1%
1-
12
#122260000000
0!
0%
b1 *
0-
02
b1 6
#122270000000
1!
1%
1-
12
#122280000000
0!
0%
b10 *
0-
02
b10 6
#122290000000
1!
1%
1-
12
#122300000000
0!
0%
b11 *
0-
02
b11 6
#122310000000
1!
1%
1-
12
15
#122320000000
0!
0%
b100 *
0-
02
b100 6
#122330000000
1!
1%
1-
12
#122340000000
0!
0%
b101 *
0-
02
b101 6
#122350000000
1!
1%
1-
12
#122360000000
0!
0%
b110 *
0-
02
b110 6
#122370000000
1!
1%
1-
12
#122380000000
0!
0%
b111 *
0-
02
b111 6
#122390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#122400000000
0!
0%
b0 *
0-
02
b0 6
#122410000000
1!
1%
1-
12
#122420000000
0!
0%
b1 *
0-
02
b1 6
#122430000000
1!
1%
1-
12
#122440000000
0!
0%
b10 *
0-
02
b10 6
#122450000000
1!
1%
1-
12
#122460000000
0!
0%
b11 *
0-
02
b11 6
#122470000000
1!
1%
1-
12
15
#122480000000
0!
0%
b100 *
0-
02
b100 6
#122490000000
1!
1%
1-
12
#122500000000
0!
0%
b101 *
0-
02
b101 6
#122510000000
1!
1%
1-
12
#122520000000
0!
0%
b110 *
0-
02
b110 6
#122530000000
1!
1%
1-
12
#122540000000
0!
0%
b111 *
0-
02
b111 6
#122550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#122560000000
0!
0%
b0 *
0-
02
b0 6
#122570000000
1!
1%
1-
12
#122580000000
0!
0%
b1 *
0-
02
b1 6
#122590000000
1!
1%
1-
12
#122600000000
0!
0%
b10 *
0-
02
b10 6
#122610000000
1!
1%
1-
12
#122620000000
0!
0%
b11 *
0-
02
b11 6
#122630000000
1!
1%
1-
12
15
#122640000000
0!
0%
b100 *
0-
02
b100 6
#122650000000
1!
1%
1-
12
#122660000000
0!
0%
b101 *
0-
02
b101 6
#122670000000
1!
1%
1-
12
#122680000000
0!
0%
b110 *
0-
02
b110 6
#122690000000
1!
1%
1-
12
#122700000000
0!
0%
b111 *
0-
02
b111 6
#122710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#122720000000
0!
0%
b0 *
0-
02
b0 6
#122730000000
1!
1%
1-
12
#122740000000
0!
0%
b1 *
0-
02
b1 6
#122750000000
1!
1%
1-
12
#122760000000
0!
0%
b10 *
0-
02
b10 6
#122770000000
1!
1%
1-
12
#122780000000
0!
0%
b11 *
0-
02
b11 6
#122790000000
1!
1%
1-
12
15
#122800000000
0!
0%
b100 *
0-
02
b100 6
#122810000000
1!
1%
1-
12
#122820000000
0!
0%
b101 *
0-
02
b101 6
#122830000000
1!
1%
1-
12
#122840000000
0!
0%
b110 *
0-
02
b110 6
#122850000000
1!
1%
1-
12
#122860000000
0!
0%
b111 *
0-
02
b111 6
#122870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#122880000000
0!
0%
b0 *
0-
02
b0 6
#122890000000
1!
1%
1-
12
#122900000000
0!
0%
b1 *
0-
02
b1 6
#122910000000
1!
1%
1-
12
#122920000000
0!
0%
b10 *
0-
02
b10 6
#122930000000
1!
1%
1-
12
#122940000000
0!
0%
b11 *
0-
02
b11 6
#122950000000
1!
1%
1-
12
15
#122960000000
0!
0%
b100 *
0-
02
b100 6
#122970000000
1!
1%
1-
12
#122980000000
0!
0%
b101 *
0-
02
b101 6
#122990000000
1!
1%
1-
12
#123000000000
0!
0%
b110 *
0-
02
b110 6
#123010000000
1!
1%
1-
12
#123020000000
0!
0%
b111 *
0-
02
b111 6
#123030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#123040000000
0!
0%
b0 *
0-
02
b0 6
#123050000000
1!
1%
1-
12
#123060000000
0!
0%
b1 *
0-
02
b1 6
#123070000000
1!
1%
1-
12
#123080000000
0!
0%
b10 *
0-
02
b10 6
#123090000000
1!
1%
1-
12
#123100000000
0!
0%
b11 *
0-
02
b11 6
#123110000000
1!
1%
1-
12
15
#123120000000
0!
0%
b100 *
0-
02
b100 6
#123130000000
1!
1%
1-
12
#123140000000
0!
0%
b101 *
0-
02
b101 6
#123150000000
1!
1%
1-
12
#123160000000
0!
0%
b110 *
0-
02
b110 6
#123170000000
1!
1%
1-
12
#123180000000
0!
0%
b111 *
0-
02
b111 6
#123190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#123200000000
0!
0%
b0 *
0-
02
b0 6
#123210000000
1!
1%
1-
12
#123220000000
0!
0%
b1 *
0-
02
b1 6
#123230000000
1!
1%
1-
12
#123240000000
0!
0%
b10 *
0-
02
b10 6
#123250000000
1!
1%
1-
12
#123260000000
0!
0%
b11 *
0-
02
b11 6
#123270000000
1!
1%
1-
12
15
#123280000000
0!
0%
b100 *
0-
02
b100 6
#123290000000
1!
1%
1-
12
#123300000000
0!
0%
b101 *
0-
02
b101 6
#123310000000
1!
1%
1-
12
#123320000000
0!
0%
b110 *
0-
02
b110 6
#123330000000
1!
1%
1-
12
#123340000000
0!
0%
b111 *
0-
02
b111 6
#123350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#123360000000
0!
0%
b0 *
0-
02
b0 6
#123370000000
1!
1%
1-
12
#123380000000
0!
0%
b1 *
0-
02
b1 6
#123390000000
1!
1%
1-
12
#123400000000
0!
0%
b10 *
0-
02
b10 6
#123410000000
1!
1%
1-
12
#123420000000
0!
0%
b11 *
0-
02
b11 6
#123430000000
1!
1%
1-
12
15
#123440000000
0!
0%
b100 *
0-
02
b100 6
#123450000000
1!
1%
1-
12
#123460000000
0!
0%
b101 *
0-
02
b101 6
#123470000000
1!
1%
1-
12
#123480000000
0!
0%
b110 *
0-
02
b110 6
#123490000000
1!
1%
1-
12
#123500000000
0!
0%
b111 *
0-
02
b111 6
#123510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#123520000000
0!
0%
b0 *
0-
02
b0 6
#123530000000
1!
1%
1-
12
#123540000000
0!
0%
b1 *
0-
02
b1 6
#123550000000
1!
1%
1-
12
#123560000000
0!
0%
b10 *
0-
02
b10 6
#123570000000
1!
1%
1-
12
#123580000000
0!
0%
b11 *
0-
02
b11 6
#123590000000
1!
1%
1-
12
15
#123600000000
0!
0%
b100 *
0-
02
b100 6
#123610000000
1!
1%
1-
12
#123620000000
0!
0%
b101 *
0-
02
b101 6
#123630000000
1!
1%
1-
12
#123640000000
0!
0%
b110 *
0-
02
b110 6
#123650000000
1!
1%
1-
12
#123660000000
0!
0%
b111 *
0-
02
b111 6
#123670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#123680000000
0!
0%
b0 *
0-
02
b0 6
#123690000000
1!
1%
1-
12
#123700000000
0!
0%
b1 *
0-
02
b1 6
#123710000000
1!
1%
1-
12
#123720000000
0!
0%
b10 *
0-
02
b10 6
#123730000000
1!
1%
1-
12
#123740000000
0!
0%
b11 *
0-
02
b11 6
#123750000000
1!
1%
1-
12
15
#123760000000
0!
0%
b100 *
0-
02
b100 6
#123770000000
1!
1%
1-
12
#123780000000
0!
0%
b101 *
0-
02
b101 6
#123790000000
1!
1%
1-
12
#123800000000
0!
0%
b110 *
0-
02
b110 6
#123810000000
1!
1%
1-
12
#123820000000
0!
0%
b111 *
0-
02
b111 6
#123830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#123840000000
0!
0%
b0 *
0-
02
b0 6
#123850000000
1!
1%
1-
12
#123860000000
0!
0%
b1 *
0-
02
b1 6
#123870000000
1!
1%
1-
12
#123880000000
0!
0%
b10 *
0-
02
b10 6
#123890000000
1!
1%
1-
12
#123900000000
0!
0%
b11 *
0-
02
b11 6
#123910000000
1!
1%
1-
12
15
#123920000000
0!
0%
b100 *
0-
02
b100 6
#123930000000
1!
1%
1-
12
#123940000000
0!
0%
b101 *
0-
02
b101 6
#123950000000
1!
1%
1-
12
#123960000000
0!
0%
b110 *
0-
02
b110 6
#123970000000
1!
1%
1-
12
#123980000000
0!
0%
b111 *
0-
02
b111 6
#123990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#124000000000
0!
0%
b0 *
0-
02
b0 6
#124010000000
1!
1%
1-
12
#124020000000
0!
0%
b1 *
0-
02
b1 6
#124030000000
1!
1%
1-
12
#124040000000
0!
0%
b10 *
0-
02
b10 6
#124050000000
1!
1%
1-
12
#124060000000
0!
0%
b11 *
0-
02
b11 6
#124070000000
1!
1%
1-
12
15
#124080000000
0!
0%
b100 *
0-
02
b100 6
#124090000000
1!
1%
1-
12
#124100000000
0!
0%
b101 *
0-
02
b101 6
#124110000000
1!
1%
1-
12
#124120000000
0!
0%
b110 *
0-
02
b110 6
#124130000000
1!
1%
1-
12
#124140000000
0!
0%
b111 *
0-
02
b111 6
#124150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#124160000000
0!
0%
b0 *
0-
02
b0 6
#124170000000
1!
1%
1-
12
#124180000000
0!
0%
b1 *
0-
02
b1 6
#124190000000
1!
1%
1-
12
#124200000000
0!
0%
b10 *
0-
02
b10 6
#124210000000
1!
1%
1-
12
#124220000000
0!
0%
b11 *
0-
02
b11 6
#124230000000
1!
1%
1-
12
15
#124240000000
0!
0%
b100 *
0-
02
b100 6
#124250000000
1!
1%
1-
12
#124260000000
0!
0%
b101 *
0-
02
b101 6
#124270000000
1!
1%
1-
12
#124280000000
0!
0%
b110 *
0-
02
b110 6
#124290000000
1!
1%
1-
12
#124300000000
0!
0%
b111 *
0-
02
b111 6
#124310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#124320000000
0!
0%
b0 *
0-
02
b0 6
#124330000000
1!
1%
1-
12
#124340000000
0!
0%
b1 *
0-
02
b1 6
#124350000000
1!
1%
1-
12
#124360000000
0!
0%
b10 *
0-
02
b10 6
#124370000000
1!
1%
1-
12
#124380000000
0!
0%
b11 *
0-
02
b11 6
#124390000000
1!
1%
1-
12
15
#124400000000
0!
0%
b100 *
0-
02
b100 6
#124410000000
1!
1%
1-
12
#124420000000
0!
0%
b101 *
0-
02
b101 6
#124430000000
1!
1%
1-
12
#124440000000
0!
0%
b110 *
0-
02
b110 6
#124450000000
1!
1%
1-
12
#124460000000
0!
0%
b111 *
0-
02
b111 6
#124470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#124480000000
0!
0%
b0 *
0-
02
b0 6
#124490000000
1!
1%
1-
12
#124500000000
0!
0%
b1 *
0-
02
b1 6
#124510000000
1!
1%
1-
12
#124520000000
0!
0%
b10 *
0-
02
b10 6
#124530000000
1!
1%
1-
12
#124540000000
0!
0%
b11 *
0-
02
b11 6
#124550000000
1!
1%
1-
12
15
#124560000000
0!
0%
b100 *
0-
02
b100 6
#124570000000
1!
1%
1-
12
#124580000000
0!
0%
b101 *
0-
02
b101 6
#124590000000
1!
1%
1-
12
#124600000000
0!
0%
b110 *
0-
02
b110 6
#124610000000
1!
1%
1-
12
#124620000000
0!
0%
b111 *
0-
02
b111 6
#124630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#124640000000
0!
0%
b0 *
0-
02
b0 6
#124650000000
1!
1%
1-
12
#124660000000
0!
0%
b1 *
0-
02
b1 6
#124670000000
1!
1%
1-
12
#124680000000
0!
0%
b10 *
0-
02
b10 6
#124690000000
1!
1%
1-
12
#124700000000
0!
0%
b11 *
0-
02
b11 6
#124710000000
1!
1%
1-
12
15
#124720000000
0!
0%
b100 *
0-
02
b100 6
#124730000000
1!
1%
1-
12
#124740000000
0!
0%
b101 *
0-
02
b101 6
#124750000000
1!
1%
1-
12
#124760000000
0!
0%
b110 *
0-
02
b110 6
#124770000000
1!
1%
1-
12
#124780000000
0!
0%
b111 *
0-
02
b111 6
#124790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#124800000000
0!
0%
b0 *
0-
02
b0 6
#124810000000
1!
1%
1-
12
#124820000000
0!
0%
b1 *
0-
02
b1 6
#124830000000
1!
1%
1-
12
#124840000000
0!
0%
b10 *
0-
02
b10 6
#124850000000
1!
1%
1-
12
#124860000000
0!
0%
b11 *
0-
02
b11 6
#124870000000
1!
1%
1-
12
15
#124880000000
0!
0%
b100 *
0-
02
b100 6
#124890000000
1!
1%
1-
12
#124900000000
0!
0%
b101 *
0-
02
b101 6
#124910000000
1!
1%
1-
12
#124920000000
0!
0%
b110 *
0-
02
b110 6
#124930000000
1!
1%
1-
12
#124940000000
0!
0%
b111 *
0-
02
b111 6
#124950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#124960000000
0!
0%
b0 *
0-
02
b0 6
#124970000000
1!
1%
1-
12
#124980000000
0!
0%
b1 *
0-
02
b1 6
#124990000000
1!
1%
1-
12
#125000000000
0!
0%
b10 *
0-
02
b10 6
#125010000000
1!
1%
1-
12
#125020000000
0!
0%
b11 *
0-
02
b11 6
#125030000000
1!
1%
1-
12
15
#125040000000
0!
0%
b100 *
0-
02
b100 6
#125050000000
1!
1%
1-
12
#125060000000
0!
0%
b101 *
0-
02
b101 6
#125070000000
1!
1%
1-
12
#125080000000
0!
0%
b110 *
0-
02
b110 6
#125090000000
1!
1%
1-
12
#125100000000
0!
0%
b111 *
0-
02
b111 6
#125110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#125120000000
0!
0%
b0 *
0-
02
b0 6
#125130000000
1!
1%
1-
12
#125140000000
0!
0%
b1 *
0-
02
b1 6
#125150000000
1!
1%
1-
12
#125160000000
0!
0%
b10 *
0-
02
b10 6
#125170000000
1!
1%
1-
12
#125180000000
0!
0%
b11 *
0-
02
b11 6
#125190000000
1!
1%
1-
12
15
#125200000000
0!
0%
b100 *
0-
02
b100 6
#125210000000
1!
1%
1-
12
#125220000000
0!
0%
b101 *
0-
02
b101 6
#125230000000
1!
1%
1-
12
#125240000000
0!
0%
b110 *
0-
02
b110 6
#125250000000
1!
1%
1-
12
#125260000000
0!
0%
b111 *
0-
02
b111 6
#125270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#125280000000
0!
0%
b0 *
0-
02
b0 6
#125290000000
1!
1%
1-
12
#125300000000
0!
0%
b1 *
0-
02
b1 6
#125310000000
1!
1%
1-
12
#125320000000
0!
0%
b10 *
0-
02
b10 6
#125330000000
1!
1%
1-
12
#125340000000
0!
0%
b11 *
0-
02
b11 6
#125350000000
1!
1%
1-
12
15
#125360000000
0!
0%
b100 *
0-
02
b100 6
#125370000000
1!
1%
1-
12
#125380000000
0!
0%
b101 *
0-
02
b101 6
#125390000000
1!
1%
1-
12
#125400000000
0!
0%
b110 *
0-
02
b110 6
#125410000000
1!
1%
1-
12
#125420000000
0!
0%
b111 *
0-
02
b111 6
#125430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#125440000000
0!
0%
b0 *
0-
02
b0 6
#125450000000
1!
1%
1-
12
#125460000000
0!
0%
b1 *
0-
02
b1 6
#125470000000
1!
1%
1-
12
#125480000000
0!
0%
b10 *
0-
02
b10 6
#125490000000
1!
1%
1-
12
#125500000000
0!
0%
b11 *
0-
02
b11 6
#125510000000
1!
1%
1-
12
15
#125520000000
0!
0%
b100 *
0-
02
b100 6
#125530000000
1!
1%
1-
12
#125540000000
0!
0%
b101 *
0-
02
b101 6
#125550000000
1!
1%
1-
12
#125560000000
0!
0%
b110 *
0-
02
b110 6
#125570000000
1!
1%
1-
12
#125580000000
0!
0%
b111 *
0-
02
b111 6
#125590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#125600000000
0!
0%
b0 *
0-
02
b0 6
#125610000000
1!
1%
1-
12
#125620000000
0!
0%
b1 *
0-
02
b1 6
#125630000000
1!
1%
1-
12
#125640000000
0!
0%
b10 *
0-
02
b10 6
#125650000000
1!
1%
1-
12
#125660000000
0!
0%
b11 *
0-
02
b11 6
#125670000000
1!
1%
1-
12
15
#125680000000
0!
0%
b100 *
0-
02
b100 6
#125690000000
1!
1%
1-
12
#125700000000
0!
0%
b101 *
0-
02
b101 6
#125710000000
1!
1%
1-
12
#125720000000
0!
0%
b110 *
0-
02
b110 6
#125730000000
1!
1%
1-
12
#125740000000
0!
0%
b111 *
0-
02
b111 6
#125750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#125760000000
0!
0%
b0 *
0-
02
b0 6
#125770000000
1!
1%
1-
12
#125780000000
0!
0%
b1 *
0-
02
b1 6
#125790000000
1!
1%
1-
12
#125800000000
0!
0%
b10 *
0-
02
b10 6
#125810000000
1!
1%
1-
12
#125820000000
0!
0%
b11 *
0-
02
b11 6
#125830000000
1!
1%
1-
12
15
#125840000000
0!
0%
b100 *
0-
02
b100 6
#125850000000
1!
1%
1-
12
#125860000000
0!
0%
b101 *
0-
02
b101 6
#125870000000
1!
1%
1-
12
#125880000000
0!
0%
b110 *
0-
02
b110 6
#125890000000
1!
1%
1-
12
#125900000000
0!
0%
b111 *
0-
02
b111 6
#125910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#125920000000
0!
0%
b0 *
0-
02
b0 6
#125930000000
1!
1%
1-
12
#125940000000
0!
0%
b1 *
0-
02
b1 6
#125950000000
1!
1%
1-
12
#125960000000
0!
0%
b10 *
0-
02
b10 6
#125970000000
1!
1%
1-
12
#125980000000
0!
0%
b11 *
0-
02
b11 6
#125990000000
1!
1%
1-
12
15
#126000000000
0!
0%
b100 *
0-
02
b100 6
#126010000000
1!
1%
1-
12
#126020000000
0!
0%
b101 *
0-
02
b101 6
#126030000000
1!
1%
1-
12
#126040000000
0!
0%
b110 *
0-
02
b110 6
#126050000000
1!
1%
1-
12
#126060000000
0!
0%
b111 *
0-
02
b111 6
#126070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#126080000000
0!
0%
b0 *
0-
02
b0 6
#126090000000
1!
1%
1-
12
#126100000000
0!
0%
b1 *
0-
02
b1 6
#126110000000
1!
1%
1-
12
#126120000000
0!
0%
b10 *
0-
02
b10 6
#126130000000
1!
1%
1-
12
#126140000000
0!
0%
b11 *
0-
02
b11 6
#126150000000
1!
1%
1-
12
15
#126160000000
0!
0%
b100 *
0-
02
b100 6
#126170000000
1!
1%
1-
12
#126180000000
0!
0%
b101 *
0-
02
b101 6
#126190000000
1!
1%
1-
12
#126200000000
0!
0%
b110 *
0-
02
b110 6
#126210000000
1!
1%
1-
12
#126220000000
0!
0%
b111 *
0-
02
b111 6
#126230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#126240000000
0!
0%
b0 *
0-
02
b0 6
#126250000000
1!
1%
1-
12
#126260000000
0!
0%
b1 *
0-
02
b1 6
#126270000000
1!
1%
1-
12
#126280000000
0!
0%
b10 *
0-
02
b10 6
#126290000000
1!
1%
1-
12
#126300000000
0!
0%
b11 *
0-
02
b11 6
#126310000000
1!
1%
1-
12
15
#126320000000
0!
0%
b100 *
0-
02
b100 6
#126330000000
1!
1%
1-
12
#126340000000
0!
0%
b101 *
0-
02
b101 6
#126350000000
1!
1%
1-
12
#126360000000
0!
0%
b110 *
0-
02
b110 6
#126370000000
1!
1%
1-
12
#126380000000
0!
0%
b111 *
0-
02
b111 6
#126390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#126400000000
0!
0%
b0 *
0-
02
b0 6
#126410000000
1!
1%
1-
12
#126420000000
0!
0%
b1 *
0-
02
b1 6
#126430000000
1!
1%
1-
12
#126440000000
0!
0%
b10 *
0-
02
b10 6
#126450000000
1!
1%
1-
12
#126460000000
0!
0%
b11 *
0-
02
b11 6
#126470000000
1!
1%
1-
12
15
#126480000000
0!
0%
b100 *
0-
02
b100 6
#126490000000
1!
1%
1-
12
#126500000000
0!
0%
b101 *
0-
02
b101 6
#126510000000
1!
1%
1-
12
#126520000000
0!
0%
b110 *
0-
02
b110 6
#126530000000
1!
1%
1-
12
#126540000000
0!
0%
b111 *
0-
02
b111 6
#126550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#126560000000
0!
0%
b0 *
0-
02
b0 6
#126570000000
1!
1%
1-
12
#126580000000
0!
0%
b1 *
0-
02
b1 6
#126590000000
1!
1%
1-
12
#126600000000
0!
0%
b10 *
0-
02
b10 6
#126610000000
1!
1%
1-
12
#126620000000
0!
0%
b11 *
0-
02
b11 6
#126630000000
1!
1%
1-
12
15
#126640000000
0!
0%
b100 *
0-
02
b100 6
#126650000000
1!
1%
1-
12
#126660000000
0!
0%
b101 *
0-
02
b101 6
#126670000000
1!
1%
1-
12
#126680000000
0!
0%
b110 *
0-
02
b110 6
#126690000000
1!
1%
1-
12
#126700000000
0!
0%
b111 *
0-
02
b111 6
#126710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#126720000000
0!
0%
b0 *
0-
02
b0 6
#126730000000
1!
1%
1-
12
#126740000000
0!
0%
b1 *
0-
02
b1 6
#126750000000
1!
1%
1-
12
#126760000000
0!
0%
b10 *
0-
02
b10 6
#126770000000
1!
1%
1-
12
#126780000000
0!
0%
b11 *
0-
02
b11 6
#126790000000
1!
1%
1-
12
15
#126800000000
0!
0%
b100 *
0-
02
b100 6
#126810000000
1!
1%
1-
12
#126820000000
0!
0%
b101 *
0-
02
b101 6
#126830000000
1!
1%
1-
12
#126840000000
0!
0%
b110 *
0-
02
b110 6
#126850000000
1!
1%
1-
12
#126860000000
0!
0%
b111 *
0-
02
b111 6
#126870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#126880000000
0!
0%
b0 *
0-
02
b0 6
#126890000000
1!
1%
1-
12
#126900000000
0!
0%
b1 *
0-
02
b1 6
#126910000000
1!
1%
1-
12
#126920000000
0!
0%
b10 *
0-
02
b10 6
#126930000000
1!
1%
1-
12
#126940000000
0!
0%
b11 *
0-
02
b11 6
#126950000000
1!
1%
1-
12
15
#126960000000
0!
0%
b100 *
0-
02
b100 6
#126970000000
1!
1%
1-
12
#126980000000
0!
0%
b101 *
0-
02
b101 6
#126990000000
1!
1%
1-
12
#127000000000
0!
0%
b110 *
0-
02
b110 6
#127010000000
1!
1%
1-
12
#127020000000
0!
0%
b111 *
0-
02
b111 6
#127030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#127040000000
0!
0%
b0 *
0-
02
b0 6
#127050000000
1!
1%
1-
12
#127060000000
0!
0%
b1 *
0-
02
b1 6
#127070000000
1!
1%
1-
12
#127080000000
0!
0%
b10 *
0-
02
b10 6
#127090000000
1!
1%
1-
12
#127100000000
0!
0%
b11 *
0-
02
b11 6
#127110000000
1!
1%
1-
12
15
#127120000000
0!
0%
b100 *
0-
02
b100 6
#127130000000
1!
1%
1-
12
#127140000000
0!
0%
b101 *
0-
02
b101 6
#127150000000
1!
1%
1-
12
#127160000000
0!
0%
b110 *
0-
02
b110 6
#127170000000
1!
1%
1-
12
#127180000000
0!
0%
b111 *
0-
02
b111 6
#127190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#127200000000
0!
0%
b0 *
0-
02
b0 6
#127210000000
1!
1%
1-
12
#127220000000
0!
0%
b1 *
0-
02
b1 6
#127230000000
1!
1%
1-
12
#127240000000
0!
0%
b10 *
0-
02
b10 6
#127250000000
1!
1%
1-
12
#127260000000
0!
0%
b11 *
0-
02
b11 6
#127270000000
1!
1%
1-
12
15
#127280000000
0!
0%
b100 *
0-
02
b100 6
#127290000000
1!
1%
1-
12
#127300000000
0!
0%
b101 *
0-
02
b101 6
#127310000000
1!
1%
1-
12
#127320000000
0!
0%
b110 *
0-
02
b110 6
#127330000000
1!
1%
1-
12
#127340000000
0!
0%
b111 *
0-
02
b111 6
#127350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#127360000000
0!
0%
b0 *
0-
02
b0 6
#127370000000
1!
1%
1-
12
#127380000000
0!
0%
b1 *
0-
02
b1 6
#127390000000
1!
1%
1-
12
#127400000000
0!
0%
b10 *
0-
02
b10 6
#127410000000
1!
1%
1-
12
#127420000000
0!
0%
b11 *
0-
02
b11 6
#127430000000
1!
1%
1-
12
15
#127440000000
0!
0%
b100 *
0-
02
b100 6
#127450000000
1!
1%
1-
12
#127460000000
0!
0%
b101 *
0-
02
b101 6
#127470000000
1!
1%
1-
12
#127480000000
0!
0%
b110 *
0-
02
b110 6
#127490000000
1!
1%
1-
12
#127500000000
0!
0%
b111 *
0-
02
b111 6
#127510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#127520000000
0!
0%
b0 *
0-
02
b0 6
#127530000000
1!
1%
1-
12
#127540000000
0!
0%
b1 *
0-
02
b1 6
#127550000000
1!
1%
1-
12
#127560000000
0!
0%
b10 *
0-
02
b10 6
#127570000000
1!
1%
1-
12
#127580000000
0!
0%
b11 *
0-
02
b11 6
#127590000000
1!
1%
1-
12
15
#127600000000
0!
0%
b100 *
0-
02
b100 6
#127610000000
1!
1%
1-
12
#127620000000
0!
0%
b101 *
0-
02
b101 6
#127630000000
1!
1%
1-
12
#127640000000
0!
0%
b110 *
0-
02
b110 6
#127650000000
1!
1%
1-
12
#127660000000
0!
0%
b111 *
0-
02
b111 6
#127670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#127680000000
0!
0%
b0 *
0-
02
b0 6
#127690000000
1!
1%
1-
12
#127700000000
0!
0%
b1 *
0-
02
b1 6
#127710000000
1!
1%
1-
12
#127720000000
0!
0%
b10 *
0-
02
b10 6
#127730000000
1!
1%
1-
12
#127740000000
0!
0%
b11 *
0-
02
b11 6
#127750000000
1!
1%
1-
12
15
#127760000000
0!
0%
b100 *
0-
02
b100 6
#127770000000
1!
1%
1-
12
#127780000000
0!
0%
b101 *
0-
02
b101 6
#127790000000
1!
1%
1-
12
#127800000000
0!
0%
b110 *
0-
02
b110 6
#127810000000
1!
1%
1-
12
#127820000000
0!
0%
b111 *
0-
02
b111 6
#127830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#127840000000
0!
0%
b0 *
0-
02
b0 6
#127850000000
1!
1%
1-
12
#127860000000
0!
0%
b1 *
0-
02
b1 6
#127870000000
1!
1%
1-
12
#127880000000
0!
0%
b10 *
0-
02
b10 6
#127890000000
1!
1%
1-
12
#127900000000
0!
0%
b11 *
0-
02
b11 6
#127910000000
1!
1%
1-
12
15
#127920000000
0!
0%
b100 *
0-
02
b100 6
#127930000000
1!
1%
1-
12
#127940000000
0!
0%
b101 *
0-
02
b101 6
#127950000000
1!
1%
1-
12
#127960000000
0!
0%
b110 *
0-
02
b110 6
#127970000000
1!
1%
1-
12
#127980000000
0!
0%
b111 *
0-
02
b111 6
#127990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#128000000000
0!
0%
b0 *
0-
02
b0 6
#128010000000
1!
1%
1-
12
#128020000000
0!
0%
b1 *
0-
02
b1 6
#128030000000
1!
1%
1-
12
#128040000000
0!
0%
b10 *
0-
02
b10 6
#128050000000
1!
1%
1-
12
#128060000000
0!
0%
b11 *
0-
02
b11 6
#128070000000
1!
1%
1-
12
15
#128080000000
0!
0%
b100 *
0-
02
b100 6
#128090000000
1!
1%
1-
12
#128100000000
0!
0%
b101 *
0-
02
b101 6
#128110000000
1!
1%
1-
12
#128120000000
0!
0%
b110 *
0-
02
b110 6
#128130000000
1!
1%
1-
12
#128140000000
0!
0%
b111 *
0-
02
b111 6
#128150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#128160000000
0!
0%
b0 *
0-
02
b0 6
#128170000000
1!
1%
1-
12
#128180000000
0!
0%
b1 *
0-
02
b1 6
#128190000000
1!
1%
1-
12
#128200000000
0!
0%
b10 *
0-
02
b10 6
#128210000000
1!
1%
1-
12
#128220000000
0!
0%
b11 *
0-
02
b11 6
#128230000000
1!
1%
1-
12
15
#128240000000
0!
0%
b100 *
0-
02
b100 6
#128250000000
1!
1%
1-
12
#128260000000
0!
0%
b101 *
0-
02
b101 6
#128270000000
1!
1%
1-
12
#128280000000
0!
0%
b110 *
0-
02
b110 6
#128290000000
1!
1%
1-
12
#128300000000
0!
0%
b111 *
0-
02
b111 6
#128310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#128320000000
0!
0%
b0 *
0-
02
b0 6
#128330000000
1!
1%
1-
12
#128340000000
0!
0%
b1 *
0-
02
b1 6
#128350000000
1!
1%
1-
12
#128360000000
0!
0%
b10 *
0-
02
b10 6
#128370000000
1!
1%
1-
12
#128380000000
0!
0%
b11 *
0-
02
b11 6
#128390000000
1!
1%
1-
12
15
#128400000000
0!
0%
b100 *
0-
02
b100 6
#128410000000
1!
1%
1-
12
#128420000000
0!
0%
b101 *
0-
02
b101 6
#128430000000
1!
1%
1-
12
#128440000000
0!
0%
b110 *
0-
02
b110 6
#128450000000
1!
1%
1-
12
#128460000000
0!
0%
b111 *
0-
02
b111 6
#128470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#128480000000
0!
0%
b0 *
0-
02
b0 6
#128490000000
1!
1%
1-
12
#128500000000
0!
0%
b1 *
0-
02
b1 6
#128510000000
1!
1%
1-
12
#128520000000
0!
0%
b10 *
0-
02
b10 6
#128530000000
1!
1%
1-
12
#128540000000
0!
0%
b11 *
0-
02
b11 6
#128550000000
1!
1%
1-
12
15
#128560000000
0!
0%
b100 *
0-
02
b100 6
#128570000000
1!
1%
1-
12
#128580000000
0!
0%
b101 *
0-
02
b101 6
#128590000000
1!
1%
1-
12
#128600000000
0!
0%
b110 *
0-
02
b110 6
#128610000000
1!
1%
1-
12
#128620000000
0!
0%
b111 *
0-
02
b111 6
#128630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#128640000000
0!
0%
b0 *
0-
02
b0 6
#128650000000
1!
1%
1-
12
#128660000000
0!
0%
b1 *
0-
02
b1 6
#128670000000
1!
1%
1-
12
#128680000000
0!
0%
b10 *
0-
02
b10 6
#128690000000
1!
1%
1-
12
#128700000000
0!
0%
b11 *
0-
02
b11 6
#128710000000
1!
1%
1-
12
15
#128720000000
0!
0%
b100 *
0-
02
b100 6
#128730000000
1!
1%
1-
12
#128740000000
0!
0%
b101 *
0-
02
b101 6
#128750000000
1!
1%
1-
12
#128760000000
0!
0%
b110 *
0-
02
b110 6
#128770000000
1!
1%
1-
12
#128780000000
0!
0%
b111 *
0-
02
b111 6
#128790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#128800000000
0!
0%
b0 *
0-
02
b0 6
#128810000000
1!
1%
1-
12
#128820000000
0!
0%
b1 *
0-
02
b1 6
#128830000000
1!
1%
1-
12
#128840000000
0!
0%
b10 *
0-
02
b10 6
#128850000000
1!
1%
1-
12
#128860000000
0!
0%
b11 *
0-
02
b11 6
#128870000000
1!
1%
1-
12
15
#128880000000
0!
0%
b100 *
0-
02
b100 6
#128890000000
1!
1%
1-
12
#128900000000
0!
0%
b101 *
0-
02
b101 6
#128910000000
1!
1%
1-
12
#128920000000
0!
0%
b110 *
0-
02
b110 6
#128930000000
1!
1%
1-
12
#128940000000
0!
0%
b111 *
0-
02
b111 6
#128950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#128960000000
0!
0%
b0 *
0-
02
b0 6
#128970000000
1!
1%
1-
12
#128980000000
0!
0%
b1 *
0-
02
b1 6
#128990000000
1!
1%
1-
12
#129000000000
0!
0%
b10 *
0-
02
b10 6
#129010000000
1!
1%
1-
12
#129020000000
0!
0%
b11 *
0-
02
b11 6
#129030000000
1!
1%
1-
12
15
#129040000000
0!
0%
b100 *
0-
02
b100 6
#129050000000
1!
1%
1-
12
#129060000000
0!
0%
b101 *
0-
02
b101 6
#129070000000
1!
1%
1-
12
#129080000000
0!
0%
b110 *
0-
02
b110 6
#129090000000
1!
1%
1-
12
#129100000000
0!
0%
b111 *
0-
02
b111 6
#129110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#129120000000
0!
0%
b0 *
0-
02
b0 6
#129130000000
1!
1%
1-
12
#129140000000
0!
0%
b1 *
0-
02
b1 6
#129150000000
1!
1%
1-
12
#129160000000
0!
0%
b10 *
0-
02
b10 6
#129170000000
1!
1%
1-
12
#129180000000
0!
0%
b11 *
0-
02
b11 6
#129190000000
1!
1%
1-
12
15
#129200000000
0!
0%
b100 *
0-
02
b100 6
#129210000000
1!
1%
1-
12
#129220000000
0!
0%
b101 *
0-
02
b101 6
#129230000000
1!
1%
1-
12
#129240000000
0!
0%
b110 *
0-
02
b110 6
#129250000000
1!
1%
1-
12
#129260000000
0!
0%
b111 *
0-
02
b111 6
#129270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#129280000000
0!
0%
b0 *
0-
02
b0 6
#129290000000
1!
1%
1-
12
#129300000000
0!
0%
b1 *
0-
02
b1 6
#129310000000
1!
1%
1-
12
#129320000000
0!
0%
b10 *
0-
02
b10 6
#129330000000
1!
1%
1-
12
#129340000000
0!
0%
b11 *
0-
02
b11 6
#129350000000
1!
1%
1-
12
15
#129360000000
0!
0%
b100 *
0-
02
b100 6
#129370000000
1!
1%
1-
12
#129380000000
0!
0%
b101 *
0-
02
b101 6
#129390000000
1!
1%
1-
12
#129400000000
0!
0%
b110 *
0-
02
b110 6
#129410000000
1!
1%
1-
12
#129420000000
0!
0%
b111 *
0-
02
b111 6
#129430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#129440000000
0!
0%
b0 *
0-
02
b0 6
#129450000000
1!
1%
1-
12
#129460000000
0!
0%
b1 *
0-
02
b1 6
#129470000000
1!
1%
1-
12
#129480000000
0!
0%
b10 *
0-
02
b10 6
#129490000000
1!
1%
1-
12
#129500000000
0!
0%
b11 *
0-
02
b11 6
#129510000000
1!
1%
1-
12
15
#129520000000
0!
0%
b100 *
0-
02
b100 6
#129530000000
1!
1%
1-
12
#129540000000
0!
0%
b101 *
0-
02
b101 6
#129550000000
1!
1%
1-
12
#129560000000
0!
0%
b110 *
0-
02
b110 6
#129570000000
1!
1%
1-
12
#129580000000
0!
0%
b111 *
0-
02
b111 6
#129590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#129600000000
0!
0%
b0 *
0-
02
b0 6
#129610000000
1!
1%
1-
12
#129620000000
0!
0%
b1 *
0-
02
b1 6
#129630000000
1!
1%
1-
12
#129640000000
0!
0%
b10 *
0-
02
b10 6
#129650000000
1!
1%
1-
12
#129660000000
0!
0%
b11 *
0-
02
b11 6
#129670000000
1!
1%
1-
12
15
#129680000000
0!
0%
b100 *
0-
02
b100 6
#129690000000
1!
1%
1-
12
#129700000000
0!
0%
b101 *
0-
02
b101 6
#129710000000
1!
1%
1-
12
#129720000000
0!
0%
b110 *
0-
02
b110 6
#129730000000
1!
1%
1-
12
#129740000000
0!
0%
b111 *
0-
02
b111 6
#129750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#129760000000
0!
0%
b0 *
0-
02
b0 6
#129770000000
1!
1%
1-
12
#129780000000
0!
0%
b1 *
0-
02
b1 6
#129790000000
1!
1%
1-
12
#129800000000
0!
0%
b10 *
0-
02
b10 6
#129810000000
1!
1%
1-
12
#129820000000
0!
0%
b11 *
0-
02
b11 6
#129830000000
1!
1%
1-
12
15
#129840000000
0!
0%
b100 *
0-
02
b100 6
#129850000000
1!
1%
1-
12
#129860000000
0!
0%
b101 *
0-
02
b101 6
#129870000000
1!
1%
1-
12
#129880000000
0!
0%
b110 *
0-
02
b110 6
#129890000000
1!
1%
1-
12
#129900000000
0!
0%
b111 *
0-
02
b111 6
#129910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#129920000000
0!
0%
b0 *
0-
02
b0 6
#129930000000
1!
1%
1-
12
#129940000000
0!
0%
b1 *
0-
02
b1 6
#129950000000
1!
1%
1-
12
#129960000000
0!
0%
b10 *
0-
02
b10 6
#129970000000
1!
1%
1-
12
#129980000000
0!
0%
b11 *
0-
02
b11 6
#129990000000
1!
1%
1-
12
15
#130000000000
0!
0%
b100 *
0-
02
b100 6
#130010000000
1!
1%
1-
12
#130020000000
0!
0%
b101 *
0-
02
b101 6
#130030000000
1!
1%
1-
12
#130040000000
0!
0%
b110 *
0-
02
b110 6
#130050000000
1!
1%
1-
12
#130060000000
0!
0%
b111 *
0-
02
b111 6
#130070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#130080000000
0!
0%
b0 *
0-
02
b0 6
#130090000000
1!
1%
1-
12
#130100000000
0!
0%
b1 *
0-
02
b1 6
#130110000000
1!
1%
1-
12
#130120000000
0!
0%
b10 *
0-
02
b10 6
#130130000000
1!
1%
1-
12
#130140000000
0!
0%
b11 *
0-
02
b11 6
#130150000000
1!
1%
1-
12
15
#130160000000
0!
0%
b100 *
0-
02
b100 6
#130170000000
1!
1%
1-
12
#130180000000
0!
0%
b101 *
0-
02
b101 6
#130190000000
1!
1%
1-
12
#130200000000
0!
0%
b110 *
0-
02
b110 6
#130210000000
1!
1%
1-
12
#130220000000
0!
0%
b111 *
0-
02
b111 6
#130230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#130240000000
0!
0%
b0 *
0-
02
b0 6
#130250000000
1!
1%
1-
12
#130260000000
0!
0%
b1 *
0-
02
b1 6
#130270000000
1!
1%
1-
12
#130280000000
0!
0%
b10 *
0-
02
b10 6
#130290000000
1!
1%
1-
12
#130300000000
0!
0%
b11 *
0-
02
b11 6
#130310000000
1!
1%
1-
12
15
#130320000000
0!
0%
b100 *
0-
02
b100 6
#130330000000
1!
1%
1-
12
#130340000000
0!
0%
b101 *
0-
02
b101 6
#130350000000
1!
1%
1-
12
#130360000000
0!
0%
b110 *
0-
02
b110 6
#130370000000
1!
1%
1-
12
#130380000000
0!
0%
b111 *
0-
02
b111 6
#130390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#130400000000
0!
0%
b0 *
0-
02
b0 6
#130410000000
1!
1%
1-
12
#130420000000
0!
0%
b1 *
0-
02
b1 6
#130430000000
1!
1%
1-
12
#130440000000
0!
0%
b10 *
0-
02
b10 6
#130450000000
1!
1%
1-
12
#130460000000
0!
0%
b11 *
0-
02
b11 6
#130470000000
1!
1%
1-
12
15
#130480000000
0!
0%
b100 *
0-
02
b100 6
#130490000000
1!
1%
1-
12
#130500000000
0!
0%
b101 *
0-
02
b101 6
#130510000000
1!
1%
1-
12
#130520000000
0!
0%
b110 *
0-
02
b110 6
#130530000000
1!
1%
1-
12
#130540000000
0!
0%
b111 *
0-
02
b111 6
#130550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#130560000000
0!
0%
b0 *
0-
02
b0 6
#130570000000
1!
1%
1-
12
#130580000000
0!
0%
b1 *
0-
02
b1 6
#130590000000
1!
1%
1-
12
#130600000000
0!
0%
b10 *
0-
02
b10 6
#130610000000
1!
1%
1-
12
#130620000000
0!
0%
b11 *
0-
02
b11 6
#130630000000
1!
1%
1-
12
15
#130640000000
0!
0%
b100 *
0-
02
b100 6
#130650000000
1!
1%
1-
12
#130660000000
0!
0%
b101 *
0-
02
b101 6
#130670000000
1!
1%
1-
12
#130680000000
0!
0%
b110 *
0-
02
b110 6
#130690000000
1!
1%
1-
12
#130700000000
0!
0%
b111 *
0-
02
b111 6
#130710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#130720000000
0!
0%
b0 *
0-
02
b0 6
#130730000000
1!
1%
1-
12
#130740000000
0!
0%
b1 *
0-
02
b1 6
#130750000000
1!
1%
1-
12
#130760000000
0!
0%
b10 *
0-
02
b10 6
#130770000000
1!
1%
1-
12
#130780000000
0!
0%
b11 *
0-
02
b11 6
#130790000000
1!
1%
1-
12
15
#130800000000
0!
0%
b100 *
0-
02
b100 6
#130810000000
1!
1%
1-
12
#130820000000
0!
0%
b101 *
0-
02
b101 6
#130830000000
1!
1%
1-
12
#130840000000
0!
0%
b110 *
0-
02
b110 6
#130850000000
1!
1%
1-
12
#130860000000
0!
0%
b111 *
0-
02
b111 6
#130870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#130880000000
0!
0%
b0 *
0-
02
b0 6
#130890000000
1!
1%
1-
12
#130900000000
0!
0%
b1 *
0-
02
b1 6
#130910000000
1!
1%
1-
12
#130920000000
0!
0%
b10 *
0-
02
b10 6
#130930000000
1!
1%
1-
12
#130940000000
0!
0%
b11 *
0-
02
b11 6
#130950000000
1!
1%
1-
12
15
#130960000000
0!
0%
b100 *
0-
02
b100 6
#130970000000
1!
1%
1-
12
#130980000000
0!
0%
b101 *
0-
02
b101 6
#130990000000
1!
1%
1-
12
#131000000000
0!
0%
b110 *
0-
02
b110 6
#131010000000
1!
1%
1-
12
#131020000000
0!
0%
b111 *
0-
02
b111 6
#131030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#131040000000
0!
0%
b0 *
0-
02
b0 6
#131050000000
1!
1%
1-
12
#131060000000
0!
0%
b1 *
0-
02
b1 6
#131070000000
1!
1%
1-
12
#131080000000
0!
0%
b10 *
0-
02
b10 6
#131090000000
1!
1%
1-
12
#131100000000
0!
0%
b11 *
0-
02
b11 6
#131110000000
1!
1%
1-
12
15
#131120000000
0!
0%
b100 *
0-
02
b100 6
#131130000000
1!
1%
1-
12
#131140000000
0!
0%
b101 *
0-
02
b101 6
#131150000000
1!
1%
1-
12
#131160000000
0!
0%
b110 *
0-
02
b110 6
#131170000000
1!
1%
1-
12
#131180000000
0!
0%
b111 *
0-
02
b111 6
#131190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#131200000000
0!
0%
b0 *
0-
02
b0 6
#131210000000
1!
1%
1-
12
#131220000000
0!
0%
b1 *
0-
02
b1 6
#131230000000
1!
1%
1-
12
#131240000000
0!
0%
b10 *
0-
02
b10 6
#131250000000
1!
1%
1-
12
#131260000000
0!
0%
b11 *
0-
02
b11 6
#131270000000
1!
1%
1-
12
15
#131280000000
0!
0%
b100 *
0-
02
b100 6
#131290000000
1!
1%
1-
12
#131300000000
0!
0%
b101 *
0-
02
b101 6
#131310000000
1!
1%
1-
12
#131320000000
0!
0%
b110 *
0-
02
b110 6
#131330000000
1!
1%
1-
12
#131340000000
0!
0%
b111 *
0-
02
b111 6
#131350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#131360000000
0!
0%
b0 *
0-
02
b0 6
#131370000000
1!
1%
1-
12
#131380000000
0!
0%
b1 *
0-
02
b1 6
#131390000000
1!
1%
1-
12
#131400000000
0!
0%
b10 *
0-
02
b10 6
#131410000000
1!
1%
1-
12
#131420000000
0!
0%
b11 *
0-
02
b11 6
#131430000000
1!
1%
1-
12
15
#131440000000
0!
0%
b100 *
0-
02
b100 6
#131450000000
1!
1%
1-
12
#131460000000
0!
0%
b101 *
0-
02
b101 6
#131470000000
1!
1%
1-
12
#131480000000
0!
0%
b110 *
0-
02
b110 6
#131490000000
1!
1%
1-
12
#131500000000
0!
0%
b111 *
0-
02
b111 6
#131510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#131520000000
0!
0%
b0 *
0-
02
b0 6
#131530000000
1!
1%
1-
12
#131540000000
0!
0%
b1 *
0-
02
b1 6
#131550000000
1!
1%
1-
12
#131560000000
0!
0%
b10 *
0-
02
b10 6
#131570000000
1!
1%
1-
12
#131580000000
0!
0%
b11 *
0-
02
b11 6
#131590000000
1!
1%
1-
12
15
#131600000000
0!
0%
b100 *
0-
02
b100 6
#131610000000
1!
1%
1-
12
#131620000000
0!
0%
b101 *
0-
02
b101 6
#131630000000
1!
1%
1-
12
#131640000000
0!
0%
b110 *
0-
02
b110 6
#131650000000
1!
1%
1-
12
#131660000000
0!
0%
b111 *
0-
02
b111 6
#131670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#131680000000
0!
0%
b0 *
0-
02
b0 6
#131690000000
1!
1%
1-
12
#131700000000
0!
0%
b1 *
0-
02
b1 6
#131710000000
1!
1%
1-
12
#131720000000
0!
0%
b10 *
0-
02
b10 6
#131730000000
1!
1%
1-
12
#131740000000
0!
0%
b11 *
0-
02
b11 6
#131750000000
1!
1%
1-
12
15
#131760000000
0!
0%
b100 *
0-
02
b100 6
#131770000000
1!
1%
1-
12
#131780000000
0!
0%
b101 *
0-
02
b101 6
#131790000000
1!
1%
1-
12
#131800000000
0!
0%
b110 *
0-
02
b110 6
#131810000000
1!
1%
1-
12
#131820000000
0!
0%
b111 *
0-
02
b111 6
#131830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#131840000000
0!
0%
b0 *
0-
02
b0 6
#131850000000
1!
1%
1-
12
#131860000000
0!
0%
b1 *
0-
02
b1 6
#131870000000
1!
1%
1-
12
#131880000000
0!
0%
b10 *
0-
02
b10 6
#131890000000
1!
1%
1-
12
#131900000000
0!
0%
b11 *
0-
02
b11 6
#131910000000
1!
1%
1-
12
15
#131920000000
0!
0%
b100 *
0-
02
b100 6
#131930000000
1!
1%
1-
12
#131940000000
0!
0%
b101 *
0-
02
b101 6
#131950000000
1!
1%
1-
12
#131960000000
0!
0%
b110 *
0-
02
b110 6
#131970000000
1!
1%
1-
12
#131980000000
0!
0%
b111 *
0-
02
b111 6
#131990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#132000000000
0!
0%
b0 *
0-
02
b0 6
#132010000000
1!
1%
1-
12
#132020000000
0!
0%
b1 *
0-
02
b1 6
#132030000000
1!
1%
1-
12
#132040000000
0!
0%
b10 *
0-
02
b10 6
#132050000000
1!
1%
1-
12
#132060000000
0!
0%
b11 *
0-
02
b11 6
#132070000000
1!
1%
1-
12
15
#132080000000
0!
0%
b100 *
0-
02
b100 6
#132090000000
1!
1%
1-
12
#132100000000
0!
0%
b101 *
0-
02
b101 6
#132110000000
1!
1%
1-
12
#132120000000
0!
0%
b110 *
0-
02
b110 6
#132130000000
1!
1%
1-
12
#132140000000
0!
0%
b111 *
0-
02
b111 6
#132150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#132160000000
0!
0%
b0 *
0-
02
b0 6
#132170000000
1!
1%
1-
12
#132180000000
0!
0%
b1 *
0-
02
b1 6
#132190000000
1!
1%
1-
12
#132200000000
0!
0%
b10 *
0-
02
b10 6
#132210000000
1!
1%
1-
12
#132220000000
0!
0%
b11 *
0-
02
b11 6
#132230000000
1!
1%
1-
12
15
#132240000000
0!
0%
b100 *
0-
02
b100 6
#132250000000
1!
1%
1-
12
#132260000000
0!
0%
b101 *
0-
02
b101 6
#132270000000
1!
1%
1-
12
#132280000000
0!
0%
b110 *
0-
02
b110 6
#132290000000
1!
1%
1-
12
#132300000000
0!
0%
b111 *
0-
02
b111 6
#132310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#132320000000
0!
0%
b0 *
0-
02
b0 6
#132330000000
1!
1%
1-
12
#132340000000
0!
0%
b1 *
0-
02
b1 6
#132350000000
1!
1%
1-
12
#132360000000
0!
0%
b10 *
0-
02
b10 6
#132370000000
1!
1%
1-
12
#132380000000
0!
0%
b11 *
0-
02
b11 6
#132390000000
1!
1%
1-
12
15
#132400000000
0!
0%
b100 *
0-
02
b100 6
#132410000000
1!
1%
1-
12
#132420000000
0!
0%
b101 *
0-
02
b101 6
#132430000000
1!
1%
1-
12
#132440000000
0!
0%
b110 *
0-
02
b110 6
#132450000000
1!
1%
1-
12
#132460000000
0!
0%
b111 *
0-
02
b111 6
#132470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#132480000000
0!
0%
b0 *
0-
02
b0 6
#132490000000
1!
1%
1-
12
#132500000000
0!
0%
b1 *
0-
02
b1 6
#132510000000
1!
1%
1-
12
#132520000000
0!
0%
b10 *
0-
02
b10 6
#132530000000
1!
1%
1-
12
#132540000000
0!
0%
b11 *
0-
02
b11 6
#132550000000
1!
1%
1-
12
15
#132560000000
0!
0%
b100 *
0-
02
b100 6
#132570000000
1!
1%
1-
12
#132580000000
0!
0%
b101 *
0-
02
b101 6
#132590000000
1!
1%
1-
12
#132600000000
0!
0%
b110 *
0-
02
b110 6
#132610000000
1!
1%
1-
12
#132620000000
0!
0%
b111 *
0-
02
b111 6
#132630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#132640000000
0!
0%
b0 *
0-
02
b0 6
#132650000000
1!
1%
1-
12
#132660000000
0!
0%
b1 *
0-
02
b1 6
#132670000000
1!
1%
1-
12
#132680000000
0!
0%
b10 *
0-
02
b10 6
#132690000000
1!
1%
1-
12
#132700000000
0!
0%
b11 *
0-
02
b11 6
#132710000000
1!
1%
1-
12
15
#132720000000
0!
0%
b100 *
0-
02
b100 6
#132730000000
1!
1%
1-
12
#132740000000
0!
0%
b101 *
0-
02
b101 6
#132750000000
1!
1%
1-
12
#132760000000
0!
0%
b110 *
0-
02
b110 6
#132770000000
1!
1%
1-
12
#132780000000
0!
0%
b111 *
0-
02
b111 6
#132790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#132800000000
0!
0%
b0 *
0-
02
b0 6
#132810000000
1!
1%
1-
12
#132820000000
0!
0%
b1 *
0-
02
b1 6
#132830000000
1!
1%
1-
12
#132840000000
0!
0%
b10 *
0-
02
b10 6
#132850000000
1!
1%
1-
12
#132860000000
0!
0%
b11 *
0-
02
b11 6
#132870000000
1!
1%
1-
12
15
#132880000000
0!
0%
b100 *
0-
02
b100 6
#132890000000
1!
1%
1-
12
#132900000000
0!
0%
b101 *
0-
02
b101 6
#132910000000
1!
1%
1-
12
#132920000000
0!
0%
b110 *
0-
02
b110 6
#132930000000
1!
1%
1-
12
#132940000000
0!
0%
b111 *
0-
02
b111 6
#132950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#132960000000
0!
0%
b0 *
0-
02
b0 6
#132970000000
1!
1%
1-
12
#132980000000
0!
0%
b1 *
0-
02
b1 6
#132990000000
1!
1%
1-
12
#133000000000
0!
0%
b10 *
0-
02
b10 6
#133010000000
1!
1%
1-
12
#133020000000
0!
0%
b11 *
0-
02
b11 6
#133030000000
1!
1%
1-
12
15
#133040000000
0!
0%
b100 *
0-
02
b100 6
#133050000000
1!
1%
1-
12
#133060000000
0!
0%
b101 *
0-
02
b101 6
#133070000000
1!
1%
1-
12
#133080000000
0!
0%
b110 *
0-
02
b110 6
#133090000000
1!
1%
1-
12
#133100000000
0!
0%
b111 *
0-
02
b111 6
#133110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#133120000000
0!
0%
b0 *
0-
02
b0 6
#133130000000
1!
1%
1-
12
#133140000000
0!
0%
b1 *
0-
02
b1 6
#133150000000
1!
1%
1-
12
#133160000000
0!
0%
b10 *
0-
02
b10 6
#133170000000
1!
1%
1-
12
#133180000000
0!
0%
b11 *
0-
02
b11 6
#133190000000
1!
1%
1-
12
15
#133200000000
0!
0%
b100 *
0-
02
b100 6
#133210000000
1!
1%
1-
12
#133220000000
0!
0%
b101 *
0-
02
b101 6
#133230000000
1!
1%
1-
12
#133240000000
0!
0%
b110 *
0-
02
b110 6
#133250000000
1!
1%
1-
12
#133260000000
0!
0%
b111 *
0-
02
b111 6
#133270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#133280000000
0!
0%
b0 *
0-
02
b0 6
#133290000000
1!
1%
1-
12
#133300000000
0!
0%
b1 *
0-
02
b1 6
#133310000000
1!
1%
1-
12
#133320000000
0!
0%
b10 *
0-
02
b10 6
#133330000000
1!
1%
1-
12
#133340000000
0!
0%
b11 *
0-
02
b11 6
#133350000000
1!
1%
1-
12
15
#133360000000
0!
0%
b100 *
0-
02
b100 6
#133370000000
1!
1%
1-
12
#133380000000
0!
0%
b101 *
0-
02
b101 6
#133390000000
1!
1%
1-
12
#133400000000
0!
0%
b110 *
0-
02
b110 6
#133410000000
1!
1%
1-
12
#133420000000
0!
0%
b111 *
0-
02
b111 6
#133430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#133440000000
0!
0%
b0 *
0-
02
b0 6
#133450000000
1!
1%
1-
12
#133460000000
0!
0%
b1 *
0-
02
b1 6
#133470000000
1!
1%
1-
12
#133480000000
0!
0%
b10 *
0-
02
b10 6
#133490000000
1!
1%
1-
12
#133500000000
0!
0%
b11 *
0-
02
b11 6
#133510000000
1!
1%
1-
12
15
#133520000000
0!
0%
b100 *
0-
02
b100 6
#133530000000
1!
1%
1-
12
#133540000000
0!
0%
b101 *
0-
02
b101 6
#133550000000
1!
1%
1-
12
#133560000000
0!
0%
b110 *
0-
02
b110 6
#133570000000
1!
1%
1-
12
#133580000000
0!
0%
b111 *
0-
02
b111 6
#133590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#133600000000
0!
0%
b0 *
0-
02
b0 6
#133610000000
1!
1%
1-
12
#133620000000
0!
0%
b1 *
0-
02
b1 6
#133630000000
1!
1%
1-
12
#133640000000
0!
0%
b10 *
0-
02
b10 6
#133650000000
1!
1%
1-
12
#133660000000
0!
0%
b11 *
0-
02
b11 6
#133670000000
1!
1%
1-
12
15
#133680000000
0!
0%
b100 *
0-
02
b100 6
#133690000000
1!
1%
1-
12
#133700000000
0!
0%
b101 *
0-
02
b101 6
#133710000000
1!
1%
1-
12
#133720000000
0!
0%
b110 *
0-
02
b110 6
#133730000000
1!
1%
1-
12
#133740000000
0!
0%
b111 *
0-
02
b111 6
#133750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#133760000000
0!
0%
b0 *
0-
02
b0 6
#133770000000
1!
1%
1-
12
#133780000000
0!
0%
b1 *
0-
02
b1 6
#133790000000
1!
1%
1-
12
#133800000000
0!
0%
b10 *
0-
02
b10 6
#133810000000
1!
1%
1-
12
#133820000000
0!
0%
b11 *
0-
02
b11 6
#133830000000
1!
1%
1-
12
15
#133840000000
0!
0%
b100 *
0-
02
b100 6
#133850000000
1!
1%
1-
12
#133860000000
0!
0%
b101 *
0-
02
b101 6
#133870000000
1!
1%
1-
12
#133880000000
0!
0%
b110 *
0-
02
b110 6
#133890000000
1!
1%
1-
12
#133900000000
0!
0%
b111 *
0-
02
b111 6
#133910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#133920000000
0!
0%
b0 *
0-
02
b0 6
#133930000000
1!
1%
1-
12
#133940000000
0!
0%
b1 *
0-
02
b1 6
#133950000000
1!
1%
1-
12
#133960000000
0!
0%
b10 *
0-
02
b10 6
#133970000000
1!
1%
1-
12
#133980000000
0!
0%
b11 *
0-
02
b11 6
#133990000000
1!
1%
1-
12
15
#134000000000
0!
0%
b100 *
0-
02
b100 6
#134010000000
1!
1%
1-
12
#134020000000
0!
0%
b101 *
0-
02
b101 6
#134030000000
1!
1%
1-
12
#134040000000
0!
0%
b110 *
0-
02
b110 6
#134050000000
1!
1%
1-
12
#134060000000
0!
0%
b111 *
0-
02
b111 6
#134070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#134080000000
0!
0%
b0 *
0-
02
b0 6
#134090000000
1!
1%
1-
12
#134100000000
0!
0%
b1 *
0-
02
b1 6
#134110000000
1!
1%
1-
12
#134120000000
0!
0%
b10 *
0-
02
b10 6
#134130000000
1!
1%
1-
12
#134140000000
0!
0%
b11 *
0-
02
b11 6
#134150000000
1!
1%
1-
12
15
#134160000000
0!
0%
b100 *
0-
02
b100 6
#134170000000
1!
1%
1-
12
#134180000000
0!
0%
b101 *
0-
02
b101 6
#134190000000
1!
1%
1-
12
#134200000000
0!
0%
b110 *
0-
02
b110 6
#134210000000
1!
1%
1-
12
#134220000000
0!
0%
b111 *
0-
02
b111 6
#134230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#134240000000
0!
0%
b0 *
0-
02
b0 6
#134250000000
1!
1%
1-
12
#134260000000
0!
0%
b1 *
0-
02
b1 6
#134270000000
1!
1%
1-
12
#134280000000
0!
0%
b10 *
0-
02
b10 6
#134290000000
1!
1%
1-
12
#134300000000
0!
0%
b11 *
0-
02
b11 6
#134310000000
1!
1%
1-
12
15
#134320000000
0!
0%
b100 *
0-
02
b100 6
#134330000000
1!
1%
1-
12
#134340000000
0!
0%
b101 *
0-
02
b101 6
#134350000000
1!
1%
1-
12
#134360000000
0!
0%
b110 *
0-
02
b110 6
#134370000000
1!
1%
1-
12
#134380000000
0!
0%
b111 *
0-
02
b111 6
#134390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#134400000000
0!
0%
b0 *
0-
02
b0 6
#134410000000
1!
1%
1-
12
#134420000000
0!
0%
b1 *
0-
02
b1 6
#134430000000
1!
1%
1-
12
#134440000000
0!
0%
b10 *
0-
02
b10 6
#134450000000
1!
1%
1-
12
#134460000000
0!
0%
b11 *
0-
02
b11 6
#134470000000
1!
1%
1-
12
15
#134480000000
0!
0%
b100 *
0-
02
b100 6
#134490000000
1!
1%
1-
12
#134500000000
0!
0%
b101 *
0-
02
b101 6
#134510000000
1!
1%
1-
12
#134520000000
0!
0%
b110 *
0-
02
b110 6
#134530000000
1!
1%
1-
12
#134540000000
0!
0%
b111 *
0-
02
b111 6
#134550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#134560000000
0!
0%
b0 *
0-
02
b0 6
#134570000000
1!
1%
1-
12
#134580000000
0!
0%
b1 *
0-
02
b1 6
#134590000000
1!
1%
1-
12
#134600000000
0!
0%
b10 *
0-
02
b10 6
#134610000000
1!
1%
1-
12
#134620000000
0!
0%
b11 *
0-
02
b11 6
#134630000000
1!
1%
1-
12
15
#134640000000
0!
0%
b100 *
0-
02
b100 6
#134650000000
1!
1%
1-
12
#134660000000
0!
0%
b101 *
0-
02
b101 6
#134670000000
1!
1%
1-
12
#134680000000
0!
0%
b110 *
0-
02
b110 6
#134690000000
1!
1%
1-
12
#134700000000
0!
0%
b111 *
0-
02
b111 6
#134710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#134720000000
0!
0%
b0 *
0-
02
b0 6
#134730000000
1!
1%
1-
12
#134740000000
0!
0%
b1 *
0-
02
b1 6
#134750000000
1!
1%
1-
12
#134760000000
0!
0%
b10 *
0-
02
b10 6
#134770000000
1!
1%
1-
12
#134780000000
0!
0%
b11 *
0-
02
b11 6
#134790000000
1!
1%
1-
12
15
#134800000000
0!
0%
b100 *
0-
02
b100 6
#134810000000
1!
1%
1-
12
#134820000000
0!
0%
b101 *
0-
02
b101 6
#134830000000
1!
1%
1-
12
#134840000000
0!
0%
b110 *
0-
02
b110 6
#134850000000
1!
1%
1-
12
#134860000000
0!
0%
b111 *
0-
02
b111 6
#134870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#134880000000
0!
0%
b0 *
0-
02
b0 6
#134890000000
1!
1%
1-
12
#134900000000
0!
0%
b1 *
0-
02
b1 6
#134910000000
1!
1%
1-
12
#134920000000
0!
0%
b10 *
0-
02
b10 6
#134930000000
1!
1%
1-
12
#134940000000
0!
0%
b11 *
0-
02
b11 6
#134950000000
1!
1%
1-
12
15
#134960000000
0!
0%
b100 *
0-
02
b100 6
#134970000000
1!
1%
1-
12
#134980000000
0!
0%
b101 *
0-
02
b101 6
#134990000000
1!
1%
1-
12
#135000000000
0!
0%
b110 *
0-
02
b110 6
#135010000000
1!
1%
1-
12
#135020000000
0!
0%
b111 *
0-
02
b111 6
#135030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#135040000000
0!
0%
b0 *
0-
02
b0 6
#135050000000
1!
1%
1-
12
#135060000000
0!
0%
b1 *
0-
02
b1 6
#135070000000
1!
1%
1-
12
#135080000000
0!
0%
b10 *
0-
02
b10 6
#135090000000
1!
1%
1-
12
#135100000000
0!
0%
b11 *
0-
02
b11 6
#135110000000
1!
1%
1-
12
15
#135120000000
0!
0%
b100 *
0-
02
b100 6
#135130000000
1!
1%
1-
12
#135140000000
0!
0%
b101 *
0-
02
b101 6
#135150000000
1!
1%
1-
12
#135160000000
0!
0%
b110 *
0-
02
b110 6
#135170000000
1!
1%
1-
12
#135180000000
0!
0%
b111 *
0-
02
b111 6
#135190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#135200000000
0!
0%
b0 *
0-
02
b0 6
#135210000000
1!
1%
1-
12
#135220000000
0!
0%
b1 *
0-
02
b1 6
#135230000000
1!
1%
1-
12
#135240000000
0!
0%
b10 *
0-
02
b10 6
#135250000000
1!
1%
1-
12
#135260000000
0!
0%
b11 *
0-
02
b11 6
#135270000000
1!
1%
1-
12
15
#135280000000
0!
0%
b100 *
0-
02
b100 6
#135290000000
1!
1%
1-
12
#135300000000
0!
0%
b101 *
0-
02
b101 6
#135310000000
1!
1%
1-
12
#135320000000
0!
0%
b110 *
0-
02
b110 6
#135330000000
1!
1%
1-
12
#135340000000
0!
0%
b111 *
0-
02
b111 6
#135350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#135360000000
0!
0%
b0 *
0-
02
b0 6
#135370000000
1!
1%
1-
12
#135380000000
0!
0%
b1 *
0-
02
b1 6
#135390000000
1!
1%
1-
12
#135400000000
0!
0%
b10 *
0-
02
b10 6
#135410000000
1!
1%
1-
12
#135420000000
0!
0%
b11 *
0-
02
b11 6
#135430000000
1!
1%
1-
12
15
#135440000000
0!
0%
b100 *
0-
02
b100 6
#135450000000
1!
1%
1-
12
#135460000000
0!
0%
b101 *
0-
02
b101 6
#135470000000
1!
1%
1-
12
#135480000000
0!
0%
b110 *
0-
02
b110 6
#135490000000
1!
1%
1-
12
#135500000000
0!
0%
b111 *
0-
02
b111 6
#135510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#135520000000
0!
0%
b0 *
0-
02
b0 6
#135530000000
1!
1%
1-
12
#135540000000
0!
0%
b1 *
0-
02
b1 6
#135550000000
1!
1%
1-
12
#135560000000
0!
0%
b10 *
0-
02
b10 6
#135570000000
1!
1%
1-
12
#135580000000
0!
0%
b11 *
0-
02
b11 6
#135590000000
1!
1%
1-
12
15
#135600000000
0!
0%
b100 *
0-
02
b100 6
#135610000000
1!
1%
1-
12
#135620000000
0!
0%
b101 *
0-
02
b101 6
#135630000000
1!
1%
1-
12
#135640000000
0!
0%
b110 *
0-
02
b110 6
#135650000000
1!
1%
1-
12
#135660000000
0!
0%
b111 *
0-
02
b111 6
#135670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#135680000000
0!
0%
b0 *
0-
02
b0 6
#135690000000
1!
1%
1-
12
#135700000000
0!
0%
b1 *
0-
02
b1 6
#135710000000
1!
1%
1-
12
#135720000000
0!
0%
b10 *
0-
02
b10 6
#135730000000
1!
1%
1-
12
#135740000000
0!
0%
b11 *
0-
02
b11 6
#135750000000
1!
1%
1-
12
15
#135760000000
0!
0%
b100 *
0-
02
b100 6
#135770000000
1!
1%
1-
12
#135780000000
0!
0%
b101 *
0-
02
b101 6
#135790000000
1!
1%
1-
12
#135800000000
0!
0%
b110 *
0-
02
b110 6
#135810000000
1!
1%
1-
12
#135820000000
0!
0%
b111 *
0-
02
b111 6
#135830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#135840000000
0!
0%
b0 *
0-
02
b0 6
#135850000000
1!
1%
1-
12
#135860000000
0!
0%
b1 *
0-
02
b1 6
#135870000000
1!
1%
1-
12
#135880000000
0!
0%
b10 *
0-
02
b10 6
#135890000000
1!
1%
1-
12
#135900000000
0!
0%
b11 *
0-
02
b11 6
#135910000000
1!
1%
1-
12
15
#135920000000
0!
0%
b100 *
0-
02
b100 6
#135930000000
1!
1%
1-
12
#135940000000
0!
0%
b101 *
0-
02
b101 6
#135950000000
1!
1%
1-
12
#135960000000
0!
0%
b110 *
0-
02
b110 6
#135970000000
1!
1%
1-
12
#135980000000
0!
0%
b111 *
0-
02
b111 6
#135990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#136000000000
0!
0%
b0 *
0-
02
b0 6
#136010000000
1!
1%
1-
12
#136020000000
0!
0%
b1 *
0-
02
b1 6
#136030000000
1!
1%
1-
12
#136040000000
0!
0%
b10 *
0-
02
b10 6
#136050000000
1!
1%
1-
12
#136060000000
0!
0%
b11 *
0-
02
b11 6
#136070000000
1!
1%
1-
12
15
#136080000000
0!
0%
b100 *
0-
02
b100 6
#136090000000
1!
1%
1-
12
#136100000000
0!
0%
b101 *
0-
02
b101 6
#136110000000
1!
1%
1-
12
#136120000000
0!
0%
b110 *
0-
02
b110 6
#136130000000
1!
1%
1-
12
#136140000000
0!
0%
b111 *
0-
02
b111 6
#136150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#136160000000
0!
0%
b0 *
0-
02
b0 6
#136170000000
1!
1%
1-
12
#136180000000
0!
0%
b1 *
0-
02
b1 6
#136190000000
1!
1%
1-
12
#136200000000
0!
0%
b10 *
0-
02
b10 6
#136210000000
1!
1%
1-
12
#136220000000
0!
0%
b11 *
0-
02
b11 6
#136230000000
1!
1%
1-
12
15
#136240000000
0!
0%
b100 *
0-
02
b100 6
#136250000000
1!
1%
1-
12
#136260000000
0!
0%
b101 *
0-
02
b101 6
#136270000000
1!
1%
1-
12
#136280000000
0!
0%
b110 *
0-
02
b110 6
#136290000000
1!
1%
1-
12
#136300000000
0!
0%
b111 *
0-
02
b111 6
#136310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#136320000000
0!
0%
b0 *
0-
02
b0 6
#136330000000
1!
1%
1-
12
#136340000000
0!
0%
b1 *
0-
02
b1 6
#136350000000
1!
1%
1-
12
#136360000000
0!
0%
b10 *
0-
02
b10 6
#136370000000
1!
1%
1-
12
#136380000000
0!
0%
b11 *
0-
02
b11 6
#136390000000
1!
1%
1-
12
15
#136400000000
0!
0%
b100 *
0-
02
b100 6
#136410000000
1!
1%
1-
12
#136420000000
0!
0%
b101 *
0-
02
b101 6
#136430000000
1!
1%
1-
12
#136440000000
0!
0%
b110 *
0-
02
b110 6
#136450000000
1!
1%
1-
12
#136460000000
0!
0%
b111 *
0-
02
b111 6
#136470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#136480000000
0!
0%
b0 *
0-
02
b0 6
#136490000000
1!
1%
1-
12
#136500000000
0!
0%
b1 *
0-
02
b1 6
#136510000000
1!
1%
1-
12
#136520000000
0!
0%
b10 *
0-
02
b10 6
#136530000000
1!
1%
1-
12
#136540000000
0!
0%
b11 *
0-
02
b11 6
#136550000000
1!
1%
1-
12
15
#136560000000
0!
0%
b100 *
0-
02
b100 6
#136570000000
1!
1%
1-
12
#136580000000
0!
0%
b101 *
0-
02
b101 6
#136590000000
1!
1%
1-
12
#136600000000
0!
0%
b110 *
0-
02
b110 6
#136610000000
1!
1%
1-
12
#136620000000
0!
0%
b111 *
0-
02
b111 6
#136630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#136640000000
0!
0%
b0 *
0-
02
b0 6
#136650000000
1!
1%
1-
12
#136660000000
0!
0%
b1 *
0-
02
b1 6
#136670000000
1!
1%
1-
12
#136680000000
0!
0%
b10 *
0-
02
b10 6
#136690000000
1!
1%
1-
12
#136700000000
0!
0%
b11 *
0-
02
b11 6
#136710000000
1!
1%
1-
12
15
#136720000000
0!
0%
b100 *
0-
02
b100 6
#136730000000
1!
1%
1-
12
#136740000000
0!
0%
b101 *
0-
02
b101 6
#136750000000
1!
1%
1-
12
#136760000000
0!
0%
b110 *
0-
02
b110 6
#136770000000
1!
1%
1-
12
#136780000000
0!
0%
b111 *
0-
02
b111 6
#136790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#136800000000
0!
0%
b0 *
0-
02
b0 6
#136810000000
1!
1%
1-
12
#136820000000
0!
0%
b1 *
0-
02
b1 6
#136830000000
1!
1%
1-
12
#136840000000
0!
0%
b10 *
0-
02
b10 6
#136850000000
1!
1%
1-
12
#136860000000
0!
0%
b11 *
0-
02
b11 6
#136870000000
1!
1%
1-
12
15
#136880000000
0!
0%
b100 *
0-
02
b100 6
#136890000000
1!
1%
1-
12
#136900000000
0!
0%
b101 *
0-
02
b101 6
#136910000000
1!
1%
1-
12
#136920000000
0!
0%
b110 *
0-
02
b110 6
#136930000000
1!
1%
1-
12
#136940000000
0!
0%
b111 *
0-
02
b111 6
#136950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#136960000000
0!
0%
b0 *
0-
02
b0 6
#136970000000
1!
1%
1-
12
#136980000000
0!
0%
b1 *
0-
02
b1 6
#136990000000
1!
1%
1-
12
#137000000000
0!
0%
b10 *
0-
02
b10 6
#137010000000
1!
1%
1-
12
#137020000000
0!
0%
b11 *
0-
02
b11 6
#137030000000
1!
1%
1-
12
15
#137040000000
0!
0%
b100 *
0-
02
b100 6
#137050000000
1!
1%
1-
12
#137060000000
0!
0%
b101 *
0-
02
b101 6
#137070000000
1!
1%
1-
12
#137080000000
0!
0%
b110 *
0-
02
b110 6
#137090000000
1!
1%
1-
12
#137100000000
0!
0%
b111 *
0-
02
b111 6
#137110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#137120000000
0!
0%
b0 *
0-
02
b0 6
#137130000000
1!
1%
1-
12
#137140000000
0!
0%
b1 *
0-
02
b1 6
#137150000000
1!
1%
1-
12
#137160000000
0!
0%
b10 *
0-
02
b10 6
#137170000000
1!
1%
1-
12
#137180000000
0!
0%
b11 *
0-
02
b11 6
#137190000000
1!
1%
1-
12
15
#137200000000
0!
0%
b100 *
0-
02
b100 6
#137210000000
1!
1%
1-
12
#137220000000
0!
0%
b101 *
0-
02
b101 6
#137230000000
1!
1%
1-
12
#137240000000
0!
0%
b110 *
0-
02
b110 6
#137250000000
1!
1%
1-
12
#137260000000
0!
0%
b111 *
0-
02
b111 6
#137270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#137280000000
0!
0%
b0 *
0-
02
b0 6
#137290000000
1!
1%
1-
12
#137300000000
0!
0%
b1 *
0-
02
b1 6
#137310000000
1!
1%
1-
12
#137320000000
0!
0%
b10 *
0-
02
b10 6
#137330000000
1!
1%
1-
12
#137340000000
0!
0%
b11 *
0-
02
b11 6
#137350000000
1!
1%
1-
12
15
#137360000000
0!
0%
b100 *
0-
02
b100 6
#137370000000
1!
1%
1-
12
#137380000000
0!
0%
b101 *
0-
02
b101 6
#137390000000
1!
1%
1-
12
#137400000000
0!
0%
b110 *
0-
02
b110 6
#137410000000
1!
1%
1-
12
#137420000000
0!
0%
b111 *
0-
02
b111 6
#137430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#137440000000
0!
0%
b0 *
0-
02
b0 6
#137450000000
1!
1%
1-
12
#137460000000
0!
0%
b1 *
0-
02
b1 6
#137470000000
1!
1%
1-
12
#137480000000
0!
0%
b10 *
0-
02
b10 6
#137490000000
1!
1%
1-
12
#137500000000
0!
0%
b11 *
0-
02
b11 6
#137510000000
1!
1%
1-
12
15
#137520000000
0!
0%
b100 *
0-
02
b100 6
#137530000000
1!
1%
1-
12
#137540000000
0!
0%
b101 *
0-
02
b101 6
#137550000000
1!
1%
1-
12
#137560000000
0!
0%
b110 *
0-
02
b110 6
#137570000000
1!
1%
1-
12
#137580000000
0!
0%
b111 *
0-
02
b111 6
#137590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#137600000000
0!
0%
b0 *
0-
02
b0 6
#137610000000
1!
1%
1-
12
#137620000000
0!
0%
b1 *
0-
02
b1 6
#137630000000
1!
1%
1-
12
#137640000000
0!
0%
b10 *
0-
02
b10 6
#137650000000
1!
1%
1-
12
#137660000000
0!
0%
b11 *
0-
02
b11 6
#137670000000
1!
1%
1-
12
15
#137680000000
0!
0%
b100 *
0-
02
b100 6
#137690000000
1!
1%
1-
12
#137700000000
0!
0%
b101 *
0-
02
b101 6
#137710000000
1!
1%
1-
12
#137720000000
0!
0%
b110 *
0-
02
b110 6
#137730000000
1!
1%
1-
12
#137740000000
0!
0%
b111 *
0-
02
b111 6
#137750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#137760000000
0!
0%
b0 *
0-
02
b0 6
#137770000000
1!
1%
1-
12
#137780000000
0!
0%
b1 *
0-
02
b1 6
#137790000000
1!
1%
1-
12
#137800000000
0!
0%
b10 *
0-
02
b10 6
#137810000000
1!
1%
1-
12
#137820000000
0!
0%
b11 *
0-
02
b11 6
#137830000000
1!
1%
1-
12
15
#137840000000
0!
0%
b100 *
0-
02
b100 6
#137850000000
1!
1%
1-
12
#137860000000
0!
0%
b101 *
0-
02
b101 6
#137870000000
1!
1%
1-
12
#137880000000
0!
0%
b110 *
0-
02
b110 6
#137890000000
1!
1%
1-
12
#137900000000
0!
0%
b111 *
0-
02
b111 6
#137910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#137920000000
0!
0%
b0 *
0-
02
b0 6
#137930000000
1!
1%
1-
12
#137940000000
0!
0%
b1 *
0-
02
b1 6
#137950000000
1!
1%
1-
12
#137960000000
0!
0%
b10 *
0-
02
b10 6
#137970000000
1!
1%
1-
12
#137980000000
0!
0%
b11 *
0-
02
b11 6
#137990000000
1!
1%
1-
12
15
#138000000000
0!
0%
b100 *
0-
02
b100 6
#138010000000
1!
1%
1-
12
#138020000000
0!
0%
b101 *
0-
02
b101 6
#138030000000
1!
1%
1-
12
#138040000000
0!
0%
b110 *
0-
02
b110 6
#138050000000
1!
1%
1-
12
#138060000000
0!
0%
b111 *
0-
02
b111 6
#138070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#138080000000
0!
0%
b0 *
0-
02
b0 6
#138090000000
1!
1%
1-
12
#138100000000
0!
0%
b1 *
0-
02
b1 6
#138110000000
1!
1%
1-
12
#138120000000
0!
0%
b10 *
0-
02
b10 6
#138130000000
1!
1%
1-
12
#138140000000
0!
0%
b11 *
0-
02
b11 6
#138150000000
1!
1%
1-
12
15
#138160000000
0!
0%
b100 *
0-
02
b100 6
#138170000000
1!
1%
1-
12
#138180000000
0!
0%
b101 *
0-
02
b101 6
#138190000000
1!
1%
1-
12
#138200000000
0!
0%
b110 *
0-
02
b110 6
#138210000000
1!
1%
1-
12
#138220000000
0!
0%
b111 *
0-
02
b111 6
#138230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#138240000000
0!
0%
b0 *
0-
02
b0 6
#138250000000
1!
1%
1-
12
#138260000000
0!
0%
b1 *
0-
02
b1 6
#138270000000
1!
1%
1-
12
#138280000000
0!
0%
b10 *
0-
02
b10 6
#138290000000
1!
1%
1-
12
#138300000000
0!
0%
b11 *
0-
02
b11 6
#138310000000
1!
1%
1-
12
15
#138320000000
0!
0%
b100 *
0-
02
b100 6
#138330000000
1!
1%
1-
12
#138340000000
0!
0%
b101 *
0-
02
b101 6
#138350000000
1!
1%
1-
12
#138360000000
0!
0%
b110 *
0-
02
b110 6
#138370000000
1!
1%
1-
12
#138380000000
0!
0%
b111 *
0-
02
b111 6
#138390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#138400000000
0!
0%
b0 *
0-
02
b0 6
#138410000000
1!
1%
1-
12
#138420000000
0!
0%
b1 *
0-
02
b1 6
#138430000000
1!
1%
1-
12
#138440000000
0!
0%
b10 *
0-
02
b10 6
#138450000000
1!
1%
1-
12
#138460000000
0!
0%
b11 *
0-
02
b11 6
#138470000000
1!
1%
1-
12
15
#138480000000
0!
0%
b100 *
0-
02
b100 6
#138490000000
1!
1%
1-
12
#138500000000
0!
0%
b101 *
0-
02
b101 6
#138510000000
1!
1%
1-
12
#138520000000
0!
0%
b110 *
0-
02
b110 6
#138530000000
1!
1%
1-
12
#138540000000
0!
0%
b111 *
0-
02
b111 6
#138550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#138560000000
0!
0%
b0 *
0-
02
b0 6
#138570000000
1!
1%
1-
12
#138580000000
0!
0%
b1 *
0-
02
b1 6
#138590000000
1!
1%
1-
12
#138600000000
0!
0%
b10 *
0-
02
b10 6
#138610000000
1!
1%
1-
12
#138620000000
0!
0%
b11 *
0-
02
b11 6
#138630000000
1!
1%
1-
12
15
#138640000000
0!
0%
b100 *
0-
02
b100 6
#138650000000
1!
1%
1-
12
#138660000000
0!
0%
b101 *
0-
02
b101 6
#138670000000
1!
1%
1-
12
#138680000000
0!
0%
b110 *
0-
02
b110 6
#138690000000
1!
1%
1-
12
#138700000000
0!
0%
b111 *
0-
02
b111 6
#138710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#138720000000
0!
0%
b0 *
0-
02
b0 6
#138730000000
1!
1%
1-
12
#138740000000
0!
0%
b1 *
0-
02
b1 6
#138750000000
1!
1%
1-
12
#138760000000
0!
0%
b10 *
0-
02
b10 6
#138770000000
1!
1%
1-
12
#138780000000
0!
0%
b11 *
0-
02
b11 6
#138790000000
1!
1%
1-
12
15
#138800000000
0!
0%
b100 *
0-
02
b100 6
#138810000000
1!
1%
1-
12
#138820000000
0!
0%
b101 *
0-
02
b101 6
#138830000000
1!
1%
1-
12
#138840000000
0!
0%
b110 *
0-
02
b110 6
#138850000000
1!
1%
1-
12
#138860000000
0!
0%
b111 *
0-
02
b111 6
#138870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#138880000000
0!
0%
b0 *
0-
02
b0 6
#138890000000
1!
1%
1-
12
#138900000000
0!
0%
b1 *
0-
02
b1 6
#138910000000
1!
1%
1-
12
#138920000000
0!
0%
b10 *
0-
02
b10 6
#138930000000
1!
1%
1-
12
#138940000000
0!
0%
b11 *
0-
02
b11 6
#138950000000
1!
1%
1-
12
15
#138960000000
0!
0%
b100 *
0-
02
b100 6
#138970000000
1!
1%
1-
12
#138980000000
0!
0%
b101 *
0-
02
b101 6
#138990000000
1!
1%
1-
12
#139000000000
0!
0%
b110 *
0-
02
b110 6
#139010000000
1!
1%
1-
12
#139020000000
0!
0%
b111 *
0-
02
b111 6
#139030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#139040000000
0!
0%
b0 *
0-
02
b0 6
#139050000000
1!
1%
1-
12
#139060000000
0!
0%
b1 *
0-
02
b1 6
#139070000000
1!
1%
1-
12
#139080000000
0!
0%
b10 *
0-
02
b10 6
#139090000000
1!
1%
1-
12
#139100000000
0!
0%
b11 *
0-
02
b11 6
#139110000000
1!
1%
1-
12
15
#139120000000
0!
0%
b100 *
0-
02
b100 6
#139130000000
1!
1%
1-
12
#139140000000
0!
0%
b101 *
0-
02
b101 6
#139150000000
1!
1%
1-
12
#139160000000
0!
0%
b110 *
0-
02
b110 6
#139170000000
1!
1%
1-
12
#139180000000
0!
0%
b111 *
0-
02
b111 6
#139190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#139200000000
0!
0%
b0 *
0-
02
b0 6
#139210000000
1!
1%
1-
12
#139220000000
0!
0%
b1 *
0-
02
b1 6
#139230000000
1!
1%
1-
12
#139240000000
0!
0%
b10 *
0-
02
b10 6
#139250000000
1!
1%
1-
12
#139260000000
0!
0%
b11 *
0-
02
b11 6
#139270000000
1!
1%
1-
12
15
#139280000000
0!
0%
b100 *
0-
02
b100 6
#139290000000
1!
1%
1-
12
#139300000000
0!
0%
b101 *
0-
02
b101 6
#139310000000
1!
1%
1-
12
#139320000000
0!
0%
b110 *
0-
02
b110 6
#139330000000
1!
1%
1-
12
#139340000000
0!
0%
b111 *
0-
02
b111 6
#139350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#139360000000
0!
0%
b0 *
0-
02
b0 6
#139370000000
1!
1%
1-
12
#139380000000
0!
0%
b1 *
0-
02
b1 6
#139390000000
1!
1%
1-
12
#139400000000
0!
0%
b10 *
0-
02
b10 6
#139410000000
1!
1%
1-
12
#139420000000
0!
0%
b11 *
0-
02
b11 6
#139430000000
1!
1%
1-
12
15
#139440000000
0!
0%
b100 *
0-
02
b100 6
#139450000000
1!
1%
1-
12
#139460000000
0!
0%
b101 *
0-
02
b101 6
#139470000000
1!
1%
1-
12
#139480000000
0!
0%
b110 *
0-
02
b110 6
#139490000000
1!
1%
1-
12
#139500000000
0!
0%
b111 *
0-
02
b111 6
#139510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#139520000000
0!
0%
b0 *
0-
02
b0 6
#139530000000
1!
1%
1-
12
#139540000000
0!
0%
b1 *
0-
02
b1 6
#139550000000
1!
1%
1-
12
#139560000000
0!
0%
b10 *
0-
02
b10 6
#139570000000
1!
1%
1-
12
#139580000000
0!
0%
b11 *
0-
02
b11 6
#139590000000
1!
1%
1-
12
15
#139600000000
0!
0%
b100 *
0-
02
b100 6
#139610000000
1!
1%
1-
12
#139620000000
0!
0%
b101 *
0-
02
b101 6
#139630000000
1!
1%
1-
12
#139640000000
0!
0%
b110 *
0-
02
b110 6
#139650000000
1!
1%
1-
12
#139660000000
0!
0%
b111 *
0-
02
b111 6
#139670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#139680000000
0!
0%
b0 *
0-
02
b0 6
#139690000000
1!
1%
1-
12
#139700000000
0!
0%
b1 *
0-
02
b1 6
#139710000000
1!
1%
1-
12
#139720000000
0!
0%
b10 *
0-
02
b10 6
#139730000000
1!
1%
1-
12
#139740000000
0!
0%
b11 *
0-
02
b11 6
#139750000000
1!
1%
1-
12
15
#139760000000
0!
0%
b100 *
0-
02
b100 6
#139770000000
1!
1%
1-
12
#139780000000
0!
0%
b101 *
0-
02
b101 6
#139790000000
1!
1%
1-
12
#139800000000
0!
0%
b110 *
0-
02
b110 6
#139810000000
1!
1%
1-
12
#139820000000
0!
0%
b111 *
0-
02
b111 6
#139830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#139840000000
0!
0%
b0 *
0-
02
b0 6
#139850000000
1!
1%
1-
12
#139860000000
0!
0%
b1 *
0-
02
b1 6
#139870000000
1!
1%
1-
12
#139880000000
0!
0%
b10 *
0-
02
b10 6
#139890000000
1!
1%
1-
12
#139900000000
0!
0%
b11 *
0-
02
b11 6
#139910000000
1!
1%
1-
12
15
#139920000000
0!
0%
b100 *
0-
02
b100 6
#139930000000
1!
1%
1-
12
#139940000000
0!
0%
b101 *
0-
02
b101 6
#139950000000
1!
1%
1-
12
#139960000000
0!
0%
b110 *
0-
02
b110 6
#139970000000
1!
1%
1-
12
#139980000000
0!
0%
b111 *
0-
02
b111 6
#139990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#140000000000
0!
0%
b0 *
0-
02
b0 6
#140010000000
1!
1%
1-
12
#140020000000
0!
0%
b1 *
0-
02
b1 6
#140030000000
1!
1%
1-
12
#140040000000
0!
0%
b10 *
0-
02
b10 6
#140050000000
1!
1%
1-
12
#140060000000
0!
0%
b11 *
0-
02
b11 6
#140070000000
1!
1%
1-
12
15
#140080000000
0!
0%
b100 *
0-
02
b100 6
#140090000000
1!
1%
1-
12
#140100000000
0!
0%
b101 *
0-
02
b101 6
#140110000000
1!
1%
1-
12
#140120000000
0!
0%
b110 *
0-
02
b110 6
#140130000000
1!
1%
1-
12
#140140000000
0!
0%
b111 *
0-
02
b111 6
#140150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#140160000000
0!
0%
b0 *
0-
02
b0 6
#140170000000
1!
1%
1-
12
#140180000000
0!
0%
b1 *
0-
02
b1 6
#140190000000
1!
1%
1-
12
#140200000000
0!
0%
b10 *
0-
02
b10 6
#140210000000
1!
1%
1-
12
#140220000000
0!
0%
b11 *
0-
02
b11 6
#140230000000
1!
1%
1-
12
15
#140240000000
0!
0%
b100 *
0-
02
b100 6
#140250000000
1!
1%
1-
12
#140260000000
0!
0%
b101 *
0-
02
b101 6
#140270000000
1!
1%
1-
12
#140280000000
0!
0%
b110 *
0-
02
b110 6
#140290000000
1!
1%
1-
12
#140300000000
0!
0%
b111 *
0-
02
b111 6
#140310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#140320000000
0!
0%
b0 *
0-
02
b0 6
#140330000000
1!
1%
1-
12
#140340000000
0!
0%
b1 *
0-
02
b1 6
#140350000000
1!
1%
1-
12
#140360000000
0!
0%
b10 *
0-
02
b10 6
#140370000000
1!
1%
1-
12
#140380000000
0!
0%
b11 *
0-
02
b11 6
#140390000000
1!
1%
1-
12
15
#140400000000
0!
0%
b100 *
0-
02
b100 6
#140410000000
1!
1%
1-
12
#140420000000
0!
0%
b101 *
0-
02
b101 6
#140430000000
1!
1%
1-
12
#140440000000
0!
0%
b110 *
0-
02
b110 6
#140450000000
1!
1%
1-
12
#140460000000
0!
0%
b111 *
0-
02
b111 6
#140470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#140480000000
0!
0%
b0 *
0-
02
b0 6
#140490000000
1!
1%
1-
12
#140500000000
0!
0%
b1 *
0-
02
b1 6
#140510000000
1!
1%
1-
12
#140520000000
0!
0%
b10 *
0-
02
b10 6
#140530000000
1!
1%
1-
12
#140540000000
0!
0%
b11 *
0-
02
b11 6
#140550000000
1!
1%
1-
12
15
#140560000000
0!
0%
b100 *
0-
02
b100 6
#140570000000
1!
1%
1-
12
#140580000000
0!
0%
b101 *
0-
02
b101 6
#140590000000
1!
1%
1-
12
#140600000000
0!
0%
b110 *
0-
02
b110 6
#140610000000
1!
1%
1-
12
#140620000000
0!
0%
b111 *
0-
02
b111 6
#140630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#140640000000
0!
0%
b0 *
0-
02
b0 6
#140650000000
1!
1%
1-
12
#140660000000
0!
0%
b1 *
0-
02
b1 6
#140670000000
1!
1%
1-
12
#140680000000
0!
0%
b10 *
0-
02
b10 6
#140690000000
1!
1%
1-
12
#140700000000
0!
0%
b11 *
0-
02
b11 6
#140710000000
1!
1%
1-
12
15
#140720000000
0!
0%
b100 *
0-
02
b100 6
#140730000000
1!
1%
1-
12
#140740000000
0!
0%
b101 *
0-
02
b101 6
#140750000000
1!
1%
1-
12
#140760000000
0!
0%
b110 *
0-
02
b110 6
#140770000000
1!
1%
1-
12
#140780000000
0!
0%
b111 *
0-
02
b111 6
#140790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#140800000000
0!
0%
b0 *
0-
02
b0 6
#140810000000
1!
1%
1-
12
#140820000000
0!
0%
b1 *
0-
02
b1 6
#140830000000
1!
1%
1-
12
#140840000000
0!
0%
b10 *
0-
02
b10 6
#140850000000
1!
1%
1-
12
#140860000000
0!
0%
b11 *
0-
02
b11 6
#140870000000
1!
1%
1-
12
15
#140880000000
0!
0%
b100 *
0-
02
b100 6
#140890000000
1!
1%
1-
12
#140900000000
0!
0%
b101 *
0-
02
b101 6
#140910000000
1!
1%
1-
12
#140920000000
0!
0%
b110 *
0-
02
b110 6
#140930000000
1!
1%
1-
12
#140940000000
0!
0%
b111 *
0-
02
b111 6
#140950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#140960000000
0!
0%
b0 *
0-
02
b0 6
#140970000000
1!
1%
1-
12
#140980000000
0!
0%
b1 *
0-
02
b1 6
#140990000000
1!
1%
1-
12
#141000000000
0!
0%
b10 *
0-
02
b10 6
#141010000000
1!
1%
1-
12
#141020000000
0!
0%
b11 *
0-
02
b11 6
#141030000000
1!
1%
1-
12
15
#141040000000
0!
0%
b100 *
0-
02
b100 6
#141050000000
1!
1%
1-
12
#141060000000
0!
0%
b101 *
0-
02
b101 6
#141070000000
1!
1%
1-
12
#141080000000
0!
0%
b110 *
0-
02
b110 6
#141090000000
1!
1%
1-
12
#141100000000
0!
0%
b111 *
0-
02
b111 6
#141110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#141120000000
0!
0%
b0 *
0-
02
b0 6
#141130000000
1!
1%
1-
12
#141140000000
0!
0%
b1 *
0-
02
b1 6
#141150000000
1!
1%
1-
12
#141160000000
0!
0%
b10 *
0-
02
b10 6
#141170000000
1!
1%
1-
12
#141180000000
0!
0%
b11 *
0-
02
b11 6
#141190000000
1!
1%
1-
12
15
#141200000000
0!
0%
b100 *
0-
02
b100 6
#141210000000
1!
1%
1-
12
#141220000000
0!
0%
b101 *
0-
02
b101 6
#141230000000
1!
1%
1-
12
#141240000000
0!
0%
b110 *
0-
02
b110 6
#141250000000
1!
1%
1-
12
#141260000000
0!
0%
b111 *
0-
02
b111 6
#141270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#141280000000
0!
0%
b0 *
0-
02
b0 6
#141290000000
1!
1%
1-
12
#141300000000
0!
0%
b1 *
0-
02
b1 6
#141310000000
1!
1%
1-
12
#141320000000
0!
0%
b10 *
0-
02
b10 6
#141330000000
1!
1%
1-
12
#141340000000
0!
0%
b11 *
0-
02
b11 6
#141350000000
1!
1%
1-
12
15
#141360000000
0!
0%
b100 *
0-
02
b100 6
#141370000000
1!
1%
1-
12
#141380000000
0!
0%
b101 *
0-
02
b101 6
#141390000000
1!
1%
1-
12
#141400000000
0!
0%
b110 *
0-
02
b110 6
#141410000000
1!
1%
1-
12
#141420000000
0!
0%
b111 *
0-
02
b111 6
#141430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#141440000000
0!
0%
b0 *
0-
02
b0 6
#141450000000
1!
1%
1-
12
#141460000000
0!
0%
b1 *
0-
02
b1 6
#141470000000
1!
1%
1-
12
#141480000000
0!
0%
b10 *
0-
02
b10 6
#141490000000
1!
1%
1-
12
#141500000000
0!
0%
b11 *
0-
02
b11 6
#141510000000
1!
1%
1-
12
15
#141520000000
0!
0%
b100 *
0-
02
b100 6
#141530000000
1!
1%
1-
12
#141540000000
0!
0%
b101 *
0-
02
b101 6
#141550000000
1!
1%
1-
12
#141560000000
0!
0%
b110 *
0-
02
b110 6
#141570000000
1!
1%
1-
12
#141580000000
0!
0%
b111 *
0-
02
b111 6
#141590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#141600000000
0!
0%
b0 *
0-
02
b0 6
#141610000000
1!
1%
1-
12
#141620000000
0!
0%
b1 *
0-
02
b1 6
#141630000000
1!
1%
1-
12
#141640000000
0!
0%
b10 *
0-
02
b10 6
#141650000000
1!
1%
1-
12
#141660000000
0!
0%
b11 *
0-
02
b11 6
#141670000000
1!
1%
1-
12
15
#141680000000
0!
0%
b100 *
0-
02
b100 6
#141690000000
1!
1%
1-
12
#141700000000
0!
0%
b101 *
0-
02
b101 6
#141710000000
1!
1%
1-
12
#141720000000
0!
0%
b110 *
0-
02
b110 6
#141730000000
1!
1%
1-
12
#141740000000
0!
0%
b111 *
0-
02
b111 6
#141750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#141760000000
0!
0%
b0 *
0-
02
b0 6
#141770000000
1!
1%
1-
12
#141780000000
0!
0%
b1 *
0-
02
b1 6
#141790000000
1!
1%
1-
12
#141800000000
0!
0%
b10 *
0-
02
b10 6
#141810000000
1!
1%
1-
12
#141820000000
0!
0%
b11 *
0-
02
b11 6
#141830000000
1!
1%
1-
12
15
#141840000000
0!
0%
b100 *
0-
02
b100 6
#141850000000
1!
1%
1-
12
#141860000000
0!
0%
b101 *
0-
02
b101 6
#141870000000
1!
1%
1-
12
#141880000000
0!
0%
b110 *
0-
02
b110 6
#141890000000
1!
1%
1-
12
#141900000000
0!
0%
b111 *
0-
02
b111 6
#141910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#141920000000
0!
0%
b0 *
0-
02
b0 6
#141930000000
1!
1%
1-
12
#141940000000
0!
0%
b1 *
0-
02
b1 6
#141950000000
1!
1%
1-
12
#141960000000
0!
0%
b10 *
0-
02
b10 6
#141970000000
1!
1%
1-
12
#141980000000
0!
0%
b11 *
0-
02
b11 6
#141990000000
1!
1%
1-
12
15
#142000000000
0!
0%
b100 *
0-
02
b100 6
#142010000000
1!
1%
1-
12
#142020000000
0!
0%
b101 *
0-
02
b101 6
#142030000000
1!
1%
1-
12
#142040000000
0!
0%
b110 *
0-
02
b110 6
#142050000000
1!
1%
1-
12
#142060000000
0!
0%
b111 *
0-
02
b111 6
#142070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#142080000000
0!
0%
b0 *
0-
02
b0 6
#142090000000
1!
1%
1-
12
#142100000000
0!
0%
b1 *
0-
02
b1 6
#142110000000
1!
1%
1-
12
#142120000000
0!
0%
b10 *
0-
02
b10 6
#142130000000
1!
1%
1-
12
#142140000000
0!
0%
b11 *
0-
02
b11 6
#142150000000
1!
1%
1-
12
15
#142160000000
0!
0%
b100 *
0-
02
b100 6
#142170000000
1!
1%
1-
12
#142180000000
0!
0%
b101 *
0-
02
b101 6
#142190000000
1!
1%
1-
12
#142200000000
0!
0%
b110 *
0-
02
b110 6
#142210000000
1!
1%
1-
12
#142220000000
0!
0%
b111 *
0-
02
b111 6
#142230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#142240000000
0!
0%
b0 *
0-
02
b0 6
#142250000000
1!
1%
1-
12
#142260000000
0!
0%
b1 *
0-
02
b1 6
#142270000000
1!
1%
1-
12
#142280000000
0!
0%
b10 *
0-
02
b10 6
#142290000000
1!
1%
1-
12
#142300000000
0!
0%
b11 *
0-
02
b11 6
#142310000000
1!
1%
1-
12
15
#142320000000
0!
0%
b100 *
0-
02
b100 6
#142330000000
1!
1%
1-
12
#142340000000
0!
0%
b101 *
0-
02
b101 6
#142350000000
1!
1%
1-
12
#142360000000
0!
0%
b110 *
0-
02
b110 6
#142370000000
1!
1%
1-
12
#142380000000
0!
0%
b111 *
0-
02
b111 6
#142390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#142400000000
0!
0%
b0 *
0-
02
b0 6
#142410000000
1!
1%
1-
12
#142420000000
0!
0%
b1 *
0-
02
b1 6
#142430000000
1!
1%
1-
12
#142440000000
0!
0%
b10 *
0-
02
b10 6
#142450000000
1!
1%
1-
12
#142460000000
0!
0%
b11 *
0-
02
b11 6
#142470000000
1!
1%
1-
12
15
#142480000000
0!
0%
b100 *
0-
02
b100 6
#142490000000
1!
1%
1-
12
#142500000000
0!
0%
b101 *
0-
02
b101 6
#142510000000
1!
1%
1-
12
#142520000000
0!
0%
b110 *
0-
02
b110 6
#142530000000
1!
1%
1-
12
#142540000000
0!
0%
b111 *
0-
02
b111 6
#142550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#142560000000
0!
0%
b0 *
0-
02
b0 6
#142570000000
1!
1%
1-
12
#142580000000
0!
0%
b1 *
0-
02
b1 6
#142590000000
1!
1%
1-
12
#142600000000
0!
0%
b10 *
0-
02
b10 6
#142610000000
1!
1%
1-
12
#142620000000
0!
0%
b11 *
0-
02
b11 6
#142630000000
1!
1%
1-
12
15
#142640000000
0!
0%
b100 *
0-
02
b100 6
#142650000000
1!
1%
1-
12
#142660000000
0!
0%
b101 *
0-
02
b101 6
#142670000000
1!
1%
1-
12
#142680000000
0!
0%
b110 *
0-
02
b110 6
#142690000000
1!
1%
1-
12
#142700000000
0!
0%
b111 *
0-
02
b111 6
#142710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#142720000000
0!
0%
b0 *
0-
02
b0 6
#142730000000
1!
1%
1-
12
#142740000000
0!
0%
b1 *
0-
02
b1 6
#142750000000
1!
1%
1-
12
#142760000000
0!
0%
b10 *
0-
02
b10 6
#142770000000
1!
1%
1-
12
#142780000000
0!
0%
b11 *
0-
02
b11 6
#142790000000
1!
1%
1-
12
15
#142800000000
0!
0%
b100 *
0-
02
b100 6
#142810000000
1!
1%
1-
12
#142820000000
0!
0%
b101 *
0-
02
b101 6
#142830000000
1!
1%
1-
12
#142840000000
0!
0%
b110 *
0-
02
b110 6
#142850000000
1!
1%
1-
12
#142860000000
0!
0%
b111 *
0-
02
b111 6
#142870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#142880000000
0!
0%
b0 *
0-
02
b0 6
#142890000000
1!
1%
1-
12
#142900000000
0!
0%
b1 *
0-
02
b1 6
#142910000000
1!
1%
1-
12
#142920000000
0!
0%
b10 *
0-
02
b10 6
#142930000000
1!
1%
1-
12
#142940000000
0!
0%
b11 *
0-
02
b11 6
#142950000000
1!
1%
1-
12
15
#142960000000
0!
0%
b100 *
0-
02
b100 6
#142970000000
1!
1%
1-
12
#142980000000
0!
0%
b101 *
0-
02
b101 6
#142990000000
1!
1%
1-
12
#143000000000
0!
0%
b110 *
0-
02
b110 6
#143010000000
1!
1%
1-
12
#143020000000
0!
0%
b111 *
0-
02
b111 6
#143030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#143040000000
0!
0%
b0 *
0-
02
b0 6
#143050000000
1!
1%
1-
12
#143060000000
0!
0%
b1 *
0-
02
b1 6
#143070000000
1!
1%
1-
12
#143080000000
0!
0%
b10 *
0-
02
b10 6
#143090000000
1!
1%
1-
12
#143100000000
0!
0%
b11 *
0-
02
b11 6
#143110000000
1!
1%
1-
12
15
#143120000000
0!
0%
b100 *
0-
02
b100 6
#143130000000
1!
1%
1-
12
#143140000000
0!
0%
b101 *
0-
02
b101 6
#143150000000
1!
1%
1-
12
#143160000000
0!
0%
b110 *
0-
02
b110 6
#143170000000
1!
1%
1-
12
#143180000000
0!
0%
b111 *
0-
02
b111 6
#143190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#143200000000
0!
0%
b0 *
0-
02
b0 6
#143210000000
1!
1%
1-
12
#143220000000
0!
0%
b1 *
0-
02
b1 6
#143230000000
1!
1%
1-
12
#143240000000
0!
0%
b10 *
0-
02
b10 6
#143250000000
1!
1%
1-
12
#143260000000
0!
0%
b11 *
0-
02
b11 6
#143270000000
1!
1%
1-
12
15
#143280000000
0!
0%
b100 *
0-
02
b100 6
#143290000000
1!
1%
1-
12
#143300000000
0!
0%
b101 *
0-
02
b101 6
#143310000000
1!
1%
1-
12
#143320000000
0!
0%
b110 *
0-
02
b110 6
#143330000000
1!
1%
1-
12
#143340000000
0!
0%
b111 *
0-
02
b111 6
#143350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#143360000000
0!
0%
b0 *
0-
02
b0 6
#143370000000
1!
1%
1-
12
#143380000000
0!
0%
b1 *
0-
02
b1 6
#143390000000
1!
1%
1-
12
#143400000000
0!
0%
b10 *
0-
02
b10 6
#143410000000
1!
1%
1-
12
#143420000000
0!
0%
b11 *
0-
02
b11 6
#143430000000
1!
1%
1-
12
15
#143440000000
0!
0%
b100 *
0-
02
b100 6
#143450000000
1!
1%
1-
12
#143460000000
0!
0%
b101 *
0-
02
b101 6
#143470000000
1!
1%
1-
12
#143480000000
0!
0%
b110 *
0-
02
b110 6
#143490000000
1!
1%
1-
12
#143500000000
0!
0%
b111 *
0-
02
b111 6
#143510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#143520000000
0!
0%
b0 *
0-
02
b0 6
#143530000000
1!
1%
1-
12
#143540000000
0!
0%
b1 *
0-
02
b1 6
#143550000000
1!
1%
1-
12
#143560000000
0!
0%
b10 *
0-
02
b10 6
#143570000000
1!
1%
1-
12
#143580000000
0!
0%
b11 *
0-
02
b11 6
#143590000000
1!
1%
1-
12
15
#143600000000
0!
0%
b100 *
0-
02
b100 6
#143610000000
1!
1%
1-
12
#143620000000
0!
0%
b101 *
0-
02
b101 6
#143630000000
1!
1%
1-
12
#143640000000
0!
0%
b110 *
0-
02
b110 6
#143650000000
1!
1%
1-
12
#143660000000
0!
0%
b111 *
0-
02
b111 6
#143670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#143680000000
0!
0%
b0 *
0-
02
b0 6
#143690000000
1!
1%
1-
12
#143700000000
0!
0%
b1 *
0-
02
b1 6
#143710000000
1!
1%
1-
12
#143720000000
0!
0%
b10 *
0-
02
b10 6
#143730000000
1!
1%
1-
12
#143740000000
0!
0%
b11 *
0-
02
b11 6
#143750000000
1!
1%
1-
12
15
#143760000000
0!
0%
b100 *
0-
02
b100 6
#143770000000
1!
1%
1-
12
#143780000000
0!
0%
b101 *
0-
02
b101 6
#143790000000
1!
1%
1-
12
#143800000000
0!
0%
b110 *
0-
02
b110 6
#143810000000
1!
1%
1-
12
#143820000000
0!
0%
b111 *
0-
02
b111 6
#143830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#143840000000
0!
0%
b0 *
0-
02
b0 6
#143850000000
1!
1%
1-
12
#143860000000
0!
0%
b1 *
0-
02
b1 6
#143870000000
1!
1%
1-
12
#143880000000
0!
0%
b10 *
0-
02
b10 6
#143890000000
1!
1%
1-
12
#143900000000
0!
0%
b11 *
0-
02
b11 6
#143910000000
1!
1%
1-
12
15
#143920000000
0!
0%
b100 *
0-
02
b100 6
#143930000000
1!
1%
1-
12
#143940000000
0!
0%
b101 *
0-
02
b101 6
#143950000000
1!
1%
1-
12
#143960000000
0!
0%
b110 *
0-
02
b110 6
#143970000000
1!
1%
1-
12
#143980000000
0!
0%
b111 *
0-
02
b111 6
#143990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#144000000000
0!
0%
b0 *
0-
02
b0 6
#144010000000
1!
1%
1-
12
#144020000000
0!
0%
b1 *
0-
02
b1 6
#144030000000
1!
1%
1-
12
#144040000000
0!
0%
b10 *
0-
02
b10 6
#144050000000
1!
1%
1-
12
#144060000000
0!
0%
b11 *
0-
02
b11 6
#144070000000
1!
1%
1-
12
15
#144080000000
0!
0%
b100 *
0-
02
b100 6
#144090000000
1!
1%
1-
12
#144100000000
0!
0%
b101 *
0-
02
b101 6
#144110000000
1!
1%
1-
12
#144120000000
0!
0%
b110 *
0-
02
b110 6
#144130000000
1!
1%
1-
12
#144140000000
0!
0%
b111 *
0-
02
b111 6
#144150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#144160000000
0!
0%
b0 *
0-
02
b0 6
#144170000000
1!
1%
1-
12
#144180000000
0!
0%
b1 *
0-
02
b1 6
#144190000000
1!
1%
1-
12
#144200000000
0!
0%
b10 *
0-
02
b10 6
#144210000000
1!
1%
1-
12
#144220000000
0!
0%
b11 *
0-
02
b11 6
#144230000000
1!
1%
1-
12
15
#144240000000
0!
0%
b100 *
0-
02
b100 6
#144250000000
1!
1%
1-
12
#144260000000
0!
0%
b101 *
0-
02
b101 6
#144270000000
1!
1%
1-
12
#144280000000
0!
0%
b110 *
0-
02
b110 6
#144290000000
1!
1%
1-
12
#144300000000
0!
0%
b111 *
0-
02
b111 6
#144310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#144320000000
0!
0%
b0 *
0-
02
b0 6
#144330000000
1!
1%
1-
12
#144340000000
0!
0%
b1 *
0-
02
b1 6
#144350000000
1!
1%
1-
12
#144360000000
0!
0%
b10 *
0-
02
b10 6
#144370000000
1!
1%
1-
12
#144380000000
0!
0%
b11 *
0-
02
b11 6
#144390000000
1!
1%
1-
12
15
#144400000000
0!
0%
b100 *
0-
02
b100 6
#144410000000
1!
1%
1-
12
#144420000000
0!
0%
b101 *
0-
02
b101 6
#144430000000
1!
1%
1-
12
#144440000000
0!
0%
b110 *
0-
02
b110 6
#144450000000
1!
1%
1-
12
#144460000000
0!
0%
b111 *
0-
02
b111 6
#144470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#144480000000
0!
0%
b0 *
0-
02
b0 6
#144490000000
1!
1%
1-
12
#144500000000
0!
0%
b1 *
0-
02
b1 6
#144510000000
1!
1%
1-
12
#144520000000
0!
0%
b10 *
0-
02
b10 6
#144530000000
1!
1%
1-
12
#144540000000
0!
0%
b11 *
0-
02
b11 6
#144550000000
1!
1%
1-
12
15
#144560000000
0!
0%
b100 *
0-
02
b100 6
#144570000000
1!
1%
1-
12
#144580000000
0!
0%
b101 *
0-
02
b101 6
#144590000000
1!
1%
1-
12
#144600000000
0!
0%
b110 *
0-
02
b110 6
#144610000000
1!
1%
1-
12
#144620000000
0!
0%
b111 *
0-
02
b111 6
#144630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#144640000000
0!
0%
b0 *
0-
02
b0 6
#144650000000
1!
1%
1-
12
#144660000000
0!
0%
b1 *
0-
02
b1 6
#144670000000
1!
1%
1-
12
#144680000000
0!
0%
b10 *
0-
02
b10 6
#144690000000
1!
1%
1-
12
#144700000000
0!
0%
b11 *
0-
02
b11 6
#144710000000
1!
1%
1-
12
15
#144720000000
0!
0%
b100 *
0-
02
b100 6
#144730000000
1!
1%
1-
12
#144740000000
0!
0%
b101 *
0-
02
b101 6
#144750000000
1!
1%
1-
12
#144760000000
0!
0%
b110 *
0-
02
b110 6
#144770000000
1!
1%
1-
12
#144780000000
0!
0%
b111 *
0-
02
b111 6
#144790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#144800000000
0!
0%
b0 *
0-
02
b0 6
#144810000000
1!
1%
1-
12
#144820000000
0!
0%
b1 *
0-
02
b1 6
#144830000000
1!
1%
1-
12
#144840000000
0!
0%
b10 *
0-
02
b10 6
#144850000000
1!
1%
1-
12
#144860000000
0!
0%
b11 *
0-
02
b11 6
#144870000000
1!
1%
1-
12
15
#144880000000
0!
0%
b100 *
0-
02
b100 6
#144890000000
1!
1%
1-
12
#144900000000
0!
0%
b101 *
0-
02
b101 6
#144910000000
1!
1%
1-
12
#144920000000
0!
0%
b110 *
0-
02
b110 6
#144930000000
1!
1%
1-
12
#144940000000
0!
0%
b111 *
0-
02
b111 6
#144950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#144960000000
0!
0%
b0 *
0-
02
b0 6
#144970000000
1!
1%
1-
12
#144980000000
0!
0%
b1 *
0-
02
b1 6
#144990000000
1!
1%
1-
12
#145000000000
0!
0%
b10 *
0-
02
b10 6
#145010000000
1!
1%
1-
12
#145020000000
0!
0%
b11 *
0-
02
b11 6
#145030000000
1!
1%
1-
12
15
#145040000000
0!
0%
b100 *
0-
02
b100 6
#145050000000
1!
1%
1-
12
#145060000000
0!
0%
b101 *
0-
02
b101 6
#145070000000
1!
1%
1-
12
#145080000000
0!
0%
b110 *
0-
02
b110 6
#145090000000
1!
1%
1-
12
#145100000000
0!
0%
b111 *
0-
02
b111 6
#145110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#145120000000
0!
0%
b0 *
0-
02
b0 6
#145130000000
1!
1%
1-
12
#145140000000
0!
0%
b1 *
0-
02
b1 6
#145150000000
1!
1%
1-
12
#145160000000
0!
0%
b10 *
0-
02
b10 6
#145170000000
1!
1%
1-
12
#145180000000
0!
0%
b11 *
0-
02
b11 6
#145190000000
1!
1%
1-
12
15
#145200000000
0!
0%
b100 *
0-
02
b100 6
#145210000000
1!
1%
1-
12
#145220000000
0!
0%
b101 *
0-
02
b101 6
#145230000000
1!
1%
1-
12
#145240000000
0!
0%
b110 *
0-
02
b110 6
#145250000000
1!
1%
1-
12
#145260000000
0!
0%
b111 *
0-
02
b111 6
#145270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#145280000000
0!
0%
b0 *
0-
02
b0 6
#145290000000
1!
1%
1-
12
#145300000000
0!
0%
b1 *
0-
02
b1 6
#145310000000
1!
1%
1-
12
#145320000000
0!
0%
b10 *
0-
02
b10 6
#145330000000
1!
1%
1-
12
#145340000000
0!
0%
b11 *
0-
02
b11 6
#145350000000
1!
1%
1-
12
15
#145360000000
0!
0%
b100 *
0-
02
b100 6
#145370000000
1!
1%
1-
12
#145380000000
0!
0%
b101 *
0-
02
b101 6
#145390000000
1!
1%
1-
12
#145400000000
0!
0%
b110 *
0-
02
b110 6
#145410000000
1!
1%
1-
12
#145420000000
0!
0%
b111 *
0-
02
b111 6
#145430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#145440000000
0!
0%
b0 *
0-
02
b0 6
#145450000000
1!
1%
1-
12
#145460000000
0!
0%
b1 *
0-
02
b1 6
#145470000000
1!
1%
1-
12
#145480000000
0!
0%
b10 *
0-
02
b10 6
#145490000000
1!
1%
1-
12
#145500000000
0!
0%
b11 *
0-
02
b11 6
#145510000000
1!
1%
1-
12
15
#145520000000
0!
0%
b100 *
0-
02
b100 6
#145530000000
1!
1%
1-
12
#145540000000
0!
0%
b101 *
0-
02
b101 6
#145550000000
1!
1%
1-
12
#145560000000
0!
0%
b110 *
0-
02
b110 6
#145570000000
1!
1%
1-
12
#145580000000
0!
0%
b111 *
0-
02
b111 6
#145590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#145600000000
0!
0%
b0 *
0-
02
b0 6
#145610000000
1!
1%
1-
12
#145620000000
0!
0%
b1 *
0-
02
b1 6
#145630000000
1!
1%
1-
12
#145640000000
0!
0%
b10 *
0-
02
b10 6
#145650000000
1!
1%
1-
12
#145660000000
0!
0%
b11 *
0-
02
b11 6
#145670000000
1!
1%
1-
12
15
#145680000000
0!
0%
b100 *
0-
02
b100 6
#145690000000
1!
1%
1-
12
#145700000000
0!
0%
b101 *
0-
02
b101 6
#145710000000
1!
1%
1-
12
#145720000000
0!
0%
b110 *
0-
02
b110 6
#145730000000
1!
1%
1-
12
#145740000000
0!
0%
b111 *
0-
02
b111 6
#145750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#145760000000
0!
0%
b0 *
0-
02
b0 6
#145770000000
1!
1%
1-
12
#145780000000
0!
0%
b1 *
0-
02
b1 6
#145790000000
1!
1%
1-
12
#145800000000
0!
0%
b10 *
0-
02
b10 6
#145810000000
1!
1%
1-
12
#145820000000
0!
0%
b11 *
0-
02
b11 6
#145830000000
1!
1%
1-
12
15
#145840000000
0!
0%
b100 *
0-
02
b100 6
#145850000000
1!
1%
1-
12
#145860000000
0!
0%
b101 *
0-
02
b101 6
#145870000000
1!
1%
1-
12
#145880000000
0!
0%
b110 *
0-
02
b110 6
#145890000000
1!
1%
1-
12
#145900000000
0!
0%
b111 *
0-
02
b111 6
#145910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#145920000000
0!
0%
b0 *
0-
02
b0 6
#145930000000
1!
1%
1-
12
#145940000000
0!
0%
b1 *
0-
02
b1 6
#145950000000
1!
1%
1-
12
#145960000000
0!
0%
b10 *
0-
02
b10 6
#145970000000
1!
1%
1-
12
#145980000000
0!
0%
b11 *
0-
02
b11 6
#145990000000
1!
1%
1-
12
15
#146000000000
0!
0%
b100 *
0-
02
b100 6
#146010000000
1!
1%
1-
12
#146020000000
0!
0%
b101 *
0-
02
b101 6
#146030000000
1!
1%
1-
12
#146040000000
0!
0%
b110 *
0-
02
b110 6
#146050000000
1!
1%
1-
12
#146060000000
0!
0%
b111 *
0-
02
b111 6
#146070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#146080000000
0!
0%
b0 *
0-
02
b0 6
#146090000000
1!
1%
1-
12
#146100000000
0!
0%
b1 *
0-
02
b1 6
#146110000000
1!
1%
1-
12
#146120000000
0!
0%
b10 *
0-
02
b10 6
#146130000000
1!
1%
1-
12
#146140000000
0!
0%
b11 *
0-
02
b11 6
#146150000000
1!
1%
1-
12
15
#146160000000
0!
0%
b100 *
0-
02
b100 6
#146170000000
1!
1%
1-
12
#146180000000
0!
0%
b101 *
0-
02
b101 6
#146190000000
1!
1%
1-
12
#146200000000
0!
0%
b110 *
0-
02
b110 6
#146210000000
1!
1%
1-
12
#146220000000
0!
0%
b111 *
0-
02
b111 6
#146230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#146240000000
0!
0%
b0 *
0-
02
b0 6
#146250000000
1!
1%
1-
12
#146260000000
0!
0%
b1 *
0-
02
b1 6
#146270000000
1!
1%
1-
12
#146280000000
0!
0%
b10 *
0-
02
b10 6
#146290000000
1!
1%
1-
12
#146300000000
0!
0%
b11 *
0-
02
b11 6
#146310000000
1!
1%
1-
12
15
#146320000000
0!
0%
b100 *
0-
02
b100 6
#146330000000
1!
1%
1-
12
#146340000000
0!
0%
b101 *
0-
02
b101 6
#146350000000
1!
1%
1-
12
#146360000000
0!
0%
b110 *
0-
02
b110 6
#146370000000
1!
1%
1-
12
#146380000000
0!
0%
b111 *
0-
02
b111 6
#146390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#146400000000
0!
0%
b0 *
0-
02
b0 6
#146410000000
1!
1%
1-
12
#146420000000
0!
0%
b1 *
0-
02
b1 6
#146430000000
1!
1%
1-
12
#146440000000
0!
0%
b10 *
0-
02
b10 6
#146450000000
1!
1%
1-
12
#146460000000
0!
0%
b11 *
0-
02
b11 6
#146470000000
1!
1%
1-
12
15
#146480000000
0!
0%
b100 *
0-
02
b100 6
#146490000000
1!
1%
1-
12
#146500000000
0!
0%
b101 *
0-
02
b101 6
#146510000000
1!
1%
1-
12
#146520000000
0!
0%
b110 *
0-
02
b110 6
#146530000000
1!
1%
1-
12
#146540000000
0!
0%
b111 *
0-
02
b111 6
#146550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#146560000000
0!
0%
b0 *
0-
02
b0 6
#146570000000
1!
1%
1-
12
#146580000000
0!
0%
b1 *
0-
02
b1 6
#146590000000
1!
1%
1-
12
#146600000000
0!
0%
b10 *
0-
02
b10 6
#146610000000
1!
1%
1-
12
#146620000000
0!
0%
b11 *
0-
02
b11 6
#146630000000
1!
1%
1-
12
15
#146640000000
0!
0%
b100 *
0-
02
b100 6
#146650000000
1!
1%
1-
12
#146660000000
0!
0%
b101 *
0-
02
b101 6
#146670000000
1!
1%
1-
12
#146680000000
0!
0%
b110 *
0-
02
b110 6
#146690000000
1!
1%
1-
12
#146700000000
0!
0%
b111 *
0-
02
b111 6
#146710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#146720000000
0!
0%
b0 *
0-
02
b0 6
#146730000000
1!
1%
1-
12
#146740000000
0!
0%
b1 *
0-
02
b1 6
#146750000000
1!
1%
1-
12
#146760000000
0!
0%
b10 *
0-
02
b10 6
#146770000000
1!
1%
1-
12
#146780000000
0!
0%
b11 *
0-
02
b11 6
#146790000000
1!
1%
1-
12
15
#146800000000
0!
0%
b100 *
0-
02
b100 6
#146810000000
1!
1%
1-
12
#146820000000
0!
0%
b101 *
0-
02
b101 6
#146830000000
1!
1%
1-
12
#146840000000
0!
0%
b110 *
0-
02
b110 6
#146850000000
1!
1%
1-
12
#146860000000
0!
0%
b111 *
0-
02
b111 6
#146870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#146880000000
0!
0%
b0 *
0-
02
b0 6
#146890000000
1!
1%
1-
12
#146900000000
0!
0%
b1 *
0-
02
b1 6
#146910000000
1!
1%
1-
12
#146920000000
0!
0%
b10 *
0-
02
b10 6
#146930000000
1!
1%
1-
12
#146940000000
0!
0%
b11 *
0-
02
b11 6
#146950000000
1!
1%
1-
12
15
#146960000000
0!
0%
b100 *
0-
02
b100 6
#146970000000
1!
1%
1-
12
#146980000000
0!
0%
b101 *
0-
02
b101 6
#146990000000
1!
1%
1-
12
#147000000000
0!
0%
b110 *
0-
02
b110 6
#147010000000
1!
1%
1-
12
#147020000000
0!
0%
b111 *
0-
02
b111 6
#147030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#147040000000
0!
0%
b0 *
0-
02
b0 6
#147050000000
1!
1%
1-
12
#147060000000
0!
0%
b1 *
0-
02
b1 6
#147070000000
1!
1%
1-
12
#147080000000
0!
0%
b10 *
0-
02
b10 6
#147090000000
1!
1%
1-
12
#147100000000
0!
0%
b11 *
0-
02
b11 6
#147110000000
1!
1%
1-
12
15
#147120000000
0!
0%
b100 *
0-
02
b100 6
#147130000000
1!
1%
1-
12
#147140000000
0!
0%
b101 *
0-
02
b101 6
#147150000000
1!
1%
1-
12
#147160000000
0!
0%
b110 *
0-
02
b110 6
#147170000000
1!
1%
1-
12
#147180000000
0!
0%
b111 *
0-
02
b111 6
#147190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#147200000000
0!
0%
b0 *
0-
02
b0 6
#147210000000
1!
1%
1-
12
#147220000000
0!
0%
b1 *
0-
02
b1 6
#147230000000
1!
1%
1-
12
#147240000000
0!
0%
b10 *
0-
02
b10 6
#147250000000
1!
1%
1-
12
#147260000000
0!
0%
b11 *
0-
02
b11 6
#147270000000
1!
1%
1-
12
15
#147280000000
0!
0%
b100 *
0-
02
b100 6
#147290000000
1!
1%
1-
12
#147300000000
0!
0%
b101 *
0-
02
b101 6
#147310000000
1!
1%
1-
12
#147320000000
0!
0%
b110 *
0-
02
b110 6
#147330000000
1!
1%
1-
12
#147340000000
0!
0%
b111 *
0-
02
b111 6
#147350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#147360000000
0!
0%
b0 *
0-
02
b0 6
#147370000000
1!
1%
1-
12
#147380000000
0!
0%
b1 *
0-
02
b1 6
#147390000000
1!
1%
1-
12
#147400000000
0!
0%
b10 *
0-
02
b10 6
#147410000000
1!
1%
1-
12
#147420000000
0!
0%
b11 *
0-
02
b11 6
#147430000000
1!
1%
1-
12
15
#147440000000
0!
0%
b100 *
0-
02
b100 6
#147450000000
1!
1%
1-
12
#147460000000
0!
0%
b101 *
0-
02
b101 6
#147470000000
1!
1%
1-
12
#147480000000
0!
0%
b110 *
0-
02
b110 6
#147490000000
1!
1%
1-
12
#147500000000
0!
0%
b111 *
0-
02
b111 6
#147510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#147520000000
0!
0%
b0 *
0-
02
b0 6
#147530000000
1!
1%
1-
12
#147540000000
0!
0%
b1 *
0-
02
b1 6
#147550000000
1!
1%
1-
12
#147560000000
0!
0%
b10 *
0-
02
b10 6
#147570000000
1!
1%
1-
12
#147580000000
0!
0%
b11 *
0-
02
b11 6
#147590000000
1!
1%
1-
12
15
#147600000000
0!
0%
b100 *
0-
02
b100 6
#147610000000
1!
1%
1-
12
#147620000000
0!
0%
b101 *
0-
02
b101 6
#147630000000
1!
1%
1-
12
#147640000000
0!
0%
b110 *
0-
02
b110 6
#147650000000
1!
1%
1-
12
#147660000000
0!
0%
b111 *
0-
02
b111 6
#147670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#147680000000
0!
0%
b0 *
0-
02
b0 6
#147690000000
1!
1%
1-
12
#147700000000
0!
0%
b1 *
0-
02
b1 6
#147710000000
1!
1%
1-
12
#147720000000
0!
0%
b10 *
0-
02
b10 6
#147730000000
1!
1%
1-
12
#147740000000
0!
0%
b11 *
0-
02
b11 6
#147750000000
1!
1%
1-
12
15
#147760000000
0!
0%
b100 *
0-
02
b100 6
#147770000000
1!
1%
1-
12
#147780000000
0!
0%
b101 *
0-
02
b101 6
#147790000000
1!
1%
1-
12
#147800000000
0!
0%
b110 *
0-
02
b110 6
#147810000000
1!
1%
1-
12
#147820000000
0!
0%
b111 *
0-
02
b111 6
#147830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#147840000000
0!
0%
b0 *
0-
02
b0 6
#147850000000
1!
1%
1-
12
#147860000000
0!
0%
b1 *
0-
02
b1 6
#147870000000
1!
1%
1-
12
#147880000000
0!
0%
b10 *
0-
02
b10 6
#147890000000
1!
1%
1-
12
#147900000000
0!
0%
b11 *
0-
02
b11 6
#147910000000
1!
1%
1-
12
15
#147920000000
0!
0%
b100 *
0-
02
b100 6
#147930000000
1!
1%
1-
12
#147940000000
0!
0%
b101 *
0-
02
b101 6
#147950000000
1!
1%
1-
12
#147960000000
0!
0%
b110 *
0-
02
b110 6
#147970000000
1!
1%
1-
12
#147980000000
0!
0%
b111 *
0-
02
b111 6
#147990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#148000000000
0!
0%
b0 *
0-
02
b0 6
#148010000000
1!
1%
1-
12
#148020000000
0!
0%
b1 *
0-
02
b1 6
#148030000000
1!
1%
1-
12
#148040000000
0!
0%
b10 *
0-
02
b10 6
#148050000000
1!
1%
1-
12
#148060000000
0!
0%
b11 *
0-
02
b11 6
#148070000000
1!
1%
1-
12
15
#148080000000
0!
0%
b100 *
0-
02
b100 6
#148090000000
1!
1%
1-
12
#148100000000
0!
0%
b101 *
0-
02
b101 6
#148110000000
1!
1%
1-
12
#148120000000
0!
0%
b110 *
0-
02
b110 6
#148130000000
1!
1%
1-
12
#148140000000
0!
0%
b111 *
0-
02
b111 6
#148150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#148160000000
0!
0%
b0 *
0-
02
b0 6
#148170000000
1!
1%
1-
12
#148180000000
0!
0%
b1 *
0-
02
b1 6
#148190000000
1!
1%
1-
12
#148200000000
0!
0%
b10 *
0-
02
b10 6
#148210000000
1!
1%
1-
12
#148220000000
0!
0%
b11 *
0-
02
b11 6
#148230000000
1!
1%
1-
12
15
#148240000000
0!
0%
b100 *
0-
02
b100 6
#148250000000
1!
1%
1-
12
#148260000000
0!
0%
b101 *
0-
02
b101 6
#148270000000
1!
1%
1-
12
#148280000000
0!
0%
b110 *
0-
02
b110 6
#148290000000
1!
1%
1-
12
#148300000000
0!
0%
b111 *
0-
02
b111 6
#148310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#148320000000
0!
0%
b0 *
0-
02
b0 6
#148330000000
1!
1%
1-
12
#148340000000
0!
0%
b1 *
0-
02
b1 6
#148350000000
1!
1%
1-
12
#148360000000
0!
0%
b10 *
0-
02
b10 6
#148370000000
1!
1%
1-
12
#148380000000
0!
0%
b11 *
0-
02
b11 6
#148390000000
1!
1%
1-
12
15
#148400000000
0!
0%
b100 *
0-
02
b100 6
#148410000000
1!
1%
1-
12
#148420000000
0!
0%
b101 *
0-
02
b101 6
#148430000000
1!
1%
1-
12
#148440000000
0!
0%
b110 *
0-
02
b110 6
#148450000000
1!
1%
1-
12
#148460000000
0!
0%
b111 *
0-
02
b111 6
#148470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#148480000000
0!
0%
b0 *
0-
02
b0 6
#148490000000
1!
1%
1-
12
#148500000000
0!
0%
b1 *
0-
02
b1 6
#148510000000
1!
1%
1-
12
#148520000000
0!
0%
b10 *
0-
02
b10 6
#148530000000
1!
1%
1-
12
#148540000000
0!
0%
b11 *
0-
02
b11 6
#148550000000
1!
1%
1-
12
15
#148560000000
0!
0%
b100 *
0-
02
b100 6
#148570000000
1!
1%
1-
12
#148580000000
0!
0%
b101 *
0-
02
b101 6
#148590000000
1!
1%
1-
12
#148600000000
0!
0%
b110 *
0-
02
b110 6
#148610000000
1!
1%
1-
12
#148620000000
0!
0%
b111 *
0-
02
b111 6
#148630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#148640000000
0!
0%
b0 *
0-
02
b0 6
#148650000000
1!
1%
1-
12
#148660000000
0!
0%
b1 *
0-
02
b1 6
#148670000000
1!
1%
1-
12
#148680000000
0!
0%
b10 *
0-
02
b10 6
#148690000000
1!
1%
1-
12
#148700000000
0!
0%
b11 *
0-
02
b11 6
#148710000000
1!
1%
1-
12
15
#148720000000
0!
0%
b100 *
0-
02
b100 6
#148730000000
1!
1%
1-
12
#148740000000
0!
0%
b101 *
0-
02
b101 6
#148750000000
1!
1%
1-
12
#148760000000
0!
0%
b110 *
0-
02
b110 6
#148770000000
1!
1%
1-
12
#148780000000
0!
0%
b111 *
0-
02
b111 6
#148790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#148800000000
0!
0%
b0 *
0-
02
b0 6
#148810000000
1!
1%
1-
12
#148820000000
0!
0%
b1 *
0-
02
b1 6
#148830000000
1!
1%
1-
12
#148840000000
0!
0%
b10 *
0-
02
b10 6
#148850000000
1!
1%
1-
12
#148860000000
0!
0%
b11 *
0-
02
b11 6
#148870000000
1!
1%
1-
12
15
#148880000000
0!
0%
b100 *
0-
02
b100 6
#148890000000
1!
1%
1-
12
#148900000000
0!
0%
b101 *
0-
02
b101 6
#148910000000
1!
1%
1-
12
#148920000000
0!
0%
b110 *
0-
02
b110 6
#148930000000
1!
1%
1-
12
#148940000000
0!
0%
b111 *
0-
02
b111 6
#148950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#148960000000
0!
0%
b0 *
0-
02
b0 6
#148970000000
1!
1%
1-
12
#148980000000
0!
0%
b1 *
0-
02
b1 6
#148990000000
1!
1%
1-
12
#149000000000
0!
0%
b10 *
0-
02
b10 6
#149010000000
1!
1%
1-
12
#149020000000
0!
0%
b11 *
0-
02
b11 6
#149030000000
1!
1%
1-
12
15
#149040000000
0!
0%
b100 *
0-
02
b100 6
#149050000000
1!
1%
1-
12
#149060000000
0!
0%
b101 *
0-
02
b101 6
#149070000000
1!
1%
1-
12
#149080000000
0!
0%
b110 *
0-
02
b110 6
#149090000000
1!
1%
1-
12
#149100000000
0!
0%
b111 *
0-
02
b111 6
#149110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#149120000000
0!
0%
b0 *
0-
02
b0 6
#149130000000
1!
1%
1-
12
#149140000000
0!
0%
b1 *
0-
02
b1 6
#149150000000
1!
1%
1-
12
#149160000000
0!
0%
b10 *
0-
02
b10 6
#149170000000
1!
1%
1-
12
#149180000000
0!
0%
b11 *
0-
02
b11 6
#149190000000
1!
1%
1-
12
15
#149200000000
0!
0%
b100 *
0-
02
b100 6
#149210000000
1!
1%
1-
12
#149220000000
0!
0%
b101 *
0-
02
b101 6
#149230000000
1!
1%
1-
12
#149240000000
0!
0%
b110 *
0-
02
b110 6
#149250000000
1!
1%
1-
12
#149260000000
0!
0%
b111 *
0-
02
b111 6
#149270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#149280000000
0!
0%
b0 *
0-
02
b0 6
#149290000000
1!
1%
1-
12
#149300000000
0!
0%
b1 *
0-
02
b1 6
#149310000000
1!
1%
1-
12
#149320000000
0!
0%
b10 *
0-
02
b10 6
#149330000000
1!
1%
1-
12
#149340000000
0!
0%
b11 *
0-
02
b11 6
#149350000000
1!
1%
1-
12
15
#149360000000
0!
0%
b100 *
0-
02
b100 6
#149370000000
1!
1%
1-
12
#149380000000
0!
0%
b101 *
0-
02
b101 6
#149390000000
1!
1%
1-
12
#149400000000
0!
0%
b110 *
0-
02
b110 6
#149410000000
1!
1%
1-
12
#149420000000
0!
0%
b111 *
0-
02
b111 6
#149430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#149440000000
0!
0%
b0 *
0-
02
b0 6
#149450000000
1!
1%
1-
12
#149460000000
0!
0%
b1 *
0-
02
b1 6
#149470000000
1!
1%
1-
12
#149480000000
0!
0%
b10 *
0-
02
b10 6
#149490000000
1!
1%
1-
12
#149500000000
0!
0%
b11 *
0-
02
b11 6
#149510000000
1!
1%
1-
12
15
#149520000000
0!
0%
b100 *
0-
02
b100 6
#149530000000
1!
1%
1-
12
#149540000000
0!
0%
b101 *
0-
02
b101 6
#149550000000
1!
1%
1-
12
#149560000000
0!
0%
b110 *
0-
02
b110 6
#149570000000
1!
1%
1-
12
#149580000000
0!
0%
b111 *
0-
02
b111 6
#149590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#149600000000
0!
0%
b0 *
0-
02
b0 6
#149610000000
1!
1%
1-
12
#149620000000
0!
0%
b1 *
0-
02
b1 6
#149630000000
1!
1%
1-
12
#149640000000
0!
0%
b10 *
0-
02
b10 6
#149650000000
1!
1%
1-
12
#149660000000
0!
0%
b11 *
0-
02
b11 6
#149670000000
1!
1%
1-
12
15
#149680000000
0!
0%
b100 *
0-
02
b100 6
#149690000000
1!
1%
1-
12
#149700000000
0!
0%
b101 *
0-
02
b101 6
#149710000000
1!
1%
1-
12
#149720000000
0!
0%
b110 *
0-
02
b110 6
#149730000000
1!
1%
1-
12
#149740000000
0!
0%
b111 *
0-
02
b111 6
#149750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#149760000000
0!
0%
b0 *
0-
02
b0 6
#149770000000
1!
1%
1-
12
#149780000000
0!
0%
b1 *
0-
02
b1 6
#149790000000
1!
1%
1-
12
#149800000000
0!
0%
b10 *
0-
02
b10 6
#149810000000
1!
1%
1-
12
#149820000000
0!
0%
b11 *
0-
02
b11 6
#149830000000
1!
1%
1-
12
15
#149840000000
0!
0%
b100 *
0-
02
b100 6
#149850000000
1!
1%
1-
12
#149860000000
0!
0%
b101 *
0-
02
b101 6
#149870000000
1!
1%
1-
12
#149880000000
0!
0%
b110 *
0-
02
b110 6
#149890000000
1!
1%
1-
12
#149900000000
0!
0%
b111 *
0-
02
b111 6
#149910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#149920000000
0!
0%
b0 *
0-
02
b0 6
#149930000000
1!
1%
1-
12
#149940000000
0!
0%
b1 *
0-
02
b1 6
#149950000000
1!
1%
1-
12
#149960000000
0!
0%
b10 *
0-
02
b10 6
#149970000000
1!
1%
1-
12
#149980000000
0!
0%
b11 *
0-
02
b11 6
#149990000000
1!
1%
1-
12
15
#150000000000
0!
0%
b100 *
0-
02
b100 6
#150010000000
1!
1%
1-
12
#150020000000
0!
0%
b101 *
0-
02
b101 6
#150030000000
1!
1%
1-
12
#150040000000
0!
0%
b110 *
0-
02
b110 6
#150050000000
1!
1%
1-
12
#150060000000
0!
0%
b111 *
0-
02
b111 6
#150070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#150080000000
0!
0%
b0 *
0-
02
b0 6
#150090000000
1!
1%
1-
12
#150100000000
0!
0%
b1 *
0-
02
b1 6
#150110000000
1!
1%
1-
12
#150120000000
0!
0%
b10 *
0-
02
b10 6
#150130000000
1!
1%
1-
12
#150140000000
0!
0%
b11 *
0-
02
b11 6
#150150000000
1!
1%
1-
12
15
#150160000000
0!
0%
b100 *
0-
02
b100 6
#150170000000
1!
1%
1-
12
#150180000000
0!
0%
b101 *
0-
02
b101 6
#150190000000
1!
1%
1-
12
#150200000000
0!
0%
b110 *
0-
02
b110 6
#150210000000
1!
1%
1-
12
#150220000000
0!
0%
b111 *
0-
02
b111 6
#150230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#150240000000
0!
0%
b0 *
0-
02
b0 6
#150250000000
1!
1%
1-
12
#150260000000
0!
0%
b1 *
0-
02
b1 6
#150270000000
1!
1%
1-
12
#150280000000
0!
0%
b10 *
0-
02
b10 6
#150290000000
1!
1%
1-
12
#150300000000
0!
0%
b11 *
0-
02
b11 6
#150310000000
1!
1%
1-
12
15
#150320000000
0!
0%
b100 *
0-
02
b100 6
#150330000000
1!
1%
1-
12
#150340000000
0!
0%
b101 *
0-
02
b101 6
#150350000000
1!
1%
1-
12
#150360000000
0!
0%
b110 *
0-
02
b110 6
#150370000000
1!
1%
1-
12
#150380000000
0!
0%
b111 *
0-
02
b111 6
#150390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#150400000000
0!
0%
b0 *
0-
02
b0 6
#150410000000
1!
1%
1-
12
#150420000000
0!
0%
b1 *
0-
02
b1 6
#150430000000
1!
1%
1-
12
#150440000000
0!
0%
b10 *
0-
02
b10 6
#150450000000
1!
1%
1-
12
#150460000000
0!
0%
b11 *
0-
02
b11 6
#150470000000
1!
1%
1-
12
15
#150480000000
0!
0%
b100 *
0-
02
b100 6
#150490000000
1!
1%
1-
12
#150500000000
0!
0%
b101 *
0-
02
b101 6
#150510000000
1!
1%
1-
12
#150520000000
0!
0%
b110 *
0-
02
b110 6
#150530000000
1!
1%
1-
12
#150540000000
0!
0%
b111 *
0-
02
b111 6
#150550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#150560000000
0!
0%
b0 *
0-
02
b0 6
#150570000000
1!
1%
1-
12
#150580000000
0!
0%
b1 *
0-
02
b1 6
#150590000000
1!
1%
1-
12
#150600000000
0!
0%
b10 *
0-
02
b10 6
#150610000000
1!
1%
1-
12
#150620000000
0!
0%
b11 *
0-
02
b11 6
#150630000000
1!
1%
1-
12
15
#150640000000
0!
0%
b100 *
0-
02
b100 6
#150650000000
1!
1%
1-
12
#150660000000
0!
0%
b101 *
0-
02
b101 6
#150670000000
1!
1%
1-
12
#150680000000
0!
0%
b110 *
0-
02
b110 6
#150690000000
1!
1%
1-
12
#150700000000
0!
0%
b111 *
0-
02
b111 6
#150710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#150720000000
0!
0%
b0 *
0-
02
b0 6
#150730000000
1!
1%
1-
12
#150740000000
0!
0%
b1 *
0-
02
b1 6
#150750000000
1!
1%
1-
12
#150760000000
0!
0%
b10 *
0-
02
b10 6
#150770000000
1!
1%
1-
12
#150780000000
0!
0%
b11 *
0-
02
b11 6
#150790000000
1!
1%
1-
12
15
#150800000000
0!
0%
b100 *
0-
02
b100 6
#150810000000
1!
1%
1-
12
#150820000000
0!
0%
b101 *
0-
02
b101 6
#150830000000
1!
1%
1-
12
#150840000000
0!
0%
b110 *
0-
02
b110 6
#150850000000
1!
1%
1-
12
#150860000000
0!
0%
b111 *
0-
02
b111 6
#150870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#150880000000
0!
0%
b0 *
0-
02
b0 6
#150890000000
1!
1%
1-
12
#150900000000
0!
0%
b1 *
0-
02
b1 6
#150910000000
1!
1%
1-
12
#150920000000
0!
0%
b10 *
0-
02
b10 6
#150930000000
1!
1%
1-
12
#150940000000
0!
0%
b11 *
0-
02
b11 6
#150950000000
1!
1%
1-
12
15
#150960000000
0!
0%
b100 *
0-
02
b100 6
#150970000000
1!
1%
1-
12
#150980000000
0!
0%
b101 *
0-
02
b101 6
#150990000000
1!
1%
1-
12
#151000000000
0!
0%
b110 *
0-
02
b110 6
#151010000000
1!
1%
1-
12
#151020000000
0!
0%
b111 *
0-
02
b111 6
#151030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#151040000000
0!
0%
b0 *
0-
02
b0 6
#151050000000
1!
1%
1-
12
#151060000000
0!
0%
b1 *
0-
02
b1 6
#151070000000
1!
1%
1-
12
#151080000000
0!
0%
b10 *
0-
02
b10 6
#151090000000
1!
1%
1-
12
#151100000000
0!
0%
b11 *
0-
02
b11 6
#151110000000
1!
1%
1-
12
15
#151120000000
0!
0%
b100 *
0-
02
b100 6
#151130000000
1!
1%
1-
12
#151140000000
0!
0%
b101 *
0-
02
b101 6
#151150000000
1!
1%
1-
12
#151160000000
0!
0%
b110 *
0-
02
b110 6
#151170000000
1!
1%
1-
12
#151180000000
0!
0%
b111 *
0-
02
b111 6
#151190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#151200000000
0!
0%
b0 *
0-
02
b0 6
#151210000000
1!
1%
1-
12
#151220000000
0!
0%
b1 *
0-
02
b1 6
#151230000000
1!
1%
1-
12
#151240000000
0!
0%
b10 *
0-
02
b10 6
#151250000000
1!
1%
1-
12
#151260000000
0!
0%
b11 *
0-
02
b11 6
#151270000000
1!
1%
1-
12
15
#151280000000
0!
0%
b100 *
0-
02
b100 6
#151290000000
1!
1%
1-
12
#151300000000
0!
0%
b101 *
0-
02
b101 6
#151310000000
1!
1%
1-
12
#151320000000
0!
0%
b110 *
0-
02
b110 6
#151330000000
1!
1%
1-
12
#151340000000
0!
0%
b111 *
0-
02
b111 6
#151350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#151360000000
0!
0%
b0 *
0-
02
b0 6
#151370000000
1!
1%
1-
12
#151380000000
0!
0%
b1 *
0-
02
b1 6
#151390000000
1!
1%
1-
12
#151400000000
0!
0%
b10 *
0-
02
b10 6
#151410000000
1!
1%
1-
12
#151420000000
0!
0%
b11 *
0-
02
b11 6
#151430000000
1!
1%
1-
12
15
#151440000000
0!
0%
b100 *
0-
02
b100 6
#151450000000
1!
1%
1-
12
#151460000000
0!
0%
b101 *
0-
02
b101 6
#151470000000
1!
1%
1-
12
#151480000000
0!
0%
b110 *
0-
02
b110 6
#151490000000
1!
1%
1-
12
#151500000000
0!
0%
b111 *
0-
02
b111 6
#151510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#151520000000
0!
0%
b0 *
0-
02
b0 6
#151530000000
1!
1%
1-
12
#151540000000
0!
0%
b1 *
0-
02
b1 6
#151550000000
1!
1%
1-
12
#151560000000
0!
0%
b10 *
0-
02
b10 6
#151570000000
1!
1%
1-
12
#151580000000
0!
0%
b11 *
0-
02
b11 6
#151590000000
1!
1%
1-
12
15
#151600000000
0!
0%
b100 *
0-
02
b100 6
#151610000000
1!
1%
1-
12
#151620000000
0!
0%
b101 *
0-
02
b101 6
#151630000000
1!
1%
1-
12
#151640000000
0!
0%
b110 *
0-
02
b110 6
#151650000000
1!
1%
1-
12
#151660000000
0!
0%
b111 *
0-
02
b111 6
#151670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#151680000000
0!
0%
b0 *
0-
02
b0 6
#151690000000
1!
1%
1-
12
#151700000000
0!
0%
b1 *
0-
02
b1 6
#151710000000
1!
1%
1-
12
#151720000000
0!
0%
b10 *
0-
02
b10 6
#151730000000
1!
1%
1-
12
#151740000000
0!
0%
b11 *
0-
02
b11 6
#151750000000
1!
1%
1-
12
15
#151760000000
0!
0%
b100 *
0-
02
b100 6
#151770000000
1!
1%
1-
12
#151780000000
0!
0%
b101 *
0-
02
b101 6
#151790000000
1!
1%
1-
12
#151800000000
0!
0%
b110 *
0-
02
b110 6
#151810000000
1!
1%
1-
12
#151820000000
0!
0%
b111 *
0-
02
b111 6
#151830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#151840000000
0!
0%
b0 *
0-
02
b0 6
#151850000000
1!
1%
1-
12
#151860000000
0!
0%
b1 *
0-
02
b1 6
#151870000000
1!
1%
1-
12
#151880000000
0!
0%
b10 *
0-
02
b10 6
#151890000000
1!
1%
1-
12
#151900000000
0!
0%
b11 *
0-
02
b11 6
#151910000000
1!
1%
1-
12
15
#151920000000
0!
0%
b100 *
0-
02
b100 6
#151930000000
1!
1%
1-
12
#151940000000
0!
0%
b101 *
0-
02
b101 6
#151950000000
1!
1%
1-
12
#151960000000
0!
0%
b110 *
0-
02
b110 6
#151970000000
1!
1%
1-
12
#151980000000
0!
0%
b111 *
0-
02
b111 6
#151990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#152000000000
0!
0%
b0 *
0-
02
b0 6
#152010000000
1!
1%
1-
12
#152020000000
0!
0%
b1 *
0-
02
b1 6
#152030000000
1!
1%
1-
12
#152040000000
0!
0%
b10 *
0-
02
b10 6
#152050000000
1!
1%
1-
12
#152060000000
0!
0%
b11 *
0-
02
b11 6
#152070000000
1!
1%
1-
12
15
#152080000000
0!
0%
b100 *
0-
02
b100 6
#152090000000
1!
1%
1-
12
#152100000000
0!
0%
b101 *
0-
02
b101 6
#152110000000
1!
1%
1-
12
#152120000000
0!
0%
b110 *
0-
02
b110 6
#152130000000
1!
1%
1-
12
#152140000000
0!
0%
b111 *
0-
02
b111 6
#152150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#152160000000
0!
0%
b0 *
0-
02
b0 6
#152170000000
1!
1%
1-
12
#152180000000
0!
0%
b1 *
0-
02
b1 6
#152190000000
1!
1%
1-
12
#152200000000
0!
0%
b10 *
0-
02
b10 6
#152210000000
1!
1%
1-
12
#152220000000
0!
0%
b11 *
0-
02
b11 6
#152230000000
1!
1%
1-
12
15
#152240000000
0!
0%
b100 *
0-
02
b100 6
#152250000000
1!
1%
1-
12
#152260000000
0!
0%
b101 *
0-
02
b101 6
#152270000000
1!
1%
1-
12
#152280000000
0!
0%
b110 *
0-
02
b110 6
#152290000000
1!
1%
1-
12
#152300000000
0!
0%
b111 *
0-
02
b111 6
#152310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#152320000000
0!
0%
b0 *
0-
02
b0 6
#152330000000
1!
1%
1-
12
#152340000000
0!
0%
b1 *
0-
02
b1 6
#152350000000
1!
1%
1-
12
#152360000000
0!
0%
b10 *
0-
02
b10 6
#152370000000
1!
1%
1-
12
#152380000000
0!
0%
b11 *
0-
02
b11 6
#152390000000
1!
1%
1-
12
15
#152400000000
0!
0%
b100 *
0-
02
b100 6
#152410000000
1!
1%
1-
12
#152420000000
0!
0%
b101 *
0-
02
b101 6
#152430000000
1!
1%
1-
12
#152440000000
0!
0%
b110 *
0-
02
b110 6
#152450000000
1!
1%
1-
12
#152460000000
0!
0%
b111 *
0-
02
b111 6
#152470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#152480000000
0!
0%
b0 *
0-
02
b0 6
#152490000000
1!
1%
1-
12
#152500000000
0!
0%
b1 *
0-
02
b1 6
#152510000000
1!
1%
1-
12
#152520000000
0!
0%
b10 *
0-
02
b10 6
#152530000000
1!
1%
1-
12
#152540000000
0!
0%
b11 *
0-
02
b11 6
#152550000000
1!
1%
1-
12
15
#152560000000
0!
0%
b100 *
0-
02
b100 6
#152570000000
1!
1%
1-
12
#152580000000
0!
0%
b101 *
0-
02
b101 6
#152590000000
1!
1%
1-
12
#152600000000
0!
0%
b110 *
0-
02
b110 6
#152610000000
1!
1%
1-
12
#152620000000
0!
0%
b111 *
0-
02
b111 6
#152630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#152640000000
0!
0%
b0 *
0-
02
b0 6
#152650000000
1!
1%
1-
12
#152660000000
0!
0%
b1 *
0-
02
b1 6
#152670000000
1!
1%
1-
12
#152680000000
0!
0%
b10 *
0-
02
b10 6
#152690000000
1!
1%
1-
12
#152700000000
0!
0%
b11 *
0-
02
b11 6
#152710000000
1!
1%
1-
12
15
#152720000000
0!
0%
b100 *
0-
02
b100 6
#152730000000
1!
1%
1-
12
#152740000000
0!
0%
b101 *
0-
02
b101 6
#152750000000
1!
1%
1-
12
#152760000000
0!
0%
b110 *
0-
02
b110 6
#152770000000
1!
1%
1-
12
#152780000000
0!
0%
b111 *
0-
02
b111 6
#152790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#152800000000
0!
0%
b0 *
0-
02
b0 6
#152810000000
1!
1%
1-
12
#152820000000
0!
0%
b1 *
0-
02
b1 6
#152830000000
1!
1%
1-
12
#152840000000
0!
0%
b10 *
0-
02
b10 6
#152850000000
1!
1%
1-
12
#152860000000
0!
0%
b11 *
0-
02
b11 6
#152870000000
1!
1%
1-
12
15
#152880000000
0!
0%
b100 *
0-
02
b100 6
#152890000000
1!
1%
1-
12
#152900000000
0!
0%
b101 *
0-
02
b101 6
#152910000000
1!
1%
1-
12
#152920000000
0!
0%
b110 *
0-
02
b110 6
#152930000000
1!
1%
1-
12
#152940000000
0!
0%
b111 *
0-
02
b111 6
#152950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#152960000000
0!
0%
b0 *
0-
02
b0 6
#152970000000
1!
1%
1-
12
#152980000000
0!
0%
b1 *
0-
02
b1 6
#152990000000
1!
1%
1-
12
#153000000000
0!
0%
b10 *
0-
02
b10 6
#153010000000
1!
1%
1-
12
#153020000000
0!
0%
b11 *
0-
02
b11 6
#153030000000
1!
1%
1-
12
15
#153040000000
0!
0%
b100 *
0-
02
b100 6
#153050000000
1!
1%
1-
12
#153060000000
0!
0%
b101 *
0-
02
b101 6
#153070000000
1!
1%
1-
12
#153080000000
0!
0%
b110 *
0-
02
b110 6
#153090000000
1!
1%
1-
12
#153100000000
0!
0%
b111 *
0-
02
b111 6
#153110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#153120000000
0!
0%
b0 *
0-
02
b0 6
#153130000000
1!
1%
1-
12
#153140000000
0!
0%
b1 *
0-
02
b1 6
#153150000000
1!
1%
1-
12
#153160000000
0!
0%
b10 *
0-
02
b10 6
#153170000000
1!
1%
1-
12
#153180000000
0!
0%
b11 *
0-
02
b11 6
#153190000000
1!
1%
1-
12
15
#153200000000
0!
0%
b100 *
0-
02
b100 6
#153210000000
1!
1%
1-
12
#153220000000
0!
0%
b101 *
0-
02
b101 6
#153230000000
1!
1%
1-
12
#153240000000
0!
0%
b110 *
0-
02
b110 6
#153250000000
1!
1%
1-
12
#153260000000
0!
0%
b111 *
0-
02
b111 6
#153270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#153280000000
0!
0%
b0 *
0-
02
b0 6
#153290000000
1!
1%
1-
12
#153300000000
0!
0%
b1 *
0-
02
b1 6
#153310000000
1!
1%
1-
12
#153320000000
0!
0%
b10 *
0-
02
b10 6
#153330000000
1!
1%
1-
12
#153340000000
0!
0%
b11 *
0-
02
b11 6
#153350000000
1!
1%
1-
12
15
#153360000000
0!
0%
b100 *
0-
02
b100 6
#153370000000
1!
1%
1-
12
#153380000000
0!
0%
b101 *
0-
02
b101 6
#153390000000
1!
1%
1-
12
#153400000000
0!
0%
b110 *
0-
02
b110 6
#153410000000
1!
1%
1-
12
#153420000000
0!
0%
b111 *
0-
02
b111 6
#153430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#153440000000
0!
0%
b0 *
0-
02
b0 6
#153450000000
1!
1%
1-
12
#153460000000
0!
0%
b1 *
0-
02
b1 6
#153470000000
1!
1%
1-
12
#153480000000
0!
0%
b10 *
0-
02
b10 6
#153490000000
1!
1%
1-
12
#153500000000
0!
0%
b11 *
0-
02
b11 6
#153510000000
1!
1%
1-
12
15
#153520000000
0!
0%
b100 *
0-
02
b100 6
#153530000000
1!
1%
1-
12
#153540000000
0!
0%
b101 *
0-
02
b101 6
#153550000000
1!
1%
1-
12
#153560000000
0!
0%
b110 *
0-
02
b110 6
#153570000000
1!
1%
1-
12
#153580000000
0!
0%
b111 *
0-
02
b111 6
#153590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#153600000000
0!
0%
b0 *
0-
02
b0 6
#153610000000
1!
1%
1-
12
#153620000000
0!
0%
b1 *
0-
02
b1 6
#153630000000
1!
1%
1-
12
#153640000000
0!
0%
b10 *
0-
02
b10 6
#153650000000
1!
1%
1-
12
#153660000000
0!
0%
b11 *
0-
02
b11 6
#153670000000
1!
1%
1-
12
15
#153680000000
0!
0%
b100 *
0-
02
b100 6
#153690000000
1!
1%
1-
12
#153700000000
0!
0%
b101 *
0-
02
b101 6
#153710000000
1!
1%
1-
12
#153720000000
0!
0%
b110 *
0-
02
b110 6
#153730000000
1!
1%
1-
12
#153740000000
0!
0%
b111 *
0-
02
b111 6
#153750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#153760000000
0!
0%
b0 *
0-
02
b0 6
#153770000000
1!
1%
1-
12
#153780000000
0!
0%
b1 *
0-
02
b1 6
#153790000000
1!
1%
1-
12
#153800000000
0!
0%
b10 *
0-
02
b10 6
#153810000000
1!
1%
1-
12
#153820000000
0!
0%
b11 *
0-
02
b11 6
#153830000000
1!
1%
1-
12
15
#153840000000
0!
0%
b100 *
0-
02
b100 6
#153850000000
1!
1%
1-
12
#153860000000
0!
0%
b101 *
0-
02
b101 6
#153870000000
1!
1%
1-
12
#153880000000
0!
0%
b110 *
0-
02
b110 6
#153890000000
1!
1%
1-
12
#153900000000
0!
0%
b111 *
0-
02
b111 6
#153910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#153920000000
0!
0%
b0 *
0-
02
b0 6
#153930000000
1!
1%
1-
12
#153940000000
0!
0%
b1 *
0-
02
b1 6
#153950000000
1!
1%
1-
12
#153960000000
0!
0%
b10 *
0-
02
b10 6
#153970000000
1!
1%
1-
12
#153980000000
0!
0%
b11 *
0-
02
b11 6
#153990000000
1!
1%
1-
12
15
#154000000000
0!
0%
b100 *
0-
02
b100 6
#154010000000
1!
1%
1-
12
#154020000000
0!
0%
b101 *
0-
02
b101 6
#154030000000
1!
1%
1-
12
#154040000000
0!
0%
b110 *
0-
02
b110 6
#154050000000
1!
1%
1-
12
#154060000000
0!
0%
b111 *
0-
02
b111 6
#154070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#154080000000
0!
0%
b0 *
0-
02
b0 6
#154090000000
1!
1%
1-
12
#154100000000
0!
0%
b1 *
0-
02
b1 6
#154110000000
1!
1%
1-
12
#154120000000
0!
0%
b10 *
0-
02
b10 6
#154130000000
1!
1%
1-
12
#154140000000
0!
0%
b11 *
0-
02
b11 6
#154150000000
1!
1%
1-
12
15
#154160000000
0!
0%
b100 *
0-
02
b100 6
#154170000000
1!
1%
1-
12
#154180000000
0!
0%
b101 *
0-
02
b101 6
#154190000000
1!
1%
1-
12
#154200000000
0!
0%
b110 *
0-
02
b110 6
#154210000000
1!
1%
1-
12
#154220000000
0!
0%
b111 *
0-
02
b111 6
#154230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#154240000000
0!
0%
b0 *
0-
02
b0 6
#154250000000
1!
1%
1-
12
#154260000000
0!
0%
b1 *
0-
02
b1 6
#154270000000
1!
1%
1-
12
#154280000000
0!
0%
b10 *
0-
02
b10 6
#154290000000
1!
1%
1-
12
#154300000000
0!
0%
b11 *
0-
02
b11 6
#154310000000
1!
1%
1-
12
15
#154320000000
0!
0%
b100 *
0-
02
b100 6
#154330000000
1!
1%
1-
12
#154340000000
0!
0%
b101 *
0-
02
b101 6
#154350000000
1!
1%
1-
12
#154360000000
0!
0%
b110 *
0-
02
b110 6
#154370000000
1!
1%
1-
12
#154380000000
0!
0%
b111 *
0-
02
b111 6
#154390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#154400000000
0!
0%
b0 *
0-
02
b0 6
#154410000000
1!
1%
1-
12
#154420000000
0!
0%
b1 *
0-
02
b1 6
#154430000000
1!
1%
1-
12
#154440000000
0!
0%
b10 *
0-
02
b10 6
#154450000000
1!
1%
1-
12
#154460000000
0!
0%
b11 *
0-
02
b11 6
#154470000000
1!
1%
1-
12
15
#154480000000
0!
0%
b100 *
0-
02
b100 6
#154490000000
1!
1%
1-
12
#154500000000
0!
0%
b101 *
0-
02
b101 6
#154510000000
1!
1%
1-
12
#154520000000
0!
0%
b110 *
0-
02
b110 6
#154530000000
1!
1%
1-
12
#154540000000
0!
0%
b111 *
0-
02
b111 6
#154550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#154560000000
0!
0%
b0 *
0-
02
b0 6
#154570000000
1!
1%
1-
12
#154580000000
0!
0%
b1 *
0-
02
b1 6
#154590000000
1!
1%
1-
12
#154600000000
0!
0%
b10 *
0-
02
b10 6
#154610000000
1!
1%
1-
12
#154620000000
0!
0%
b11 *
0-
02
b11 6
#154630000000
1!
1%
1-
12
15
#154640000000
0!
0%
b100 *
0-
02
b100 6
#154650000000
1!
1%
1-
12
#154660000000
0!
0%
b101 *
0-
02
b101 6
#154670000000
1!
1%
1-
12
#154680000000
0!
0%
b110 *
0-
02
b110 6
#154690000000
1!
1%
1-
12
#154700000000
0!
0%
b111 *
0-
02
b111 6
#154710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#154720000000
0!
0%
b0 *
0-
02
b0 6
#154730000000
1!
1%
1-
12
#154740000000
0!
0%
b1 *
0-
02
b1 6
#154750000000
1!
1%
1-
12
#154760000000
0!
0%
b10 *
0-
02
b10 6
#154770000000
1!
1%
1-
12
#154780000000
0!
0%
b11 *
0-
02
b11 6
#154790000000
1!
1%
1-
12
15
#154800000000
0!
0%
b100 *
0-
02
b100 6
#154810000000
1!
1%
1-
12
#154820000000
0!
0%
b101 *
0-
02
b101 6
#154830000000
1!
1%
1-
12
#154840000000
0!
0%
b110 *
0-
02
b110 6
#154850000000
1!
1%
1-
12
#154860000000
0!
0%
b111 *
0-
02
b111 6
#154870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#154880000000
0!
0%
b0 *
0-
02
b0 6
#154890000000
1!
1%
1-
12
#154900000000
0!
0%
b1 *
0-
02
b1 6
#154910000000
1!
1%
1-
12
#154920000000
0!
0%
b10 *
0-
02
b10 6
#154930000000
1!
1%
1-
12
#154940000000
0!
0%
b11 *
0-
02
b11 6
#154950000000
1!
1%
1-
12
15
#154960000000
0!
0%
b100 *
0-
02
b100 6
#154970000000
1!
1%
1-
12
#154980000000
0!
0%
b101 *
0-
02
b101 6
#154990000000
1!
1%
1-
12
#155000000000
0!
0%
b110 *
0-
02
b110 6
#155010000000
1!
1%
1-
12
#155020000000
0!
0%
b111 *
0-
02
b111 6
#155030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#155040000000
0!
0%
b0 *
0-
02
b0 6
#155050000000
1!
1%
1-
12
#155060000000
0!
0%
b1 *
0-
02
b1 6
#155070000000
1!
1%
1-
12
#155080000000
0!
0%
b10 *
0-
02
b10 6
#155090000000
1!
1%
1-
12
#155100000000
0!
0%
b11 *
0-
02
b11 6
#155110000000
1!
1%
1-
12
15
#155120000000
0!
0%
b100 *
0-
02
b100 6
#155130000000
1!
1%
1-
12
#155140000000
0!
0%
b101 *
0-
02
b101 6
#155150000000
1!
1%
1-
12
#155160000000
0!
0%
b110 *
0-
02
b110 6
#155170000000
1!
1%
1-
12
#155180000000
0!
0%
b111 *
0-
02
b111 6
#155190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#155200000000
0!
0%
b0 *
0-
02
b0 6
#155210000000
1!
1%
1-
12
#155220000000
0!
0%
b1 *
0-
02
b1 6
#155230000000
1!
1%
1-
12
#155240000000
0!
0%
b10 *
0-
02
b10 6
#155250000000
1!
1%
1-
12
#155260000000
0!
0%
b11 *
0-
02
b11 6
#155270000000
1!
1%
1-
12
15
#155280000000
0!
0%
b100 *
0-
02
b100 6
#155290000000
1!
1%
1-
12
#155300000000
0!
0%
b101 *
0-
02
b101 6
#155310000000
1!
1%
1-
12
#155320000000
0!
0%
b110 *
0-
02
b110 6
#155330000000
1!
1%
1-
12
#155340000000
0!
0%
b111 *
0-
02
b111 6
#155350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#155360000000
0!
0%
b0 *
0-
02
b0 6
#155370000000
1!
1%
1-
12
#155380000000
0!
0%
b1 *
0-
02
b1 6
#155390000000
1!
1%
1-
12
#155400000000
0!
0%
b10 *
0-
02
b10 6
#155410000000
1!
1%
1-
12
#155420000000
0!
0%
b11 *
0-
02
b11 6
#155430000000
1!
1%
1-
12
15
#155440000000
0!
0%
b100 *
0-
02
b100 6
#155450000000
1!
1%
1-
12
#155460000000
0!
0%
b101 *
0-
02
b101 6
#155470000000
1!
1%
1-
12
#155480000000
0!
0%
b110 *
0-
02
b110 6
#155490000000
1!
1%
1-
12
#155500000000
0!
0%
b111 *
0-
02
b111 6
#155510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#155520000000
0!
0%
b0 *
0-
02
b0 6
#155530000000
1!
1%
1-
12
#155540000000
0!
0%
b1 *
0-
02
b1 6
#155550000000
1!
1%
1-
12
#155560000000
0!
0%
b10 *
0-
02
b10 6
#155570000000
1!
1%
1-
12
#155580000000
0!
0%
b11 *
0-
02
b11 6
#155590000000
1!
1%
1-
12
15
#155600000000
0!
0%
b100 *
0-
02
b100 6
#155610000000
1!
1%
1-
12
#155620000000
0!
0%
b101 *
0-
02
b101 6
#155630000000
1!
1%
1-
12
#155640000000
0!
0%
b110 *
0-
02
b110 6
#155650000000
1!
1%
1-
12
#155660000000
0!
0%
b111 *
0-
02
b111 6
#155670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#155680000000
0!
0%
b0 *
0-
02
b0 6
#155690000000
1!
1%
1-
12
#155700000000
0!
0%
b1 *
0-
02
b1 6
#155710000000
1!
1%
1-
12
#155720000000
0!
0%
b10 *
0-
02
b10 6
#155730000000
1!
1%
1-
12
#155740000000
0!
0%
b11 *
0-
02
b11 6
#155750000000
1!
1%
1-
12
15
#155760000000
0!
0%
b100 *
0-
02
b100 6
#155770000000
1!
1%
1-
12
#155780000000
0!
0%
b101 *
0-
02
b101 6
#155790000000
1!
1%
1-
12
#155800000000
0!
0%
b110 *
0-
02
b110 6
#155810000000
1!
1%
1-
12
#155820000000
0!
0%
b111 *
0-
02
b111 6
#155830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#155840000000
0!
0%
b0 *
0-
02
b0 6
#155850000000
1!
1%
1-
12
#155860000000
0!
0%
b1 *
0-
02
b1 6
#155870000000
1!
1%
1-
12
#155880000000
0!
0%
b10 *
0-
02
b10 6
#155890000000
1!
1%
1-
12
#155900000000
0!
0%
b11 *
0-
02
b11 6
#155910000000
1!
1%
1-
12
15
#155920000000
0!
0%
b100 *
0-
02
b100 6
#155930000000
1!
1%
1-
12
#155940000000
0!
0%
b101 *
0-
02
b101 6
#155950000000
1!
1%
1-
12
#155960000000
0!
0%
b110 *
0-
02
b110 6
#155970000000
1!
1%
1-
12
#155980000000
0!
0%
b111 *
0-
02
b111 6
#155990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#156000000000
0!
0%
b0 *
0-
02
b0 6
#156010000000
1!
1%
1-
12
#156020000000
0!
0%
b1 *
0-
02
b1 6
#156030000000
1!
1%
1-
12
#156040000000
0!
0%
b10 *
0-
02
b10 6
#156050000000
1!
1%
1-
12
#156060000000
0!
0%
b11 *
0-
02
b11 6
#156070000000
1!
1%
1-
12
15
#156080000000
0!
0%
b100 *
0-
02
b100 6
#156090000000
1!
1%
1-
12
#156100000000
0!
0%
b101 *
0-
02
b101 6
#156110000000
1!
1%
1-
12
#156120000000
0!
0%
b110 *
0-
02
b110 6
#156130000000
1!
1%
1-
12
#156140000000
0!
0%
b111 *
0-
02
b111 6
#156150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#156160000000
0!
0%
b0 *
0-
02
b0 6
#156170000000
1!
1%
1-
12
#156180000000
0!
0%
b1 *
0-
02
b1 6
#156190000000
1!
1%
1-
12
#156200000000
0!
0%
b10 *
0-
02
b10 6
#156210000000
1!
1%
1-
12
#156220000000
0!
0%
b11 *
0-
02
b11 6
#156230000000
1!
1%
1-
12
15
#156240000000
0!
0%
b100 *
0-
02
b100 6
#156250000000
1!
1%
1-
12
#156260000000
0!
0%
b101 *
0-
02
b101 6
#156270000000
1!
1%
1-
12
#156280000000
0!
0%
b110 *
0-
02
b110 6
#156290000000
1!
1%
1-
12
#156300000000
0!
0%
b111 *
0-
02
b111 6
#156310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#156320000000
0!
0%
b0 *
0-
02
b0 6
#156330000000
1!
1%
1-
12
#156340000000
0!
0%
b1 *
0-
02
b1 6
#156350000000
1!
1%
1-
12
#156360000000
0!
0%
b10 *
0-
02
b10 6
#156370000000
1!
1%
1-
12
#156380000000
0!
0%
b11 *
0-
02
b11 6
#156390000000
1!
1%
1-
12
15
#156400000000
0!
0%
b100 *
0-
02
b100 6
#156410000000
1!
1%
1-
12
#156420000000
0!
0%
b101 *
0-
02
b101 6
#156430000000
1!
1%
1-
12
#156440000000
0!
0%
b110 *
0-
02
b110 6
#156450000000
1!
1%
1-
12
#156460000000
0!
0%
b111 *
0-
02
b111 6
#156470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#156480000000
0!
0%
b0 *
0-
02
b0 6
#156490000000
1!
1%
1-
12
#156500000000
0!
0%
b1 *
0-
02
b1 6
#156510000000
1!
1%
1-
12
#156520000000
0!
0%
b10 *
0-
02
b10 6
#156530000000
1!
1%
1-
12
#156540000000
0!
0%
b11 *
0-
02
b11 6
#156550000000
1!
1%
1-
12
15
#156560000000
0!
0%
b100 *
0-
02
b100 6
#156570000000
1!
1%
1-
12
#156580000000
0!
0%
b101 *
0-
02
b101 6
#156590000000
1!
1%
1-
12
#156600000000
0!
0%
b110 *
0-
02
b110 6
#156610000000
1!
1%
1-
12
#156620000000
0!
0%
b111 *
0-
02
b111 6
#156630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#156640000000
0!
0%
b0 *
0-
02
b0 6
#156650000000
1!
1%
1-
12
#156660000000
0!
0%
b1 *
0-
02
b1 6
#156670000000
1!
1%
1-
12
#156680000000
0!
0%
b10 *
0-
02
b10 6
#156690000000
1!
1%
1-
12
#156700000000
0!
0%
b11 *
0-
02
b11 6
#156710000000
1!
1%
1-
12
15
#156720000000
0!
0%
b100 *
0-
02
b100 6
#156730000000
1!
1%
1-
12
#156740000000
0!
0%
b101 *
0-
02
b101 6
#156750000000
1!
1%
1-
12
#156760000000
0!
0%
b110 *
0-
02
b110 6
#156770000000
1!
1%
1-
12
#156780000000
0!
0%
b111 *
0-
02
b111 6
#156790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#156800000000
0!
0%
b0 *
0-
02
b0 6
#156810000000
1!
1%
1-
12
#156820000000
0!
0%
b1 *
0-
02
b1 6
#156830000000
1!
1%
1-
12
#156840000000
0!
0%
b10 *
0-
02
b10 6
#156850000000
1!
1%
1-
12
#156860000000
0!
0%
b11 *
0-
02
b11 6
#156870000000
1!
1%
1-
12
15
#156880000000
0!
0%
b100 *
0-
02
b100 6
#156890000000
1!
1%
1-
12
#156900000000
0!
0%
b101 *
0-
02
b101 6
#156910000000
1!
1%
1-
12
#156920000000
0!
0%
b110 *
0-
02
b110 6
#156930000000
1!
1%
1-
12
#156940000000
0!
0%
b111 *
0-
02
b111 6
#156950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#156960000000
0!
0%
b0 *
0-
02
b0 6
#156970000000
1!
1%
1-
12
#156980000000
0!
0%
b1 *
0-
02
b1 6
#156990000000
1!
1%
1-
12
#157000000000
0!
0%
b10 *
0-
02
b10 6
#157010000000
1!
1%
1-
12
#157020000000
0!
0%
b11 *
0-
02
b11 6
#157030000000
1!
1%
1-
12
15
#157040000000
0!
0%
b100 *
0-
02
b100 6
#157050000000
1!
1%
1-
12
#157060000000
0!
0%
b101 *
0-
02
b101 6
#157070000000
1!
1%
1-
12
#157080000000
0!
0%
b110 *
0-
02
b110 6
#157090000000
1!
1%
1-
12
#157100000000
0!
0%
b111 *
0-
02
b111 6
#157110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#157120000000
0!
0%
b0 *
0-
02
b0 6
#157130000000
1!
1%
1-
12
#157140000000
0!
0%
b1 *
0-
02
b1 6
#157150000000
1!
1%
1-
12
#157160000000
0!
0%
b10 *
0-
02
b10 6
#157170000000
1!
1%
1-
12
#157180000000
0!
0%
b11 *
0-
02
b11 6
#157190000000
1!
1%
1-
12
15
#157200000000
0!
0%
b100 *
0-
02
b100 6
#157210000000
1!
1%
1-
12
#157220000000
0!
0%
b101 *
0-
02
b101 6
#157230000000
1!
1%
1-
12
#157240000000
0!
0%
b110 *
0-
02
b110 6
#157250000000
1!
1%
1-
12
#157260000000
0!
0%
b111 *
0-
02
b111 6
#157270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#157280000000
0!
0%
b0 *
0-
02
b0 6
#157290000000
1!
1%
1-
12
#157300000000
0!
0%
b1 *
0-
02
b1 6
#157310000000
1!
1%
1-
12
#157320000000
0!
0%
b10 *
0-
02
b10 6
#157330000000
1!
1%
1-
12
#157340000000
0!
0%
b11 *
0-
02
b11 6
#157350000000
1!
1%
1-
12
15
#157360000000
0!
0%
b100 *
0-
02
b100 6
#157370000000
1!
1%
1-
12
#157380000000
0!
0%
b101 *
0-
02
b101 6
#157390000000
1!
1%
1-
12
#157400000000
0!
0%
b110 *
0-
02
b110 6
#157410000000
1!
1%
1-
12
#157420000000
0!
0%
b111 *
0-
02
b111 6
#157430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#157440000000
0!
0%
b0 *
0-
02
b0 6
#157450000000
1!
1%
1-
12
#157460000000
0!
0%
b1 *
0-
02
b1 6
#157470000000
1!
1%
1-
12
#157480000000
0!
0%
b10 *
0-
02
b10 6
#157490000000
1!
1%
1-
12
#157500000000
0!
0%
b11 *
0-
02
b11 6
#157510000000
1!
1%
1-
12
15
#157520000000
0!
0%
b100 *
0-
02
b100 6
#157530000000
1!
1%
1-
12
#157540000000
0!
0%
b101 *
0-
02
b101 6
#157550000000
1!
1%
1-
12
#157560000000
0!
0%
b110 *
0-
02
b110 6
#157570000000
1!
1%
1-
12
#157580000000
0!
0%
b111 *
0-
02
b111 6
#157590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#157600000000
0!
0%
b0 *
0-
02
b0 6
#157610000000
1!
1%
1-
12
#157620000000
0!
0%
b1 *
0-
02
b1 6
#157630000000
1!
1%
1-
12
#157640000000
0!
0%
b10 *
0-
02
b10 6
#157650000000
1!
1%
1-
12
#157660000000
0!
0%
b11 *
0-
02
b11 6
#157670000000
1!
1%
1-
12
15
#157680000000
0!
0%
b100 *
0-
02
b100 6
#157690000000
1!
1%
1-
12
#157700000000
0!
0%
b101 *
0-
02
b101 6
#157710000000
1!
1%
1-
12
#157720000000
0!
0%
b110 *
0-
02
b110 6
#157730000000
1!
1%
1-
12
#157740000000
0!
0%
b111 *
0-
02
b111 6
#157750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#157760000000
0!
0%
b0 *
0-
02
b0 6
#157770000000
1!
1%
1-
12
#157780000000
0!
0%
b1 *
0-
02
b1 6
#157790000000
1!
1%
1-
12
#157800000000
0!
0%
b10 *
0-
02
b10 6
#157810000000
1!
1%
1-
12
#157820000000
0!
0%
b11 *
0-
02
b11 6
#157830000000
1!
1%
1-
12
15
#157840000000
0!
0%
b100 *
0-
02
b100 6
#157850000000
1!
1%
1-
12
#157860000000
0!
0%
b101 *
0-
02
b101 6
#157870000000
1!
1%
1-
12
#157880000000
0!
0%
b110 *
0-
02
b110 6
#157890000000
1!
1%
1-
12
#157900000000
0!
0%
b111 *
0-
02
b111 6
#157910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#157920000000
0!
0%
b0 *
0-
02
b0 6
#157930000000
1!
1%
1-
12
#157940000000
0!
0%
b1 *
0-
02
b1 6
#157950000000
1!
1%
1-
12
#157960000000
0!
0%
b10 *
0-
02
b10 6
#157970000000
1!
1%
1-
12
#157980000000
0!
0%
b11 *
0-
02
b11 6
#157990000000
1!
1%
1-
12
15
#158000000000
0!
0%
b100 *
0-
02
b100 6
#158010000000
1!
1%
1-
12
#158020000000
0!
0%
b101 *
0-
02
b101 6
#158030000000
1!
1%
1-
12
#158040000000
0!
0%
b110 *
0-
02
b110 6
#158050000000
1!
1%
1-
12
#158060000000
0!
0%
b111 *
0-
02
b111 6
#158070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#158080000000
0!
0%
b0 *
0-
02
b0 6
#158090000000
1!
1%
1-
12
#158100000000
0!
0%
b1 *
0-
02
b1 6
#158110000000
1!
1%
1-
12
#158120000000
0!
0%
b10 *
0-
02
b10 6
#158130000000
1!
1%
1-
12
#158140000000
0!
0%
b11 *
0-
02
b11 6
#158150000000
1!
1%
1-
12
15
#158160000000
0!
0%
b100 *
0-
02
b100 6
#158170000000
1!
1%
1-
12
#158180000000
0!
0%
b101 *
0-
02
b101 6
#158190000000
1!
1%
1-
12
#158200000000
0!
0%
b110 *
0-
02
b110 6
#158210000000
1!
1%
1-
12
#158220000000
0!
0%
b111 *
0-
02
b111 6
#158230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#158240000000
0!
0%
b0 *
0-
02
b0 6
#158250000000
1!
1%
1-
12
#158260000000
0!
0%
b1 *
0-
02
b1 6
#158270000000
1!
1%
1-
12
#158280000000
0!
0%
b10 *
0-
02
b10 6
#158290000000
1!
1%
1-
12
#158300000000
0!
0%
b11 *
0-
02
b11 6
#158310000000
1!
1%
1-
12
15
#158320000000
0!
0%
b100 *
0-
02
b100 6
#158330000000
1!
1%
1-
12
#158340000000
0!
0%
b101 *
0-
02
b101 6
#158350000000
1!
1%
1-
12
#158360000000
0!
0%
b110 *
0-
02
b110 6
#158370000000
1!
1%
1-
12
#158380000000
0!
0%
b111 *
0-
02
b111 6
#158390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#158400000000
0!
0%
b0 *
0-
02
b0 6
#158410000000
1!
1%
1-
12
#158420000000
0!
0%
b1 *
0-
02
b1 6
#158430000000
1!
1%
1-
12
#158440000000
0!
0%
b10 *
0-
02
b10 6
#158450000000
1!
1%
1-
12
#158460000000
0!
0%
b11 *
0-
02
b11 6
#158470000000
1!
1%
1-
12
15
#158480000000
0!
0%
b100 *
0-
02
b100 6
#158490000000
1!
1%
1-
12
#158500000000
0!
0%
b101 *
0-
02
b101 6
#158510000000
1!
1%
1-
12
#158520000000
0!
0%
b110 *
0-
02
b110 6
#158530000000
1!
1%
1-
12
#158540000000
0!
0%
b111 *
0-
02
b111 6
#158550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#158560000000
0!
0%
b0 *
0-
02
b0 6
#158570000000
1!
1%
1-
12
#158580000000
0!
0%
b1 *
0-
02
b1 6
#158590000000
1!
1%
1-
12
#158600000000
0!
0%
b10 *
0-
02
b10 6
#158610000000
1!
1%
1-
12
#158620000000
0!
0%
b11 *
0-
02
b11 6
#158630000000
1!
1%
1-
12
15
#158640000000
0!
0%
b100 *
0-
02
b100 6
#158650000000
1!
1%
1-
12
#158660000000
0!
0%
b101 *
0-
02
b101 6
#158670000000
1!
1%
1-
12
#158680000000
0!
0%
b110 *
0-
02
b110 6
#158690000000
1!
1%
1-
12
#158700000000
0!
0%
b111 *
0-
02
b111 6
#158710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#158720000000
0!
0%
b0 *
0-
02
b0 6
#158730000000
1!
1%
1-
12
#158740000000
0!
0%
b1 *
0-
02
b1 6
#158750000000
1!
1%
1-
12
#158760000000
0!
0%
b10 *
0-
02
b10 6
#158770000000
1!
1%
1-
12
#158780000000
0!
0%
b11 *
0-
02
b11 6
#158790000000
1!
1%
1-
12
15
#158800000000
0!
0%
b100 *
0-
02
b100 6
#158810000000
1!
1%
1-
12
#158820000000
0!
0%
b101 *
0-
02
b101 6
#158830000000
1!
1%
1-
12
#158840000000
0!
0%
b110 *
0-
02
b110 6
#158850000000
1!
1%
1-
12
#158860000000
0!
0%
b111 *
0-
02
b111 6
#158870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#158880000000
0!
0%
b0 *
0-
02
b0 6
#158890000000
1!
1%
1-
12
#158900000000
0!
0%
b1 *
0-
02
b1 6
#158910000000
1!
1%
1-
12
#158920000000
0!
0%
b10 *
0-
02
b10 6
#158930000000
1!
1%
1-
12
#158940000000
0!
0%
b11 *
0-
02
b11 6
#158950000000
1!
1%
1-
12
15
#158960000000
0!
0%
b100 *
0-
02
b100 6
#158970000000
1!
1%
1-
12
#158980000000
0!
0%
b101 *
0-
02
b101 6
#158990000000
1!
1%
1-
12
#159000000000
0!
0%
b110 *
0-
02
b110 6
#159010000000
1!
1%
1-
12
#159020000000
0!
0%
b111 *
0-
02
b111 6
#159030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#159040000000
0!
0%
b0 *
0-
02
b0 6
#159050000000
1!
1%
1-
12
#159060000000
0!
0%
b1 *
0-
02
b1 6
#159070000000
1!
1%
1-
12
#159080000000
0!
0%
b10 *
0-
02
b10 6
#159090000000
1!
1%
1-
12
#159100000000
0!
0%
b11 *
0-
02
b11 6
#159110000000
1!
1%
1-
12
15
#159120000000
0!
0%
b100 *
0-
02
b100 6
#159130000000
1!
1%
1-
12
#159140000000
0!
0%
b101 *
0-
02
b101 6
#159150000000
1!
1%
1-
12
#159160000000
0!
0%
b110 *
0-
02
b110 6
#159170000000
1!
1%
1-
12
#159180000000
0!
0%
b111 *
0-
02
b111 6
#159190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#159200000000
0!
0%
b0 *
0-
02
b0 6
#159210000000
1!
1%
1-
12
#159220000000
0!
0%
b1 *
0-
02
b1 6
#159230000000
1!
1%
1-
12
#159240000000
0!
0%
b10 *
0-
02
b10 6
#159250000000
1!
1%
1-
12
#159260000000
0!
0%
b11 *
0-
02
b11 6
#159270000000
1!
1%
1-
12
15
#159280000000
0!
0%
b100 *
0-
02
b100 6
#159290000000
1!
1%
1-
12
#159300000000
0!
0%
b101 *
0-
02
b101 6
#159310000000
1!
1%
1-
12
#159320000000
0!
0%
b110 *
0-
02
b110 6
#159330000000
1!
1%
1-
12
#159340000000
0!
0%
b111 *
0-
02
b111 6
#159350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#159360000000
0!
0%
b0 *
0-
02
b0 6
#159370000000
1!
1%
1-
12
#159380000000
0!
0%
b1 *
0-
02
b1 6
#159390000000
1!
1%
1-
12
#159400000000
0!
0%
b10 *
0-
02
b10 6
#159410000000
1!
1%
1-
12
#159420000000
0!
0%
b11 *
0-
02
b11 6
#159430000000
1!
1%
1-
12
15
#159440000000
0!
0%
b100 *
0-
02
b100 6
#159450000000
1!
1%
1-
12
#159460000000
0!
0%
b101 *
0-
02
b101 6
#159470000000
1!
1%
1-
12
#159480000000
0!
0%
b110 *
0-
02
b110 6
#159490000000
1!
1%
1-
12
#159500000000
0!
0%
b111 *
0-
02
b111 6
#159510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#159520000000
0!
0%
b0 *
0-
02
b0 6
#159530000000
1!
1%
1-
12
#159540000000
0!
0%
b1 *
0-
02
b1 6
#159550000000
1!
1%
1-
12
#159560000000
0!
0%
b10 *
0-
02
b10 6
#159570000000
1!
1%
1-
12
#159580000000
0!
0%
b11 *
0-
02
b11 6
#159590000000
1!
1%
1-
12
15
#159600000000
0!
0%
b100 *
0-
02
b100 6
#159610000000
1!
1%
1-
12
#159620000000
0!
0%
b101 *
0-
02
b101 6
#159630000000
1!
1%
1-
12
#159640000000
0!
0%
b110 *
0-
02
b110 6
#159650000000
1!
1%
1-
12
#159660000000
0!
0%
b111 *
0-
02
b111 6
#159670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#159680000000
0!
0%
b0 *
0-
02
b0 6
#159690000000
1!
1%
1-
12
#159700000000
0!
0%
b1 *
0-
02
b1 6
#159710000000
1!
1%
1-
12
#159720000000
0!
0%
b10 *
0-
02
b10 6
#159730000000
1!
1%
1-
12
#159740000000
0!
0%
b11 *
0-
02
b11 6
#159750000000
1!
1%
1-
12
15
#159760000000
0!
0%
b100 *
0-
02
b100 6
#159770000000
1!
1%
1-
12
#159780000000
0!
0%
b101 *
0-
02
b101 6
#159790000000
1!
1%
1-
12
#159800000000
0!
0%
b110 *
0-
02
b110 6
#159810000000
1!
1%
1-
12
#159820000000
0!
0%
b111 *
0-
02
b111 6
#159830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#159840000000
0!
0%
b0 *
0-
02
b0 6
#159850000000
1!
1%
1-
12
#159860000000
0!
0%
b1 *
0-
02
b1 6
#159870000000
1!
1%
1-
12
#159880000000
0!
0%
b10 *
0-
02
b10 6
#159890000000
1!
1%
1-
12
#159900000000
0!
0%
b11 *
0-
02
b11 6
#159910000000
1!
1%
1-
12
15
#159920000000
0!
0%
b100 *
0-
02
b100 6
#159930000000
1!
1%
1-
12
#159940000000
0!
0%
b101 *
0-
02
b101 6
#159950000000
1!
1%
1-
12
#159960000000
0!
0%
b110 *
0-
02
b110 6
#159970000000
1!
1%
1-
12
#159980000000
0!
0%
b111 *
0-
02
b111 6
#159990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#160000000000
0!
0%
b0 *
0-
02
b0 6
#160010000000
1!
1%
1-
12
#160020000000
0!
0%
b1 *
0-
02
b1 6
#160030000000
1!
1%
1-
12
#160040000000
0!
0%
b10 *
0-
02
b10 6
#160050000000
1!
1%
1-
12
#160060000000
0!
0%
b11 *
0-
02
b11 6
#160070000000
1!
1%
1-
12
15
#160080000000
0!
0%
b100 *
0-
02
b100 6
#160090000000
1!
1%
1-
12
#160100000000
0!
0%
b101 *
0-
02
b101 6
#160110000000
1!
1%
1-
12
#160120000000
0!
0%
b110 *
0-
02
b110 6
#160130000000
1!
1%
1-
12
#160140000000
0!
0%
b111 *
0-
02
b111 6
#160150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#160160000000
0!
0%
b0 *
0-
02
b0 6
#160170000000
1!
1%
1-
12
#160180000000
0!
0%
b1 *
0-
02
b1 6
#160190000000
1!
1%
1-
12
#160200000000
0!
0%
b10 *
0-
02
b10 6
#160210000000
1!
1%
1-
12
#160220000000
0!
0%
b11 *
0-
02
b11 6
#160230000000
1!
1%
1-
12
15
#160240000000
0!
0%
b100 *
0-
02
b100 6
#160250000000
1!
1%
1-
12
#160260000000
0!
0%
b101 *
0-
02
b101 6
#160270000000
1!
1%
1-
12
#160280000000
0!
0%
b110 *
0-
02
b110 6
#160290000000
1!
1%
1-
12
#160300000000
0!
0%
b111 *
0-
02
b111 6
#160310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#160320000000
0!
0%
b0 *
0-
02
b0 6
#160330000000
1!
1%
1-
12
#160340000000
0!
0%
b1 *
0-
02
b1 6
#160350000000
1!
1%
1-
12
#160360000000
0!
0%
b10 *
0-
02
b10 6
#160370000000
1!
1%
1-
12
#160380000000
0!
0%
b11 *
0-
02
b11 6
#160390000000
1!
1%
1-
12
15
#160400000000
0!
0%
b100 *
0-
02
b100 6
#160410000000
1!
1%
1-
12
#160420000000
0!
0%
b101 *
0-
02
b101 6
#160430000000
1!
1%
1-
12
#160440000000
0!
0%
b110 *
0-
02
b110 6
#160450000000
1!
1%
1-
12
#160460000000
0!
0%
b111 *
0-
02
b111 6
#160470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#160480000000
0!
0%
b0 *
0-
02
b0 6
#160490000000
1!
1%
1-
12
#160500000000
0!
0%
b1 *
0-
02
b1 6
#160510000000
1!
1%
1-
12
#160520000000
0!
0%
b10 *
0-
02
b10 6
#160530000000
1!
1%
1-
12
#160540000000
0!
0%
b11 *
0-
02
b11 6
#160550000000
1!
1%
1-
12
15
#160560000000
0!
0%
b100 *
0-
02
b100 6
#160570000000
1!
1%
1-
12
#160580000000
0!
0%
b101 *
0-
02
b101 6
#160590000000
1!
1%
1-
12
#160600000000
0!
0%
b110 *
0-
02
b110 6
#160610000000
1!
1%
1-
12
#160620000000
0!
0%
b111 *
0-
02
b111 6
#160630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#160640000000
0!
0%
b0 *
0-
02
b0 6
#160650000000
1!
1%
1-
12
#160660000000
0!
0%
b1 *
0-
02
b1 6
#160670000000
1!
1%
1-
12
#160680000000
0!
0%
b10 *
0-
02
b10 6
#160690000000
1!
1%
1-
12
#160700000000
0!
0%
b11 *
0-
02
b11 6
#160710000000
1!
1%
1-
12
15
#160720000000
0!
0%
b100 *
0-
02
b100 6
#160730000000
1!
1%
1-
12
#160740000000
0!
0%
b101 *
0-
02
b101 6
#160750000000
1!
1%
1-
12
#160760000000
0!
0%
b110 *
0-
02
b110 6
#160770000000
1!
1%
1-
12
#160780000000
0!
0%
b111 *
0-
02
b111 6
#160790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#160800000000
0!
0%
b0 *
0-
02
b0 6
#160810000000
1!
1%
1-
12
#160820000000
0!
0%
b1 *
0-
02
b1 6
#160830000000
1!
1%
1-
12
#160840000000
0!
0%
b10 *
0-
02
b10 6
#160850000000
1!
1%
1-
12
#160860000000
0!
0%
b11 *
0-
02
b11 6
#160870000000
1!
1%
1-
12
15
#160880000000
0!
0%
b100 *
0-
02
b100 6
#160890000000
1!
1%
1-
12
#160900000000
0!
0%
b101 *
0-
02
b101 6
#160910000000
1!
1%
1-
12
#160920000000
0!
0%
b110 *
0-
02
b110 6
#160930000000
1!
1%
1-
12
#160940000000
0!
0%
b111 *
0-
02
b111 6
#160950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#160960000000
0!
0%
b0 *
0-
02
b0 6
#160970000000
1!
1%
1-
12
#160980000000
0!
0%
b1 *
0-
02
b1 6
#160990000000
1!
1%
1-
12
#161000000000
0!
0%
b10 *
0-
02
b10 6
#161010000000
1!
1%
1-
12
#161020000000
0!
0%
b11 *
0-
02
b11 6
#161030000000
1!
1%
1-
12
15
#161040000000
0!
0%
b100 *
0-
02
b100 6
#161050000000
1!
1%
1-
12
#161060000000
0!
0%
b101 *
0-
02
b101 6
#161070000000
1!
1%
1-
12
#161080000000
0!
0%
b110 *
0-
02
b110 6
#161090000000
1!
1%
1-
12
#161100000000
0!
0%
b111 *
0-
02
b111 6
#161110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#161120000000
0!
0%
b0 *
0-
02
b0 6
#161130000000
1!
1%
1-
12
#161140000000
0!
0%
b1 *
0-
02
b1 6
#161150000000
1!
1%
1-
12
#161160000000
0!
0%
b10 *
0-
02
b10 6
#161170000000
1!
1%
1-
12
#161180000000
0!
0%
b11 *
0-
02
b11 6
#161190000000
1!
1%
1-
12
15
#161200000000
0!
0%
b100 *
0-
02
b100 6
#161210000000
1!
1%
1-
12
#161220000000
0!
0%
b101 *
0-
02
b101 6
#161230000000
1!
1%
1-
12
#161240000000
0!
0%
b110 *
0-
02
b110 6
#161250000000
1!
1%
1-
12
#161260000000
0!
0%
b111 *
0-
02
b111 6
#161270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#161280000000
0!
0%
b0 *
0-
02
b0 6
#161290000000
1!
1%
1-
12
#161300000000
0!
0%
b1 *
0-
02
b1 6
#161310000000
1!
1%
1-
12
#161320000000
0!
0%
b10 *
0-
02
b10 6
#161330000000
1!
1%
1-
12
#161340000000
0!
0%
b11 *
0-
02
b11 6
#161350000000
1!
1%
1-
12
15
#161360000000
0!
0%
b100 *
0-
02
b100 6
#161370000000
1!
1%
1-
12
#161380000000
0!
0%
b101 *
0-
02
b101 6
#161390000000
1!
1%
1-
12
#161400000000
0!
0%
b110 *
0-
02
b110 6
#161410000000
1!
1%
1-
12
#161420000000
0!
0%
b111 *
0-
02
b111 6
#161430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#161440000000
0!
0%
b0 *
0-
02
b0 6
#161450000000
1!
1%
1-
12
#161460000000
0!
0%
b1 *
0-
02
b1 6
#161470000000
1!
1%
1-
12
#161480000000
0!
0%
b10 *
0-
02
b10 6
#161490000000
1!
1%
1-
12
#161500000000
0!
0%
b11 *
0-
02
b11 6
#161510000000
1!
1%
1-
12
15
#161520000000
0!
0%
b100 *
0-
02
b100 6
#161530000000
1!
1%
1-
12
#161540000000
0!
0%
b101 *
0-
02
b101 6
#161550000000
1!
1%
1-
12
#161560000000
0!
0%
b110 *
0-
02
b110 6
#161570000000
1!
1%
1-
12
#161580000000
0!
0%
b111 *
0-
02
b111 6
#161590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#161600000000
0!
0%
b0 *
0-
02
b0 6
#161610000000
1!
1%
1-
12
#161620000000
0!
0%
b1 *
0-
02
b1 6
#161630000000
1!
1%
1-
12
#161640000000
0!
0%
b10 *
0-
02
b10 6
#161650000000
1!
1%
1-
12
#161660000000
0!
0%
b11 *
0-
02
b11 6
#161670000000
1!
1%
1-
12
15
#161680000000
0!
0%
b100 *
0-
02
b100 6
#161690000000
1!
1%
1-
12
#161700000000
0!
0%
b101 *
0-
02
b101 6
#161710000000
1!
1%
1-
12
#161720000000
0!
0%
b110 *
0-
02
b110 6
#161730000000
1!
1%
1-
12
#161740000000
0!
0%
b111 *
0-
02
b111 6
#161750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#161760000000
0!
0%
b0 *
0-
02
b0 6
#161770000000
1!
1%
1-
12
#161780000000
0!
0%
b1 *
0-
02
b1 6
#161790000000
1!
1%
1-
12
#161800000000
0!
0%
b10 *
0-
02
b10 6
#161810000000
1!
1%
1-
12
#161820000000
0!
0%
b11 *
0-
02
b11 6
#161830000000
1!
1%
1-
12
15
#161840000000
0!
0%
b100 *
0-
02
b100 6
#161850000000
1!
1%
1-
12
#161860000000
0!
0%
b101 *
0-
02
b101 6
#161870000000
1!
1%
1-
12
#161880000000
0!
0%
b110 *
0-
02
b110 6
#161890000000
1!
1%
1-
12
#161900000000
0!
0%
b111 *
0-
02
b111 6
#161910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#161920000000
0!
0%
b0 *
0-
02
b0 6
#161930000000
1!
1%
1-
12
#161940000000
0!
0%
b1 *
0-
02
b1 6
#161950000000
1!
1%
1-
12
#161960000000
0!
0%
b10 *
0-
02
b10 6
#161970000000
1!
1%
1-
12
#161980000000
0!
0%
b11 *
0-
02
b11 6
#161990000000
1!
1%
1-
12
15
#162000000000
0!
0%
b100 *
0-
02
b100 6
#162010000000
1!
1%
1-
12
#162020000000
0!
0%
b101 *
0-
02
b101 6
#162030000000
1!
1%
1-
12
#162040000000
0!
0%
b110 *
0-
02
b110 6
#162050000000
1!
1%
1-
12
#162060000000
0!
0%
b111 *
0-
02
b111 6
#162070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#162080000000
0!
0%
b0 *
0-
02
b0 6
#162090000000
1!
1%
1-
12
#162100000000
0!
0%
b1 *
0-
02
b1 6
#162110000000
1!
1%
1-
12
#162120000000
0!
0%
b10 *
0-
02
b10 6
#162130000000
1!
1%
1-
12
#162140000000
0!
0%
b11 *
0-
02
b11 6
#162150000000
1!
1%
1-
12
15
#162160000000
0!
0%
b100 *
0-
02
b100 6
#162170000000
1!
1%
1-
12
#162180000000
0!
0%
b101 *
0-
02
b101 6
#162190000000
1!
1%
1-
12
#162200000000
0!
0%
b110 *
0-
02
b110 6
#162210000000
1!
1%
1-
12
#162220000000
0!
0%
b111 *
0-
02
b111 6
#162230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#162240000000
0!
0%
b0 *
0-
02
b0 6
#162250000000
1!
1%
1-
12
#162260000000
0!
0%
b1 *
0-
02
b1 6
#162270000000
1!
1%
1-
12
#162280000000
0!
0%
b10 *
0-
02
b10 6
#162290000000
1!
1%
1-
12
#162300000000
0!
0%
b11 *
0-
02
b11 6
#162310000000
1!
1%
1-
12
15
#162320000000
0!
0%
b100 *
0-
02
b100 6
#162330000000
1!
1%
1-
12
#162340000000
0!
0%
b101 *
0-
02
b101 6
#162350000000
1!
1%
1-
12
#162360000000
0!
0%
b110 *
0-
02
b110 6
#162370000000
1!
1%
1-
12
#162380000000
0!
0%
b111 *
0-
02
b111 6
#162390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#162400000000
0!
0%
b0 *
0-
02
b0 6
#162410000000
1!
1%
1-
12
#162420000000
0!
0%
b1 *
0-
02
b1 6
#162430000000
1!
1%
1-
12
#162440000000
0!
0%
b10 *
0-
02
b10 6
#162450000000
1!
1%
1-
12
#162460000000
0!
0%
b11 *
0-
02
b11 6
#162470000000
1!
1%
1-
12
15
#162480000000
0!
0%
b100 *
0-
02
b100 6
#162490000000
1!
1%
1-
12
#162500000000
0!
0%
b101 *
0-
02
b101 6
#162510000000
1!
1%
1-
12
#162520000000
0!
0%
b110 *
0-
02
b110 6
#162530000000
1!
1%
1-
12
#162540000000
0!
0%
b111 *
0-
02
b111 6
#162550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#162560000000
0!
0%
b0 *
0-
02
b0 6
#162570000000
1!
1%
1-
12
#162580000000
0!
0%
b1 *
0-
02
b1 6
#162590000000
1!
1%
1-
12
#162600000000
0!
0%
b10 *
0-
02
b10 6
#162610000000
1!
1%
1-
12
#162620000000
0!
0%
b11 *
0-
02
b11 6
#162630000000
1!
1%
1-
12
15
#162640000000
0!
0%
b100 *
0-
02
b100 6
#162650000000
1!
1%
1-
12
#162660000000
0!
0%
b101 *
0-
02
b101 6
#162670000000
1!
1%
1-
12
#162680000000
0!
0%
b110 *
0-
02
b110 6
#162690000000
1!
1%
1-
12
#162700000000
0!
0%
b111 *
0-
02
b111 6
#162710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#162720000000
0!
0%
b0 *
0-
02
b0 6
#162730000000
1!
1%
1-
12
#162740000000
0!
0%
b1 *
0-
02
b1 6
#162750000000
1!
1%
1-
12
#162760000000
0!
0%
b10 *
0-
02
b10 6
#162770000000
1!
1%
1-
12
#162780000000
0!
0%
b11 *
0-
02
b11 6
#162790000000
1!
1%
1-
12
15
#162800000000
0!
0%
b100 *
0-
02
b100 6
#162810000000
1!
1%
1-
12
#162820000000
0!
0%
b101 *
0-
02
b101 6
#162830000000
1!
1%
1-
12
#162840000000
0!
0%
b110 *
0-
02
b110 6
#162850000000
1!
1%
1-
12
#162860000000
0!
0%
b111 *
0-
02
b111 6
#162870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#162880000000
0!
0%
b0 *
0-
02
b0 6
#162890000000
1!
1%
1-
12
#162900000000
0!
0%
b1 *
0-
02
b1 6
#162910000000
1!
1%
1-
12
#162920000000
0!
0%
b10 *
0-
02
b10 6
#162930000000
1!
1%
1-
12
#162940000000
0!
0%
b11 *
0-
02
b11 6
#162950000000
1!
1%
1-
12
15
#162960000000
0!
0%
b100 *
0-
02
b100 6
#162970000000
1!
1%
1-
12
#162980000000
0!
0%
b101 *
0-
02
b101 6
#162990000000
1!
1%
1-
12
#163000000000
0!
0%
b110 *
0-
02
b110 6
#163010000000
1!
1%
1-
12
#163020000000
0!
0%
b111 *
0-
02
b111 6
#163030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#163040000000
0!
0%
b0 *
0-
02
b0 6
#163050000000
1!
1%
1-
12
#163060000000
0!
0%
b1 *
0-
02
b1 6
#163070000000
1!
1%
1-
12
#163080000000
0!
0%
b10 *
0-
02
b10 6
#163090000000
1!
1%
1-
12
#163100000000
0!
0%
b11 *
0-
02
b11 6
#163110000000
1!
1%
1-
12
15
#163120000000
0!
0%
b100 *
0-
02
b100 6
#163130000000
1!
1%
1-
12
#163140000000
0!
0%
b101 *
0-
02
b101 6
#163150000000
1!
1%
1-
12
#163160000000
0!
0%
b110 *
0-
02
b110 6
#163170000000
1!
1%
1-
12
#163180000000
0!
0%
b111 *
0-
02
b111 6
#163190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#163200000000
0!
0%
b0 *
0-
02
b0 6
#163210000000
1!
1%
1-
12
#163220000000
0!
0%
b1 *
0-
02
b1 6
#163230000000
1!
1%
1-
12
#163240000000
0!
0%
b10 *
0-
02
b10 6
#163250000000
1!
1%
1-
12
#163260000000
0!
0%
b11 *
0-
02
b11 6
#163270000000
1!
1%
1-
12
15
#163280000000
0!
0%
b100 *
0-
02
b100 6
#163290000000
1!
1%
1-
12
#163300000000
0!
0%
b101 *
0-
02
b101 6
#163310000000
1!
1%
1-
12
#163320000000
0!
0%
b110 *
0-
02
b110 6
#163330000000
1!
1%
1-
12
#163340000000
0!
0%
b111 *
0-
02
b111 6
#163350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#163360000000
0!
0%
b0 *
0-
02
b0 6
#163370000000
1!
1%
1-
12
#163380000000
0!
0%
b1 *
0-
02
b1 6
#163390000000
1!
1%
1-
12
#163400000000
0!
0%
b10 *
0-
02
b10 6
#163410000000
1!
1%
1-
12
#163420000000
0!
0%
b11 *
0-
02
b11 6
#163430000000
1!
1%
1-
12
15
#163440000000
0!
0%
b100 *
0-
02
b100 6
#163450000000
1!
1%
1-
12
#163460000000
0!
0%
b101 *
0-
02
b101 6
#163470000000
1!
1%
1-
12
#163480000000
0!
0%
b110 *
0-
02
b110 6
#163490000000
1!
1%
1-
12
#163500000000
0!
0%
b111 *
0-
02
b111 6
#163510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#163520000000
0!
0%
b0 *
0-
02
b0 6
#163530000000
1!
1%
1-
12
#163540000000
0!
0%
b1 *
0-
02
b1 6
#163550000000
1!
1%
1-
12
#163560000000
0!
0%
b10 *
0-
02
b10 6
#163570000000
1!
1%
1-
12
#163580000000
0!
0%
b11 *
0-
02
b11 6
#163590000000
1!
1%
1-
12
15
#163600000000
0!
0%
b100 *
0-
02
b100 6
#163610000000
1!
1%
1-
12
#163620000000
0!
0%
b101 *
0-
02
b101 6
#163630000000
1!
1%
1-
12
#163640000000
0!
0%
b110 *
0-
02
b110 6
#163650000000
1!
1%
1-
12
#163660000000
0!
0%
b111 *
0-
02
b111 6
#163670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#163680000000
0!
0%
b0 *
0-
02
b0 6
#163690000000
1!
1%
1-
12
#163700000000
0!
0%
b1 *
0-
02
b1 6
#163710000000
1!
1%
1-
12
#163720000000
0!
0%
b10 *
0-
02
b10 6
#163730000000
1!
1%
1-
12
#163740000000
0!
0%
b11 *
0-
02
b11 6
#163750000000
1!
1%
1-
12
15
#163760000000
0!
0%
b100 *
0-
02
b100 6
#163770000000
1!
1%
1-
12
#163780000000
0!
0%
b101 *
0-
02
b101 6
#163790000000
1!
1%
1-
12
#163800000000
0!
0%
b110 *
0-
02
b110 6
#163810000000
1!
1%
1-
12
#163820000000
0!
0%
b111 *
0-
02
b111 6
#163830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#163840000000
0!
0%
b0 *
0-
02
b0 6
#163850000000
1!
1%
1-
12
#163860000000
0!
0%
b1 *
0-
02
b1 6
#163870000000
1!
1%
1-
12
#163880000000
0!
0%
b10 *
0-
02
b10 6
#163890000000
1!
1%
1-
12
#163900000000
0!
0%
b11 *
0-
02
b11 6
#163910000000
1!
1%
1-
12
15
#163920000000
0!
0%
b100 *
0-
02
b100 6
#163930000000
1!
1%
1-
12
#163940000000
0!
0%
b101 *
0-
02
b101 6
#163950000000
1!
1%
1-
12
#163960000000
0!
0%
b110 *
0-
02
b110 6
#163970000000
1!
1%
1-
12
#163980000000
0!
0%
b111 *
0-
02
b111 6
#163990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#164000000000
0!
0%
b0 *
0-
02
b0 6
#164010000000
1!
1%
1-
12
#164020000000
0!
0%
b1 *
0-
02
b1 6
#164030000000
1!
1%
1-
12
#164040000000
0!
0%
b10 *
0-
02
b10 6
#164050000000
1!
1%
1-
12
#164060000000
0!
0%
b11 *
0-
02
b11 6
#164070000000
1!
1%
1-
12
15
#164080000000
0!
0%
b100 *
0-
02
b100 6
#164090000000
1!
1%
1-
12
#164100000000
0!
0%
b101 *
0-
02
b101 6
#164110000000
1!
1%
1-
12
#164120000000
0!
0%
b110 *
0-
02
b110 6
#164130000000
1!
1%
1-
12
#164140000000
0!
0%
b111 *
0-
02
b111 6
#164150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#164160000000
0!
0%
b0 *
0-
02
b0 6
#164170000000
1!
1%
1-
12
#164180000000
0!
0%
b1 *
0-
02
b1 6
#164190000000
1!
1%
1-
12
#164200000000
0!
0%
b10 *
0-
02
b10 6
#164210000000
1!
1%
1-
12
#164220000000
0!
0%
b11 *
0-
02
b11 6
#164230000000
1!
1%
1-
12
15
#164240000000
0!
0%
b100 *
0-
02
b100 6
#164250000000
1!
1%
1-
12
#164260000000
0!
0%
b101 *
0-
02
b101 6
#164270000000
1!
1%
1-
12
#164280000000
0!
0%
b110 *
0-
02
b110 6
#164290000000
1!
1%
1-
12
#164300000000
0!
0%
b111 *
0-
02
b111 6
#164310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#164320000000
0!
0%
b0 *
0-
02
b0 6
#164330000000
1!
1%
1-
12
#164340000000
0!
0%
b1 *
0-
02
b1 6
#164350000000
1!
1%
1-
12
#164360000000
0!
0%
b10 *
0-
02
b10 6
#164370000000
1!
1%
1-
12
#164380000000
0!
0%
b11 *
0-
02
b11 6
#164390000000
1!
1%
1-
12
15
#164400000000
0!
0%
b100 *
0-
02
b100 6
#164410000000
1!
1%
1-
12
#164420000000
0!
0%
b101 *
0-
02
b101 6
#164430000000
1!
1%
1-
12
#164440000000
0!
0%
b110 *
0-
02
b110 6
#164450000000
1!
1%
1-
12
#164460000000
0!
0%
b111 *
0-
02
b111 6
#164470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#164480000000
0!
0%
b0 *
0-
02
b0 6
#164490000000
1!
1%
1-
12
#164500000000
0!
0%
b1 *
0-
02
b1 6
#164510000000
1!
1%
1-
12
#164520000000
0!
0%
b10 *
0-
02
b10 6
#164530000000
1!
1%
1-
12
#164540000000
0!
0%
b11 *
0-
02
b11 6
#164550000000
1!
1%
1-
12
15
#164560000000
0!
0%
b100 *
0-
02
b100 6
#164570000000
1!
1%
1-
12
#164580000000
0!
0%
b101 *
0-
02
b101 6
#164590000000
1!
1%
1-
12
#164600000000
0!
0%
b110 *
0-
02
b110 6
#164610000000
1!
1%
1-
12
#164620000000
0!
0%
b111 *
0-
02
b111 6
#164630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#164640000000
0!
0%
b0 *
0-
02
b0 6
#164650000000
1!
1%
1-
12
#164660000000
0!
0%
b1 *
0-
02
b1 6
#164670000000
1!
1%
1-
12
#164680000000
0!
0%
b10 *
0-
02
b10 6
#164690000000
1!
1%
1-
12
#164700000000
0!
0%
b11 *
0-
02
b11 6
#164710000000
1!
1%
1-
12
15
#164720000000
0!
0%
b100 *
0-
02
b100 6
#164730000000
1!
1%
1-
12
#164740000000
0!
0%
b101 *
0-
02
b101 6
#164750000000
1!
1%
1-
12
#164760000000
0!
0%
b110 *
0-
02
b110 6
#164770000000
1!
1%
1-
12
#164780000000
0!
0%
b111 *
0-
02
b111 6
#164790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#164800000000
0!
0%
b0 *
0-
02
b0 6
#164810000000
1!
1%
1-
12
#164820000000
0!
0%
b1 *
0-
02
b1 6
#164830000000
1!
1%
1-
12
#164840000000
0!
0%
b10 *
0-
02
b10 6
#164850000000
1!
1%
1-
12
#164860000000
0!
0%
b11 *
0-
02
b11 6
#164870000000
1!
1%
1-
12
15
#164880000000
0!
0%
b100 *
0-
02
b100 6
#164890000000
1!
1%
1-
12
#164900000000
0!
0%
b101 *
0-
02
b101 6
#164910000000
1!
1%
1-
12
#164920000000
0!
0%
b110 *
0-
02
b110 6
#164930000000
1!
1%
1-
12
#164940000000
0!
0%
b111 *
0-
02
b111 6
#164950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#164960000000
0!
0%
b0 *
0-
02
b0 6
#164970000000
1!
1%
1-
12
#164980000000
0!
0%
b1 *
0-
02
b1 6
#164990000000
1!
1%
1-
12
#165000000000
0!
0%
b10 *
0-
02
b10 6
#165010000000
1!
1%
1-
12
#165020000000
0!
0%
b11 *
0-
02
b11 6
#165030000000
1!
1%
1-
12
15
#165040000000
0!
0%
b100 *
0-
02
b100 6
#165050000000
1!
1%
1-
12
#165060000000
0!
0%
b101 *
0-
02
b101 6
#165070000000
1!
1%
1-
12
#165080000000
0!
0%
b110 *
0-
02
b110 6
#165090000000
1!
1%
1-
12
#165100000000
0!
0%
b111 *
0-
02
b111 6
#165110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#165120000000
0!
0%
b0 *
0-
02
b0 6
#165130000000
1!
1%
1-
12
#165140000000
0!
0%
b1 *
0-
02
b1 6
#165150000000
1!
1%
1-
12
#165160000000
0!
0%
b10 *
0-
02
b10 6
#165170000000
1!
1%
1-
12
#165180000000
0!
0%
b11 *
0-
02
b11 6
#165190000000
1!
1%
1-
12
15
#165200000000
0!
0%
b100 *
0-
02
b100 6
#165210000000
1!
1%
1-
12
#165220000000
0!
0%
b101 *
0-
02
b101 6
#165230000000
1!
1%
1-
12
#165240000000
0!
0%
b110 *
0-
02
b110 6
#165250000000
1!
1%
1-
12
#165260000000
0!
0%
b111 *
0-
02
b111 6
#165270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#165280000000
0!
0%
b0 *
0-
02
b0 6
#165290000000
1!
1%
1-
12
#165300000000
0!
0%
b1 *
0-
02
b1 6
#165310000000
1!
1%
1-
12
#165320000000
0!
0%
b10 *
0-
02
b10 6
#165330000000
1!
1%
1-
12
#165340000000
0!
0%
b11 *
0-
02
b11 6
#165350000000
1!
1%
1-
12
15
#165360000000
0!
0%
b100 *
0-
02
b100 6
#165370000000
1!
1%
1-
12
#165380000000
0!
0%
b101 *
0-
02
b101 6
#165390000000
1!
1%
1-
12
#165400000000
0!
0%
b110 *
0-
02
b110 6
#165410000000
1!
1%
1-
12
#165420000000
0!
0%
b111 *
0-
02
b111 6
#165430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#165440000000
0!
0%
b0 *
0-
02
b0 6
#165450000000
1!
1%
1-
12
#165460000000
0!
0%
b1 *
0-
02
b1 6
#165470000000
1!
1%
1-
12
#165480000000
0!
0%
b10 *
0-
02
b10 6
#165490000000
1!
1%
1-
12
#165500000000
0!
0%
b11 *
0-
02
b11 6
#165510000000
1!
1%
1-
12
15
#165520000000
0!
0%
b100 *
0-
02
b100 6
#165530000000
1!
1%
1-
12
#165540000000
0!
0%
b101 *
0-
02
b101 6
#165550000000
1!
1%
1-
12
#165560000000
0!
0%
b110 *
0-
02
b110 6
#165570000000
1!
1%
1-
12
#165580000000
0!
0%
b111 *
0-
02
b111 6
#165590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#165600000000
0!
0%
b0 *
0-
02
b0 6
#165610000000
1!
1%
1-
12
#165620000000
0!
0%
b1 *
0-
02
b1 6
#165630000000
1!
1%
1-
12
#165640000000
0!
0%
b10 *
0-
02
b10 6
#165650000000
1!
1%
1-
12
#165660000000
0!
0%
b11 *
0-
02
b11 6
#165670000000
1!
1%
1-
12
15
#165680000000
0!
0%
b100 *
0-
02
b100 6
#165690000000
1!
1%
1-
12
#165700000000
0!
0%
b101 *
0-
02
b101 6
#165710000000
1!
1%
1-
12
#165720000000
0!
0%
b110 *
0-
02
b110 6
#165730000000
1!
1%
1-
12
#165740000000
0!
0%
b111 *
0-
02
b111 6
#165750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#165760000000
0!
0%
b0 *
0-
02
b0 6
#165770000000
1!
1%
1-
12
#165780000000
0!
0%
b1 *
0-
02
b1 6
#165790000000
1!
1%
1-
12
#165800000000
0!
0%
b10 *
0-
02
b10 6
#165810000000
1!
1%
1-
12
#165820000000
0!
0%
b11 *
0-
02
b11 6
#165830000000
1!
1%
1-
12
15
#165840000000
0!
0%
b100 *
0-
02
b100 6
#165850000000
1!
1%
1-
12
#165860000000
0!
0%
b101 *
0-
02
b101 6
#165870000000
1!
1%
1-
12
#165880000000
0!
0%
b110 *
0-
02
b110 6
#165890000000
1!
1%
1-
12
#165900000000
0!
0%
b111 *
0-
02
b111 6
#165910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#165920000000
0!
0%
b0 *
0-
02
b0 6
#165930000000
1!
1%
1-
12
#165940000000
0!
0%
b1 *
0-
02
b1 6
#165950000000
1!
1%
1-
12
#165960000000
0!
0%
b10 *
0-
02
b10 6
#165970000000
1!
1%
1-
12
#165980000000
0!
0%
b11 *
0-
02
b11 6
#165990000000
1!
1%
1-
12
15
#166000000000
0!
0%
b100 *
0-
02
b100 6
#166010000000
1!
1%
1-
12
#166020000000
0!
0%
b101 *
0-
02
b101 6
#166030000000
1!
1%
1-
12
#166040000000
0!
0%
b110 *
0-
02
b110 6
#166050000000
1!
1%
1-
12
#166060000000
0!
0%
b111 *
0-
02
b111 6
#166070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#166080000000
0!
0%
b0 *
0-
02
b0 6
#166090000000
1!
1%
1-
12
#166100000000
0!
0%
b1 *
0-
02
b1 6
#166110000000
1!
1%
1-
12
#166120000000
0!
0%
b10 *
0-
02
b10 6
#166130000000
1!
1%
1-
12
#166140000000
0!
0%
b11 *
0-
02
b11 6
#166150000000
1!
1%
1-
12
15
#166160000000
0!
0%
b100 *
0-
02
b100 6
#166170000000
1!
1%
1-
12
#166180000000
0!
0%
b101 *
0-
02
b101 6
#166190000000
1!
1%
1-
12
#166200000000
0!
0%
b110 *
0-
02
b110 6
#166210000000
1!
1%
1-
12
#166220000000
0!
0%
b111 *
0-
02
b111 6
#166230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#166240000000
0!
0%
b0 *
0-
02
b0 6
#166250000000
1!
1%
1-
12
#166260000000
0!
0%
b1 *
0-
02
b1 6
#166270000000
1!
1%
1-
12
#166280000000
0!
0%
b10 *
0-
02
b10 6
#166290000000
1!
1%
1-
12
#166300000000
0!
0%
b11 *
0-
02
b11 6
#166310000000
1!
1%
1-
12
15
#166320000000
0!
0%
b100 *
0-
02
b100 6
#166330000000
1!
1%
1-
12
#166340000000
0!
0%
b101 *
0-
02
b101 6
#166350000000
1!
1%
1-
12
#166360000000
0!
0%
b110 *
0-
02
b110 6
#166370000000
1!
1%
1-
12
#166380000000
0!
0%
b111 *
0-
02
b111 6
#166390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#166400000000
0!
0%
b0 *
0-
02
b0 6
#166410000000
1!
1%
1-
12
#166420000000
0!
0%
b1 *
0-
02
b1 6
#166430000000
1!
1%
1-
12
#166440000000
0!
0%
b10 *
0-
02
b10 6
#166450000000
1!
1%
1-
12
#166460000000
0!
0%
b11 *
0-
02
b11 6
#166470000000
1!
1%
1-
12
15
#166480000000
0!
0%
b100 *
0-
02
b100 6
#166490000000
1!
1%
1-
12
#166500000000
0!
0%
b101 *
0-
02
b101 6
#166510000000
1!
1%
1-
12
#166520000000
0!
0%
b110 *
0-
02
b110 6
#166530000000
1!
1%
1-
12
#166540000000
0!
0%
b111 *
0-
02
b111 6
#166550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#166560000000
0!
0%
b0 *
0-
02
b0 6
#166570000000
1!
1%
1-
12
#166580000000
0!
0%
b1 *
0-
02
b1 6
#166590000000
1!
1%
1-
12
#166600000000
0!
0%
b10 *
0-
02
b10 6
#166610000000
1!
1%
1-
12
#166620000000
0!
0%
b11 *
0-
02
b11 6
#166630000000
1!
1%
1-
12
15
#166640000000
0!
0%
b100 *
0-
02
b100 6
#166650000000
1!
1%
1-
12
#166660000000
0!
0%
b101 *
0-
02
b101 6
#166670000000
1!
1%
1-
12
#166680000000
0!
0%
b110 *
0-
02
b110 6
#166690000000
1!
1%
1-
12
#166700000000
0!
0%
b111 *
0-
02
b111 6
#166710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#166720000000
0!
0%
b0 *
0-
02
b0 6
#166730000000
1!
1%
1-
12
#166740000000
0!
0%
b1 *
0-
02
b1 6
#166750000000
1!
1%
1-
12
#166760000000
0!
0%
b10 *
0-
02
b10 6
#166770000000
1!
1%
1-
12
#166780000000
0!
0%
b11 *
0-
02
b11 6
#166790000000
1!
1%
1-
12
15
#166800000000
0!
0%
b100 *
0-
02
b100 6
#166810000000
1!
1%
1-
12
#166820000000
0!
0%
b101 *
0-
02
b101 6
#166830000000
1!
1%
1-
12
#166840000000
0!
0%
b110 *
0-
02
b110 6
#166850000000
1!
1%
1-
12
#166860000000
0!
0%
b111 *
0-
02
b111 6
#166870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#166880000000
0!
0%
b0 *
0-
02
b0 6
#166890000000
1!
1%
1-
12
#166900000000
0!
0%
b1 *
0-
02
b1 6
#166910000000
1!
1%
1-
12
#166920000000
0!
0%
b10 *
0-
02
b10 6
#166930000000
1!
1%
1-
12
#166940000000
0!
0%
b11 *
0-
02
b11 6
#166950000000
1!
1%
1-
12
15
#166960000000
0!
0%
b100 *
0-
02
b100 6
#166970000000
1!
1%
1-
12
#166980000000
0!
0%
b101 *
0-
02
b101 6
#166990000000
1!
1%
1-
12
#167000000000
0!
0%
b110 *
0-
02
b110 6
#167010000000
1!
1%
1-
12
#167020000000
0!
0%
b111 *
0-
02
b111 6
#167030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#167040000000
0!
0%
b0 *
0-
02
b0 6
#167050000000
1!
1%
1-
12
#167060000000
0!
0%
b1 *
0-
02
b1 6
#167070000000
1!
1%
1-
12
#167080000000
0!
0%
b10 *
0-
02
b10 6
#167090000000
1!
1%
1-
12
#167100000000
0!
0%
b11 *
0-
02
b11 6
#167110000000
1!
1%
1-
12
15
#167120000000
0!
0%
b100 *
0-
02
b100 6
#167130000000
1!
1%
1-
12
#167140000000
0!
0%
b101 *
0-
02
b101 6
#167150000000
1!
1%
1-
12
#167160000000
0!
0%
b110 *
0-
02
b110 6
#167170000000
1!
1%
1-
12
#167180000000
0!
0%
b111 *
0-
02
b111 6
#167190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#167200000000
0!
0%
b0 *
0-
02
b0 6
#167210000000
1!
1%
1-
12
#167220000000
0!
0%
b1 *
0-
02
b1 6
#167230000000
1!
1%
1-
12
#167240000000
0!
0%
b10 *
0-
02
b10 6
#167250000000
1!
1%
1-
12
#167260000000
0!
0%
b11 *
0-
02
b11 6
#167270000000
1!
1%
1-
12
15
#167280000000
0!
0%
b100 *
0-
02
b100 6
#167290000000
1!
1%
1-
12
#167300000000
0!
0%
b101 *
0-
02
b101 6
#167310000000
1!
1%
1-
12
#167320000000
0!
0%
b110 *
0-
02
b110 6
#167330000000
1!
1%
1-
12
#167340000000
0!
0%
b111 *
0-
02
b111 6
#167350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#167360000000
0!
0%
b0 *
0-
02
b0 6
#167370000000
1!
1%
1-
12
#167380000000
0!
0%
b1 *
0-
02
b1 6
#167390000000
1!
1%
1-
12
#167400000000
0!
0%
b10 *
0-
02
b10 6
#167410000000
1!
1%
1-
12
#167420000000
0!
0%
b11 *
0-
02
b11 6
#167430000000
1!
1%
1-
12
15
#167440000000
0!
0%
b100 *
0-
02
b100 6
#167450000000
1!
1%
1-
12
#167460000000
0!
0%
b101 *
0-
02
b101 6
#167470000000
1!
1%
1-
12
#167480000000
0!
0%
b110 *
0-
02
b110 6
#167490000000
1!
1%
1-
12
#167500000000
0!
0%
b111 *
0-
02
b111 6
#167510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#167520000000
0!
0%
b0 *
0-
02
b0 6
#167530000000
1!
1%
1-
12
#167540000000
0!
0%
b1 *
0-
02
b1 6
#167550000000
1!
1%
1-
12
#167560000000
0!
0%
b10 *
0-
02
b10 6
#167570000000
1!
1%
1-
12
#167580000000
0!
0%
b11 *
0-
02
b11 6
#167590000000
1!
1%
1-
12
15
#167600000000
0!
0%
b100 *
0-
02
b100 6
#167610000000
1!
1%
1-
12
#167620000000
0!
0%
b101 *
0-
02
b101 6
#167630000000
1!
1%
1-
12
#167640000000
0!
0%
b110 *
0-
02
b110 6
#167650000000
1!
1%
1-
12
#167660000000
0!
0%
b111 *
0-
02
b111 6
#167670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#167680000000
0!
0%
b0 *
0-
02
b0 6
#167690000000
1!
1%
1-
12
#167700000000
0!
0%
b1 *
0-
02
b1 6
#167710000000
1!
1%
1-
12
#167720000000
0!
0%
b10 *
0-
02
b10 6
#167730000000
1!
1%
1-
12
#167740000000
0!
0%
b11 *
0-
02
b11 6
#167750000000
1!
1%
1-
12
15
#167760000000
0!
0%
b100 *
0-
02
b100 6
#167770000000
1!
1%
1-
12
#167780000000
0!
0%
b101 *
0-
02
b101 6
#167790000000
1!
1%
1-
12
#167800000000
0!
0%
b110 *
0-
02
b110 6
#167810000000
1!
1%
1-
12
#167820000000
0!
0%
b111 *
0-
02
b111 6
#167830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#167840000000
0!
0%
b0 *
0-
02
b0 6
#167850000000
1!
1%
1-
12
#167860000000
0!
0%
b1 *
0-
02
b1 6
#167870000000
1!
1%
1-
12
#167880000000
0!
0%
b10 *
0-
02
b10 6
#167890000000
1!
1%
1-
12
#167900000000
0!
0%
b11 *
0-
02
b11 6
#167910000000
1!
1%
1-
12
15
#167920000000
0!
0%
b100 *
0-
02
b100 6
#167930000000
1!
1%
1-
12
#167940000000
0!
0%
b101 *
0-
02
b101 6
#167950000000
1!
1%
1-
12
#167960000000
0!
0%
b110 *
0-
02
b110 6
#167970000000
1!
1%
1-
12
#167980000000
0!
0%
b111 *
0-
02
b111 6
#167990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#168000000000
0!
0%
b0 *
0-
02
b0 6
#168010000000
1!
1%
1-
12
#168020000000
0!
0%
b1 *
0-
02
b1 6
#168030000000
1!
1%
1-
12
#168040000000
0!
0%
b10 *
0-
02
b10 6
#168050000000
1!
1%
1-
12
#168060000000
0!
0%
b11 *
0-
02
b11 6
#168070000000
1!
1%
1-
12
15
#168080000000
0!
0%
b100 *
0-
02
b100 6
#168090000000
1!
1%
1-
12
#168100000000
0!
0%
b101 *
0-
02
b101 6
#168110000000
1!
1%
1-
12
#168120000000
0!
0%
b110 *
0-
02
b110 6
#168130000000
1!
1%
1-
12
#168140000000
0!
0%
b111 *
0-
02
b111 6
#168150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#168160000000
0!
0%
b0 *
0-
02
b0 6
#168170000000
1!
1%
1-
12
#168180000000
0!
0%
b1 *
0-
02
b1 6
#168190000000
1!
1%
1-
12
#168200000000
0!
0%
b10 *
0-
02
b10 6
#168210000000
1!
1%
1-
12
#168220000000
0!
0%
b11 *
0-
02
b11 6
#168230000000
1!
1%
1-
12
15
#168240000000
0!
0%
b100 *
0-
02
b100 6
#168250000000
1!
1%
1-
12
#168260000000
0!
0%
b101 *
0-
02
b101 6
#168270000000
1!
1%
1-
12
#168280000000
0!
0%
b110 *
0-
02
b110 6
#168290000000
1!
1%
1-
12
#168300000000
0!
0%
b111 *
0-
02
b111 6
#168310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#168320000000
0!
0%
b0 *
0-
02
b0 6
#168330000000
1!
1%
1-
12
#168340000000
0!
0%
b1 *
0-
02
b1 6
#168350000000
1!
1%
1-
12
#168360000000
0!
0%
b10 *
0-
02
b10 6
#168370000000
1!
1%
1-
12
#168380000000
0!
0%
b11 *
0-
02
b11 6
#168390000000
1!
1%
1-
12
15
#168400000000
0!
0%
b100 *
0-
02
b100 6
#168410000000
1!
1%
1-
12
#168420000000
0!
0%
b101 *
0-
02
b101 6
#168430000000
1!
1%
1-
12
#168440000000
0!
0%
b110 *
0-
02
b110 6
#168450000000
1!
1%
1-
12
#168460000000
0!
0%
b111 *
0-
02
b111 6
#168470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#168480000000
0!
0%
b0 *
0-
02
b0 6
#168490000000
1!
1%
1-
12
#168500000000
0!
0%
b1 *
0-
02
b1 6
#168510000000
1!
1%
1-
12
#168520000000
0!
0%
b10 *
0-
02
b10 6
#168530000000
1!
1%
1-
12
#168540000000
0!
0%
b11 *
0-
02
b11 6
#168550000000
1!
1%
1-
12
15
#168560000000
0!
0%
b100 *
0-
02
b100 6
#168570000000
1!
1%
1-
12
#168580000000
0!
0%
b101 *
0-
02
b101 6
#168590000000
1!
1%
1-
12
#168600000000
0!
0%
b110 *
0-
02
b110 6
#168610000000
1!
1%
1-
12
#168620000000
0!
0%
b111 *
0-
02
b111 6
#168630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#168640000000
0!
0%
b0 *
0-
02
b0 6
#168650000000
1!
1%
1-
12
#168660000000
0!
0%
b1 *
0-
02
b1 6
#168670000000
1!
1%
1-
12
#168680000000
0!
0%
b10 *
0-
02
b10 6
#168690000000
1!
1%
1-
12
#168700000000
0!
0%
b11 *
0-
02
b11 6
#168710000000
1!
1%
1-
12
15
#168720000000
0!
0%
b100 *
0-
02
b100 6
#168730000000
1!
1%
1-
12
#168740000000
0!
0%
b101 *
0-
02
b101 6
#168750000000
1!
1%
1-
12
#168760000000
0!
0%
b110 *
0-
02
b110 6
#168770000000
1!
1%
1-
12
#168780000000
0!
0%
b111 *
0-
02
b111 6
#168790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#168800000000
0!
0%
b0 *
0-
02
b0 6
#168810000000
1!
1%
1-
12
#168820000000
0!
0%
b1 *
0-
02
b1 6
#168830000000
1!
1%
1-
12
#168840000000
0!
0%
b10 *
0-
02
b10 6
#168850000000
1!
1%
1-
12
#168860000000
0!
0%
b11 *
0-
02
b11 6
#168870000000
1!
1%
1-
12
15
#168880000000
0!
0%
b100 *
0-
02
b100 6
#168890000000
1!
1%
1-
12
#168900000000
0!
0%
b101 *
0-
02
b101 6
#168910000000
1!
1%
1-
12
#168920000000
0!
0%
b110 *
0-
02
b110 6
#168930000000
1!
1%
1-
12
#168940000000
0!
0%
b111 *
0-
02
b111 6
#168950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#168960000000
0!
0%
b0 *
0-
02
b0 6
#168970000000
1!
1%
1-
12
#168980000000
0!
0%
b1 *
0-
02
b1 6
#168990000000
1!
1%
1-
12
#169000000000
0!
0%
b10 *
0-
02
b10 6
#169010000000
1!
1%
1-
12
#169020000000
0!
0%
b11 *
0-
02
b11 6
#169030000000
1!
1%
1-
12
15
#169040000000
0!
0%
b100 *
0-
02
b100 6
#169050000000
1!
1%
1-
12
#169060000000
0!
0%
b101 *
0-
02
b101 6
#169070000000
1!
1%
1-
12
#169080000000
0!
0%
b110 *
0-
02
b110 6
#169090000000
1!
1%
1-
12
#169100000000
0!
0%
b111 *
0-
02
b111 6
#169110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#169120000000
0!
0%
b0 *
0-
02
b0 6
#169130000000
1!
1%
1-
12
#169140000000
0!
0%
b1 *
0-
02
b1 6
#169150000000
1!
1%
1-
12
#169160000000
0!
0%
b10 *
0-
02
b10 6
#169170000000
1!
1%
1-
12
#169180000000
0!
0%
b11 *
0-
02
b11 6
#169190000000
1!
1%
1-
12
15
#169200000000
0!
0%
b100 *
0-
02
b100 6
#169210000000
1!
1%
1-
12
#169220000000
0!
0%
b101 *
0-
02
b101 6
#169230000000
1!
1%
1-
12
#169240000000
0!
0%
b110 *
0-
02
b110 6
#169250000000
1!
1%
1-
12
#169260000000
0!
0%
b111 *
0-
02
b111 6
#169270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#169280000000
0!
0%
b0 *
0-
02
b0 6
#169290000000
1!
1%
1-
12
#169300000000
0!
0%
b1 *
0-
02
b1 6
#169310000000
1!
1%
1-
12
#169320000000
0!
0%
b10 *
0-
02
b10 6
#169330000000
1!
1%
1-
12
#169340000000
0!
0%
b11 *
0-
02
b11 6
#169350000000
1!
1%
1-
12
15
#169360000000
0!
0%
b100 *
0-
02
b100 6
#169370000000
1!
1%
1-
12
#169380000000
0!
0%
b101 *
0-
02
b101 6
#169390000000
1!
1%
1-
12
#169400000000
0!
0%
b110 *
0-
02
b110 6
#169410000000
1!
1%
1-
12
#169420000000
0!
0%
b111 *
0-
02
b111 6
#169430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#169440000000
0!
0%
b0 *
0-
02
b0 6
#169450000000
1!
1%
1-
12
#169460000000
0!
0%
b1 *
0-
02
b1 6
#169470000000
1!
1%
1-
12
#169480000000
0!
0%
b10 *
0-
02
b10 6
#169490000000
1!
1%
1-
12
#169500000000
0!
0%
b11 *
0-
02
b11 6
#169510000000
1!
1%
1-
12
15
#169520000000
0!
0%
b100 *
0-
02
b100 6
#169530000000
1!
1%
1-
12
#169540000000
0!
0%
b101 *
0-
02
b101 6
#169550000000
1!
1%
1-
12
#169560000000
0!
0%
b110 *
0-
02
b110 6
#169570000000
1!
1%
1-
12
#169580000000
0!
0%
b111 *
0-
02
b111 6
#169590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#169600000000
0!
0%
b0 *
0-
02
b0 6
#169610000000
1!
1%
1-
12
#169620000000
0!
0%
b1 *
0-
02
b1 6
#169630000000
1!
1%
1-
12
#169640000000
0!
0%
b10 *
0-
02
b10 6
#169650000000
1!
1%
1-
12
#169660000000
0!
0%
b11 *
0-
02
b11 6
#169670000000
1!
1%
1-
12
15
#169680000000
0!
0%
b100 *
0-
02
b100 6
#169690000000
1!
1%
1-
12
#169700000000
0!
0%
b101 *
0-
02
b101 6
#169710000000
1!
1%
1-
12
#169720000000
0!
0%
b110 *
0-
02
b110 6
#169730000000
1!
1%
1-
12
#169740000000
0!
0%
b111 *
0-
02
b111 6
#169750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#169760000000
0!
0%
b0 *
0-
02
b0 6
#169770000000
1!
1%
1-
12
#169780000000
0!
0%
b1 *
0-
02
b1 6
#169790000000
1!
1%
1-
12
#169800000000
0!
0%
b10 *
0-
02
b10 6
#169810000000
1!
1%
1-
12
#169820000000
0!
0%
b11 *
0-
02
b11 6
#169830000000
1!
1%
1-
12
15
#169840000000
0!
0%
b100 *
0-
02
b100 6
#169850000000
1!
1%
1-
12
#169860000000
0!
0%
b101 *
0-
02
b101 6
#169870000000
1!
1%
1-
12
#169880000000
0!
0%
b110 *
0-
02
b110 6
#169890000000
1!
1%
1-
12
#169900000000
0!
0%
b111 *
0-
02
b111 6
#169910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#169920000000
0!
0%
b0 *
0-
02
b0 6
#169930000000
1!
1%
1-
12
#169940000000
0!
0%
b1 *
0-
02
b1 6
#169950000000
1!
1%
1-
12
#169960000000
0!
0%
b10 *
0-
02
b10 6
#169970000000
1!
1%
1-
12
#169980000000
0!
0%
b11 *
0-
02
b11 6
#169990000000
1!
1%
1-
12
15
#170000000000
0!
0%
b100 *
0-
02
b100 6
#170010000000
1!
1%
1-
12
#170020000000
0!
0%
b101 *
0-
02
b101 6
#170030000000
1!
1%
1-
12
#170040000000
0!
0%
b110 *
0-
02
b110 6
#170050000000
1!
1%
1-
12
#170060000000
0!
0%
b111 *
0-
02
b111 6
#170070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#170080000000
0!
0%
b0 *
0-
02
b0 6
#170090000000
1!
1%
1-
12
#170100000000
0!
0%
b1 *
0-
02
b1 6
#170110000000
1!
1%
1-
12
#170120000000
0!
0%
b10 *
0-
02
b10 6
#170130000000
1!
1%
1-
12
#170140000000
0!
0%
b11 *
0-
02
b11 6
#170150000000
1!
1%
1-
12
15
#170160000000
0!
0%
b100 *
0-
02
b100 6
#170170000000
1!
1%
1-
12
#170180000000
0!
0%
b101 *
0-
02
b101 6
#170190000000
1!
1%
1-
12
#170200000000
0!
0%
b110 *
0-
02
b110 6
#170210000000
1!
1%
1-
12
#170220000000
0!
0%
b111 *
0-
02
b111 6
#170230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#170240000000
0!
0%
b0 *
0-
02
b0 6
#170250000000
1!
1%
1-
12
#170260000000
0!
0%
b1 *
0-
02
b1 6
#170270000000
1!
1%
1-
12
#170280000000
0!
0%
b10 *
0-
02
b10 6
#170290000000
1!
1%
1-
12
#170300000000
0!
0%
b11 *
0-
02
b11 6
#170310000000
1!
1%
1-
12
15
#170320000000
0!
0%
b100 *
0-
02
b100 6
#170330000000
1!
1%
1-
12
#170340000000
0!
0%
b101 *
0-
02
b101 6
#170350000000
1!
1%
1-
12
#170360000000
0!
0%
b110 *
0-
02
b110 6
#170370000000
1!
1%
1-
12
#170380000000
0!
0%
b111 *
0-
02
b111 6
#170390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#170400000000
0!
0%
b0 *
0-
02
b0 6
#170410000000
1!
1%
1-
12
#170420000000
0!
0%
b1 *
0-
02
b1 6
#170430000000
1!
1%
1-
12
#170440000000
0!
0%
b10 *
0-
02
b10 6
#170450000000
1!
1%
1-
12
#170460000000
0!
0%
b11 *
0-
02
b11 6
#170470000000
1!
1%
1-
12
15
#170480000000
0!
0%
b100 *
0-
02
b100 6
#170490000000
1!
1%
1-
12
#170500000000
0!
0%
b101 *
0-
02
b101 6
#170510000000
1!
1%
1-
12
#170520000000
0!
0%
b110 *
0-
02
b110 6
#170530000000
1!
1%
1-
12
#170540000000
0!
0%
b111 *
0-
02
b111 6
#170550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#170560000000
0!
0%
b0 *
0-
02
b0 6
#170570000000
1!
1%
1-
12
#170580000000
0!
0%
b1 *
0-
02
b1 6
#170590000000
1!
1%
1-
12
#170600000000
0!
0%
b10 *
0-
02
b10 6
#170610000000
1!
1%
1-
12
#170620000000
0!
0%
b11 *
0-
02
b11 6
#170630000000
1!
1%
1-
12
15
#170640000000
0!
0%
b100 *
0-
02
b100 6
#170650000000
1!
1%
1-
12
#170660000000
0!
0%
b101 *
0-
02
b101 6
#170670000000
1!
1%
1-
12
#170680000000
0!
0%
b110 *
0-
02
b110 6
#170690000000
1!
1%
1-
12
#170700000000
0!
0%
b111 *
0-
02
b111 6
#170710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#170720000000
0!
0%
b0 *
0-
02
b0 6
#170730000000
1!
1%
1-
12
#170740000000
0!
0%
b1 *
0-
02
b1 6
#170750000000
1!
1%
1-
12
#170760000000
0!
0%
b10 *
0-
02
b10 6
#170770000000
1!
1%
1-
12
#170780000000
0!
0%
b11 *
0-
02
b11 6
#170790000000
1!
1%
1-
12
15
#170800000000
0!
0%
b100 *
0-
02
b100 6
#170810000000
1!
1%
1-
12
#170820000000
0!
0%
b101 *
0-
02
b101 6
#170830000000
1!
1%
1-
12
#170840000000
0!
0%
b110 *
0-
02
b110 6
#170850000000
1!
1%
1-
12
#170860000000
0!
0%
b111 *
0-
02
b111 6
#170870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#170880000000
0!
0%
b0 *
0-
02
b0 6
#170890000000
1!
1%
1-
12
#170900000000
0!
0%
b1 *
0-
02
b1 6
#170910000000
1!
1%
1-
12
#170920000000
0!
0%
b10 *
0-
02
b10 6
#170930000000
1!
1%
1-
12
#170940000000
0!
0%
b11 *
0-
02
b11 6
#170950000000
1!
1%
1-
12
15
#170960000000
0!
0%
b100 *
0-
02
b100 6
#170970000000
1!
1%
1-
12
#170980000000
0!
0%
b101 *
0-
02
b101 6
#170990000000
1!
1%
1-
12
#171000000000
0!
0%
b110 *
0-
02
b110 6
#171010000000
1!
1%
1-
12
#171020000000
0!
0%
b111 *
0-
02
b111 6
#171030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#171040000000
0!
0%
b0 *
0-
02
b0 6
#171050000000
1!
1%
1-
12
#171060000000
0!
0%
b1 *
0-
02
b1 6
#171070000000
1!
1%
1-
12
#171080000000
0!
0%
b10 *
0-
02
b10 6
#171090000000
1!
1%
1-
12
#171100000000
0!
0%
b11 *
0-
02
b11 6
#171110000000
1!
1%
1-
12
15
#171120000000
0!
0%
b100 *
0-
02
b100 6
#171130000000
1!
1%
1-
12
#171140000000
0!
0%
b101 *
0-
02
b101 6
#171150000000
1!
1%
1-
12
#171160000000
0!
0%
b110 *
0-
02
b110 6
#171170000000
1!
1%
1-
12
#171180000000
0!
0%
b111 *
0-
02
b111 6
#171190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#171200000000
0!
0%
b0 *
0-
02
b0 6
#171210000000
1!
1%
1-
12
#171220000000
0!
0%
b1 *
0-
02
b1 6
#171230000000
1!
1%
1-
12
#171240000000
0!
0%
b10 *
0-
02
b10 6
#171250000000
1!
1%
1-
12
#171260000000
0!
0%
b11 *
0-
02
b11 6
#171270000000
1!
1%
1-
12
15
#171280000000
0!
0%
b100 *
0-
02
b100 6
#171290000000
1!
1%
1-
12
#171300000000
0!
0%
b101 *
0-
02
b101 6
#171310000000
1!
1%
1-
12
#171320000000
0!
0%
b110 *
0-
02
b110 6
#171330000000
1!
1%
1-
12
#171340000000
0!
0%
b111 *
0-
02
b111 6
#171350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#171360000000
0!
0%
b0 *
0-
02
b0 6
#171370000000
1!
1%
1-
12
#171380000000
0!
0%
b1 *
0-
02
b1 6
#171390000000
1!
1%
1-
12
#171400000000
0!
0%
b10 *
0-
02
b10 6
#171410000000
1!
1%
1-
12
#171420000000
0!
0%
b11 *
0-
02
b11 6
#171430000000
1!
1%
1-
12
15
#171440000000
0!
0%
b100 *
0-
02
b100 6
#171450000000
1!
1%
1-
12
#171460000000
0!
0%
b101 *
0-
02
b101 6
#171470000000
1!
1%
1-
12
#171480000000
0!
0%
b110 *
0-
02
b110 6
#171490000000
1!
1%
1-
12
#171500000000
0!
0%
b111 *
0-
02
b111 6
#171510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#171520000000
0!
0%
b0 *
0-
02
b0 6
#171530000000
1!
1%
1-
12
#171540000000
0!
0%
b1 *
0-
02
b1 6
#171550000000
1!
1%
1-
12
#171560000000
0!
0%
b10 *
0-
02
b10 6
#171570000000
1!
1%
1-
12
#171580000000
0!
0%
b11 *
0-
02
b11 6
#171590000000
1!
1%
1-
12
15
#171600000000
0!
0%
b100 *
0-
02
b100 6
#171610000000
1!
1%
1-
12
#171620000000
0!
0%
b101 *
0-
02
b101 6
#171630000000
1!
1%
1-
12
#171640000000
0!
0%
b110 *
0-
02
b110 6
#171650000000
1!
1%
1-
12
#171660000000
0!
0%
b111 *
0-
02
b111 6
#171670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#171680000000
0!
0%
b0 *
0-
02
b0 6
#171690000000
1!
1%
1-
12
#171700000000
0!
0%
b1 *
0-
02
b1 6
#171710000000
1!
1%
1-
12
#171720000000
0!
0%
b10 *
0-
02
b10 6
#171730000000
1!
1%
1-
12
#171740000000
0!
0%
b11 *
0-
02
b11 6
#171750000000
1!
1%
1-
12
15
#171760000000
0!
0%
b100 *
0-
02
b100 6
#171770000000
1!
1%
1-
12
#171780000000
0!
0%
b101 *
0-
02
b101 6
#171790000000
1!
1%
1-
12
#171800000000
0!
0%
b110 *
0-
02
b110 6
#171810000000
1!
1%
1-
12
#171820000000
0!
0%
b111 *
0-
02
b111 6
#171830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#171840000000
0!
0%
b0 *
0-
02
b0 6
#171850000000
1!
1%
1-
12
#171860000000
0!
0%
b1 *
0-
02
b1 6
#171870000000
1!
1%
1-
12
#171880000000
0!
0%
b10 *
0-
02
b10 6
#171890000000
1!
1%
1-
12
#171900000000
0!
0%
b11 *
0-
02
b11 6
#171910000000
1!
1%
1-
12
15
#171920000000
0!
0%
b100 *
0-
02
b100 6
#171930000000
1!
1%
1-
12
#171940000000
0!
0%
b101 *
0-
02
b101 6
#171950000000
1!
1%
1-
12
#171960000000
0!
0%
b110 *
0-
02
b110 6
#171970000000
1!
1%
1-
12
#171980000000
0!
0%
b111 *
0-
02
b111 6
#171990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#172000000000
0!
0%
b0 *
0-
02
b0 6
#172010000000
1!
1%
1-
12
#172020000000
0!
0%
b1 *
0-
02
b1 6
#172030000000
1!
1%
1-
12
#172040000000
0!
0%
b10 *
0-
02
b10 6
#172050000000
1!
1%
1-
12
#172060000000
0!
0%
b11 *
0-
02
b11 6
#172070000000
1!
1%
1-
12
15
#172080000000
0!
0%
b100 *
0-
02
b100 6
#172090000000
1!
1%
1-
12
#172100000000
0!
0%
b101 *
0-
02
b101 6
#172110000000
1!
1%
1-
12
#172120000000
0!
0%
b110 *
0-
02
b110 6
#172130000000
1!
1%
1-
12
#172140000000
0!
0%
b111 *
0-
02
b111 6
#172150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#172160000000
0!
0%
b0 *
0-
02
b0 6
#172170000000
1!
1%
1-
12
#172180000000
0!
0%
b1 *
0-
02
b1 6
#172190000000
1!
1%
1-
12
#172200000000
0!
0%
b10 *
0-
02
b10 6
#172210000000
1!
1%
1-
12
#172220000000
0!
0%
b11 *
0-
02
b11 6
#172230000000
1!
1%
1-
12
15
#172240000000
0!
0%
b100 *
0-
02
b100 6
#172250000000
1!
1%
1-
12
#172260000000
0!
0%
b101 *
0-
02
b101 6
#172270000000
1!
1%
1-
12
#172280000000
0!
0%
b110 *
0-
02
b110 6
#172290000000
1!
1%
1-
12
#172300000000
0!
0%
b111 *
0-
02
b111 6
#172310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#172320000000
0!
0%
b0 *
0-
02
b0 6
#172330000000
1!
1%
1-
12
#172340000000
0!
0%
b1 *
0-
02
b1 6
#172350000000
1!
1%
1-
12
#172360000000
0!
0%
b10 *
0-
02
b10 6
#172370000000
1!
1%
1-
12
#172380000000
0!
0%
b11 *
0-
02
b11 6
#172390000000
1!
1%
1-
12
15
#172400000000
0!
0%
b100 *
0-
02
b100 6
#172410000000
1!
1%
1-
12
#172420000000
0!
0%
b101 *
0-
02
b101 6
#172430000000
1!
1%
1-
12
#172440000000
0!
0%
b110 *
0-
02
b110 6
#172450000000
1!
1%
1-
12
#172460000000
0!
0%
b111 *
0-
02
b111 6
#172470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#172480000000
0!
0%
b0 *
0-
02
b0 6
#172490000000
1!
1%
1-
12
#172500000000
0!
0%
b1 *
0-
02
b1 6
#172510000000
1!
1%
1-
12
#172520000000
0!
0%
b10 *
0-
02
b10 6
#172530000000
1!
1%
1-
12
#172540000000
0!
0%
b11 *
0-
02
b11 6
#172550000000
1!
1%
1-
12
15
#172560000000
0!
0%
b100 *
0-
02
b100 6
#172570000000
1!
1%
1-
12
#172580000000
0!
0%
b101 *
0-
02
b101 6
#172590000000
1!
1%
1-
12
#172600000000
0!
0%
b110 *
0-
02
b110 6
#172610000000
1!
1%
1-
12
#172620000000
0!
0%
b111 *
0-
02
b111 6
#172630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#172640000000
0!
0%
b0 *
0-
02
b0 6
#172650000000
1!
1%
1-
12
#172660000000
0!
0%
b1 *
0-
02
b1 6
#172670000000
1!
1%
1-
12
#172680000000
0!
0%
b10 *
0-
02
b10 6
#172690000000
1!
1%
1-
12
#172700000000
0!
0%
b11 *
0-
02
b11 6
#172710000000
1!
1%
1-
12
15
#172720000000
0!
0%
b100 *
0-
02
b100 6
#172730000000
1!
1%
1-
12
#172740000000
0!
0%
b101 *
0-
02
b101 6
#172750000000
1!
1%
1-
12
#172760000000
0!
0%
b110 *
0-
02
b110 6
#172770000000
1!
1%
1-
12
#172780000000
0!
0%
b111 *
0-
02
b111 6
#172790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#172800000000
0!
0%
b0 *
0-
02
b0 6
#172810000000
1!
1%
1-
12
#172820000000
0!
0%
b1 *
0-
02
b1 6
#172830000000
1!
1%
1-
12
#172840000000
0!
0%
b10 *
0-
02
b10 6
#172850000000
1!
1%
1-
12
#172860000000
0!
0%
b11 *
0-
02
b11 6
#172870000000
1!
1%
1-
12
15
#172880000000
0!
0%
b100 *
0-
02
b100 6
#172890000000
1!
1%
1-
12
#172900000000
0!
0%
b101 *
0-
02
b101 6
#172910000000
1!
1%
1-
12
#172920000000
0!
0%
b110 *
0-
02
b110 6
#172930000000
1!
1%
1-
12
#172940000000
0!
0%
b111 *
0-
02
b111 6
#172950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#172960000000
0!
0%
b0 *
0-
02
b0 6
#172970000000
1!
1%
1-
12
#172980000000
0!
0%
b1 *
0-
02
b1 6
#172990000000
1!
1%
1-
12
#173000000000
0!
0%
b10 *
0-
02
b10 6
#173010000000
1!
1%
1-
12
#173020000000
0!
0%
b11 *
0-
02
b11 6
#173030000000
1!
1%
1-
12
15
#173040000000
0!
0%
b100 *
0-
02
b100 6
#173050000000
1!
1%
1-
12
#173060000000
0!
0%
b101 *
0-
02
b101 6
#173070000000
1!
1%
1-
12
#173080000000
0!
0%
b110 *
0-
02
b110 6
#173090000000
1!
1%
1-
12
#173100000000
0!
0%
b111 *
0-
02
b111 6
#173110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#173120000000
0!
0%
b0 *
0-
02
b0 6
#173130000000
1!
1%
1-
12
#173140000000
0!
0%
b1 *
0-
02
b1 6
#173150000000
1!
1%
1-
12
#173160000000
0!
0%
b10 *
0-
02
b10 6
#173170000000
1!
1%
1-
12
#173180000000
0!
0%
b11 *
0-
02
b11 6
#173190000000
1!
1%
1-
12
15
#173200000000
0!
0%
b100 *
0-
02
b100 6
#173210000000
1!
1%
1-
12
#173220000000
0!
0%
b101 *
0-
02
b101 6
#173230000000
1!
1%
1-
12
#173240000000
0!
0%
b110 *
0-
02
b110 6
#173250000000
1!
1%
1-
12
#173260000000
0!
0%
b111 *
0-
02
b111 6
#173270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#173280000000
0!
0%
b0 *
0-
02
b0 6
#173290000000
1!
1%
1-
12
#173300000000
0!
0%
b1 *
0-
02
b1 6
#173310000000
1!
1%
1-
12
#173320000000
0!
0%
b10 *
0-
02
b10 6
#173330000000
1!
1%
1-
12
#173340000000
0!
0%
b11 *
0-
02
b11 6
#173350000000
1!
1%
1-
12
15
#173360000000
0!
0%
b100 *
0-
02
b100 6
#173370000000
1!
1%
1-
12
#173380000000
0!
0%
b101 *
0-
02
b101 6
#173390000000
1!
1%
1-
12
#173400000000
0!
0%
b110 *
0-
02
b110 6
#173410000000
1!
1%
1-
12
#173420000000
0!
0%
b111 *
0-
02
b111 6
#173430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#173440000000
0!
0%
b0 *
0-
02
b0 6
#173450000000
1!
1%
1-
12
#173460000000
0!
0%
b1 *
0-
02
b1 6
#173470000000
1!
1%
1-
12
#173480000000
0!
0%
b10 *
0-
02
b10 6
#173490000000
1!
1%
1-
12
#173500000000
0!
0%
b11 *
0-
02
b11 6
#173510000000
1!
1%
1-
12
15
#173520000000
0!
0%
b100 *
0-
02
b100 6
#173530000000
1!
1%
1-
12
#173540000000
0!
0%
b101 *
0-
02
b101 6
#173550000000
1!
1%
1-
12
#173560000000
0!
0%
b110 *
0-
02
b110 6
#173570000000
1!
1%
1-
12
#173580000000
0!
0%
b111 *
0-
02
b111 6
#173590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#173600000000
0!
0%
b0 *
0-
02
b0 6
#173610000000
1!
1%
1-
12
#173620000000
0!
0%
b1 *
0-
02
b1 6
#173630000000
1!
1%
1-
12
#173640000000
0!
0%
b10 *
0-
02
b10 6
#173650000000
1!
1%
1-
12
#173660000000
0!
0%
b11 *
0-
02
b11 6
#173670000000
1!
1%
1-
12
15
#173680000000
0!
0%
b100 *
0-
02
b100 6
#173690000000
1!
1%
1-
12
#173700000000
0!
0%
b101 *
0-
02
b101 6
#173710000000
1!
1%
1-
12
#173720000000
0!
0%
b110 *
0-
02
b110 6
#173730000000
1!
1%
1-
12
#173740000000
0!
0%
b111 *
0-
02
b111 6
#173750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#173760000000
0!
0%
b0 *
0-
02
b0 6
#173770000000
1!
1%
1-
12
#173780000000
0!
0%
b1 *
0-
02
b1 6
#173790000000
1!
1%
1-
12
#173800000000
0!
0%
b10 *
0-
02
b10 6
#173810000000
1!
1%
1-
12
#173820000000
0!
0%
b11 *
0-
02
b11 6
#173830000000
1!
1%
1-
12
15
#173840000000
0!
0%
b100 *
0-
02
b100 6
#173850000000
1!
1%
1-
12
#173860000000
0!
0%
b101 *
0-
02
b101 6
#173870000000
1!
1%
1-
12
#173880000000
0!
0%
b110 *
0-
02
b110 6
#173890000000
1!
1%
1-
12
#173900000000
0!
0%
b111 *
0-
02
b111 6
#173910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#173920000000
0!
0%
b0 *
0-
02
b0 6
#173930000000
1!
1%
1-
12
#173940000000
0!
0%
b1 *
0-
02
b1 6
#173950000000
1!
1%
1-
12
#173960000000
0!
0%
b10 *
0-
02
b10 6
#173970000000
1!
1%
1-
12
#173980000000
0!
0%
b11 *
0-
02
b11 6
#173990000000
1!
1%
1-
12
15
#174000000000
0!
0%
b100 *
0-
02
b100 6
#174010000000
1!
1%
1-
12
#174020000000
0!
0%
b101 *
0-
02
b101 6
#174030000000
1!
1%
1-
12
#174040000000
0!
0%
b110 *
0-
02
b110 6
#174050000000
1!
1%
1-
12
#174060000000
0!
0%
b111 *
0-
02
b111 6
#174070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#174080000000
0!
0%
b0 *
0-
02
b0 6
#174090000000
1!
1%
1-
12
#174100000000
0!
0%
b1 *
0-
02
b1 6
#174110000000
1!
1%
1-
12
#174120000000
0!
0%
b10 *
0-
02
b10 6
#174130000000
1!
1%
1-
12
#174140000000
0!
0%
b11 *
0-
02
b11 6
#174150000000
1!
1%
1-
12
15
#174160000000
0!
0%
b100 *
0-
02
b100 6
#174170000000
1!
1%
1-
12
#174180000000
0!
0%
b101 *
0-
02
b101 6
#174190000000
1!
1%
1-
12
#174200000000
0!
0%
b110 *
0-
02
b110 6
#174210000000
1!
1%
1-
12
#174220000000
0!
0%
b111 *
0-
02
b111 6
#174230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#174240000000
0!
0%
b0 *
0-
02
b0 6
#174250000000
1!
1%
1-
12
#174260000000
0!
0%
b1 *
0-
02
b1 6
#174270000000
1!
1%
1-
12
#174280000000
0!
0%
b10 *
0-
02
b10 6
#174290000000
1!
1%
1-
12
#174300000000
0!
0%
b11 *
0-
02
b11 6
#174310000000
1!
1%
1-
12
15
#174320000000
0!
0%
b100 *
0-
02
b100 6
#174330000000
1!
1%
1-
12
#174340000000
0!
0%
b101 *
0-
02
b101 6
#174350000000
1!
1%
1-
12
#174360000000
0!
0%
b110 *
0-
02
b110 6
#174370000000
1!
1%
1-
12
#174380000000
0!
0%
b111 *
0-
02
b111 6
#174390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#174400000000
0!
0%
b0 *
0-
02
b0 6
#174410000000
1!
1%
1-
12
#174420000000
0!
0%
b1 *
0-
02
b1 6
#174430000000
1!
1%
1-
12
#174440000000
0!
0%
b10 *
0-
02
b10 6
#174450000000
1!
1%
1-
12
#174460000000
0!
0%
b11 *
0-
02
b11 6
#174470000000
1!
1%
1-
12
15
#174480000000
0!
0%
b100 *
0-
02
b100 6
#174490000000
1!
1%
1-
12
#174500000000
0!
0%
b101 *
0-
02
b101 6
#174510000000
1!
1%
1-
12
#174520000000
0!
0%
b110 *
0-
02
b110 6
#174530000000
1!
1%
1-
12
#174540000000
0!
0%
b111 *
0-
02
b111 6
#174550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#174560000000
0!
0%
b0 *
0-
02
b0 6
#174570000000
1!
1%
1-
12
#174580000000
0!
0%
b1 *
0-
02
b1 6
#174590000000
1!
1%
1-
12
#174600000000
0!
0%
b10 *
0-
02
b10 6
#174610000000
1!
1%
1-
12
#174620000000
0!
0%
b11 *
0-
02
b11 6
#174630000000
1!
1%
1-
12
15
#174640000000
0!
0%
b100 *
0-
02
b100 6
#174650000000
1!
1%
1-
12
#174660000000
0!
0%
b101 *
0-
02
b101 6
#174670000000
1!
1%
1-
12
#174680000000
0!
0%
b110 *
0-
02
b110 6
#174690000000
1!
1%
1-
12
#174700000000
0!
0%
b111 *
0-
02
b111 6
#174710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#174720000000
0!
0%
b0 *
0-
02
b0 6
#174730000000
1!
1%
1-
12
#174740000000
0!
0%
b1 *
0-
02
b1 6
#174750000000
1!
1%
1-
12
#174760000000
0!
0%
b10 *
0-
02
b10 6
#174770000000
1!
1%
1-
12
#174780000000
0!
0%
b11 *
0-
02
b11 6
#174790000000
1!
1%
1-
12
15
#174800000000
0!
0%
b100 *
0-
02
b100 6
#174810000000
1!
1%
1-
12
#174820000000
0!
0%
b101 *
0-
02
b101 6
#174830000000
1!
1%
1-
12
#174840000000
0!
0%
b110 *
0-
02
b110 6
#174850000000
1!
1%
1-
12
#174860000000
0!
0%
b111 *
0-
02
b111 6
#174870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#174880000000
0!
0%
b0 *
0-
02
b0 6
#174890000000
1!
1%
1-
12
#174900000000
0!
0%
b1 *
0-
02
b1 6
#174910000000
1!
1%
1-
12
#174920000000
0!
0%
b10 *
0-
02
b10 6
#174930000000
1!
1%
1-
12
#174940000000
0!
0%
b11 *
0-
02
b11 6
#174950000000
1!
1%
1-
12
15
#174960000000
0!
0%
b100 *
0-
02
b100 6
#174970000000
1!
1%
1-
12
#174980000000
0!
0%
b101 *
0-
02
b101 6
#174990000000
1!
1%
1-
12
#175000000000
0!
0%
b110 *
0-
02
b110 6
#175010000000
1!
1%
1-
12
#175020000000
0!
0%
b111 *
0-
02
b111 6
#175030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#175040000000
0!
0%
b0 *
0-
02
b0 6
#175050000000
1!
1%
1-
12
#175060000000
0!
0%
b1 *
0-
02
b1 6
#175070000000
1!
1%
1-
12
#175080000000
0!
0%
b10 *
0-
02
b10 6
#175090000000
1!
1%
1-
12
#175100000000
0!
0%
b11 *
0-
02
b11 6
#175110000000
1!
1%
1-
12
15
#175120000000
0!
0%
b100 *
0-
02
b100 6
#175130000000
1!
1%
1-
12
#175140000000
0!
0%
b101 *
0-
02
b101 6
#175150000000
1!
1%
1-
12
#175160000000
0!
0%
b110 *
0-
02
b110 6
#175170000000
1!
1%
1-
12
#175180000000
0!
0%
b111 *
0-
02
b111 6
#175190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#175200000000
0!
0%
b0 *
0-
02
b0 6
#175210000000
1!
1%
1-
12
#175220000000
0!
0%
b1 *
0-
02
b1 6
#175230000000
1!
1%
1-
12
#175240000000
0!
0%
b10 *
0-
02
b10 6
#175250000000
1!
1%
1-
12
#175260000000
0!
0%
b11 *
0-
02
b11 6
#175270000000
1!
1%
1-
12
15
#175280000000
0!
0%
b100 *
0-
02
b100 6
#175290000000
1!
1%
1-
12
#175300000000
0!
0%
b101 *
0-
02
b101 6
#175310000000
1!
1%
1-
12
#175320000000
0!
0%
b110 *
0-
02
b110 6
#175330000000
1!
1%
1-
12
#175340000000
0!
0%
b111 *
0-
02
b111 6
#175350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#175360000000
0!
0%
b0 *
0-
02
b0 6
#175370000000
1!
1%
1-
12
#175380000000
0!
0%
b1 *
0-
02
b1 6
#175390000000
1!
1%
1-
12
#175400000000
0!
0%
b10 *
0-
02
b10 6
#175410000000
1!
1%
1-
12
#175420000000
0!
0%
b11 *
0-
02
b11 6
#175430000000
1!
1%
1-
12
15
#175440000000
0!
0%
b100 *
0-
02
b100 6
#175450000000
1!
1%
1-
12
#175460000000
0!
0%
b101 *
0-
02
b101 6
#175470000000
1!
1%
1-
12
#175480000000
0!
0%
b110 *
0-
02
b110 6
#175490000000
1!
1%
1-
12
#175500000000
0!
0%
b111 *
0-
02
b111 6
#175510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#175520000000
0!
0%
b0 *
0-
02
b0 6
#175530000000
1!
1%
1-
12
#175540000000
0!
0%
b1 *
0-
02
b1 6
#175550000000
1!
1%
1-
12
#175560000000
0!
0%
b10 *
0-
02
b10 6
#175570000000
1!
1%
1-
12
#175580000000
0!
0%
b11 *
0-
02
b11 6
#175590000000
1!
1%
1-
12
15
#175600000000
0!
0%
b100 *
0-
02
b100 6
#175610000000
1!
1%
1-
12
#175620000000
0!
0%
b101 *
0-
02
b101 6
#175630000000
1!
1%
1-
12
#175640000000
0!
0%
b110 *
0-
02
b110 6
#175650000000
1!
1%
1-
12
#175660000000
0!
0%
b111 *
0-
02
b111 6
#175670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#175680000000
0!
0%
b0 *
0-
02
b0 6
#175690000000
1!
1%
1-
12
#175700000000
0!
0%
b1 *
0-
02
b1 6
#175710000000
1!
1%
1-
12
#175720000000
0!
0%
b10 *
0-
02
b10 6
#175730000000
1!
1%
1-
12
#175740000000
0!
0%
b11 *
0-
02
b11 6
#175750000000
1!
1%
1-
12
15
#175760000000
0!
0%
b100 *
0-
02
b100 6
#175770000000
1!
1%
1-
12
#175780000000
0!
0%
b101 *
0-
02
b101 6
#175790000000
1!
1%
1-
12
#175800000000
0!
0%
b110 *
0-
02
b110 6
#175810000000
1!
1%
1-
12
#175820000000
0!
0%
b111 *
0-
02
b111 6
#175830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#175840000000
0!
0%
b0 *
0-
02
b0 6
#175850000000
1!
1%
1-
12
#175860000000
0!
0%
b1 *
0-
02
b1 6
#175870000000
1!
1%
1-
12
#175880000000
0!
0%
b10 *
0-
02
b10 6
#175890000000
1!
1%
1-
12
#175900000000
0!
0%
b11 *
0-
02
b11 6
#175910000000
1!
1%
1-
12
15
#175920000000
0!
0%
b100 *
0-
02
b100 6
#175930000000
1!
1%
1-
12
#175940000000
0!
0%
b101 *
0-
02
b101 6
#175950000000
1!
1%
1-
12
#175960000000
0!
0%
b110 *
0-
02
b110 6
#175970000000
1!
1%
1-
12
#175980000000
0!
0%
b111 *
0-
02
b111 6
#175990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#176000000000
0!
0%
b0 *
0-
02
b0 6
#176010000000
1!
1%
1-
12
#176020000000
0!
0%
b1 *
0-
02
b1 6
#176030000000
1!
1%
1-
12
#176040000000
0!
0%
b10 *
0-
02
b10 6
#176050000000
1!
1%
1-
12
#176060000000
0!
0%
b11 *
0-
02
b11 6
#176070000000
1!
1%
1-
12
15
#176080000000
0!
0%
b100 *
0-
02
b100 6
#176090000000
1!
1%
1-
12
#176100000000
0!
0%
b101 *
0-
02
b101 6
#176110000000
1!
1%
1-
12
#176120000000
0!
0%
b110 *
0-
02
b110 6
#176130000000
1!
1%
1-
12
#176140000000
0!
0%
b111 *
0-
02
b111 6
#176150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#176160000000
0!
0%
b0 *
0-
02
b0 6
#176170000000
1!
1%
1-
12
#176180000000
0!
0%
b1 *
0-
02
b1 6
#176190000000
1!
1%
1-
12
#176200000000
0!
0%
b10 *
0-
02
b10 6
#176210000000
1!
1%
1-
12
#176220000000
0!
0%
b11 *
0-
02
b11 6
#176230000000
1!
1%
1-
12
15
#176240000000
0!
0%
b100 *
0-
02
b100 6
#176250000000
1!
1%
1-
12
#176260000000
0!
0%
b101 *
0-
02
b101 6
#176270000000
1!
1%
1-
12
#176280000000
0!
0%
b110 *
0-
02
b110 6
#176290000000
1!
1%
1-
12
#176300000000
0!
0%
b111 *
0-
02
b111 6
#176310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#176320000000
0!
0%
b0 *
0-
02
b0 6
#176330000000
1!
1%
1-
12
#176340000000
0!
0%
b1 *
0-
02
b1 6
#176350000000
1!
1%
1-
12
#176360000000
0!
0%
b10 *
0-
02
b10 6
#176370000000
1!
1%
1-
12
#176380000000
0!
0%
b11 *
0-
02
b11 6
#176390000000
1!
1%
1-
12
15
#176400000000
0!
0%
b100 *
0-
02
b100 6
#176410000000
1!
1%
1-
12
#176420000000
0!
0%
b101 *
0-
02
b101 6
#176430000000
1!
1%
1-
12
#176440000000
0!
0%
b110 *
0-
02
b110 6
#176450000000
1!
1%
1-
12
#176460000000
0!
0%
b111 *
0-
02
b111 6
#176470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#176480000000
0!
0%
b0 *
0-
02
b0 6
#176490000000
1!
1%
1-
12
#176500000000
0!
0%
b1 *
0-
02
b1 6
#176510000000
1!
1%
1-
12
#176520000000
0!
0%
b10 *
0-
02
b10 6
#176530000000
1!
1%
1-
12
#176540000000
0!
0%
b11 *
0-
02
b11 6
#176550000000
1!
1%
1-
12
15
#176560000000
0!
0%
b100 *
0-
02
b100 6
#176570000000
1!
1%
1-
12
#176580000000
0!
0%
b101 *
0-
02
b101 6
#176590000000
1!
1%
1-
12
#176600000000
0!
0%
b110 *
0-
02
b110 6
#176610000000
1!
1%
1-
12
#176620000000
0!
0%
b111 *
0-
02
b111 6
#176630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#176640000000
0!
0%
b0 *
0-
02
b0 6
#176650000000
1!
1%
1-
12
#176660000000
0!
0%
b1 *
0-
02
b1 6
#176670000000
1!
1%
1-
12
#176680000000
0!
0%
b10 *
0-
02
b10 6
#176690000000
1!
1%
1-
12
#176700000000
0!
0%
b11 *
0-
02
b11 6
#176710000000
1!
1%
1-
12
15
#176720000000
0!
0%
b100 *
0-
02
b100 6
#176730000000
1!
1%
1-
12
#176740000000
0!
0%
b101 *
0-
02
b101 6
#176750000000
1!
1%
1-
12
#176760000000
0!
0%
b110 *
0-
02
b110 6
#176770000000
1!
1%
1-
12
#176780000000
0!
0%
b111 *
0-
02
b111 6
#176790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#176800000000
0!
0%
b0 *
0-
02
b0 6
#176810000000
1!
1%
1-
12
#176820000000
0!
0%
b1 *
0-
02
b1 6
#176830000000
1!
1%
1-
12
#176840000000
0!
0%
b10 *
0-
02
b10 6
#176850000000
1!
1%
1-
12
#176860000000
0!
0%
b11 *
0-
02
b11 6
#176870000000
1!
1%
1-
12
15
#176880000000
0!
0%
b100 *
0-
02
b100 6
#176890000000
1!
1%
1-
12
#176900000000
0!
0%
b101 *
0-
02
b101 6
#176910000000
1!
1%
1-
12
#176920000000
0!
0%
b110 *
0-
02
b110 6
#176930000000
1!
1%
1-
12
#176940000000
0!
0%
b111 *
0-
02
b111 6
#176950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#176960000000
0!
0%
b0 *
0-
02
b0 6
#176970000000
1!
1%
1-
12
#176980000000
0!
0%
b1 *
0-
02
b1 6
#176990000000
1!
1%
1-
12
#177000000000
0!
0%
b10 *
0-
02
b10 6
#177010000000
1!
1%
1-
12
#177020000000
0!
0%
b11 *
0-
02
b11 6
#177030000000
1!
1%
1-
12
15
#177040000000
0!
0%
b100 *
0-
02
b100 6
#177050000000
1!
1%
1-
12
#177060000000
0!
0%
b101 *
0-
02
b101 6
#177070000000
1!
1%
1-
12
#177080000000
0!
0%
b110 *
0-
02
b110 6
#177090000000
1!
1%
1-
12
#177100000000
0!
0%
b111 *
0-
02
b111 6
#177110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#177120000000
0!
0%
b0 *
0-
02
b0 6
#177130000000
1!
1%
1-
12
#177140000000
0!
0%
b1 *
0-
02
b1 6
#177150000000
1!
1%
1-
12
#177160000000
0!
0%
b10 *
0-
02
b10 6
#177170000000
1!
1%
1-
12
#177180000000
0!
0%
b11 *
0-
02
b11 6
#177190000000
1!
1%
1-
12
15
#177200000000
0!
0%
b100 *
0-
02
b100 6
#177210000000
1!
1%
1-
12
#177220000000
0!
0%
b101 *
0-
02
b101 6
#177230000000
1!
1%
1-
12
#177240000000
0!
0%
b110 *
0-
02
b110 6
#177250000000
1!
1%
1-
12
#177260000000
0!
0%
b111 *
0-
02
b111 6
#177270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#177280000000
0!
0%
b0 *
0-
02
b0 6
#177290000000
1!
1%
1-
12
#177300000000
0!
0%
b1 *
0-
02
b1 6
#177310000000
1!
1%
1-
12
#177320000000
0!
0%
b10 *
0-
02
b10 6
#177330000000
1!
1%
1-
12
#177340000000
0!
0%
b11 *
0-
02
b11 6
#177350000000
1!
1%
1-
12
15
#177360000000
0!
0%
b100 *
0-
02
b100 6
#177370000000
1!
1%
1-
12
#177380000000
0!
0%
b101 *
0-
02
b101 6
#177390000000
1!
1%
1-
12
#177400000000
0!
0%
b110 *
0-
02
b110 6
#177410000000
1!
1%
1-
12
#177420000000
0!
0%
b111 *
0-
02
b111 6
#177430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#177440000000
0!
0%
b0 *
0-
02
b0 6
#177450000000
1!
1%
1-
12
#177460000000
0!
0%
b1 *
0-
02
b1 6
#177470000000
1!
1%
1-
12
#177480000000
0!
0%
b10 *
0-
02
b10 6
#177490000000
1!
1%
1-
12
#177500000000
0!
0%
b11 *
0-
02
b11 6
#177510000000
1!
1%
1-
12
15
#177520000000
0!
0%
b100 *
0-
02
b100 6
#177530000000
1!
1%
1-
12
#177540000000
0!
0%
b101 *
0-
02
b101 6
#177550000000
1!
1%
1-
12
#177560000000
0!
0%
b110 *
0-
02
b110 6
#177570000000
1!
1%
1-
12
#177580000000
0!
0%
b111 *
0-
02
b111 6
#177590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#177600000000
0!
0%
b0 *
0-
02
b0 6
#177610000000
1!
1%
1-
12
#177620000000
0!
0%
b1 *
0-
02
b1 6
#177630000000
1!
1%
1-
12
#177640000000
0!
0%
b10 *
0-
02
b10 6
#177650000000
1!
1%
1-
12
#177660000000
0!
0%
b11 *
0-
02
b11 6
#177670000000
1!
1%
1-
12
15
#177680000000
0!
0%
b100 *
0-
02
b100 6
#177690000000
1!
1%
1-
12
#177700000000
0!
0%
b101 *
0-
02
b101 6
#177710000000
1!
1%
1-
12
#177720000000
0!
0%
b110 *
0-
02
b110 6
#177730000000
1!
1%
1-
12
#177740000000
0!
0%
b111 *
0-
02
b111 6
#177750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#177760000000
0!
0%
b0 *
0-
02
b0 6
#177770000000
1!
1%
1-
12
#177780000000
0!
0%
b1 *
0-
02
b1 6
#177790000000
1!
1%
1-
12
#177800000000
0!
0%
b10 *
0-
02
b10 6
#177810000000
1!
1%
1-
12
#177820000000
0!
0%
b11 *
0-
02
b11 6
#177830000000
1!
1%
1-
12
15
#177840000000
0!
0%
b100 *
0-
02
b100 6
#177850000000
1!
1%
1-
12
#177860000000
0!
0%
b101 *
0-
02
b101 6
#177870000000
1!
1%
1-
12
#177880000000
0!
0%
b110 *
0-
02
b110 6
#177890000000
1!
1%
1-
12
#177900000000
0!
0%
b111 *
0-
02
b111 6
#177910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#177920000000
0!
0%
b0 *
0-
02
b0 6
#177930000000
1!
1%
1-
12
#177940000000
0!
0%
b1 *
0-
02
b1 6
#177950000000
1!
1%
1-
12
#177960000000
0!
0%
b10 *
0-
02
b10 6
#177970000000
1!
1%
1-
12
#177980000000
0!
0%
b11 *
0-
02
b11 6
#177990000000
1!
1%
1-
12
15
#178000000000
0!
0%
b100 *
0-
02
b100 6
#178010000000
1!
1%
1-
12
#178020000000
0!
0%
b101 *
0-
02
b101 6
#178030000000
1!
1%
1-
12
#178040000000
0!
0%
b110 *
0-
02
b110 6
#178050000000
1!
1%
1-
12
#178060000000
0!
0%
b111 *
0-
02
b111 6
#178070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#178080000000
0!
0%
b0 *
0-
02
b0 6
#178090000000
1!
1%
1-
12
#178100000000
0!
0%
b1 *
0-
02
b1 6
#178110000000
1!
1%
1-
12
#178120000000
0!
0%
b10 *
0-
02
b10 6
#178130000000
1!
1%
1-
12
#178140000000
0!
0%
b11 *
0-
02
b11 6
#178150000000
1!
1%
1-
12
15
#178160000000
0!
0%
b100 *
0-
02
b100 6
#178170000000
1!
1%
1-
12
#178180000000
0!
0%
b101 *
0-
02
b101 6
#178190000000
1!
1%
1-
12
#178200000000
0!
0%
b110 *
0-
02
b110 6
#178210000000
1!
1%
1-
12
#178220000000
0!
0%
b111 *
0-
02
b111 6
#178230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#178240000000
0!
0%
b0 *
0-
02
b0 6
#178250000000
1!
1%
1-
12
#178260000000
0!
0%
b1 *
0-
02
b1 6
#178270000000
1!
1%
1-
12
#178280000000
0!
0%
b10 *
0-
02
b10 6
#178290000000
1!
1%
1-
12
#178300000000
0!
0%
b11 *
0-
02
b11 6
#178310000000
1!
1%
1-
12
15
#178320000000
0!
0%
b100 *
0-
02
b100 6
#178330000000
1!
1%
1-
12
#178340000000
0!
0%
b101 *
0-
02
b101 6
#178350000000
1!
1%
1-
12
#178360000000
0!
0%
b110 *
0-
02
b110 6
#178370000000
1!
1%
1-
12
#178380000000
0!
0%
b111 *
0-
02
b111 6
#178390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#178400000000
0!
0%
b0 *
0-
02
b0 6
#178410000000
1!
1%
1-
12
#178420000000
0!
0%
b1 *
0-
02
b1 6
#178430000000
1!
1%
1-
12
#178440000000
0!
0%
b10 *
0-
02
b10 6
#178450000000
1!
1%
1-
12
#178460000000
0!
0%
b11 *
0-
02
b11 6
#178470000000
1!
1%
1-
12
15
#178480000000
0!
0%
b100 *
0-
02
b100 6
#178490000000
1!
1%
1-
12
#178500000000
0!
0%
b101 *
0-
02
b101 6
#178510000000
1!
1%
1-
12
#178520000000
0!
0%
b110 *
0-
02
b110 6
#178530000000
1!
1%
1-
12
#178540000000
0!
0%
b111 *
0-
02
b111 6
#178550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#178560000000
0!
0%
b0 *
0-
02
b0 6
#178570000000
1!
1%
1-
12
#178580000000
0!
0%
b1 *
0-
02
b1 6
#178590000000
1!
1%
1-
12
#178600000000
0!
0%
b10 *
0-
02
b10 6
#178610000000
1!
1%
1-
12
#178620000000
0!
0%
b11 *
0-
02
b11 6
#178630000000
1!
1%
1-
12
15
#178640000000
0!
0%
b100 *
0-
02
b100 6
#178650000000
1!
1%
1-
12
#178660000000
0!
0%
b101 *
0-
02
b101 6
#178670000000
1!
1%
1-
12
#178680000000
0!
0%
b110 *
0-
02
b110 6
#178690000000
1!
1%
1-
12
#178700000000
0!
0%
b111 *
0-
02
b111 6
#178710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#178720000000
0!
0%
b0 *
0-
02
b0 6
#178730000000
1!
1%
1-
12
#178740000000
0!
0%
b1 *
0-
02
b1 6
#178750000000
1!
1%
1-
12
#178760000000
0!
0%
b10 *
0-
02
b10 6
#178770000000
1!
1%
1-
12
#178780000000
0!
0%
b11 *
0-
02
b11 6
#178790000000
1!
1%
1-
12
15
#178800000000
0!
0%
b100 *
0-
02
b100 6
#178810000000
1!
1%
1-
12
#178820000000
0!
0%
b101 *
0-
02
b101 6
#178830000000
1!
1%
1-
12
#178840000000
0!
0%
b110 *
0-
02
b110 6
#178850000000
1!
1%
1-
12
#178860000000
0!
0%
b111 *
0-
02
b111 6
#178870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#178880000000
0!
0%
b0 *
0-
02
b0 6
#178890000000
1!
1%
1-
12
#178900000000
0!
0%
b1 *
0-
02
b1 6
#178910000000
1!
1%
1-
12
#178920000000
0!
0%
b10 *
0-
02
b10 6
#178930000000
1!
1%
1-
12
#178940000000
0!
0%
b11 *
0-
02
b11 6
#178950000000
1!
1%
1-
12
15
#178960000000
0!
0%
b100 *
0-
02
b100 6
#178970000000
1!
1%
1-
12
#178980000000
0!
0%
b101 *
0-
02
b101 6
#178990000000
1!
1%
1-
12
#179000000000
0!
0%
b110 *
0-
02
b110 6
#179010000000
1!
1%
1-
12
#179020000000
0!
0%
b111 *
0-
02
b111 6
#179030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#179040000000
0!
0%
b0 *
0-
02
b0 6
#179050000000
1!
1%
1-
12
#179060000000
0!
0%
b1 *
0-
02
b1 6
#179070000000
1!
1%
1-
12
#179080000000
0!
0%
b10 *
0-
02
b10 6
#179090000000
1!
1%
1-
12
#179100000000
0!
0%
b11 *
0-
02
b11 6
#179110000000
1!
1%
1-
12
15
#179120000000
0!
0%
b100 *
0-
02
b100 6
#179130000000
1!
1%
1-
12
#179140000000
0!
0%
b101 *
0-
02
b101 6
#179150000000
1!
1%
1-
12
#179160000000
0!
0%
b110 *
0-
02
b110 6
#179170000000
1!
1%
1-
12
#179180000000
0!
0%
b111 *
0-
02
b111 6
#179190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#179200000000
0!
0%
b0 *
0-
02
b0 6
#179210000000
1!
1%
1-
12
#179220000000
0!
0%
b1 *
0-
02
b1 6
#179230000000
1!
1%
1-
12
#179240000000
0!
0%
b10 *
0-
02
b10 6
#179250000000
1!
1%
1-
12
#179260000000
0!
0%
b11 *
0-
02
b11 6
#179270000000
1!
1%
1-
12
15
#179280000000
0!
0%
b100 *
0-
02
b100 6
#179290000000
1!
1%
1-
12
#179300000000
0!
0%
b101 *
0-
02
b101 6
#179310000000
1!
1%
1-
12
#179320000000
0!
0%
b110 *
0-
02
b110 6
#179330000000
1!
1%
1-
12
#179340000000
0!
0%
b111 *
0-
02
b111 6
#179350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#179360000000
0!
0%
b0 *
0-
02
b0 6
#179370000000
1!
1%
1-
12
#179380000000
0!
0%
b1 *
0-
02
b1 6
#179390000000
1!
1%
1-
12
#179400000000
0!
0%
b10 *
0-
02
b10 6
#179410000000
1!
1%
1-
12
#179420000000
0!
0%
b11 *
0-
02
b11 6
#179430000000
1!
1%
1-
12
15
#179440000000
0!
0%
b100 *
0-
02
b100 6
#179450000000
1!
1%
1-
12
#179460000000
0!
0%
b101 *
0-
02
b101 6
#179470000000
1!
1%
1-
12
#179480000000
0!
0%
b110 *
0-
02
b110 6
#179490000000
1!
1%
1-
12
#179500000000
0!
0%
b111 *
0-
02
b111 6
#179510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#179520000000
0!
0%
b0 *
0-
02
b0 6
#179530000000
1!
1%
1-
12
#179540000000
0!
0%
b1 *
0-
02
b1 6
#179550000000
1!
1%
1-
12
#179560000000
0!
0%
b10 *
0-
02
b10 6
#179570000000
1!
1%
1-
12
#179580000000
0!
0%
b11 *
0-
02
b11 6
#179590000000
1!
1%
1-
12
15
#179600000000
0!
0%
b100 *
0-
02
b100 6
#179610000000
1!
1%
1-
12
#179620000000
0!
0%
b101 *
0-
02
b101 6
#179630000000
1!
1%
1-
12
#179640000000
0!
0%
b110 *
0-
02
b110 6
#179650000000
1!
1%
1-
12
#179660000000
0!
0%
b111 *
0-
02
b111 6
#179670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#179680000000
0!
0%
b0 *
0-
02
b0 6
#179690000000
1!
1%
1-
12
#179700000000
0!
0%
b1 *
0-
02
b1 6
#179710000000
1!
1%
1-
12
#179720000000
0!
0%
b10 *
0-
02
b10 6
#179730000000
1!
1%
1-
12
#179740000000
0!
0%
b11 *
0-
02
b11 6
#179750000000
1!
1%
1-
12
15
#179760000000
0!
0%
b100 *
0-
02
b100 6
#179770000000
1!
1%
1-
12
#179780000000
0!
0%
b101 *
0-
02
b101 6
#179790000000
1!
1%
1-
12
#179800000000
0!
0%
b110 *
0-
02
b110 6
#179810000000
1!
1%
1-
12
#179820000000
0!
0%
b111 *
0-
02
b111 6
#179830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#179840000000
0!
0%
b0 *
0-
02
b0 6
#179850000000
1!
1%
1-
12
#179860000000
0!
0%
b1 *
0-
02
b1 6
#179870000000
1!
1%
1-
12
#179880000000
0!
0%
b10 *
0-
02
b10 6
#179890000000
1!
1%
1-
12
#179900000000
0!
0%
b11 *
0-
02
b11 6
#179910000000
1!
1%
1-
12
15
#179920000000
0!
0%
b100 *
0-
02
b100 6
#179930000000
1!
1%
1-
12
#179940000000
0!
0%
b101 *
0-
02
b101 6
#179950000000
1!
1%
1-
12
#179960000000
0!
0%
b110 *
0-
02
b110 6
#179970000000
1!
1%
1-
12
#179980000000
0!
0%
b111 *
0-
02
b111 6
#179990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#180000000000
0!
0%
b0 *
0-
02
b0 6
#180010000000
1!
1%
1-
12
#180020000000
0!
0%
b1 *
0-
02
b1 6
#180030000000
1!
1%
1-
12
#180040000000
0!
0%
b10 *
0-
02
b10 6
#180050000000
1!
1%
1-
12
#180060000000
0!
0%
b11 *
0-
02
b11 6
#180070000000
1!
1%
1-
12
15
#180080000000
0!
0%
b100 *
0-
02
b100 6
#180090000000
1!
1%
1-
12
#180100000000
0!
0%
b101 *
0-
02
b101 6
#180110000000
1!
1%
1-
12
#180120000000
0!
0%
b110 *
0-
02
b110 6
#180130000000
1!
1%
1-
12
#180140000000
0!
0%
b111 *
0-
02
b111 6
#180150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#180160000000
0!
0%
b0 *
0-
02
b0 6
#180170000000
1!
1%
1-
12
#180180000000
0!
0%
b1 *
0-
02
b1 6
#180190000000
1!
1%
1-
12
#180200000000
0!
0%
b10 *
0-
02
b10 6
#180210000000
1!
1%
1-
12
#180220000000
0!
0%
b11 *
0-
02
b11 6
#180230000000
1!
1%
1-
12
15
#180240000000
0!
0%
b100 *
0-
02
b100 6
#180250000000
1!
1%
1-
12
#180260000000
0!
0%
b101 *
0-
02
b101 6
#180270000000
1!
1%
1-
12
#180280000000
0!
0%
b110 *
0-
02
b110 6
#180290000000
1!
1%
1-
12
#180300000000
0!
0%
b111 *
0-
02
b111 6
#180310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#180320000000
0!
0%
b0 *
0-
02
b0 6
#180330000000
1!
1%
1-
12
#180340000000
0!
0%
b1 *
0-
02
b1 6
#180350000000
1!
1%
1-
12
#180360000000
0!
0%
b10 *
0-
02
b10 6
#180370000000
1!
1%
1-
12
#180380000000
0!
0%
b11 *
0-
02
b11 6
#180390000000
1!
1%
1-
12
15
#180400000000
0!
0%
b100 *
0-
02
b100 6
#180410000000
1!
1%
1-
12
#180420000000
0!
0%
b101 *
0-
02
b101 6
#180430000000
1!
1%
1-
12
#180440000000
0!
0%
b110 *
0-
02
b110 6
#180450000000
1!
1%
1-
12
#180460000000
0!
0%
b111 *
0-
02
b111 6
#180470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#180480000000
0!
0%
b0 *
0-
02
b0 6
#180490000000
1!
1%
1-
12
#180500000000
0!
0%
b1 *
0-
02
b1 6
#180510000000
1!
1%
1-
12
#180520000000
0!
0%
b10 *
0-
02
b10 6
#180530000000
1!
1%
1-
12
#180540000000
0!
0%
b11 *
0-
02
b11 6
#180550000000
1!
1%
1-
12
15
#180560000000
0!
0%
b100 *
0-
02
b100 6
#180570000000
1!
1%
1-
12
#180580000000
0!
0%
b101 *
0-
02
b101 6
#180590000000
1!
1%
1-
12
#180600000000
0!
0%
b110 *
0-
02
b110 6
#180610000000
1!
1%
1-
12
#180620000000
0!
0%
b111 *
0-
02
b111 6
#180630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#180640000000
0!
0%
b0 *
0-
02
b0 6
#180650000000
1!
1%
1-
12
#180660000000
0!
0%
b1 *
0-
02
b1 6
#180670000000
1!
1%
1-
12
#180680000000
0!
0%
b10 *
0-
02
b10 6
#180690000000
1!
1%
1-
12
#180700000000
0!
0%
b11 *
0-
02
b11 6
#180710000000
1!
1%
1-
12
15
#180720000000
0!
0%
b100 *
0-
02
b100 6
#180730000000
1!
1%
1-
12
#180740000000
0!
0%
b101 *
0-
02
b101 6
#180750000000
1!
1%
1-
12
#180760000000
0!
0%
b110 *
0-
02
b110 6
#180770000000
1!
1%
1-
12
#180780000000
0!
0%
b111 *
0-
02
b111 6
#180790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#180800000000
0!
0%
b0 *
0-
02
b0 6
#180810000000
1!
1%
1-
12
#180820000000
0!
0%
b1 *
0-
02
b1 6
#180830000000
1!
1%
1-
12
#180840000000
0!
0%
b10 *
0-
02
b10 6
#180850000000
1!
1%
1-
12
#180860000000
0!
0%
b11 *
0-
02
b11 6
#180870000000
1!
1%
1-
12
15
#180880000000
0!
0%
b100 *
0-
02
b100 6
#180890000000
1!
1%
1-
12
#180900000000
0!
0%
b101 *
0-
02
b101 6
#180910000000
1!
1%
1-
12
#180920000000
0!
0%
b110 *
0-
02
b110 6
#180930000000
1!
1%
1-
12
#180940000000
0!
0%
b111 *
0-
02
b111 6
#180950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#180960000000
0!
0%
b0 *
0-
02
b0 6
#180970000000
1!
1%
1-
12
#180980000000
0!
0%
b1 *
0-
02
b1 6
#180990000000
1!
1%
1-
12
#181000000000
0!
0%
b10 *
0-
02
b10 6
#181010000000
1!
1%
1-
12
#181020000000
0!
0%
b11 *
0-
02
b11 6
#181030000000
1!
1%
1-
12
15
#181040000000
0!
0%
b100 *
0-
02
b100 6
#181050000000
1!
1%
1-
12
#181060000000
0!
0%
b101 *
0-
02
b101 6
#181070000000
1!
1%
1-
12
#181080000000
0!
0%
b110 *
0-
02
b110 6
#181090000000
1!
1%
1-
12
#181100000000
0!
0%
b111 *
0-
02
b111 6
#181110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#181120000000
0!
0%
b0 *
0-
02
b0 6
#181130000000
1!
1%
1-
12
#181140000000
0!
0%
b1 *
0-
02
b1 6
#181150000000
1!
1%
1-
12
#181160000000
0!
0%
b10 *
0-
02
b10 6
#181170000000
1!
1%
1-
12
#181180000000
0!
0%
b11 *
0-
02
b11 6
#181190000000
1!
1%
1-
12
15
#181200000000
0!
0%
b100 *
0-
02
b100 6
#181210000000
1!
1%
1-
12
#181220000000
0!
0%
b101 *
0-
02
b101 6
#181230000000
1!
1%
1-
12
#181240000000
0!
0%
b110 *
0-
02
b110 6
#181250000000
1!
1%
1-
12
#181260000000
0!
0%
b111 *
0-
02
b111 6
#181270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#181280000000
0!
0%
b0 *
0-
02
b0 6
#181290000000
1!
1%
1-
12
#181300000000
0!
0%
b1 *
0-
02
b1 6
#181310000000
1!
1%
1-
12
#181320000000
0!
0%
b10 *
0-
02
b10 6
#181330000000
1!
1%
1-
12
#181340000000
0!
0%
b11 *
0-
02
b11 6
#181350000000
1!
1%
1-
12
15
#181360000000
0!
0%
b100 *
0-
02
b100 6
#181370000000
1!
1%
1-
12
#181380000000
0!
0%
b101 *
0-
02
b101 6
#181390000000
1!
1%
1-
12
#181400000000
0!
0%
b110 *
0-
02
b110 6
#181410000000
1!
1%
1-
12
#181420000000
0!
0%
b111 *
0-
02
b111 6
#181430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#181440000000
0!
0%
b0 *
0-
02
b0 6
#181450000000
1!
1%
1-
12
#181460000000
0!
0%
b1 *
0-
02
b1 6
#181470000000
1!
1%
1-
12
#181480000000
0!
0%
b10 *
0-
02
b10 6
#181490000000
1!
1%
1-
12
#181500000000
0!
0%
b11 *
0-
02
b11 6
#181510000000
1!
1%
1-
12
15
#181520000000
0!
0%
b100 *
0-
02
b100 6
#181530000000
1!
1%
1-
12
#181540000000
0!
0%
b101 *
0-
02
b101 6
#181550000000
1!
1%
1-
12
#181560000000
0!
0%
b110 *
0-
02
b110 6
#181570000000
1!
1%
1-
12
#181580000000
0!
0%
b111 *
0-
02
b111 6
#181590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#181600000000
0!
0%
b0 *
0-
02
b0 6
#181610000000
1!
1%
1-
12
#181620000000
0!
0%
b1 *
0-
02
b1 6
#181630000000
1!
1%
1-
12
#181640000000
0!
0%
b10 *
0-
02
b10 6
#181650000000
1!
1%
1-
12
#181660000000
0!
0%
b11 *
0-
02
b11 6
#181670000000
1!
1%
1-
12
15
#181680000000
0!
0%
b100 *
0-
02
b100 6
#181690000000
1!
1%
1-
12
#181700000000
0!
0%
b101 *
0-
02
b101 6
#181710000000
1!
1%
1-
12
#181720000000
0!
0%
b110 *
0-
02
b110 6
#181730000000
1!
1%
1-
12
#181740000000
0!
0%
b111 *
0-
02
b111 6
#181750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#181760000000
0!
0%
b0 *
0-
02
b0 6
#181770000000
1!
1%
1-
12
#181780000000
0!
0%
b1 *
0-
02
b1 6
#181790000000
1!
1%
1-
12
#181800000000
0!
0%
b10 *
0-
02
b10 6
#181810000000
1!
1%
1-
12
#181820000000
0!
0%
b11 *
0-
02
b11 6
#181830000000
1!
1%
1-
12
15
#181840000000
0!
0%
b100 *
0-
02
b100 6
#181850000000
1!
1%
1-
12
#181860000000
0!
0%
b101 *
0-
02
b101 6
#181870000000
1!
1%
1-
12
#181880000000
0!
0%
b110 *
0-
02
b110 6
#181890000000
1!
1%
1-
12
#181900000000
0!
0%
b111 *
0-
02
b111 6
#181910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#181920000000
0!
0%
b0 *
0-
02
b0 6
#181930000000
1!
1%
1-
12
#181940000000
0!
0%
b1 *
0-
02
b1 6
#181950000000
1!
1%
1-
12
#181960000000
0!
0%
b10 *
0-
02
b10 6
#181970000000
1!
1%
1-
12
#181980000000
0!
0%
b11 *
0-
02
b11 6
#181990000000
1!
1%
1-
12
15
#182000000000
0!
0%
b100 *
0-
02
b100 6
#182010000000
1!
1%
1-
12
#182020000000
0!
0%
b101 *
0-
02
b101 6
#182030000000
1!
1%
1-
12
#182040000000
0!
0%
b110 *
0-
02
b110 6
#182050000000
1!
1%
1-
12
#182060000000
0!
0%
b111 *
0-
02
b111 6
#182070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#182080000000
0!
0%
b0 *
0-
02
b0 6
#182090000000
1!
1%
1-
12
#182100000000
0!
0%
b1 *
0-
02
b1 6
#182110000000
1!
1%
1-
12
#182120000000
0!
0%
b10 *
0-
02
b10 6
#182130000000
1!
1%
1-
12
#182140000000
0!
0%
b11 *
0-
02
b11 6
#182150000000
1!
1%
1-
12
15
#182160000000
0!
0%
b100 *
0-
02
b100 6
#182170000000
1!
1%
1-
12
#182180000000
0!
0%
b101 *
0-
02
b101 6
#182190000000
1!
1%
1-
12
#182200000000
0!
0%
b110 *
0-
02
b110 6
#182210000000
1!
1%
1-
12
#182220000000
0!
0%
b111 *
0-
02
b111 6
#182230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#182240000000
0!
0%
b0 *
0-
02
b0 6
#182250000000
1!
1%
1-
12
#182260000000
0!
0%
b1 *
0-
02
b1 6
#182270000000
1!
1%
1-
12
#182280000000
0!
0%
b10 *
0-
02
b10 6
#182290000000
1!
1%
1-
12
#182300000000
0!
0%
b11 *
0-
02
b11 6
#182310000000
1!
1%
1-
12
15
#182320000000
0!
0%
b100 *
0-
02
b100 6
#182330000000
1!
1%
1-
12
#182340000000
0!
0%
b101 *
0-
02
b101 6
#182350000000
1!
1%
1-
12
#182360000000
0!
0%
b110 *
0-
02
b110 6
#182370000000
1!
1%
1-
12
#182380000000
0!
0%
b111 *
0-
02
b111 6
#182390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#182400000000
0!
0%
b0 *
0-
02
b0 6
#182410000000
1!
1%
1-
12
#182420000000
0!
0%
b1 *
0-
02
b1 6
#182430000000
1!
1%
1-
12
#182440000000
0!
0%
b10 *
0-
02
b10 6
#182450000000
1!
1%
1-
12
#182460000000
0!
0%
b11 *
0-
02
b11 6
#182470000000
1!
1%
1-
12
15
#182480000000
0!
0%
b100 *
0-
02
b100 6
#182490000000
1!
1%
1-
12
#182500000000
0!
0%
b101 *
0-
02
b101 6
#182510000000
1!
1%
1-
12
#182520000000
0!
0%
b110 *
0-
02
b110 6
#182530000000
1!
1%
1-
12
#182540000000
0!
0%
b111 *
0-
02
b111 6
#182550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#182560000000
0!
0%
b0 *
0-
02
b0 6
#182570000000
1!
1%
1-
12
#182580000000
0!
0%
b1 *
0-
02
b1 6
#182590000000
1!
1%
1-
12
#182600000000
0!
0%
b10 *
0-
02
b10 6
#182610000000
1!
1%
1-
12
#182620000000
0!
0%
b11 *
0-
02
b11 6
#182630000000
1!
1%
1-
12
15
#182640000000
0!
0%
b100 *
0-
02
b100 6
#182650000000
1!
1%
1-
12
#182660000000
0!
0%
b101 *
0-
02
b101 6
#182670000000
1!
1%
1-
12
#182680000000
0!
0%
b110 *
0-
02
b110 6
#182690000000
1!
1%
1-
12
#182700000000
0!
0%
b111 *
0-
02
b111 6
#182710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#182720000000
0!
0%
b0 *
0-
02
b0 6
#182730000000
1!
1%
1-
12
#182740000000
0!
0%
b1 *
0-
02
b1 6
#182750000000
1!
1%
1-
12
#182760000000
0!
0%
b10 *
0-
02
b10 6
#182770000000
1!
1%
1-
12
#182780000000
0!
0%
b11 *
0-
02
b11 6
#182790000000
1!
1%
1-
12
15
#182800000000
0!
0%
b100 *
0-
02
b100 6
#182810000000
1!
1%
1-
12
#182820000000
0!
0%
b101 *
0-
02
b101 6
#182830000000
1!
1%
1-
12
#182840000000
0!
0%
b110 *
0-
02
b110 6
#182850000000
1!
1%
1-
12
#182860000000
0!
0%
b111 *
0-
02
b111 6
#182870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#182880000000
0!
0%
b0 *
0-
02
b0 6
#182890000000
1!
1%
1-
12
#182900000000
0!
0%
b1 *
0-
02
b1 6
#182910000000
1!
1%
1-
12
#182920000000
0!
0%
b10 *
0-
02
b10 6
#182930000000
1!
1%
1-
12
#182940000000
0!
0%
b11 *
0-
02
b11 6
#182950000000
1!
1%
1-
12
15
#182960000000
0!
0%
b100 *
0-
02
b100 6
#182970000000
1!
1%
1-
12
#182980000000
0!
0%
b101 *
0-
02
b101 6
#182990000000
1!
1%
1-
12
#183000000000
0!
0%
b110 *
0-
02
b110 6
#183010000000
1!
1%
1-
12
#183020000000
0!
0%
b111 *
0-
02
b111 6
#183030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#183040000000
0!
0%
b0 *
0-
02
b0 6
#183050000000
1!
1%
1-
12
#183060000000
0!
0%
b1 *
0-
02
b1 6
#183070000000
1!
1%
1-
12
#183080000000
0!
0%
b10 *
0-
02
b10 6
#183090000000
1!
1%
1-
12
#183100000000
0!
0%
b11 *
0-
02
b11 6
#183110000000
1!
1%
1-
12
15
#183120000000
0!
0%
b100 *
0-
02
b100 6
#183130000000
1!
1%
1-
12
#183140000000
0!
0%
b101 *
0-
02
b101 6
#183150000000
1!
1%
1-
12
#183160000000
0!
0%
b110 *
0-
02
b110 6
#183170000000
1!
1%
1-
12
#183180000000
0!
0%
b111 *
0-
02
b111 6
#183190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#183200000000
0!
0%
b0 *
0-
02
b0 6
#183210000000
1!
1%
1-
12
#183220000000
0!
0%
b1 *
0-
02
b1 6
#183230000000
1!
1%
1-
12
#183240000000
0!
0%
b10 *
0-
02
b10 6
#183250000000
1!
1%
1-
12
#183260000000
0!
0%
b11 *
0-
02
b11 6
#183270000000
1!
1%
1-
12
15
#183280000000
0!
0%
b100 *
0-
02
b100 6
#183290000000
1!
1%
1-
12
#183300000000
0!
0%
b101 *
0-
02
b101 6
#183310000000
1!
1%
1-
12
#183320000000
0!
0%
b110 *
0-
02
b110 6
#183330000000
1!
1%
1-
12
#183340000000
0!
0%
b111 *
0-
02
b111 6
#183350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#183360000000
0!
0%
b0 *
0-
02
b0 6
#183370000000
1!
1%
1-
12
#183380000000
0!
0%
b1 *
0-
02
b1 6
#183390000000
1!
1%
1-
12
#183400000000
0!
0%
b10 *
0-
02
b10 6
#183410000000
1!
1%
1-
12
#183420000000
0!
0%
b11 *
0-
02
b11 6
#183430000000
1!
1%
1-
12
15
#183440000000
0!
0%
b100 *
0-
02
b100 6
#183450000000
1!
1%
1-
12
#183460000000
0!
0%
b101 *
0-
02
b101 6
#183470000000
1!
1%
1-
12
#183480000000
0!
0%
b110 *
0-
02
b110 6
#183490000000
1!
1%
1-
12
#183500000000
0!
0%
b111 *
0-
02
b111 6
#183510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#183520000000
0!
0%
b0 *
0-
02
b0 6
#183530000000
1!
1%
1-
12
#183540000000
0!
0%
b1 *
0-
02
b1 6
#183550000000
1!
1%
1-
12
#183560000000
0!
0%
b10 *
0-
02
b10 6
#183570000000
1!
1%
1-
12
#183580000000
0!
0%
b11 *
0-
02
b11 6
#183590000000
1!
1%
1-
12
15
#183600000000
0!
0%
b100 *
0-
02
b100 6
#183610000000
1!
1%
1-
12
#183620000000
0!
0%
b101 *
0-
02
b101 6
#183630000000
1!
1%
1-
12
#183640000000
0!
0%
b110 *
0-
02
b110 6
#183650000000
1!
1%
1-
12
#183660000000
0!
0%
b111 *
0-
02
b111 6
#183670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#183680000000
0!
0%
b0 *
0-
02
b0 6
#183690000000
1!
1%
1-
12
#183700000000
0!
0%
b1 *
0-
02
b1 6
#183710000000
1!
1%
1-
12
#183720000000
0!
0%
b10 *
0-
02
b10 6
#183730000000
1!
1%
1-
12
#183740000000
0!
0%
b11 *
0-
02
b11 6
#183750000000
1!
1%
1-
12
15
#183760000000
0!
0%
b100 *
0-
02
b100 6
#183770000000
1!
1%
1-
12
#183780000000
0!
0%
b101 *
0-
02
b101 6
#183790000000
1!
1%
1-
12
#183800000000
0!
0%
b110 *
0-
02
b110 6
#183810000000
1!
1%
1-
12
#183820000000
0!
0%
b111 *
0-
02
b111 6
#183830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#183840000000
0!
0%
b0 *
0-
02
b0 6
#183850000000
1!
1%
1-
12
#183860000000
0!
0%
b1 *
0-
02
b1 6
#183870000000
1!
1%
1-
12
#183880000000
0!
0%
b10 *
0-
02
b10 6
#183890000000
1!
1%
1-
12
#183900000000
0!
0%
b11 *
0-
02
b11 6
#183910000000
1!
1%
1-
12
15
#183920000000
0!
0%
b100 *
0-
02
b100 6
#183930000000
1!
1%
1-
12
#183940000000
0!
0%
b101 *
0-
02
b101 6
#183950000000
1!
1%
1-
12
#183960000000
0!
0%
b110 *
0-
02
b110 6
#183970000000
1!
1%
1-
12
#183980000000
0!
0%
b111 *
0-
02
b111 6
#183990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#184000000000
0!
0%
b0 *
0-
02
b0 6
#184010000000
1!
1%
1-
12
#184020000000
0!
0%
b1 *
0-
02
b1 6
#184030000000
1!
1%
1-
12
#184040000000
0!
0%
b10 *
0-
02
b10 6
#184050000000
1!
1%
1-
12
#184060000000
0!
0%
b11 *
0-
02
b11 6
#184070000000
1!
1%
1-
12
15
#184080000000
0!
0%
b100 *
0-
02
b100 6
#184090000000
1!
1%
1-
12
#184100000000
0!
0%
b101 *
0-
02
b101 6
#184110000000
1!
1%
1-
12
#184120000000
0!
0%
b110 *
0-
02
b110 6
#184130000000
1!
1%
1-
12
#184140000000
0!
0%
b111 *
0-
02
b111 6
#184150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#184160000000
0!
0%
b0 *
0-
02
b0 6
#184170000000
1!
1%
1-
12
#184180000000
0!
0%
b1 *
0-
02
b1 6
#184190000000
1!
1%
1-
12
#184200000000
0!
0%
b10 *
0-
02
b10 6
#184210000000
1!
1%
1-
12
#184220000000
0!
0%
b11 *
0-
02
b11 6
#184230000000
1!
1%
1-
12
15
#184240000000
0!
0%
b100 *
0-
02
b100 6
#184250000000
1!
1%
1-
12
#184260000000
0!
0%
b101 *
0-
02
b101 6
#184270000000
1!
1%
1-
12
#184280000000
0!
0%
b110 *
0-
02
b110 6
#184290000000
1!
1%
1-
12
#184300000000
0!
0%
b111 *
0-
02
b111 6
#184310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#184320000000
0!
0%
b0 *
0-
02
b0 6
#184330000000
1!
1%
1-
12
#184340000000
0!
0%
b1 *
0-
02
b1 6
#184350000000
1!
1%
1-
12
#184360000000
0!
0%
b10 *
0-
02
b10 6
#184370000000
1!
1%
1-
12
#184380000000
0!
0%
b11 *
0-
02
b11 6
#184390000000
1!
1%
1-
12
15
#184400000000
0!
0%
b100 *
0-
02
b100 6
#184410000000
1!
1%
1-
12
#184420000000
0!
0%
b101 *
0-
02
b101 6
#184430000000
1!
1%
1-
12
#184440000000
0!
0%
b110 *
0-
02
b110 6
#184450000000
1!
1%
1-
12
#184460000000
0!
0%
b111 *
0-
02
b111 6
#184470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#184480000000
0!
0%
b0 *
0-
02
b0 6
#184490000000
1!
1%
1-
12
#184500000000
0!
0%
b1 *
0-
02
b1 6
#184510000000
1!
1%
1-
12
#184520000000
0!
0%
b10 *
0-
02
b10 6
#184530000000
1!
1%
1-
12
#184540000000
0!
0%
b11 *
0-
02
b11 6
#184550000000
1!
1%
1-
12
15
#184560000000
0!
0%
b100 *
0-
02
b100 6
#184570000000
1!
1%
1-
12
#184580000000
0!
0%
b101 *
0-
02
b101 6
#184590000000
1!
1%
1-
12
#184600000000
0!
0%
b110 *
0-
02
b110 6
#184610000000
1!
1%
1-
12
#184620000000
0!
0%
b111 *
0-
02
b111 6
#184630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#184640000000
0!
0%
b0 *
0-
02
b0 6
#184650000000
1!
1%
1-
12
#184660000000
0!
0%
b1 *
0-
02
b1 6
#184670000000
1!
1%
1-
12
#184680000000
0!
0%
b10 *
0-
02
b10 6
#184690000000
1!
1%
1-
12
#184700000000
0!
0%
b11 *
0-
02
b11 6
#184710000000
1!
1%
1-
12
15
#184720000000
0!
0%
b100 *
0-
02
b100 6
#184730000000
1!
1%
1-
12
#184740000000
0!
0%
b101 *
0-
02
b101 6
#184750000000
1!
1%
1-
12
#184760000000
0!
0%
b110 *
0-
02
b110 6
#184770000000
1!
1%
1-
12
#184780000000
0!
0%
b111 *
0-
02
b111 6
#184790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#184800000000
0!
0%
b0 *
0-
02
b0 6
#184810000000
1!
1%
1-
12
#184820000000
0!
0%
b1 *
0-
02
b1 6
#184830000000
1!
1%
1-
12
#184840000000
0!
0%
b10 *
0-
02
b10 6
#184850000000
1!
1%
1-
12
#184860000000
0!
0%
b11 *
0-
02
b11 6
#184870000000
1!
1%
1-
12
15
#184880000000
0!
0%
b100 *
0-
02
b100 6
#184890000000
1!
1%
1-
12
#184900000000
0!
0%
b101 *
0-
02
b101 6
#184910000000
1!
1%
1-
12
#184920000000
0!
0%
b110 *
0-
02
b110 6
#184930000000
1!
1%
1-
12
#184940000000
0!
0%
b111 *
0-
02
b111 6
#184950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#184960000000
0!
0%
b0 *
0-
02
b0 6
#184970000000
1!
1%
1-
12
#184980000000
0!
0%
b1 *
0-
02
b1 6
#184990000000
1!
1%
1-
12
#185000000000
0!
0%
b10 *
0-
02
b10 6
#185010000000
1!
1%
1-
12
#185020000000
0!
0%
b11 *
0-
02
b11 6
#185030000000
1!
1%
1-
12
15
#185040000000
0!
0%
b100 *
0-
02
b100 6
#185050000000
1!
1%
1-
12
#185060000000
0!
0%
b101 *
0-
02
b101 6
#185070000000
1!
1%
1-
12
#185080000000
0!
0%
b110 *
0-
02
b110 6
#185090000000
1!
1%
1-
12
#185100000000
0!
0%
b111 *
0-
02
b111 6
#185110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#185120000000
0!
0%
b0 *
0-
02
b0 6
#185130000000
1!
1%
1-
12
#185140000000
0!
0%
b1 *
0-
02
b1 6
#185150000000
1!
1%
1-
12
#185160000000
0!
0%
b10 *
0-
02
b10 6
#185170000000
1!
1%
1-
12
#185180000000
0!
0%
b11 *
0-
02
b11 6
#185190000000
1!
1%
1-
12
15
#185200000000
0!
0%
b100 *
0-
02
b100 6
#185210000000
1!
1%
1-
12
#185220000000
0!
0%
b101 *
0-
02
b101 6
#185230000000
1!
1%
1-
12
#185240000000
0!
0%
b110 *
0-
02
b110 6
#185250000000
1!
1%
1-
12
#185260000000
0!
0%
b111 *
0-
02
b111 6
#185270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#185280000000
0!
0%
b0 *
0-
02
b0 6
#185290000000
1!
1%
1-
12
#185300000000
0!
0%
b1 *
0-
02
b1 6
#185310000000
1!
1%
1-
12
#185320000000
0!
0%
b10 *
0-
02
b10 6
#185330000000
1!
1%
1-
12
#185340000000
0!
0%
b11 *
0-
02
b11 6
#185350000000
1!
1%
1-
12
15
#185360000000
0!
0%
b100 *
0-
02
b100 6
#185370000000
1!
1%
1-
12
#185380000000
0!
0%
b101 *
0-
02
b101 6
#185390000000
1!
1%
1-
12
#185400000000
0!
0%
b110 *
0-
02
b110 6
#185410000000
1!
1%
1-
12
#185420000000
0!
0%
b111 *
0-
02
b111 6
#185430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#185440000000
0!
0%
b0 *
0-
02
b0 6
#185450000000
1!
1%
1-
12
#185460000000
0!
0%
b1 *
0-
02
b1 6
#185470000000
1!
1%
1-
12
#185480000000
0!
0%
b10 *
0-
02
b10 6
#185490000000
1!
1%
1-
12
#185500000000
0!
0%
b11 *
0-
02
b11 6
#185510000000
1!
1%
1-
12
15
#185520000000
0!
0%
b100 *
0-
02
b100 6
#185530000000
1!
1%
1-
12
#185540000000
0!
0%
b101 *
0-
02
b101 6
#185550000000
1!
1%
1-
12
#185560000000
0!
0%
b110 *
0-
02
b110 6
#185570000000
1!
1%
1-
12
#185580000000
0!
0%
b111 *
0-
02
b111 6
#185590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#185600000000
0!
0%
b0 *
0-
02
b0 6
#185610000000
1!
1%
1-
12
#185620000000
0!
0%
b1 *
0-
02
b1 6
#185630000000
1!
1%
1-
12
#185640000000
0!
0%
b10 *
0-
02
b10 6
#185650000000
1!
1%
1-
12
#185660000000
0!
0%
b11 *
0-
02
b11 6
#185670000000
1!
1%
1-
12
15
#185680000000
0!
0%
b100 *
0-
02
b100 6
#185690000000
1!
1%
1-
12
#185700000000
0!
0%
b101 *
0-
02
b101 6
#185710000000
1!
1%
1-
12
#185720000000
0!
0%
b110 *
0-
02
b110 6
#185730000000
1!
1%
1-
12
#185740000000
0!
0%
b111 *
0-
02
b111 6
#185750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#185760000000
0!
0%
b0 *
0-
02
b0 6
#185770000000
1!
1%
1-
12
#185780000000
0!
0%
b1 *
0-
02
b1 6
#185790000000
1!
1%
1-
12
#185800000000
0!
0%
b10 *
0-
02
b10 6
#185810000000
1!
1%
1-
12
#185820000000
0!
0%
b11 *
0-
02
b11 6
#185830000000
1!
1%
1-
12
15
#185840000000
0!
0%
b100 *
0-
02
b100 6
#185850000000
1!
1%
1-
12
#185860000000
0!
0%
b101 *
0-
02
b101 6
#185870000000
1!
1%
1-
12
#185880000000
0!
0%
b110 *
0-
02
b110 6
#185890000000
1!
1%
1-
12
#185900000000
0!
0%
b111 *
0-
02
b111 6
#185910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#185920000000
0!
0%
b0 *
0-
02
b0 6
#185930000000
1!
1%
1-
12
#185940000000
0!
0%
b1 *
0-
02
b1 6
#185950000000
1!
1%
1-
12
#185960000000
0!
0%
b10 *
0-
02
b10 6
#185970000000
1!
1%
1-
12
#185980000000
0!
0%
b11 *
0-
02
b11 6
#185990000000
1!
1%
1-
12
15
#186000000000
0!
0%
b100 *
0-
02
b100 6
#186010000000
1!
1%
1-
12
#186020000000
0!
0%
b101 *
0-
02
b101 6
#186030000000
1!
1%
1-
12
#186040000000
0!
0%
b110 *
0-
02
b110 6
#186050000000
1!
1%
1-
12
#186060000000
0!
0%
b111 *
0-
02
b111 6
#186070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#186080000000
0!
0%
b0 *
0-
02
b0 6
#186090000000
1!
1%
1-
12
#186100000000
0!
0%
b1 *
0-
02
b1 6
#186110000000
1!
1%
1-
12
#186120000000
0!
0%
b10 *
0-
02
b10 6
#186130000000
1!
1%
1-
12
#186140000000
0!
0%
b11 *
0-
02
b11 6
#186150000000
1!
1%
1-
12
15
#186160000000
0!
0%
b100 *
0-
02
b100 6
#186170000000
1!
1%
1-
12
#186180000000
0!
0%
b101 *
0-
02
b101 6
#186190000000
1!
1%
1-
12
#186200000000
0!
0%
b110 *
0-
02
b110 6
#186210000000
1!
1%
1-
12
#186220000000
0!
0%
b111 *
0-
02
b111 6
#186230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#186240000000
0!
0%
b0 *
0-
02
b0 6
#186250000000
1!
1%
1-
12
#186260000000
0!
0%
b1 *
0-
02
b1 6
#186270000000
1!
1%
1-
12
#186280000000
0!
0%
b10 *
0-
02
b10 6
#186290000000
1!
1%
1-
12
#186300000000
0!
0%
b11 *
0-
02
b11 6
#186310000000
1!
1%
1-
12
15
#186320000000
0!
0%
b100 *
0-
02
b100 6
#186330000000
1!
1%
1-
12
#186340000000
0!
0%
b101 *
0-
02
b101 6
#186350000000
1!
1%
1-
12
#186360000000
0!
0%
b110 *
0-
02
b110 6
#186370000000
1!
1%
1-
12
#186380000000
0!
0%
b111 *
0-
02
b111 6
#186390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#186400000000
0!
0%
b0 *
0-
02
b0 6
#186410000000
1!
1%
1-
12
#186420000000
0!
0%
b1 *
0-
02
b1 6
#186430000000
1!
1%
1-
12
#186440000000
0!
0%
b10 *
0-
02
b10 6
#186450000000
1!
1%
1-
12
#186460000000
0!
0%
b11 *
0-
02
b11 6
#186470000000
1!
1%
1-
12
15
#186480000000
0!
0%
b100 *
0-
02
b100 6
#186490000000
1!
1%
1-
12
#186500000000
0!
0%
b101 *
0-
02
b101 6
#186510000000
1!
1%
1-
12
#186520000000
0!
0%
b110 *
0-
02
b110 6
#186530000000
1!
1%
1-
12
#186540000000
0!
0%
b111 *
0-
02
b111 6
#186550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#186560000000
0!
0%
b0 *
0-
02
b0 6
#186570000000
1!
1%
1-
12
#186580000000
0!
0%
b1 *
0-
02
b1 6
#186590000000
1!
1%
1-
12
#186600000000
0!
0%
b10 *
0-
02
b10 6
#186610000000
1!
1%
1-
12
#186620000000
0!
0%
b11 *
0-
02
b11 6
#186630000000
1!
1%
1-
12
15
#186640000000
0!
0%
b100 *
0-
02
b100 6
#186650000000
1!
1%
1-
12
#186660000000
0!
0%
b101 *
0-
02
b101 6
#186670000000
1!
1%
1-
12
#186680000000
0!
0%
b110 *
0-
02
b110 6
#186690000000
1!
1%
1-
12
#186700000000
0!
0%
b111 *
0-
02
b111 6
#186710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#186720000000
0!
0%
b0 *
0-
02
b0 6
#186730000000
1!
1%
1-
12
#186740000000
0!
0%
b1 *
0-
02
b1 6
#186750000000
1!
1%
1-
12
#186760000000
0!
0%
b10 *
0-
02
b10 6
#186770000000
1!
1%
1-
12
#186780000000
0!
0%
b11 *
0-
02
b11 6
#186790000000
1!
1%
1-
12
15
#186800000000
0!
0%
b100 *
0-
02
b100 6
#186810000000
1!
1%
1-
12
#186820000000
0!
0%
b101 *
0-
02
b101 6
#186830000000
1!
1%
1-
12
#186840000000
0!
0%
b110 *
0-
02
b110 6
#186850000000
1!
1%
1-
12
#186860000000
0!
0%
b111 *
0-
02
b111 6
#186870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#186880000000
0!
0%
b0 *
0-
02
b0 6
#186890000000
1!
1%
1-
12
#186900000000
0!
0%
b1 *
0-
02
b1 6
#186910000000
1!
1%
1-
12
#186920000000
0!
0%
b10 *
0-
02
b10 6
#186930000000
1!
1%
1-
12
#186940000000
0!
0%
b11 *
0-
02
b11 6
#186950000000
1!
1%
1-
12
15
#186960000000
0!
0%
b100 *
0-
02
b100 6
#186970000000
1!
1%
1-
12
#186980000000
0!
0%
b101 *
0-
02
b101 6
#186990000000
1!
1%
1-
12
#187000000000
0!
0%
b110 *
0-
02
b110 6
#187010000000
1!
1%
1-
12
#187020000000
0!
0%
b111 *
0-
02
b111 6
#187030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#187040000000
0!
0%
b0 *
0-
02
b0 6
#187050000000
1!
1%
1-
12
#187060000000
0!
0%
b1 *
0-
02
b1 6
#187070000000
1!
1%
1-
12
#187080000000
0!
0%
b10 *
0-
02
b10 6
#187090000000
1!
1%
1-
12
#187100000000
0!
0%
b11 *
0-
02
b11 6
#187110000000
1!
1%
1-
12
15
#187120000000
0!
0%
b100 *
0-
02
b100 6
#187130000000
1!
1%
1-
12
#187140000000
0!
0%
b101 *
0-
02
b101 6
#187150000000
1!
1%
1-
12
#187160000000
0!
0%
b110 *
0-
02
b110 6
#187170000000
1!
1%
1-
12
#187180000000
0!
0%
b111 *
0-
02
b111 6
#187190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#187200000000
0!
0%
b0 *
0-
02
b0 6
#187210000000
1!
1%
1-
12
#187220000000
0!
0%
b1 *
0-
02
b1 6
#187230000000
1!
1%
1-
12
#187240000000
0!
0%
b10 *
0-
02
b10 6
#187250000000
1!
1%
1-
12
#187260000000
0!
0%
b11 *
0-
02
b11 6
#187270000000
1!
1%
1-
12
15
#187280000000
0!
0%
b100 *
0-
02
b100 6
#187290000000
1!
1%
1-
12
#187300000000
0!
0%
b101 *
0-
02
b101 6
#187310000000
1!
1%
1-
12
#187320000000
0!
0%
b110 *
0-
02
b110 6
#187330000000
1!
1%
1-
12
#187340000000
0!
0%
b111 *
0-
02
b111 6
#187350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#187360000000
0!
0%
b0 *
0-
02
b0 6
#187370000000
1!
1%
1-
12
#187380000000
0!
0%
b1 *
0-
02
b1 6
#187390000000
1!
1%
1-
12
#187400000000
0!
0%
b10 *
0-
02
b10 6
#187410000000
1!
1%
1-
12
#187420000000
0!
0%
b11 *
0-
02
b11 6
#187430000000
1!
1%
1-
12
15
#187440000000
0!
0%
b100 *
0-
02
b100 6
#187450000000
1!
1%
1-
12
#187460000000
0!
0%
b101 *
0-
02
b101 6
#187470000000
1!
1%
1-
12
#187480000000
0!
0%
b110 *
0-
02
b110 6
#187490000000
1!
1%
1-
12
#187500000000
0!
0%
b111 *
0-
02
b111 6
#187510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#187520000000
0!
0%
b0 *
0-
02
b0 6
#187530000000
1!
1%
1-
12
#187540000000
0!
0%
b1 *
0-
02
b1 6
#187550000000
1!
1%
1-
12
#187560000000
0!
0%
b10 *
0-
02
b10 6
#187570000000
1!
1%
1-
12
#187580000000
0!
0%
b11 *
0-
02
b11 6
#187590000000
1!
1%
1-
12
15
#187600000000
0!
0%
b100 *
0-
02
b100 6
#187610000000
1!
1%
1-
12
#187620000000
0!
0%
b101 *
0-
02
b101 6
#187630000000
1!
1%
1-
12
#187640000000
0!
0%
b110 *
0-
02
b110 6
#187650000000
1!
1%
1-
12
#187660000000
0!
0%
b111 *
0-
02
b111 6
#187670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#187680000000
0!
0%
b0 *
0-
02
b0 6
#187690000000
1!
1%
1-
12
#187700000000
0!
0%
b1 *
0-
02
b1 6
#187710000000
1!
1%
1-
12
#187720000000
0!
0%
b10 *
0-
02
b10 6
#187730000000
1!
1%
1-
12
#187740000000
0!
0%
b11 *
0-
02
b11 6
#187750000000
1!
1%
1-
12
15
#187760000000
0!
0%
b100 *
0-
02
b100 6
#187770000000
1!
1%
1-
12
#187780000000
0!
0%
b101 *
0-
02
b101 6
#187790000000
1!
1%
1-
12
#187800000000
0!
0%
b110 *
0-
02
b110 6
#187810000000
1!
1%
1-
12
#187820000000
0!
0%
b111 *
0-
02
b111 6
#187830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#187840000000
0!
0%
b0 *
0-
02
b0 6
#187850000000
1!
1%
1-
12
#187860000000
0!
0%
b1 *
0-
02
b1 6
#187870000000
1!
1%
1-
12
#187880000000
0!
0%
b10 *
0-
02
b10 6
#187890000000
1!
1%
1-
12
#187900000000
0!
0%
b11 *
0-
02
b11 6
#187910000000
1!
1%
1-
12
15
#187920000000
0!
0%
b100 *
0-
02
b100 6
#187930000000
1!
1%
1-
12
#187940000000
0!
0%
b101 *
0-
02
b101 6
#187950000000
1!
1%
1-
12
#187960000000
0!
0%
b110 *
0-
02
b110 6
#187970000000
1!
1%
1-
12
#187980000000
0!
0%
b111 *
0-
02
b111 6
#187990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#188000000000
0!
0%
b0 *
0-
02
b0 6
#188010000000
1!
1%
1-
12
#188020000000
0!
0%
b1 *
0-
02
b1 6
#188030000000
1!
1%
1-
12
#188040000000
0!
0%
b10 *
0-
02
b10 6
#188050000000
1!
1%
1-
12
#188060000000
0!
0%
b11 *
0-
02
b11 6
#188070000000
1!
1%
1-
12
15
#188080000000
0!
0%
b100 *
0-
02
b100 6
#188090000000
1!
1%
1-
12
#188100000000
0!
0%
b101 *
0-
02
b101 6
#188110000000
1!
1%
1-
12
#188120000000
0!
0%
b110 *
0-
02
b110 6
#188130000000
1!
1%
1-
12
#188140000000
0!
0%
b111 *
0-
02
b111 6
#188150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#188160000000
0!
0%
b0 *
0-
02
b0 6
#188170000000
1!
1%
1-
12
#188180000000
0!
0%
b1 *
0-
02
b1 6
#188190000000
1!
1%
1-
12
#188200000000
0!
0%
b10 *
0-
02
b10 6
#188210000000
1!
1%
1-
12
#188220000000
0!
0%
b11 *
0-
02
b11 6
#188230000000
1!
1%
1-
12
15
#188240000000
0!
0%
b100 *
0-
02
b100 6
#188250000000
1!
1%
1-
12
#188260000000
0!
0%
b101 *
0-
02
b101 6
#188270000000
1!
1%
1-
12
#188280000000
0!
0%
b110 *
0-
02
b110 6
#188290000000
1!
1%
1-
12
#188300000000
0!
0%
b111 *
0-
02
b111 6
#188310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#188320000000
0!
0%
b0 *
0-
02
b0 6
#188330000000
1!
1%
1-
12
#188340000000
0!
0%
b1 *
0-
02
b1 6
#188350000000
1!
1%
1-
12
#188360000000
0!
0%
b10 *
0-
02
b10 6
#188370000000
1!
1%
1-
12
#188380000000
0!
0%
b11 *
0-
02
b11 6
#188390000000
1!
1%
1-
12
15
#188400000000
0!
0%
b100 *
0-
02
b100 6
#188410000000
1!
1%
1-
12
#188420000000
0!
0%
b101 *
0-
02
b101 6
#188430000000
1!
1%
1-
12
#188440000000
0!
0%
b110 *
0-
02
b110 6
#188450000000
1!
1%
1-
12
#188460000000
0!
0%
b111 *
0-
02
b111 6
#188470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#188480000000
0!
0%
b0 *
0-
02
b0 6
#188490000000
1!
1%
1-
12
#188500000000
0!
0%
b1 *
0-
02
b1 6
#188510000000
1!
1%
1-
12
#188520000000
0!
0%
b10 *
0-
02
b10 6
#188530000000
1!
1%
1-
12
#188540000000
0!
0%
b11 *
0-
02
b11 6
#188550000000
1!
1%
1-
12
15
#188560000000
0!
0%
b100 *
0-
02
b100 6
#188570000000
1!
1%
1-
12
#188580000000
0!
0%
b101 *
0-
02
b101 6
#188590000000
1!
1%
1-
12
#188600000000
0!
0%
b110 *
0-
02
b110 6
#188610000000
1!
1%
1-
12
#188620000000
0!
0%
b111 *
0-
02
b111 6
#188630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#188640000000
0!
0%
b0 *
0-
02
b0 6
#188650000000
1!
1%
1-
12
#188660000000
0!
0%
b1 *
0-
02
b1 6
#188670000000
1!
1%
1-
12
#188680000000
0!
0%
b10 *
0-
02
b10 6
#188690000000
1!
1%
1-
12
#188700000000
0!
0%
b11 *
0-
02
b11 6
#188710000000
1!
1%
1-
12
15
#188720000000
0!
0%
b100 *
0-
02
b100 6
#188730000000
1!
1%
1-
12
#188740000000
0!
0%
b101 *
0-
02
b101 6
#188750000000
1!
1%
1-
12
#188760000000
0!
0%
b110 *
0-
02
b110 6
#188770000000
1!
1%
1-
12
#188780000000
0!
0%
b111 *
0-
02
b111 6
#188790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#188800000000
0!
0%
b0 *
0-
02
b0 6
#188810000000
1!
1%
1-
12
#188820000000
0!
0%
b1 *
0-
02
b1 6
#188830000000
1!
1%
1-
12
#188840000000
0!
0%
b10 *
0-
02
b10 6
#188850000000
1!
1%
1-
12
#188860000000
0!
0%
b11 *
0-
02
b11 6
#188870000000
1!
1%
1-
12
15
#188880000000
0!
0%
b100 *
0-
02
b100 6
#188890000000
1!
1%
1-
12
#188900000000
0!
0%
b101 *
0-
02
b101 6
#188910000000
1!
1%
1-
12
#188920000000
0!
0%
b110 *
0-
02
b110 6
#188930000000
1!
1%
1-
12
#188940000000
0!
0%
b111 *
0-
02
b111 6
#188950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#188960000000
0!
0%
b0 *
0-
02
b0 6
#188970000000
1!
1%
1-
12
#188980000000
0!
0%
b1 *
0-
02
b1 6
#188990000000
1!
1%
1-
12
#189000000000
0!
0%
b10 *
0-
02
b10 6
#189010000000
1!
1%
1-
12
#189020000000
0!
0%
b11 *
0-
02
b11 6
#189030000000
1!
1%
1-
12
15
#189040000000
0!
0%
b100 *
0-
02
b100 6
#189050000000
1!
1%
1-
12
#189060000000
0!
0%
b101 *
0-
02
b101 6
#189070000000
1!
1%
1-
12
#189080000000
0!
0%
b110 *
0-
02
b110 6
#189090000000
1!
1%
1-
12
#189100000000
0!
0%
b111 *
0-
02
b111 6
#189110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#189120000000
0!
0%
b0 *
0-
02
b0 6
#189130000000
1!
1%
1-
12
#189140000000
0!
0%
b1 *
0-
02
b1 6
#189150000000
1!
1%
1-
12
#189160000000
0!
0%
b10 *
0-
02
b10 6
#189170000000
1!
1%
1-
12
#189180000000
0!
0%
b11 *
0-
02
b11 6
#189190000000
1!
1%
1-
12
15
#189200000000
0!
0%
b100 *
0-
02
b100 6
#189210000000
1!
1%
1-
12
#189220000000
0!
0%
b101 *
0-
02
b101 6
#189230000000
1!
1%
1-
12
#189240000000
0!
0%
b110 *
0-
02
b110 6
#189250000000
1!
1%
1-
12
#189260000000
0!
0%
b111 *
0-
02
b111 6
#189270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#189280000000
0!
0%
b0 *
0-
02
b0 6
#189290000000
1!
1%
1-
12
#189300000000
0!
0%
b1 *
0-
02
b1 6
#189310000000
1!
1%
1-
12
#189320000000
0!
0%
b10 *
0-
02
b10 6
#189330000000
1!
1%
1-
12
#189340000000
0!
0%
b11 *
0-
02
b11 6
#189350000000
1!
1%
1-
12
15
#189360000000
0!
0%
b100 *
0-
02
b100 6
#189370000000
1!
1%
1-
12
#189380000000
0!
0%
b101 *
0-
02
b101 6
#189390000000
1!
1%
1-
12
#189400000000
0!
0%
b110 *
0-
02
b110 6
#189410000000
1!
1%
1-
12
#189420000000
0!
0%
b111 *
0-
02
b111 6
#189430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#189440000000
0!
0%
b0 *
0-
02
b0 6
#189450000000
1!
1%
1-
12
#189460000000
0!
0%
b1 *
0-
02
b1 6
#189470000000
1!
1%
1-
12
#189480000000
0!
0%
b10 *
0-
02
b10 6
#189490000000
1!
1%
1-
12
#189500000000
0!
0%
b11 *
0-
02
b11 6
#189510000000
1!
1%
1-
12
15
#189520000000
0!
0%
b100 *
0-
02
b100 6
#189530000000
1!
1%
1-
12
#189540000000
0!
0%
b101 *
0-
02
b101 6
#189550000000
1!
1%
1-
12
#189560000000
0!
0%
b110 *
0-
02
b110 6
#189570000000
1!
1%
1-
12
#189580000000
0!
0%
b111 *
0-
02
b111 6
#189590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#189600000000
0!
0%
b0 *
0-
02
b0 6
#189610000000
1!
1%
1-
12
#189620000000
0!
0%
b1 *
0-
02
b1 6
#189630000000
1!
1%
1-
12
#189640000000
0!
0%
b10 *
0-
02
b10 6
#189650000000
1!
1%
1-
12
#189660000000
0!
0%
b11 *
0-
02
b11 6
#189670000000
1!
1%
1-
12
15
#189680000000
0!
0%
b100 *
0-
02
b100 6
#189690000000
1!
1%
1-
12
#189700000000
0!
0%
b101 *
0-
02
b101 6
#189710000000
1!
1%
1-
12
#189720000000
0!
0%
b110 *
0-
02
b110 6
#189730000000
1!
1%
1-
12
#189740000000
0!
0%
b111 *
0-
02
b111 6
#189750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#189760000000
0!
0%
b0 *
0-
02
b0 6
#189770000000
1!
1%
1-
12
#189780000000
0!
0%
b1 *
0-
02
b1 6
#189790000000
1!
1%
1-
12
#189800000000
0!
0%
b10 *
0-
02
b10 6
#189810000000
1!
1%
1-
12
#189820000000
0!
0%
b11 *
0-
02
b11 6
#189830000000
1!
1%
1-
12
15
#189840000000
0!
0%
b100 *
0-
02
b100 6
#189850000000
1!
1%
1-
12
#189860000000
0!
0%
b101 *
0-
02
b101 6
#189870000000
1!
1%
1-
12
#189880000000
0!
0%
b110 *
0-
02
b110 6
#189890000000
1!
1%
1-
12
#189900000000
0!
0%
b111 *
0-
02
b111 6
#189910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#189920000000
0!
0%
b0 *
0-
02
b0 6
#189930000000
1!
1%
1-
12
#189940000000
0!
0%
b1 *
0-
02
b1 6
#189950000000
1!
1%
1-
12
#189960000000
0!
0%
b10 *
0-
02
b10 6
#189970000000
1!
1%
1-
12
#189980000000
0!
0%
b11 *
0-
02
b11 6
#189990000000
1!
1%
1-
12
15
#190000000000
0!
0%
b100 *
0-
02
b100 6
#190010000000
1!
1%
1-
12
#190020000000
0!
0%
b101 *
0-
02
b101 6
#190030000000
1!
1%
1-
12
#190040000000
0!
0%
b110 *
0-
02
b110 6
#190050000000
1!
1%
1-
12
#190060000000
0!
0%
b111 *
0-
02
b111 6
#190070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#190080000000
0!
0%
b0 *
0-
02
b0 6
#190090000000
1!
1%
1-
12
#190100000000
0!
0%
b1 *
0-
02
b1 6
#190110000000
1!
1%
1-
12
#190120000000
0!
0%
b10 *
0-
02
b10 6
#190130000000
1!
1%
1-
12
#190140000000
0!
0%
b11 *
0-
02
b11 6
#190150000000
1!
1%
1-
12
15
#190160000000
0!
0%
b100 *
0-
02
b100 6
#190170000000
1!
1%
1-
12
#190180000000
0!
0%
b101 *
0-
02
b101 6
#190190000000
1!
1%
1-
12
#190200000000
0!
0%
b110 *
0-
02
b110 6
#190210000000
1!
1%
1-
12
#190220000000
0!
0%
b111 *
0-
02
b111 6
#190230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#190240000000
0!
0%
b0 *
0-
02
b0 6
#190250000000
1!
1%
1-
12
#190260000000
0!
0%
b1 *
0-
02
b1 6
#190270000000
1!
1%
1-
12
#190280000000
0!
0%
b10 *
0-
02
b10 6
#190290000000
1!
1%
1-
12
#190300000000
0!
0%
b11 *
0-
02
b11 6
#190310000000
1!
1%
1-
12
15
#190320000000
0!
0%
b100 *
0-
02
b100 6
#190330000000
1!
1%
1-
12
#190340000000
0!
0%
b101 *
0-
02
b101 6
#190350000000
1!
1%
1-
12
#190360000000
0!
0%
b110 *
0-
02
b110 6
#190370000000
1!
1%
1-
12
#190380000000
0!
0%
b111 *
0-
02
b111 6
#190390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#190400000000
0!
0%
b0 *
0-
02
b0 6
#190410000000
1!
1%
1-
12
#190420000000
0!
0%
b1 *
0-
02
b1 6
#190430000000
1!
1%
1-
12
#190440000000
0!
0%
b10 *
0-
02
b10 6
#190450000000
1!
1%
1-
12
#190460000000
0!
0%
b11 *
0-
02
b11 6
#190470000000
1!
1%
1-
12
15
#190480000000
0!
0%
b100 *
0-
02
b100 6
#190490000000
1!
1%
1-
12
#190500000000
0!
0%
b101 *
0-
02
b101 6
#190510000000
1!
1%
1-
12
#190520000000
0!
0%
b110 *
0-
02
b110 6
#190530000000
1!
1%
1-
12
#190540000000
0!
0%
b111 *
0-
02
b111 6
#190550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#190560000000
0!
0%
b0 *
0-
02
b0 6
#190570000000
1!
1%
1-
12
#190580000000
0!
0%
b1 *
0-
02
b1 6
#190590000000
1!
1%
1-
12
#190600000000
0!
0%
b10 *
0-
02
b10 6
#190610000000
1!
1%
1-
12
#190620000000
0!
0%
b11 *
0-
02
b11 6
#190630000000
1!
1%
1-
12
15
#190640000000
0!
0%
b100 *
0-
02
b100 6
#190650000000
1!
1%
1-
12
#190660000000
0!
0%
b101 *
0-
02
b101 6
#190670000000
1!
1%
1-
12
#190680000000
0!
0%
b110 *
0-
02
b110 6
#190690000000
1!
1%
1-
12
#190700000000
0!
0%
b111 *
0-
02
b111 6
#190710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#190720000000
0!
0%
b0 *
0-
02
b0 6
#190730000000
1!
1%
1-
12
#190740000000
0!
0%
b1 *
0-
02
b1 6
#190750000000
1!
1%
1-
12
#190760000000
0!
0%
b10 *
0-
02
b10 6
#190770000000
1!
1%
1-
12
#190780000000
0!
0%
b11 *
0-
02
b11 6
#190790000000
1!
1%
1-
12
15
#190800000000
0!
0%
b100 *
0-
02
b100 6
#190810000000
1!
1%
1-
12
#190820000000
0!
0%
b101 *
0-
02
b101 6
#190830000000
1!
1%
1-
12
#190840000000
0!
0%
b110 *
0-
02
b110 6
#190850000000
1!
1%
1-
12
#190860000000
0!
0%
b111 *
0-
02
b111 6
#190870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#190880000000
0!
0%
b0 *
0-
02
b0 6
#190890000000
1!
1%
1-
12
#190900000000
0!
0%
b1 *
0-
02
b1 6
#190910000000
1!
1%
1-
12
#190920000000
0!
0%
b10 *
0-
02
b10 6
#190930000000
1!
1%
1-
12
#190940000000
0!
0%
b11 *
0-
02
b11 6
#190950000000
1!
1%
1-
12
15
#190960000000
0!
0%
b100 *
0-
02
b100 6
#190970000000
1!
1%
1-
12
#190980000000
0!
0%
b101 *
0-
02
b101 6
#190990000000
1!
1%
1-
12
#191000000000
0!
0%
b110 *
0-
02
b110 6
#191010000000
1!
1%
1-
12
#191020000000
0!
0%
b111 *
0-
02
b111 6
#191030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#191040000000
0!
0%
b0 *
0-
02
b0 6
#191050000000
1!
1%
1-
12
#191060000000
0!
0%
b1 *
0-
02
b1 6
#191070000000
1!
1%
1-
12
#191080000000
0!
0%
b10 *
0-
02
b10 6
#191090000000
1!
1%
1-
12
#191100000000
0!
0%
b11 *
0-
02
b11 6
#191110000000
1!
1%
1-
12
15
#191120000000
0!
0%
b100 *
0-
02
b100 6
#191130000000
1!
1%
1-
12
#191140000000
0!
0%
b101 *
0-
02
b101 6
#191150000000
1!
1%
1-
12
#191160000000
0!
0%
b110 *
0-
02
b110 6
#191170000000
1!
1%
1-
12
#191180000000
0!
0%
b111 *
0-
02
b111 6
#191190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#191200000000
0!
0%
b0 *
0-
02
b0 6
#191210000000
1!
1%
1-
12
#191220000000
0!
0%
b1 *
0-
02
b1 6
#191230000000
1!
1%
1-
12
#191240000000
0!
0%
b10 *
0-
02
b10 6
#191250000000
1!
1%
1-
12
#191260000000
0!
0%
b11 *
0-
02
b11 6
#191270000000
1!
1%
1-
12
15
#191280000000
0!
0%
b100 *
0-
02
b100 6
#191290000000
1!
1%
1-
12
#191300000000
0!
0%
b101 *
0-
02
b101 6
#191310000000
1!
1%
1-
12
#191320000000
0!
0%
b110 *
0-
02
b110 6
#191330000000
1!
1%
1-
12
#191340000000
0!
0%
b111 *
0-
02
b111 6
#191350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#191360000000
0!
0%
b0 *
0-
02
b0 6
#191370000000
1!
1%
1-
12
#191380000000
0!
0%
b1 *
0-
02
b1 6
#191390000000
1!
1%
1-
12
#191400000000
0!
0%
b10 *
0-
02
b10 6
#191410000000
1!
1%
1-
12
#191420000000
0!
0%
b11 *
0-
02
b11 6
#191430000000
1!
1%
1-
12
15
#191440000000
0!
0%
b100 *
0-
02
b100 6
#191450000000
1!
1%
1-
12
#191460000000
0!
0%
b101 *
0-
02
b101 6
#191470000000
1!
1%
1-
12
#191480000000
0!
0%
b110 *
0-
02
b110 6
#191490000000
1!
1%
1-
12
#191500000000
0!
0%
b111 *
0-
02
b111 6
#191510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#191520000000
0!
0%
b0 *
0-
02
b0 6
#191530000000
1!
1%
1-
12
#191540000000
0!
0%
b1 *
0-
02
b1 6
#191550000000
1!
1%
1-
12
#191560000000
0!
0%
b10 *
0-
02
b10 6
#191570000000
1!
1%
1-
12
#191580000000
0!
0%
b11 *
0-
02
b11 6
#191590000000
1!
1%
1-
12
15
#191600000000
0!
0%
b100 *
0-
02
b100 6
#191610000000
1!
1%
1-
12
#191620000000
0!
0%
b101 *
0-
02
b101 6
#191630000000
1!
1%
1-
12
#191640000000
0!
0%
b110 *
0-
02
b110 6
#191650000000
1!
1%
1-
12
#191660000000
0!
0%
b111 *
0-
02
b111 6
#191670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#191680000000
0!
0%
b0 *
0-
02
b0 6
#191690000000
1!
1%
1-
12
#191700000000
0!
0%
b1 *
0-
02
b1 6
#191710000000
1!
1%
1-
12
#191720000000
0!
0%
b10 *
0-
02
b10 6
#191730000000
1!
1%
1-
12
#191740000000
0!
0%
b11 *
0-
02
b11 6
#191750000000
1!
1%
1-
12
15
#191760000000
0!
0%
b100 *
0-
02
b100 6
#191770000000
1!
1%
1-
12
#191780000000
0!
0%
b101 *
0-
02
b101 6
#191790000000
1!
1%
1-
12
#191800000000
0!
0%
b110 *
0-
02
b110 6
#191810000000
1!
1%
1-
12
#191820000000
0!
0%
b111 *
0-
02
b111 6
#191830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#191840000000
0!
0%
b0 *
0-
02
b0 6
#191850000000
1!
1%
1-
12
#191860000000
0!
0%
b1 *
0-
02
b1 6
#191870000000
1!
1%
1-
12
#191880000000
0!
0%
b10 *
0-
02
b10 6
#191890000000
1!
1%
1-
12
#191900000000
0!
0%
b11 *
0-
02
b11 6
#191910000000
1!
1%
1-
12
15
#191920000000
0!
0%
b100 *
0-
02
b100 6
#191930000000
1!
1%
1-
12
#191940000000
0!
0%
b101 *
0-
02
b101 6
#191950000000
1!
1%
1-
12
#191960000000
0!
0%
b110 *
0-
02
b110 6
#191970000000
1!
1%
1-
12
#191980000000
0!
0%
b111 *
0-
02
b111 6
#191990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#192000000000
0!
0%
b0 *
0-
02
b0 6
#192010000000
1!
1%
1-
12
#192020000000
0!
0%
b1 *
0-
02
b1 6
#192030000000
1!
1%
1-
12
#192040000000
0!
0%
b10 *
0-
02
b10 6
#192050000000
1!
1%
1-
12
#192060000000
0!
0%
b11 *
0-
02
b11 6
#192070000000
1!
1%
1-
12
15
#192080000000
0!
0%
b100 *
0-
02
b100 6
#192090000000
1!
1%
1-
12
#192100000000
0!
0%
b101 *
0-
02
b101 6
#192110000000
1!
1%
1-
12
#192120000000
0!
0%
b110 *
0-
02
b110 6
#192130000000
1!
1%
1-
12
#192140000000
0!
0%
b111 *
0-
02
b111 6
#192150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#192160000000
0!
0%
b0 *
0-
02
b0 6
#192170000000
1!
1%
1-
12
#192180000000
0!
0%
b1 *
0-
02
b1 6
#192190000000
1!
1%
1-
12
#192200000000
0!
0%
b10 *
0-
02
b10 6
#192210000000
1!
1%
1-
12
#192220000000
0!
0%
b11 *
0-
02
b11 6
#192230000000
1!
1%
1-
12
15
#192240000000
0!
0%
b100 *
0-
02
b100 6
#192250000000
1!
1%
1-
12
#192260000000
0!
0%
b101 *
0-
02
b101 6
#192270000000
1!
1%
1-
12
#192280000000
0!
0%
b110 *
0-
02
b110 6
#192290000000
1!
1%
1-
12
#192300000000
0!
0%
b111 *
0-
02
b111 6
#192310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#192320000000
0!
0%
b0 *
0-
02
b0 6
#192330000000
1!
1%
1-
12
#192340000000
0!
0%
b1 *
0-
02
b1 6
#192350000000
1!
1%
1-
12
#192360000000
0!
0%
b10 *
0-
02
b10 6
#192370000000
1!
1%
1-
12
#192380000000
0!
0%
b11 *
0-
02
b11 6
#192390000000
1!
1%
1-
12
15
#192400000000
0!
0%
b100 *
0-
02
b100 6
#192410000000
1!
1%
1-
12
#192420000000
0!
0%
b101 *
0-
02
b101 6
#192430000000
1!
1%
1-
12
#192440000000
0!
0%
b110 *
0-
02
b110 6
#192450000000
1!
1%
1-
12
#192460000000
0!
0%
b111 *
0-
02
b111 6
#192470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#192480000000
0!
0%
b0 *
0-
02
b0 6
#192490000000
1!
1%
1-
12
#192500000000
0!
0%
b1 *
0-
02
b1 6
#192510000000
1!
1%
1-
12
#192520000000
0!
0%
b10 *
0-
02
b10 6
#192530000000
1!
1%
1-
12
#192540000000
0!
0%
b11 *
0-
02
b11 6
#192550000000
1!
1%
1-
12
15
#192560000000
0!
0%
b100 *
0-
02
b100 6
#192570000000
1!
1%
1-
12
#192580000000
0!
0%
b101 *
0-
02
b101 6
#192590000000
1!
1%
1-
12
#192600000000
0!
0%
b110 *
0-
02
b110 6
#192610000000
1!
1%
1-
12
#192620000000
0!
0%
b111 *
0-
02
b111 6
#192630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#192640000000
0!
0%
b0 *
0-
02
b0 6
#192650000000
1!
1%
1-
12
#192660000000
0!
0%
b1 *
0-
02
b1 6
#192670000000
1!
1%
1-
12
#192680000000
0!
0%
b10 *
0-
02
b10 6
#192690000000
1!
1%
1-
12
#192700000000
0!
0%
b11 *
0-
02
b11 6
#192710000000
1!
1%
1-
12
15
#192720000000
0!
0%
b100 *
0-
02
b100 6
#192730000000
1!
1%
1-
12
#192740000000
0!
0%
b101 *
0-
02
b101 6
#192750000000
1!
1%
1-
12
#192760000000
0!
0%
b110 *
0-
02
b110 6
#192770000000
1!
1%
1-
12
#192780000000
0!
0%
b111 *
0-
02
b111 6
#192790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#192800000000
0!
0%
b0 *
0-
02
b0 6
#192810000000
1!
1%
1-
12
#192820000000
0!
0%
b1 *
0-
02
b1 6
#192830000000
1!
1%
1-
12
#192840000000
0!
0%
b10 *
0-
02
b10 6
#192850000000
1!
1%
1-
12
#192860000000
0!
0%
b11 *
0-
02
b11 6
#192870000000
1!
1%
1-
12
15
#192880000000
0!
0%
b100 *
0-
02
b100 6
#192890000000
1!
1%
1-
12
#192900000000
0!
0%
b101 *
0-
02
b101 6
#192910000000
1!
1%
1-
12
#192920000000
0!
0%
b110 *
0-
02
b110 6
#192930000000
1!
1%
1-
12
#192940000000
0!
0%
b111 *
0-
02
b111 6
#192950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#192960000000
0!
0%
b0 *
0-
02
b0 6
#192970000000
1!
1%
1-
12
#192980000000
0!
0%
b1 *
0-
02
b1 6
#192990000000
1!
1%
1-
12
#193000000000
0!
0%
b10 *
0-
02
b10 6
#193010000000
1!
1%
1-
12
#193020000000
0!
0%
b11 *
0-
02
b11 6
#193030000000
1!
1%
1-
12
15
#193040000000
0!
0%
b100 *
0-
02
b100 6
#193050000000
1!
1%
1-
12
#193060000000
0!
0%
b101 *
0-
02
b101 6
#193070000000
1!
1%
1-
12
#193080000000
0!
0%
b110 *
0-
02
b110 6
#193090000000
1!
1%
1-
12
#193100000000
0!
0%
b111 *
0-
02
b111 6
#193110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#193120000000
0!
0%
b0 *
0-
02
b0 6
#193130000000
1!
1%
1-
12
#193140000000
0!
0%
b1 *
0-
02
b1 6
#193150000000
1!
1%
1-
12
#193160000000
0!
0%
b10 *
0-
02
b10 6
#193170000000
1!
1%
1-
12
#193180000000
0!
0%
b11 *
0-
02
b11 6
#193190000000
1!
1%
1-
12
15
#193200000000
0!
0%
b100 *
0-
02
b100 6
#193210000000
1!
1%
1-
12
#193220000000
0!
0%
b101 *
0-
02
b101 6
#193230000000
1!
1%
1-
12
#193240000000
0!
0%
b110 *
0-
02
b110 6
#193250000000
1!
1%
1-
12
#193260000000
0!
0%
b111 *
0-
02
b111 6
#193270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#193280000000
0!
0%
b0 *
0-
02
b0 6
#193290000000
1!
1%
1-
12
#193300000000
0!
0%
b1 *
0-
02
b1 6
#193310000000
1!
1%
1-
12
#193320000000
0!
0%
b10 *
0-
02
b10 6
#193330000000
1!
1%
1-
12
#193340000000
0!
0%
b11 *
0-
02
b11 6
#193350000000
1!
1%
1-
12
15
#193360000000
0!
0%
b100 *
0-
02
b100 6
#193370000000
1!
1%
1-
12
#193380000000
0!
0%
b101 *
0-
02
b101 6
#193390000000
1!
1%
1-
12
#193400000000
0!
0%
b110 *
0-
02
b110 6
#193410000000
1!
1%
1-
12
#193420000000
0!
0%
b111 *
0-
02
b111 6
#193430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#193440000000
0!
0%
b0 *
0-
02
b0 6
#193450000000
1!
1%
1-
12
#193460000000
0!
0%
b1 *
0-
02
b1 6
#193470000000
1!
1%
1-
12
#193480000000
0!
0%
b10 *
0-
02
b10 6
#193490000000
1!
1%
1-
12
#193500000000
0!
0%
b11 *
0-
02
b11 6
#193510000000
1!
1%
1-
12
15
#193520000000
0!
0%
b100 *
0-
02
b100 6
#193530000000
1!
1%
1-
12
#193540000000
0!
0%
b101 *
0-
02
b101 6
#193550000000
1!
1%
1-
12
#193560000000
0!
0%
b110 *
0-
02
b110 6
#193570000000
1!
1%
1-
12
#193580000000
0!
0%
b111 *
0-
02
b111 6
#193590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#193600000000
0!
0%
b0 *
0-
02
b0 6
#193610000000
1!
1%
1-
12
#193620000000
0!
0%
b1 *
0-
02
b1 6
#193630000000
1!
1%
1-
12
#193640000000
0!
0%
b10 *
0-
02
b10 6
#193650000000
1!
1%
1-
12
#193660000000
0!
0%
b11 *
0-
02
b11 6
#193670000000
1!
1%
1-
12
15
#193680000000
0!
0%
b100 *
0-
02
b100 6
#193690000000
1!
1%
1-
12
#193700000000
0!
0%
b101 *
0-
02
b101 6
#193710000000
1!
1%
1-
12
#193720000000
0!
0%
b110 *
0-
02
b110 6
#193730000000
1!
1%
1-
12
#193740000000
0!
0%
b111 *
0-
02
b111 6
#193750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#193760000000
0!
0%
b0 *
0-
02
b0 6
#193770000000
1!
1%
1-
12
#193780000000
0!
0%
b1 *
0-
02
b1 6
#193790000000
1!
1%
1-
12
#193800000000
0!
0%
b10 *
0-
02
b10 6
#193810000000
1!
1%
1-
12
#193820000000
0!
0%
b11 *
0-
02
b11 6
#193830000000
1!
1%
1-
12
15
#193840000000
0!
0%
b100 *
0-
02
b100 6
#193850000000
1!
1%
1-
12
#193860000000
0!
0%
b101 *
0-
02
b101 6
#193870000000
1!
1%
1-
12
#193880000000
0!
0%
b110 *
0-
02
b110 6
#193890000000
1!
1%
1-
12
#193900000000
0!
0%
b111 *
0-
02
b111 6
#193910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#193920000000
0!
0%
b0 *
0-
02
b0 6
#193930000000
1!
1%
1-
12
#193940000000
0!
0%
b1 *
0-
02
b1 6
#193950000000
1!
1%
1-
12
#193960000000
0!
0%
b10 *
0-
02
b10 6
#193970000000
1!
1%
1-
12
#193980000000
0!
0%
b11 *
0-
02
b11 6
#193990000000
1!
1%
1-
12
15
#194000000000
0!
0%
b100 *
0-
02
b100 6
#194010000000
1!
1%
1-
12
#194020000000
0!
0%
b101 *
0-
02
b101 6
#194030000000
1!
1%
1-
12
#194040000000
0!
0%
b110 *
0-
02
b110 6
#194050000000
1!
1%
1-
12
#194060000000
0!
0%
b111 *
0-
02
b111 6
#194070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#194080000000
0!
0%
b0 *
0-
02
b0 6
#194090000000
1!
1%
1-
12
#194100000000
0!
0%
b1 *
0-
02
b1 6
#194110000000
1!
1%
1-
12
#194120000000
0!
0%
b10 *
0-
02
b10 6
#194130000000
1!
1%
1-
12
#194140000000
0!
0%
b11 *
0-
02
b11 6
#194150000000
1!
1%
1-
12
15
#194160000000
0!
0%
b100 *
0-
02
b100 6
#194170000000
1!
1%
1-
12
#194180000000
0!
0%
b101 *
0-
02
b101 6
#194190000000
1!
1%
1-
12
#194200000000
0!
0%
b110 *
0-
02
b110 6
#194210000000
1!
1%
1-
12
#194220000000
0!
0%
b111 *
0-
02
b111 6
#194230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#194240000000
0!
0%
b0 *
0-
02
b0 6
#194250000000
1!
1%
1-
12
#194260000000
0!
0%
b1 *
0-
02
b1 6
#194270000000
1!
1%
1-
12
#194280000000
0!
0%
b10 *
0-
02
b10 6
#194290000000
1!
1%
1-
12
#194300000000
0!
0%
b11 *
0-
02
b11 6
#194310000000
1!
1%
1-
12
15
#194320000000
0!
0%
b100 *
0-
02
b100 6
#194330000000
1!
1%
1-
12
#194340000000
0!
0%
b101 *
0-
02
b101 6
#194350000000
1!
1%
1-
12
#194360000000
0!
0%
b110 *
0-
02
b110 6
#194370000000
1!
1%
1-
12
#194380000000
0!
0%
b111 *
0-
02
b111 6
#194390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#194400000000
0!
0%
b0 *
0-
02
b0 6
#194410000000
1!
1%
1-
12
#194420000000
0!
0%
b1 *
0-
02
b1 6
#194430000000
1!
1%
1-
12
#194440000000
0!
0%
b10 *
0-
02
b10 6
#194450000000
1!
1%
1-
12
#194460000000
0!
0%
b11 *
0-
02
b11 6
#194470000000
1!
1%
1-
12
15
#194480000000
0!
0%
b100 *
0-
02
b100 6
#194490000000
1!
1%
1-
12
#194500000000
0!
0%
b101 *
0-
02
b101 6
#194510000000
1!
1%
1-
12
#194520000000
0!
0%
b110 *
0-
02
b110 6
#194530000000
1!
1%
1-
12
#194540000000
0!
0%
b111 *
0-
02
b111 6
#194550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#194560000000
0!
0%
b0 *
0-
02
b0 6
#194570000000
1!
1%
1-
12
#194580000000
0!
0%
b1 *
0-
02
b1 6
#194590000000
1!
1%
1-
12
#194600000000
0!
0%
b10 *
0-
02
b10 6
#194610000000
1!
1%
1-
12
#194620000000
0!
0%
b11 *
0-
02
b11 6
#194630000000
1!
1%
1-
12
15
#194640000000
0!
0%
b100 *
0-
02
b100 6
#194650000000
1!
1%
1-
12
#194660000000
0!
0%
b101 *
0-
02
b101 6
#194670000000
1!
1%
1-
12
#194680000000
0!
0%
b110 *
0-
02
b110 6
#194690000000
1!
1%
1-
12
#194700000000
0!
0%
b111 *
0-
02
b111 6
#194710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#194720000000
0!
0%
b0 *
0-
02
b0 6
#194730000000
1!
1%
1-
12
#194740000000
0!
0%
b1 *
0-
02
b1 6
#194750000000
1!
1%
1-
12
#194760000000
0!
0%
b10 *
0-
02
b10 6
#194770000000
1!
1%
1-
12
#194780000000
0!
0%
b11 *
0-
02
b11 6
#194790000000
1!
1%
1-
12
15
#194800000000
0!
0%
b100 *
0-
02
b100 6
#194810000000
1!
1%
1-
12
#194820000000
0!
0%
b101 *
0-
02
b101 6
#194830000000
1!
1%
1-
12
#194840000000
0!
0%
b110 *
0-
02
b110 6
#194850000000
1!
1%
1-
12
#194860000000
0!
0%
b111 *
0-
02
b111 6
#194870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#194880000000
0!
0%
b0 *
0-
02
b0 6
#194890000000
1!
1%
1-
12
#194900000000
0!
0%
b1 *
0-
02
b1 6
#194910000000
1!
1%
1-
12
#194920000000
0!
0%
b10 *
0-
02
b10 6
#194930000000
1!
1%
1-
12
#194940000000
0!
0%
b11 *
0-
02
b11 6
#194950000000
1!
1%
1-
12
15
#194960000000
0!
0%
b100 *
0-
02
b100 6
#194970000000
1!
1%
1-
12
#194980000000
0!
0%
b101 *
0-
02
b101 6
#194990000000
1!
1%
1-
12
#195000000000
0!
0%
b110 *
0-
02
b110 6
#195010000000
1!
1%
1-
12
#195020000000
0!
0%
b111 *
0-
02
b111 6
#195030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#195040000000
0!
0%
b0 *
0-
02
b0 6
#195050000000
1!
1%
1-
12
#195060000000
0!
0%
b1 *
0-
02
b1 6
#195070000000
1!
1%
1-
12
#195080000000
0!
0%
b10 *
0-
02
b10 6
#195090000000
1!
1%
1-
12
#195100000000
0!
0%
b11 *
0-
02
b11 6
#195110000000
1!
1%
1-
12
15
#195120000000
0!
0%
b100 *
0-
02
b100 6
#195130000000
1!
1%
1-
12
#195140000000
0!
0%
b101 *
0-
02
b101 6
#195150000000
1!
1%
1-
12
#195160000000
0!
0%
b110 *
0-
02
b110 6
#195170000000
1!
1%
1-
12
#195180000000
0!
0%
b111 *
0-
02
b111 6
#195190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#195200000000
0!
0%
b0 *
0-
02
b0 6
#195210000000
1!
1%
1-
12
#195220000000
0!
0%
b1 *
0-
02
b1 6
#195230000000
1!
1%
1-
12
#195240000000
0!
0%
b10 *
0-
02
b10 6
#195250000000
1!
1%
1-
12
#195260000000
0!
0%
b11 *
0-
02
b11 6
#195270000000
1!
1%
1-
12
15
#195280000000
0!
0%
b100 *
0-
02
b100 6
#195290000000
1!
1%
1-
12
#195300000000
0!
0%
b101 *
0-
02
b101 6
#195310000000
1!
1%
1-
12
#195320000000
0!
0%
b110 *
0-
02
b110 6
#195330000000
1!
1%
1-
12
#195340000000
0!
0%
b111 *
0-
02
b111 6
#195350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#195360000000
0!
0%
b0 *
0-
02
b0 6
#195370000000
1!
1%
1-
12
#195380000000
0!
0%
b1 *
0-
02
b1 6
#195390000000
1!
1%
1-
12
#195400000000
0!
0%
b10 *
0-
02
b10 6
#195410000000
1!
1%
1-
12
#195420000000
0!
0%
b11 *
0-
02
b11 6
#195430000000
1!
1%
1-
12
15
#195440000000
0!
0%
b100 *
0-
02
b100 6
#195450000000
1!
1%
1-
12
#195460000000
0!
0%
b101 *
0-
02
b101 6
#195470000000
1!
1%
1-
12
#195480000000
0!
0%
b110 *
0-
02
b110 6
#195490000000
1!
1%
1-
12
#195500000000
0!
0%
b111 *
0-
02
b111 6
#195510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#195520000000
0!
0%
b0 *
0-
02
b0 6
#195530000000
1!
1%
1-
12
#195540000000
0!
0%
b1 *
0-
02
b1 6
#195550000000
1!
1%
1-
12
#195560000000
0!
0%
b10 *
0-
02
b10 6
#195570000000
1!
1%
1-
12
#195580000000
0!
0%
b11 *
0-
02
b11 6
#195590000000
1!
1%
1-
12
15
#195600000000
0!
0%
b100 *
0-
02
b100 6
#195610000000
1!
1%
1-
12
#195620000000
0!
0%
b101 *
0-
02
b101 6
#195630000000
1!
1%
1-
12
#195640000000
0!
0%
b110 *
0-
02
b110 6
#195650000000
1!
1%
1-
12
#195660000000
0!
0%
b111 *
0-
02
b111 6
#195670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#195680000000
0!
0%
b0 *
0-
02
b0 6
#195690000000
1!
1%
1-
12
#195700000000
0!
0%
b1 *
0-
02
b1 6
#195710000000
1!
1%
1-
12
#195720000000
0!
0%
b10 *
0-
02
b10 6
#195730000000
1!
1%
1-
12
#195740000000
0!
0%
b11 *
0-
02
b11 6
#195750000000
1!
1%
1-
12
15
#195760000000
0!
0%
b100 *
0-
02
b100 6
#195770000000
1!
1%
1-
12
#195780000000
0!
0%
b101 *
0-
02
b101 6
#195790000000
1!
1%
1-
12
#195800000000
0!
0%
b110 *
0-
02
b110 6
#195810000000
1!
1%
1-
12
#195820000000
0!
0%
b111 *
0-
02
b111 6
#195830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#195840000000
0!
0%
b0 *
0-
02
b0 6
#195850000000
1!
1%
1-
12
#195860000000
0!
0%
b1 *
0-
02
b1 6
#195870000000
1!
1%
1-
12
#195880000000
0!
0%
b10 *
0-
02
b10 6
#195890000000
1!
1%
1-
12
#195900000000
0!
0%
b11 *
0-
02
b11 6
#195910000000
1!
1%
1-
12
15
#195920000000
0!
0%
b100 *
0-
02
b100 6
#195930000000
1!
1%
1-
12
#195940000000
0!
0%
b101 *
0-
02
b101 6
#195950000000
1!
1%
1-
12
#195960000000
0!
0%
b110 *
0-
02
b110 6
#195970000000
1!
1%
1-
12
#195980000000
0!
0%
b111 *
0-
02
b111 6
#195990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#196000000000
0!
0%
b0 *
0-
02
b0 6
#196010000000
1!
1%
1-
12
#196020000000
0!
0%
b1 *
0-
02
b1 6
#196030000000
1!
1%
1-
12
#196040000000
0!
0%
b10 *
0-
02
b10 6
#196050000000
1!
1%
1-
12
#196060000000
0!
0%
b11 *
0-
02
b11 6
#196070000000
1!
1%
1-
12
15
#196080000000
0!
0%
b100 *
0-
02
b100 6
#196090000000
1!
1%
1-
12
#196100000000
0!
0%
b101 *
0-
02
b101 6
#196110000000
1!
1%
1-
12
#196120000000
0!
0%
b110 *
0-
02
b110 6
#196130000000
1!
1%
1-
12
#196140000000
0!
0%
b111 *
0-
02
b111 6
#196150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#196160000000
0!
0%
b0 *
0-
02
b0 6
#196170000000
1!
1%
1-
12
#196180000000
0!
0%
b1 *
0-
02
b1 6
#196190000000
1!
1%
1-
12
#196200000000
0!
0%
b10 *
0-
02
b10 6
#196210000000
1!
1%
1-
12
#196220000000
0!
0%
b11 *
0-
02
b11 6
#196230000000
1!
1%
1-
12
15
#196240000000
0!
0%
b100 *
0-
02
b100 6
#196250000000
1!
1%
1-
12
#196260000000
0!
0%
b101 *
0-
02
b101 6
#196270000000
1!
1%
1-
12
#196280000000
0!
0%
b110 *
0-
02
b110 6
#196290000000
1!
1%
1-
12
#196300000000
0!
0%
b111 *
0-
02
b111 6
#196310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#196320000000
0!
0%
b0 *
0-
02
b0 6
#196330000000
1!
1%
1-
12
#196340000000
0!
0%
b1 *
0-
02
b1 6
#196350000000
1!
1%
1-
12
#196360000000
0!
0%
b10 *
0-
02
b10 6
#196370000000
1!
1%
1-
12
#196380000000
0!
0%
b11 *
0-
02
b11 6
#196390000000
1!
1%
1-
12
15
#196400000000
0!
0%
b100 *
0-
02
b100 6
#196410000000
1!
1%
1-
12
#196420000000
0!
0%
b101 *
0-
02
b101 6
#196430000000
1!
1%
1-
12
#196440000000
0!
0%
b110 *
0-
02
b110 6
#196450000000
1!
1%
1-
12
#196460000000
0!
0%
b111 *
0-
02
b111 6
#196470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#196480000000
0!
0%
b0 *
0-
02
b0 6
#196490000000
1!
1%
1-
12
#196500000000
0!
0%
b1 *
0-
02
b1 6
#196510000000
1!
1%
1-
12
#196520000000
0!
0%
b10 *
0-
02
b10 6
#196530000000
1!
1%
1-
12
#196540000000
0!
0%
b11 *
0-
02
b11 6
#196550000000
1!
1%
1-
12
15
#196560000000
0!
0%
b100 *
0-
02
b100 6
#196570000000
1!
1%
1-
12
#196580000000
0!
0%
b101 *
0-
02
b101 6
#196590000000
1!
1%
1-
12
#196600000000
0!
0%
b110 *
0-
02
b110 6
#196610000000
1!
1%
1-
12
#196620000000
0!
0%
b111 *
0-
02
b111 6
#196630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#196640000000
0!
0%
b0 *
0-
02
b0 6
#196650000000
1!
1%
1-
12
#196660000000
0!
0%
b1 *
0-
02
b1 6
#196670000000
1!
1%
1-
12
#196680000000
0!
0%
b10 *
0-
02
b10 6
#196690000000
1!
1%
1-
12
#196700000000
0!
0%
b11 *
0-
02
b11 6
#196710000000
1!
1%
1-
12
15
#196720000000
0!
0%
b100 *
0-
02
b100 6
#196730000000
1!
1%
1-
12
#196740000000
0!
0%
b101 *
0-
02
b101 6
#196750000000
1!
1%
1-
12
#196760000000
0!
0%
b110 *
0-
02
b110 6
#196770000000
1!
1%
1-
12
#196780000000
0!
0%
b111 *
0-
02
b111 6
#196790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#196800000000
0!
0%
b0 *
0-
02
b0 6
#196810000000
1!
1%
1-
12
#196820000000
0!
0%
b1 *
0-
02
b1 6
#196830000000
1!
1%
1-
12
#196840000000
0!
0%
b10 *
0-
02
b10 6
#196850000000
1!
1%
1-
12
#196860000000
0!
0%
b11 *
0-
02
b11 6
#196870000000
1!
1%
1-
12
15
#196880000000
0!
0%
b100 *
0-
02
b100 6
#196890000000
1!
1%
1-
12
#196900000000
0!
0%
b101 *
0-
02
b101 6
#196910000000
1!
1%
1-
12
#196920000000
0!
0%
b110 *
0-
02
b110 6
#196930000000
1!
1%
1-
12
#196940000000
0!
0%
b111 *
0-
02
b111 6
#196950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#196960000000
0!
0%
b0 *
0-
02
b0 6
#196970000000
1!
1%
1-
12
#196980000000
0!
0%
b1 *
0-
02
b1 6
#196990000000
1!
1%
1-
12
#197000000000
0!
0%
b10 *
0-
02
b10 6
#197010000000
1!
1%
1-
12
#197020000000
0!
0%
b11 *
0-
02
b11 6
#197030000000
1!
1%
1-
12
15
#197040000000
0!
0%
b100 *
0-
02
b100 6
#197050000000
1!
1%
1-
12
#197060000000
0!
0%
b101 *
0-
02
b101 6
#197070000000
1!
1%
1-
12
#197080000000
0!
0%
b110 *
0-
02
b110 6
#197090000000
1!
1%
1-
12
#197100000000
0!
0%
b111 *
0-
02
b111 6
#197110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#197120000000
0!
0%
b0 *
0-
02
b0 6
#197130000000
1!
1%
1-
12
#197140000000
0!
0%
b1 *
0-
02
b1 6
#197150000000
1!
1%
1-
12
#197160000000
0!
0%
b10 *
0-
02
b10 6
#197170000000
1!
1%
1-
12
#197180000000
0!
0%
b11 *
0-
02
b11 6
#197190000000
1!
1%
1-
12
15
#197200000000
0!
0%
b100 *
0-
02
b100 6
#197210000000
1!
1%
1-
12
#197220000000
0!
0%
b101 *
0-
02
b101 6
#197230000000
1!
1%
1-
12
#197240000000
0!
0%
b110 *
0-
02
b110 6
#197250000000
1!
1%
1-
12
#197260000000
0!
0%
b111 *
0-
02
b111 6
#197270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#197280000000
0!
0%
b0 *
0-
02
b0 6
#197290000000
1!
1%
1-
12
#197300000000
0!
0%
b1 *
0-
02
b1 6
#197310000000
1!
1%
1-
12
#197320000000
0!
0%
b10 *
0-
02
b10 6
#197330000000
1!
1%
1-
12
#197340000000
0!
0%
b11 *
0-
02
b11 6
#197350000000
1!
1%
1-
12
15
#197360000000
0!
0%
b100 *
0-
02
b100 6
#197370000000
1!
1%
1-
12
#197380000000
0!
0%
b101 *
0-
02
b101 6
#197390000000
1!
1%
1-
12
#197400000000
0!
0%
b110 *
0-
02
b110 6
#197410000000
1!
1%
1-
12
#197420000000
0!
0%
b111 *
0-
02
b111 6
#197430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#197440000000
0!
0%
b0 *
0-
02
b0 6
#197450000000
1!
1%
1-
12
#197460000000
0!
0%
b1 *
0-
02
b1 6
#197470000000
1!
1%
1-
12
#197480000000
0!
0%
b10 *
0-
02
b10 6
#197490000000
1!
1%
1-
12
#197500000000
0!
0%
b11 *
0-
02
b11 6
#197510000000
1!
1%
1-
12
15
#197520000000
0!
0%
b100 *
0-
02
b100 6
#197530000000
1!
1%
1-
12
#197540000000
0!
0%
b101 *
0-
02
b101 6
#197550000000
1!
1%
1-
12
#197560000000
0!
0%
b110 *
0-
02
b110 6
#197570000000
1!
1%
1-
12
#197580000000
0!
0%
b111 *
0-
02
b111 6
#197590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#197600000000
0!
0%
b0 *
0-
02
b0 6
#197610000000
1!
1%
1-
12
#197620000000
0!
0%
b1 *
0-
02
b1 6
#197630000000
1!
1%
1-
12
#197640000000
0!
0%
b10 *
0-
02
b10 6
#197650000000
1!
1%
1-
12
#197660000000
0!
0%
b11 *
0-
02
b11 6
#197670000000
1!
1%
1-
12
15
#197680000000
0!
0%
b100 *
0-
02
b100 6
#197690000000
1!
1%
1-
12
#197700000000
0!
0%
b101 *
0-
02
b101 6
#197710000000
1!
1%
1-
12
#197720000000
0!
0%
b110 *
0-
02
b110 6
#197730000000
1!
1%
1-
12
#197740000000
0!
0%
b111 *
0-
02
b111 6
#197750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#197760000000
0!
0%
b0 *
0-
02
b0 6
#197770000000
1!
1%
1-
12
#197780000000
0!
0%
b1 *
0-
02
b1 6
#197790000000
1!
1%
1-
12
#197800000000
0!
0%
b10 *
0-
02
b10 6
#197810000000
1!
1%
1-
12
#197820000000
0!
0%
b11 *
0-
02
b11 6
#197830000000
1!
1%
1-
12
15
#197840000000
0!
0%
b100 *
0-
02
b100 6
#197850000000
1!
1%
1-
12
#197860000000
0!
0%
b101 *
0-
02
b101 6
#197870000000
1!
1%
1-
12
#197880000000
0!
0%
b110 *
0-
02
b110 6
#197890000000
1!
1%
1-
12
#197900000000
0!
0%
b111 *
0-
02
b111 6
#197910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#197920000000
0!
0%
b0 *
0-
02
b0 6
#197930000000
1!
1%
1-
12
#197940000000
0!
0%
b1 *
0-
02
b1 6
#197950000000
1!
1%
1-
12
#197960000000
0!
0%
b10 *
0-
02
b10 6
#197970000000
1!
1%
1-
12
#197980000000
0!
0%
b11 *
0-
02
b11 6
#197990000000
1!
1%
1-
12
15
#198000000000
0!
0%
b100 *
0-
02
b100 6
#198010000000
1!
1%
1-
12
#198020000000
0!
0%
b101 *
0-
02
b101 6
#198030000000
1!
1%
1-
12
#198040000000
0!
0%
b110 *
0-
02
b110 6
#198050000000
1!
1%
1-
12
#198060000000
0!
0%
b111 *
0-
02
b111 6
#198070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#198080000000
0!
0%
b0 *
0-
02
b0 6
#198090000000
1!
1%
1-
12
#198100000000
0!
0%
b1 *
0-
02
b1 6
#198110000000
1!
1%
1-
12
#198120000000
0!
0%
b10 *
0-
02
b10 6
#198130000000
1!
1%
1-
12
#198140000000
0!
0%
b11 *
0-
02
b11 6
#198150000000
1!
1%
1-
12
15
#198160000000
0!
0%
b100 *
0-
02
b100 6
#198170000000
1!
1%
1-
12
#198180000000
0!
0%
b101 *
0-
02
b101 6
#198190000000
1!
1%
1-
12
#198200000000
0!
0%
b110 *
0-
02
b110 6
#198210000000
1!
1%
1-
12
#198220000000
0!
0%
b111 *
0-
02
b111 6
#198230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#198240000000
0!
0%
b0 *
0-
02
b0 6
#198250000000
1!
1%
1-
12
#198260000000
0!
0%
b1 *
0-
02
b1 6
#198270000000
1!
1%
1-
12
#198280000000
0!
0%
b10 *
0-
02
b10 6
#198290000000
1!
1%
1-
12
#198300000000
0!
0%
b11 *
0-
02
b11 6
#198310000000
1!
1%
1-
12
15
#198320000000
0!
0%
b100 *
0-
02
b100 6
#198330000000
1!
1%
1-
12
#198340000000
0!
0%
b101 *
0-
02
b101 6
#198350000000
1!
1%
1-
12
#198360000000
0!
0%
b110 *
0-
02
b110 6
#198370000000
1!
1%
1-
12
#198380000000
0!
0%
b111 *
0-
02
b111 6
#198390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#198400000000
0!
0%
b0 *
0-
02
b0 6
#198410000000
1!
1%
1-
12
#198420000000
0!
0%
b1 *
0-
02
b1 6
#198430000000
1!
1%
1-
12
#198440000000
0!
0%
b10 *
0-
02
b10 6
#198450000000
1!
1%
1-
12
#198460000000
0!
0%
b11 *
0-
02
b11 6
#198470000000
1!
1%
1-
12
15
#198480000000
0!
0%
b100 *
0-
02
b100 6
#198490000000
1!
1%
1-
12
#198500000000
0!
0%
b101 *
0-
02
b101 6
#198510000000
1!
1%
1-
12
#198520000000
0!
0%
b110 *
0-
02
b110 6
#198530000000
1!
1%
1-
12
#198540000000
0!
0%
b111 *
0-
02
b111 6
#198550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#198560000000
0!
0%
b0 *
0-
02
b0 6
#198570000000
1!
1%
1-
12
#198580000000
0!
0%
b1 *
0-
02
b1 6
#198590000000
1!
1%
1-
12
#198600000000
0!
0%
b10 *
0-
02
b10 6
#198610000000
1!
1%
1-
12
#198620000000
0!
0%
b11 *
0-
02
b11 6
#198630000000
1!
1%
1-
12
15
#198640000000
0!
0%
b100 *
0-
02
b100 6
#198650000000
1!
1%
1-
12
#198660000000
0!
0%
b101 *
0-
02
b101 6
#198670000000
1!
1%
1-
12
#198680000000
0!
0%
b110 *
0-
02
b110 6
#198690000000
1!
1%
1-
12
#198700000000
0!
0%
b111 *
0-
02
b111 6
#198710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#198720000000
0!
0%
b0 *
0-
02
b0 6
#198730000000
1!
1%
1-
12
#198740000000
0!
0%
b1 *
0-
02
b1 6
#198750000000
1!
1%
1-
12
#198760000000
0!
0%
b10 *
0-
02
b10 6
#198770000000
1!
1%
1-
12
#198780000000
0!
0%
b11 *
0-
02
b11 6
#198790000000
1!
1%
1-
12
15
#198800000000
0!
0%
b100 *
0-
02
b100 6
#198810000000
1!
1%
1-
12
#198820000000
0!
0%
b101 *
0-
02
b101 6
#198830000000
1!
1%
1-
12
#198840000000
0!
0%
b110 *
0-
02
b110 6
#198850000000
1!
1%
1-
12
#198860000000
0!
0%
b111 *
0-
02
b111 6
#198870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#198880000000
0!
0%
b0 *
0-
02
b0 6
#198890000000
1!
1%
1-
12
#198900000000
0!
0%
b1 *
0-
02
b1 6
#198910000000
1!
1%
1-
12
#198920000000
0!
0%
b10 *
0-
02
b10 6
#198930000000
1!
1%
1-
12
#198940000000
0!
0%
b11 *
0-
02
b11 6
#198950000000
1!
1%
1-
12
15
#198960000000
0!
0%
b100 *
0-
02
b100 6
#198970000000
1!
1%
1-
12
#198980000000
0!
0%
b101 *
0-
02
b101 6
#198990000000
1!
1%
1-
12
#199000000000
0!
0%
b110 *
0-
02
b110 6
#199010000000
1!
1%
1-
12
#199020000000
0!
0%
b111 *
0-
02
b111 6
#199030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#199040000000
0!
0%
b0 *
0-
02
b0 6
#199050000000
1!
1%
1-
12
#199060000000
0!
0%
b1 *
0-
02
b1 6
#199070000000
1!
1%
1-
12
#199080000000
0!
0%
b10 *
0-
02
b10 6
#199090000000
1!
1%
1-
12
#199100000000
0!
0%
b11 *
0-
02
b11 6
#199110000000
1!
1%
1-
12
15
#199120000000
0!
0%
b100 *
0-
02
b100 6
#199130000000
1!
1%
1-
12
#199140000000
0!
0%
b101 *
0-
02
b101 6
#199150000000
1!
1%
1-
12
#199160000000
0!
0%
b110 *
0-
02
b110 6
#199170000000
1!
1%
1-
12
#199180000000
0!
0%
b111 *
0-
02
b111 6
#199190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#199200000000
0!
0%
b0 *
0-
02
b0 6
#199210000000
1!
1%
1-
12
#199220000000
0!
0%
b1 *
0-
02
b1 6
#199230000000
1!
1%
1-
12
#199240000000
0!
0%
b10 *
0-
02
b10 6
#199250000000
1!
1%
1-
12
#199260000000
0!
0%
b11 *
0-
02
b11 6
#199270000000
1!
1%
1-
12
15
#199280000000
0!
0%
b100 *
0-
02
b100 6
#199290000000
1!
1%
1-
12
#199300000000
0!
0%
b101 *
0-
02
b101 6
#199310000000
1!
1%
1-
12
#199320000000
0!
0%
b110 *
0-
02
b110 6
#199330000000
1!
1%
1-
12
#199340000000
0!
0%
b111 *
0-
02
b111 6
#199350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#199360000000
0!
0%
b0 *
0-
02
b0 6
#199370000000
1!
1%
1-
12
#199380000000
0!
0%
b1 *
0-
02
b1 6
#199390000000
1!
1%
1-
12
#199400000000
0!
0%
b10 *
0-
02
b10 6
#199410000000
1!
1%
1-
12
#199420000000
0!
0%
b11 *
0-
02
b11 6
#199430000000
1!
1%
1-
12
15
#199440000000
0!
0%
b100 *
0-
02
b100 6
#199450000000
1!
1%
1-
12
#199460000000
0!
0%
b101 *
0-
02
b101 6
#199470000000
1!
1%
1-
12
#199480000000
0!
0%
b110 *
0-
02
b110 6
#199490000000
1!
1%
1-
12
#199500000000
0!
0%
b111 *
0-
02
b111 6
#199510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#199520000000
0!
0%
b0 *
0-
02
b0 6
#199530000000
1!
1%
1-
12
#199540000000
0!
0%
b1 *
0-
02
b1 6
#199550000000
1!
1%
1-
12
#199560000000
0!
0%
b10 *
0-
02
b10 6
#199570000000
1!
1%
1-
12
#199580000000
0!
0%
b11 *
0-
02
b11 6
#199590000000
1!
1%
1-
12
15
#199600000000
0!
0%
b100 *
0-
02
b100 6
#199610000000
1!
1%
1-
12
#199620000000
0!
0%
b101 *
0-
02
b101 6
#199630000000
1!
1%
1-
12
#199640000000
0!
0%
b110 *
0-
02
b110 6
#199650000000
1!
1%
1-
12
#199660000000
0!
0%
b111 *
0-
02
b111 6
#199670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#199680000000
0!
0%
b0 *
0-
02
b0 6
#199690000000
1!
1%
1-
12
#199700000000
0!
0%
b1 *
0-
02
b1 6
#199710000000
1!
1%
1-
12
#199720000000
0!
0%
b10 *
0-
02
b10 6
#199730000000
1!
1%
1-
12
#199740000000
0!
0%
b11 *
0-
02
b11 6
#199750000000
1!
1%
1-
12
15
#199760000000
0!
0%
b100 *
0-
02
b100 6
#199770000000
1!
1%
1-
12
#199780000000
0!
0%
b101 *
0-
02
b101 6
#199790000000
1!
1%
1-
12
#199800000000
0!
0%
b110 *
0-
02
b110 6
#199810000000
1!
1%
1-
12
#199820000000
0!
0%
b111 *
0-
02
b111 6
#199830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#199840000000
0!
0%
b0 *
0-
02
b0 6
#199850000000
1!
1%
1-
12
#199860000000
0!
0%
b1 *
0-
02
b1 6
#199870000000
1!
1%
1-
12
#199880000000
0!
0%
b10 *
0-
02
b10 6
#199890000000
1!
1%
1-
12
#199900000000
0!
0%
b11 *
0-
02
b11 6
#199910000000
1!
1%
1-
12
15
#199920000000
0!
0%
b100 *
0-
02
b100 6
#199930000000
1!
1%
1-
12
#199940000000
0!
0%
b101 *
0-
02
b101 6
#199950000000
1!
1%
1-
12
#199960000000
0!
0%
b110 *
0-
02
b110 6
#199970000000
1!
1%
1-
12
#199980000000
0!
0%
b111 *
0-
02
b111 6
#199990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#200000000000
0!
0%
b0 *
0-
02
b0 6
#200010000000
1!
1%
1-
12
#200020000000
0!
0%
b1 *
0-
02
b1 6
#200030000000
1!
1%
1-
12
#200040000000
0!
0%
b10 *
0-
02
b10 6
#200050000000
1!
1%
1-
12
#200060000000
0!
0%
b11 *
0-
02
b11 6
#200070000000
1!
1%
1-
12
15
#200080000000
0!
0%
b100 *
0-
02
b100 6
#200090000000
1!
1%
1-
12
#200100000000
0!
0%
b101 *
0-
02
b101 6
#200110000000
1!
1%
1-
12
#200120000000
0!
0%
b110 *
0-
02
b110 6
#200130000000
1!
1%
1-
12
#200140000000
0!
0%
b111 *
0-
02
b111 6
#200150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#200160000000
0!
0%
b0 *
0-
02
b0 6
#200170000000
1!
1%
1-
12
#200180000000
0!
0%
b1 *
0-
02
b1 6
#200190000000
1!
1%
1-
12
#200200000000
0!
0%
b10 *
0-
02
b10 6
#200210000000
1!
1%
1-
12
#200220000000
0!
0%
b11 *
0-
02
b11 6
#200230000000
1!
1%
1-
12
15
#200240000000
0!
0%
b100 *
0-
02
b100 6
#200250000000
1!
1%
1-
12
#200260000000
0!
0%
b101 *
0-
02
b101 6
#200270000000
1!
1%
1-
12
#200280000000
0!
0%
b110 *
0-
02
b110 6
#200290000000
1!
1%
1-
12
#200300000000
0!
0%
b111 *
0-
02
b111 6
#200310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#200320000000
0!
0%
b0 *
0-
02
b0 6
#200330000000
1!
1%
1-
12
#200340000000
0!
0%
b1 *
0-
02
b1 6
#200350000000
1!
1%
1-
12
#200360000000
0!
0%
b10 *
0-
02
b10 6
#200370000000
1!
1%
1-
12
#200380000000
0!
0%
b11 *
0-
02
b11 6
#200390000000
1!
1%
1-
12
15
#200400000000
0!
0%
b100 *
0-
02
b100 6
#200410000000
1!
1%
1-
12
#200420000000
0!
0%
b101 *
0-
02
b101 6
#200430000000
1!
1%
1-
12
#200440000000
0!
0%
b110 *
0-
02
b110 6
#200450000000
1!
1%
1-
12
#200460000000
0!
0%
b111 *
0-
02
b111 6
#200470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#200480000000
0!
0%
b0 *
0-
02
b0 6
#200490000000
1!
1%
1-
12
#200500000000
0!
0%
b1 *
0-
02
b1 6
#200510000000
1!
1%
1-
12
#200520000000
0!
0%
b10 *
0-
02
b10 6
#200530000000
1!
1%
1-
12
#200540000000
0!
0%
b11 *
0-
02
b11 6
#200550000000
1!
1%
1-
12
15
#200560000000
0!
0%
b100 *
0-
02
b100 6
#200570000000
1!
1%
1-
12
#200580000000
0!
0%
b101 *
0-
02
b101 6
#200590000000
1!
1%
1-
12
#200600000000
0!
0%
b110 *
0-
02
b110 6
#200610000000
1!
1%
1-
12
#200620000000
0!
0%
b111 *
0-
02
b111 6
#200630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#200640000000
0!
0%
b0 *
0-
02
b0 6
#200650000000
1!
1%
1-
12
#200660000000
0!
0%
b1 *
0-
02
b1 6
#200670000000
1!
1%
1-
12
#200680000000
0!
0%
b10 *
0-
02
b10 6
#200690000000
1!
1%
1-
12
#200700000000
0!
0%
b11 *
0-
02
b11 6
#200710000000
1!
1%
1-
12
15
#200720000000
0!
0%
b100 *
0-
02
b100 6
#200730000000
1!
1%
1-
12
#200740000000
0!
0%
b101 *
0-
02
b101 6
#200750000000
1!
1%
1-
12
#200760000000
0!
0%
b110 *
0-
02
b110 6
#200770000000
1!
1%
1-
12
#200780000000
0!
0%
b111 *
0-
02
b111 6
#200790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#200800000000
0!
0%
b0 *
0-
02
b0 6
#200810000000
1!
1%
1-
12
#200820000000
0!
0%
b1 *
0-
02
b1 6
#200830000000
1!
1%
1-
12
#200840000000
0!
0%
b10 *
0-
02
b10 6
#200850000000
1!
1%
1-
12
#200860000000
0!
0%
b11 *
0-
02
b11 6
#200870000000
1!
1%
1-
12
15
#200880000000
0!
0%
b100 *
0-
02
b100 6
#200890000000
1!
1%
1-
12
#200900000000
0!
0%
b101 *
0-
02
b101 6
#200910000000
1!
1%
1-
12
#200920000000
0!
0%
b110 *
0-
02
b110 6
#200930000000
1!
1%
1-
12
#200940000000
0!
0%
b111 *
0-
02
b111 6
#200950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#200960000000
0!
0%
b0 *
0-
02
b0 6
#200970000000
1!
1%
1-
12
#200980000000
0!
0%
b1 *
0-
02
b1 6
#200990000000
1!
1%
1-
12
#201000000000
0!
0%
b10 *
0-
02
b10 6
#201010000000
1!
1%
1-
12
#201020000000
0!
0%
b11 *
0-
02
b11 6
#201030000000
1!
1%
1-
12
15
#201040000000
0!
0%
b100 *
0-
02
b100 6
#201050000000
1!
1%
1-
12
#201060000000
0!
0%
b101 *
0-
02
b101 6
#201070000000
1!
1%
1-
12
#201080000000
0!
0%
b110 *
0-
02
b110 6
#201090000000
1!
1%
1-
12
#201100000000
0!
0%
b111 *
0-
02
b111 6
#201110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#201120000000
0!
0%
b0 *
0-
02
b0 6
#201130000000
1!
1%
1-
12
#201140000000
0!
0%
b1 *
0-
02
b1 6
#201150000000
1!
1%
1-
12
#201160000000
0!
0%
b10 *
0-
02
b10 6
#201170000000
1!
1%
1-
12
#201180000000
0!
0%
b11 *
0-
02
b11 6
#201190000000
1!
1%
1-
12
15
#201200000000
0!
0%
b100 *
0-
02
b100 6
#201210000000
1!
1%
1-
12
#201220000000
0!
0%
b101 *
0-
02
b101 6
#201230000000
1!
1%
1-
12
#201240000000
0!
0%
b110 *
0-
02
b110 6
#201250000000
1!
1%
1-
12
#201260000000
0!
0%
b111 *
0-
02
b111 6
#201270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#201280000000
0!
0%
b0 *
0-
02
b0 6
#201290000000
1!
1%
1-
12
#201300000000
0!
0%
b1 *
0-
02
b1 6
#201310000000
1!
1%
1-
12
#201320000000
0!
0%
b10 *
0-
02
b10 6
#201330000000
1!
1%
1-
12
#201340000000
0!
0%
b11 *
0-
02
b11 6
#201350000000
1!
1%
1-
12
15
#201360000000
0!
0%
b100 *
0-
02
b100 6
#201370000000
1!
1%
1-
12
#201380000000
0!
0%
b101 *
0-
02
b101 6
#201390000000
1!
1%
1-
12
#201400000000
0!
0%
b110 *
0-
02
b110 6
#201410000000
1!
1%
1-
12
#201420000000
0!
0%
b111 *
0-
02
b111 6
#201430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#201440000000
0!
0%
b0 *
0-
02
b0 6
#201450000000
1!
1%
1-
12
#201460000000
0!
0%
b1 *
0-
02
b1 6
#201470000000
1!
1%
1-
12
#201480000000
0!
0%
b10 *
0-
02
b10 6
#201490000000
1!
1%
1-
12
#201500000000
0!
0%
b11 *
0-
02
b11 6
#201510000000
1!
1%
1-
12
15
#201520000000
0!
0%
b100 *
0-
02
b100 6
#201530000000
1!
1%
1-
12
#201540000000
0!
0%
b101 *
0-
02
b101 6
#201550000000
1!
1%
1-
12
#201560000000
0!
0%
b110 *
0-
02
b110 6
#201570000000
1!
1%
1-
12
#201580000000
0!
0%
b111 *
0-
02
b111 6
#201590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#201600000000
0!
0%
b0 *
0-
02
b0 6
#201610000000
1!
1%
1-
12
#201620000000
0!
0%
b1 *
0-
02
b1 6
#201630000000
1!
1%
1-
12
#201640000000
0!
0%
b10 *
0-
02
b10 6
#201650000000
1!
1%
1-
12
#201660000000
0!
0%
b11 *
0-
02
b11 6
#201670000000
1!
1%
1-
12
15
#201680000000
0!
0%
b100 *
0-
02
b100 6
#201690000000
1!
1%
1-
12
#201700000000
0!
0%
b101 *
0-
02
b101 6
#201710000000
1!
1%
1-
12
#201720000000
0!
0%
b110 *
0-
02
b110 6
#201730000000
1!
1%
1-
12
#201740000000
0!
0%
b111 *
0-
02
b111 6
#201750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#201760000000
0!
0%
b0 *
0-
02
b0 6
#201770000000
1!
1%
1-
12
#201780000000
0!
0%
b1 *
0-
02
b1 6
#201790000000
1!
1%
1-
12
#201800000000
0!
0%
b10 *
0-
02
b10 6
#201810000000
1!
1%
1-
12
#201820000000
0!
0%
b11 *
0-
02
b11 6
#201830000000
1!
1%
1-
12
15
#201840000000
0!
0%
b100 *
0-
02
b100 6
#201850000000
1!
1%
1-
12
#201860000000
0!
0%
b101 *
0-
02
b101 6
#201870000000
1!
1%
1-
12
#201880000000
0!
0%
b110 *
0-
02
b110 6
#201890000000
1!
1%
1-
12
#201900000000
0!
0%
b111 *
0-
02
b111 6
#201910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#201920000000
0!
0%
b0 *
0-
02
b0 6
#201930000000
1!
1%
1-
12
#201940000000
0!
0%
b1 *
0-
02
b1 6
#201950000000
1!
1%
1-
12
#201960000000
0!
0%
b10 *
0-
02
b10 6
#201970000000
1!
1%
1-
12
#201980000000
0!
0%
b11 *
0-
02
b11 6
#201990000000
1!
1%
1-
12
15
#202000000000
0!
0%
b100 *
0-
02
b100 6
#202010000000
1!
1%
1-
12
#202020000000
0!
0%
b101 *
0-
02
b101 6
#202030000000
1!
1%
1-
12
#202040000000
0!
0%
b110 *
0-
02
b110 6
#202050000000
1!
1%
1-
12
#202060000000
0!
0%
b111 *
0-
02
b111 6
#202070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#202080000000
0!
0%
b0 *
0-
02
b0 6
#202090000000
1!
1%
1-
12
#202100000000
0!
0%
b1 *
0-
02
b1 6
#202110000000
1!
1%
1-
12
#202120000000
0!
0%
b10 *
0-
02
b10 6
#202130000000
1!
1%
1-
12
#202140000000
0!
0%
b11 *
0-
02
b11 6
#202150000000
1!
1%
1-
12
15
#202160000000
0!
0%
b100 *
0-
02
b100 6
#202170000000
1!
1%
1-
12
#202180000000
0!
0%
b101 *
0-
02
b101 6
#202190000000
1!
1%
1-
12
#202200000000
0!
0%
b110 *
0-
02
b110 6
#202210000000
1!
1%
1-
12
#202220000000
0!
0%
b111 *
0-
02
b111 6
#202230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#202240000000
0!
0%
b0 *
0-
02
b0 6
#202250000000
1!
1%
1-
12
#202260000000
0!
0%
b1 *
0-
02
b1 6
#202270000000
1!
1%
1-
12
#202280000000
0!
0%
b10 *
0-
02
b10 6
#202290000000
1!
1%
1-
12
#202300000000
0!
0%
b11 *
0-
02
b11 6
#202310000000
1!
1%
1-
12
15
#202320000000
0!
0%
b100 *
0-
02
b100 6
#202330000000
1!
1%
1-
12
#202340000000
0!
0%
b101 *
0-
02
b101 6
#202350000000
1!
1%
1-
12
#202360000000
0!
0%
b110 *
0-
02
b110 6
#202370000000
1!
1%
1-
12
#202380000000
0!
0%
b111 *
0-
02
b111 6
#202390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#202400000000
0!
0%
b0 *
0-
02
b0 6
#202410000000
1!
1%
1-
12
#202420000000
0!
0%
b1 *
0-
02
b1 6
#202430000000
1!
1%
1-
12
#202440000000
0!
0%
b10 *
0-
02
b10 6
#202450000000
1!
1%
1-
12
#202460000000
0!
0%
b11 *
0-
02
b11 6
#202470000000
1!
1%
1-
12
15
#202480000000
0!
0%
b100 *
0-
02
b100 6
#202490000000
1!
1%
1-
12
#202500000000
0!
0%
b101 *
0-
02
b101 6
#202510000000
1!
1%
1-
12
#202520000000
0!
0%
b110 *
0-
02
b110 6
#202530000000
1!
1%
1-
12
#202540000000
0!
0%
b111 *
0-
02
b111 6
#202550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#202560000000
0!
0%
b0 *
0-
02
b0 6
#202570000000
1!
1%
1-
12
#202580000000
0!
0%
b1 *
0-
02
b1 6
#202590000000
1!
1%
1-
12
#202600000000
0!
0%
b10 *
0-
02
b10 6
#202610000000
1!
1%
1-
12
#202620000000
0!
0%
b11 *
0-
02
b11 6
#202630000000
1!
1%
1-
12
15
#202640000000
0!
0%
b100 *
0-
02
b100 6
#202650000000
1!
1%
1-
12
#202660000000
0!
0%
b101 *
0-
02
b101 6
#202670000000
1!
1%
1-
12
#202680000000
0!
0%
b110 *
0-
02
b110 6
#202690000000
1!
1%
1-
12
#202700000000
0!
0%
b111 *
0-
02
b111 6
#202710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#202720000000
0!
0%
b0 *
0-
02
b0 6
#202730000000
1!
1%
1-
12
#202740000000
0!
0%
b1 *
0-
02
b1 6
#202750000000
1!
1%
1-
12
#202760000000
0!
0%
b10 *
0-
02
b10 6
#202770000000
1!
1%
1-
12
#202780000000
0!
0%
b11 *
0-
02
b11 6
#202790000000
1!
1%
1-
12
15
#202800000000
0!
0%
b100 *
0-
02
b100 6
#202810000000
1!
1%
1-
12
#202820000000
0!
0%
b101 *
0-
02
b101 6
#202830000000
1!
1%
1-
12
#202840000000
0!
0%
b110 *
0-
02
b110 6
#202850000000
1!
1%
1-
12
#202860000000
0!
0%
b111 *
0-
02
b111 6
#202870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#202880000000
0!
0%
b0 *
0-
02
b0 6
#202890000000
1!
1%
1-
12
#202900000000
0!
0%
b1 *
0-
02
b1 6
#202910000000
1!
1%
1-
12
#202920000000
0!
0%
b10 *
0-
02
b10 6
#202930000000
1!
1%
1-
12
#202940000000
0!
0%
b11 *
0-
02
b11 6
#202950000000
1!
1%
1-
12
15
#202960000000
0!
0%
b100 *
0-
02
b100 6
#202970000000
1!
1%
1-
12
#202980000000
0!
0%
b101 *
0-
02
b101 6
#202990000000
1!
1%
1-
12
#203000000000
0!
0%
b110 *
0-
02
b110 6
#203010000000
1!
1%
1-
12
#203020000000
0!
0%
b111 *
0-
02
b111 6
#203030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#203040000000
0!
0%
b0 *
0-
02
b0 6
#203050000000
1!
1%
1-
12
#203060000000
0!
0%
b1 *
0-
02
b1 6
#203070000000
1!
1%
1-
12
#203080000000
0!
0%
b10 *
0-
02
b10 6
#203090000000
1!
1%
1-
12
#203100000000
0!
0%
b11 *
0-
02
b11 6
#203110000000
1!
1%
1-
12
15
#203120000000
0!
0%
b100 *
0-
02
b100 6
#203130000000
1!
1%
1-
12
#203140000000
0!
0%
b101 *
0-
02
b101 6
#203150000000
1!
1%
1-
12
#203160000000
0!
0%
b110 *
0-
02
b110 6
#203170000000
1!
1%
1-
12
#203180000000
0!
0%
b111 *
0-
02
b111 6
#203190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#203200000000
0!
0%
b0 *
0-
02
b0 6
#203210000000
1!
1%
1-
12
#203220000000
0!
0%
b1 *
0-
02
b1 6
#203230000000
1!
1%
1-
12
#203240000000
0!
0%
b10 *
0-
02
b10 6
#203250000000
1!
1%
1-
12
#203260000000
0!
0%
b11 *
0-
02
b11 6
#203270000000
1!
1%
1-
12
15
#203280000000
0!
0%
b100 *
0-
02
b100 6
#203290000000
1!
1%
1-
12
#203300000000
0!
0%
b101 *
0-
02
b101 6
#203310000000
1!
1%
1-
12
#203320000000
0!
0%
b110 *
0-
02
b110 6
#203330000000
1!
1%
1-
12
#203340000000
0!
0%
b111 *
0-
02
b111 6
#203350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#203360000000
0!
0%
b0 *
0-
02
b0 6
#203370000000
1!
1%
1-
12
#203380000000
0!
0%
b1 *
0-
02
b1 6
#203390000000
1!
1%
1-
12
#203400000000
0!
0%
b10 *
0-
02
b10 6
#203410000000
1!
1%
1-
12
#203420000000
0!
0%
b11 *
0-
02
b11 6
#203430000000
1!
1%
1-
12
15
#203440000000
0!
0%
b100 *
0-
02
b100 6
#203450000000
1!
1%
1-
12
#203460000000
0!
0%
b101 *
0-
02
b101 6
#203470000000
1!
1%
1-
12
#203480000000
0!
0%
b110 *
0-
02
b110 6
#203490000000
1!
1%
1-
12
#203500000000
0!
0%
b111 *
0-
02
b111 6
#203510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#203520000000
0!
0%
b0 *
0-
02
b0 6
#203530000000
1!
1%
1-
12
#203540000000
0!
0%
b1 *
0-
02
b1 6
#203550000000
1!
1%
1-
12
#203560000000
0!
0%
b10 *
0-
02
b10 6
#203570000000
1!
1%
1-
12
#203580000000
0!
0%
b11 *
0-
02
b11 6
#203590000000
1!
1%
1-
12
15
#203600000000
0!
0%
b100 *
0-
02
b100 6
#203610000000
1!
1%
1-
12
#203620000000
0!
0%
b101 *
0-
02
b101 6
#203630000000
1!
1%
1-
12
#203640000000
0!
0%
b110 *
0-
02
b110 6
#203650000000
1!
1%
1-
12
#203660000000
0!
0%
b111 *
0-
02
b111 6
#203670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#203680000000
0!
0%
b0 *
0-
02
b0 6
#203690000000
1!
1%
1-
12
#203700000000
0!
0%
b1 *
0-
02
b1 6
#203710000000
1!
1%
1-
12
#203720000000
0!
0%
b10 *
0-
02
b10 6
#203730000000
1!
1%
1-
12
#203740000000
0!
0%
b11 *
0-
02
b11 6
#203750000000
1!
1%
1-
12
15
#203760000000
0!
0%
b100 *
0-
02
b100 6
#203770000000
1!
1%
1-
12
#203780000000
0!
0%
b101 *
0-
02
b101 6
#203790000000
1!
1%
1-
12
#203800000000
0!
0%
b110 *
0-
02
b110 6
#203810000000
1!
1%
1-
12
#203820000000
0!
0%
b111 *
0-
02
b111 6
#203830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#203840000000
0!
0%
b0 *
0-
02
b0 6
#203850000000
1!
1%
1-
12
#203860000000
0!
0%
b1 *
0-
02
b1 6
#203870000000
1!
1%
1-
12
#203880000000
0!
0%
b10 *
0-
02
b10 6
#203890000000
1!
1%
1-
12
#203900000000
0!
0%
b11 *
0-
02
b11 6
#203910000000
1!
1%
1-
12
15
#203920000000
0!
0%
b100 *
0-
02
b100 6
#203930000000
1!
1%
1-
12
#203940000000
0!
0%
b101 *
0-
02
b101 6
#203950000000
1!
1%
1-
12
#203960000000
0!
0%
b110 *
0-
02
b110 6
#203970000000
1!
1%
1-
12
#203980000000
0!
0%
b111 *
0-
02
b111 6
#203990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#204000000000
0!
0%
b0 *
0-
02
b0 6
#204010000000
1!
1%
1-
12
#204020000000
0!
0%
b1 *
0-
02
b1 6
#204030000000
1!
1%
1-
12
#204040000000
0!
0%
b10 *
0-
02
b10 6
#204050000000
1!
1%
1-
12
#204060000000
0!
0%
b11 *
0-
02
b11 6
#204070000000
1!
1%
1-
12
15
#204080000000
0!
0%
b100 *
0-
02
b100 6
#204090000000
1!
1%
1-
12
#204100000000
0!
0%
b101 *
0-
02
b101 6
#204110000000
1!
1%
1-
12
#204120000000
0!
0%
b110 *
0-
02
b110 6
#204130000000
1!
1%
1-
12
#204140000000
0!
0%
b111 *
0-
02
b111 6
#204150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#204160000000
0!
0%
b0 *
0-
02
b0 6
#204170000000
1!
1%
1-
12
#204180000000
0!
0%
b1 *
0-
02
b1 6
#204190000000
1!
1%
1-
12
#204200000000
0!
0%
b10 *
0-
02
b10 6
#204210000000
1!
1%
1-
12
#204220000000
0!
0%
b11 *
0-
02
b11 6
#204230000000
1!
1%
1-
12
15
#204240000000
0!
0%
b100 *
0-
02
b100 6
#204250000000
1!
1%
1-
12
#204260000000
0!
0%
b101 *
0-
02
b101 6
#204270000000
1!
1%
1-
12
#204280000000
0!
0%
b110 *
0-
02
b110 6
#204290000000
1!
1%
1-
12
#204300000000
0!
0%
b111 *
0-
02
b111 6
#204310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#204320000000
0!
0%
b0 *
0-
02
b0 6
#204330000000
1!
1%
1-
12
#204340000000
0!
0%
b1 *
0-
02
b1 6
#204350000000
1!
1%
1-
12
#204360000000
0!
0%
b10 *
0-
02
b10 6
#204370000000
1!
1%
1-
12
#204380000000
0!
0%
b11 *
0-
02
b11 6
#204390000000
1!
1%
1-
12
15
#204400000000
0!
0%
b100 *
0-
02
b100 6
#204410000000
1!
1%
1-
12
#204420000000
0!
0%
b101 *
0-
02
b101 6
#204430000000
1!
1%
1-
12
#204440000000
0!
0%
b110 *
0-
02
b110 6
#204450000000
1!
1%
1-
12
#204460000000
0!
0%
b111 *
0-
02
b111 6
#204470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#204480000000
0!
0%
b0 *
0-
02
b0 6
#204490000000
1!
1%
1-
12
#204500000000
0!
0%
b1 *
0-
02
b1 6
#204510000000
1!
1%
1-
12
#204520000000
0!
0%
b10 *
0-
02
b10 6
#204530000000
1!
1%
1-
12
#204540000000
0!
0%
b11 *
0-
02
b11 6
#204550000000
1!
1%
1-
12
15
#204560000000
0!
0%
b100 *
0-
02
b100 6
#204570000000
1!
1%
1-
12
#204580000000
0!
0%
b101 *
0-
02
b101 6
#204590000000
1!
1%
1-
12
#204600000000
0!
0%
b110 *
0-
02
b110 6
#204610000000
1!
1%
1-
12
#204620000000
0!
0%
b111 *
0-
02
b111 6
#204630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#204640000000
0!
0%
b0 *
0-
02
b0 6
#204650000000
1!
1%
1-
12
#204660000000
0!
0%
b1 *
0-
02
b1 6
#204670000000
1!
1%
1-
12
#204680000000
0!
0%
b10 *
0-
02
b10 6
#204690000000
1!
1%
1-
12
#204700000000
0!
0%
b11 *
0-
02
b11 6
#204710000000
1!
1%
1-
12
15
#204720000000
0!
0%
b100 *
0-
02
b100 6
#204730000000
1!
1%
1-
12
#204740000000
0!
0%
b101 *
0-
02
b101 6
#204750000000
1!
1%
1-
12
#204760000000
0!
0%
b110 *
0-
02
b110 6
#204770000000
1!
1%
1-
12
#204780000000
0!
0%
b111 *
0-
02
b111 6
#204790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#204800000000
0!
0%
b0 *
0-
02
b0 6
#204810000000
1!
1%
1-
12
#204820000000
0!
0%
b1 *
0-
02
b1 6
#204830000000
1!
1%
1-
12
#204840000000
0!
0%
b10 *
0-
02
b10 6
#204850000000
1!
1%
1-
12
#204860000000
0!
0%
b11 *
0-
02
b11 6
#204870000000
1!
1%
1-
12
15
#204880000000
0!
0%
b100 *
0-
02
b100 6
#204890000000
1!
1%
1-
12
#204900000000
0!
0%
b101 *
0-
02
b101 6
#204910000000
1!
1%
1-
12
#204920000000
0!
0%
b110 *
0-
02
b110 6
#204930000000
1!
1%
1-
12
#204940000000
0!
0%
b111 *
0-
02
b111 6
#204950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#204960000000
0!
0%
b0 *
0-
02
b0 6
#204970000000
1!
1%
1-
12
#204980000000
0!
0%
b1 *
0-
02
b1 6
#204990000000
1!
1%
1-
12
#205000000000
0!
0%
b10 *
0-
02
b10 6
#205010000000
1!
1%
1-
12
#205020000000
0!
0%
b11 *
0-
02
b11 6
#205030000000
1!
1%
1-
12
15
#205040000000
0!
0%
b100 *
0-
02
b100 6
#205050000000
1!
1%
1-
12
#205060000000
0!
0%
b101 *
0-
02
b101 6
#205070000000
1!
1%
1-
12
#205080000000
0!
0%
b110 *
0-
02
b110 6
#205090000000
1!
1%
1-
12
#205100000000
0!
0%
b111 *
0-
02
b111 6
#205110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#205120000000
0!
0%
b0 *
0-
02
b0 6
#205130000000
1!
1%
1-
12
#205140000000
0!
0%
b1 *
0-
02
b1 6
#205150000000
1!
1%
1-
12
#205160000000
0!
0%
b10 *
0-
02
b10 6
#205170000000
1!
1%
1-
12
#205180000000
0!
0%
b11 *
0-
02
b11 6
#205190000000
1!
1%
1-
12
15
#205200000000
0!
0%
b100 *
0-
02
b100 6
#205210000000
1!
1%
1-
12
#205220000000
0!
0%
b101 *
0-
02
b101 6
#205230000000
1!
1%
1-
12
#205240000000
0!
0%
b110 *
0-
02
b110 6
#205250000000
1!
1%
1-
12
#205260000000
0!
0%
b111 *
0-
02
b111 6
#205270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#205280000000
0!
0%
b0 *
0-
02
b0 6
#205290000000
1!
1%
1-
12
#205300000000
0!
0%
b1 *
0-
02
b1 6
#205310000000
1!
1%
1-
12
#205320000000
0!
0%
b10 *
0-
02
b10 6
#205330000000
1!
1%
1-
12
#205340000000
0!
0%
b11 *
0-
02
b11 6
#205350000000
1!
1%
1-
12
15
#205360000000
0!
0%
b100 *
0-
02
b100 6
#205370000000
1!
1%
1-
12
#205380000000
0!
0%
b101 *
0-
02
b101 6
#205390000000
1!
1%
1-
12
#205400000000
0!
0%
b110 *
0-
02
b110 6
#205410000000
1!
1%
1-
12
#205420000000
0!
0%
b111 *
0-
02
b111 6
#205430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#205440000000
0!
0%
b0 *
0-
02
b0 6
#205450000000
1!
1%
1-
12
#205460000000
0!
0%
b1 *
0-
02
b1 6
#205470000000
1!
1%
1-
12
#205480000000
0!
0%
b10 *
0-
02
b10 6
#205490000000
1!
1%
1-
12
#205500000000
0!
0%
b11 *
0-
02
b11 6
#205510000000
1!
1%
1-
12
15
#205520000000
0!
0%
b100 *
0-
02
b100 6
#205530000000
1!
1%
1-
12
#205540000000
0!
0%
b101 *
0-
02
b101 6
#205550000000
1!
1%
1-
12
#205560000000
0!
0%
b110 *
0-
02
b110 6
#205570000000
1!
1%
1-
12
#205580000000
0!
0%
b111 *
0-
02
b111 6
#205590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#205600000000
0!
0%
b0 *
0-
02
b0 6
#205610000000
1!
1%
1-
12
#205620000000
0!
0%
b1 *
0-
02
b1 6
#205630000000
1!
1%
1-
12
#205640000000
0!
0%
b10 *
0-
02
b10 6
#205650000000
1!
1%
1-
12
#205660000000
0!
0%
b11 *
0-
02
b11 6
#205670000000
1!
1%
1-
12
15
#205680000000
0!
0%
b100 *
0-
02
b100 6
#205690000000
1!
1%
1-
12
#205700000000
0!
0%
b101 *
0-
02
b101 6
#205710000000
1!
1%
1-
12
#205720000000
0!
0%
b110 *
0-
02
b110 6
#205730000000
1!
1%
1-
12
#205740000000
0!
0%
b111 *
0-
02
b111 6
#205750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#205760000000
0!
0%
b0 *
0-
02
b0 6
#205770000000
1!
1%
1-
12
#205780000000
0!
0%
b1 *
0-
02
b1 6
#205790000000
1!
1%
1-
12
#205800000000
0!
0%
b10 *
0-
02
b10 6
#205810000000
1!
1%
1-
12
#205820000000
0!
0%
b11 *
0-
02
b11 6
#205830000000
1!
1%
1-
12
15
#205840000000
0!
0%
b100 *
0-
02
b100 6
#205850000000
1!
1%
1-
12
#205860000000
0!
0%
b101 *
0-
02
b101 6
#205870000000
1!
1%
1-
12
#205880000000
0!
0%
b110 *
0-
02
b110 6
#205890000000
1!
1%
1-
12
#205900000000
0!
0%
b111 *
0-
02
b111 6
#205910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#205920000000
0!
0%
b0 *
0-
02
b0 6
#205930000000
1!
1%
1-
12
#205940000000
0!
0%
b1 *
0-
02
b1 6
#205950000000
1!
1%
1-
12
#205960000000
0!
0%
b10 *
0-
02
b10 6
#205970000000
1!
1%
1-
12
#205980000000
0!
0%
b11 *
0-
02
b11 6
#205990000000
1!
1%
1-
12
15
#206000000000
0!
0%
b100 *
0-
02
b100 6
#206010000000
1!
1%
1-
12
#206020000000
0!
0%
b101 *
0-
02
b101 6
#206030000000
1!
1%
1-
12
#206040000000
0!
0%
b110 *
0-
02
b110 6
#206050000000
1!
1%
1-
12
#206060000000
0!
0%
b111 *
0-
02
b111 6
#206070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#206080000000
0!
0%
b0 *
0-
02
b0 6
#206090000000
1!
1%
1-
12
#206100000000
0!
0%
b1 *
0-
02
b1 6
#206110000000
1!
1%
1-
12
#206120000000
0!
0%
b10 *
0-
02
b10 6
#206130000000
1!
1%
1-
12
#206140000000
0!
0%
b11 *
0-
02
b11 6
#206150000000
1!
1%
1-
12
15
#206160000000
0!
0%
b100 *
0-
02
b100 6
#206170000000
1!
1%
1-
12
#206180000000
0!
0%
b101 *
0-
02
b101 6
#206190000000
1!
1%
1-
12
#206200000000
0!
0%
b110 *
0-
02
b110 6
#206210000000
1!
1%
1-
12
#206220000000
0!
0%
b111 *
0-
02
b111 6
#206230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#206240000000
0!
0%
b0 *
0-
02
b0 6
#206250000000
1!
1%
1-
12
#206260000000
0!
0%
b1 *
0-
02
b1 6
#206270000000
1!
1%
1-
12
#206280000000
0!
0%
b10 *
0-
02
b10 6
#206290000000
1!
1%
1-
12
#206300000000
0!
0%
b11 *
0-
02
b11 6
#206310000000
1!
1%
1-
12
15
#206320000000
0!
0%
b100 *
0-
02
b100 6
#206330000000
1!
1%
1-
12
#206340000000
0!
0%
b101 *
0-
02
b101 6
#206350000000
1!
1%
1-
12
#206360000000
0!
0%
b110 *
0-
02
b110 6
#206370000000
1!
1%
1-
12
#206380000000
0!
0%
b111 *
0-
02
b111 6
#206390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#206400000000
0!
0%
b0 *
0-
02
b0 6
#206410000000
1!
1%
1-
12
#206420000000
0!
0%
b1 *
0-
02
b1 6
#206430000000
1!
1%
1-
12
#206440000000
0!
0%
b10 *
0-
02
b10 6
#206450000000
1!
1%
1-
12
#206460000000
0!
0%
b11 *
0-
02
b11 6
#206470000000
1!
1%
1-
12
15
#206480000000
0!
0%
b100 *
0-
02
b100 6
#206490000000
1!
1%
1-
12
#206500000000
0!
0%
b101 *
0-
02
b101 6
#206510000000
1!
1%
1-
12
#206520000000
0!
0%
b110 *
0-
02
b110 6
#206530000000
1!
1%
1-
12
#206540000000
0!
0%
b111 *
0-
02
b111 6
#206550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#206560000000
0!
0%
b0 *
0-
02
b0 6
#206570000000
1!
1%
1-
12
#206580000000
0!
0%
b1 *
0-
02
b1 6
#206590000000
1!
1%
1-
12
#206600000000
0!
0%
b10 *
0-
02
b10 6
#206610000000
1!
1%
1-
12
#206620000000
0!
0%
b11 *
0-
02
b11 6
#206630000000
1!
1%
1-
12
15
#206640000000
0!
0%
b100 *
0-
02
b100 6
#206650000000
1!
1%
1-
12
#206660000000
0!
0%
b101 *
0-
02
b101 6
#206670000000
1!
1%
1-
12
#206680000000
0!
0%
b110 *
0-
02
b110 6
#206690000000
1!
1%
1-
12
#206700000000
0!
0%
b111 *
0-
02
b111 6
#206710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#206720000000
0!
0%
b0 *
0-
02
b0 6
#206730000000
1!
1%
1-
12
#206740000000
0!
0%
b1 *
0-
02
b1 6
#206750000000
1!
1%
1-
12
#206760000000
0!
0%
b10 *
0-
02
b10 6
#206770000000
1!
1%
1-
12
#206780000000
0!
0%
b11 *
0-
02
b11 6
#206790000000
1!
1%
1-
12
15
#206800000000
0!
0%
b100 *
0-
02
b100 6
#206810000000
1!
1%
1-
12
#206820000000
0!
0%
b101 *
0-
02
b101 6
#206830000000
1!
1%
1-
12
#206840000000
0!
0%
b110 *
0-
02
b110 6
#206850000000
1!
1%
1-
12
#206860000000
0!
0%
b111 *
0-
02
b111 6
#206870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#206880000000
0!
0%
b0 *
0-
02
b0 6
#206890000000
1!
1%
1-
12
#206900000000
0!
0%
b1 *
0-
02
b1 6
#206910000000
1!
1%
1-
12
#206920000000
0!
0%
b10 *
0-
02
b10 6
#206930000000
1!
1%
1-
12
#206940000000
0!
0%
b11 *
0-
02
b11 6
#206950000000
1!
1%
1-
12
15
#206960000000
0!
0%
b100 *
0-
02
b100 6
#206970000000
1!
1%
1-
12
#206980000000
0!
0%
b101 *
0-
02
b101 6
#206990000000
1!
1%
1-
12
#207000000000
0!
0%
b110 *
0-
02
b110 6
#207010000000
1!
1%
1-
12
#207020000000
0!
0%
b111 *
0-
02
b111 6
#207030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#207040000000
0!
0%
b0 *
0-
02
b0 6
#207050000000
1!
1%
1-
12
#207060000000
0!
0%
b1 *
0-
02
b1 6
#207070000000
1!
1%
1-
12
#207080000000
0!
0%
b10 *
0-
02
b10 6
#207090000000
1!
1%
1-
12
#207100000000
0!
0%
b11 *
0-
02
b11 6
#207110000000
1!
1%
1-
12
15
#207120000000
0!
0%
b100 *
0-
02
b100 6
#207130000000
1!
1%
1-
12
#207140000000
0!
0%
b101 *
0-
02
b101 6
#207150000000
1!
1%
1-
12
#207160000000
0!
0%
b110 *
0-
02
b110 6
#207170000000
1!
1%
1-
12
#207180000000
0!
0%
b111 *
0-
02
b111 6
#207190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#207200000000
0!
0%
b0 *
0-
02
b0 6
#207210000000
1!
1%
1-
12
#207220000000
0!
0%
b1 *
0-
02
b1 6
#207230000000
1!
1%
1-
12
#207240000000
0!
0%
b10 *
0-
02
b10 6
#207250000000
1!
1%
1-
12
#207260000000
0!
0%
b11 *
0-
02
b11 6
#207270000000
1!
1%
1-
12
15
#207280000000
0!
0%
b100 *
0-
02
b100 6
#207290000000
1!
1%
1-
12
#207300000000
0!
0%
b101 *
0-
02
b101 6
#207310000000
1!
1%
1-
12
#207320000000
0!
0%
b110 *
0-
02
b110 6
#207330000000
1!
1%
1-
12
#207340000000
0!
0%
b111 *
0-
02
b111 6
#207350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#207360000000
0!
0%
b0 *
0-
02
b0 6
#207370000000
1!
1%
1-
12
#207380000000
0!
0%
b1 *
0-
02
b1 6
#207390000000
1!
1%
1-
12
#207400000000
0!
0%
b10 *
0-
02
b10 6
#207410000000
1!
1%
1-
12
#207420000000
0!
0%
b11 *
0-
02
b11 6
#207430000000
1!
1%
1-
12
15
#207440000000
0!
0%
b100 *
0-
02
b100 6
#207450000000
1!
1%
1-
12
#207460000000
0!
0%
b101 *
0-
02
b101 6
#207470000000
1!
1%
1-
12
#207480000000
0!
0%
b110 *
0-
02
b110 6
#207490000000
1!
1%
1-
12
#207500000000
0!
0%
b111 *
0-
02
b111 6
#207510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#207520000000
0!
0%
b0 *
0-
02
b0 6
#207530000000
1!
1%
1-
12
#207540000000
0!
0%
b1 *
0-
02
b1 6
#207550000000
1!
1%
1-
12
#207560000000
0!
0%
b10 *
0-
02
b10 6
#207570000000
1!
1%
1-
12
#207580000000
0!
0%
b11 *
0-
02
b11 6
#207590000000
1!
1%
1-
12
15
#207600000000
0!
0%
b100 *
0-
02
b100 6
#207610000000
1!
1%
1-
12
#207620000000
0!
0%
b101 *
0-
02
b101 6
#207630000000
1!
1%
1-
12
#207640000000
0!
0%
b110 *
0-
02
b110 6
#207650000000
1!
1%
1-
12
#207660000000
0!
0%
b111 *
0-
02
b111 6
#207670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#207680000000
0!
0%
b0 *
0-
02
b0 6
#207690000000
1!
1%
1-
12
#207700000000
0!
0%
b1 *
0-
02
b1 6
#207710000000
1!
1%
1-
12
#207720000000
0!
0%
b10 *
0-
02
b10 6
#207730000000
1!
1%
1-
12
#207740000000
0!
0%
b11 *
0-
02
b11 6
#207750000000
1!
1%
1-
12
15
#207760000000
0!
0%
b100 *
0-
02
b100 6
#207770000000
1!
1%
1-
12
#207780000000
0!
0%
b101 *
0-
02
b101 6
#207790000000
1!
1%
1-
12
#207800000000
0!
0%
b110 *
0-
02
b110 6
#207810000000
1!
1%
1-
12
#207820000000
0!
0%
b111 *
0-
02
b111 6
#207830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#207840000000
0!
0%
b0 *
0-
02
b0 6
#207850000000
1!
1%
1-
12
#207860000000
0!
0%
b1 *
0-
02
b1 6
#207870000000
1!
1%
1-
12
#207880000000
0!
0%
b10 *
0-
02
b10 6
#207890000000
1!
1%
1-
12
#207900000000
0!
0%
b11 *
0-
02
b11 6
#207910000000
1!
1%
1-
12
15
#207920000000
0!
0%
b100 *
0-
02
b100 6
#207930000000
1!
1%
1-
12
#207940000000
0!
0%
b101 *
0-
02
b101 6
#207950000000
1!
1%
1-
12
#207960000000
0!
0%
b110 *
0-
02
b110 6
#207970000000
1!
1%
1-
12
#207980000000
0!
0%
b111 *
0-
02
b111 6
#207990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#208000000000
0!
0%
b0 *
0-
02
b0 6
#208010000000
1!
1%
1-
12
#208020000000
0!
0%
b1 *
0-
02
b1 6
#208030000000
1!
1%
1-
12
#208040000000
0!
0%
b10 *
0-
02
b10 6
#208050000000
1!
1%
1-
12
#208060000000
0!
0%
b11 *
0-
02
b11 6
#208070000000
1!
1%
1-
12
15
#208080000000
0!
0%
b100 *
0-
02
b100 6
#208090000000
1!
1%
1-
12
#208100000000
0!
0%
b101 *
0-
02
b101 6
#208110000000
1!
1%
1-
12
#208120000000
0!
0%
b110 *
0-
02
b110 6
#208130000000
1!
1%
1-
12
#208140000000
0!
0%
b111 *
0-
02
b111 6
#208150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#208160000000
0!
0%
b0 *
0-
02
b0 6
#208170000000
1!
1%
1-
12
#208180000000
0!
0%
b1 *
0-
02
b1 6
#208190000000
1!
1%
1-
12
#208200000000
0!
0%
b10 *
0-
02
b10 6
#208210000000
1!
1%
1-
12
#208220000000
0!
0%
b11 *
0-
02
b11 6
#208230000000
1!
1%
1-
12
15
#208240000000
0!
0%
b100 *
0-
02
b100 6
#208250000000
1!
1%
1-
12
#208260000000
0!
0%
b101 *
0-
02
b101 6
#208270000000
1!
1%
1-
12
#208280000000
0!
0%
b110 *
0-
02
b110 6
#208290000000
1!
1%
1-
12
#208300000000
0!
0%
b111 *
0-
02
b111 6
#208310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#208320000000
0!
0%
b0 *
0-
02
b0 6
#208330000000
1!
1%
1-
12
#208340000000
0!
0%
b1 *
0-
02
b1 6
#208350000000
1!
1%
1-
12
#208360000000
0!
0%
b10 *
0-
02
b10 6
#208370000000
1!
1%
1-
12
#208380000000
0!
0%
b11 *
0-
02
b11 6
#208390000000
1!
1%
1-
12
15
#208400000000
0!
0%
b100 *
0-
02
b100 6
#208410000000
1!
1%
1-
12
#208420000000
0!
0%
b101 *
0-
02
b101 6
#208430000000
1!
1%
1-
12
#208440000000
0!
0%
b110 *
0-
02
b110 6
#208450000000
1!
1%
1-
12
#208460000000
0!
0%
b111 *
0-
02
b111 6
#208470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#208480000000
0!
0%
b0 *
0-
02
b0 6
#208490000000
1!
1%
1-
12
#208500000000
0!
0%
b1 *
0-
02
b1 6
#208510000000
1!
1%
1-
12
#208520000000
0!
0%
b10 *
0-
02
b10 6
#208530000000
1!
1%
1-
12
#208540000000
0!
0%
b11 *
0-
02
b11 6
#208550000000
1!
1%
1-
12
15
#208560000000
0!
0%
b100 *
0-
02
b100 6
#208570000000
1!
1%
1-
12
#208580000000
0!
0%
b101 *
0-
02
b101 6
#208590000000
1!
1%
1-
12
#208600000000
0!
0%
b110 *
0-
02
b110 6
#208610000000
1!
1%
1-
12
#208620000000
0!
0%
b111 *
0-
02
b111 6
#208630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#208640000000
0!
0%
b0 *
0-
02
b0 6
#208650000000
1!
1%
1-
12
#208660000000
0!
0%
b1 *
0-
02
b1 6
#208670000000
1!
1%
1-
12
#208680000000
0!
0%
b10 *
0-
02
b10 6
#208690000000
1!
1%
1-
12
#208700000000
0!
0%
b11 *
0-
02
b11 6
#208710000000
1!
1%
1-
12
15
#208720000000
0!
0%
b100 *
0-
02
b100 6
#208730000000
1!
1%
1-
12
#208740000000
0!
0%
b101 *
0-
02
b101 6
#208750000000
1!
1%
1-
12
#208760000000
0!
0%
b110 *
0-
02
b110 6
#208770000000
1!
1%
1-
12
#208780000000
0!
0%
b111 *
0-
02
b111 6
#208790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#208800000000
0!
0%
b0 *
0-
02
b0 6
#208810000000
1!
1%
1-
12
#208820000000
0!
0%
b1 *
0-
02
b1 6
#208830000000
1!
1%
1-
12
#208840000000
0!
0%
b10 *
0-
02
b10 6
#208850000000
1!
1%
1-
12
#208860000000
0!
0%
b11 *
0-
02
b11 6
#208870000000
1!
1%
1-
12
15
#208880000000
0!
0%
b100 *
0-
02
b100 6
#208890000000
1!
1%
1-
12
#208900000000
0!
0%
b101 *
0-
02
b101 6
#208910000000
1!
1%
1-
12
#208920000000
0!
0%
b110 *
0-
02
b110 6
#208930000000
1!
1%
1-
12
#208940000000
0!
0%
b111 *
0-
02
b111 6
#208950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#208960000000
0!
0%
b0 *
0-
02
b0 6
#208970000000
1!
1%
1-
12
#208980000000
0!
0%
b1 *
0-
02
b1 6
#208990000000
1!
1%
1-
12
#209000000000
0!
0%
b10 *
0-
02
b10 6
#209010000000
1!
1%
1-
12
#209020000000
0!
0%
b11 *
0-
02
b11 6
#209030000000
1!
1%
1-
12
15
#209040000000
0!
0%
b100 *
0-
02
b100 6
#209050000000
1!
1%
1-
12
#209060000000
0!
0%
b101 *
0-
02
b101 6
#209070000000
1!
1%
1-
12
#209080000000
0!
0%
b110 *
0-
02
b110 6
#209090000000
1!
1%
1-
12
#209100000000
0!
0%
b111 *
0-
02
b111 6
#209110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#209120000000
0!
0%
b0 *
0-
02
b0 6
#209130000000
1!
1%
1-
12
#209140000000
0!
0%
b1 *
0-
02
b1 6
#209150000000
1!
1%
1-
12
#209160000000
0!
0%
b10 *
0-
02
b10 6
#209170000000
1!
1%
1-
12
#209180000000
0!
0%
b11 *
0-
02
b11 6
#209190000000
1!
1%
1-
12
15
#209200000000
0!
0%
b100 *
0-
02
b100 6
#209210000000
1!
1%
1-
12
#209220000000
0!
0%
b101 *
0-
02
b101 6
#209230000000
1!
1%
1-
12
#209240000000
0!
0%
b110 *
0-
02
b110 6
#209250000000
1!
1%
1-
12
#209260000000
0!
0%
b111 *
0-
02
b111 6
#209270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#209280000000
0!
0%
b0 *
0-
02
b0 6
#209290000000
1!
1%
1-
12
#209300000000
0!
0%
b1 *
0-
02
b1 6
#209310000000
1!
1%
1-
12
#209320000000
0!
0%
b10 *
0-
02
b10 6
#209330000000
1!
1%
1-
12
#209340000000
0!
0%
b11 *
0-
02
b11 6
#209350000000
1!
1%
1-
12
15
#209360000000
0!
0%
b100 *
0-
02
b100 6
#209370000000
1!
1%
1-
12
#209380000000
0!
0%
b101 *
0-
02
b101 6
#209390000000
1!
1%
1-
12
#209400000000
0!
0%
b110 *
0-
02
b110 6
#209410000000
1!
1%
1-
12
#209420000000
0!
0%
b111 *
0-
02
b111 6
#209430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#209440000000
0!
0%
b0 *
0-
02
b0 6
#209450000000
1!
1%
1-
12
#209460000000
0!
0%
b1 *
0-
02
b1 6
#209470000000
1!
1%
1-
12
#209480000000
0!
0%
b10 *
0-
02
b10 6
#209490000000
1!
1%
1-
12
#209500000000
0!
0%
b11 *
0-
02
b11 6
#209510000000
1!
1%
1-
12
15
#209520000000
0!
0%
b100 *
0-
02
b100 6
#209530000000
1!
1%
1-
12
#209540000000
0!
0%
b101 *
0-
02
b101 6
#209550000000
1!
1%
1-
12
#209560000000
0!
0%
b110 *
0-
02
b110 6
#209570000000
1!
1%
1-
12
#209580000000
0!
0%
b111 *
0-
02
b111 6
#209590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#209600000000
0!
0%
b0 *
0-
02
b0 6
#209610000000
1!
1%
1-
12
#209620000000
0!
0%
b1 *
0-
02
b1 6
#209630000000
1!
1%
1-
12
#209640000000
0!
0%
b10 *
0-
02
b10 6
#209650000000
1!
1%
1-
12
#209660000000
0!
0%
b11 *
0-
02
b11 6
#209670000000
1!
1%
1-
12
15
#209680000000
0!
0%
b100 *
0-
02
b100 6
#209690000000
1!
1%
1-
12
#209700000000
0!
0%
b101 *
0-
02
b101 6
#209710000000
1!
1%
1-
12
#209720000000
0!
0%
b110 *
0-
02
b110 6
#209730000000
1!
1%
1-
12
#209740000000
0!
0%
b111 *
0-
02
b111 6
#209750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#209760000000
0!
0%
b0 *
0-
02
b0 6
#209770000000
1!
1%
1-
12
#209780000000
0!
0%
b1 *
0-
02
b1 6
#209790000000
1!
1%
1-
12
#209800000000
0!
0%
b10 *
0-
02
b10 6
#209810000000
1!
1%
1-
12
#209820000000
0!
0%
b11 *
0-
02
b11 6
#209830000000
1!
1%
1-
12
15
#209840000000
0!
0%
b100 *
0-
02
b100 6
#209850000000
1!
1%
1-
12
#209860000000
0!
0%
b101 *
0-
02
b101 6
#209870000000
1!
1%
1-
12
#209880000000
0!
0%
b110 *
0-
02
b110 6
#209890000000
1!
1%
1-
12
#209900000000
0!
0%
b111 *
0-
02
b111 6
#209910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#209920000000
0!
0%
b0 *
0-
02
b0 6
#209930000000
1!
1%
1-
12
#209940000000
0!
0%
b1 *
0-
02
b1 6
#209950000000
1!
1%
1-
12
#209960000000
0!
0%
b10 *
0-
02
b10 6
#209970000000
1!
1%
1-
12
#209980000000
0!
0%
b11 *
0-
02
b11 6
#209990000000
1!
1%
1-
12
15
#210000000000
0!
0%
b100 *
0-
02
b100 6
#210010000000
1!
1%
1-
12
#210020000000
0!
0%
b101 *
0-
02
b101 6
#210030000000
1!
1%
1-
12
#210040000000
0!
0%
b110 *
0-
02
b110 6
#210050000000
1!
1%
1-
12
#210060000000
0!
0%
b111 *
0-
02
b111 6
#210070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#210080000000
0!
0%
b0 *
0-
02
b0 6
#210090000000
1!
1%
1-
12
#210100000000
0!
0%
b1 *
0-
02
b1 6
#210110000000
1!
1%
1-
12
#210120000000
0!
0%
b10 *
0-
02
b10 6
#210130000000
1!
1%
1-
12
#210140000000
0!
0%
b11 *
0-
02
b11 6
#210150000000
1!
1%
1-
12
15
#210160000000
0!
0%
b100 *
0-
02
b100 6
#210170000000
1!
1%
1-
12
#210180000000
0!
0%
b101 *
0-
02
b101 6
#210190000000
1!
1%
1-
12
#210200000000
0!
0%
b110 *
0-
02
b110 6
#210210000000
1!
1%
1-
12
#210220000000
0!
0%
b111 *
0-
02
b111 6
#210230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#210240000000
0!
0%
b0 *
0-
02
b0 6
#210250000000
1!
1%
1-
12
#210260000000
0!
0%
b1 *
0-
02
b1 6
#210270000000
1!
1%
1-
12
#210280000000
0!
0%
b10 *
0-
02
b10 6
#210290000000
1!
1%
1-
12
#210300000000
0!
0%
b11 *
0-
02
b11 6
#210310000000
1!
1%
1-
12
15
#210320000000
0!
0%
b100 *
0-
02
b100 6
#210330000000
1!
1%
1-
12
#210340000000
0!
0%
b101 *
0-
02
b101 6
#210350000000
1!
1%
1-
12
#210360000000
0!
0%
b110 *
0-
02
b110 6
#210370000000
1!
1%
1-
12
#210380000000
0!
0%
b111 *
0-
02
b111 6
#210390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#210400000000
0!
0%
b0 *
0-
02
b0 6
#210410000000
1!
1%
1-
12
#210420000000
0!
0%
b1 *
0-
02
b1 6
#210430000000
1!
1%
1-
12
#210440000000
0!
0%
b10 *
0-
02
b10 6
#210450000000
1!
1%
1-
12
#210460000000
0!
0%
b11 *
0-
02
b11 6
#210470000000
1!
1%
1-
12
15
#210480000000
0!
0%
b100 *
0-
02
b100 6
#210490000000
1!
1%
1-
12
#210500000000
0!
0%
b101 *
0-
02
b101 6
#210510000000
1!
1%
1-
12
#210520000000
0!
0%
b110 *
0-
02
b110 6
#210530000000
1!
1%
1-
12
#210540000000
0!
0%
b111 *
0-
02
b111 6
#210550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#210560000000
0!
0%
b0 *
0-
02
b0 6
#210570000000
1!
1%
1-
12
#210580000000
0!
0%
b1 *
0-
02
b1 6
#210590000000
1!
1%
1-
12
#210600000000
0!
0%
b10 *
0-
02
b10 6
#210610000000
1!
1%
1-
12
#210620000000
0!
0%
b11 *
0-
02
b11 6
#210630000000
1!
1%
1-
12
15
#210640000000
0!
0%
b100 *
0-
02
b100 6
#210650000000
1!
1%
1-
12
#210660000000
0!
0%
b101 *
0-
02
b101 6
#210670000000
1!
1%
1-
12
#210680000000
0!
0%
b110 *
0-
02
b110 6
#210690000000
1!
1%
1-
12
#210700000000
0!
0%
b111 *
0-
02
b111 6
#210710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#210720000000
0!
0%
b0 *
0-
02
b0 6
#210730000000
1!
1%
1-
12
#210740000000
0!
0%
b1 *
0-
02
b1 6
#210750000000
1!
1%
1-
12
#210760000000
0!
0%
b10 *
0-
02
b10 6
#210770000000
1!
1%
1-
12
#210780000000
0!
0%
b11 *
0-
02
b11 6
#210790000000
1!
1%
1-
12
15
#210800000000
0!
0%
b100 *
0-
02
b100 6
#210810000000
1!
1%
1-
12
#210820000000
0!
0%
b101 *
0-
02
b101 6
#210830000000
1!
1%
1-
12
#210840000000
0!
0%
b110 *
0-
02
b110 6
#210850000000
1!
1%
1-
12
#210860000000
0!
0%
b111 *
0-
02
b111 6
#210870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#210880000000
0!
0%
b0 *
0-
02
b0 6
#210890000000
1!
1%
1-
12
#210900000000
0!
0%
b1 *
0-
02
b1 6
#210910000000
1!
1%
1-
12
#210920000000
0!
0%
b10 *
0-
02
b10 6
#210930000000
1!
1%
1-
12
#210940000000
0!
0%
b11 *
0-
02
b11 6
#210950000000
1!
1%
1-
12
15
#210960000000
0!
0%
b100 *
0-
02
b100 6
#210970000000
1!
1%
1-
12
#210980000000
0!
0%
b101 *
0-
02
b101 6
#210990000000
1!
1%
1-
12
#211000000000
0!
0%
b110 *
0-
02
b110 6
#211010000000
1!
1%
1-
12
#211020000000
0!
0%
b111 *
0-
02
b111 6
#211030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#211040000000
0!
0%
b0 *
0-
02
b0 6
#211050000000
1!
1%
1-
12
#211060000000
0!
0%
b1 *
0-
02
b1 6
#211070000000
1!
1%
1-
12
#211080000000
0!
0%
b10 *
0-
02
b10 6
#211090000000
1!
1%
1-
12
#211100000000
0!
0%
b11 *
0-
02
b11 6
#211110000000
1!
1%
1-
12
15
#211120000000
0!
0%
b100 *
0-
02
b100 6
#211130000000
1!
1%
1-
12
#211140000000
0!
0%
b101 *
0-
02
b101 6
#211150000000
1!
1%
1-
12
#211160000000
0!
0%
b110 *
0-
02
b110 6
#211170000000
1!
1%
1-
12
#211180000000
0!
0%
b111 *
0-
02
b111 6
#211190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#211200000000
0!
0%
b0 *
0-
02
b0 6
#211210000000
1!
1%
1-
12
#211220000000
0!
0%
b1 *
0-
02
b1 6
#211230000000
1!
1%
1-
12
#211240000000
0!
0%
b10 *
0-
02
b10 6
#211250000000
1!
1%
1-
12
#211260000000
0!
0%
b11 *
0-
02
b11 6
#211270000000
1!
1%
1-
12
15
#211280000000
0!
0%
b100 *
0-
02
b100 6
#211290000000
1!
1%
1-
12
#211300000000
0!
0%
b101 *
0-
02
b101 6
#211310000000
1!
1%
1-
12
#211320000000
0!
0%
b110 *
0-
02
b110 6
#211330000000
1!
1%
1-
12
#211340000000
0!
0%
b111 *
0-
02
b111 6
#211350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#211360000000
0!
0%
b0 *
0-
02
b0 6
#211370000000
1!
1%
1-
12
#211380000000
0!
0%
b1 *
0-
02
b1 6
#211390000000
1!
1%
1-
12
#211400000000
0!
0%
b10 *
0-
02
b10 6
#211410000000
1!
1%
1-
12
#211420000000
0!
0%
b11 *
0-
02
b11 6
#211430000000
1!
1%
1-
12
15
#211440000000
0!
0%
b100 *
0-
02
b100 6
#211450000000
1!
1%
1-
12
#211460000000
0!
0%
b101 *
0-
02
b101 6
#211470000000
1!
1%
1-
12
#211480000000
0!
0%
b110 *
0-
02
b110 6
#211490000000
1!
1%
1-
12
#211500000000
0!
0%
b111 *
0-
02
b111 6
#211510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#211520000000
0!
0%
b0 *
0-
02
b0 6
#211530000000
1!
1%
1-
12
#211540000000
0!
0%
b1 *
0-
02
b1 6
#211550000000
1!
1%
1-
12
#211560000000
0!
0%
b10 *
0-
02
b10 6
#211570000000
1!
1%
1-
12
#211580000000
0!
0%
b11 *
0-
02
b11 6
#211590000000
1!
1%
1-
12
15
#211600000000
0!
0%
b100 *
0-
02
b100 6
#211610000000
1!
1%
1-
12
#211620000000
0!
0%
b101 *
0-
02
b101 6
#211630000000
1!
1%
1-
12
#211640000000
0!
0%
b110 *
0-
02
b110 6
#211650000000
1!
1%
1-
12
#211660000000
0!
0%
b111 *
0-
02
b111 6
#211670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#211680000000
0!
0%
b0 *
0-
02
b0 6
#211690000000
1!
1%
1-
12
#211700000000
0!
0%
b1 *
0-
02
b1 6
#211710000000
1!
1%
1-
12
#211720000000
0!
0%
b10 *
0-
02
b10 6
#211730000000
1!
1%
1-
12
#211740000000
0!
0%
b11 *
0-
02
b11 6
#211750000000
1!
1%
1-
12
15
#211760000000
0!
0%
b100 *
0-
02
b100 6
#211770000000
1!
1%
1-
12
#211780000000
0!
0%
b101 *
0-
02
b101 6
#211790000000
1!
1%
1-
12
#211800000000
0!
0%
b110 *
0-
02
b110 6
#211810000000
1!
1%
1-
12
#211820000000
0!
0%
b111 *
0-
02
b111 6
#211830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#211840000000
0!
0%
b0 *
0-
02
b0 6
#211850000000
1!
1%
1-
12
#211860000000
0!
0%
b1 *
0-
02
b1 6
#211870000000
1!
1%
1-
12
#211880000000
0!
0%
b10 *
0-
02
b10 6
#211890000000
1!
1%
1-
12
#211900000000
0!
0%
b11 *
0-
02
b11 6
#211910000000
1!
1%
1-
12
15
#211920000000
0!
0%
b100 *
0-
02
b100 6
#211930000000
1!
1%
1-
12
#211940000000
0!
0%
b101 *
0-
02
b101 6
#211950000000
1!
1%
1-
12
#211960000000
0!
0%
b110 *
0-
02
b110 6
#211970000000
1!
1%
1-
12
#211980000000
0!
0%
b111 *
0-
02
b111 6
#211990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#212000000000
0!
0%
b0 *
0-
02
b0 6
#212010000000
1!
1%
1-
12
#212020000000
0!
0%
b1 *
0-
02
b1 6
#212030000000
1!
1%
1-
12
#212040000000
0!
0%
b10 *
0-
02
b10 6
#212050000000
1!
1%
1-
12
#212060000000
0!
0%
b11 *
0-
02
b11 6
#212070000000
1!
1%
1-
12
15
#212080000000
0!
0%
b100 *
0-
02
b100 6
#212090000000
1!
1%
1-
12
#212100000000
0!
0%
b101 *
0-
02
b101 6
#212110000000
1!
1%
1-
12
#212120000000
0!
0%
b110 *
0-
02
b110 6
#212130000000
1!
1%
1-
12
#212140000000
0!
0%
b111 *
0-
02
b111 6
#212150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#212160000000
0!
0%
b0 *
0-
02
b0 6
#212170000000
1!
1%
1-
12
#212180000000
0!
0%
b1 *
0-
02
b1 6
#212190000000
1!
1%
1-
12
#212200000000
0!
0%
b10 *
0-
02
b10 6
#212210000000
1!
1%
1-
12
#212220000000
0!
0%
b11 *
0-
02
b11 6
#212230000000
1!
1%
1-
12
15
#212240000000
0!
0%
b100 *
0-
02
b100 6
#212250000000
1!
1%
1-
12
#212260000000
0!
0%
b101 *
0-
02
b101 6
#212270000000
1!
1%
1-
12
#212280000000
0!
0%
b110 *
0-
02
b110 6
#212290000000
1!
1%
1-
12
#212300000000
0!
0%
b111 *
0-
02
b111 6
#212310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#212320000000
0!
0%
b0 *
0-
02
b0 6
#212330000000
1!
1%
1-
12
#212340000000
0!
0%
b1 *
0-
02
b1 6
#212350000000
1!
1%
1-
12
#212360000000
0!
0%
b10 *
0-
02
b10 6
#212370000000
1!
1%
1-
12
#212380000000
0!
0%
b11 *
0-
02
b11 6
#212390000000
1!
1%
1-
12
15
#212400000000
0!
0%
b100 *
0-
02
b100 6
#212410000000
1!
1%
1-
12
#212420000000
0!
0%
b101 *
0-
02
b101 6
#212430000000
1!
1%
1-
12
#212440000000
0!
0%
b110 *
0-
02
b110 6
#212450000000
1!
1%
1-
12
#212460000000
0!
0%
b111 *
0-
02
b111 6
#212470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#212480000000
0!
0%
b0 *
0-
02
b0 6
#212490000000
1!
1%
1-
12
#212500000000
0!
0%
b1 *
0-
02
b1 6
#212510000000
1!
1%
1-
12
#212520000000
0!
0%
b10 *
0-
02
b10 6
#212530000000
1!
1%
1-
12
#212540000000
0!
0%
b11 *
0-
02
b11 6
#212550000000
1!
1%
1-
12
15
#212560000000
0!
0%
b100 *
0-
02
b100 6
#212570000000
1!
1%
1-
12
#212580000000
0!
0%
b101 *
0-
02
b101 6
#212590000000
1!
1%
1-
12
#212600000000
0!
0%
b110 *
0-
02
b110 6
#212610000000
1!
1%
1-
12
#212620000000
0!
0%
b111 *
0-
02
b111 6
#212630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#212640000000
0!
0%
b0 *
0-
02
b0 6
#212650000000
1!
1%
1-
12
#212660000000
0!
0%
b1 *
0-
02
b1 6
#212670000000
1!
1%
1-
12
#212680000000
0!
0%
b10 *
0-
02
b10 6
#212690000000
1!
1%
1-
12
#212700000000
0!
0%
b11 *
0-
02
b11 6
#212710000000
1!
1%
1-
12
15
#212720000000
0!
0%
b100 *
0-
02
b100 6
#212730000000
1!
1%
1-
12
#212740000000
0!
0%
b101 *
0-
02
b101 6
#212750000000
1!
1%
1-
12
#212760000000
0!
0%
b110 *
0-
02
b110 6
#212770000000
1!
1%
1-
12
#212780000000
0!
0%
b111 *
0-
02
b111 6
#212790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#212800000000
0!
0%
b0 *
0-
02
b0 6
#212810000000
1!
1%
1-
12
#212820000000
0!
0%
b1 *
0-
02
b1 6
#212830000000
1!
1%
1-
12
#212840000000
0!
0%
b10 *
0-
02
b10 6
#212850000000
1!
1%
1-
12
#212860000000
0!
0%
b11 *
0-
02
b11 6
#212870000000
1!
1%
1-
12
15
#212880000000
0!
0%
b100 *
0-
02
b100 6
#212890000000
1!
1%
1-
12
#212900000000
0!
0%
b101 *
0-
02
b101 6
#212910000000
1!
1%
1-
12
#212920000000
0!
0%
b110 *
0-
02
b110 6
#212930000000
1!
1%
1-
12
#212940000000
0!
0%
b111 *
0-
02
b111 6
#212950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#212960000000
0!
0%
b0 *
0-
02
b0 6
#212970000000
1!
1%
1-
12
#212980000000
0!
0%
b1 *
0-
02
b1 6
#212990000000
1!
1%
1-
12
#213000000000
0!
0%
b10 *
0-
02
b10 6
#213010000000
1!
1%
1-
12
#213020000000
0!
0%
b11 *
0-
02
b11 6
#213030000000
1!
1%
1-
12
15
#213040000000
0!
0%
b100 *
0-
02
b100 6
#213050000000
1!
1%
1-
12
#213060000000
0!
0%
b101 *
0-
02
b101 6
#213070000000
1!
1%
1-
12
#213080000000
0!
0%
b110 *
0-
02
b110 6
#213090000000
1!
1%
1-
12
#213100000000
0!
0%
b111 *
0-
02
b111 6
#213110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#213120000000
0!
0%
b0 *
0-
02
b0 6
#213130000000
1!
1%
1-
12
#213140000000
0!
0%
b1 *
0-
02
b1 6
#213150000000
1!
1%
1-
12
#213160000000
0!
0%
b10 *
0-
02
b10 6
#213170000000
1!
1%
1-
12
#213180000000
0!
0%
b11 *
0-
02
b11 6
#213190000000
1!
1%
1-
12
15
#213200000000
0!
0%
b100 *
0-
02
b100 6
#213210000000
1!
1%
1-
12
#213220000000
0!
0%
b101 *
0-
02
b101 6
#213230000000
1!
1%
1-
12
#213240000000
0!
0%
b110 *
0-
02
b110 6
#213250000000
1!
1%
1-
12
#213260000000
0!
0%
b111 *
0-
02
b111 6
#213270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#213280000000
0!
0%
b0 *
0-
02
b0 6
#213290000000
1!
1%
1-
12
#213300000000
0!
0%
b1 *
0-
02
b1 6
#213310000000
1!
1%
1-
12
#213320000000
0!
0%
b10 *
0-
02
b10 6
#213330000000
1!
1%
1-
12
#213340000000
0!
0%
b11 *
0-
02
b11 6
#213350000000
1!
1%
1-
12
15
#213360000000
0!
0%
b100 *
0-
02
b100 6
#213370000000
1!
1%
1-
12
#213380000000
0!
0%
b101 *
0-
02
b101 6
#213390000000
1!
1%
1-
12
#213400000000
0!
0%
b110 *
0-
02
b110 6
#213410000000
1!
1%
1-
12
#213420000000
0!
0%
b111 *
0-
02
b111 6
#213430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#213440000000
0!
0%
b0 *
0-
02
b0 6
#213450000000
1!
1%
1-
12
#213460000000
0!
0%
b1 *
0-
02
b1 6
#213470000000
1!
1%
1-
12
#213480000000
0!
0%
b10 *
0-
02
b10 6
#213490000000
1!
1%
1-
12
#213500000000
0!
0%
b11 *
0-
02
b11 6
#213510000000
1!
1%
1-
12
15
#213520000000
0!
0%
b100 *
0-
02
b100 6
#213530000000
1!
1%
1-
12
#213540000000
0!
0%
b101 *
0-
02
b101 6
#213550000000
1!
1%
1-
12
#213560000000
0!
0%
b110 *
0-
02
b110 6
#213570000000
1!
1%
1-
12
#213580000000
0!
0%
b111 *
0-
02
b111 6
#213590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#213600000000
0!
0%
b0 *
0-
02
b0 6
#213610000000
1!
1%
1-
12
#213620000000
0!
0%
b1 *
0-
02
b1 6
#213630000000
1!
1%
1-
12
#213640000000
0!
0%
b10 *
0-
02
b10 6
#213650000000
1!
1%
1-
12
#213660000000
0!
0%
b11 *
0-
02
b11 6
#213670000000
1!
1%
1-
12
15
#213680000000
0!
0%
b100 *
0-
02
b100 6
#213690000000
1!
1%
1-
12
#213700000000
0!
0%
b101 *
0-
02
b101 6
#213710000000
1!
1%
1-
12
#213720000000
0!
0%
b110 *
0-
02
b110 6
#213730000000
1!
1%
1-
12
#213740000000
0!
0%
b111 *
0-
02
b111 6
#213750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#213760000000
0!
0%
b0 *
0-
02
b0 6
#213770000000
1!
1%
1-
12
#213780000000
0!
0%
b1 *
0-
02
b1 6
#213790000000
1!
1%
1-
12
#213800000000
0!
0%
b10 *
0-
02
b10 6
#213810000000
1!
1%
1-
12
#213820000000
0!
0%
b11 *
0-
02
b11 6
#213830000000
1!
1%
1-
12
15
#213840000000
0!
0%
b100 *
0-
02
b100 6
#213850000000
1!
1%
1-
12
#213860000000
0!
0%
b101 *
0-
02
b101 6
#213870000000
1!
1%
1-
12
#213880000000
0!
0%
b110 *
0-
02
b110 6
#213890000000
1!
1%
1-
12
#213900000000
0!
0%
b111 *
0-
02
b111 6
#213910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#213920000000
0!
0%
b0 *
0-
02
b0 6
#213930000000
1!
1%
1-
12
#213940000000
0!
0%
b1 *
0-
02
b1 6
#213950000000
1!
1%
1-
12
#213960000000
0!
0%
b10 *
0-
02
b10 6
#213970000000
1!
1%
1-
12
#213980000000
0!
0%
b11 *
0-
02
b11 6
#213990000000
1!
1%
1-
12
15
#214000000000
0!
0%
b100 *
0-
02
b100 6
#214010000000
1!
1%
1-
12
#214020000000
0!
0%
b101 *
0-
02
b101 6
#214030000000
1!
1%
1-
12
#214040000000
0!
0%
b110 *
0-
02
b110 6
#214050000000
1!
1%
1-
12
#214060000000
0!
0%
b111 *
0-
02
b111 6
#214070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#214080000000
0!
0%
b0 *
0-
02
b0 6
#214090000000
1!
1%
1-
12
#214100000000
0!
0%
b1 *
0-
02
b1 6
#214110000000
1!
1%
1-
12
#214120000000
0!
0%
b10 *
0-
02
b10 6
#214130000000
1!
1%
1-
12
#214140000000
0!
0%
b11 *
0-
02
b11 6
#214150000000
1!
1%
1-
12
15
#214160000000
0!
0%
b100 *
0-
02
b100 6
#214170000000
1!
1%
1-
12
#214180000000
0!
0%
b101 *
0-
02
b101 6
#214190000000
1!
1%
1-
12
#214200000000
0!
0%
b110 *
0-
02
b110 6
#214210000000
1!
1%
1-
12
#214220000000
0!
0%
b111 *
0-
02
b111 6
#214230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#214240000000
0!
0%
b0 *
0-
02
b0 6
#214250000000
1!
1%
1-
12
#214260000000
0!
0%
b1 *
0-
02
b1 6
#214270000000
1!
1%
1-
12
#214280000000
0!
0%
b10 *
0-
02
b10 6
#214290000000
1!
1%
1-
12
#214300000000
0!
0%
b11 *
0-
02
b11 6
#214310000000
1!
1%
1-
12
15
#214320000000
0!
0%
b100 *
0-
02
b100 6
#214330000000
1!
1%
1-
12
#214340000000
0!
0%
b101 *
0-
02
b101 6
#214350000000
1!
1%
1-
12
#214360000000
0!
0%
b110 *
0-
02
b110 6
#214370000000
1!
1%
1-
12
#214380000000
0!
0%
b111 *
0-
02
b111 6
#214390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#214400000000
0!
0%
b0 *
0-
02
b0 6
#214410000000
1!
1%
1-
12
#214420000000
0!
0%
b1 *
0-
02
b1 6
#214430000000
1!
1%
1-
12
#214440000000
0!
0%
b10 *
0-
02
b10 6
#214450000000
1!
1%
1-
12
#214460000000
0!
0%
b11 *
0-
02
b11 6
#214470000000
1!
1%
1-
12
15
#214480000000
0!
0%
b100 *
0-
02
b100 6
#214490000000
1!
1%
1-
12
#214500000000
0!
0%
b101 *
0-
02
b101 6
#214510000000
1!
1%
1-
12
#214520000000
0!
0%
b110 *
0-
02
b110 6
#214530000000
1!
1%
1-
12
#214540000000
0!
0%
b111 *
0-
02
b111 6
#214550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#214560000000
0!
0%
b0 *
0-
02
b0 6
#214570000000
1!
1%
1-
12
#214580000000
0!
0%
b1 *
0-
02
b1 6
#214590000000
1!
1%
1-
12
#214600000000
0!
0%
b10 *
0-
02
b10 6
#214610000000
1!
1%
1-
12
#214620000000
0!
0%
b11 *
0-
02
b11 6
#214630000000
1!
1%
1-
12
15
#214640000000
0!
0%
b100 *
0-
02
b100 6
#214650000000
1!
1%
1-
12
#214660000000
0!
0%
b101 *
0-
02
b101 6
#214670000000
1!
1%
1-
12
#214680000000
0!
0%
b110 *
0-
02
b110 6
#214690000000
1!
1%
1-
12
#214700000000
0!
0%
b111 *
0-
02
b111 6
#214710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#214720000000
0!
0%
b0 *
0-
02
b0 6
#214730000000
1!
1%
1-
12
#214740000000
0!
0%
b1 *
0-
02
b1 6
#214750000000
1!
1%
1-
12
#214760000000
0!
0%
b10 *
0-
02
b10 6
#214770000000
1!
1%
1-
12
#214780000000
0!
0%
b11 *
0-
02
b11 6
#214790000000
1!
1%
1-
12
15
#214800000000
0!
0%
b100 *
0-
02
b100 6
#214810000000
1!
1%
1-
12
#214820000000
0!
0%
b101 *
0-
02
b101 6
#214830000000
1!
1%
1-
12
#214840000000
0!
0%
b110 *
0-
02
b110 6
#214850000000
1!
1%
1-
12
#214860000000
0!
0%
b111 *
0-
02
b111 6
#214870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#214880000000
0!
0%
b0 *
0-
02
b0 6
#214890000000
1!
1%
1-
12
#214900000000
0!
0%
b1 *
0-
02
b1 6
#214910000000
1!
1%
1-
12
#214920000000
0!
0%
b10 *
0-
02
b10 6
#214930000000
1!
1%
1-
12
#214940000000
0!
0%
b11 *
0-
02
b11 6
#214950000000
1!
1%
1-
12
15
#214960000000
0!
0%
b100 *
0-
02
b100 6
#214970000000
1!
1%
1-
12
#214980000000
0!
0%
b101 *
0-
02
b101 6
#214990000000
1!
1%
1-
12
#215000000000
0!
0%
b110 *
0-
02
b110 6
#215010000000
1!
1%
1-
12
#215020000000
0!
0%
b111 *
0-
02
b111 6
#215030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#215040000000
0!
0%
b0 *
0-
02
b0 6
#215050000000
1!
1%
1-
12
#215060000000
0!
0%
b1 *
0-
02
b1 6
#215070000000
1!
1%
1-
12
#215080000000
0!
0%
b10 *
0-
02
b10 6
#215090000000
1!
1%
1-
12
#215100000000
0!
0%
b11 *
0-
02
b11 6
#215110000000
1!
1%
1-
12
15
#215120000000
0!
0%
b100 *
0-
02
b100 6
#215130000000
1!
1%
1-
12
#215140000000
0!
0%
b101 *
0-
02
b101 6
#215150000000
1!
1%
1-
12
#215160000000
0!
0%
b110 *
0-
02
b110 6
#215170000000
1!
1%
1-
12
#215180000000
0!
0%
b111 *
0-
02
b111 6
#215190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#215200000000
0!
0%
b0 *
0-
02
b0 6
#215210000000
1!
1%
1-
12
#215220000000
0!
0%
b1 *
0-
02
b1 6
#215230000000
1!
1%
1-
12
#215240000000
0!
0%
b10 *
0-
02
b10 6
#215250000000
1!
1%
1-
12
#215260000000
0!
0%
b11 *
0-
02
b11 6
#215270000000
1!
1%
1-
12
15
#215280000000
0!
0%
b100 *
0-
02
b100 6
#215290000000
1!
1%
1-
12
#215300000000
0!
0%
b101 *
0-
02
b101 6
#215310000000
1!
1%
1-
12
#215320000000
0!
0%
b110 *
0-
02
b110 6
#215330000000
1!
1%
1-
12
#215340000000
0!
0%
b111 *
0-
02
b111 6
#215350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#215360000000
0!
0%
b0 *
0-
02
b0 6
#215370000000
1!
1%
1-
12
#215380000000
0!
0%
b1 *
0-
02
b1 6
#215390000000
1!
1%
1-
12
#215400000000
0!
0%
b10 *
0-
02
b10 6
#215410000000
1!
1%
1-
12
#215420000000
0!
0%
b11 *
0-
02
b11 6
#215430000000
1!
1%
1-
12
15
#215440000000
0!
0%
b100 *
0-
02
b100 6
#215450000000
1!
1%
1-
12
#215460000000
0!
0%
b101 *
0-
02
b101 6
#215470000000
1!
1%
1-
12
#215480000000
0!
0%
b110 *
0-
02
b110 6
#215490000000
1!
1%
1-
12
#215500000000
0!
0%
b111 *
0-
02
b111 6
#215510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#215520000000
0!
0%
b0 *
0-
02
b0 6
#215530000000
1!
1%
1-
12
#215540000000
0!
0%
b1 *
0-
02
b1 6
#215550000000
1!
1%
1-
12
#215560000000
0!
0%
b10 *
0-
02
b10 6
#215570000000
1!
1%
1-
12
#215580000000
0!
0%
b11 *
0-
02
b11 6
#215590000000
1!
1%
1-
12
15
#215600000000
0!
0%
b100 *
0-
02
b100 6
#215610000000
1!
1%
1-
12
#215620000000
0!
0%
b101 *
0-
02
b101 6
#215630000000
1!
1%
1-
12
#215640000000
0!
0%
b110 *
0-
02
b110 6
#215650000000
1!
1%
1-
12
#215660000000
0!
0%
b111 *
0-
02
b111 6
#215670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#215680000000
0!
0%
b0 *
0-
02
b0 6
#215690000000
1!
1%
1-
12
#215700000000
0!
0%
b1 *
0-
02
b1 6
#215710000000
1!
1%
1-
12
#215720000000
0!
0%
b10 *
0-
02
b10 6
#215730000000
1!
1%
1-
12
#215740000000
0!
0%
b11 *
0-
02
b11 6
#215750000000
1!
1%
1-
12
15
#215760000000
0!
0%
b100 *
0-
02
b100 6
#215770000000
1!
1%
1-
12
#215780000000
0!
0%
b101 *
0-
02
b101 6
#215790000000
1!
1%
1-
12
#215800000000
0!
0%
b110 *
0-
02
b110 6
#215810000000
1!
1%
1-
12
#215820000000
0!
0%
b111 *
0-
02
b111 6
#215830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#215840000000
0!
0%
b0 *
0-
02
b0 6
#215850000000
1!
1%
1-
12
#215860000000
0!
0%
b1 *
0-
02
b1 6
#215870000000
1!
1%
1-
12
#215880000000
0!
0%
b10 *
0-
02
b10 6
#215890000000
1!
1%
1-
12
#215900000000
0!
0%
b11 *
0-
02
b11 6
#215910000000
1!
1%
1-
12
15
#215920000000
0!
0%
b100 *
0-
02
b100 6
#215930000000
1!
1%
1-
12
#215940000000
0!
0%
b101 *
0-
02
b101 6
#215950000000
1!
1%
1-
12
#215960000000
0!
0%
b110 *
0-
02
b110 6
#215970000000
1!
1%
1-
12
#215980000000
0!
0%
b111 *
0-
02
b111 6
#215990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#216000000000
0!
0%
b0 *
0-
02
b0 6
#216010000000
1!
1%
1-
12
#216020000000
0!
0%
b1 *
0-
02
b1 6
#216030000000
1!
1%
1-
12
#216040000000
0!
0%
b10 *
0-
02
b10 6
#216050000000
1!
1%
1-
12
#216060000000
0!
0%
b11 *
0-
02
b11 6
#216070000000
1!
1%
1-
12
15
#216080000000
0!
0%
b100 *
0-
02
b100 6
#216090000000
1!
1%
1-
12
#216100000000
0!
0%
b101 *
0-
02
b101 6
#216110000000
1!
1%
1-
12
#216120000000
0!
0%
b110 *
0-
02
b110 6
#216130000000
1!
1%
1-
12
#216140000000
0!
0%
b111 *
0-
02
b111 6
#216150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#216160000000
0!
0%
b0 *
0-
02
b0 6
#216170000000
1!
1%
1-
12
#216180000000
0!
0%
b1 *
0-
02
b1 6
#216190000000
1!
1%
1-
12
#216200000000
0!
0%
b10 *
0-
02
b10 6
#216210000000
1!
1%
1-
12
#216220000000
0!
0%
b11 *
0-
02
b11 6
#216230000000
1!
1%
1-
12
15
#216240000000
0!
0%
b100 *
0-
02
b100 6
#216250000000
1!
1%
1-
12
#216260000000
0!
0%
b101 *
0-
02
b101 6
#216270000000
1!
1%
1-
12
#216280000000
0!
0%
b110 *
0-
02
b110 6
#216290000000
1!
1%
1-
12
#216300000000
0!
0%
b111 *
0-
02
b111 6
#216310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#216320000000
0!
0%
b0 *
0-
02
b0 6
#216330000000
1!
1%
1-
12
#216340000000
0!
0%
b1 *
0-
02
b1 6
#216350000000
1!
1%
1-
12
#216360000000
0!
0%
b10 *
0-
02
b10 6
#216370000000
1!
1%
1-
12
#216380000000
0!
0%
b11 *
0-
02
b11 6
#216390000000
1!
1%
1-
12
15
#216400000000
0!
0%
b100 *
0-
02
b100 6
#216410000000
1!
1%
1-
12
#216420000000
0!
0%
b101 *
0-
02
b101 6
#216430000000
1!
1%
1-
12
#216440000000
0!
0%
b110 *
0-
02
b110 6
#216450000000
1!
1%
1-
12
#216460000000
0!
0%
b111 *
0-
02
b111 6
#216470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#216480000000
0!
0%
b0 *
0-
02
b0 6
#216490000000
1!
1%
1-
12
#216500000000
0!
0%
b1 *
0-
02
b1 6
#216510000000
1!
1%
1-
12
#216520000000
0!
0%
b10 *
0-
02
b10 6
#216530000000
1!
1%
1-
12
#216540000000
0!
0%
b11 *
0-
02
b11 6
#216550000000
1!
1%
1-
12
15
#216560000000
0!
0%
b100 *
0-
02
b100 6
#216570000000
1!
1%
1-
12
#216580000000
0!
0%
b101 *
0-
02
b101 6
#216590000000
1!
1%
1-
12
#216600000000
0!
0%
b110 *
0-
02
b110 6
#216610000000
1!
1%
1-
12
#216620000000
0!
0%
b111 *
0-
02
b111 6
#216630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#216640000000
0!
0%
b0 *
0-
02
b0 6
#216650000000
1!
1%
1-
12
#216660000000
0!
0%
b1 *
0-
02
b1 6
#216670000000
1!
1%
1-
12
#216680000000
0!
0%
b10 *
0-
02
b10 6
#216690000000
1!
1%
1-
12
#216700000000
0!
0%
b11 *
0-
02
b11 6
#216710000000
1!
1%
1-
12
15
#216720000000
0!
0%
b100 *
0-
02
b100 6
#216730000000
1!
1%
1-
12
#216740000000
0!
0%
b101 *
0-
02
b101 6
#216750000000
1!
1%
1-
12
#216760000000
0!
0%
b110 *
0-
02
b110 6
#216770000000
1!
1%
1-
12
#216780000000
0!
0%
b111 *
0-
02
b111 6
#216790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#216800000000
0!
0%
b0 *
0-
02
b0 6
#216810000000
1!
1%
1-
12
#216820000000
0!
0%
b1 *
0-
02
b1 6
#216830000000
1!
1%
1-
12
#216840000000
0!
0%
b10 *
0-
02
b10 6
#216850000000
1!
1%
1-
12
#216860000000
0!
0%
b11 *
0-
02
b11 6
#216870000000
1!
1%
1-
12
15
#216880000000
0!
0%
b100 *
0-
02
b100 6
#216890000000
1!
1%
1-
12
#216900000000
0!
0%
b101 *
0-
02
b101 6
#216910000000
1!
1%
1-
12
#216920000000
0!
0%
b110 *
0-
02
b110 6
#216930000000
1!
1%
1-
12
#216940000000
0!
0%
b111 *
0-
02
b111 6
#216950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#216960000000
0!
0%
b0 *
0-
02
b0 6
#216970000000
1!
1%
1-
12
#216980000000
0!
0%
b1 *
0-
02
b1 6
#216990000000
1!
1%
1-
12
#217000000000
0!
0%
b10 *
0-
02
b10 6
#217010000000
1!
1%
1-
12
#217020000000
0!
0%
b11 *
0-
02
b11 6
#217030000000
1!
1%
1-
12
15
#217040000000
0!
0%
b100 *
0-
02
b100 6
#217050000000
1!
1%
1-
12
#217060000000
0!
0%
b101 *
0-
02
b101 6
#217070000000
1!
1%
1-
12
#217080000000
0!
0%
b110 *
0-
02
b110 6
#217090000000
1!
1%
1-
12
#217100000000
0!
0%
b111 *
0-
02
b111 6
#217110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#217120000000
0!
0%
b0 *
0-
02
b0 6
#217130000000
1!
1%
1-
12
#217140000000
0!
0%
b1 *
0-
02
b1 6
#217150000000
1!
1%
1-
12
#217160000000
0!
0%
b10 *
0-
02
b10 6
#217170000000
1!
1%
1-
12
#217180000000
0!
0%
b11 *
0-
02
b11 6
#217190000000
1!
1%
1-
12
15
#217200000000
0!
0%
b100 *
0-
02
b100 6
#217210000000
1!
1%
1-
12
#217220000000
0!
0%
b101 *
0-
02
b101 6
#217230000000
1!
1%
1-
12
#217240000000
0!
0%
b110 *
0-
02
b110 6
#217250000000
1!
1%
1-
12
#217260000000
0!
0%
b111 *
0-
02
b111 6
#217270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#217280000000
0!
0%
b0 *
0-
02
b0 6
#217290000000
1!
1%
1-
12
#217300000000
0!
0%
b1 *
0-
02
b1 6
#217310000000
1!
1%
1-
12
#217320000000
0!
0%
b10 *
0-
02
b10 6
#217330000000
1!
1%
1-
12
#217340000000
0!
0%
b11 *
0-
02
b11 6
#217350000000
1!
1%
1-
12
15
#217360000000
0!
0%
b100 *
0-
02
b100 6
#217370000000
1!
1%
1-
12
#217380000000
0!
0%
b101 *
0-
02
b101 6
#217390000000
1!
1%
1-
12
#217400000000
0!
0%
b110 *
0-
02
b110 6
#217410000000
1!
1%
1-
12
#217420000000
0!
0%
b111 *
0-
02
b111 6
#217430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#217440000000
0!
0%
b0 *
0-
02
b0 6
#217450000000
1!
1%
1-
12
#217460000000
0!
0%
b1 *
0-
02
b1 6
#217470000000
1!
1%
1-
12
#217480000000
0!
0%
b10 *
0-
02
b10 6
#217490000000
1!
1%
1-
12
#217500000000
0!
0%
b11 *
0-
02
b11 6
#217510000000
1!
1%
1-
12
15
#217520000000
0!
0%
b100 *
0-
02
b100 6
#217530000000
1!
1%
1-
12
#217540000000
0!
0%
b101 *
0-
02
b101 6
#217550000000
1!
1%
1-
12
#217560000000
0!
0%
b110 *
0-
02
b110 6
#217570000000
1!
1%
1-
12
#217580000000
0!
0%
b111 *
0-
02
b111 6
#217590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#217600000000
0!
0%
b0 *
0-
02
b0 6
#217610000000
1!
1%
1-
12
#217620000000
0!
0%
b1 *
0-
02
b1 6
#217630000000
1!
1%
1-
12
#217640000000
0!
0%
b10 *
0-
02
b10 6
#217650000000
1!
1%
1-
12
#217660000000
0!
0%
b11 *
0-
02
b11 6
#217670000000
1!
1%
1-
12
15
#217680000000
0!
0%
b100 *
0-
02
b100 6
#217690000000
1!
1%
1-
12
#217700000000
0!
0%
b101 *
0-
02
b101 6
#217710000000
1!
1%
1-
12
#217720000000
0!
0%
b110 *
0-
02
b110 6
#217730000000
1!
1%
1-
12
#217740000000
0!
0%
b111 *
0-
02
b111 6
#217750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#217760000000
0!
0%
b0 *
0-
02
b0 6
#217770000000
1!
1%
1-
12
#217780000000
0!
0%
b1 *
0-
02
b1 6
#217790000000
1!
1%
1-
12
#217800000000
0!
0%
b10 *
0-
02
b10 6
#217810000000
1!
1%
1-
12
#217820000000
0!
0%
b11 *
0-
02
b11 6
#217830000000
1!
1%
1-
12
15
#217840000000
0!
0%
b100 *
0-
02
b100 6
#217850000000
1!
1%
1-
12
#217860000000
0!
0%
b101 *
0-
02
b101 6
#217870000000
1!
1%
1-
12
#217880000000
0!
0%
b110 *
0-
02
b110 6
#217890000000
1!
1%
1-
12
#217900000000
0!
0%
b111 *
0-
02
b111 6
#217910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#217920000000
0!
0%
b0 *
0-
02
b0 6
#217930000000
1!
1%
1-
12
#217940000000
0!
0%
b1 *
0-
02
b1 6
#217950000000
1!
1%
1-
12
#217960000000
0!
0%
b10 *
0-
02
b10 6
#217970000000
1!
1%
1-
12
#217980000000
0!
0%
b11 *
0-
02
b11 6
#217990000000
1!
1%
1-
12
15
#218000000000
0!
0%
b100 *
0-
02
b100 6
#218010000000
1!
1%
1-
12
#218020000000
0!
0%
b101 *
0-
02
b101 6
#218030000000
1!
1%
1-
12
#218040000000
0!
0%
b110 *
0-
02
b110 6
#218050000000
1!
1%
1-
12
#218060000000
0!
0%
b111 *
0-
02
b111 6
#218070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#218080000000
0!
0%
b0 *
0-
02
b0 6
#218090000000
1!
1%
1-
12
#218100000000
0!
0%
b1 *
0-
02
b1 6
#218110000000
1!
1%
1-
12
#218120000000
0!
0%
b10 *
0-
02
b10 6
#218130000000
1!
1%
1-
12
#218140000000
0!
0%
b11 *
0-
02
b11 6
#218150000000
1!
1%
1-
12
15
#218160000000
0!
0%
b100 *
0-
02
b100 6
#218170000000
1!
1%
1-
12
#218180000000
0!
0%
b101 *
0-
02
b101 6
#218190000000
1!
1%
1-
12
#218200000000
0!
0%
b110 *
0-
02
b110 6
#218210000000
1!
1%
1-
12
#218220000000
0!
0%
b111 *
0-
02
b111 6
#218230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#218240000000
0!
0%
b0 *
0-
02
b0 6
#218250000000
1!
1%
1-
12
#218260000000
0!
0%
b1 *
0-
02
b1 6
#218270000000
1!
1%
1-
12
#218280000000
0!
0%
b10 *
0-
02
b10 6
#218290000000
1!
1%
1-
12
#218300000000
0!
0%
b11 *
0-
02
b11 6
#218310000000
1!
1%
1-
12
15
#218320000000
0!
0%
b100 *
0-
02
b100 6
#218330000000
1!
1%
1-
12
#218340000000
0!
0%
b101 *
0-
02
b101 6
#218350000000
1!
1%
1-
12
#218360000000
0!
0%
b110 *
0-
02
b110 6
#218370000000
1!
1%
1-
12
#218380000000
0!
0%
b111 *
0-
02
b111 6
#218390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#218400000000
0!
0%
b0 *
0-
02
b0 6
#218410000000
1!
1%
1-
12
#218420000000
0!
0%
b1 *
0-
02
b1 6
#218430000000
1!
1%
1-
12
#218440000000
0!
0%
b10 *
0-
02
b10 6
#218450000000
1!
1%
1-
12
#218460000000
0!
0%
b11 *
0-
02
b11 6
#218470000000
1!
1%
1-
12
15
#218480000000
0!
0%
b100 *
0-
02
b100 6
#218490000000
1!
1%
1-
12
#218500000000
0!
0%
b101 *
0-
02
b101 6
#218510000000
1!
1%
1-
12
#218520000000
0!
0%
b110 *
0-
02
b110 6
#218530000000
1!
1%
1-
12
#218540000000
0!
0%
b111 *
0-
02
b111 6
#218550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#218560000000
0!
0%
b0 *
0-
02
b0 6
#218570000000
1!
1%
1-
12
#218580000000
0!
0%
b1 *
0-
02
b1 6
#218590000000
1!
1%
1-
12
#218600000000
0!
0%
b10 *
0-
02
b10 6
#218610000000
1!
1%
1-
12
#218620000000
0!
0%
b11 *
0-
02
b11 6
#218630000000
1!
1%
1-
12
15
#218640000000
0!
0%
b100 *
0-
02
b100 6
#218650000000
1!
1%
1-
12
#218660000000
0!
0%
b101 *
0-
02
b101 6
#218670000000
1!
1%
1-
12
#218680000000
0!
0%
b110 *
0-
02
b110 6
#218690000000
1!
1%
1-
12
#218700000000
0!
0%
b111 *
0-
02
b111 6
#218710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#218720000000
0!
0%
b0 *
0-
02
b0 6
#218730000000
1!
1%
1-
12
#218740000000
0!
0%
b1 *
0-
02
b1 6
#218750000000
1!
1%
1-
12
#218760000000
0!
0%
b10 *
0-
02
b10 6
#218770000000
1!
1%
1-
12
#218780000000
0!
0%
b11 *
0-
02
b11 6
#218790000000
1!
1%
1-
12
15
#218800000000
0!
0%
b100 *
0-
02
b100 6
#218810000000
1!
1%
1-
12
#218820000000
0!
0%
b101 *
0-
02
b101 6
#218830000000
1!
1%
1-
12
#218840000000
0!
0%
b110 *
0-
02
b110 6
#218850000000
1!
1%
1-
12
#218860000000
0!
0%
b111 *
0-
02
b111 6
#218870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#218880000000
0!
0%
b0 *
0-
02
b0 6
#218890000000
1!
1%
1-
12
#218900000000
0!
0%
b1 *
0-
02
b1 6
#218910000000
1!
1%
1-
12
#218920000000
0!
0%
b10 *
0-
02
b10 6
#218930000000
1!
1%
1-
12
#218940000000
0!
0%
b11 *
0-
02
b11 6
#218950000000
1!
1%
1-
12
15
#218960000000
0!
0%
b100 *
0-
02
b100 6
#218970000000
1!
1%
1-
12
#218980000000
0!
0%
b101 *
0-
02
b101 6
#218990000000
1!
1%
1-
12
#219000000000
0!
0%
b110 *
0-
02
b110 6
#219010000000
1!
1%
1-
12
#219020000000
0!
0%
b111 *
0-
02
b111 6
#219030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#219040000000
0!
0%
b0 *
0-
02
b0 6
#219050000000
1!
1%
1-
12
#219060000000
0!
0%
b1 *
0-
02
b1 6
#219070000000
1!
1%
1-
12
#219080000000
0!
0%
b10 *
0-
02
b10 6
#219090000000
1!
1%
1-
12
#219100000000
0!
0%
b11 *
0-
02
b11 6
#219110000000
1!
1%
1-
12
15
#219120000000
0!
0%
b100 *
0-
02
b100 6
#219130000000
1!
1%
1-
12
#219140000000
0!
0%
b101 *
0-
02
b101 6
#219150000000
1!
1%
1-
12
#219160000000
0!
0%
b110 *
0-
02
b110 6
#219170000000
1!
1%
1-
12
#219180000000
0!
0%
b111 *
0-
02
b111 6
#219190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#219200000000
0!
0%
b0 *
0-
02
b0 6
#219210000000
1!
1%
1-
12
#219220000000
0!
0%
b1 *
0-
02
b1 6
#219230000000
1!
1%
1-
12
#219240000000
0!
0%
b10 *
0-
02
b10 6
#219250000000
1!
1%
1-
12
#219260000000
0!
0%
b11 *
0-
02
b11 6
#219270000000
1!
1%
1-
12
15
#219280000000
0!
0%
b100 *
0-
02
b100 6
#219290000000
1!
1%
1-
12
#219300000000
0!
0%
b101 *
0-
02
b101 6
#219310000000
1!
1%
1-
12
#219320000000
0!
0%
b110 *
0-
02
b110 6
#219330000000
1!
1%
1-
12
#219340000000
0!
0%
b111 *
0-
02
b111 6
#219350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#219360000000
0!
0%
b0 *
0-
02
b0 6
#219370000000
1!
1%
1-
12
#219380000000
0!
0%
b1 *
0-
02
b1 6
#219390000000
1!
1%
1-
12
#219400000000
0!
0%
b10 *
0-
02
b10 6
#219410000000
1!
1%
1-
12
#219420000000
0!
0%
b11 *
0-
02
b11 6
#219430000000
1!
1%
1-
12
15
#219440000000
0!
0%
b100 *
0-
02
b100 6
#219450000000
1!
1%
1-
12
#219460000000
0!
0%
b101 *
0-
02
b101 6
#219470000000
1!
1%
1-
12
#219480000000
0!
0%
b110 *
0-
02
b110 6
#219490000000
1!
1%
1-
12
#219500000000
0!
0%
b111 *
0-
02
b111 6
#219510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#219520000000
0!
0%
b0 *
0-
02
b0 6
#219530000000
1!
1%
1-
12
#219540000000
0!
0%
b1 *
0-
02
b1 6
#219550000000
1!
1%
1-
12
#219560000000
0!
0%
b10 *
0-
02
b10 6
#219570000000
1!
1%
1-
12
#219580000000
0!
0%
b11 *
0-
02
b11 6
#219590000000
1!
1%
1-
12
15
#219600000000
0!
0%
b100 *
0-
02
b100 6
#219610000000
1!
1%
1-
12
#219620000000
0!
0%
b101 *
0-
02
b101 6
#219630000000
1!
1%
1-
12
#219640000000
0!
0%
b110 *
0-
02
b110 6
#219650000000
1!
1%
1-
12
#219660000000
0!
0%
b111 *
0-
02
b111 6
#219670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#219680000000
0!
0%
b0 *
0-
02
b0 6
#219690000000
1!
1%
1-
12
#219700000000
0!
0%
b1 *
0-
02
b1 6
#219710000000
1!
1%
1-
12
#219720000000
0!
0%
b10 *
0-
02
b10 6
#219730000000
1!
1%
1-
12
#219740000000
0!
0%
b11 *
0-
02
b11 6
#219750000000
1!
1%
1-
12
15
#219760000000
0!
0%
b100 *
0-
02
b100 6
#219770000000
1!
1%
1-
12
#219780000000
0!
0%
b101 *
0-
02
b101 6
#219790000000
1!
1%
1-
12
#219800000000
0!
0%
b110 *
0-
02
b110 6
#219810000000
1!
1%
1-
12
#219820000000
0!
0%
b111 *
0-
02
b111 6
#219830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#219840000000
0!
0%
b0 *
0-
02
b0 6
#219850000000
1!
1%
1-
12
#219860000000
0!
0%
b1 *
0-
02
b1 6
#219870000000
1!
1%
1-
12
#219880000000
0!
0%
b10 *
0-
02
b10 6
#219890000000
1!
1%
1-
12
#219900000000
0!
0%
b11 *
0-
02
b11 6
#219910000000
1!
1%
1-
12
15
#219920000000
0!
0%
b100 *
0-
02
b100 6
#219930000000
1!
1%
1-
12
#219940000000
0!
0%
b101 *
0-
02
b101 6
#219950000000
1!
1%
1-
12
#219960000000
0!
0%
b110 *
0-
02
b110 6
#219970000000
1!
1%
1-
12
#219980000000
0!
0%
b111 *
0-
02
b111 6
#219990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#220000000000
0!
0%
b0 *
0-
02
b0 6
#220010000000
1!
1%
1-
12
#220020000000
0!
0%
b1 *
0-
02
b1 6
#220030000000
1!
1%
1-
12
#220040000000
0!
0%
b10 *
0-
02
b10 6
#220050000000
1!
1%
1-
12
#220060000000
0!
0%
b11 *
0-
02
b11 6
#220070000000
1!
1%
1-
12
15
#220080000000
0!
0%
b100 *
0-
02
b100 6
#220090000000
1!
1%
1-
12
#220100000000
0!
0%
b101 *
0-
02
b101 6
#220110000000
1!
1%
1-
12
#220120000000
0!
0%
b110 *
0-
02
b110 6
#220130000000
1!
1%
1-
12
#220140000000
0!
0%
b111 *
0-
02
b111 6
#220150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#220160000000
0!
0%
b0 *
0-
02
b0 6
#220170000000
1!
1%
1-
12
#220180000000
0!
0%
b1 *
0-
02
b1 6
#220190000000
1!
1%
1-
12
#220200000000
0!
0%
b10 *
0-
02
b10 6
#220210000000
1!
1%
1-
12
#220220000000
0!
0%
b11 *
0-
02
b11 6
#220230000000
1!
1%
1-
12
15
#220240000000
0!
0%
b100 *
0-
02
b100 6
#220250000000
1!
1%
1-
12
#220260000000
0!
0%
b101 *
0-
02
b101 6
#220270000000
1!
1%
1-
12
#220280000000
0!
0%
b110 *
0-
02
b110 6
#220290000000
1!
1%
1-
12
#220300000000
0!
0%
b111 *
0-
02
b111 6
#220310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#220320000000
0!
0%
b0 *
0-
02
b0 6
#220330000000
1!
1%
1-
12
#220340000000
0!
0%
b1 *
0-
02
b1 6
#220350000000
1!
1%
1-
12
#220360000000
0!
0%
b10 *
0-
02
b10 6
#220370000000
1!
1%
1-
12
#220380000000
0!
0%
b11 *
0-
02
b11 6
#220390000000
1!
1%
1-
12
15
#220400000000
0!
0%
b100 *
0-
02
b100 6
#220410000000
1!
1%
1-
12
#220420000000
0!
0%
b101 *
0-
02
b101 6
#220430000000
1!
1%
1-
12
#220440000000
0!
0%
b110 *
0-
02
b110 6
#220450000000
1!
1%
1-
12
#220460000000
0!
0%
b111 *
0-
02
b111 6
#220470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#220480000000
0!
0%
b0 *
0-
02
b0 6
#220490000000
1!
1%
1-
12
#220500000000
0!
0%
b1 *
0-
02
b1 6
#220510000000
1!
1%
1-
12
#220520000000
0!
0%
b10 *
0-
02
b10 6
#220530000000
1!
1%
1-
12
#220540000000
0!
0%
b11 *
0-
02
b11 6
#220550000000
1!
1%
1-
12
15
#220560000000
0!
0%
b100 *
0-
02
b100 6
#220570000000
1!
1%
1-
12
#220580000000
0!
0%
b101 *
0-
02
b101 6
#220590000000
1!
1%
1-
12
#220600000000
0!
0%
b110 *
0-
02
b110 6
#220610000000
1!
1%
1-
12
#220620000000
0!
0%
b111 *
0-
02
b111 6
#220630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#220640000000
0!
0%
b0 *
0-
02
b0 6
#220650000000
1!
1%
1-
12
#220660000000
0!
0%
b1 *
0-
02
b1 6
#220670000000
1!
1%
1-
12
#220680000000
0!
0%
b10 *
0-
02
b10 6
#220690000000
1!
1%
1-
12
#220700000000
0!
0%
b11 *
0-
02
b11 6
#220710000000
1!
1%
1-
12
15
#220720000000
0!
0%
b100 *
0-
02
b100 6
#220730000000
1!
1%
1-
12
#220740000000
0!
0%
b101 *
0-
02
b101 6
#220750000000
1!
1%
1-
12
#220760000000
0!
0%
b110 *
0-
02
b110 6
#220770000000
1!
1%
1-
12
#220780000000
0!
0%
b111 *
0-
02
b111 6
#220790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#220800000000
0!
0%
b0 *
0-
02
b0 6
#220810000000
1!
1%
1-
12
#220820000000
0!
0%
b1 *
0-
02
b1 6
#220830000000
1!
1%
1-
12
#220840000000
0!
0%
b10 *
0-
02
b10 6
#220850000000
1!
1%
1-
12
#220860000000
0!
0%
b11 *
0-
02
b11 6
#220870000000
1!
1%
1-
12
15
#220880000000
0!
0%
b100 *
0-
02
b100 6
#220890000000
1!
1%
1-
12
#220900000000
0!
0%
b101 *
0-
02
b101 6
#220910000000
1!
1%
1-
12
#220920000000
0!
0%
b110 *
0-
02
b110 6
#220930000000
1!
1%
1-
12
#220940000000
0!
0%
b111 *
0-
02
b111 6
#220950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#220960000000
0!
0%
b0 *
0-
02
b0 6
#220970000000
1!
1%
1-
12
#220980000000
0!
0%
b1 *
0-
02
b1 6
#220990000000
1!
1%
1-
12
#221000000000
0!
0%
b10 *
0-
02
b10 6
#221010000000
1!
1%
1-
12
#221020000000
0!
0%
b11 *
0-
02
b11 6
#221030000000
1!
1%
1-
12
15
#221040000000
0!
0%
b100 *
0-
02
b100 6
#221050000000
1!
1%
1-
12
#221060000000
0!
0%
b101 *
0-
02
b101 6
#221070000000
1!
1%
1-
12
#221080000000
0!
0%
b110 *
0-
02
b110 6
#221090000000
1!
1%
1-
12
#221100000000
0!
0%
b111 *
0-
02
b111 6
#221110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#221120000000
0!
0%
b0 *
0-
02
b0 6
#221130000000
1!
1%
1-
12
#221140000000
0!
0%
b1 *
0-
02
b1 6
#221150000000
1!
1%
1-
12
#221160000000
0!
0%
b10 *
0-
02
b10 6
#221170000000
1!
1%
1-
12
#221180000000
0!
0%
b11 *
0-
02
b11 6
#221190000000
1!
1%
1-
12
15
#221200000000
0!
0%
b100 *
0-
02
b100 6
#221210000000
1!
1%
1-
12
#221220000000
0!
0%
b101 *
0-
02
b101 6
#221230000000
1!
1%
1-
12
#221240000000
0!
0%
b110 *
0-
02
b110 6
#221250000000
1!
1%
1-
12
#221260000000
0!
0%
b111 *
0-
02
b111 6
#221270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#221280000000
0!
0%
b0 *
0-
02
b0 6
#221290000000
1!
1%
1-
12
#221300000000
0!
0%
b1 *
0-
02
b1 6
#221310000000
1!
1%
1-
12
#221320000000
0!
0%
b10 *
0-
02
b10 6
#221330000000
1!
1%
1-
12
#221340000000
0!
0%
b11 *
0-
02
b11 6
#221350000000
1!
1%
1-
12
15
#221360000000
0!
0%
b100 *
0-
02
b100 6
#221370000000
1!
1%
1-
12
#221380000000
0!
0%
b101 *
0-
02
b101 6
#221390000000
1!
1%
1-
12
#221400000000
0!
0%
b110 *
0-
02
b110 6
#221410000000
1!
1%
1-
12
#221420000000
0!
0%
b111 *
0-
02
b111 6
#221430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#221440000000
0!
0%
b0 *
0-
02
b0 6
#221450000000
1!
1%
1-
12
#221460000000
0!
0%
b1 *
0-
02
b1 6
#221470000000
1!
1%
1-
12
#221480000000
0!
0%
b10 *
0-
02
b10 6
#221490000000
1!
1%
1-
12
#221500000000
0!
0%
b11 *
0-
02
b11 6
#221510000000
1!
1%
1-
12
15
#221520000000
0!
0%
b100 *
0-
02
b100 6
#221530000000
1!
1%
1-
12
#221540000000
0!
0%
b101 *
0-
02
b101 6
#221550000000
1!
1%
1-
12
#221560000000
0!
0%
b110 *
0-
02
b110 6
#221570000000
1!
1%
1-
12
#221580000000
0!
0%
b111 *
0-
02
b111 6
#221590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#221600000000
0!
0%
b0 *
0-
02
b0 6
#221610000000
1!
1%
1-
12
#221620000000
0!
0%
b1 *
0-
02
b1 6
#221630000000
1!
1%
1-
12
#221640000000
0!
0%
b10 *
0-
02
b10 6
#221650000000
1!
1%
1-
12
#221660000000
0!
0%
b11 *
0-
02
b11 6
#221670000000
1!
1%
1-
12
15
#221680000000
0!
0%
b100 *
0-
02
b100 6
#221690000000
1!
1%
1-
12
#221700000000
0!
0%
b101 *
0-
02
b101 6
#221710000000
1!
1%
1-
12
#221720000000
0!
0%
b110 *
0-
02
b110 6
#221730000000
1!
1%
1-
12
#221740000000
0!
0%
b111 *
0-
02
b111 6
#221750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#221760000000
0!
0%
b0 *
0-
02
b0 6
#221770000000
1!
1%
1-
12
#221780000000
0!
0%
b1 *
0-
02
b1 6
#221790000000
1!
1%
1-
12
#221800000000
0!
0%
b10 *
0-
02
b10 6
#221810000000
1!
1%
1-
12
#221820000000
0!
0%
b11 *
0-
02
b11 6
#221830000000
1!
1%
1-
12
15
#221840000000
0!
0%
b100 *
0-
02
b100 6
#221850000000
1!
1%
1-
12
#221860000000
0!
0%
b101 *
0-
02
b101 6
#221870000000
1!
1%
1-
12
#221880000000
0!
0%
b110 *
0-
02
b110 6
#221890000000
1!
1%
1-
12
#221900000000
0!
0%
b111 *
0-
02
b111 6
#221910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#221920000000
0!
0%
b0 *
0-
02
b0 6
#221930000000
1!
1%
1-
12
#221940000000
0!
0%
b1 *
0-
02
b1 6
#221950000000
1!
1%
1-
12
#221960000000
0!
0%
b10 *
0-
02
b10 6
#221970000000
1!
1%
1-
12
#221980000000
0!
0%
b11 *
0-
02
b11 6
#221990000000
1!
1%
1-
12
15
#222000000000
0!
0%
b100 *
0-
02
b100 6
#222010000000
1!
1%
1-
12
#222020000000
0!
0%
b101 *
0-
02
b101 6
#222030000000
1!
1%
1-
12
#222040000000
0!
0%
b110 *
0-
02
b110 6
#222050000000
1!
1%
1-
12
#222060000000
0!
0%
b111 *
0-
02
b111 6
#222070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#222080000000
0!
0%
b0 *
0-
02
b0 6
#222090000000
1!
1%
1-
12
#222100000000
0!
0%
b1 *
0-
02
b1 6
#222110000000
1!
1%
1-
12
#222120000000
0!
0%
b10 *
0-
02
b10 6
#222130000000
1!
1%
1-
12
#222140000000
0!
0%
b11 *
0-
02
b11 6
#222150000000
1!
1%
1-
12
15
#222160000000
0!
0%
b100 *
0-
02
b100 6
#222170000000
1!
1%
1-
12
#222180000000
0!
0%
b101 *
0-
02
b101 6
#222190000000
1!
1%
1-
12
#222200000000
0!
0%
b110 *
0-
02
b110 6
#222210000000
1!
1%
1-
12
#222220000000
0!
0%
b111 *
0-
02
b111 6
#222230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#222240000000
0!
0%
b0 *
0-
02
b0 6
#222250000000
1!
1%
1-
12
#222260000000
0!
0%
b1 *
0-
02
b1 6
#222270000000
1!
1%
1-
12
#222280000000
0!
0%
b10 *
0-
02
b10 6
#222290000000
1!
1%
1-
12
#222300000000
0!
0%
b11 *
0-
02
b11 6
#222310000000
1!
1%
1-
12
15
#222320000000
0!
0%
b100 *
0-
02
b100 6
#222330000000
1!
1%
1-
12
#222340000000
0!
0%
b101 *
0-
02
b101 6
#222350000000
1!
1%
1-
12
#222360000000
0!
0%
b110 *
0-
02
b110 6
#222370000000
1!
1%
1-
12
#222380000000
0!
0%
b111 *
0-
02
b111 6
#222390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#222400000000
0!
0%
b0 *
0-
02
b0 6
#222410000000
1!
1%
1-
12
#222420000000
0!
0%
b1 *
0-
02
b1 6
#222430000000
1!
1%
1-
12
#222440000000
0!
0%
b10 *
0-
02
b10 6
#222450000000
1!
1%
1-
12
#222460000000
0!
0%
b11 *
0-
02
b11 6
#222470000000
1!
1%
1-
12
15
#222480000000
0!
0%
b100 *
0-
02
b100 6
#222490000000
1!
1%
1-
12
#222500000000
0!
0%
b101 *
0-
02
b101 6
#222510000000
1!
1%
1-
12
#222520000000
0!
0%
b110 *
0-
02
b110 6
#222530000000
1!
1%
1-
12
#222540000000
0!
0%
b111 *
0-
02
b111 6
#222550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#222560000000
0!
0%
b0 *
0-
02
b0 6
#222570000000
1!
1%
1-
12
#222580000000
0!
0%
b1 *
0-
02
b1 6
#222590000000
1!
1%
1-
12
#222600000000
0!
0%
b10 *
0-
02
b10 6
#222610000000
1!
1%
1-
12
#222620000000
0!
0%
b11 *
0-
02
b11 6
#222630000000
1!
1%
1-
12
15
#222640000000
0!
0%
b100 *
0-
02
b100 6
#222650000000
1!
1%
1-
12
#222660000000
0!
0%
b101 *
0-
02
b101 6
#222670000000
1!
1%
1-
12
#222680000000
0!
0%
b110 *
0-
02
b110 6
#222690000000
1!
1%
1-
12
#222700000000
0!
0%
b111 *
0-
02
b111 6
#222710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#222720000000
0!
0%
b0 *
0-
02
b0 6
#222730000000
1!
1%
1-
12
#222740000000
0!
0%
b1 *
0-
02
b1 6
#222750000000
1!
1%
1-
12
#222760000000
0!
0%
b10 *
0-
02
b10 6
#222770000000
1!
1%
1-
12
#222780000000
0!
0%
b11 *
0-
02
b11 6
#222790000000
1!
1%
1-
12
15
#222800000000
0!
0%
b100 *
0-
02
b100 6
#222810000000
1!
1%
1-
12
#222820000000
0!
0%
b101 *
0-
02
b101 6
#222830000000
1!
1%
1-
12
#222840000000
0!
0%
b110 *
0-
02
b110 6
#222850000000
1!
1%
1-
12
#222860000000
0!
0%
b111 *
0-
02
b111 6
#222870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#222880000000
0!
0%
b0 *
0-
02
b0 6
#222890000000
1!
1%
1-
12
#222900000000
0!
0%
b1 *
0-
02
b1 6
#222910000000
1!
1%
1-
12
#222920000000
0!
0%
b10 *
0-
02
b10 6
#222930000000
1!
1%
1-
12
#222940000000
0!
0%
b11 *
0-
02
b11 6
#222950000000
1!
1%
1-
12
15
#222960000000
0!
0%
b100 *
0-
02
b100 6
#222970000000
1!
1%
1-
12
#222980000000
0!
0%
b101 *
0-
02
b101 6
#222990000000
1!
1%
1-
12
#223000000000
0!
0%
b110 *
0-
02
b110 6
#223010000000
1!
1%
1-
12
#223020000000
0!
0%
b111 *
0-
02
b111 6
#223030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#223040000000
0!
0%
b0 *
0-
02
b0 6
#223050000000
1!
1%
1-
12
#223060000000
0!
0%
b1 *
0-
02
b1 6
#223070000000
1!
1%
1-
12
#223080000000
0!
0%
b10 *
0-
02
b10 6
#223090000000
1!
1%
1-
12
#223100000000
0!
0%
b11 *
0-
02
b11 6
#223110000000
1!
1%
1-
12
15
#223120000000
0!
0%
b100 *
0-
02
b100 6
#223130000000
1!
1%
1-
12
#223140000000
0!
0%
b101 *
0-
02
b101 6
#223150000000
1!
1%
1-
12
#223160000000
0!
0%
b110 *
0-
02
b110 6
#223170000000
1!
1%
1-
12
#223180000000
0!
0%
b111 *
0-
02
b111 6
#223190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#223200000000
0!
0%
b0 *
0-
02
b0 6
#223210000000
1!
1%
1-
12
#223220000000
0!
0%
b1 *
0-
02
b1 6
#223230000000
1!
1%
1-
12
#223240000000
0!
0%
b10 *
0-
02
b10 6
#223250000000
1!
1%
1-
12
#223260000000
0!
0%
b11 *
0-
02
b11 6
#223270000000
1!
1%
1-
12
15
#223280000000
0!
0%
b100 *
0-
02
b100 6
#223290000000
1!
1%
1-
12
#223300000000
0!
0%
b101 *
0-
02
b101 6
#223310000000
1!
1%
1-
12
#223320000000
0!
0%
b110 *
0-
02
b110 6
#223330000000
1!
1%
1-
12
#223340000000
0!
0%
b111 *
0-
02
b111 6
#223350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#223360000000
0!
0%
b0 *
0-
02
b0 6
#223370000000
1!
1%
1-
12
#223380000000
0!
0%
b1 *
0-
02
b1 6
#223390000000
1!
1%
1-
12
#223400000000
0!
0%
b10 *
0-
02
b10 6
#223410000000
1!
1%
1-
12
#223420000000
0!
0%
b11 *
0-
02
b11 6
#223430000000
1!
1%
1-
12
15
#223440000000
0!
0%
b100 *
0-
02
b100 6
#223450000000
1!
1%
1-
12
#223460000000
0!
0%
b101 *
0-
02
b101 6
#223470000000
1!
1%
1-
12
#223480000000
0!
0%
b110 *
0-
02
b110 6
#223490000000
1!
1%
1-
12
#223500000000
0!
0%
b111 *
0-
02
b111 6
#223510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#223520000000
0!
0%
b0 *
0-
02
b0 6
#223530000000
1!
1%
1-
12
#223540000000
0!
0%
b1 *
0-
02
b1 6
#223550000000
1!
1%
1-
12
#223560000000
0!
0%
b10 *
0-
02
b10 6
#223570000000
1!
1%
1-
12
#223580000000
0!
0%
b11 *
0-
02
b11 6
#223590000000
1!
1%
1-
12
15
#223600000000
0!
0%
b100 *
0-
02
b100 6
#223610000000
1!
1%
1-
12
#223620000000
0!
0%
b101 *
0-
02
b101 6
#223630000000
1!
1%
1-
12
#223640000000
0!
0%
b110 *
0-
02
b110 6
#223650000000
1!
1%
1-
12
#223660000000
0!
0%
b111 *
0-
02
b111 6
#223670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#223680000000
0!
0%
b0 *
0-
02
b0 6
#223690000000
1!
1%
1-
12
#223700000000
0!
0%
b1 *
0-
02
b1 6
#223710000000
1!
1%
1-
12
#223720000000
0!
0%
b10 *
0-
02
b10 6
#223730000000
1!
1%
1-
12
#223740000000
0!
0%
b11 *
0-
02
b11 6
#223750000000
1!
1%
1-
12
15
#223760000000
0!
0%
b100 *
0-
02
b100 6
#223770000000
1!
1%
1-
12
#223780000000
0!
0%
b101 *
0-
02
b101 6
#223790000000
1!
1%
1-
12
#223800000000
0!
0%
b110 *
0-
02
b110 6
#223810000000
1!
1%
1-
12
#223820000000
0!
0%
b111 *
0-
02
b111 6
#223830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#223840000000
0!
0%
b0 *
0-
02
b0 6
#223850000000
1!
1%
1-
12
#223860000000
0!
0%
b1 *
0-
02
b1 6
#223870000000
1!
1%
1-
12
#223880000000
0!
0%
b10 *
0-
02
b10 6
#223890000000
1!
1%
1-
12
#223900000000
0!
0%
b11 *
0-
02
b11 6
#223910000000
1!
1%
1-
12
15
#223920000000
0!
0%
b100 *
0-
02
b100 6
#223930000000
1!
1%
1-
12
#223940000000
0!
0%
b101 *
0-
02
b101 6
#223950000000
1!
1%
1-
12
#223960000000
0!
0%
b110 *
0-
02
b110 6
#223970000000
1!
1%
1-
12
#223980000000
0!
0%
b111 *
0-
02
b111 6
#223990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#224000000000
0!
0%
b0 *
0-
02
b0 6
#224010000000
1!
1%
1-
12
#224020000000
0!
0%
b1 *
0-
02
b1 6
#224030000000
1!
1%
1-
12
#224040000000
0!
0%
b10 *
0-
02
b10 6
#224050000000
1!
1%
1-
12
#224060000000
0!
0%
b11 *
0-
02
b11 6
#224070000000
1!
1%
1-
12
15
#224080000000
0!
0%
b100 *
0-
02
b100 6
#224090000000
1!
1%
1-
12
#224100000000
0!
0%
b101 *
0-
02
b101 6
#224110000000
1!
1%
1-
12
#224120000000
0!
0%
b110 *
0-
02
b110 6
#224130000000
1!
1%
1-
12
#224140000000
0!
0%
b111 *
0-
02
b111 6
#224150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#224160000000
0!
0%
b0 *
0-
02
b0 6
#224170000000
1!
1%
1-
12
#224180000000
0!
0%
b1 *
0-
02
b1 6
#224190000000
1!
1%
1-
12
#224200000000
0!
0%
b10 *
0-
02
b10 6
#224210000000
1!
1%
1-
12
#224220000000
0!
0%
b11 *
0-
02
b11 6
#224230000000
1!
1%
1-
12
15
#224240000000
0!
0%
b100 *
0-
02
b100 6
#224250000000
1!
1%
1-
12
#224260000000
0!
0%
b101 *
0-
02
b101 6
#224270000000
1!
1%
1-
12
#224280000000
0!
0%
b110 *
0-
02
b110 6
#224290000000
1!
1%
1-
12
#224300000000
0!
0%
b111 *
0-
02
b111 6
#224310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#224320000000
0!
0%
b0 *
0-
02
b0 6
#224330000000
1!
1%
1-
12
#224340000000
0!
0%
b1 *
0-
02
b1 6
#224350000000
1!
1%
1-
12
#224360000000
0!
0%
b10 *
0-
02
b10 6
#224370000000
1!
1%
1-
12
#224380000000
0!
0%
b11 *
0-
02
b11 6
#224390000000
1!
1%
1-
12
15
#224400000000
0!
0%
b100 *
0-
02
b100 6
#224410000000
1!
1%
1-
12
#224420000000
0!
0%
b101 *
0-
02
b101 6
#224430000000
1!
1%
1-
12
#224440000000
0!
0%
b110 *
0-
02
b110 6
#224450000000
1!
1%
1-
12
#224460000000
0!
0%
b111 *
0-
02
b111 6
#224470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#224480000000
0!
0%
b0 *
0-
02
b0 6
#224490000000
1!
1%
1-
12
#224500000000
0!
0%
b1 *
0-
02
b1 6
#224510000000
1!
1%
1-
12
#224520000000
0!
0%
b10 *
0-
02
b10 6
#224530000000
1!
1%
1-
12
#224540000000
0!
0%
b11 *
0-
02
b11 6
#224550000000
1!
1%
1-
12
15
#224560000000
0!
0%
b100 *
0-
02
b100 6
#224570000000
1!
1%
1-
12
#224580000000
0!
0%
b101 *
0-
02
b101 6
#224590000000
1!
1%
1-
12
#224600000000
0!
0%
b110 *
0-
02
b110 6
#224610000000
1!
1%
1-
12
#224620000000
0!
0%
b111 *
0-
02
b111 6
#224630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#224640000000
0!
0%
b0 *
0-
02
b0 6
#224650000000
1!
1%
1-
12
#224660000000
0!
0%
b1 *
0-
02
b1 6
#224670000000
1!
1%
1-
12
#224680000000
0!
0%
b10 *
0-
02
b10 6
#224690000000
1!
1%
1-
12
#224700000000
0!
0%
b11 *
0-
02
b11 6
#224710000000
1!
1%
1-
12
15
#224720000000
0!
0%
b100 *
0-
02
b100 6
#224730000000
1!
1%
1-
12
#224740000000
0!
0%
b101 *
0-
02
b101 6
#224750000000
1!
1%
1-
12
#224760000000
0!
0%
b110 *
0-
02
b110 6
#224770000000
1!
1%
1-
12
#224780000000
0!
0%
b111 *
0-
02
b111 6
#224790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#224800000000
0!
0%
b0 *
0-
02
b0 6
#224810000000
1!
1%
1-
12
#224820000000
0!
0%
b1 *
0-
02
b1 6
#224830000000
1!
1%
1-
12
#224840000000
0!
0%
b10 *
0-
02
b10 6
#224850000000
1!
1%
1-
12
#224860000000
0!
0%
b11 *
0-
02
b11 6
#224870000000
1!
1%
1-
12
15
#224880000000
0!
0%
b100 *
0-
02
b100 6
#224890000000
1!
1%
1-
12
#224900000000
0!
0%
b101 *
0-
02
b101 6
#224910000000
1!
1%
1-
12
#224920000000
0!
0%
b110 *
0-
02
b110 6
#224930000000
1!
1%
1-
12
#224940000000
0!
0%
b111 *
0-
02
b111 6
#224950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#224960000000
0!
0%
b0 *
0-
02
b0 6
#224970000000
1!
1%
1-
12
#224980000000
0!
0%
b1 *
0-
02
b1 6
#224990000000
1!
1%
1-
12
#225000000000
0!
0%
b10 *
0-
02
b10 6
#225010000000
1!
1%
1-
12
#225020000000
0!
0%
b11 *
0-
02
b11 6
#225030000000
1!
1%
1-
12
15
#225040000000
0!
0%
b100 *
0-
02
b100 6
#225050000000
1!
1%
1-
12
#225060000000
0!
0%
b101 *
0-
02
b101 6
#225070000000
1!
1%
1-
12
#225080000000
0!
0%
b110 *
0-
02
b110 6
#225090000000
1!
1%
1-
12
#225100000000
0!
0%
b111 *
0-
02
b111 6
#225110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#225120000000
0!
0%
b0 *
0-
02
b0 6
#225130000000
1!
1%
1-
12
#225140000000
0!
0%
b1 *
0-
02
b1 6
#225150000000
1!
1%
1-
12
#225160000000
0!
0%
b10 *
0-
02
b10 6
#225170000000
1!
1%
1-
12
#225180000000
0!
0%
b11 *
0-
02
b11 6
#225190000000
1!
1%
1-
12
15
#225200000000
0!
0%
b100 *
0-
02
b100 6
#225210000000
1!
1%
1-
12
#225220000000
0!
0%
b101 *
0-
02
b101 6
#225230000000
1!
1%
1-
12
#225240000000
0!
0%
b110 *
0-
02
b110 6
#225250000000
1!
1%
1-
12
#225260000000
0!
0%
b111 *
0-
02
b111 6
#225270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#225280000000
0!
0%
b0 *
0-
02
b0 6
#225290000000
1!
1%
1-
12
#225300000000
0!
0%
b1 *
0-
02
b1 6
#225310000000
1!
1%
1-
12
#225320000000
0!
0%
b10 *
0-
02
b10 6
#225330000000
1!
1%
1-
12
#225340000000
0!
0%
b11 *
0-
02
b11 6
#225350000000
1!
1%
1-
12
15
#225360000000
0!
0%
b100 *
0-
02
b100 6
#225370000000
1!
1%
1-
12
#225380000000
0!
0%
b101 *
0-
02
b101 6
#225390000000
1!
1%
1-
12
#225400000000
0!
0%
b110 *
0-
02
b110 6
#225410000000
1!
1%
1-
12
#225420000000
0!
0%
b111 *
0-
02
b111 6
#225430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#225440000000
0!
0%
b0 *
0-
02
b0 6
#225450000000
1!
1%
1-
12
#225460000000
0!
0%
b1 *
0-
02
b1 6
#225470000000
1!
1%
1-
12
#225480000000
0!
0%
b10 *
0-
02
b10 6
#225490000000
1!
1%
1-
12
#225500000000
0!
0%
b11 *
0-
02
b11 6
#225510000000
1!
1%
1-
12
15
#225520000000
0!
0%
b100 *
0-
02
b100 6
#225530000000
1!
1%
1-
12
#225540000000
0!
0%
b101 *
0-
02
b101 6
#225550000000
1!
1%
1-
12
#225560000000
0!
0%
b110 *
0-
02
b110 6
#225570000000
1!
1%
1-
12
#225580000000
0!
0%
b111 *
0-
02
b111 6
#225590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#225600000000
0!
0%
b0 *
0-
02
b0 6
#225610000000
1!
1%
1-
12
#225620000000
0!
0%
b1 *
0-
02
b1 6
#225630000000
1!
1%
1-
12
#225640000000
0!
0%
b10 *
0-
02
b10 6
#225650000000
1!
1%
1-
12
#225660000000
0!
0%
b11 *
0-
02
b11 6
#225670000000
1!
1%
1-
12
15
#225680000000
0!
0%
b100 *
0-
02
b100 6
#225690000000
1!
1%
1-
12
#225700000000
0!
0%
b101 *
0-
02
b101 6
#225710000000
1!
1%
1-
12
#225720000000
0!
0%
b110 *
0-
02
b110 6
#225730000000
1!
1%
1-
12
#225740000000
0!
0%
b111 *
0-
02
b111 6
#225750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#225760000000
0!
0%
b0 *
0-
02
b0 6
#225770000000
1!
1%
1-
12
#225780000000
0!
0%
b1 *
0-
02
b1 6
#225790000000
1!
1%
1-
12
#225800000000
0!
0%
b10 *
0-
02
b10 6
#225810000000
1!
1%
1-
12
#225820000000
0!
0%
b11 *
0-
02
b11 6
#225830000000
1!
1%
1-
12
15
#225840000000
0!
0%
b100 *
0-
02
b100 6
#225850000000
1!
1%
1-
12
#225860000000
0!
0%
b101 *
0-
02
b101 6
#225870000000
1!
1%
1-
12
#225880000000
0!
0%
b110 *
0-
02
b110 6
#225890000000
1!
1%
1-
12
#225900000000
0!
0%
b111 *
0-
02
b111 6
#225910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#225920000000
0!
0%
b0 *
0-
02
b0 6
#225930000000
1!
1%
1-
12
#225940000000
0!
0%
b1 *
0-
02
b1 6
#225950000000
1!
1%
1-
12
#225960000000
0!
0%
b10 *
0-
02
b10 6
#225970000000
1!
1%
1-
12
#225980000000
0!
0%
b11 *
0-
02
b11 6
#225990000000
1!
1%
1-
12
15
#226000000000
0!
0%
b100 *
0-
02
b100 6
#226010000000
1!
1%
1-
12
#226020000000
0!
0%
b101 *
0-
02
b101 6
#226030000000
1!
1%
1-
12
#226040000000
0!
0%
b110 *
0-
02
b110 6
#226050000000
1!
1%
1-
12
#226060000000
0!
0%
b111 *
0-
02
b111 6
#226070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#226080000000
0!
0%
b0 *
0-
02
b0 6
#226090000000
1!
1%
1-
12
#226100000000
0!
0%
b1 *
0-
02
b1 6
#226110000000
1!
1%
1-
12
#226120000000
0!
0%
b10 *
0-
02
b10 6
#226130000000
1!
1%
1-
12
#226140000000
0!
0%
b11 *
0-
02
b11 6
#226150000000
1!
1%
1-
12
15
#226160000000
0!
0%
b100 *
0-
02
b100 6
#226170000000
1!
1%
1-
12
#226180000000
0!
0%
b101 *
0-
02
b101 6
#226190000000
1!
1%
1-
12
#226200000000
0!
0%
b110 *
0-
02
b110 6
#226210000000
1!
1%
1-
12
#226220000000
0!
0%
b111 *
0-
02
b111 6
#226230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#226240000000
0!
0%
b0 *
0-
02
b0 6
#226250000000
1!
1%
1-
12
#226260000000
0!
0%
b1 *
0-
02
b1 6
#226270000000
1!
1%
1-
12
#226280000000
0!
0%
b10 *
0-
02
b10 6
#226290000000
1!
1%
1-
12
#226300000000
0!
0%
b11 *
0-
02
b11 6
#226310000000
1!
1%
1-
12
15
#226320000000
0!
0%
b100 *
0-
02
b100 6
#226330000000
1!
1%
1-
12
#226340000000
0!
0%
b101 *
0-
02
b101 6
#226350000000
1!
1%
1-
12
#226360000000
0!
0%
b110 *
0-
02
b110 6
#226370000000
1!
1%
1-
12
#226380000000
0!
0%
b111 *
0-
02
b111 6
#226390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#226400000000
0!
0%
b0 *
0-
02
b0 6
#226410000000
1!
1%
1-
12
#226420000000
0!
0%
b1 *
0-
02
b1 6
#226430000000
1!
1%
1-
12
#226440000000
0!
0%
b10 *
0-
02
b10 6
#226450000000
1!
1%
1-
12
#226460000000
0!
0%
b11 *
0-
02
b11 6
#226470000000
1!
1%
1-
12
15
#226480000000
0!
0%
b100 *
0-
02
b100 6
#226490000000
1!
1%
1-
12
#226500000000
0!
0%
b101 *
0-
02
b101 6
#226510000000
1!
1%
1-
12
#226520000000
0!
0%
b110 *
0-
02
b110 6
#226530000000
1!
1%
1-
12
#226540000000
0!
0%
b111 *
0-
02
b111 6
#226550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#226560000000
0!
0%
b0 *
0-
02
b0 6
#226570000000
1!
1%
1-
12
#226580000000
0!
0%
b1 *
0-
02
b1 6
#226590000000
1!
1%
1-
12
#226600000000
0!
0%
b10 *
0-
02
b10 6
#226610000000
1!
1%
1-
12
#226620000000
0!
0%
b11 *
0-
02
b11 6
#226630000000
1!
1%
1-
12
15
#226640000000
0!
0%
b100 *
0-
02
b100 6
#226650000000
1!
1%
1-
12
#226660000000
0!
0%
b101 *
0-
02
b101 6
#226670000000
1!
1%
1-
12
#226680000000
0!
0%
b110 *
0-
02
b110 6
#226690000000
1!
1%
1-
12
#226700000000
0!
0%
b111 *
0-
02
b111 6
#226710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#226720000000
0!
0%
b0 *
0-
02
b0 6
#226730000000
1!
1%
1-
12
#226740000000
0!
0%
b1 *
0-
02
b1 6
#226750000000
1!
1%
1-
12
#226760000000
0!
0%
b10 *
0-
02
b10 6
#226770000000
1!
1%
1-
12
#226780000000
0!
0%
b11 *
0-
02
b11 6
#226790000000
1!
1%
1-
12
15
#226800000000
0!
0%
b100 *
0-
02
b100 6
#226810000000
1!
1%
1-
12
#226820000000
0!
0%
b101 *
0-
02
b101 6
#226830000000
1!
1%
1-
12
#226840000000
0!
0%
b110 *
0-
02
b110 6
#226850000000
1!
1%
1-
12
#226860000000
0!
0%
b111 *
0-
02
b111 6
#226870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#226880000000
0!
0%
b0 *
0-
02
b0 6
#226890000000
1!
1%
1-
12
#226900000000
0!
0%
b1 *
0-
02
b1 6
#226910000000
1!
1%
1-
12
#226920000000
0!
0%
b10 *
0-
02
b10 6
#226930000000
1!
1%
1-
12
#226940000000
0!
0%
b11 *
0-
02
b11 6
#226950000000
1!
1%
1-
12
15
#226960000000
0!
0%
b100 *
0-
02
b100 6
#226970000000
1!
1%
1-
12
#226980000000
0!
0%
b101 *
0-
02
b101 6
#226990000000
1!
1%
1-
12
#227000000000
0!
0%
b110 *
0-
02
b110 6
#227010000000
1!
1%
1-
12
#227020000000
0!
0%
b111 *
0-
02
b111 6
#227030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#227040000000
0!
0%
b0 *
0-
02
b0 6
#227050000000
1!
1%
1-
12
#227060000000
0!
0%
b1 *
0-
02
b1 6
#227070000000
1!
1%
1-
12
#227080000000
0!
0%
b10 *
0-
02
b10 6
#227090000000
1!
1%
1-
12
#227100000000
0!
0%
b11 *
0-
02
b11 6
#227110000000
1!
1%
1-
12
15
#227120000000
0!
0%
b100 *
0-
02
b100 6
#227130000000
1!
1%
1-
12
#227140000000
0!
0%
b101 *
0-
02
b101 6
#227150000000
1!
1%
1-
12
#227160000000
0!
0%
b110 *
0-
02
b110 6
#227170000000
1!
1%
1-
12
#227180000000
0!
0%
b111 *
0-
02
b111 6
#227190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#227200000000
0!
0%
b0 *
0-
02
b0 6
#227210000000
1!
1%
1-
12
#227220000000
0!
0%
b1 *
0-
02
b1 6
#227230000000
1!
1%
1-
12
#227240000000
0!
0%
b10 *
0-
02
b10 6
#227250000000
1!
1%
1-
12
#227260000000
0!
0%
b11 *
0-
02
b11 6
#227270000000
1!
1%
1-
12
15
#227280000000
0!
0%
b100 *
0-
02
b100 6
#227290000000
1!
1%
1-
12
#227300000000
0!
0%
b101 *
0-
02
b101 6
#227310000000
1!
1%
1-
12
#227320000000
0!
0%
b110 *
0-
02
b110 6
#227330000000
1!
1%
1-
12
#227340000000
0!
0%
b111 *
0-
02
b111 6
#227350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#227360000000
0!
0%
b0 *
0-
02
b0 6
#227370000000
1!
1%
1-
12
#227380000000
0!
0%
b1 *
0-
02
b1 6
#227390000000
1!
1%
1-
12
#227400000000
0!
0%
b10 *
0-
02
b10 6
#227410000000
1!
1%
1-
12
#227420000000
0!
0%
b11 *
0-
02
b11 6
#227430000000
1!
1%
1-
12
15
#227440000000
0!
0%
b100 *
0-
02
b100 6
#227450000000
1!
1%
1-
12
#227460000000
0!
0%
b101 *
0-
02
b101 6
#227470000000
1!
1%
1-
12
#227480000000
0!
0%
b110 *
0-
02
b110 6
#227490000000
1!
1%
1-
12
#227500000000
0!
0%
b111 *
0-
02
b111 6
#227510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#227520000000
0!
0%
b0 *
0-
02
b0 6
#227530000000
1!
1%
1-
12
#227540000000
0!
0%
b1 *
0-
02
b1 6
#227550000000
1!
1%
1-
12
#227560000000
0!
0%
b10 *
0-
02
b10 6
#227570000000
1!
1%
1-
12
#227580000000
0!
0%
b11 *
0-
02
b11 6
#227590000000
1!
1%
1-
12
15
#227600000000
0!
0%
b100 *
0-
02
b100 6
#227610000000
1!
1%
1-
12
#227620000000
0!
0%
b101 *
0-
02
b101 6
#227630000000
1!
1%
1-
12
#227640000000
0!
0%
b110 *
0-
02
b110 6
#227650000000
1!
1%
1-
12
#227660000000
0!
0%
b111 *
0-
02
b111 6
#227670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#227680000000
0!
0%
b0 *
0-
02
b0 6
#227690000000
1!
1%
1-
12
#227700000000
0!
0%
b1 *
0-
02
b1 6
#227710000000
1!
1%
1-
12
#227720000000
0!
0%
b10 *
0-
02
b10 6
#227730000000
1!
1%
1-
12
#227740000000
0!
0%
b11 *
0-
02
b11 6
#227750000000
1!
1%
1-
12
15
#227760000000
0!
0%
b100 *
0-
02
b100 6
#227770000000
1!
1%
1-
12
#227780000000
0!
0%
b101 *
0-
02
b101 6
#227790000000
1!
1%
1-
12
#227800000000
0!
0%
b110 *
0-
02
b110 6
#227810000000
1!
1%
1-
12
#227820000000
0!
0%
b111 *
0-
02
b111 6
#227830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#227840000000
0!
0%
b0 *
0-
02
b0 6
#227850000000
1!
1%
1-
12
#227860000000
0!
0%
b1 *
0-
02
b1 6
#227870000000
1!
1%
1-
12
#227880000000
0!
0%
b10 *
0-
02
b10 6
#227890000000
1!
1%
1-
12
#227900000000
0!
0%
b11 *
0-
02
b11 6
#227910000000
1!
1%
1-
12
15
#227920000000
0!
0%
b100 *
0-
02
b100 6
#227930000000
1!
1%
1-
12
#227940000000
0!
0%
b101 *
0-
02
b101 6
#227950000000
1!
1%
1-
12
#227960000000
0!
0%
b110 *
0-
02
b110 6
#227970000000
1!
1%
1-
12
#227980000000
0!
0%
b111 *
0-
02
b111 6
#227990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#228000000000
0!
0%
b0 *
0-
02
b0 6
#228010000000
1!
1%
1-
12
#228020000000
0!
0%
b1 *
0-
02
b1 6
#228030000000
1!
1%
1-
12
#228040000000
0!
0%
b10 *
0-
02
b10 6
#228050000000
1!
1%
1-
12
#228060000000
0!
0%
b11 *
0-
02
b11 6
#228070000000
1!
1%
1-
12
15
#228080000000
0!
0%
b100 *
0-
02
b100 6
#228090000000
1!
1%
1-
12
#228100000000
0!
0%
b101 *
0-
02
b101 6
#228110000000
1!
1%
1-
12
#228120000000
0!
0%
b110 *
0-
02
b110 6
#228130000000
1!
1%
1-
12
#228140000000
0!
0%
b111 *
0-
02
b111 6
#228150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#228160000000
0!
0%
b0 *
0-
02
b0 6
#228170000000
1!
1%
1-
12
#228180000000
0!
0%
b1 *
0-
02
b1 6
#228190000000
1!
1%
1-
12
#228200000000
0!
0%
b10 *
0-
02
b10 6
#228210000000
1!
1%
1-
12
#228220000000
0!
0%
b11 *
0-
02
b11 6
#228230000000
1!
1%
1-
12
15
#228240000000
0!
0%
b100 *
0-
02
b100 6
#228250000000
1!
1%
1-
12
#228260000000
0!
0%
b101 *
0-
02
b101 6
#228270000000
1!
1%
1-
12
#228280000000
0!
0%
b110 *
0-
02
b110 6
#228290000000
1!
1%
1-
12
#228300000000
0!
0%
b111 *
0-
02
b111 6
#228310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#228320000000
0!
0%
b0 *
0-
02
b0 6
#228330000000
1!
1%
1-
12
#228340000000
0!
0%
b1 *
0-
02
b1 6
#228350000000
1!
1%
1-
12
#228360000000
0!
0%
b10 *
0-
02
b10 6
#228370000000
1!
1%
1-
12
#228380000000
0!
0%
b11 *
0-
02
b11 6
#228390000000
1!
1%
1-
12
15
#228400000000
0!
0%
b100 *
0-
02
b100 6
#228410000000
1!
1%
1-
12
#228420000000
0!
0%
b101 *
0-
02
b101 6
#228430000000
1!
1%
1-
12
#228440000000
0!
0%
b110 *
0-
02
b110 6
#228450000000
1!
1%
1-
12
#228460000000
0!
0%
b111 *
0-
02
b111 6
#228470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#228480000000
0!
0%
b0 *
0-
02
b0 6
#228490000000
1!
1%
1-
12
#228500000000
0!
0%
b1 *
0-
02
b1 6
#228510000000
1!
1%
1-
12
#228520000000
0!
0%
b10 *
0-
02
b10 6
#228530000000
1!
1%
1-
12
#228540000000
0!
0%
b11 *
0-
02
b11 6
#228550000000
1!
1%
1-
12
15
#228560000000
0!
0%
b100 *
0-
02
b100 6
#228570000000
1!
1%
1-
12
#228580000000
0!
0%
b101 *
0-
02
b101 6
#228590000000
1!
1%
1-
12
#228600000000
0!
0%
b110 *
0-
02
b110 6
#228610000000
1!
1%
1-
12
#228620000000
0!
0%
b111 *
0-
02
b111 6
#228630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#228640000000
0!
0%
b0 *
0-
02
b0 6
#228650000000
1!
1%
1-
12
#228660000000
0!
0%
b1 *
0-
02
b1 6
#228670000000
1!
1%
1-
12
#228680000000
0!
0%
b10 *
0-
02
b10 6
#228690000000
1!
1%
1-
12
#228700000000
0!
0%
b11 *
0-
02
b11 6
#228710000000
1!
1%
1-
12
15
#228720000000
0!
0%
b100 *
0-
02
b100 6
#228730000000
1!
1%
1-
12
#228740000000
0!
0%
b101 *
0-
02
b101 6
#228750000000
1!
1%
1-
12
#228760000000
0!
0%
b110 *
0-
02
b110 6
#228770000000
1!
1%
1-
12
#228780000000
0!
0%
b111 *
0-
02
b111 6
#228790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#228800000000
0!
0%
b0 *
0-
02
b0 6
#228810000000
1!
1%
1-
12
#228820000000
0!
0%
b1 *
0-
02
b1 6
#228830000000
1!
1%
1-
12
#228840000000
0!
0%
b10 *
0-
02
b10 6
#228850000000
1!
1%
1-
12
#228860000000
0!
0%
b11 *
0-
02
b11 6
#228870000000
1!
1%
1-
12
15
#228880000000
0!
0%
b100 *
0-
02
b100 6
#228890000000
1!
1%
1-
12
#228900000000
0!
0%
b101 *
0-
02
b101 6
#228910000000
1!
1%
1-
12
#228920000000
0!
0%
b110 *
0-
02
b110 6
#228930000000
1!
1%
1-
12
#228940000000
0!
0%
b111 *
0-
02
b111 6
#228950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#228960000000
0!
0%
b0 *
0-
02
b0 6
#228970000000
1!
1%
1-
12
#228980000000
0!
0%
b1 *
0-
02
b1 6
#228990000000
1!
1%
1-
12
#229000000000
0!
0%
b10 *
0-
02
b10 6
#229010000000
1!
1%
1-
12
#229020000000
0!
0%
b11 *
0-
02
b11 6
#229030000000
1!
1%
1-
12
15
#229040000000
0!
0%
b100 *
0-
02
b100 6
#229050000000
1!
1%
1-
12
#229060000000
0!
0%
b101 *
0-
02
b101 6
#229070000000
1!
1%
1-
12
#229080000000
0!
0%
b110 *
0-
02
b110 6
#229090000000
1!
1%
1-
12
#229100000000
0!
0%
b111 *
0-
02
b111 6
#229110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#229120000000
0!
0%
b0 *
0-
02
b0 6
#229130000000
1!
1%
1-
12
#229140000000
0!
0%
b1 *
0-
02
b1 6
#229150000000
1!
1%
1-
12
#229160000000
0!
0%
b10 *
0-
02
b10 6
#229170000000
1!
1%
1-
12
#229180000000
0!
0%
b11 *
0-
02
b11 6
#229190000000
1!
1%
1-
12
15
#229200000000
0!
0%
b100 *
0-
02
b100 6
#229210000000
1!
1%
1-
12
#229220000000
0!
0%
b101 *
0-
02
b101 6
#229230000000
1!
1%
1-
12
#229240000000
0!
0%
b110 *
0-
02
b110 6
#229250000000
1!
1%
1-
12
#229260000000
0!
0%
b111 *
0-
02
b111 6
#229270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#229280000000
0!
0%
b0 *
0-
02
b0 6
#229290000000
1!
1%
1-
12
#229300000000
0!
0%
b1 *
0-
02
b1 6
#229310000000
1!
1%
1-
12
#229320000000
0!
0%
b10 *
0-
02
b10 6
#229330000000
1!
1%
1-
12
#229340000000
0!
0%
b11 *
0-
02
b11 6
#229350000000
1!
1%
1-
12
15
#229360000000
0!
0%
b100 *
0-
02
b100 6
#229370000000
1!
1%
1-
12
#229380000000
0!
0%
b101 *
0-
02
b101 6
#229390000000
1!
1%
1-
12
#229400000000
0!
0%
b110 *
0-
02
b110 6
#229410000000
1!
1%
1-
12
#229420000000
0!
0%
b111 *
0-
02
b111 6
#229430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#229440000000
0!
0%
b0 *
0-
02
b0 6
#229450000000
1!
1%
1-
12
#229460000000
0!
0%
b1 *
0-
02
b1 6
#229470000000
1!
1%
1-
12
#229480000000
0!
0%
b10 *
0-
02
b10 6
#229490000000
1!
1%
1-
12
#229500000000
0!
0%
b11 *
0-
02
b11 6
#229510000000
1!
1%
1-
12
15
#229520000000
0!
0%
b100 *
0-
02
b100 6
#229530000000
1!
1%
1-
12
#229540000000
0!
0%
b101 *
0-
02
b101 6
#229550000000
1!
1%
1-
12
#229560000000
0!
0%
b110 *
0-
02
b110 6
#229570000000
1!
1%
1-
12
#229580000000
0!
0%
b111 *
0-
02
b111 6
#229590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#229600000000
0!
0%
b0 *
0-
02
b0 6
#229610000000
1!
1%
1-
12
#229620000000
0!
0%
b1 *
0-
02
b1 6
#229630000000
1!
1%
1-
12
#229640000000
0!
0%
b10 *
0-
02
b10 6
#229650000000
1!
1%
1-
12
#229660000000
0!
0%
b11 *
0-
02
b11 6
#229670000000
1!
1%
1-
12
15
#229680000000
0!
0%
b100 *
0-
02
b100 6
#229690000000
1!
1%
1-
12
#229700000000
0!
0%
b101 *
0-
02
b101 6
#229710000000
1!
1%
1-
12
#229720000000
0!
0%
b110 *
0-
02
b110 6
#229730000000
1!
1%
1-
12
#229740000000
0!
0%
b111 *
0-
02
b111 6
#229750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#229760000000
0!
0%
b0 *
0-
02
b0 6
#229770000000
1!
1%
1-
12
#229780000000
0!
0%
b1 *
0-
02
b1 6
#229790000000
1!
1%
1-
12
#229800000000
0!
0%
b10 *
0-
02
b10 6
#229810000000
1!
1%
1-
12
#229820000000
0!
0%
b11 *
0-
02
b11 6
#229830000000
1!
1%
1-
12
15
#229840000000
0!
0%
b100 *
0-
02
b100 6
#229850000000
1!
1%
1-
12
#229860000000
0!
0%
b101 *
0-
02
b101 6
#229870000000
1!
1%
1-
12
#229880000000
0!
0%
b110 *
0-
02
b110 6
#229890000000
1!
1%
1-
12
#229900000000
0!
0%
b111 *
0-
02
b111 6
#229910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#229920000000
0!
0%
b0 *
0-
02
b0 6
#229930000000
1!
1%
1-
12
#229940000000
0!
0%
b1 *
0-
02
b1 6
#229950000000
1!
1%
1-
12
#229960000000
0!
0%
b10 *
0-
02
b10 6
#229970000000
1!
1%
1-
12
#229980000000
0!
0%
b11 *
0-
02
b11 6
#229990000000
1!
1%
1-
12
15
#230000000000
0!
0%
b100 *
0-
02
b100 6
#230010000000
1!
1%
1-
12
#230020000000
0!
0%
b101 *
0-
02
b101 6
#230030000000
1!
1%
1-
12
#230040000000
0!
0%
b110 *
0-
02
b110 6
#230050000000
1!
1%
1-
12
#230060000000
0!
0%
b111 *
0-
02
b111 6
#230070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#230080000000
0!
0%
b0 *
0-
02
b0 6
#230090000000
1!
1%
1-
12
#230100000000
0!
0%
b1 *
0-
02
b1 6
#230110000000
1!
1%
1-
12
#230120000000
0!
0%
b10 *
0-
02
b10 6
#230130000000
1!
1%
1-
12
#230140000000
0!
0%
b11 *
0-
02
b11 6
#230150000000
1!
1%
1-
12
15
#230160000000
0!
0%
b100 *
0-
02
b100 6
#230170000000
1!
1%
1-
12
#230180000000
0!
0%
b101 *
0-
02
b101 6
#230190000000
1!
1%
1-
12
#230200000000
0!
0%
b110 *
0-
02
b110 6
#230210000000
1!
1%
1-
12
#230220000000
0!
0%
b111 *
0-
02
b111 6
#230230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#230240000000
0!
0%
b0 *
0-
02
b0 6
#230250000000
1!
1%
1-
12
#230260000000
0!
0%
b1 *
0-
02
b1 6
#230270000000
1!
1%
1-
12
#230280000000
0!
0%
b10 *
0-
02
b10 6
#230290000000
1!
1%
1-
12
#230300000000
0!
0%
b11 *
0-
02
b11 6
#230310000000
1!
1%
1-
12
15
#230320000000
0!
0%
b100 *
0-
02
b100 6
#230330000000
1!
1%
1-
12
#230340000000
0!
0%
b101 *
0-
02
b101 6
#230350000000
1!
1%
1-
12
#230360000000
0!
0%
b110 *
0-
02
b110 6
#230370000000
1!
1%
1-
12
#230380000000
0!
0%
b111 *
0-
02
b111 6
#230390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#230400000000
0!
0%
b0 *
0-
02
b0 6
#230410000000
1!
1%
1-
12
#230420000000
0!
0%
b1 *
0-
02
b1 6
#230430000000
1!
1%
1-
12
#230440000000
0!
0%
b10 *
0-
02
b10 6
#230450000000
1!
1%
1-
12
#230460000000
0!
0%
b11 *
0-
02
b11 6
#230470000000
1!
1%
1-
12
15
#230480000000
0!
0%
b100 *
0-
02
b100 6
#230490000000
1!
1%
1-
12
#230500000000
0!
0%
b101 *
0-
02
b101 6
#230510000000
1!
1%
1-
12
#230520000000
0!
0%
b110 *
0-
02
b110 6
#230530000000
1!
1%
1-
12
#230540000000
0!
0%
b111 *
0-
02
b111 6
#230550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#230560000000
0!
0%
b0 *
0-
02
b0 6
#230570000000
1!
1%
1-
12
#230580000000
0!
0%
b1 *
0-
02
b1 6
#230590000000
1!
1%
1-
12
#230600000000
0!
0%
b10 *
0-
02
b10 6
#230610000000
1!
1%
1-
12
#230620000000
0!
0%
b11 *
0-
02
b11 6
#230630000000
1!
1%
1-
12
15
#230640000000
0!
0%
b100 *
0-
02
b100 6
#230650000000
1!
1%
1-
12
#230660000000
0!
0%
b101 *
0-
02
b101 6
#230670000000
1!
1%
1-
12
#230680000000
0!
0%
b110 *
0-
02
b110 6
#230690000000
1!
1%
1-
12
#230700000000
0!
0%
b111 *
0-
02
b111 6
#230710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#230720000000
0!
0%
b0 *
0-
02
b0 6
#230730000000
1!
1%
1-
12
#230740000000
0!
0%
b1 *
0-
02
b1 6
#230750000000
1!
1%
1-
12
#230760000000
0!
0%
b10 *
0-
02
b10 6
#230770000000
1!
1%
1-
12
#230780000000
0!
0%
b11 *
0-
02
b11 6
#230790000000
1!
1%
1-
12
15
#230800000000
0!
0%
b100 *
0-
02
b100 6
#230810000000
1!
1%
1-
12
#230820000000
0!
0%
b101 *
0-
02
b101 6
#230830000000
1!
1%
1-
12
#230840000000
0!
0%
b110 *
0-
02
b110 6
#230850000000
1!
1%
1-
12
#230860000000
0!
0%
b111 *
0-
02
b111 6
#230870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#230880000000
0!
0%
b0 *
0-
02
b0 6
#230890000000
1!
1%
1-
12
#230900000000
0!
0%
b1 *
0-
02
b1 6
#230910000000
1!
1%
1-
12
#230920000000
0!
0%
b10 *
0-
02
b10 6
#230930000000
1!
1%
1-
12
#230940000000
0!
0%
b11 *
0-
02
b11 6
#230950000000
1!
1%
1-
12
15
#230960000000
0!
0%
b100 *
0-
02
b100 6
#230970000000
1!
1%
1-
12
#230980000000
0!
0%
b101 *
0-
02
b101 6
#230990000000
1!
1%
1-
12
#231000000000
0!
0%
b110 *
0-
02
b110 6
#231010000000
1!
1%
1-
12
#231020000000
0!
0%
b111 *
0-
02
b111 6
#231030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#231040000000
0!
0%
b0 *
0-
02
b0 6
#231050000000
1!
1%
1-
12
#231060000000
0!
0%
b1 *
0-
02
b1 6
#231070000000
1!
1%
1-
12
#231080000000
0!
0%
b10 *
0-
02
b10 6
#231090000000
1!
1%
1-
12
#231100000000
0!
0%
b11 *
0-
02
b11 6
#231110000000
1!
1%
1-
12
15
#231120000000
0!
0%
b100 *
0-
02
b100 6
#231130000000
1!
1%
1-
12
#231140000000
0!
0%
b101 *
0-
02
b101 6
#231150000000
1!
1%
1-
12
#231160000000
0!
0%
b110 *
0-
02
b110 6
#231170000000
1!
1%
1-
12
#231180000000
0!
0%
b111 *
0-
02
b111 6
#231190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#231200000000
0!
0%
b0 *
0-
02
b0 6
#231210000000
1!
1%
1-
12
#231220000000
0!
0%
b1 *
0-
02
b1 6
#231230000000
1!
1%
1-
12
#231240000000
0!
0%
b10 *
0-
02
b10 6
#231250000000
1!
1%
1-
12
#231260000000
0!
0%
b11 *
0-
02
b11 6
#231270000000
1!
1%
1-
12
15
#231280000000
0!
0%
b100 *
0-
02
b100 6
#231290000000
1!
1%
1-
12
#231300000000
0!
0%
b101 *
0-
02
b101 6
#231310000000
1!
1%
1-
12
#231320000000
0!
0%
b110 *
0-
02
b110 6
#231330000000
1!
1%
1-
12
#231340000000
0!
0%
b111 *
0-
02
b111 6
#231350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#231360000000
0!
0%
b0 *
0-
02
b0 6
#231370000000
1!
1%
1-
12
#231380000000
0!
0%
b1 *
0-
02
b1 6
#231390000000
1!
1%
1-
12
#231400000000
0!
0%
b10 *
0-
02
b10 6
#231410000000
1!
1%
1-
12
#231420000000
0!
0%
b11 *
0-
02
b11 6
#231430000000
1!
1%
1-
12
15
#231440000000
0!
0%
b100 *
0-
02
b100 6
#231450000000
1!
1%
1-
12
#231460000000
0!
0%
b101 *
0-
02
b101 6
#231470000000
1!
1%
1-
12
#231480000000
0!
0%
b110 *
0-
02
b110 6
#231490000000
1!
1%
1-
12
#231500000000
0!
0%
b111 *
0-
02
b111 6
#231510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#231520000000
0!
0%
b0 *
0-
02
b0 6
#231530000000
1!
1%
1-
12
#231540000000
0!
0%
b1 *
0-
02
b1 6
#231550000000
1!
1%
1-
12
#231560000000
0!
0%
b10 *
0-
02
b10 6
#231570000000
1!
1%
1-
12
#231580000000
0!
0%
b11 *
0-
02
b11 6
#231590000000
1!
1%
1-
12
15
#231600000000
0!
0%
b100 *
0-
02
b100 6
#231610000000
1!
1%
1-
12
#231620000000
0!
0%
b101 *
0-
02
b101 6
#231630000000
1!
1%
1-
12
#231640000000
0!
0%
b110 *
0-
02
b110 6
#231650000000
1!
1%
1-
12
#231660000000
0!
0%
b111 *
0-
02
b111 6
#231670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#231680000000
0!
0%
b0 *
0-
02
b0 6
#231690000000
1!
1%
1-
12
#231700000000
0!
0%
b1 *
0-
02
b1 6
#231710000000
1!
1%
1-
12
#231720000000
0!
0%
b10 *
0-
02
b10 6
#231730000000
1!
1%
1-
12
#231740000000
0!
0%
b11 *
0-
02
b11 6
#231750000000
1!
1%
1-
12
15
#231760000000
0!
0%
b100 *
0-
02
b100 6
#231770000000
1!
1%
1-
12
#231780000000
0!
0%
b101 *
0-
02
b101 6
#231790000000
1!
1%
1-
12
#231800000000
0!
0%
b110 *
0-
02
b110 6
#231810000000
1!
1%
1-
12
#231820000000
0!
0%
b111 *
0-
02
b111 6
#231830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#231840000000
0!
0%
b0 *
0-
02
b0 6
#231850000000
1!
1%
1-
12
#231860000000
0!
0%
b1 *
0-
02
b1 6
#231870000000
1!
1%
1-
12
#231880000000
0!
0%
b10 *
0-
02
b10 6
#231890000000
1!
1%
1-
12
#231900000000
0!
0%
b11 *
0-
02
b11 6
#231910000000
1!
1%
1-
12
15
#231920000000
0!
0%
b100 *
0-
02
b100 6
#231930000000
1!
1%
1-
12
#231940000000
0!
0%
b101 *
0-
02
b101 6
#231950000000
1!
1%
1-
12
#231960000000
0!
0%
b110 *
0-
02
b110 6
#231970000000
1!
1%
1-
12
#231980000000
0!
0%
b111 *
0-
02
b111 6
#231990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#232000000000
0!
0%
b0 *
0-
02
b0 6
#232010000000
1!
1%
1-
12
#232020000000
0!
0%
b1 *
0-
02
b1 6
#232030000000
1!
1%
1-
12
#232040000000
0!
0%
b10 *
0-
02
b10 6
#232050000000
1!
1%
1-
12
#232060000000
0!
0%
b11 *
0-
02
b11 6
#232070000000
1!
1%
1-
12
15
#232080000000
0!
0%
b100 *
0-
02
b100 6
#232090000000
1!
1%
1-
12
#232100000000
0!
0%
b101 *
0-
02
b101 6
#232110000000
1!
1%
1-
12
#232120000000
0!
0%
b110 *
0-
02
b110 6
#232130000000
1!
1%
1-
12
#232140000000
0!
0%
b111 *
0-
02
b111 6
#232150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#232160000000
0!
0%
b0 *
0-
02
b0 6
#232170000000
1!
1%
1-
12
#232180000000
0!
0%
b1 *
0-
02
b1 6
#232190000000
1!
1%
1-
12
#232200000000
0!
0%
b10 *
0-
02
b10 6
#232210000000
1!
1%
1-
12
#232220000000
0!
0%
b11 *
0-
02
b11 6
#232230000000
1!
1%
1-
12
15
#232240000000
0!
0%
b100 *
0-
02
b100 6
#232250000000
1!
1%
1-
12
#232260000000
0!
0%
b101 *
0-
02
b101 6
#232270000000
1!
1%
1-
12
#232280000000
0!
0%
b110 *
0-
02
b110 6
#232290000000
1!
1%
1-
12
#232300000000
0!
0%
b111 *
0-
02
b111 6
#232310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#232320000000
0!
0%
b0 *
0-
02
b0 6
#232330000000
1!
1%
1-
12
#232340000000
0!
0%
b1 *
0-
02
b1 6
#232350000000
1!
1%
1-
12
#232360000000
0!
0%
b10 *
0-
02
b10 6
#232370000000
1!
1%
1-
12
#232380000000
0!
0%
b11 *
0-
02
b11 6
#232390000000
1!
1%
1-
12
15
#232400000000
0!
0%
b100 *
0-
02
b100 6
#232410000000
1!
1%
1-
12
#232420000000
0!
0%
b101 *
0-
02
b101 6
#232430000000
1!
1%
1-
12
#232440000000
0!
0%
b110 *
0-
02
b110 6
#232450000000
1!
1%
1-
12
#232460000000
0!
0%
b111 *
0-
02
b111 6
#232470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#232480000000
0!
0%
b0 *
0-
02
b0 6
#232490000000
1!
1%
1-
12
#232500000000
0!
0%
b1 *
0-
02
b1 6
#232510000000
1!
1%
1-
12
#232520000000
0!
0%
b10 *
0-
02
b10 6
#232530000000
1!
1%
1-
12
#232540000000
0!
0%
b11 *
0-
02
b11 6
#232550000000
1!
1%
1-
12
15
#232560000000
0!
0%
b100 *
0-
02
b100 6
#232570000000
1!
1%
1-
12
#232580000000
0!
0%
b101 *
0-
02
b101 6
#232590000000
1!
1%
1-
12
#232600000000
0!
0%
b110 *
0-
02
b110 6
#232610000000
1!
1%
1-
12
#232620000000
0!
0%
b111 *
0-
02
b111 6
#232630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#232640000000
0!
0%
b0 *
0-
02
b0 6
#232650000000
1!
1%
1-
12
#232660000000
0!
0%
b1 *
0-
02
b1 6
#232670000000
1!
1%
1-
12
#232680000000
0!
0%
b10 *
0-
02
b10 6
#232690000000
1!
1%
1-
12
#232700000000
0!
0%
b11 *
0-
02
b11 6
#232710000000
1!
1%
1-
12
15
#232720000000
0!
0%
b100 *
0-
02
b100 6
#232730000000
1!
1%
1-
12
#232740000000
0!
0%
b101 *
0-
02
b101 6
#232750000000
1!
1%
1-
12
#232760000000
0!
0%
b110 *
0-
02
b110 6
#232770000000
1!
1%
1-
12
#232780000000
0!
0%
b111 *
0-
02
b111 6
#232790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#232800000000
0!
0%
b0 *
0-
02
b0 6
#232810000000
1!
1%
1-
12
#232820000000
0!
0%
b1 *
0-
02
b1 6
#232830000000
1!
1%
1-
12
#232840000000
0!
0%
b10 *
0-
02
b10 6
#232850000000
1!
1%
1-
12
#232860000000
0!
0%
b11 *
0-
02
b11 6
#232870000000
1!
1%
1-
12
15
#232880000000
0!
0%
b100 *
0-
02
b100 6
#232890000000
1!
1%
1-
12
#232900000000
0!
0%
b101 *
0-
02
b101 6
#232910000000
1!
1%
1-
12
#232920000000
0!
0%
b110 *
0-
02
b110 6
#232930000000
1!
1%
1-
12
#232940000000
0!
0%
b111 *
0-
02
b111 6
#232950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#232960000000
0!
0%
b0 *
0-
02
b0 6
#232970000000
1!
1%
1-
12
#232980000000
0!
0%
b1 *
0-
02
b1 6
#232990000000
1!
1%
1-
12
#233000000000
0!
0%
b10 *
0-
02
b10 6
#233010000000
1!
1%
1-
12
#233020000000
0!
0%
b11 *
0-
02
b11 6
#233030000000
1!
1%
1-
12
15
#233040000000
0!
0%
b100 *
0-
02
b100 6
#233050000000
1!
1%
1-
12
#233060000000
0!
0%
b101 *
0-
02
b101 6
#233070000000
1!
1%
1-
12
#233080000000
0!
0%
b110 *
0-
02
b110 6
#233090000000
1!
1%
1-
12
#233100000000
0!
0%
b111 *
0-
02
b111 6
#233110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#233120000000
0!
0%
b0 *
0-
02
b0 6
#233130000000
1!
1%
1-
12
#233140000000
0!
0%
b1 *
0-
02
b1 6
#233150000000
1!
1%
1-
12
#233160000000
0!
0%
b10 *
0-
02
b10 6
#233170000000
1!
1%
1-
12
#233180000000
0!
0%
b11 *
0-
02
b11 6
#233190000000
1!
1%
1-
12
15
#233200000000
0!
0%
b100 *
0-
02
b100 6
#233210000000
1!
1%
1-
12
#233220000000
0!
0%
b101 *
0-
02
b101 6
#233230000000
1!
1%
1-
12
#233240000000
0!
0%
b110 *
0-
02
b110 6
#233250000000
1!
1%
1-
12
#233260000000
0!
0%
b111 *
0-
02
b111 6
#233270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#233280000000
0!
0%
b0 *
0-
02
b0 6
#233290000000
1!
1%
1-
12
#233300000000
0!
0%
b1 *
0-
02
b1 6
#233310000000
1!
1%
1-
12
#233320000000
0!
0%
b10 *
0-
02
b10 6
#233330000000
1!
1%
1-
12
#233340000000
0!
0%
b11 *
0-
02
b11 6
#233350000000
1!
1%
1-
12
15
#233360000000
0!
0%
b100 *
0-
02
b100 6
#233370000000
1!
1%
1-
12
#233380000000
0!
0%
b101 *
0-
02
b101 6
#233390000000
1!
1%
1-
12
#233400000000
0!
0%
b110 *
0-
02
b110 6
#233410000000
1!
1%
1-
12
#233420000000
0!
0%
b111 *
0-
02
b111 6
#233430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#233440000000
0!
0%
b0 *
0-
02
b0 6
#233450000000
1!
1%
1-
12
#233460000000
0!
0%
b1 *
0-
02
b1 6
#233470000000
1!
1%
1-
12
#233480000000
0!
0%
b10 *
0-
02
b10 6
#233490000000
1!
1%
1-
12
#233500000000
0!
0%
b11 *
0-
02
b11 6
#233510000000
1!
1%
1-
12
15
#233520000000
0!
0%
b100 *
0-
02
b100 6
#233530000000
1!
1%
1-
12
#233540000000
0!
0%
b101 *
0-
02
b101 6
#233550000000
1!
1%
1-
12
#233560000000
0!
0%
b110 *
0-
02
b110 6
#233570000000
1!
1%
1-
12
#233580000000
0!
0%
b111 *
0-
02
b111 6
#233590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#233600000000
0!
0%
b0 *
0-
02
b0 6
#233610000000
1!
1%
1-
12
#233620000000
0!
0%
b1 *
0-
02
b1 6
#233630000000
1!
1%
1-
12
#233640000000
0!
0%
b10 *
0-
02
b10 6
#233650000000
1!
1%
1-
12
#233660000000
0!
0%
b11 *
0-
02
b11 6
#233670000000
1!
1%
1-
12
15
#233680000000
0!
0%
b100 *
0-
02
b100 6
#233690000000
1!
1%
1-
12
#233700000000
0!
0%
b101 *
0-
02
b101 6
#233710000000
1!
1%
1-
12
#233720000000
0!
0%
b110 *
0-
02
b110 6
#233730000000
1!
1%
1-
12
#233740000000
0!
0%
b111 *
0-
02
b111 6
#233750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#233760000000
0!
0%
b0 *
0-
02
b0 6
#233770000000
1!
1%
1-
12
#233780000000
0!
0%
b1 *
0-
02
b1 6
#233790000000
1!
1%
1-
12
#233800000000
0!
0%
b10 *
0-
02
b10 6
#233810000000
1!
1%
1-
12
#233820000000
0!
0%
b11 *
0-
02
b11 6
#233830000000
1!
1%
1-
12
15
#233840000000
0!
0%
b100 *
0-
02
b100 6
#233850000000
1!
1%
1-
12
#233860000000
0!
0%
b101 *
0-
02
b101 6
#233870000000
1!
1%
1-
12
#233880000000
0!
0%
b110 *
0-
02
b110 6
#233890000000
1!
1%
1-
12
#233900000000
0!
0%
b111 *
0-
02
b111 6
#233910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#233920000000
0!
0%
b0 *
0-
02
b0 6
#233930000000
1!
1%
1-
12
#233940000000
0!
0%
b1 *
0-
02
b1 6
#233950000000
1!
1%
1-
12
#233960000000
0!
0%
b10 *
0-
02
b10 6
#233970000000
1!
1%
1-
12
#233980000000
0!
0%
b11 *
0-
02
b11 6
#233990000000
1!
1%
1-
12
15
#234000000000
0!
0%
b100 *
0-
02
b100 6
#234010000000
1!
1%
1-
12
#234020000000
0!
0%
b101 *
0-
02
b101 6
#234030000000
1!
1%
1-
12
#234040000000
0!
0%
b110 *
0-
02
b110 6
#234050000000
1!
1%
1-
12
#234060000000
0!
0%
b111 *
0-
02
b111 6
#234070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#234080000000
0!
0%
b0 *
0-
02
b0 6
#234090000000
1!
1%
1-
12
#234100000000
0!
0%
b1 *
0-
02
b1 6
#234110000000
1!
1%
1-
12
#234120000000
0!
0%
b10 *
0-
02
b10 6
#234130000000
1!
1%
1-
12
#234140000000
0!
0%
b11 *
0-
02
b11 6
#234150000000
1!
1%
1-
12
15
#234160000000
0!
0%
b100 *
0-
02
b100 6
#234170000000
1!
1%
1-
12
#234180000000
0!
0%
b101 *
0-
02
b101 6
#234190000000
1!
1%
1-
12
#234200000000
0!
0%
b110 *
0-
02
b110 6
#234210000000
1!
1%
1-
12
#234220000000
0!
0%
b111 *
0-
02
b111 6
#234230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#234240000000
0!
0%
b0 *
0-
02
b0 6
#234250000000
1!
1%
1-
12
#234260000000
0!
0%
b1 *
0-
02
b1 6
#234270000000
1!
1%
1-
12
#234280000000
0!
0%
b10 *
0-
02
b10 6
#234290000000
1!
1%
1-
12
#234300000000
0!
0%
b11 *
0-
02
b11 6
#234310000000
1!
1%
1-
12
15
#234320000000
0!
0%
b100 *
0-
02
b100 6
#234330000000
1!
1%
1-
12
#234340000000
0!
0%
b101 *
0-
02
b101 6
#234350000000
1!
1%
1-
12
#234360000000
0!
0%
b110 *
0-
02
b110 6
#234370000000
1!
1%
1-
12
#234380000000
0!
0%
b111 *
0-
02
b111 6
#234390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#234400000000
0!
0%
b0 *
0-
02
b0 6
#234410000000
1!
1%
1-
12
#234420000000
0!
0%
b1 *
0-
02
b1 6
#234430000000
1!
1%
1-
12
#234440000000
0!
0%
b10 *
0-
02
b10 6
#234450000000
1!
1%
1-
12
#234460000000
0!
0%
b11 *
0-
02
b11 6
#234470000000
1!
1%
1-
12
15
#234480000000
0!
0%
b100 *
0-
02
b100 6
#234490000000
1!
1%
1-
12
#234500000000
0!
0%
b101 *
0-
02
b101 6
#234510000000
1!
1%
1-
12
#234520000000
0!
0%
b110 *
0-
02
b110 6
#234530000000
1!
1%
1-
12
#234540000000
0!
0%
b111 *
0-
02
b111 6
#234550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#234560000000
0!
0%
b0 *
0-
02
b0 6
#234570000000
1!
1%
1-
12
#234580000000
0!
0%
b1 *
0-
02
b1 6
#234590000000
1!
1%
1-
12
#234600000000
0!
0%
b10 *
0-
02
b10 6
#234610000000
1!
1%
1-
12
#234620000000
0!
0%
b11 *
0-
02
b11 6
#234630000000
1!
1%
1-
12
15
#234640000000
0!
0%
b100 *
0-
02
b100 6
#234650000000
1!
1%
1-
12
#234660000000
0!
0%
b101 *
0-
02
b101 6
#234670000000
1!
1%
1-
12
#234680000000
0!
0%
b110 *
0-
02
b110 6
#234690000000
1!
1%
1-
12
#234700000000
0!
0%
b111 *
0-
02
b111 6
#234710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#234720000000
0!
0%
b0 *
0-
02
b0 6
#234730000000
1!
1%
1-
12
#234740000000
0!
0%
b1 *
0-
02
b1 6
#234750000000
1!
1%
1-
12
#234760000000
0!
0%
b10 *
0-
02
b10 6
#234770000000
1!
1%
1-
12
#234780000000
0!
0%
b11 *
0-
02
b11 6
#234790000000
1!
1%
1-
12
15
#234800000000
0!
0%
b100 *
0-
02
b100 6
#234810000000
1!
1%
1-
12
#234820000000
0!
0%
b101 *
0-
02
b101 6
#234830000000
1!
1%
1-
12
#234840000000
0!
0%
b110 *
0-
02
b110 6
#234850000000
1!
1%
1-
12
#234860000000
0!
0%
b111 *
0-
02
b111 6
#234870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#234880000000
0!
0%
b0 *
0-
02
b0 6
#234890000000
1!
1%
1-
12
#234900000000
0!
0%
b1 *
0-
02
b1 6
#234910000000
1!
1%
1-
12
#234920000000
0!
0%
b10 *
0-
02
b10 6
#234930000000
1!
1%
1-
12
#234940000000
0!
0%
b11 *
0-
02
b11 6
#234950000000
1!
1%
1-
12
15
#234960000000
0!
0%
b100 *
0-
02
b100 6
#234970000000
1!
1%
1-
12
#234980000000
0!
0%
b101 *
0-
02
b101 6
#234990000000
1!
1%
1-
12
#235000000000
0!
0%
b110 *
0-
02
b110 6
#235010000000
1!
1%
1-
12
#235020000000
0!
0%
b111 *
0-
02
b111 6
#235030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#235040000000
0!
0%
b0 *
0-
02
b0 6
#235050000000
1!
1%
1-
12
#235060000000
0!
0%
b1 *
0-
02
b1 6
#235070000000
1!
1%
1-
12
#235080000000
0!
0%
b10 *
0-
02
b10 6
#235090000000
1!
1%
1-
12
#235100000000
0!
0%
b11 *
0-
02
b11 6
#235110000000
1!
1%
1-
12
15
#235120000000
0!
0%
b100 *
0-
02
b100 6
#235130000000
1!
1%
1-
12
#235140000000
0!
0%
b101 *
0-
02
b101 6
#235150000000
1!
1%
1-
12
#235160000000
0!
0%
b110 *
0-
02
b110 6
#235170000000
1!
1%
1-
12
#235180000000
0!
0%
b111 *
0-
02
b111 6
#235190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#235200000000
0!
0%
b0 *
0-
02
b0 6
#235210000000
1!
1%
1-
12
#235220000000
0!
0%
b1 *
0-
02
b1 6
#235230000000
1!
1%
1-
12
#235240000000
0!
0%
b10 *
0-
02
b10 6
#235250000000
1!
1%
1-
12
#235260000000
0!
0%
b11 *
0-
02
b11 6
#235270000000
1!
1%
1-
12
15
#235280000000
0!
0%
b100 *
0-
02
b100 6
#235290000000
1!
1%
1-
12
#235300000000
0!
0%
b101 *
0-
02
b101 6
#235310000000
1!
1%
1-
12
#235320000000
0!
0%
b110 *
0-
02
b110 6
#235330000000
1!
1%
1-
12
#235340000000
0!
0%
b111 *
0-
02
b111 6
#235350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#235360000000
0!
0%
b0 *
0-
02
b0 6
#235370000000
1!
1%
1-
12
#235380000000
0!
0%
b1 *
0-
02
b1 6
#235390000000
1!
1%
1-
12
#235400000000
0!
0%
b10 *
0-
02
b10 6
#235410000000
1!
1%
1-
12
#235420000000
0!
0%
b11 *
0-
02
b11 6
#235430000000
1!
1%
1-
12
15
#235440000000
0!
0%
b100 *
0-
02
b100 6
#235450000000
1!
1%
1-
12
#235460000000
0!
0%
b101 *
0-
02
b101 6
#235470000000
1!
1%
1-
12
#235480000000
0!
0%
b110 *
0-
02
b110 6
#235490000000
1!
1%
1-
12
#235500000000
0!
0%
b111 *
0-
02
b111 6
#235510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#235520000000
0!
0%
b0 *
0-
02
b0 6
#235530000000
1!
1%
1-
12
#235540000000
0!
0%
b1 *
0-
02
b1 6
#235550000000
1!
1%
1-
12
#235560000000
0!
0%
b10 *
0-
02
b10 6
#235570000000
1!
1%
1-
12
#235580000000
0!
0%
b11 *
0-
02
b11 6
#235590000000
1!
1%
1-
12
15
#235600000000
0!
0%
b100 *
0-
02
b100 6
#235610000000
1!
1%
1-
12
#235620000000
0!
0%
b101 *
0-
02
b101 6
#235630000000
1!
1%
1-
12
#235640000000
0!
0%
b110 *
0-
02
b110 6
#235650000000
1!
1%
1-
12
#235660000000
0!
0%
b111 *
0-
02
b111 6
#235670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#235680000000
0!
0%
b0 *
0-
02
b0 6
#235690000000
1!
1%
1-
12
#235700000000
0!
0%
b1 *
0-
02
b1 6
#235710000000
1!
1%
1-
12
#235720000000
0!
0%
b10 *
0-
02
b10 6
#235730000000
1!
1%
1-
12
#235740000000
0!
0%
b11 *
0-
02
b11 6
#235750000000
1!
1%
1-
12
15
#235760000000
0!
0%
b100 *
0-
02
b100 6
#235770000000
1!
1%
1-
12
#235780000000
0!
0%
b101 *
0-
02
b101 6
#235790000000
1!
1%
1-
12
#235800000000
0!
0%
b110 *
0-
02
b110 6
#235810000000
1!
1%
1-
12
#235820000000
0!
0%
b111 *
0-
02
b111 6
#235830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#235840000000
0!
0%
b0 *
0-
02
b0 6
#235850000000
1!
1%
1-
12
#235860000000
0!
0%
b1 *
0-
02
b1 6
#235870000000
1!
1%
1-
12
#235880000000
0!
0%
b10 *
0-
02
b10 6
#235890000000
1!
1%
1-
12
#235900000000
0!
0%
b11 *
0-
02
b11 6
#235910000000
1!
1%
1-
12
15
#235920000000
0!
0%
b100 *
0-
02
b100 6
#235930000000
1!
1%
1-
12
#235940000000
0!
0%
b101 *
0-
02
b101 6
#235950000000
1!
1%
1-
12
#235960000000
0!
0%
b110 *
0-
02
b110 6
#235970000000
1!
1%
1-
12
#235980000000
0!
0%
b111 *
0-
02
b111 6
#235990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#236000000000
0!
0%
b0 *
0-
02
b0 6
#236010000000
1!
1%
1-
12
#236020000000
0!
0%
b1 *
0-
02
b1 6
#236030000000
1!
1%
1-
12
#236040000000
0!
0%
b10 *
0-
02
b10 6
#236050000000
1!
1%
1-
12
#236060000000
0!
0%
b11 *
0-
02
b11 6
#236070000000
1!
1%
1-
12
15
#236080000000
0!
0%
b100 *
0-
02
b100 6
#236090000000
1!
1%
1-
12
#236100000000
0!
0%
b101 *
0-
02
b101 6
#236110000000
1!
1%
1-
12
#236120000000
0!
0%
b110 *
0-
02
b110 6
#236130000000
1!
1%
1-
12
#236140000000
0!
0%
b111 *
0-
02
b111 6
#236150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#236160000000
0!
0%
b0 *
0-
02
b0 6
#236170000000
1!
1%
1-
12
#236180000000
0!
0%
b1 *
0-
02
b1 6
#236190000000
1!
1%
1-
12
#236200000000
0!
0%
b10 *
0-
02
b10 6
#236210000000
1!
1%
1-
12
#236220000000
0!
0%
b11 *
0-
02
b11 6
#236230000000
1!
1%
1-
12
15
#236240000000
0!
0%
b100 *
0-
02
b100 6
#236250000000
1!
1%
1-
12
#236260000000
0!
0%
b101 *
0-
02
b101 6
#236270000000
1!
1%
1-
12
#236280000000
0!
0%
b110 *
0-
02
b110 6
#236290000000
1!
1%
1-
12
#236300000000
0!
0%
b111 *
0-
02
b111 6
#236310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#236320000000
0!
0%
b0 *
0-
02
b0 6
#236330000000
1!
1%
1-
12
#236340000000
0!
0%
b1 *
0-
02
b1 6
#236350000000
1!
1%
1-
12
#236360000000
0!
0%
b10 *
0-
02
b10 6
#236370000000
1!
1%
1-
12
#236380000000
0!
0%
b11 *
0-
02
b11 6
#236390000000
1!
1%
1-
12
15
#236400000000
0!
0%
b100 *
0-
02
b100 6
#236410000000
1!
1%
1-
12
#236420000000
0!
0%
b101 *
0-
02
b101 6
#236430000000
1!
1%
1-
12
#236440000000
0!
0%
b110 *
0-
02
b110 6
#236450000000
1!
1%
1-
12
#236460000000
0!
0%
b111 *
0-
02
b111 6
#236470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#236480000000
0!
0%
b0 *
0-
02
b0 6
#236490000000
1!
1%
1-
12
#236500000000
0!
0%
b1 *
0-
02
b1 6
#236510000000
1!
1%
1-
12
#236520000000
0!
0%
b10 *
0-
02
b10 6
#236530000000
1!
1%
1-
12
#236540000000
0!
0%
b11 *
0-
02
b11 6
#236550000000
1!
1%
1-
12
15
#236560000000
0!
0%
b100 *
0-
02
b100 6
#236570000000
1!
1%
1-
12
#236580000000
0!
0%
b101 *
0-
02
b101 6
#236590000000
1!
1%
1-
12
#236600000000
0!
0%
b110 *
0-
02
b110 6
#236610000000
1!
1%
1-
12
#236620000000
0!
0%
b111 *
0-
02
b111 6
#236630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#236640000000
0!
0%
b0 *
0-
02
b0 6
#236650000000
1!
1%
1-
12
#236660000000
0!
0%
b1 *
0-
02
b1 6
#236670000000
1!
1%
1-
12
#236680000000
0!
0%
b10 *
0-
02
b10 6
#236690000000
1!
1%
1-
12
#236700000000
0!
0%
b11 *
0-
02
b11 6
#236710000000
1!
1%
1-
12
15
#236720000000
0!
0%
b100 *
0-
02
b100 6
#236730000000
1!
1%
1-
12
#236740000000
0!
0%
b101 *
0-
02
b101 6
#236750000000
1!
1%
1-
12
#236760000000
0!
0%
b110 *
0-
02
b110 6
#236770000000
1!
1%
1-
12
#236780000000
0!
0%
b111 *
0-
02
b111 6
#236790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#236800000000
0!
0%
b0 *
0-
02
b0 6
#236810000000
1!
1%
1-
12
#236820000000
0!
0%
b1 *
0-
02
b1 6
#236830000000
1!
1%
1-
12
#236840000000
0!
0%
b10 *
0-
02
b10 6
#236850000000
1!
1%
1-
12
#236860000000
0!
0%
b11 *
0-
02
b11 6
#236870000000
1!
1%
1-
12
15
#236880000000
0!
0%
b100 *
0-
02
b100 6
#236890000000
1!
1%
1-
12
#236900000000
0!
0%
b101 *
0-
02
b101 6
#236910000000
1!
1%
1-
12
#236920000000
0!
0%
b110 *
0-
02
b110 6
#236930000000
1!
1%
1-
12
#236940000000
0!
0%
b111 *
0-
02
b111 6
#236950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#236960000000
0!
0%
b0 *
0-
02
b0 6
#236970000000
1!
1%
1-
12
#236980000000
0!
0%
b1 *
0-
02
b1 6
#236990000000
1!
1%
1-
12
#237000000000
0!
0%
b10 *
0-
02
b10 6
#237010000000
1!
1%
1-
12
#237020000000
0!
0%
b11 *
0-
02
b11 6
#237030000000
1!
1%
1-
12
15
#237040000000
0!
0%
b100 *
0-
02
b100 6
#237050000000
1!
1%
1-
12
#237060000000
0!
0%
b101 *
0-
02
b101 6
#237070000000
1!
1%
1-
12
#237080000000
0!
0%
b110 *
0-
02
b110 6
#237090000000
1!
1%
1-
12
#237100000000
0!
0%
b111 *
0-
02
b111 6
#237110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#237120000000
0!
0%
b0 *
0-
02
b0 6
#237130000000
1!
1%
1-
12
#237140000000
0!
0%
b1 *
0-
02
b1 6
#237150000000
1!
1%
1-
12
#237160000000
0!
0%
b10 *
0-
02
b10 6
#237170000000
1!
1%
1-
12
#237180000000
0!
0%
b11 *
0-
02
b11 6
#237190000000
1!
1%
1-
12
15
#237200000000
0!
0%
b100 *
0-
02
b100 6
#237210000000
1!
1%
1-
12
#237220000000
0!
0%
b101 *
0-
02
b101 6
#237230000000
1!
1%
1-
12
#237240000000
0!
0%
b110 *
0-
02
b110 6
#237250000000
1!
1%
1-
12
#237260000000
0!
0%
b111 *
0-
02
b111 6
#237270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#237280000000
0!
0%
b0 *
0-
02
b0 6
#237290000000
1!
1%
1-
12
#237300000000
0!
0%
b1 *
0-
02
b1 6
#237310000000
1!
1%
1-
12
#237320000000
0!
0%
b10 *
0-
02
b10 6
#237330000000
1!
1%
1-
12
#237340000000
0!
0%
b11 *
0-
02
b11 6
#237350000000
1!
1%
1-
12
15
#237360000000
0!
0%
b100 *
0-
02
b100 6
#237370000000
1!
1%
1-
12
#237380000000
0!
0%
b101 *
0-
02
b101 6
#237390000000
1!
1%
1-
12
#237400000000
0!
0%
b110 *
0-
02
b110 6
#237410000000
1!
1%
1-
12
#237420000000
0!
0%
b111 *
0-
02
b111 6
#237430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#237440000000
0!
0%
b0 *
0-
02
b0 6
#237450000000
1!
1%
1-
12
#237460000000
0!
0%
b1 *
0-
02
b1 6
#237470000000
1!
1%
1-
12
#237480000000
0!
0%
b10 *
0-
02
b10 6
#237490000000
1!
1%
1-
12
#237500000000
0!
0%
b11 *
0-
02
b11 6
#237510000000
1!
1%
1-
12
15
#237520000000
0!
0%
b100 *
0-
02
b100 6
#237530000000
1!
1%
1-
12
#237540000000
0!
0%
b101 *
0-
02
b101 6
#237550000000
1!
1%
1-
12
#237560000000
0!
0%
b110 *
0-
02
b110 6
#237570000000
1!
1%
1-
12
#237580000000
0!
0%
b111 *
0-
02
b111 6
#237590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#237600000000
0!
0%
b0 *
0-
02
b0 6
#237610000000
1!
1%
1-
12
#237620000000
0!
0%
b1 *
0-
02
b1 6
#237630000000
1!
1%
1-
12
#237640000000
0!
0%
b10 *
0-
02
b10 6
#237650000000
1!
1%
1-
12
#237660000000
0!
0%
b11 *
0-
02
b11 6
#237670000000
1!
1%
1-
12
15
#237680000000
0!
0%
b100 *
0-
02
b100 6
#237690000000
1!
1%
1-
12
#237700000000
0!
0%
b101 *
0-
02
b101 6
#237710000000
1!
1%
1-
12
#237720000000
0!
0%
b110 *
0-
02
b110 6
#237730000000
1!
1%
1-
12
#237740000000
0!
0%
b111 *
0-
02
b111 6
#237750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#237760000000
0!
0%
b0 *
0-
02
b0 6
#237770000000
1!
1%
1-
12
#237780000000
0!
0%
b1 *
0-
02
b1 6
#237790000000
1!
1%
1-
12
#237800000000
0!
0%
b10 *
0-
02
b10 6
#237810000000
1!
1%
1-
12
#237820000000
0!
0%
b11 *
0-
02
b11 6
#237830000000
1!
1%
1-
12
15
#237840000000
0!
0%
b100 *
0-
02
b100 6
#237850000000
1!
1%
1-
12
#237860000000
0!
0%
b101 *
0-
02
b101 6
#237870000000
1!
1%
1-
12
#237880000000
0!
0%
b110 *
0-
02
b110 6
#237890000000
1!
1%
1-
12
#237900000000
0!
0%
b111 *
0-
02
b111 6
#237910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#237920000000
0!
0%
b0 *
0-
02
b0 6
#237930000000
1!
1%
1-
12
#237940000000
0!
0%
b1 *
0-
02
b1 6
#237950000000
1!
1%
1-
12
#237960000000
0!
0%
b10 *
0-
02
b10 6
#237970000000
1!
1%
1-
12
#237980000000
0!
0%
b11 *
0-
02
b11 6
#237990000000
1!
1%
1-
12
15
#238000000000
0!
0%
b100 *
0-
02
b100 6
#238010000000
1!
1%
1-
12
#238020000000
0!
0%
b101 *
0-
02
b101 6
#238030000000
1!
1%
1-
12
#238040000000
0!
0%
b110 *
0-
02
b110 6
#238050000000
1!
1%
1-
12
#238060000000
0!
0%
b111 *
0-
02
b111 6
#238070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#238080000000
0!
0%
b0 *
0-
02
b0 6
#238090000000
1!
1%
1-
12
#238100000000
0!
0%
b1 *
0-
02
b1 6
#238110000000
1!
1%
1-
12
#238120000000
0!
0%
b10 *
0-
02
b10 6
#238130000000
1!
1%
1-
12
#238140000000
0!
0%
b11 *
0-
02
b11 6
#238150000000
1!
1%
1-
12
15
#238160000000
0!
0%
b100 *
0-
02
b100 6
#238170000000
1!
1%
1-
12
#238180000000
0!
0%
b101 *
0-
02
b101 6
#238190000000
1!
1%
1-
12
#238200000000
0!
0%
b110 *
0-
02
b110 6
#238210000000
1!
1%
1-
12
#238220000000
0!
0%
b111 *
0-
02
b111 6
#238230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#238240000000
0!
0%
b0 *
0-
02
b0 6
#238250000000
1!
1%
1-
12
#238260000000
0!
0%
b1 *
0-
02
b1 6
#238270000000
1!
1%
1-
12
#238280000000
0!
0%
b10 *
0-
02
b10 6
#238290000000
1!
1%
1-
12
#238300000000
0!
0%
b11 *
0-
02
b11 6
#238310000000
1!
1%
1-
12
15
#238320000000
0!
0%
b100 *
0-
02
b100 6
#238330000000
1!
1%
1-
12
#238340000000
0!
0%
b101 *
0-
02
b101 6
#238350000000
1!
1%
1-
12
#238360000000
0!
0%
b110 *
0-
02
b110 6
#238370000000
1!
1%
1-
12
#238380000000
0!
0%
b111 *
0-
02
b111 6
#238390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#238400000000
0!
0%
b0 *
0-
02
b0 6
#238410000000
1!
1%
1-
12
#238420000000
0!
0%
b1 *
0-
02
b1 6
#238430000000
1!
1%
1-
12
#238440000000
0!
0%
b10 *
0-
02
b10 6
#238450000000
1!
1%
1-
12
#238460000000
0!
0%
b11 *
0-
02
b11 6
#238470000000
1!
1%
1-
12
15
#238480000000
0!
0%
b100 *
0-
02
b100 6
#238490000000
1!
1%
1-
12
#238500000000
0!
0%
b101 *
0-
02
b101 6
#238510000000
1!
1%
1-
12
#238520000000
0!
0%
b110 *
0-
02
b110 6
#238530000000
1!
1%
1-
12
#238540000000
0!
0%
b111 *
0-
02
b111 6
#238550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#238560000000
0!
0%
b0 *
0-
02
b0 6
#238570000000
1!
1%
1-
12
#238580000000
0!
0%
b1 *
0-
02
b1 6
#238590000000
1!
1%
1-
12
#238600000000
0!
0%
b10 *
0-
02
b10 6
#238610000000
1!
1%
1-
12
#238620000000
0!
0%
b11 *
0-
02
b11 6
#238630000000
1!
1%
1-
12
15
#238640000000
0!
0%
b100 *
0-
02
b100 6
#238650000000
1!
1%
1-
12
#238660000000
0!
0%
b101 *
0-
02
b101 6
#238670000000
1!
1%
1-
12
#238680000000
0!
0%
b110 *
0-
02
b110 6
#238690000000
1!
1%
1-
12
#238700000000
0!
0%
b111 *
0-
02
b111 6
#238710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#238720000000
0!
0%
b0 *
0-
02
b0 6
#238730000000
1!
1%
1-
12
#238740000000
0!
0%
b1 *
0-
02
b1 6
#238750000000
1!
1%
1-
12
#238760000000
0!
0%
b10 *
0-
02
b10 6
#238770000000
1!
1%
1-
12
#238780000000
0!
0%
b11 *
0-
02
b11 6
#238790000000
1!
1%
1-
12
15
#238800000000
0!
0%
b100 *
0-
02
b100 6
#238810000000
1!
1%
1-
12
#238820000000
0!
0%
b101 *
0-
02
b101 6
#238830000000
1!
1%
1-
12
#238840000000
0!
0%
b110 *
0-
02
b110 6
#238850000000
1!
1%
1-
12
#238860000000
0!
0%
b111 *
0-
02
b111 6
#238870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#238880000000
0!
0%
b0 *
0-
02
b0 6
#238890000000
1!
1%
1-
12
#238900000000
0!
0%
b1 *
0-
02
b1 6
#238910000000
1!
1%
1-
12
#238920000000
0!
0%
b10 *
0-
02
b10 6
#238930000000
1!
1%
1-
12
#238940000000
0!
0%
b11 *
0-
02
b11 6
#238950000000
1!
1%
1-
12
15
#238960000000
0!
0%
b100 *
0-
02
b100 6
#238970000000
1!
1%
1-
12
#238980000000
0!
0%
b101 *
0-
02
b101 6
#238990000000
1!
1%
1-
12
#239000000000
0!
0%
b110 *
0-
02
b110 6
#239010000000
1!
1%
1-
12
#239020000000
0!
0%
b111 *
0-
02
b111 6
#239030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#239040000000
0!
0%
b0 *
0-
02
b0 6
#239050000000
1!
1%
1-
12
#239060000000
0!
0%
b1 *
0-
02
b1 6
#239070000000
1!
1%
1-
12
#239080000000
0!
0%
b10 *
0-
02
b10 6
#239090000000
1!
1%
1-
12
#239100000000
0!
0%
b11 *
0-
02
b11 6
#239110000000
1!
1%
1-
12
15
#239120000000
0!
0%
b100 *
0-
02
b100 6
#239130000000
1!
1%
1-
12
#239140000000
0!
0%
b101 *
0-
02
b101 6
#239150000000
1!
1%
1-
12
#239160000000
0!
0%
b110 *
0-
02
b110 6
#239170000000
1!
1%
1-
12
#239180000000
0!
0%
b111 *
0-
02
b111 6
#239190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#239200000000
0!
0%
b0 *
0-
02
b0 6
#239210000000
1!
1%
1-
12
#239220000000
0!
0%
b1 *
0-
02
b1 6
#239230000000
1!
1%
1-
12
#239240000000
0!
0%
b10 *
0-
02
b10 6
#239250000000
1!
1%
1-
12
#239260000000
0!
0%
b11 *
0-
02
b11 6
#239270000000
1!
1%
1-
12
15
#239280000000
0!
0%
b100 *
0-
02
b100 6
#239290000000
1!
1%
1-
12
#239300000000
0!
0%
b101 *
0-
02
b101 6
#239310000000
1!
1%
1-
12
#239320000000
0!
0%
b110 *
0-
02
b110 6
#239330000000
1!
1%
1-
12
#239340000000
0!
0%
b111 *
0-
02
b111 6
#239350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#239360000000
0!
0%
b0 *
0-
02
b0 6
#239370000000
1!
1%
1-
12
#239380000000
0!
0%
b1 *
0-
02
b1 6
#239390000000
1!
1%
1-
12
#239400000000
0!
0%
b10 *
0-
02
b10 6
#239410000000
1!
1%
1-
12
#239420000000
0!
0%
b11 *
0-
02
b11 6
#239430000000
1!
1%
1-
12
15
#239440000000
0!
0%
b100 *
0-
02
b100 6
#239450000000
1!
1%
1-
12
#239460000000
0!
0%
b101 *
0-
02
b101 6
#239470000000
1!
1%
1-
12
#239480000000
0!
0%
b110 *
0-
02
b110 6
#239490000000
1!
1%
1-
12
#239500000000
0!
0%
b111 *
0-
02
b111 6
#239510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#239520000000
0!
0%
b0 *
0-
02
b0 6
#239530000000
1!
1%
1-
12
#239540000000
0!
0%
b1 *
0-
02
b1 6
#239550000000
1!
1%
1-
12
#239560000000
0!
0%
b10 *
0-
02
b10 6
#239570000000
1!
1%
1-
12
#239580000000
0!
0%
b11 *
0-
02
b11 6
#239590000000
1!
1%
1-
12
15
#239600000000
0!
0%
b100 *
0-
02
b100 6
#239610000000
1!
1%
1-
12
#239620000000
0!
0%
b101 *
0-
02
b101 6
#239630000000
1!
1%
1-
12
#239640000000
0!
0%
b110 *
0-
02
b110 6
#239650000000
1!
1%
1-
12
#239660000000
0!
0%
b111 *
0-
02
b111 6
#239670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#239680000000
0!
0%
b0 *
0-
02
b0 6
#239690000000
1!
1%
1-
12
#239700000000
0!
0%
b1 *
0-
02
b1 6
#239710000000
1!
1%
1-
12
#239720000000
0!
0%
b10 *
0-
02
b10 6
#239730000000
1!
1%
1-
12
#239740000000
0!
0%
b11 *
0-
02
b11 6
#239750000000
1!
1%
1-
12
15
#239760000000
0!
0%
b100 *
0-
02
b100 6
#239770000000
1!
1%
1-
12
#239780000000
0!
0%
b101 *
0-
02
b101 6
#239790000000
1!
1%
1-
12
#239800000000
0!
0%
b110 *
0-
02
b110 6
#239810000000
1!
1%
1-
12
#239820000000
0!
0%
b111 *
0-
02
b111 6
#239830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#239840000000
0!
0%
b0 *
0-
02
b0 6
#239850000000
1!
1%
1-
12
#239860000000
0!
0%
b1 *
0-
02
b1 6
#239870000000
1!
1%
1-
12
#239880000000
0!
0%
b10 *
0-
02
b10 6
#239890000000
1!
1%
1-
12
#239900000000
0!
0%
b11 *
0-
02
b11 6
#239910000000
1!
1%
1-
12
15
#239920000000
0!
0%
b100 *
0-
02
b100 6
#239930000000
1!
1%
1-
12
#239940000000
0!
0%
b101 *
0-
02
b101 6
#239950000000
1!
1%
1-
12
#239960000000
0!
0%
b110 *
0-
02
b110 6
#239970000000
1!
1%
1-
12
#239980000000
0!
0%
b111 *
0-
02
b111 6
#239990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#240000000000
0!
0%
b0 *
0-
02
b0 6
#240010000000
1!
1%
1-
12
#240020000000
0!
0%
b1 *
0-
02
b1 6
#240030000000
1!
1%
1-
12
#240040000000
0!
0%
b10 *
0-
02
b10 6
#240050000000
1!
1%
1-
12
#240060000000
0!
0%
b11 *
0-
02
b11 6
#240070000000
1!
1%
1-
12
15
#240080000000
0!
0%
b100 *
0-
02
b100 6
#240090000000
1!
1%
1-
12
#240100000000
0!
0%
b101 *
0-
02
b101 6
#240110000000
1!
1%
1-
12
#240120000000
0!
0%
b110 *
0-
02
b110 6
#240130000000
1!
1%
1-
12
#240140000000
0!
0%
b111 *
0-
02
b111 6
#240150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#240160000000
0!
0%
b0 *
0-
02
b0 6
#240170000000
1!
1%
1-
12
#240180000000
0!
0%
b1 *
0-
02
b1 6
#240190000000
1!
1%
1-
12
#240200000000
0!
0%
b10 *
0-
02
b10 6
#240210000000
1!
1%
1-
12
#240220000000
0!
0%
b11 *
0-
02
b11 6
#240230000000
1!
1%
1-
12
15
#240240000000
0!
0%
b100 *
0-
02
b100 6
#240250000000
1!
1%
1-
12
#240260000000
0!
0%
b101 *
0-
02
b101 6
#240270000000
1!
1%
1-
12
#240280000000
0!
0%
b110 *
0-
02
b110 6
#240290000000
1!
1%
1-
12
#240300000000
0!
0%
b111 *
0-
02
b111 6
#240310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#240320000000
0!
0%
b0 *
0-
02
b0 6
#240330000000
1!
1%
1-
12
#240340000000
0!
0%
b1 *
0-
02
b1 6
#240350000000
1!
1%
1-
12
#240360000000
0!
0%
b10 *
0-
02
b10 6
#240370000000
1!
1%
1-
12
#240380000000
0!
0%
b11 *
0-
02
b11 6
#240390000000
1!
1%
1-
12
15
#240400000000
0!
0%
b100 *
0-
02
b100 6
#240410000000
1!
1%
1-
12
#240420000000
0!
0%
b101 *
0-
02
b101 6
#240430000000
1!
1%
1-
12
#240440000000
0!
0%
b110 *
0-
02
b110 6
#240450000000
1!
1%
1-
12
#240460000000
0!
0%
b111 *
0-
02
b111 6
#240470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#240480000000
0!
0%
b0 *
0-
02
b0 6
#240490000000
1!
1%
1-
12
#240500000000
0!
0%
b1 *
0-
02
b1 6
#240510000000
1!
1%
1-
12
#240520000000
0!
0%
b10 *
0-
02
b10 6
#240530000000
1!
1%
1-
12
#240540000000
0!
0%
b11 *
0-
02
b11 6
#240550000000
1!
1%
1-
12
15
#240560000000
0!
0%
b100 *
0-
02
b100 6
#240570000000
1!
1%
1-
12
#240580000000
0!
0%
b101 *
0-
02
b101 6
#240590000000
1!
1%
1-
12
#240600000000
0!
0%
b110 *
0-
02
b110 6
#240610000000
1!
1%
1-
12
#240620000000
0!
0%
b111 *
0-
02
b111 6
#240630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#240640000000
0!
0%
b0 *
0-
02
b0 6
#240650000000
1!
1%
1-
12
#240660000000
0!
0%
b1 *
0-
02
b1 6
#240670000000
1!
1%
1-
12
#240680000000
0!
0%
b10 *
0-
02
b10 6
#240690000000
1!
1%
1-
12
#240700000000
0!
0%
b11 *
0-
02
b11 6
#240710000000
1!
1%
1-
12
15
#240720000000
0!
0%
b100 *
0-
02
b100 6
#240730000000
1!
1%
1-
12
#240740000000
0!
0%
b101 *
0-
02
b101 6
#240750000000
1!
1%
1-
12
#240760000000
0!
0%
b110 *
0-
02
b110 6
#240770000000
1!
1%
1-
12
#240780000000
0!
0%
b111 *
0-
02
b111 6
#240790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#240800000000
0!
0%
b0 *
0-
02
b0 6
#240810000000
1!
1%
1-
12
#240820000000
0!
0%
b1 *
0-
02
b1 6
#240830000000
1!
1%
1-
12
#240840000000
0!
0%
b10 *
0-
02
b10 6
#240850000000
1!
1%
1-
12
#240860000000
0!
0%
b11 *
0-
02
b11 6
#240870000000
1!
1%
1-
12
15
#240880000000
0!
0%
b100 *
0-
02
b100 6
#240890000000
1!
1%
1-
12
#240900000000
0!
0%
b101 *
0-
02
b101 6
#240910000000
1!
1%
1-
12
#240920000000
0!
0%
b110 *
0-
02
b110 6
#240930000000
1!
1%
1-
12
#240940000000
0!
0%
b111 *
0-
02
b111 6
#240950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#240960000000
0!
0%
b0 *
0-
02
b0 6
#240970000000
1!
1%
1-
12
#240980000000
0!
0%
b1 *
0-
02
b1 6
#240990000000
1!
1%
1-
12
#241000000000
0!
0%
b10 *
0-
02
b10 6
#241010000000
1!
1%
1-
12
#241020000000
0!
0%
b11 *
0-
02
b11 6
#241030000000
1!
1%
1-
12
15
#241040000000
0!
0%
b100 *
0-
02
b100 6
#241050000000
1!
1%
1-
12
#241060000000
0!
0%
b101 *
0-
02
b101 6
#241070000000
1!
1%
1-
12
#241080000000
0!
0%
b110 *
0-
02
b110 6
#241090000000
1!
1%
1-
12
#241100000000
0!
0%
b111 *
0-
02
b111 6
#241110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#241120000000
0!
0%
b0 *
0-
02
b0 6
#241130000000
1!
1%
1-
12
#241140000000
0!
0%
b1 *
0-
02
b1 6
#241150000000
1!
1%
1-
12
#241160000000
0!
0%
b10 *
0-
02
b10 6
#241170000000
1!
1%
1-
12
#241180000000
0!
0%
b11 *
0-
02
b11 6
#241190000000
1!
1%
1-
12
15
#241200000000
0!
0%
b100 *
0-
02
b100 6
#241210000000
1!
1%
1-
12
#241220000000
0!
0%
b101 *
0-
02
b101 6
#241230000000
1!
1%
1-
12
#241240000000
0!
0%
b110 *
0-
02
b110 6
#241250000000
1!
1%
1-
12
#241260000000
0!
0%
b111 *
0-
02
b111 6
#241270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#241280000000
0!
0%
b0 *
0-
02
b0 6
#241290000000
1!
1%
1-
12
#241300000000
0!
0%
b1 *
0-
02
b1 6
#241310000000
1!
1%
1-
12
#241320000000
0!
0%
b10 *
0-
02
b10 6
#241330000000
1!
1%
1-
12
#241340000000
0!
0%
b11 *
0-
02
b11 6
#241350000000
1!
1%
1-
12
15
#241360000000
0!
0%
b100 *
0-
02
b100 6
#241370000000
1!
1%
1-
12
#241380000000
0!
0%
b101 *
0-
02
b101 6
#241390000000
1!
1%
1-
12
#241400000000
0!
0%
b110 *
0-
02
b110 6
#241410000000
1!
1%
1-
12
#241420000000
0!
0%
b111 *
0-
02
b111 6
#241430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#241440000000
0!
0%
b0 *
0-
02
b0 6
#241450000000
1!
1%
1-
12
#241460000000
0!
0%
b1 *
0-
02
b1 6
#241470000000
1!
1%
1-
12
#241480000000
0!
0%
b10 *
0-
02
b10 6
#241490000000
1!
1%
1-
12
#241500000000
0!
0%
b11 *
0-
02
b11 6
#241510000000
1!
1%
1-
12
15
#241520000000
0!
0%
b100 *
0-
02
b100 6
#241530000000
1!
1%
1-
12
#241540000000
0!
0%
b101 *
0-
02
b101 6
#241550000000
1!
1%
1-
12
#241560000000
0!
0%
b110 *
0-
02
b110 6
#241570000000
1!
1%
1-
12
#241580000000
0!
0%
b111 *
0-
02
b111 6
#241590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#241600000000
0!
0%
b0 *
0-
02
b0 6
#241610000000
1!
1%
1-
12
#241620000000
0!
0%
b1 *
0-
02
b1 6
#241630000000
1!
1%
1-
12
#241640000000
0!
0%
b10 *
0-
02
b10 6
#241650000000
1!
1%
1-
12
#241660000000
0!
0%
b11 *
0-
02
b11 6
#241670000000
1!
1%
1-
12
15
#241680000000
0!
0%
b100 *
0-
02
b100 6
#241690000000
1!
1%
1-
12
#241700000000
0!
0%
b101 *
0-
02
b101 6
#241710000000
1!
1%
1-
12
#241720000000
0!
0%
b110 *
0-
02
b110 6
#241730000000
1!
1%
1-
12
#241740000000
0!
0%
b111 *
0-
02
b111 6
#241750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#241760000000
0!
0%
b0 *
0-
02
b0 6
#241770000000
1!
1%
1-
12
#241780000000
0!
0%
b1 *
0-
02
b1 6
#241790000000
1!
1%
1-
12
#241800000000
0!
0%
b10 *
0-
02
b10 6
#241810000000
1!
1%
1-
12
#241820000000
0!
0%
b11 *
0-
02
b11 6
#241830000000
1!
1%
1-
12
15
#241840000000
0!
0%
b100 *
0-
02
b100 6
#241850000000
1!
1%
1-
12
#241860000000
0!
0%
b101 *
0-
02
b101 6
#241870000000
1!
1%
1-
12
#241880000000
0!
0%
b110 *
0-
02
b110 6
#241890000000
1!
1%
1-
12
#241900000000
0!
0%
b111 *
0-
02
b111 6
#241910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#241920000000
0!
0%
b0 *
0-
02
b0 6
#241930000000
1!
1%
1-
12
#241940000000
0!
0%
b1 *
0-
02
b1 6
#241950000000
1!
1%
1-
12
#241960000000
0!
0%
b10 *
0-
02
b10 6
#241970000000
1!
1%
1-
12
#241980000000
0!
0%
b11 *
0-
02
b11 6
#241990000000
1!
1%
1-
12
15
#242000000000
0!
0%
b100 *
0-
02
b100 6
#242010000000
1!
1%
1-
12
#242020000000
0!
0%
b101 *
0-
02
b101 6
#242030000000
1!
1%
1-
12
#242040000000
0!
0%
b110 *
0-
02
b110 6
#242050000000
1!
1%
1-
12
#242060000000
0!
0%
b111 *
0-
02
b111 6
#242070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#242080000000
0!
0%
b0 *
0-
02
b0 6
#242090000000
1!
1%
1-
12
#242100000000
0!
0%
b1 *
0-
02
b1 6
#242110000000
1!
1%
1-
12
#242120000000
0!
0%
b10 *
0-
02
b10 6
#242130000000
1!
1%
1-
12
#242140000000
0!
0%
b11 *
0-
02
b11 6
#242150000000
1!
1%
1-
12
15
#242160000000
0!
0%
b100 *
0-
02
b100 6
#242170000000
1!
1%
1-
12
#242180000000
0!
0%
b101 *
0-
02
b101 6
#242190000000
1!
1%
1-
12
#242200000000
0!
0%
b110 *
0-
02
b110 6
#242210000000
1!
1%
1-
12
#242220000000
0!
0%
b111 *
0-
02
b111 6
#242230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#242240000000
0!
0%
b0 *
0-
02
b0 6
#242250000000
1!
1%
1-
12
#242260000000
0!
0%
b1 *
0-
02
b1 6
#242270000000
1!
1%
1-
12
#242280000000
0!
0%
b10 *
0-
02
b10 6
#242290000000
1!
1%
1-
12
#242300000000
0!
0%
b11 *
0-
02
b11 6
#242310000000
1!
1%
1-
12
15
#242320000000
0!
0%
b100 *
0-
02
b100 6
#242330000000
1!
1%
1-
12
#242340000000
0!
0%
b101 *
0-
02
b101 6
#242350000000
1!
1%
1-
12
#242360000000
0!
0%
b110 *
0-
02
b110 6
#242370000000
1!
1%
1-
12
#242380000000
0!
0%
b111 *
0-
02
b111 6
#242390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#242400000000
0!
0%
b0 *
0-
02
b0 6
#242410000000
1!
1%
1-
12
#242420000000
0!
0%
b1 *
0-
02
b1 6
#242430000000
1!
1%
1-
12
#242440000000
0!
0%
b10 *
0-
02
b10 6
#242450000000
1!
1%
1-
12
#242460000000
0!
0%
b11 *
0-
02
b11 6
#242470000000
1!
1%
1-
12
15
#242480000000
0!
0%
b100 *
0-
02
b100 6
#242490000000
1!
1%
1-
12
#242500000000
0!
0%
b101 *
0-
02
b101 6
#242510000000
1!
1%
1-
12
#242520000000
0!
0%
b110 *
0-
02
b110 6
#242530000000
1!
1%
1-
12
#242540000000
0!
0%
b111 *
0-
02
b111 6
#242550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#242560000000
0!
0%
b0 *
0-
02
b0 6
#242570000000
1!
1%
1-
12
#242580000000
0!
0%
b1 *
0-
02
b1 6
#242590000000
1!
1%
1-
12
#242600000000
0!
0%
b10 *
0-
02
b10 6
#242610000000
1!
1%
1-
12
#242620000000
0!
0%
b11 *
0-
02
b11 6
#242630000000
1!
1%
1-
12
15
#242640000000
0!
0%
b100 *
0-
02
b100 6
#242650000000
1!
1%
1-
12
#242660000000
0!
0%
b101 *
0-
02
b101 6
#242670000000
1!
1%
1-
12
#242680000000
0!
0%
b110 *
0-
02
b110 6
#242690000000
1!
1%
1-
12
#242700000000
0!
0%
b111 *
0-
02
b111 6
#242710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#242720000000
0!
0%
b0 *
0-
02
b0 6
#242730000000
1!
1%
1-
12
#242740000000
0!
0%
b1 *
0-
02
b1 6
#242750000000
1!
1%
1-
12
#242760000000
0!
0%
b10 *
0-
02
b10 6
#242770000000
1!
1%
1-
12
#242780000000
0!
0%
b11 *
0-
02
b11 6
#242790000000
1!
1%
1-
12
15
#242800000000
0!
0%
b100 *
0-
02
b100 6
#242810000000
1!
1%
1-
12
#242820000000
0!
0%
b101 *
0-
02
b101 6
#242830000000
1!
1%
1-
12
#242840000000
0!
0%
b110 *
0-
02
b110 6
#242850000000
1!
1%
1-
12
#242860000000
0!
0%
b111 *
0-
02
b111 6
#242870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#242880000000
0!
0%
b0 *
0-
02
b0 6
#242890000000
1!
1%
1-
12
#242900000000
0!
0%
b1 *
0-
02
b1 6
#242910000000
1!
1%
1-
12
#242920000000
0!
0%
b10 *
0-
02
b10 6
#242930000000
1!
1%
1-
12
#242940000000
0!
0%
b11 *
0-
02
b11 6
#242950000000
1!
1%
1-
12
15
#242960000000
0!
0%
b100 *
0-
02
b100 6
#242970000000
1!
1%
1-
12
#242980000000
0!
0%
b101 *
0-
02
b101 6
#242990000000
1!
1%
1-
12
#243000000000
0!
0%
b110 *
0-
02
b110 6
#243010000000
1!
1%
1-
12
#243020000000
0!
0%
b111 *
0-
02
b111 6
#243030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#243040000000
0!
0%
b0 *
0-
02
b0 6
#243050000000
1!
1%
1-
12
#243060000000
0!
0%
b1 *
0-
02
b1 6
#243070000000
1!
1%
1-
12
#243080000000
0!
0%
b10 *
0-
02
b10 6
#243090000000
1!
1%
1-
12
#243100000000
0!
0%
b11 *
0-
02
b11 6
#243110000000
1!
1%
1-
12
15
#243120000000
0!
0%
b100 *
0-
02
b100 6
#243130000000
1!
1%
1-
12
#243140000000
0!
0%
b101 *
0-
02
b101 6
#243150000000
1!
1%
1-
12
#243160000000
0!
0%
b110 *
0-
02
b110 6
#243170000000
1!
1%
1-
12
#243180000000
0!
0%
b111 *
0-
02
b111 6
#243190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#243200000000
0!
0%
b0 *
0-
02
b0 6
#243210000000
1!
1%
1-
12
#243220000000
0!
0%
b1 *
0-
02
b1 6
#243230000000
1!
1%
1-
12
#243240000000
0!
0%
b10 *
0-
02
b10 6
#243250000000
1!
1%
1-
12
#243260000000
0!
0%
b11 *
0-
02
b11 6
#243270000000
1!
1%
1-
12
15
#243280000000
0!
0%
b100 *
0-
02
b100 6
#243290000000
1!
1%
1-
12
#243300000000
0!
0%
b101 *
0-
02
b101 6
#243310000000
1!
1%
1-
12
#243320000000
0!
0%
b110 *
0-
02
b110 6
#243330000000
1!
1%
1-
12
#243340000000
0!
0%
b111 *
0-
02
b111 6
#243350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#243360000000
0!
0%
b0 *
0-
02
b0 6
#243370000000
1!
1%
1-
12
#243380000000
0!
0%
b1 *
0-
02
b1 6
#243390000000
1!
1%
1-
12
#243400000000
0!
0%
b10 *
0-
02
b10 6
#243410000000
1!
1%
1-
12
#243420000000
0!
0%
b11 *
0-
02
b11 6
#243430000000
1!
1%
1-
12
15
#243440000000
0!
0%
b100 *
0-
02
b100 6
#243450000000
1!
1%
1-
12
#243460000000
0!
0%
b101 *
0-
02
b101 6
#243470000000
1!
1%
1-
12
#243480000000
0!
0%
b110 *
0-
02
b110 6
#243490000000
1!
1%
1-
12
#243500000000
0!
0%
b111 *
0-
02
b111 6
#243510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#243520000000
0!
0%
b0 *
0-
02
b0 6
#243530000000
1!
1%
1-
12
#243540000000
0!
0%
b1 *
0-
02
b1 6
#243550000000
1!
1%
1-
12
#243560000000
0!
0%
b10 *
0-
02
b10 6
#243570000000
1!
1%
1-
12
#243580000000
0!
0%
b11 *
0-
02
b11 6
#243590000000
1!
1%
1-
12
15
#243600000000
0!
0%
b100 *
0-
02
b100 6
#243610000000
1!
1%
1-
12
#243620000000
0!
0%
b101 *
0-
02
b101 6
#243630000000
1!
1%
1-
12
#243640000000
0!
0%
b110 *
0-
02
b110 6
#243650000000
1!
1%
1-
12
#243660000000
0!
0%
b111 *
0-
02
b111 6
#243670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#243680000000
0!
0%
b0 *
0-
02
b0 6
#243690000000
1!
1%
1-
12
#243700000000
0!
0%
b1 *
0-
02
b1 6
#243710000000
1!
1%
1-
12
#243720000000
0!
0%
b10 *
0-
02
b10 6
#243730000000
1!
1%
1-
12
#243740000000
0!
0%
b11 *
0-
02
b11 6
#243750000000
1!
1%
1-
12
15
#243760000000
0!
0%
b100 *
0-
02
b100 6
#243770000000
1!
1%
1-
12
#243780000000
0!
0%
b101 *
0-
02
b101 6
#243790000000
1!
1%
1-
12
#243800000000
0!
0%
b110 *
0-
02
b110 6
#243810000000
1!
1%
1-
12
#243820000000
0!
0%
b111 *
0-
02
b111 6
#243830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#243840000000
0!
0%
b0 *
0-
02
b0 6
#243850000000
1!
1%
1-
12
#243860000000
0!
0%
b1 *
0-
02
b1 6
#243870000000
1!
1%
1-
12
#243880000000
0!
0%
b10 *
0-
02
b10 6
#243890000000
1!
1%
1-
12
#243900000000
0!
0%
b11 *
0-
02
b11 6
#243910000000
1!
1%
1-
12
15
#243920000000
0!
0%
b100 *
0-
02
b100 6
#243930000000
1!
1%
1-
12
#243940000000
0!
0%
b101 *
0-
02
b101 6
#243950000000
1!
1%
1-
12
#243960000000
0!
0%
b110 *
0-
02
b110 6
#243970000000
1!
1%
1-
12
#243980000000
0!
0%
b111 *
0-
02
b111 6
#243990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#244000000000
0!
0%
b0 *
0-
02
b0 6
#244010000000
1!
1%
1-
12
#244020000000
0!
0%
b1 *
0-
02
b1 6
#244030000000
1!
1%
1-
12
#244040000000
0!
0%
b10 *
0-
02
b10 6
#244050000000
1!
1%
1-
12
#244060000000
0!
0%
b11 *
0-
02
b11 6
#244070000000
1!
1%
1-
12
15
#244080000000
0!
0%
b100 *
0-
02
b100 6
#244090000000
1!
1%
1-
12
#244100000000
0!
0%
b101 *
0-
02
b101 6
#244110000000
1!
1%
1-
12
#244120000000
0!
0%
b110 *
0-
02
b110 6
#244130000000
1!
1%
1-
12
#244140000000
0!
0%
b111 *
0-
02
b111 6
#244150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#244160000000
0!
0%
b0 *
0-
02
b0 6
#244170000000
1!
1%
1-
12
#244180000000
0!
0%
b1 *
0-
02
b1 6
#244190000000
1!
1%
1-
12
#244200000000
0!
0%
b10 *
0-
02
b10 6
#244210000000
1!
1%
1-
12
#244220000000
0!
0%
b11 *
0-
02
b11 6
#244230000000
1!
1%
1-
12
15
#244240000000
0!
0%
b100 *
0-
02
b100 6
#244250000000
1!
1%
1-
12
#244260000000
0!
0%
b101 *
0-
02
b101 6
#244270000000
1!
1%
1-
12
#244280000000
0!
0%
b110 *
0-
02
b110 6
#244290000000
1!
1%
1-
12
#244300000000
0!
0%
b111 *
0-
02
b111 6
#244310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#244320000000
0!
0%
b0 *
0-
02
b0 6
#244330000000
1!
1%
1-
12
#244340000000
0!
0%
b1 *
0-
02
b1 6
#244350000000
1!
1%
1-
12
#244360000000
0!
0%
b10 *
0-
02
b10 6
#244370000000
1!
1%
1-
12
#244380000000
0!
0%
b11 *
0-
02
b11 6
#244390000000
1!
1%
1-
12
15
#244400000000
0!
0%
b100 *
0-
02
b100 6
#244410000000
1!
1%
1-
12
#244420000000
0!
0%
b101 *
0-
02
b101 6
#244430000000
1!
1%
1-
12
#244440000000
0!
0%
b110 *
0-
02
b110 6
#244450000000
1!
1%
1-
12
#244460000000
0!
0%
b111 *
0-
02
b111 6
#244470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#244480000000
0!
0%
b0 *
0-
02
b0 6
#244490000000
1!
1%
1-
12
#244500000000
0!
0%
b1 *
0-
02
b1 6
#244510000000
1!
1%
1-
12
#244520000000
0!
0%
b10 *
0-
02
b10 6
#244530000000
1!
1%
1-
12
#244540000000
0!
0%
b11 *
0-
02
b11 6
#244550000000
1!
1%
1-
12
15
#244560000000
0!
0%
b100 *
0-
02
b100 6
#244570000000
1!
1%
1-
12
#244580000000
0!
0%
b101 *
0-
02
b101 6
#244590000000
1!
1%
1-
12
#244600000000
0!
0%
b110 *
0-
02
b110 6
#244610000000
1!
1%
1-
12
#244620000000
0!
0%
b111 *
0-
02
b111 6
#244630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#244640000000
0!
0%
b0 *
0-
02
b0 6
#244650000000
1!
1%
1-
12
#244660000000
0!
0%
b1 *
0-
02
b1 6
#244670000000
1!
1%
1-
12
#244680000000
0!
0%
b10 *
0-
02
b10 6
#244690000000
1!
1%
1-
12
#244700000000
0!
0%
b11 *
0-
02
b11 6
#244710000000
1!
1%
1-
12
15
#244720000000
0!
0%
b100 *
0-
02
b100 6
#244730000000
1!
1%
1-
12
#244740000000
0!
0%
b101 *
0-
02
b101 6
#244750000000
1!
1%
1-
12
#244760000000
0!
0%
b110 *
0-
02
b110 6
#244770000000
1!
1%
1-
12
#244780000000
0!
0%
b111 *
0-
02
b111 6
#244790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#244800000000
0!
0%
b0 *
0-
02
b0 6
#244810000000
1!
1%
1-
12
#244820000000
0!
0%
b1 *
0-
02
b1 6
#244830000000
1!
1%
1-
12
#244840000000
0!
0%
b10 *
0-
02
b10 6
#244850000000
1!
1%
1-
12
#244860000000
0!
0%
b11 *
0-
02
b11 6
#244870000000
1!
1%
1-
12
15
#244880000000
0!
0%
b100 *
0-
02
b100 6
#244890000000
1!
1%
1-
12
#244900000000
0!
0%
b101 *
0-
02
b101 6
#244910000000
1!
1%
1-
12
#244920000000
0!
0%
b110 *
0-
02
b110 6
#244930000000
1!
1%
1-
12
#244940000000
0!
0%
b111 *
0-
02
b111 6
#244950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#244960000000
0!
0%
b0 *
0-
02
b0 6
#244970000000
1!
1%
1-
12
#244980000000
0!
0%
b1 *
0-
02
b1 6
#244990000000
1!
1%
1-
12
#245000000000
0!
0%
b10 *
0-
02
b10 6
#245010000000
1!
1%
1-
12
#245020000000
0!
0%
b11 *
0-
02
b11 6
#245030000000
1!
1%
1-
12
15
#245040000000
0!
0%
b100 *
0-
02
b100 6
#245050000000
1!
1%
1-
12
#245060000000
0!
0%
b101 *
0-
02
b101 6
#245070000000
1!
1%
1-
12
#245080000000
0!
0%
b110 *
0-
02
b110 6
#245090000000
1!
1%
1-
12
#245100000000
0!
0%
b111 *
0-
02
b111 6
#245110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#245120000000
0!
0%
b0 *
0-
02
b0 6
#245130000000
1!
1%
1-
12
#245140000000
0!
0%
b1 *
0-
02
b1 6
#245150000000
1!
1%
1-
12
#245160000000
0!
0%
b10 *
0-
02
b10 6
#245170000000
1!
1%
1-
12
#245180000000
0!
0%
b11 *
0-
02
b11 6
#245190000000
1!
1%
1-
12
15
#245200000000
0!
0%
b100 *
0-
02
b100 6
#245210000000
1!
1%
1-
12
#245220000000
0!
0%
b101 *
0-
02
b101 6
#245230000000
1!
1%
1-
12
#245240000000
0!
0%
b110 *
0-
02
b110 6
#245250000000
1!
1%
1-
12
#245260000000
0!
0%
b111 *
0-
02
b111 6
#245270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#245280000000
0!
0%
b0 *
0-
02
b0 6
#245290000000
1!
1%
1-
12
#245300000000
0!
0%
b1 *
0-
02
b1 6
#245310000000
1!
1%
1-
12
#245320000000
0!
0%
b10 *
0-
02
b10 6
#245330000000
1!
1%
1-
12
#245340000000
0!
0%
b11 *
0-
02
b11 6
#245350000000
1!
1%
1-
12
15
#245360000000
0!
0%
b100 *
0-
02
b100 6
#245370000000
1!
1%
1-
12
#245380000000
0!
0%
b101 *
0-
02
b101 6
#245390000000
1!
1%
1-
12
#245400000000
0!
0%
b110 *
0-
02
b110 6
#245410000000
1!
1%
1-
12
#245420000000
0!
0%
b111 *
0-
02
b111 6
#245430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#245440000000
0!
0%
b0 *
0-
02
b0 6
#245450000000
1!
1%
1-
12
#245460000000
0!
0%
b1 *
0-
02
b1 6
#245470000000
1!
1%
1-
12
#245480000000
0!
0%
b10 *
0-
02
b10 6
#245490000000
1!
1%
1-
12
#245500000000
0!
0%
b11 *
0-
02
b11 6
#245510000000
1!
1%
1-
12
15
#245520000000
0!
0%
b100 *
0-
02
b100 6
#245530000000
1!
1%
1-
12
#245540000000
0!
0%
b101 *
0-
02
b101 6
#245550000000
1!
1%
1-
12
#245560000000
0!
0%
b110 *
0-
02
b110 6
#245570000000
1!
1%
1-
12
#245580000000
0!
0%
b111 *
0-
02
b111 6
#245590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#245600000000
0!
0%
b0 *
0-
02
b0 6
#245610000000
1!
1%
1-
12
#245620000000
0!
0%
b1 *
0-
02
b1 6
#245630000000
1!
1%
1-
12
#245640000000
0!
0%
b10 *
0-
02
b10 6
#245650000000
1!
1%
1-
12
#245660000000
0!
0%
b11 *
0-
02
b11 6
#245670000000
1!
1%
1-
12
15
#245680000000
0!
0%
b100 *
0-
02
b100 6
#245690000000
1!
1%
1-
12
#245700000000
0!
0%
b101 *
0-
02
b101 6
#245710000000
1!
1%
1-
12
#245720000000
0!
0%
b110 *
0-
02
b110 6
#245730000000
1!
1%
1-
12
#245740000000
0!
0%
b111 *
0-
02
b111 6
#245750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#245760000000
0!
0%
b0 *
0-
02
b0 6
#245770000000
1!
1%
1-
12
#245780000000
0!
0%
b1 *
0-
02
b1 6
#245790000000
1!
1%
1-
12
#245800000000
0!
0%
b10 *
0-
02
b10 6
#245810000000
1!
1%
1-
12
#245820000000
0!
0%
b11 *
0-
02
b11 6
#245830000000
1!
1%
1-
12
15
#245840000000
0!
0%
b100 *
0-
02
b100 6
#245850000000
1!
1%
1-
12
#245860000000
0!
0%
b101 *
0-
02
b101 6
#245870000000
1!
1%
1-
12
#245880000000
0!
0%
b110 *
0-
02
b110 6
#245890000000
1!
1%
1-
12
#245900000000
0!
0%
b111 *
0-
02
b111 6
#245910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#245920000000
0!
0%
b0 *
0-
02
b0 6
#245930000000
1!
1%
1-
12
#245940000000
0!
0%
b1 *
0-
02
b1 6
#245950000000
1!
1%
1-
12
#245960000000
0!
0%
b10 *
0-
02
b10 6
#245970000000
1!
1%
1-
12
#245980000000
0!
0%
b11 *
0-
02
b11 6
#245990000000
1!
1%
1-
12
15
#246000000000
0!
0%
b100 *
0-
02
b100 6
#246010000000
1!
1%
1-
12
#246020000000
0!
0%
b101 *
0-
02
b101 6
#246030000000
1!
1%
1-
12
#246040000000
0!
0%
b110 *
0-
02
b110 6
#246050000000
1!
1%
1-
12
#246060000000
0!
0%
b111 *
0-
02
b111 6
#246070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#246080000000
0!
0%
b0 *
0-
02
b0 6
#246090000000
1!
1%
1-
12
#246100000000
0!
0%
b1 *
0-
02
b1 6
#246110000000
1!
1%
1-
12
#246120000000
0!
0%
b10 *
0-
02
b10 6
#246130000000
1!
1%
1-
12
#246140000000
0!
0%
b11 *
0-
02
b11 6
#246150000000
1!
1%
1-
12
15
#246160000000
0!
0%
b100 *
0-
02
b100 6
#246170000000
1!
1%
1-
12
#246180000000
0!
0%
b101 *
0-
02
b101 6
#246190000000
1!
1%
1-
12
#246200000000
0!
0%
b110 *
0-
02
b110 6
#246210000000
1!
1%
1-
12
#246220000000
0!
0%
b111 *
0-
02
b111 6
#246230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#246240000000
0!
0%
b0 *
0-
02
b0 6
#246250000000
1!
1%
1-
12
#246260000000
0!
0%
b1 *
0-
02
b1 6
#246270000000
1!
1%
1-
12
#246280000000
0!
0%
b10 *
0-
02
b10 6
#246290000000
1!
1%
1-
12
#246300000000
0!
0%
b11 *
0-
02
b11 6
#246310000000
1!
1%
1-
12
15
#246320000000
0!
0%
b100 *
0-
02
b100 6
#246330000000
1!
1%
1-
12
#246340000000
0!
0%
b101 *
0-
02
b101 6
#246350000000
1!
1%
1-
12
#246360000000
0!
0%
b110 *
0-
02
b110 6
#246370000000
1!
1%
1-
12
#246380000000
0!
0%
b111 *
0-
02
b111 6
#246390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#246400000000
0!
0%
b0 *
0-
02
b0 6
#246410000000
1!
1%
1-
12
#246420000000
0!
0%
b1 *
0-
02
b1 6
#246430000000
1!
1%
1-
12
#246440000000
0!
0%
b10 *
0-
02
b10 6
#246450000000
1!
1%
1-
12
#246460000000
0!
0%
b11 *
0-
02
b11 6
#246470000000
1!
1%
1-
12
15
#246480000000
0!
0%
b100 *
0-
02
b100 6
#246490000000
1!
1%
1-
12
#246500000000
0!
0%
b101 *
0-
02
b101 6
#246510000000
1!
1%
1-
12
#246520000000
0!
0%
b110 *
0-
02
b110 6
#246530000000
1!
1%
1-
12
#246540000000
0!
0%
b111 *
0-
02
b111 6
#246550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#246560000000
0!
0%
b0 *
0-
02
b0 6
#246570000000
1!
1%
1-
12
#246580000000
0!
0%
b1 *
0-
02
b1 6
#246590000000
1!
1%
1-
12
#246600000000
0!
0%
b10 *
0-
02
b10 6
#246610000000
1!
1%
1-
12
#246620000000
0!
0%
b11 *
0-
02
b11 6
#246630000000
1!
1%
1-
12
15
#246640000000
0!
0%
b100 *
0-
02
b100 6
#246650000000
1!
1%
1-
12
#246660000000
0!
0%
b101 *
0-
02
b101 6
#246670000000
1!
1%
1-
12
#246680000000
0!
0%
b110 *
0-
02
b110 6
#246690000000
1!
1%
1-
12
#246700000000
0!
0%
b111 *
0-
02
b111 6
#246710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#246720000000
0!
0%
b0 *
0-
02
b0 6
#246730000000
1!
1%
1-
12
#246740000000
0!
0%
b1 *
0-
02
b1 6
#246750000000
1!
1%
1-
12
#246760000000
0!
0%
b10 *
0-
02
b10 6
#246770000000
1!
1%
1-
12
#246780000000
0!
0%
b11 *
0-
02
b11 6
#246790000000
1!
1%
1-
12
15
#246800000000
0!
0%
b100 *
0-
02
b100 6
#246810000000
1!
1%
1-
12
#246820000000
0!
0%
b101 *
0-
02
b101 6
#246830000000
1!
1%
1-
12
#246840000000
0!
0%
b110 *
0-
02
b110 6
#246850000000
1!
1%
1-
12
#246860000000
0!
0%
b111 *
0-
02
b111 6
#246870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#246880000000
0!
0%
b0 *
0-
02
b0 6
#246890000000
1!
1%
1-
12
#246900000000
0!
0%
b1 *
0-
02
b1 6
#246910000000
1!
1%
1-
12
#246920000000
0!
0%
b10 *
0-
02
b10 6
#246930000000
1!
1%
1-
12
#246940000000
0!
0%
b11 *
0-
02
b11 6
#246950000000
1!
1%
1-
12
15
#246960000000
0!
0%
b100 *
0-
02
b100 6
#246970000000
1!
1%
1-
12
#246980000000
0!
0%
b101 *
0-
02
b101 6
#246990000000
1!
1%
1-
12
#247000000000
0!
0%
b110 *
0-
02
b110 6
#247010000000
1!
1%
1-
12
#247020000000
0!
0%
b111 *
0-
02
b111 6
#247030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#247040000000
0!
0%
b0 *
0-
02
b0 6
#247050000000
1!
1%
1-
12
#247060000000
0!
0%
b1 *
0-
02
b1 6
#247070000000
1!
1%
1-
12
#247080000000
0!
0%
b10 *
0-
02
b10 6
#247090000000
1!
1%
1-
12
#247100000000
0!
0%
b11 *
0-
02
b11 6
#247110000000
1!
1%
1-
12
15
#247120000000
0!
0%
b100 *
0-
02
b100 6
#247130000000
1!
1%
1-
12
#247140000000
0!
0%
b101 *
0-
02
b101 6
#247150000000
1!
1%
1-
12
#247160000000
0!
0%
b110 *
0-
02
b110 6
#247170000000
1!
1%
1-
12
#247180000000
0!
0%
b111 *
0-
02
b111 6
#247190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#247200000000
0!
0%
b0 *
0-
02
b0 6
#247210000000
1!
1%
1-
12
#247220000000
0!
0%
b1 *
0-
02
b1 6
#247230000000
1!
1%
1-
12
#247240000000
0!
0%
b10 *
0-
02
b10 6
#247250000000
1!
1%
1-
12
#247260000000
0!
0%
b11 *
0-
02
b11 6
#247270000000
1!
1%
1-
12
15
#247280000000
0!
0%
b100 *
0-
02
b100 6
#247290000000
1!
1%
1-
12
#247300000000
0!
0%
b101 *
0-
02
b101 6
#247310000000
1!
1%
1-
12
#247320000000
0!
0%
b110 *
0-
02
b110 6
#247330000000
1!
1%
1-
12
#247340000000
0!
0%
b111 *
0-
02
b111 6
#247350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#247360000000
0!
0%
b0 *
0-
02
b0 6
#247370000000
1!
1%
1-
12
#247380000000
0!
0%
b1 *
0-
02
b1 6
#247390000000
1!
1%
1-
12
#247400000000
0!
0%
b10 *
0-
02
b10 6
#247410000000
1!
1%
1-
12
#247420000000
0!
0%
b11 *
0-
02
b11 6
#247430000000
1!
1%
1-
12
15
#247440000000
0!
0%
b100 *
0-
02
b100 6
#247450000000
1!
1%
1-
12
#247460000000
0!
0%
b101 *
0-
02
b101 6
#247470000000
1!
1%
1-
12
#247480000000
0!
0%
b110 *
0-
02
b110 6
#247490000000
1!
1%
1-
12
#247500000000
0!
0%
b111 *
0-
02
b111 6
#247510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#247520000000
0!
0%
b0 *
0-
02
b0 6
#247530000000
1!
1%
1-
12
#247540000000
0!
0%
b1 *
0-
02
b1 6
#247550000000
1!
1%
1-
12
#247560000000
0!
0%
b10 *
0-
02
b10 6
#247570000000
1!
1%
1-
12
#247580000000
0!
0%
b11 *
0-
02
b11 6
#247590000000
1!
1%
1-
12
15
#247600000000
0!
0%
b100 *
0-
02
b100 6
#247610000000
1!
1%
1-
12
#247620000000
0!
0%
b101 *
0-
02
b101 6
#247630000000
1!
1%
1-
12
#247640000000
0!
0%
b110 *
0-
02
b110 6
#247650000000
1!
1%
1-
12
#247660000000
0!
0%
b111 *
0-
02
b111 6
#247670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#247680000000
0!
0%
b0 *
0-
02
b0 6
#247690000000
1!
1%
1-
12
#247700000000
0!
0%
b1 *
0-
02
b1 6
#247710000000
1!
1%
1-
12
#247720000000
0!
0%
b10 *
0-
02
b10 6
#247730000000
1!
1%
1-
12
#247740000000
0!
0%
b11 *
0-
02
b11 6
#247750000000
1!
1%
1-
12
15
#247760000000
0!
0%
b100 *
0-
02
b100 6
#247770000000
1!
1%
1-
12
#247780000000
0!
0%
b101 *
0-
02
b101 6
#247790000000
1!
1%
1-
12
#247800000000
0!
0%
b110 *
0-
02
b110 6
#247810000000
1!
1%
1-
12
#247820000000
0!
0%
b111 *
0-
02
b111 6
#247830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#247840000000
0!
0%
b0 *
0-
02
b0 6
#247850000000
1!
1%
1-
12
#247860000000
0!
0%
b1 *
0-
02
b1 6
#247870000000
1!
1%
1-
12
#247880000000
0!
0%
b10 *
0-
02
b10 6
#247890000000
1!
1%
1-
12
#247900000000
0!
0%
b11 *
0-
02
b11 6
#247910000000
1!
1%
1-
12
15
#247920000000
0!
0%
b100 *
0-
02
b100 6
#247930000000
1!
1%
1-
12
#247940000000
0!
0%
b101 *
0-
02
b101 6
#247950000000
1!
1%
1-
12
#247960000000
0!
0%
b110 *
0-
02
b110 6
#247970000000
1!
1%
1-
12
#247980000000
0!
0%
b111 *
0-
02
b111 6
#247990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#248000000000
0!
0%
b0 *
0-
02
b0 6
#248010000000
1!
1%
1-
12
#248020000000
0!
0%
b1 *
0-
02
b1 6
#248030000000
1!
1%
1-
12
#248040000000
0!
0%
b10 *
0-
02
b10 6
#248050000000
1!
1%
1-
12
#248060000000
0!
0%
b11 *
0-
02
b11 6
#248070000000
1!
1%
1-
12
15
#248080000000
0!
0%
b100 *
0-
02
b100 6
#248090000000
1!
1%
1-
12
#248100000000
0!
0%
b101 *
0-
02
b101 6
#248110000000
1!
1%
1-
12
#248120000000
0!
0%
b110 *
0-
02
b110 6
#248130000000
1!
1%
1-
12
#248140000000
0!
0%
b111 *
0-
02
b111 6
#248150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#248160000000
0!
0%
b0 *
0-
02
b0 6
#248170000000
1!
1%
1-
12
#248180000000
0!
0%
b1 *
0-
02
b1 6
#248190000000
1!
1%
1-
12
#248200000000
0!
0%
b10 *
0-
02
b10 6
#248210000000
1!
1%
1-
12
#248220000000
0!
0%
b11 *
0-
02
b11 6
#248230000000
1!
1%
1-
12
15
#248240000000
0!
0%
b100 *
0-
02
b100 6
#248250000000
1!
1%
1-
12
#248260000000
0!
0%
b101 *
0-
02
b101 6
#248270000000
1!
1%
1-
12
#248280000000
0!
0%
b110 *
0-
02
b110 6
#248290000000
1!
1%
1-
12
#248300000000
0!
0%
b111 *
0-
02
b111 6
#248310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#248320000000
0!
0%
b0 *
0-
02
b0 6
#248330000000
1!
1%
1-
12
#248340000000
0!
0%
b1 *
0-
02
b1 6
#248350000000
1!
1%
1-
12
#248360000000
0!
0%
b10 *
0-
02
b10 6
#248370000000
1!
1%
1-
12
#248380000000
0!
0%
b11 *
0-
02
b11 6
#248390000000
1!
1%
1-
12
15
#248400000000
0!
0%
b100 *
0-
02
b100 6
#248410000000
1!
1%
1-
12
#248420000000
0!
0%
b101 *
0-
02
b101 6
#248430000000
1!
1%
1-
12
#248440000000
0!
0%
b110 *
0-
02
b110 6
#248450000000
1!
1%
1-
12
#248460000000
0!
0%
b111 *
0-
02
b111 6
#248470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#248480000000
0!
0%
b0 *
0-
02
b0 6
#248490000000
1!
1%
1-
12
#248500000000
0!
0%
b1 *
0-
02
b1 6
#248510000000
1!
1%
1-
12
#248520000000
0!
0%
b10 *
0-
02
b10 6
#248530000000
1!
1%
1-
12
#248540000000
0!
0%
b11 *
0-
02
b11 6
#248550000000
1!
1%
1-
12
15
#248560000000
0!
0%
b100 *
0-
02
b100 6
#248570000000
1!
1%
1-
12
#248580000000
0!
0%
b101 *
0-
02
b101 6
#248590000000
1!
1%
1-
12
#248600000000
0!
0%
b110 *
0-
02
b110 6
#248610000000
1!
1%
1-
12
#248620000000
0!
0%
b111 *
0-
02
b111 6
#248630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#248640000000
0!
0%
b0 *
0-
02
b0 6
#248650000000
1!
1%
1-
12
#248660000000
0!
0%
b1 *
0-
02
b1 6
#248670000000
1!
1%
1-
12
#248680000000
0!
0%
b10 *
0-
02
b10 6
#248690000000
1!
1%
1-
12
#248700000000
0!
0%
b11 *
0-
02
b11 6
#248710000000
1!
1%
1-
12
15
#248720000000
0!
0%
b100 *
0-
02
b100 6
#248730000000
1!
1%
1-
12
#248740000000
0!
0%
b101 *
0-
02
b101 6
#248750000000
1!
1%
1-
12
#248760000000
0!
0%
b110 *
0-
02
b110 6
#248770000000
1!
1%
1-
12
#248780000000
0!
0%
b111 *
0-
02
b111 6
#248790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#248800000000
0!
0%
b0 *
0-
02
b0 6
#248810000000
1!
1%
1-
12
#248820000000
0!
0%
b1 *
0-
02
b1 6
#248830000000
1!
1%
1-
12
#248840000000
0!
0%
b10 *
0-
02
b10 6
#248850000000
1!
1%
1-
12
#248860000000
0!
0%
b11 *
0-
02
b11 6
#248870000000
1!
1%
1-
12
15
#248880000000
0!
0%
b100 *
0-
02
b100 6
#248890000000
1!
1%
1-
12
#248900000000
0!
0%
b101 *
0-
02
b101 6
#248910000000
1!
1%
1-
12
#248920000000
0!
0%
b110 *
0-
02
b110 6
#248930000000
1!
1%
1-
12
#248940000000
0!
0%
b111 *
0-
02
b111 6
#248950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#248960000000
0!
0%
b0 *
0-
02
b0 6
#248970000000
1!
1%
1-
12
#248980000000
0!
0%
b1 *
0-
02
b1 6
#248990000000
1!
1%
1-
12
#249000000000
0!
0%
b10 *
0-
02
b10 6
#249010000000
1!
1%
1-
12
#249020000000
0!
0%
b11 *
0-
02
b11 6
#249030000000
1!
1%
1-
12
15
#249040000000
0!
0%
b100 *
0-
02
b100 6
#249050000000
1!
1%
1-
12
#249060000000
0!
0%
b101 *
0-
02
b101 6
#249070000000
1!
1%
1-
12
#249080000000
0!
0%
b110 *
0-
02
b110 6
#249090000000
1!
1%
1-
12
#249100000000
0!
0%
b111 *
0-
02
b111 6
#249110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#249120000000
0!
0%
b0 *
0-
02
b0 6
#249130000000
1!
1%
1-
12
#249140000000
0!
0%
b1 *
0-
02
b1 6
#249150000000
1!
1%
1-
12
#249160000000
0!
0%
b10 *
0-
02
b10 6
#249170000000
1!
1%
1-
12
#249180000000
0!
0%
b11 *
0-
02
b11 6
#249190000000
1!
1%
1-
12
15
#249200000000
0!
0%
b100 *
0-
02
b100 6
#249210000000
1!
1%
1-
12
#249220000000
0!
0%
b101 *
0-
02
b101 6
#249230000000
1!
1%
1-
12
#249240000000
0!
0%
b110 *
0-
02
b110 6
#249250000000
1!
1%
1-
12
#249260000000
0!
0%
b111 *
0-
02
b111 6
#249270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#249280000000
0!
0%
b0 *
0-
02
b0 6
#249290000000
1!
1%
1-
12
#249300000000
0!
0%
b1 *
0-
02
b1 6
#249310000000
1!
1%
1-
12
#249320000000
0!
0%
b10 *
0-
02
b10 6
#249330000000
1!
1%
1-
12
#249340000000
0!
0%
b11 *
0-
02
b11 6
#249350000000
1!
1%
1-
12
15
#249360000000
0!
0%
b100 *
0-
02
b100 6
#249370000000
1!
1%
1-
12
#249380000000
0!
0%
b101 *
0-
02
b101 6
#249390000000
1!
1%
1-
12
#249400000000
0!
0%
b110 *
0-
02
b110 6
#249410000000
1!
1%
1-
12
#249420000000
0!
0%
b111 *
0-
02
b111 6
#249430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#249440000000
0!
0%
b0 *
0-
02
b0 6
#249450000000
1!
1%
1-
12
#249460000000
0!
0%
b1 *
0-
02
b1 6
#249470000000
1!
1%
1-
12
#249480000000
0!
0%
b10 *
0-
02
b10 6
#249490000000
1!
1%
1-
12
#249500000000
0!
0%
b11 *
0-
02
b11 6
#249510000000
1!
1%
1-
12
15
#249520000000
0!
0%
b100 *
0-
02
b100 6
#249530000000
1!
1%
1-
12
#249540000000
0!
0%
b101 *
0-
02
b101 6
#249550000000
1!
1%
1-
12
#249560000000
0!
0%
b110 *
0-
02
b110 6
#249570000000
1!
1%
1-
12
#249580000000
0!
0%
b111 *
0-
02
b111 6
#249590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#249600000000
0!
0%
b0 *
0-
02
b0 6
#249610000000
1!
1%
1-
12
#249620000000
0!
0%
b1 *
0-
02
b1 6
#249630000000
1!
1%
1-
12
#249640000000
0!
0%
b10 *
0-
02
b10 6
#249650000000
1!
1%
1-
12
#249660000000
0!
0%
b11 *
0-
02
b11 6
#249670000000
1!
1%
1-
12
15
#249680000000
0!
0%
b100 *
0-
02
b100 6
#249690000000
1!
1%
1-
12
#249700000000
0!
0%
b101 *
0-
02
b101 6
#249710000000
1!
1%
1-
12
#249720000000
0!
0%
b110 *
0-
02
b110 6
#249730000000
1!
1%
1-
12
#249740000000
0!
0%
b111 *
0-
02
b111 6
#249750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#249760000000
0!
0%
b0 *
0-
02
b0 6
#249770000000
1!
1%
1-
12
#249780000000
0!
0%
b1 *
0-
02
b1 6
#249790000000
1!
1%
1-
12
#249800000000
0!
0%
b10 *
0-
02
b10 6
#249810000000
1!
1%
1-
12
#249820000000
0!
0%
b11 *
0-
02
b11 6
#249830000000
1!
1%
1-
12
15
#249840000000
0!
0%
b100 *
0-
02
b100 6
#249850000000
1!
1%
1-
12
#249860000000
0!
0%
b101 *
0-
02
b101 6
#249870000000
1!
1%
1-
12
#249880000000
0!
0%
b110 *
0-
02
b110 6
#249890000000
1!
1%
1-
12
#249900000000
0!
0%
b111 *
0-
02
b111 6
#249910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#249920000000
0!
0%
b0 *
0-
02
b0 6
#249930000000
1!
1%
1-
12
#249940000000
0!
0%
b1 *
0-
02
b1 6
#249950000000
1!
1%
1-
12
#249960000000
0!
0%
b10 *
0-
02
b10 6
#249970000000
1!
1%
1-
12
#249980000000
0!
0%
b11 *
0-
02
b11 6
#249990000000
1!
1%
1-
12
15
#250000000000
0!
0%
b100 *
0-
02
b100 6
#250010000000
1!
1%
1-
12
#250020000000
0!
0%
b101 *
0-
02
b101 6
#250030000000
1!
1%
1-
12
#250040000000
0!
0%
b110 *
0-
02
b110 6
#250050000000
1!
1%
1-
12
#250060000000
0!
0%
b111 *
0-
02
b111 6
#250070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#250080000000
0!
0%
b0 *
0-
02
b0 6
#250090000000
1!
1%
1-
12
#250100000000
0!
0%
b1 *
0-
02
b1 6
#250110000000
1!
1%
1-
12
#250120000000
0!
0%
b10 *
0-
02
b10 6
#250130000000
1!
1%
1-
12
#250140000000
0!
0%
b11 *
0-
02
b11 6
#250150000000
1!
1%
1-
12
15
#250160000000
0!
0%
b100 *
0-
02
b100 6
#250170000000
1!
1%
1-
12
#250180000000
0!
0%
b101 *
0-
02
b101 6
#250190000000
1!
1%
1-
12
#250200000000
0!
0%
b110 *
0-
02
b110 6
#250210000000
1!
1%
1-
12
#250220000000
0!
0%
b111 *
0-
02
b111 6
#250230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#250240000000
0!
0%
b0 *
0-
02
b0 6
#250250000000
1!
1%
1-
12
#250260000000
0!
0%
b1 *
0-
02
b1 6
#250270000000
1!
1%
1-
12
#250280000000
0!
0%
b10 *
0-
02
b10 6
#250290000000
1!
1%
1-
12
#250300000000
0!
0%
b11 *
0-
02
b11 6
#250310000000
1!
1%
1-
12
15
#250320000000
0!
0%
b100 *
0-
02
b100 6
#250330000000
1!
1%
1-
12
#250340000000
0!
0%
b101 *
0-
02
b101 6
#250350000000
1!
1%
1-
12
#250360000000
0!
0%
b110 *
0-
02
b110 6
#250370000000
1!
1%
1-
12
#250380000000
0!
0%
b111 *
0-
02
b111 6
#250390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#250400000000
0!
0%
b0 *
0-
02
b0 6
#250410000000
1!
1%
1-
12
#250420000000
0!
0%
b1 *
0-
02
b1 6
#250430000000
1!
1%
1-
12
#250440000000
0!
0%
b10 *
0-
02
b10 6
#250450000000
1!
1%
1-
12
#250460000000
0!
0%
b11 *
0-
02
b11 6
#250470000000
1!
1%
1-
12
15
#250480000000
0!
0%
b100 *
0-
02
b100 6
#250490000000
1!
1%
1-
12
#250500000000
0!
0%
b101 *
0-
02
b101 6
#250510000000
1!
1%
1-
12
#250520000000
0!
0%
b110 *
0-
02
b110 6
#250530000000
1!
1%
1-
12
#250540000000
0!
0%
b111 *
0-
02
b111 6
#250550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#250560000000
0!
0%
b0 *
0-
02
b0 6
#250570000000
1!
1%
1-
12
#250580000000
0!
0%
b1 *
0-
02
b1 6
#250590000000
1!
1%
1-
12
#250600000000
0!
0%
b10 *
0-
02
b10 6
#250610000000
1!
1%
1-
12
#250620000000
0!
0%
b11 *
0-
02
b11 6
#250630000000
1!
1%
1-
12
15
#250640000000
0!
0%
b100 *
0-
02
b100 6
#250650000000
1!
1%
1-
12
#250660000000
0!
0%
b101 *
0-
02
b101 6
#250670000000
1!
1%
1-
12
#250680000000
0!
0%
b110 *
0-
02
b110 6
#250690000000
1!
1%
1-
12
#250700000000
0!
0%
b111 *
0-
02
b111 6
#250710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#250720000000
0!
0%
b0 *
0-
02
b0 6
#250730000000
1!
1%
1-
12
#250740000000
0!
0%
b1 *
0-
02
b1 6
#250750000000
1!
1%
1-
12
#250760000000
0!
0%
b10 *
0-
02
b10 6
#250770000000
1!
1%
1-
12
#250780000000
0!
0%
b11 *
0-
02
b11 6
#250790000000
1!
1%
1-
12
15
#250800000000
0!
0%
b100 *
0-
02
b100 6
#250810000000
1!
1%
1-
12
#250820000000
0!
0%
b101 *
0-
02
b101 6
#250830000000
1!
1%
1-
12
#250840000000
0!
0%
b110 *
0-
02
b110 6
#250850000000
1!
1%
1-
12
#250860000000
0!
0%
b111 *
0-
02
b111 6
#250870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#250880000000
0!
0%
b0 *
0-
02
b0 6
#250890000000
1!
1%
1-
12
#250900000000
0!
0%
b1 *
0-
02
b1 6
#250910000000
1!
1%
1-
12
#250920000000
0!
0%
b10 *
0-
02
b10 6
#250930000000
1!
1%
1-
12
#250940000000
0!
0%
b11 *
0-
02
b11 6
#250950000000
1!
1%
1-
12
15
#250960000000
0!
0%
b100 *
0-
02
b100 6
#250970000000
1!
1%
1-
12
#250980000000
0!
0%
b101 *
0-
02
b101 6
#250990000000
1!
1%
1-
12
#251000000000
0!
0%
b110 *
0-
02
b110 6
#251010000000
1!
1%
1-
12
#251020000000
0!
0%
b111 *
0-
02
b111 6
#251030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#251040000000
0!
0%
b0 *
0-
02
b0 6
#251050000000
1!
1%
1-
12
#251060000000
0!
0%
b1 *
0-
02
b1 6
#251070000000
1!
1%
1-
12
#251080000000
0!
0%
b10 *
0-
02
b10 6
#251090000000
1!
1%
1-
12
#251100000000
0!
0%
b11 *
0-
02
b11 6
#251110000000
1!
1%
1-
12
15
#251120000000
0!
0%
b100 *
0-
02
b100 6
#251130000000
1!
1%
1-
12
#251140000000
0!
0%
b101 *
0-
02
b101 6
#251150000000
1!
1%
1-
12
#251160000000
0!
0%
b110 *
0-
02
b110 6
#251170000000
1!
1%
1-
12
#251180000000
0!
0%
b111 *
0-
02
b111 6
#251190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#251200000000
0!
0%
b0 *
0-
02
b0 6
#251210000000
1!
1%
1-
12
#251220000000
0!
0%
b1 *
0-
02
b1 6
#251230000000
1!
1%
1-
12
#251240000000
0!
0%
b10 *
0-
02
b10 6
#251250000000
1!
1%
1-
12
#251260000000
0!
0%
b11 *
0-
02
b11 6
#251270000000
1!
1%
1-
12
15
#251280000000
0!
0%
b100 *
0-
02
b100 6
#251290000000
1!
1%
1-
12
#251300000000
0!
0%
b101 *
0-
02
b101 6
#251310000000
1!
1%
1-
12
#251320000000
0!
0%
b110 *
0-
02
b110 6
#251330000000
1!
1%
1-
12
#251340000000
0!
0%
b111 *
0-
02
b111 6
#251350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#251360000000
0!
0%
b0 *
0-
02
b0 6
#251370000000
1!
1%
1-
12
#251380000000
0!
0%
b1 *
0-
02
b1 6
#251390000000
1!
1%
1-
12
#251400000000
0!
0%
b10 *
0-
02
b10 6
#251410000000
1!
1%
1-
12
#251420000000
0!
0%
b11 *
0-
02
b11 6
#251430000000
1!
1%
1-
12
15
#251440000000
0!
0%
b100 *
0-
02
b100 6
#251450000000
1!
1%
1-
12
#251460000000
0!
0%
b101 *
0-
02
b101 6
#251470000000
1!
1%
1-
12
#251480000000
0!
0%
b110 *
0-
02
b110 6
#251490000000
1!
1%
1-
12
#251500000000
0!
0%
b111 *
0-
02
b111 6
#251510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#251520000000
0!
0%
b0 *
0-
02
b0 6
#251530000000
1!
1%
1-
12
#251540000000
0!
0%
b1 *
0-
02
b1 6
#251550000000
1!
1%
1-
12
#251560000000
0!
0%
b10 *
0-
02
b10 6
#251570000000
1!
1%
1-
12
#251580000000
0!
0%
b11 *
0-
02
b11 6
#251590000000
1!
1%
1-
12
15
#251600000000
0!
0%
b100 *
0-
02
b100 6
#251610000000
1!
1%
1-
12
#251620000000
0!
0%
b101 *
0-
02
b101 6
#251630000000
1!
1%
1-
12
#251640000000
0!
0%
b110 *
0-
02
b110 6
#251650000000
1!
1%
1-
12
#251660000000
0!
0%
b111 *
0-
02
b111 6
#251670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#251680000000
0!
0%
b0 *
0-
02
b0 6
#251690000000
1!
1%
1-
12
#251700000000
0!
0%
b1 *
0-
02
b1 6
#251710000000
1!
1%
1-
12
#251720000000
0!
0%
b10 *
0-
02
b10 6
#251730000000
1!
1%
1-
12
#251740000000
0!
0%
b11 *
0-
02
b11 6
#251750000000
1!
1%
1-
12
15
#251760000000
0!
0%
b100 *
0-
02
b100 6
#251770000000
1!
1%
1-
12
#251780000000
0!
0%
b101 *
0-
02
b101 6
#251790000000
1!
1%
1-
12
#251800000000
0!
0%
b110 *
0-
02
b110 6
#251810000000
1!
1%
1-
12
#251820000000
0!
0%
b111 *
0-
02
b111 6
#251830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#251840000000
0!
0%
b0 *
0-
02
b0 6
#251850000000
1!
1%
1-
12
#251860000000
0!
0%
b1 *
0-
02
b1 6
#251870000000
1!
1%
1-
12
#251880000000
0!
0%
b10 *
0-
02
b10 6
#251890000000
1!
1%
1-
12
#251900000000
0!
0%
b11 *
0-
02
b11 6
#251910000000
1!
1%
1-
12
15
#251920000000
0!
0%
b100 *
0-
02
b100 6
#251930000000
1!
1%
1-
12
#251940000000
0!
0%
b101 *
0-
02
b101 6
#251950000000
1!
1%
1-
12
#251960000000
0!
0%
b110 *
0-
02
b110 6
#251970000000
1!
1%
1-
12
#251980000000
0!
0%
b111 *
0-
02
b111 6
#251990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#252000000000
0!
0%
b0 *
0-
02
b0 6
#252010000000
1!
1%
1-
12
#252020000000
0!
0%
b1 *
0-
02
b1 6
#252030000000
1!
1%
1-
12
#252040000000
0!
0%
b10 *
0-
02
b10 6
#252050000000
1!
1%
1-
12
#252060000000
0!
0%
b11 *
0-
02
b11 6
#252070000000
1!
1%
1-
12
15
#252080000000
0!
0%
b100 *
0-
02
b100 6
#252090000000
1!
1%
1-
12
#252100000000
0!
0%
b101 *
0-
02
b101 6
#252110000000
1!
1%
1-
12
#252120000000
0!
0%
b110 *
0-
02
b110 6
#252130000000
1!
1%
1-
12
#252140000000
0!
0%
b111 *
0-
02
b111 6
#252150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#252160000000
0!
0%
b0 *
0-
02
b0 6
#252170000000
1!
1%
1-
12
#252180000000
0!
0%
b1 *
0-
02
b1 6
#252190000000
1!
1%
1-
12
#252200000000
0!
0%
b10 *
0-
02
b10 6
#252210000000
1!
1%
1-
12
#252220000000
0!
0%
b11 *
0-
02
b11 6
#252230000000
1!
1%
1-
12
15
#252240000000
0!
0%
b100 *
0-
02
b100 6
#252250000000
1!
1%
1-
12
#252260000000
0!
0%
b101 *
0-
02
b101 6
#252270000000
1!
1%
1-
12
#252280000000
0!
0%
b110 *
0-
02
b110 6
#252290000000
1!
1%
1-
12
#252300000000
0!
0%
b111 *
0-
02
b111 6
#252310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#252320000000
0!
0%
b0 *
0-
02
b0 6
#252330000000
1!
1%
1-
12
#252340000000
0!
0%
b1 *
0-
02
b1 6
#252350000000
1!
1%
1-
12
#252360000000
0!
0%
b10 *
0-
02
b10 6
#252370000000
1!
1%
1-
12
#252380000000
0!
0%
b11 *
0-
02
b11 6
#252390000000
1!
1%
1-
12
15
#252400000000
0!
0%
b100 *
0-
02
b100 6
#252410000000
1!
1%
1-
12
#252420000000
0!
0%
b101 *
0-
02
b101 6
#252430000000
1!
1%
1-
12
#252440000000
0!
0%
b110 *
0-
02
b110 6
#252450000000
1!
1%
1-
12
#252460000000
0!
0%
b111 *
0-
02
b111 6
#252470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#252480000000
0!
0%
b0 *
0-
02
b0 6
#252490000000
1!
1%
1-
12
#252500000000
0!
0%
b1 *
0-
02
b1 6
#252510000000
1!
1%
1-
12
#252520000000
0!
0%
b10 *
0-
02
b10 6
#252530000000
1!
1%
1-
12
#252540000000
0!
0%
b11 *
0-
02
b11 6
#252550000000
1!
1%
1-
12
15
#252560000000
0!
0%
b100 *
0-
02
b100 6
#252570000000
1!
1%
1-
12
#252580000000
0!
0%
b101 *
0-
02
b101 6
#252590000000
1!
1%
1-
12
#252600000000
0!
0%
b110 *
0-
02
b110 6
#252610000000
1!
1%
1-
12
#252620000000
0!
0%
b111 *
0-
02
b111 6
#252630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#252640000000
0!
0%
b0 *
0-
02
b0 6
#252650000000
1!
1%
1-
12
#252660000000
0!
0%
b1 *
0-
02
b1 6
#252670000000
1!
1%
1-
12
#252680000000
0!
0%
b10 *
0-
02
b10 6
#252690000000
1!
1%
1-
12
#252700000000
0!
0%
b11 *
0-
02
b11 6
#252710000000
1!
1%
1-
12
15
#252720000000
0!
0%
b100 *
0-
02
b100 6
#252730000000
1!
1%
1-
12
#252740000000
0!
0%
b101 *
0-
02
b101 6
#252750000000
1!
1%
1-
12
#252760000000
0!
0%
b110 *
0-
02
b110 6
#252770000000
1!
1%
1-
12
#252780000000
0!
0%
b111 *
0-
02
b111 6
#252790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#252800000000
0!
0%
b0 *
0-
02
b0 6
#252810000000
1!
1%
1-
12
#252820000000
0!
0%
b1 *
0-
02
b1 6
#252830000000
1!
1%
1-
12
#252840000000
0!
0%
b10 *
0-
02
b10 6
#252850000000
1!
1%
1-
12
#252860000000
0!
0%
b11 *
0-
02
b11 6
#252870000000
1!
1%
1-
12
15
#252880000000
0!
0%
b100 *
0-
02
b100 6
#252890000000
1!
1%
1-
12
#252900000000
0!
0%
b101 *
0-
02
b101 6
#252910000000
1!
1%
1-
12
#252920000000
0!
0%
b110 *
0-
02
b110 6
#252930000000
1!
1%
1-
12
#252940000000
0!
0%
b111 *
0-
02
b111 6
#252950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#252960000000
0!
0%
b0 *
0-
02
b0 6
#252970000000
1!
1%
1-
12
#252980000000
0!
0%
b1 *
0-
02
b1 6
#252990000000
1!
1%
1-
12
#253000000000
0!
0%
b10 *
0-
02
b10 6
#253010000000
1!
1%
1-
12
#253020000000
0!
0%
b11 *
0-
02
b11 6
#253030000000
1!
1%
1-
12
15
#253040000000
0!
0%
b100 *
0-
02
b100 6
#253050000000
1!
1%
1-
12
#253060000000
0!
0%
b101 *
0-
02
b101 6
#253070000000
1!
1%
1-
12
#253080000000
0!
0%
b110 *
0-
02
b110 6
#253090000000
1!
1%
1-
12
#253100000000
0!
0%
b111 *
0-
02
b111 6
#253110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#253120000000
0!
0%
b0 *
0-
02
b0 6
#253130000000
1!
1%
1-
12
#253140000000
0!
0%
b1 *
0-
02
b1 6
#253150000000
1!
1%
1-
12
#253160000000
0!
0%
b10 *
0-
02
b10 6
#253170000000
1!
1%
1-
12
#253180000000
0!
0%
b11 *
0-
02
b11 6
#253190000000
1!
1%
1-
12
15
#253200000000
0!
0%
b100 *
0-
02
b100 6
#253210000000
1!
1%
1-
12
#253220000000
0!
0%
b101 *
0-
02
b101 6
#253230000000
1!
1%
1-
12
#253240000000
0!
0%
b110 *
0-
02
b110 6
#253250000000
1!
1%
1-
12
#253260000000
0!
0%
b111 *
0-
02
b111 6
#253270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#253280000000
0!
0%
b0 *
0-
02
b0 6
#253290000000
1!
1%
1-
12
#253300000000
0!
0%
b1 *
0-
02
b1 6
#253310000000
1!
1%
1-
12
#253320000000
0!
0%
b10 *
0-
02
b10 6
#253330000000
1!
1%
1-
12
#253340000000
0!
0%
b11 *
0-
02
b11 6
#253350000000
1!
1%
1-
12
15
#253360000000
0!
0%
b100 *
0-
02
b100 6
#253370000000
1!
1%
1-
12
#253380000000
0!
0%
b101 *
0-
02
b101 6
#253390000000
1!
1%
1-
12
#253400000000
0!
0%
b110 *
0-
02
b110 6
#253410000000
1!
1%
1-
12
#253420000000
0!
0%
b111 *
0-
02
b111 6
#253430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#253440000000
0!
0%
b0 *
0-
02
b0 6
#253450000000
1!
1%
1-
12
#253460000000
0!
0%
b1 *
0-
02
b1 6
#253470000000
1!
1%
1-
12
#253480000000
0!
0%
b10 *
0-
02
b10 6
#253490000000
1!
1%
1-
12
#253500000000
0!
0%
b11 *
0-
02
b11 6
#253510000000
1!
1%
1-
12
15
#253520000000
0!
0%
b100 *
0-
02
b100 6
#253530000000
1!
1%
1-
12
#253540000000
0!
0%
b101 *
0-
02
b101 6
#253550000000
1!
1%
1-
12
#253560000000
0!
0%
b110 *
0-
02
b110 6
#253570000000
1!
1%
1-
12
#253580000000
0!
0%
b111 *
0-
02
b111 6
#253590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#253600000000
0!
0%
b0 *
0-
02
b0 6
#253610000000
1!
1%
1-
12
#253620000000
0!
0%
b1 *
0-
02
b1 6
#253630000000
1!
1%
1-
12
#253640000000
0!
0%
b10 *
0-
02
b10 6
#253650000000
1!
1%
1-
12
#253660000000
0!
0%
b11 *
0-
02
b11 6
#253670000000
1!
1%
1-
12
15
#253680000000
0!
0%
b100 *
0-
02
b100 6
#253690000000
1!
1%
1-
12
#253700000000
0!
0%
b101 *
0-
02
b101 6
#253710000000
1!
1%
1-
12
#253720000000
0!
0%
b110 *
0-
02
b110 6
#253730000000
1!
1%
1-
12
#253740000000
0!
0%
b111 *
0-
02
b111 6
#253750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#253760000000
0!
0%
b0 *
0-
02
b0 6
#253770000000
1!
1%
1-
12
#253780000000
0!
0%
b1 *
0-
02
b1 6
#253790000000
1!
1%
1-
12
#253800000000
0!
0%
b10 *
0-
02
b10 6
#253810000000
1!
1%
1-
12
#253820000000
0!
0%
b11 *
0-
02
b11 6
#253830000000
1!
1%
1-
12
15
#253840000000
0!
0%
b100 *
0-
02
b100 6
#253850000000
1!
1%
1-
12
#253860000000
0!
0%
b101 *
0-
02
b101 6
#253870000000
1!
1%
1-
12
#253880000000
0!
0%
b110 *
0-
02
b110 6
#253890000000
1!
1%
1-
12
#253900000000
0!
0%
b111 *
0-
02
b111 6
#253910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#253920000000
0!
0%
b0 *
0-
02
b0 6
#253930000000
1!
1%
1-
12
#253940000000
0!
0%
b1 *
0-
02
b1 6
#253950000000
1!
1%
1-
12
#253960000000
0!
0%
b10 *
0-
02
b10 6
#253970000000
1!
1%
1-
12
#253980000000
0!
0%
b11 *
0-
02
b11 6
#253990000000
1!
1%
1-
12
15
#254000000000
0!
0%
b100 *
0-
02
b100 6
#254010000000
1!
1%
1-
12
#254020000000
0!
0%
b101 *
0-
02
b101 6
#254030000000
1!
1%
1-
12
#254040000000
0!
0%
b110 *
0-
02
b110 6
#254050000000
1!
1%
1-
12
#254060000000
0!
0%
b111 *
0-
02
b111 6
#254070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#254080000000
0!
0%
b0 *
0-
02
b0 6
#254090000000
1!
1%
1-
12
#254100000000
0!
0%
b1 *
0-
02
b1 6
#254110000000
1!
1%
1-
12
#254120000000
0!
0%
b10 *
0-
02
b10 6
#254130000000
1!
1%
1-
12
#254140000000
0!
0%
b11 *
0-
02
b11 6
#254150000000
1!
1%
1-
12
15
#254160000000
0!
0%
b100 *
0-
02
b100 6
#254170000000
1!
1%
1-
12
#254180000000
0!
0%
b101 *
0-
02
b101 6
#254190000000
1!
1%
1-
12
#254200000000
0!
0%
b110 *
0-
02
b110 6
#254210000000
1!
1%
1-
12
#254220000000
0!
0%
b111 *
0-
02
b111 6
#254230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#254240000000
0!
0%
b0 *
0-
02
b0 6
#254250000000
1!
1%
1-
12
#254260000000
0!
0%
b1 *
0-
02
b1 6
#254270000000
1!
1%
1-
12
#254280000000
0!
0%
b10 *
0-
02
b10 6
#254290000000
1!
1%
1-
12
#254300000000
0!
0%
b11 *
0-
02
b11 6
#254310000000
1!
1%
1-
12
15
#254320000000
0!
0%
b100 *
0-
02
b100 6
#254330000000
1!
1%
1-
12
#254340000000
0!
0%
b101 *
0-
02
b101 6
#254350000000
1!
1%
1-
12
#254360000000
0!
0%
b110 *
0-
02
b110 6
#254370000000
1!
1%
1-
12
#254380000000
0!
0%
b111 *
0-
02
b111 6
#254390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#254400000000
0!
0%
b0 *
0-
02
b0 6
#254410000000
1!
1%
1-
12
#254420000000
0!
0%
b1 *
0-
02
b1 6
#254430000000
1!
1%
1-
12
#254440000000
0!
0%
b10 *
0-
02
b10 6
#254450000000
1!
1%
1-
12
#254460000000
0!
0%
b11 *
0-
02
b11 6
#254470000000
1!
1%
1-
12
15
#254480000000
0!
0%
b100 *
0-
02
b100 6
#254490000000
1!
1%
1-
12
#254500000000
0!
0%
b101 *
0-
02
b101 6
#254510000000
1!
1%
1-
12
#254520000000
0!
0%
b110 *
0-
02
b110 6
#254530000000
1!
1%
1-
12
#254540000000
0!
0%
b111 *
0-
02
b111 6
#254550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#254560000000
0!
0%
b0 *
0-
02
b0 6
#254570000000
1!
1%
1-
12
#254580000000
0!
0%
b1 *
0-
02
b1 6
#254590000000
1!
1%
1-
12
#254600000000
0!
0%
b10 *
0-
02
b10 6
#254610000000
1!
1%
1-
12
#254620000000
0!
0%
b11 *
0-
02
b11 6
#254630000000
1!
1%
1-
12
15
#254640000000
0!
0%
b100 *
0-
02
b100 6
#254650000000
1!
1%
1-
12
#254660000000
0!
0%
b101 *
0-
02
b101 6
#254670000000
1!
1%
1-
12
#254680000000
0!
0%
b110 *
0-
02
b110 6
#254690000000
1!
1%
1-
12
#254700000000
0!
0%
b111 *
0-
02
b111 6
#254710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#254720000000
0!
0%
b0 *
0-
02
b0 6
#254730000000
1!
1%
1-
12
#254740000000
0!
0%
b1 *
0-
02
b1 6
#254750000000
1!
1%
1-
12
#254760000000
0!
0%
b10 *
0-
02
b10 6
#254770000000
1!
1%
1-
12
#254780000000
0!
0%
b11 *
0-
02
b11 6
#254790000000
1!
1%
1-
12
15
#254800000000
0!
0%
b100 *
0-
02
b100 6
#254810000000
1!
1%
1-
12
#254820000000
0!
0%
b101 *
0-
02
b101 6
#254830000000
1!
1%
1-
12
#254840000000
0!
0%
b110 *
0-
02
b110 6
#254850000000
1!
1%
1-
12
#254860000000
0!
0%
b111 *
0-
02
b111 6
#254870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#254880000000
0!
0%
b0 *
0-
02
b0 6
#254890000000
1!
1%
1-
12
#254900000000
0!
0%
b1 *
0-
02
b1 6
#254910000000
1!
1%
1-
12
#254920000000
0!
0%
b10 *
0-
02
b10 6
#254930000000
1!
1%
1-
12
#254940000000
0!
0%
b11 *
0-
02
b11 6
#254950000000
1!
1%
1-
12
15
#254960000000
0!
0%
b100 *
0-
02
b100 6
#254970000000
1!
1%
1-
12
#254980000000
0!
0%
b101 *
0-
02
b101 6
#254990000000
1!
1%
1-
12
#255000000000
0!
0%
b110 *
0-
02
b110 6
#255010000000
1!
1%
1-
12
#255020000000
0!
0%
b111 *
0-
02
b111 6
#255030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#255040000000
0!
0%
b0 *
0-
02
b0 6
#255050000000
1!
1%
1-
12
#255060000000
0!
0%
b1 *
0-
02
b1 6
#255070000000
1!
1%
1-
12
#255080000000
0!
0%
b10 *
0-
02
b10 6
#255090000000
1!
1%
1-
12
#255100000000
0!
0%
b11 *
0-
02
b11 6
#255110000000
1!
1%
1-
12
15
#255120000000
0!
0%
b100 *
0-
02
b100 6
#255130000000
1!
1%
1-
12
#255140000000
0!
0%
b101 *
0-
02
b101 6
#255150000000
1!
1%
1-
12
#255160000000
0!
0%
b110 *
0-
02
b110 6
#255170000000
1!
1%
1-
12
#255180000000
0!
0%
b111 *
0-
02
b111 6
#255190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#255200000000
0!
0%
b0 *
0-
02
b0 6
#255210000000
1!
1%
1-
12
#255220000000
0!
0%
b1 *
0-
02
b1 6
#255230000000
1!
1%
1-
12
#255240000000
0!
0%
b10 *
0-
02
b10 6
#255250000000
1!
1%
1-
12
#255260000000
0!
0%
b11 *
0-
02
b11 6
#255270000000
1!
1%
1-
12
15
#255280000000
0!
0%
b100 *
0-
02
b100 6
#255290000000
1!
1%
1-
12
#255300000000
0!
0%
b101 *
0-
02
b101 6
#255310000000
1!
1%
1-
12
#255320000000
0!
0%
b110 *
0-
02
b110 6
#255330000000
1!
1%
1-
12
#255340000000
0!
0%
b111 *
0-
02
b111 6
#255350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#255360000000
0!
0%
b0 *
0-
02
b0 6
#255370000000
1!
1%
1-
12
#255380000000
0!
0%
b1 *
0-
02
b1 6
#255390000000
1!
1%
1-
12
#255400000000
0!
0%
b10 *
0-
02
b10 6
#255410000000
1!
1%
1-
12
#255420000000
0!
0%
b11 *
0-
02
b11 6
#255430000000
1!
1%
1-
12
15
#255440000000
0!
0%
b100 *
0-
02
b100 6
#255450000000
1!
1%
1-
12
#255460000000
0!
0%
b101 *
0-
02
b101 6
#255470000000
1!
1%
1-
12
#255480000000
0!
0%
b110 *
0-
02
b110 6
#255490000000
1!
1%
1-
12
#255500000000
0!
0%
b111 *
0-
02
b111 6
#255510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#255520000000
0!
0%
b0 *
0-
02
b0 6
#255530000000
1!
1%
1-
12
#255540000000
0!
0%
b1 *
0-
02
b1 6
#255550000000
1!
1%
1-
12
#255560000000
0!
0%
b10 *
0-
02
b10 6
#255570000000
1!
1%
1-
12
#255580000000
0!
0%
b11 *
0-
02
b11 6
#255590000000
1!
1%
1-
12
15
#255600000000
0!
0%
b100 *
0-
02
b100 6
#255610000000
1!
1%
1-
12
#255620000000
0!
0%
b101 *
0-
02
b101 6
#255630000000
1!
1%
1-
12
#255640000000
0!
0%
b110 *
0-
02
b110 6
#255650000000
1!
1%
1-
12
#255660000000
0!
0%
b111 *
0-
02
b111 6
#255670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#255680000000
0!
0%
b0 *
0-
02
b0 6
#255690000000
1!
1%
1-
12
#255700000000
0!
0%
b1 *
0-
02
b1 6
#255710000000
1!
1%
1-
12
#255720000000
0!
0%
b10 *
0-
02
b10 6
#255730000000
1!
1%
1-
12
#255740000000
0!
0%
b11 *
0-
02
b11 6
#255750000000
1!
1%
1-
12
15
#255760000000
0!
0%
b100 *
0-
02
b100 6
#255770000000
1!
1%
1-
12
#255780000000
0!
0%
b101 *
0-
02
b101 6
#255790000000
1!
1%
1-
12
#255800000000
0!
0%
b110 *
0-
02
b110 6
#255810000000
1!
1%
1-
12
#255820000000
0!
0%
b111 *
0-
02
b111 6
#255830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#255840000000
0!
0%
b0 *
0-
02
b0 6
#255850000000
1!
1%
1-
12
#255860000000
0!
0%
b1 *
0-
02
b1 6
#255870000000
1!
1%
1-
12
#255880000000
0!
0%
b10 *
0-
02
b10 6
#255890000000
1!
1%
1-
12
#255900000000
0!
0%
b11 *
0-
02
b11 6
#255910000000
1!
1%
1-
12
15
#255920000000
0!
0%
b100 *
0-
02
b100 6
#255930000000
1!
1%
1-
12
#255940000000
0!
0%
b101 *
0-
02
b101 6
#255950000000
1!
1%
1-
12
#255960000000
0!
0%
b110 *
0-
02
b110 6
#255970000000
1!
1%
1-
12
#255980000000
0!
0%
b111 *
0-
02
b111 6
#255990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#256000000000
0!
0%
b0 *
0-
02
b0 6
#256010000000
1!
1%
1-
12
#256020000000
0!
0%
b1 *
0-
02
b1 6
#256030000000
1!
1%
1-
12
#256040000000
0!
0%
b10 *
0-
02
b10 6
#256050000000
1!
1%
1-
12
#256060000000
0!
0%
b11 *
0-
02
b11 6
#256070000000
1!
1%
1-
12
15
#256080000000
0!
0%
b100 *
0-
02
b100 6
#256090000000
1!
1%
1-
12
#256100000000
0!
0%
b101 *
0-
02
b101 6
#256110000000
1!
1%
1-
12
#256120000000
0!
0%
b110 *
0-
02
b110 6
#256130000000
1!
1%
1-
12
#256140000000
0!
0%
b111 *
0-
02
b111 6
#256150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#256160000000
0!
0%
b0 *
0-
02
b0 6
#256170000000
1!
1%
1-
12
#256180000000
0!
0%
b1 *
0-
02
b1 6
#256190000000
1!
1%
1-
12
#256200000000
0!
0%
b10 *
0-
02
b10 6
#256210000000
1!
1%
1-
12
#256220000000
0!
0%
b11 *
0-
02
b11 6
#256230000000
1!
1%
1-
12
15
#256240000000
0!
0%
b100 *
0-
02
b100 6
#256250000000
1!
1%
1-
12
#256260000000
0!
0%
b101 *
0-
02
b101 6
#256270000000
1!
1%
1-
12
#256280000000
0!
0%
b110 *
0-
02
b110 6
#256290000000
1!
1%
1-
12
#256300000000
0!
0%
b111 *
0-
02
b111 6
#256310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#256320000000
0!
0%
b0 *
0-
02
b0 6
#256330000000
1!
1%
1-
12
#256340000000
0!
0%
b1 *
0-
02
b1 6
#256350000000
1!
1%
1-
12
#256360000000
0!
0%
b10 *
0-
02
b10 6
#256370000000
1!
1%
1-
12
#256380000000
0!
0%
b11 *
0-
02
b11 6
#256390000000
1!
1%
1-
12
15
#256400000000
0!
0%
b100 *
0-
02
b100 6
#256410000000
1!
1%
1-
12
#256420000000
0!
0%
b101 *
0-
02
b101 6
#256430000000
1!
1%
1-
12
#256440000000
0!
0%
b110 *
0-
02
b110 6
#256450000000
1!
1%
1-
12
#256460000000
0!
0%
b111 *
0-
02
b111 6
#256470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#256480000000
0!
0%
b0 *
0-
02
b0 6
#256490000000
1!
1%
1-
12
#256500000000
0!
0%
b1 *
0-
02
b1 6
#256510000000
1!
1%
1-
12
#256520000000
0!
0%
b10 *
0-
02
b10 6
#256530000000
1!
1%
1-
12
#256540000000
0!
0%
b11 *
0-
02
b11 6
#256550000000
1!
1%
1-
12
15
#256560000000
0!
0%
b100 *
0-
02
b100 6
#256570000000
1!
1%
1-
12
#256580000000
0!
0%
b101 *
0-
02
b101 6
#256590000000
1!
1%
1-
12
#256600000000
0!
0%
b110 *
0-
02
b110 6
#256610000000
1!
1%
1-
12
#256620000000
0!
0%
b111 *
0-
02
b111 6
#256630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#256640000000
0!
0%
b0 *
0-
02
b0 6
#256650000000
1!
1%
1-
12
#256660000000
0!
0%
b1 *
0-
02
b1 6
#256670000000
1!
1%
1-
12
#256680000000
0!
0%
b10 *
0-
02
b10 6
#256690000000
1!
1%
1-
12
#256700000000
0!
0%
b11 *
0-
02
b11 6
#256710000000
1!
1%
1-
12
15
#256720000000
0!
0%
b100 *
0-
02
b100 6
#256730000000
1!
1%
1-
12
#256740000000
0!
0%
b101 *
0-
02
b101 6
#256750000000
1!
1%
1-
12
#256760000000
0!
0%
b110 *
0-
02
b110 6
#256770000000
1!
1%
1-
12
#256780000000
0!
0%
b111 *
0-
02
b111 6
#256790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#256800000000
0!
0%
b0 *
0-
02
b0 6
#256810000000
1!
1%
1-
12
#256820000000
0!
0%
b1 *
0-
02
b1 6
#256830000000
1!
1%
1-
12
#256840000000
0!
0%
b10 *
0-
02
b10 6
#256850000000
1!
1%
1-
12
#256860000000
0!
0%
b11 *
0-
02
b11 6
#256870000000
1!
1%
1-
12
15
#256880000000
0!
0%
b100 *
0-
02
b100 6
#256890000000
1!
1%
1-
12
#256900000000
0!
0%
b101 *
0-
02
b101 6
#256910000000
1!
1%
1-
12
#256920000000
0!
0%
b110 *
0-
02
b110 6
#256930000000
1!
1%
1-
12
#256940000000
0!
0%
b111 *
0-
02
b111 6
#256950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#256960000000
0!
0%
b0 *
0-
02
b0 6
#256970000000
1!
1%
1-
12
#256980000000
0!
0%
b1 *
0-
02
b1 6
#256990000000
1!
1%
1-
12
#257000000000
0!
0%
b10 *
0-
02
b10 6
#257010000000
1!
1%
1-
12
#257020000000
0!
0%
b11 *
0-
02
b11 6
#257030000000
1!
1%
1-
12
15
#257040000000
0!
0%
b100 *
0-
02
b100 6
#257050000000
1!
1%
1-
12
#257060000000
0!
0%
b101 *
0-
02
b101 6
#257070000000
1!
1%
1-
12
#257080000000
0!
0%
b110 *
0-
02
b110 6
#257090000000
1!
1%
1-
12
#257100000000
0!
0%
b111 *
0-
02
b111 6
#257110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#257120000000
0!
0%
b0 *
0-
02
b0 6
#257130000000
1!
1%
1-
12
#257140000000
0!
0%
b1 *
0-
02
b1 6
#257150000000
1!
1%
1-
12
#257160000000
0!
0%
b10 *
0-
02
b10 6
#257170000000
1!
1%
1-
12
#257180000000
0!
0%
b11 *
0-
02
b11 6
#257190000000
1!
1%
1-
12
15
#257200000000
0!
0%
b100 *
0-
02
b100 6
#257210000000
1!
1%
1-
12
#257220000000
0!
0%
b101 *
0-
02
b101 6
#257230000000
1!
1%
1-
12
#257240000000
0!
0%
b110 *
0-
02
b110 6
#257250000000
1!
1%
1-
12
#257260000000
0!
0%
b111 *
0-
02
b111 6
#257270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#257280000000
0!
0%
b0 *
0-
02
b0 6
#257290000000
1!
1%
1-
12
#257300000000
0!
0%
b1 *
0-
02
b1 6
#257310000000
1!
1%
1-
12
#257320000000
0!
0%
b10 *
0-
02
b10 6
#257330000000
1!
1%
1-
12
#257340000000
0!
0%
b11 *
0-
02
b11 6
#257350000000
1!
1%
1-
12
15
#257360000000
0!
0%
b100 *
0-
02
b100 6
#257370000000
1!
1%
1-
12
#257380000000
0!
0%
b101 *
0-
02
b101 6
#257390000000
1!
1%
1-
12
#257400000000
0!
0%
b110 *
0-
02
b110 6
#257410000000
1!
1%
1-
12
#257420000000
0!
0%
b111 *
0-
02
b111 6
#257430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#257440000000
0!
0%
b0 *
0-
02
b0 6
#257450000000
1!
1%
1-
12
#257460000000
0!
0%
b1 *
0-
02
b1 6
#257470000000
1!
1%
1-
12
#257480000000
0!
0%
b10 *
0-
02
b10 6
#257490000000
1!
1%
1-
12
#257500000000
0!
0%
b11 *
0-
02
b11 6
#257510000000
1!
1%
1-
12
15
#257520000000
0!
0%
b100 *
0-
02
b100 6
#257530000000
1!
1%
1-
12
#257540000000
0!
0%
b101 *
0-
02
b101 6
#257550000000
1!
1%
1-
12
#257560000000
0!
0%
b110 *
0-
02
b110 6
#257570000000
1!
1%
1-
12
#257580000000
0!
0%
b111 *
0-
02
b111 6
#257590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#257600000000
0!
0%
b0 *
0-
02
b0 6
#257610000000
1!
1%
1-
12
#257620000000
0!
0%
b1 *
0-
02
b1 6
#257630000000
1!
1%
1-
12
#257640000000
0!
0%
b10 *
0-
02
b10 6
#257650000000
1!
1%
1-
12
#257660000000
0!
0%
b11 *
0-
02
b11 6
#257670000000
1!
1%
1-
12
15
#257680000000
0!
0%
b100 *
0-
02
b100 6
#257690000000
1!
1%
1-
12
#257700000000
0!
0%
b101 *
0-
02
b101 6
#257710000000
1!
1%
1-
12
#257720000000
0!
0%
b110 *
0-
02
b110 6
#257730000000
1!
1%
1-
12
#257740000000
0!
0%
b111 *
0-
02
b111 6
#257750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#257760000000
0!
0%
b0 *
0-
02
b0 6
#257770000000
1!
1%
1-
12
#257780000000
0!
0%
b1 *
0-
02
b1 6
#257790000000
1!
1%
1-
12
#257800000000
0!
0%
b10 *
0-
02
b10 6
#257810000000
1!
1%
1-
12
#257820000000
0!
0%
b11 *
0-
02
b11 6
#257830000000
1!
1%
1-
12
15
#257840000000
0!
0%
b100 *
0-
02
b100 6
#257850000000
1!
1%
1-
12
#257860000000
0!
0%
b101 *
0-
02
b101 6
#257870000000
1!
1%
1-
12
#257880000000
0!
0%
b110 *
0-
02
b110 6
#257890000000
1!
1%
1-
12
#257900000000
0!
0%
b111 *
0-
02
b111 6
#257910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#257920000000
0!
0%
b0 *
0-
02
b0 6
#257930000000
1!
1%
1-
12
#257940000000
0!
0%
b1 *
0-
02
b1 6
#257950000000
1!
1%
1-
12
#257960000000
0!
0%
b10 *
0-
02
b10 6
#257970000000
1!
1%
1-
12
#257980000000
0!
0%
b11 *
0-
02
b11 6
#257990000000
1!
1%
1-
12
15
#258000000000
0!
0%
b100 *
0-
02
b100 6
#258010000000
1!
1%
1-
12
#258020000000
0!
0%
b101 *
0-
02
b101 6
#258030000000
1!
1%
1-
12
#258040000000
0!
0%
b110 *
0-
02
b110 6
#258050000000
1!
1%
1-
12
#258060000000
0!
0%
b111 *
0-
02
b111 6
#258070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#258080000000
0!
0%
b0 *
0-
02
b0 6
#258090000000
1!
1%
1-
12
#258100000000
0!
0%
b1 *
0-
02
b1 6
#258110000000
1!
1%
1-
12
#258120000000
0!
0%
b10 *
0-
02
b10 6
#258130000000
1!
1%
1-
12
#258140000000
0!
0%
b11 *
0-
02
b11 6
#258150000000
1!
1%
1-
12
15
#258160000000
0!
0%
b100 *
0-
02
b100 6
#258170000000
1!
1%
1-
12
#258180000000
0!
0%
b101 *
0-
02
b101 6
#258190000000
1!
1%
1-
12
#258200000000
0!
0%
b110 *
0-
02
b110 6
#258210000000
1!
1%
1-
12
#258220000000
0!
0%
b111 *
0-
02
b111 6
#258230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#258240000000
0!
0%
b0 *
0-
02
b0 6
#258250000000
1!
1%
1-
12
#258260000000
0!
0%
b1 *
0-
02
b1 6
#258270000000
1!
1%
1-
12
#258280000000
0!
0%
b10 *
0-
02
b10 6
#258290000000
1!
1%
1-
12
#258300000000
0!
0%
b11 *
0-
02
b11 6
#258310000000
1!
1%
1-
12
15
#258320000000
0!
0%
b100 *
0-
02
b100 6
#258330000000
1!
1%
1-
12
#258340000000
0!
0%
b101 *
0-
02
b101 6
#258350000000
1!
1%
1-
12
#258360000000
0!
0%
b110 *
0-
02
b110 6
#258370000000
1!
1%
1-
12
#258380000000
0!
0%
b111 *
0-
02
b111 6
#258390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#258400000000
0!
0%
b0 *
0-
02
b0 6
#258410000000
1!
1%
1-
12
#258420000000
0!
0%
b1 *
0-
02
b1 6
#258430000000
1!
1%
1-
12
#258440000000
0!
0%
b10 *
0-
02
b10 6
#258450000000
1!
1%
1-
12
#258460000000
0!
0%
b11 *
0-
02
b11 6
#258470000000
1!
1%
1-
12
15
#258480000000
0!
0%
b100 *
0-
02
b100 6
#258490000000
1!
1%
1-
12
#258500000000
0!
0%
b101 *
0-
02
b101 6
#258510000000
1!
1%
1-
12
#258520000000
0!
0%
b110 *
0-
02
b110 6
#258530000000
1!
1%
1-
12
#258540000000
0!
0%
b111 *
0-
02
b111 6
#258550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#258560000000
0!
0%
b0 *
0-
02
b0 6
#258570000000
1!
1%
1-
12
#258580000000
0!
0%
b1 *
0-
02
b1 6
#258590000000
1!
1%
1-
12
#258600000000
0!
0%
b10 *
0-
02
b10 6
#258610000000
1!
1%
1-
12
#258620000000
0!
0%
b11 *
0-
02
b11 6
#258630000000
1!
1%
1-
12
15
#258640000000
0!
0%
b100 *
0-
02
b100 6
#258650000000
1!
1%
1-
12
#258660000000
0!
0%
b101 *
0-
02
b101 6
#258670000000
1!
1%
1-
12
#258680000000
0!
0%
b110 *
0-
02
b110 6
#258690000000
1!
1%
1-
12
#258700000000
0!
0%
b111 *
0-
02
b111 6
#258710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#258720000000
0!
0%
b0 *
0-
02
b0 6
#258730000000
1!
1%
1-
12
#258740000000
0!
0%
b1 *
0-
02
b1 6
#258750000000
1!
1%
1-
12
#258760000000
0!
0%
b10 *
0-
02
b10 6
#258770000000
1!
1%
1-
12
#258780000000
0!
0%
b11 *
0-
02
b11 6
#258790000000
1!
1%
1-
12
15
#258800000000
0!
0%
b100 *
0-
02
b100 6
#258810000000
1!
1%
1-
12
#258820000000
0!
0%
b101 *
0-
02
b101 6
#258830000000
1!
1%
1-
12
#258840000000
0!
0%
b110 *
0-
02
b110 6
#258850000000
1!
1%
1-
12
#258860000000
0!
0%
b111 *
0-
02
b111 6
#258870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#258880000000
0!
0%
b0 *
0-
02
b0 6
#258890000000
1!
1%
1-
12
#258900000000
0!
0%
b1 *
0-
02
b1 6
#258910000000
1!
1%
1-
12
#258920000000
0!
0%
b10 *
0-
02
b10 6
#258930000000
1!
1%
1-
12
#258940000000
0!
0%
b11 *
0-
02
b11 6
#258950000000
1!
1%
1-
12
15
#258960000000
0!
0%
b100 *
0-
02
b100 6
#258970000000
1!
1%
1-
12
#258980000000
0!
0%
b101 *
0-
02
b101 6
#258990000000
1!
1%
1-
12
#259000000000
0!
0%
b110 *
0-
02
b110 6
#259010000000
1!
1%
1-
12
#259020000000
0!
0%
b111 *
0-
02
b111 6
#259030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#259040000000
0!
0%
b0 *
0-
02
b0 6
#259050000000
1!
1%
1-
12
#259060000000
0!
0%
b1 *
0-
02
b1 6
#259070000000
1!
1%
1-
12
#259080000000
0!
0%
b10 *
0-
02
b10 6
#259090000000
1!
1%
1-
12
#259100000000
0!
0%
b11 *
0-
02
b11 6
#259110000000
1!
1%
1-
12
15
#259120000000
0!
0%
b100 *
0-
02
b100 6
#259130000000
1!
1%
1-
12
#259140000000
0!
0%
b101 *
0-
02
b101 6
#259150000000
1!
1%
1-
12
#259160000000
0!
0%
b110 *
0-
02
b110 6
#259170000000
1!
1%
1-
12
#259180000000
0!
0%
b111 *
0-
02
b111 6
#259190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#259200000000
0!
0%
b0 *
0-
02
b0 6
#259210000000
1!
1%
1-
12
#259220000000
0!
0%
b1 *
0-
02
b1 6
#259230000000
1!
1%
1-
12
#259240000000
0!
0%
b10 *
0-
02
b10 6
#259250000000
1!
1%
1-
12
#259260000000
0!
0%
b11 *
0-
02
b11 6
#259270000000
1!
1%
1-
12
15
#259280000000
0!
0%
b100 *
0-
02
b100 6
#259290000000
1!
1%
1-
12
#259300000000
0!
0%
b101 *
0-
02
b101 6
#259310000000
1!
1%
1-
12
#259320000000
0!
0%
b110 *
0-
02
b110 6
#259330000000
1!
1%
1-
12
#259340000000
0!
0%
b111 *
0-
02
b111 6
#259350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#259360000000
0!
0%
b0 *
0-
02
b0 6
#259370000000
1!
1%
1-
12
#259380000000
0!
0%
b1 *
0-
02
b1 6
#259390000000
1!
1%
1-
12
#259400000000
0!
0%
b10 *
0-
02
b10 6
#259410000000
1!
1%
1-
12
#259420000000
0!
0%
b11 *
0-
02
b11 6
#259430000000
1!
1%
1-
12
15
#259440000000
0!
0%
b100 *
0-
02
b100 6
#259450000000
1!
1%
1-
12
#259460000000
0!
0%
b101 *
0-
02
b101 6
#259470000000
1!
1%
1-
12
#259480000000
0!
0%
b110 *
0-
02
b110 6
#259490000000
1!
1%
1-
12
#259500000000
0!
0%
b111 *
0-
02
b111 6
#259510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#259520000000
0!
0%
b0 *
0-
02
b0 6
#259530000000
1!
1%
1-
12
#259540000000
0!
0%
b1 *
0-
02
b1 6
#259550000000
1!
1%
1-
12
#259560000000
0!
0%
b10 *
0-
02
b10 6
#259570000000
1!
1%
1-
12
#259580000000
0!
0%
b11 *
0-
02
b11 6
#259590000000
1!
1%
1-
12
15
#259600000000
0!
0%
b100 *
0-
02
b100 6
#259610000000
1!
1%
1-
12
#259620000000
0!
0%
b101 *
0-
02
b101 6
#259630000000
1!
1%
1-
12
#259640000000
0!
0%
b110 *
0-
02
b110 6
#259650000000
1!
1%
1-
12
#259660000000
0!
0%
b111 *
0-
02
b111 6
#259670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#259680000000
0!
0%
b0 *
0-
02
b0 6
#259690000000
1!
1%
1-
12
#259700000000
0!
0%
b1 *
0-
02
b1 6
#259710000000
1!
1%
1-
12
#259720000000
0!
0%
b10 *
0-
02
b10 6
#259730000000
1!
1%
1-
12
#259740000000
0!
0%
b11 *
0-
02
b11 6
#259750000000
1!
1%
1-
12
15
#259760000000
0!
0%
b100 *
0-
02
b100 6
#259770000000
1!
1%
1-
12
#259780000000
0!
0%
b101 *
0-
02
b101 6
#259790000000
1!
1%
1-
12
#259800000000
0!
0%
b110 *
0-
02
b110 6
#259810000000
1!
1%
1-
12
#259820000000
0!
0%
b111 *
0-
02
b111 6
#259830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#259840000000
0!
0%
b0 *
0-
02
b0 6
#259850000000
1!
1%
1-
12
#259860000000
0!
0%
b1 *
0-
02
b1 6
#259870000000
1!
1%
1-
12
#259880000000
0!
0%
b10 *
0-
02
b10 6
#259890000000
1!
1%
1-
12
#259900000000
0!
0%
b11 *
0-
02
b11 6
#259910000000
1!
1%
1-
12
15
#259920000000
0!
0%
b100 *
0-
02
b100 6
#259930000000
1!
1%
1-
12
#259940000000
0!
0%
b101 *
0-
02
b101 6
#259950000000
1!
1%
1-
12
#259960000000
0!
0%
b110 *
0-
02
b110 6
#259970000000
1!
1%
1-
12
#259980000000
0!
0%
b111 *
0-
02
b111 6
#259990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#260000000000
0!
0%
b0 *
0-
02
b0 6
#260010000000
1!
1%
1-
12
#260020000000
0!
0%
b1 *
0-
02
b1 6
#260030000000
1!
1%
1-
12
#260040000000
0!
0%
b10 *
0-
02
b10 6
#260050000000
1!
1%
1-
12
#260060000000
0!
0%
b11 *
0-
02
b11 6
#260070000000
1!
1%
1-
12
15
#260080000000
0!
0%
b100 *
0-
02
b100 6
#260090000000
1!
1%
1-
12
#260100000000
0!
0%
b101 *
0-
02
b101 6
#260110000000
1!
1%
1-
12
#260120000000
0!
0%
b110 *
0-
02
b110 6
#260130000000
1!
1%
1-
12
#260140000000
0!
0%
b111 *
0-
02
b111 6
#260150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#260160000000
0!
0%
b0 *
0-
02
b0 6
#260170000000
1!
1%
1-
12
#260180000000
0!
0%
b1 *
0-
02
b1 6
#260190000000
1!
1%
1-
12
#260200000000
0!
0%
b10 *
0-
02
b10 6
#260210000000
1!
1%
1-
12
#260220000000
0!
0%
b11 *
0-
02
b11 6
#260230000000
1!
1%
1-
12
15
#260240000000
0!
0%
b100 *
0-
02
b100 6
#260250000000
1!
1%
1-
12
#260260000000
0!
0%
b101 *
0-
02
b101 6
#260270000000
1!
1%
1-
12
#260280000000
0!
0%
b110 *
0-
02
b110 6
#260290000000
1!
1%
1-
12
#260300000000
0!
0%
b111 *
0-
02
b111 6
#260310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#260320000000
0!
0%
b0 *
0-
02
b0 6
#260330000000
1!
1%
1-
12
#260340000000
0!
0%
b1 *
0-
02
b1 6
#260350000000
1!
1%
1-
12
#260360000000
0!
0%
b10 *
0-
02
b10 6
#260370000000
1!
1%
1-
12
#260380000000
0!
0%
b11 *
0-
02
b11 6
#260390000000
1!
1%
1-
12
15
#260400000000
0!
0%
b100 *
0-
02
b100 6
#260410000000
1!
1%
1-
12
#260420000000
0!
0%
b101 *
0-
02
b101 6
#260430000000
1!
1%
1-
12
#260440000000
0!
0%
b110 *
0-
02
b110 6
#260450000000
1!
1%
1-
12
#260460000000
0!
0%
b111 *
0-
02
b111 6
#260470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#260480000000
0!
0%
b0 *
0-
02
b0 6
#260490000000
1!
1%
1-
12
#260500000000
0!
0%
b1 *
0-
02
b1 6
#260510000000
1!
1%
1-
12
#260520000000
0!
0%
b10 *
0-
02
b10 6
#260530000000
1!
1%
1-
12
#260540000000
0!
0%
b11 *
0-
02
b11 6
#260550000000
1!
1%
1-
12
15
#260560000000
0!
0%
b100 *
0-
02
b100 6
#260570000000
1!
1%
1-
12
#260580000000
0!
0%
b101 *
0-
02
b101 6
#260590000000
1!
1%
1-
12
#260600000000
0!
0%
b110 *
0-
02
b110 6
#260610000000
1!
1%
1-
12
#260620000000
0!
0%
b111 *
0-
02
b111 6
#260630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#260640000000
0!
0%
b0 *
0-
02
b0 6
#260650000000
1!
1%
1-
12
#260660000000
0!
0%
b1 *
0-
02
b1 6
#260670000000
1!
1%
1-
12
#260680000000
0!
0%
b10 *
0-
02
b10 6
#260690000000
1!
1%
1-
12
#260700000000
0!
0%
b11 *
0-
02
b11 6
#260710000000
1!
1%
1-
12
15
#260720000000
0!
0%
b100 *
0-
02
b100 6
#260730000000
1!
1%
1-
12
#260740000000
0!
0%
b101 *
0-
02
b101 6
#260750000000
1!
1%
1-
12
#260760000000
0!
0%
b110 *
0-
02
b110 6
#260770000000
1!
1%
1-
12
#260780000000
0!
0%
b111 *
0-
02
b111 6
#260790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#260800000000
0!
0%
b0 *
0-
02
b0 6
#260810000000
1!
1%
1-
12
#260820000000
0!
0%
b1 *
0-
02
b1 6
#260830000000
1!
1%
1-
12
#260840000000
0!
0%
b10 *
0-
02
b10 6
#260850000000
1!
1%
1-
12
#260860000000
0!
0%
b11 *
0-
02
b11 6
#260870000000
1!
1%
1-
12
15
#260880000000
0!
0%
b100 *
0-
02
b100 6
#260890000000
1!
1%
1-
12
#260900000000
0!
0%
b101 *
0-
02
b101 6
#260910000000
1!
1%
1-
12
#260920000000
0!
0%
b110 *
0-
02
b110 6
#260930000000
1!
1%
1-
12
#260940000000
0!
0%
b111 *
0-
02
b111 6
#260950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#260960000000
0!
0%
b0 *
0-
02
b0 6
#260970000000
1!
1%
1-
12
#260980000000
0!
0%
b1 *
0-
02
b1 6
#260990000000
1!
1%
1-
12
#261000000000
0!
0%
b10 *
0-
02
b10 6
#261010000000
1!
1%
1-
12
#261020000000
0!
0%
b11 *
0-
02
b11 6
#261030000000
1!
1%
1-
12
15
#261040000000
0!
0%
b100 *
0-
02
b100 6
#261050000000
1!
1%
1-
12
#261060000000
0!
0%
b101 *
0-
02
b101 6
#261070000000
1!
1%
1-
12
#261080000000
0!
0%
b110 *
0-
02
b110 6
#261090000000
1!
1%
1-
12
#261100000000
0!
0%
b111 *
0-
02
b111 6
#261110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#261120000000
0!
0%
b0 *
0-
02
b0 6
#261130000000
1!
1%
1-
12
#261140000000
0!
0%
b1 *
0-
02
b1 6
#261150000000
1!
1%
1-
12
#261160000000
0!
0%
b10 *
0-
02
b10 6
#261170000000
1!
1%
1-
12
#261180000000
0!
0%
b11 *
0-
02
b11 6
#261190000000
1!
1%
1-
12
15
#261200000000
0!
0%
b100 *
0-
02
b100 6
#261210000000
1!
1%
1-
12
#261220000000
0!
0%
b101 *
0-
02
b101 6
#261230000000
1!
1%
1-
12
#261240000000
0!
0%
b110 *
0-
02
b110 6
#261250000000
1!
1%
1-
12
#261260000000
0!
0%
b111 *
0-
02
b111 6
#261270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#261280000000
0!
0%
b0 *
0-
02
b0 6
#261290000000
1!
1%
1-
12
#261300000000
0!
0%
b1 *
0-
02
b1 6
#261310000000
1!
1%
1-
12
#261320000000
0!
0%
b10 *
0-
02
b10 6
#261330000000
1!
1%
1-
12
#261340000000
0!
0%
b11 *
0-
02
b11 6
#261350000000
1!
1%
1-
12
15
#261360000000
0!
0%
b100 *
0-
02
b100 6
#261370000000
1!
1%
1-
12
#261380000000
0!
0%
b101 *
0-
02
b101 6
#261390000000
1!
1%
1-
12
#261400000000
0!
0%
b110 *
0-
02
b110 6
#261410000000
1!
1%
1-
12
#261420000000
0!
0%
b111 *
0-
02
b111 6
#261430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#261440000000
0!
0%
b0 *
0-
02
b0 6
#261450000000
1!
1%
1-
12
#261460000000
0!
0%
b1 *
0-
02
b1 6
#261470000000
1!
1%
1-
12
#261480000000
0!
0%
b10 *
0-
02
b10 6
#261490000000
1!
1%
1-
12
#261500000000
0!
0%
b11 *
0-
02
b11 6
#261510000000
1!
1%
1-
12
15
#261520000000
0!
0%
b100 *
0-
02
b100 6
#261530000000
1!
1%
1-
12
#261540000000
0!
0%
b101 *
0-
02
b101 6
#261550000000
1!
1%
1-
12
#261560000000
0!
0%
b110 *
0-
02
b110 6
#261570000000
1!
1%
1-
12
#261580000000
0!
0%
b111 *
0-
02
b111 6
#261590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#261600000000
0!
0%
b0 *
0-
02
b0 6
#261610000000
1!
1%
1-
12
#261620000000
0!
0%
b1 *
0-
02
b1 6
#261630000000
1!
1%
1-
12
#261640000000
0!
0%
b10 *
0-
02
b10 6
#261650000000
1!
1%
1-
12
#261660000000
0!
0%
b11 *
0-
02
b11 6
#261670000000
1!
1%
1-
12
15
#261680000000
0!
0%
b100 *
0-
02
b100 6
#261690000000
1!
1%
1-
12
#261700000000
0!
0%
b101 *
0-
02
b101 6
#261710000000
1!
1%
1-
12
#261720000000
0!
0%
b110 *
0-
02
b110 6
#261730000000
1!
1%
1-
12
#261740000000
0!
0%
b111 *
0-
02
b111 6
#261750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#261760000000
0!
0%
b0 *
0-
02
b0 6
#261770000000
1!
1%
1-
12
#261780000000
0!
0%
b1 *
0-
02
b1 6
#261790000000
1!
1%
1-
12
#261800000000
0!
0%
b10 *
0-
02
b10 6
#261810000000
1!
1%
1-
12
#261820000000
0!
0%
b11 *
0-
02
b11 6
#261830000000
1!
1%
1-
12
15
#261840000000
0!
0%
b100 *
0-
02
b100 6
#261850000000
1!
1%
1-
12
#261860000000
0!
0%
b101 *
0-
02
b101 6
#261870000000
1!
1%
1-
12
#261880000000
0!
0%
b110 *
0-
02
b110 6
#261890000000
1!
1%
1-
12
#261900000000
0!
0%
b111 *
0-
02
b111 6
#261910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#261920000000
0!
0%
b0 *
0-
02
b0 6
#261930000000
1!
1%
1-
12
#261940000000
0!
0%
b1 *
0-
02
b1 6
#261950000000
1!
1%
1-
12
#261960000000
0!
0%
b10 *
0-
02
b10 6
#261970000000
1!
1%
1-
12
#261980000000
0!
0%
b11 *
0-
02
b11 6
#261990000000
1!
1%
1-
12
15
#262000000000
0!
0%
b100 *
0-
02
b100 6
#262010000000
1!
1%
1-
12
#262020000000
0!
0%
b101 *
0-
02
b101 6
#262030000000
1!
1%
1-
12
#262040000000
0!
0%
b110 *
0-
02
b110 6
#262050000000
1!
1%
1-
12
#262060000000
0!
0%
b111 *
0-
02
b111 6
#262070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#262080000000
0!
0%
b0 *
0-
02
b0 6
#262090000000
1!
1%
1-
12
#262100000000
0!
0%
b1 *
0-
02
b1 6
#262110000000
1!
1%
1-
12
#262120000000
0!
0%
b10 *
0-
02
b10 6
#262130000000
1!
1%
1-
12
#262140000000
0!
0%
b11 *
0-
02
b11 6
#262150000000
1!
1%
1-
12
15
#262160000000
0!
0%
b100 *
0-
02
b100 6
#262170000000
1!
1%
1-
12
#262180000000
0!
0%
b101 *
0-
02
b101 6
#262190000000
1!
1%
1-
12
#262200000000
0!
0%
b110 *
0-
02
b110 6
#262210000000
1!
1%
1-
12
#262220000000
0!
0%
b111 *
0-
02
b111 6
#262230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#262240000000
0!
0%
b0 *
0-
02
b0 6
#262250000000
1!
1%
1-
12
#262260000000
0!
0%
b1 *
0-
02
b1 6
#262270000000
1!
1%
1-
12
#262280000000
0!
0%
b10 *
0-
02
b10 6
#262290000000
1!
1%
1-
12
#262300000000
0!
0%
b11 *
0-
02
b11 6
#262310000000
1!
1%
1-
12
15
#262320000000
0!
0%
b100 *
0-
02
b100 6
#262330000000
1!
1%
1-
12
#262340000000
0!
0%
b101 *
0-
02
b101 6
#262350000000
1!
1%
1-
12
#262360000000
0!
0%
b110 *
0-
02
b110 6
#262370000000
1!
1%
1-
12
#262380000000
0!
0%
b111 *
0-
02
b111 6
#262390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#262400000000
0!
0%
b0 *
0-
02
b0 6
#262410000000
1!
1%
1-
12
#262420000000
0!
0%
b1 *
0-
02
b1 6
#262430000000
1!
1%
1-
12
#262440000000
0!
0%
b10 *
0-
02
b10 6
#262450000000
1!
1%
1-
12
#262460000000
0!
0%
b11 *
0-
02
b11 6
#262470000000
1!
1%
1-
12
15
#262480000000
0!
0%
b100 *
0-
02
b100 6
#262490000000
1!
1%
1-
12
#262500000000
0!
0%
b101 *
0-
02
b101 6
#262510000000
1!
1%
1-
12
#262520000000
0!
0%
b110 *
0-
02
b110 6
#262530000000
1!
1%
1-
12
#262540000000
0!
0%
b111 *
0-
02
b111 6
#262550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#262560000000
0!
0%
b0 *
0-
02
b0 6
#262570000000
1!
1%
1-
12
#262580000000
0!
0%
b1 *
0-
02
b1 6
#262590000000
1!
1%
1-
12
#262600000000
0!
0%
b10 *
0-
02
b10 6
#262610000000
1!
1%
1-
12
#262620000000
0!
0%
b11 *
0-
02
b11 6
#262630000000
1!
1%
1-
12
15
#262640000000
0!
0%
b100 *
0-
02
b100 6
#262650000000
1!
1%
1-
12
#262660000000
0!
0%
b101 *
0-
02
b101 6
#262670000000
1!
1%
1-
12
#262680000000
0!
0%
b110 *
0-
02
b110 6
#262690000000
1!
1%
1-
12
#262700000000
0!
0%
b111 *
0-
02
b111 6
#262710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#262720000000
0!
0%
b0 *
0-
02
b0 6
#262730000000
1!
1%
1-
12
#262740000000
0!
0%
b1 *
0-
02
b1 6
#262750000000
1!
1%
1-
12
#262760000000
0!
0%
b10 *
0-
02
b10 6
#262770000000
1!
1%
1-
12
#262780000000
0!
0%
b11 *
0-
02
b11 6
#262790000000
1!
1%
1-
12
15
#262800000000
0!
0%
b100 *
0-
02
b100 6
#262810000000
1!
1%
1-
12
#262820000000
0!
0%
b101 *
0-
02
b101 6
#262830000000
1!
1%
1-
12
#262840000000
0!
0%
b110 *
0-
02
b110 6
#262850000000
1!
1%
1-
12
#262860000000
0!
0%
b111 *
0-
02
b111 6
#262870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#262880000000
0!
0%
b0 *
0-
02
b0 6
#262890000000
1!
1%
1-
12
#262900000000
0!
0%
b1 *
0-
02
b1 6
#262910000000
1!
1%
1-
12
#262920000000
0!
0%
b10 *
0-
02
b10 6
#262930000000
1!
1%
1-
12
#262940000000
0!
0%
b11 *
0-
02
b11 6
#262950000000
1!
1%
1-
12
15
#262960000000
0!
0%
b100 *
0-
02
b100 6
#262970000000
1!
1%
1-
12
#262980000000
0!
0%
b101 *
0-
02
b101 6
#262990000000
1!
1%
1-
12
#263000000000
0!
0%
b110 *
0-
02
b110 6
#263010000000
1!
1%
1-
12
#263020000000
0!
0%
b111 *
0-
02
b111 6
#263030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#263040000000
0!
0%
b0 *
0-
02
b0 6
#263050000000
1!
1%
1-
12
#263060000000
0!
0%
b1 *
0-
02
b1 6
#263070000000
1!
1%
1-
12
#263080000000
0!
0%
b10 *
0-
02
b10 6
#263090000000
1!
1%
1-
12
#263100000000
0!
0%
b11 *
0-
02
b11 6
#263110000000
1!
1%
1-
12
15
#263120000000
0!
0%
b100 *
0-
02
b100 6
#263130000000
1!
1%
1-
12
#263140000000
0!
0%
b101 *
0-
02
b101 6
#263150000000
1!
1%
1-
12
#263160000000
0!
0%
b110 *
0-
02
b110 6
#263170000000
1!
1%
1-
12
#263180000000
0!
0%
b111 *
0-
02
b111 6
#263190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#263200000000
0!
0%
b0 *
0-
02
b0 6
#263210000000
1!
1%
1-
12
#263220000000
0!
0%
b1 *
0-
02
b1 6
#263230000000
1!
1%
1-
12
#263240000000
0!
0%
b10 *
0-
02
b10 6
#263250000000
1!
1%
1-
12
#263260000000
0!
0%
b11 *
0-
02
b11 6
#263270000000
1!
1%
1-
12
15
#263280000000
0!
0%
b100 *
0-
02
b100 6
#263290000000
1!
1%
1-
12
#263300000000
0!
0%
b101 *
0-
02
b101 6
#263310000000
1!
1%
1-
12
#263320000000
0!
0%
b110 *
0-
02
b110 6
#263330000000
1!
1%
1-
12
#263340000000
0!
0%
b111 *
0-
02
b111 6
#263350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#263360000000
0!
0%
b0 *
0-
02
b0 6
#263370000000
1!
1%
1-
12
#263380000000
0!
0%
b1 *
0-
02
b1 6
#263390000000
1!
1%
1-
12
#263400000000
0!
0%
b10 *
0-
02
b10 6
#263410000000
1!
1%
1-
12
#263420000000
0!
0%
b11 *
0-
02
b11 6
#263430000000
1!
1%
1-
12
15
#263440000000
0!
0%
b100 *
0-
02
b100 6
#263450000000
1!
1%
1-
12
#263460000000
0!
0%
b101 *
0-
02
b101 6
#263470000000
1!
1%
1-
12
#263480000000
0!
0%
b110 *
0-
02
b110 6
#263490000000
1!
1%
1-
12
#263500000000
0!
0%
b111 *
0-
02
b111 6
#263510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#263520000000
0!
0%
b0 *
0-
02
b0 6
#263530000000
1!
1%
1-
12
#263540000000
0!
0%
b1 *
0-
02
b1 6
#263550000000
1!
1%
1-
12
#263560000000
0!
0%
b10 *
0-
02
b10 6
#263570000000
1!
1%
1-
12
#263580000000
0!
0%
b11 *
0-
02
b11 6
#263590000000
1!
1%
1-
12
15
#263600000000
0!
0%
b100 *
0-
02
b100 6
#263610000000
1!
1%
1-
12
#263620000000
0!
0%
b101 *
0-
02
b101 6
#263630000000
1!
1%
1-
12
#263640000000
0!
0%
b110 *
0-
02
b110 6
#263650000000
1!
1%
1-
12
#263660000000
0!
0%
b111 *
0-
02
b111 6
#263670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#263680000000
0!
0%
b0 *
0-
02
b0 6
#263690000000
1!
1%
1-
12
#263700000000
0!
0%
b1 *
0-
02
b1 6
#263710000000
1!
1%
1-
12
#263720000000
0!
0%
b10 *
0-
02
b10 6
#263730000000
1!
1%
1-
12
#263740000000
0!
0%
b11 *
0-
02
b11 6
#263750000000
1!
1%
1-
12
15
#263760000000
0!
0%
b100 *
0-
02
b100 6
#263770000000
1!
1%
1-
12
#263780000000
0!
0%
b101 *
0-
02
b101 6
#263790000000
1!
1%
1-
12
#263800000000
0!
0%
b110 *
0-
02
b110 6
#263810000000
1!
1%
1-
12
#263820000000
0!
0%
b111 *
0-
02
b111 6
#263830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#263840000000
0!
0%
b0 *
0-
02
b0 6
#263850000000
1!
1%
1-
12
#263860000000
0!
0%
b1 *
0-
02
b1 6
#263870000000
1!
1%
1-
12
#263880000000
0!
0%
b10 *
0-
02
b10 6
#263890000000
1!
1%
1-
12
#263900000000
0!
0%
b11 *
0-
02
b11 6
#263910000000
1!
1%
1-
12
15
#263920000000
0!
0%
b100 *
0-
02
b100 6
#263930000000
1!
1%
1-
12
#263940000000
0!
0%
b101 *
0-
02
b101 6
#263950000000
1!
1%
1-
12
#263960000000
0!
0%
b110 *
0-
02
b110 6
#263970000000
1!
1%
1-
12
#263980000000
0!
0%
b111 *
0-
02
b111 6
#263990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#264000000000
0!
0%
b0 *
0-
02
b0 6
#264010000000
1!
1%
1-
12
#264020000000
0!
0%
b1 *
0-
02
b1 6
#264030000000
1!
1%
1-
12
#264040000000
0!
0%
b10 *
0-
02
b10 6
#264050000000
1!
1%
1-
12
#264060000000
0!
0%
b11 *
0-
02
b11 6
#264070000000
1!
1%
1-
12
15
#264080000000
0!
0%
b100 *
0-
02
b100 6
#264090000000
1!
1%
1-
12
#264100000000
0!
0%
b101 *
0-
02
b101 6
#264110000000
1!
1%
1-
12
#264120000000
0!
0%
b110 *
0-
02
b110 6
#264130000000
1!
1%
1-
12
#264140000000
0!
0%
b111 *
0-
02
b111 6
#264150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#264160000000
0!
0%
b0 *
0-
02
b0 6
#264170000000
1!
1%
1-
12
#264180000000
0!
0%
b1 *
0-
02
b1 6
#264190000000
1!
1%
1-
12
#264200000000
0!
0%
b10 *
0-
02
b10 6
#264210000000
1!
1%
1-
12
#264220000000
0!
0%
b11 *
0-
02
b11 6
#264230000000
1!
1%
1-
12
15
#264240000000
0!
0%
b100 *
0-
02
b100 6
#264250000000
1!
1%
1-
12
#264260000000
0!
0%
b101 *
0-
02
b101 6
#264270000000
1!
1%
1-
12
#264280000000
0!
0%
b110 *
0-
02
b110 6
#264290000000
1!
1%
1-
12
#264300000000
0!
0%
b111 *
0-
02
b111 6
#264310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#264320000000
0!
0%
b0 *
0-
02
b0 6
#264330000000
1!
1%
1-
12
#264340000000
0!
0%
b1 *
0-
02
b1 6
#264350000000
1!
1%
1-
12
#264360000000
0!
0%
b10 *
0-
02
b10 6
#264370000000
1!
1%
1-
12
#264380000000
0!
0%
b11 *
0-
02
b11 6
#264390000000
1!
1%
1-
12
15
#264400000000
0!
0%
b100 *
0-
02
b100 6
#264410000000
1!
1%
1-
12
#264420000000
0!
0%
b101 *
0-
02
b101 6
#264430000000
1!
1%
1-
12
#264440000000
0!
0%
b110 *
0-
02
b110 6
#264450000000
1!
1%
1-
12
#264460000000
0!
0%
b111 *
0-
02
b111 6
#264470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#264480000000
0!
0%
b0 *
0-
02
b0 6
#264490000000
1!
1%
1-
12
#264500000000
0!
0%
b1 *
0-
02
b1 6
#264510000000
1!
1%
1-
12
#264520000000
0!
0%
b10 *
0-
02
b10 6
#264530000000
1!
1%
1-
12
#264540000000
0!
0%
b11 *
0-
02
b11 6
#264550000000
1!
1%
1-
12
15
#264560000000
0!
0%
b100 *
0-
02
b100 6
#264570000000
1!
1%
1-
12
#264580000000
0!
0%
b101 *
0-
02
b101 6
#264590000000
1!
1%
1-
12
#264600000000
0!
0%
b110 *
0-
02
b110 6
#264610000000
1!
1%
1-
12
#264620000000
0!
0%
b111 *
0-
02
b111 6
#264630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#264640000000
0!
0%
b0 *
0-
02
b0 6
#264650000000
1!
1%
1-
12
#264660000000
0!
0%
b1 *
0-
02
b1 6
#264670000000
1!
1%
1-
12
#264680000000
0!
0%
b10 *
0-
02
b10 6
#264690000000
1!
1%
1-
12
#264700000000
0!
0%
b11 *
0-
02
b11 6
#264710000000
1!
1%
1-
12
15
#264720000000
0!
0%
b100 *
0-
02
b100 6
#264730000000
1!
1%
1-
12
#264740000000
0!
0%
b101 *
0-
02
b101 6
#264750000000
1!
1%
1-
12
#264760000000
0!
0%
b110 *
0-
02
b110 6
#264770000000
1!
1%
1-
12
#264780000000
0!
0%
b111 *
0-
02
b111 6
#264790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#264800000000
0!
0%
b0 *
0-
02
b0 6
#264810000000
1!
1%
1-
12
#264820000000
0!
0%
b1 *
0-
02
b1 6
#264830000000
1!
1%
1-
12
#264840000000
0!
0%
b10 *
0-
02
b10 6
#264850000000
1!
1%
1-
12
#264860000000
0!
0%
b11 *
0-
02
b11 6
#264870000000
1!
1%
1-
12
15
#264880000000
0!
0%
b100 *
0-
02
b100 6
#264890000000
1!
1%
1-
12
#264900000000
0!
0%
b101 *
0-
02
b101 6
#264910000000
1!
1%
1-
12
#264920000000
0!
0%
b110 *
0-
02
b110 6
#264930000000
1!
1%
1-
12
#264940000000
0!
0%
b111 *
0-
02
b111 6
#264950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#264960000000
0!
0%
b0 *
0-
02
b0 6
#264970000000
1!
1%
1-
12
#264980000000
0!
0%
b1 *
0-
02
b1 6
#264990000000
1!
1%
1-
12
#265000000000
0!
0%
b10 *
0-
02
b10 6
#265010000000
1!
1%
1-
12
#265020000000
0!
0%
b11 *
0-
02
b11 6
#265030000000
1!
1%
1-
12
15
#265040000000
0!
0%
b100 *
0-
02
b100 6
#265050000000
1!
1%
1-
12
#265060000000
0!
0%
b101 *
0-
02
b101 6
#265070000000
1!
1%
1-
12
#265080000000
0!
0%
b110 *
0-
02
b110 6
#265090000000
1!
1%
1-
12
#265100000000
0!
0%
b111 *
0-
02
b111 6
#265110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#265120000000
0!
0%
b0 *
0-
02
b0 6
#265130000000
1!
1%
1-
12
#265140000000
0!
0%
b1 *
0-
02
b1 6
#265150000000
1!
1%
1-
12
#265160000000
0!
0%
b10 *
0-
02
b10 6
#265170000000
1!
1%
1-
12
#265180000000
0!
0%
b11 *
0-
02
b11 6
#265190000000
1!
1%
1-
12
15
#265200000000
0!
0%
b100 *
0-
02
b100 6
#265210000000
1!
1%
1-
12
#265220000000
0!
0%
b101 *
0-
02
b101 6
#265230000000
1!
1%
1-
12
#265240000000
0!
0%
b110 *
0-
02
b110 6
#265250000000
1!
1%
1-
12
#265260000000
0!
0%
b111 *
0-
02
b111 6
#265270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#265280000000
0!
0%
b0 *
0-
02
b0 6
#265290000000
1!
1%
1-
12
#265300000000
0!
0%
b1 *
0-
02
b1 6
#265310000000
1!
1%
1-
12
#265320000000
0!
0%
b10 *
0-
02
b10 6
#265330000000
1!
1%
1-
12
#265340000000
0!
0%
b11 *
0-
02
b11 6
#265350000000
1!
1%
1-
12
15
#265360000000
0!
0%
b100 *
0-
02
b100 6
#265370000000
1!
1%
1-
12
#265380000000
0!
0%
b101 *
0-
02
b101 6
#265390000000
1!
1%
1-
12
#265400000000
0!
0%
b110 *
0-
02
b110 6
#265410000000
1!
1%
1-
12
#265420000000
0!
0%
b111 *
0-
02
b111 6
#265430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#265440000000
0!
0%
b0 *
0-
02
b0 6
#265450000000
1!
1%
1-
12
#265460000000
0!
0%
b1 *
0-
02
b1 6
#265470000000
1!
1%
1-
12
#265480000000
0!
0%
b10 *
0-
02
b10 6
#265490000000
1!
1%
1-
12
#265500000000
0!
0%
b11 *
0-
02
b11 6
#265510000000
1!
1%
1-
12
15
#265520000000
0!
0%
b100 *
0-
02
b100 6
#265530000000
1!
1%
1-
12
#265540000000
0!
0%
b101 *
0-
02
b101 6
#265550000000
1!
1%
1-
12
#265560000000
0!
0%
b110 *
0-
02
b110 6
#265570000000
1!
1%
1-
12
#265580000000
0!
0%
b111 *
0-
02
b111 6
#265590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#265600000000
0!
0%
b0 *
0-
02
b0 6
#265610000000
1!
1%
1-
12
#265620000000
0!
0%
b1 *
0-
02
b1 6
#265630000000
1!
1%
1-
12
#265640000000
0!
0%
b10 *
0-
02
b10 6
#265650000000
1!
1%
1-
12
#265660000000
0!
0%
b11 *
0-
02
b11 6
#265670000000
1!
1%
1-
12
15
#265680000000
0!
0%
b100 *
0-
02
b100 6
#265690000000
1!
1%
1-
12
#265700000000
0!
0%
b101 *
0-
02
b101 6
#265710000000
1!
1%
1-
12
#265720000000
0!
0%
b110 *
0-
02
b110 6
#265730000000
1!
1%
1-
12
#265740000000
0!
0%
b111 *
0-
02
b111 6
#265750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#265760000000
0!
0%
b0 *
0-
02
b0 6
#265770000000
1!
1%
1-
12
#265780000000
0!
0%
b1 *
0-
02
b1 6
#265790000000
1!
1%
1-
12
#265800000000
0!
0%
b10 *
0-
02
b10 6
#265810000000
1!
1%
1-
12
#265820000000
0!
0%
b11 *
0-
02
b11 6
#265830000000
1!
1%
1-
12
15
#265840000000
0!
0%
b100 *
0-
02
b100 6
#265850000000
1!
1%
1-
12
#265860000000
0!
0%
b101 *
0-
02
b101 6
#265870000000
1!
1%
1-
12
#265880000000
0!
0%
b110 *
0-
02
b110 6
#265890000000
1!
1%
1-
12
#265900000000
0!
0%
b111 *
0-
02
b111 6
#265910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#265920000000
0!
0%
b0 *
0-
02
b0 6
#265930000000
1!
1%
1-
12
#265940000000
0!
0%
b1 *
0-
02
b1 6
#265950000000
1!
1%
1-
12
#265960000000
0!
0%
b10 *
0-
02
b10 6
#265970000000
1!
1%
1-
12
#265980000000
0!
0%
b11 *
0-
02
b11 6
#265990000000
1!
1%
1-
12
15
#266000000000
0!
0%
b100 *
0-
02
b100 6
#266010000000
1!
1%
1-
12
#266020000000
0!
0%
b101 *
0-
02
b101 6
#266030000000
1!
1%
1-
12
#266040000000
0!
0%
b110 *
0-
02
b110 6
#266050000000
1!
1%
1-
12
#266060000000
0!
0%
b111 *
0-
02
b111 6
#266070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#266080000000
0!
0%
b0 *
0-
02
b0 6
#266090000000
1!
1%
1-
12
#266100000000
0!
0%
b1 *
0-
02
b1 6
#266110000000
1!
1%
1-
12
#266120000000
0!
0%
b10 *
0-
02
b10 6
#266130000000
1!
1%
1-
12
#266140000000
0!
0%
b11 *
0-
02
b11 6
#266150000000
1!
1%
1-
12
15
#266160000000
0!
0%
b100 *
0-
02
b100 6
#266170000000
1!
1%
1-
12
#266180000000
0!
0%
b101 *
0-
02
b101 6
#266190000000
1!
1%
1-
12
#266200000000
0!
0%
b110 *
0-
02
b110 6
#266210000000
1!
1%
1-
12
#266220000000
0!
0%
b111 *
0-
02
b111 6
#266230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#266240000000
0!
0%
b0 *
0-
02
b0 6
#266250000000
1!
1%
1-
12
#266260000000
0!
0%
b1 *
0-
02
b1 6
#266270000000
1!
1%
1-
12
#266280000000
0!
0%
b10 *
0-
02
b10 6
#266290000000
1!
1%
1-
12
#266300000000
0!
0%
b11 *
0-
02
b11 6
#266310000000
1!
1%
1-
12
15
#266320000000
0!
0%
b100 *
0-
02
b100 6
#266330000000
1!
1%
1-
12
#266340000000
0!
0%
b101 *
0-
02
b101 6
#266350000000
1!
1%
1-
12
#266360000000
0!
0%
b110 *
0-
02
b110 6
#266370000000
1!
1%
1-
12
#266380000000
0!
0%
b111 *
0-
02
b111 6
#266390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#266400000000
0!
0%
b0 *
0-
02
b0 6
#266410000000
1!
1%
1-
12
#266420000000
0!
0%
b1 *
0-
02
b1 6
#266430000000
1!
1%
1-
12
#266440000000
0!
0%
b10 *
0-
02
b10 6
#266450000000
1!
1%
1-
12
#266460000000
0!
0%
b11 *
0-
02
b11 6
#266470000000
1!
1%
1-
12
15
#266480000000
0!
0%
b100 *
0-
02
b100 6
#266490000000
1!
1%
1-
12
#266500000000
0!
0%
b101 *
0-
02
b101 6
#266510000000
1!
1%
1-
12
#266520000000
0!
0%
b110 *
0-
02
b110 6
#266530000000
1!
1%
1-
12
#266540000000
0!
0%
b111 *
0-
02
b111 6
#266550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#266560000000
0!
0%
b0 *
0-
02
b0 6
#266570000000
1!
1%
1-
12
#266580000000
0!
0%
b1 *
0-
02
b1 6
#266590000000
1!
1%
1-
12
#266600000000
0!
0%
b10 *
0-
02
b10 6
#266610000000
1!
1%
1-
12
#266620000000
0!
0%
b11 *
0-
02
b11 6
#266630000000
1!
1%
1-
12
15
#266640000000
0!
0%
b100 *
0-
02
b100 6
#266650000000
1!
1%
1-
12
#266660000000
0!
0%
b101 *
0-
02
b101 6
#266670000000
1!
1%
1-
12
#266680000000
0!
0%
b110 *
0-
02
b110 6
#266690000000
1!
1%
1-
12
#266700000000
0!
0%
b111 *
0-
02
b111 6
#266710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#266720000000
0!
0%
b0 *
0-
02
b0 6
#266730000000
1!
1%
1-
12
#266740000000
0!
0%
b1 *
0-
02
b1 6
#266750000000
1!
1%
1-
12
#266760000000
0!
0%
b10 *
0-
02
b10 6
#266770000000
1!
1%
1-
12
#266780000000
0!
0%
b11 *
0-
02
b11 6
#266790000000
1!
1%
1-
12
15
#266800000000
0!
0%
b100 *
0-
02
b100 6
#266810000000
1!
1%
1-
12
#266820000000
0!
0%
b101 *
0-
02
b101 6
#266830000000
1!
1%
1-
12
#266840000000
0!
0%
b110 *
0-
02
b110 6
#266850000000
1!
1%
1-
12
#266860000000
0!
0%
b111 *
0-
02
b111 6
#266870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#266880000000
0!
0%
b0 *
0-
02
b0 6
#266890000000
1!
1%
1-
12
#266900000000
0!
0%
b1 *
0-
02
b1 6
#266910000000
1!
1%
1-
12
#266920000000
0!
0%
b10 *
0-
02
b10 6
#266930000000
1!
1%
1-
12
#266940000000
0!
0%
b11 *
0-
02
b11 6
#266950000000
1!
1%
1-
12
15
#266960000000
0!
0%
b100 *
0-
02
b100 6
#266970000000
1!
1%
1-
12
#266980000000
0!
0%
b101 *
0-
02
b101 6
#266990000000
1!
1%
1-
12
#267000000000
0!
0%
b110 *
0-
02
b110 6
#267010000000
1!
1%
1-
12
#267020000000
0!
0%
b111 *
0-
02
b111 6
#267030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#267040000000
0!
0%
b0 *
0-
02
b0 6
#267050000000
1!
1%
1-
12
#267060000000
0!
0%
b1 *
0-
02
b1 6
#267070000000
1!
1%
1-
12
#267080000000
0!
0%
b10 *
0-
02
b10 6
#267090000000
1!
1%
1-
12
#267100000000
0!
0%
b11 *
0-
02
b11 6
#267110000000
1!
1%
1-
12
15
#267120000000
0!
0%
b100 *
0-
02
b100 6
#267130000000
1!
1%
1-
12
#267140000000
0!
0%
b101 *
0-
02
b101 6
#267150000000
1!
1%
1-
12
#267160000000
0!
0%
b110 *
0-
02
b110 6
#267170000000
1!
1%
1-
12
#267180000000
0!
0%
b111 *
0-
02
b111 6
#267190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#267200000000
0!
0%
b0 *
0-
02
b0 6
#267210000000
1!
1%
1-
12
#267220000000
0!
0%
b1 *
0-
02
b1 6
#267230000000
1!
1%
1-
12
#267240000000
0!
0%
b10 *
0-
02
b10 6
#267250000000
1!
1%
1-
12
#267260000000
0!
0%
b11 *
0-
02
b11 6
#267270000000
1!
1%
1-
12
15
#267280000000
0!
0%
b100 *
0-
02
b100 6
#267290000000
1!
1%
1-
12
#267300000000
0!
0%
b101 *
0-
02
b101 6
#267310000000
1!
1%
1-
12
#267320000000
0!
0%
b110 *
0-
02
b110 6
#267330000000
1!
1%
1-
12
#267340000000
0!
0%
b111 *
0-
02
b111 6
#267350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#267360000000
0!
0%
b0 *
0-
02
b0 6
#267370000000
1!
1%
1-
12
#267380000000
0!
0%
b1 *
0-
02
b1 6
#267390000000
1!
1%
1-
12
#267400000000
0!
0%
b10 *
0-
02
b10 6
#267410000000
1!
1%
1-
12
#267420000000
0!
0%
b11 *
0-
02
b11 6
#267430000000
1!
1%
1-
12
15
#267440000000
0!
0%
b100 *
0-
02
b100 6
#267450000000
1!
1%
1-
12
#267460000000
0!
0%
b101 *
0-
02
b101 6
#267470000000
1!
1%
1-
12
#267480000000
0!
0%
b110 *
0-
02
b110 6
#267490000000
1!
1%
1-
12
#267500000000
0!
0%
b111 *
0-
02
b111 6
#267510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#267520000000
0!
0%
b0 *
0-
02
b0 6
#267530000000
1!
1%
1-
12
#267540000000
0!
0%
b1 *
0-
02
b1 6
#267550000000
1!
1%
1-
12
#267560000000
0!
0%
b10 *
0-
02
b10 6
#267570000000
1!
1%
1-
12
#267580000000
0!
0%
b11 *
0-
02
b11 6
#267590000000
1!
1%
1-
12
15
#267600000000
0!
0%
b100 *
0-
02
b100 6
#267610000000
1!
1%
1-
12
#267620000000
0!
0%
b101 *
0-
02
b101 6
#267630000000
1!
1%
1-
12
#267640000000
0!
0%
b110 *
0-
02
b110 6
#267650000000
1!
1%
1-
12
#267660000000
0!
0%
b111 *
0-
02
b111 6
#267670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#267680000000
0!
0%
b0 *
0-
02
b0 6
#267690000000
1!
1%
1-
12
#267700000000
0!
0%
b1 *
0-
02
b1 6
#267710000000
1!
1%
1-
12
#267720000000
0!
0%
b10 *
0-
02
b10 6
#267730000000
1!
1%
1-
12
#267740000000
0!
0%
b11 *
0-
02
b11 6
#267750000000
1!
1%
1-
12
15
#267760000000
0!
0%
b100 *
0-
02
b100 6
#267770000000
1!
1%
1-
12
#267780000000
0!
0%
b101 *
0-
02
b101 6
#267790000000
1!
1%
1-
12
#267800000000
0!
0%
b110 *
0-
02
b110 6
#267810000000
1!
1%
1-
12
#267820000000
0!
0%
b111 *
0-
02
b111 6
#267830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#267840000000
0!
0%
b0 *
0-
02
b0 6
#267850000000
1!
1%
1-
12
#267860000000
0!
0%
b1 *
0-
02
b1 6
#267870000000
1!
1%
1-
12
#267880000000
0!
0%
b10 *
0-
02
b10 6
#267890000000
1!
1%
1-
12
#267900000000
0!
0%
b11 *
0-
02
b11 6
#267910000000
1!
1%
1-
12
15
#267920000000
0!
0%
b100 *
0-
02
b100 6
#267930000000
1!
1%
1-
12
#267940000000
0!
0%
b101 *
0-
02
b101 6
#267950000000
1!
1%
1-
12
#267960000000
0!
0%
b110 *
0-
02
b110 6
#267970000000
1!
1%
1-
12
#267980000000
0!
0%
b111 *
0-
02
b111 6
#267990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#268000000000
0!
0%
b0 *
0-
02
b0 6
#268010000000
1!
1%
1-
12
#268020000000
0!
0%
b1 *
0-
02
b1 6
#268030000000
1!
1%
1-
12
#268040000000
0!
0%
b10 *
0-
02
b10 6
#268050000000
1!
1%
1-
12
#268060000000
0!
0%
b11 *
0-
02
b11 6
#268070000000
1!
1%
1-
12
15
#268080000000
0!
0%
b100 *
0-
02
b100 6
#268090000000
1!
1%
1-
12
#268100000000
0!
0%
b101 *
0-
02
b101 6
#268110000000
1!
1%
1-
12
#268120000000
0!
0%
b110 *
0-
02
b110 6
#268130000000
1!
1%
1-
12
#268140000000
0!
0%
b111 *
0-
02
b111 6
#268150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#268160000000
0!
0%
b0 *
0-
02
b0 6
#268170000000
1!
1%
1-
12
#268180000000
0!
0%
b1 *
0-
02
b1 6
#268190000000
1!
1%
1-
12
#268200000000
0!
0%
b10 *
0-
02
b10 6
#268210000000
1!
1%
1-
12
#268220000000
0!
0%
b11 *
0-
02
b11 6
#268230000000
1!
1%
1-
12
15
#268240000000
0!
0%
b100 *
0-
02
b100 6
#268250000000
1!
1%
1-
12
#268260000000
0!
0%
b101 *
0-
02
b101 6
#268270000000
1!
1%
1-
12
#268280000000
0!
0%
b110 *
0-
02
b110 6
#268290000000
1!
1%
1-
12
#268300000000
0!
0%
b111 *
0-
02
b111 6
#268310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#268320000000
0!
0%
b0 *
0-
02
b0 6
#268330000000
1!
1%
1-
12
#268340000000
0!
0%
b1 *
0-
02
b1 6
#268350000000
1!
1%
1-
12
#268360000000
0!
0%
b10 *
0-
02
b10 6
#268370000000
1!
1%
1-
12
#268380000000
0!
0%
b11 *
0-
02
b11 6
#268390000000
1!
1%
1-
12
15
#268400000000
0!
0%
b100 *
0-
02
b100 6
#268410000000
1!
1%
1-
12
#268420000000
0!
0%
b101 *
0-
02
b101 6
#268430000000
1!
1%
1-
12
#268440000000
0!
0%
b110 *
0-
02
b110 6
#268450000000
1!
1%
1-
12
#268460000000
0!
0%
b111 *
0-
02
b111 6
#268470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#268480000000
0!
0%
b0 *
0-
02
b0 6
#268490000000
1!
1%
1-
12
#268500000000
0!
0%
b1 *
0-
02
b1 6
#268510000000
1!
1%
1-
12
#268520000000
0!
0%
b10 *
0-
02
b10 6
#268530000000
1!
1%
1-
12
#268540000000
0!
0%
b11 *
0-
02
b11 6
#268550000000
1!
1%
1-
12
15
#268560000000
0!
0%
b100 *
0-
02
b100 6
#268570000000
1!
1%
1-
12
#268580000000
0!
0%
b101 *
0-
02
b101 6
#268590000000
1!
1%
1-
12
#268600000000
0!
0%
b110 *
0-
02
b110 6
#268610000000
1!
1%
1-
12
#268620000000
0!
0%
b111 *
0-
02
b111 6
#268630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#268640000000
0!
0%
b0 *
0-
02
b0 6
#268650000000
1!
1%
1-
12
#268660000000
0!
0%
b1 *
0-
02
b1 6
#268670000000
1!
1%
1-
12
#268680000000
0!
0%
b10 *
0-
02
b10 6
#268690000000
1!
1%
1-
12
#268700000000
0!
0%
b11 *
0-
02
b11 6
#268710000000
1!
1%
1-
12
15
#268720000000
0!
0%
b100 *
0-
02
b100 6
#268730000000
1!
1%
1-
12
#268740000000
0!
0%
b101 *
0-
02
b101 6
#268750000000
1!
1%
1-
12
#268760000000
0!
0%
b110 *
0-
02
b110 6
#268770000000
1!
1%
1-
12
#268780000000
0!
0%
b111 *
0-
02
b111 6
#268790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#268800000000
0!
0%
b0 *
0-
02
b0 6
#268810000000
1!
1%
1-
12
#268820000000
0!
0%
b1 *
0-
02
b1 6
#268830000000
1!
1%
1-
12
#268840000000
0!
0%
b10 *
0-
02
b10 6
#268850000000
1!
1%
1-
12
#268860000000
0!
0%
b11 *
0-
02
b11 6
#268870000000
1!
1%
1-
12
15
#268880000000
0!
0%
b100 *
0-
02
b100 6
#268890000000
1!
1%
1-
12
#268900000000
0!
0%
b101 *
0-
02
b101 6
#268910000000
1!
1%
1-
12
#268920000000
0!
0%
b110 *
0-
02
b110 6
#268930000000
1!
1%
1-
12
#268940000000
0!
0%
b111 *
0-
02
b111 6
#268950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#268960000000
0!
0%
b0 *
0-
02
b0 6
#268970000000
1!
1%
1-
12
#268980000000
0!
0%
b1 *
0-
02
b1 6
#268990000000
1!
1%
1-
12
#269000000000
0!
0%
b10 *
0-
02
b10 6
#269010000000
1!
1%
1-
12
#269020000000
0!
0%
b11 *
0-
02
b11 6
#269030000000
1!
1%
1-
12
15
#269040000000
0!
0%
b100 *
0-
02
b100 6
#269050000000
1!
1%
1-
12
#269060000000
0!
0%
b101 *
0-
02
b101 6
#269070000000
1!
1%
1-
12
#269080000000
0!
0%
b110 *
0-
02
b110 6
#269090000000
1!
1%
1-
12
#269100000000
0!
0%
b111 *
0-
02
b111 6
#269110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#269120000000
0!
0%
b0 *
0-
02
b0 6
#269130000000
1!
1%
1-
12
#269140000000
0!
0%
b1 *
0-
02
b1 6
#269150000000
1!
1%
1-
12
#269160000000
0!
0%
b10 *
0-
02
b10 6
#269170000000
1!
1%
1-
12
#269180000000
0!
0%
b11 *
0-
02
b11 6
#269190000000
1!
1%
1-
12
15
#269200000000
0!
0%
b100 *
0-
02
b100 6
#269210000000
1!
1%
1-
12
#269220000000
0!
0%
b101 *
0-
02
b101 6
#269230000000
1!
1%
1-
12
#269240000000
0!
0%
b110 *
0-
02
b110 6
#269250000000
1!
1%
1-
12
#269260000000
0!
0%
b111 *
0-
02
b111 6
#269270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#269280000000
0!
0%
b0 *
0-
02
b0 6
#269290000000
1!
1%
1-
12
#269300000000
0!
0%
b1 *
0-
02
b1 6
#269310000000
1!
1%
1-
12
#269320000000
0!
0%
b10 *
0-
02
b10 6
#269330000000
1!
1%
1-
12
#269340000000
0!
0%
b11 *
0-
02
b11 6
#269350000000
1!
1%
1-
12
15
#269360000000
0!
0%
b100 *
0-
02
b100 6
#269370000000
1!
1%
1-
12
#269380000000
0!
0%
b101 *
0-
02
b101 6
#269390000000
1!
1%
1-
12
#269400000000
0!
0%
b110 *
0-
02
b110 6
#269410000000
1!
1%
1-
12
#269420000000
0!
0%
b111 *
0-
02
b111 6
#269430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#269440000000
0!
0%
b0 *
0-
02
b0 6
#269450000000
1!
1%
1-
12
#269460000000
0!
0%
b1 *
0-
02
b1 6
#269470000000
1!
1%
1-
12
#269480000000
0!
0%
b10 *
0-
02
b10 6
#269490000000
1!
1%
1-
12
#269500000000
0!
0%
b11 *
0-
02
b11 6
#269510000000
1!
1%
1-
12
15
#269520000000
0!
0%
b100 *
0-
02
b100 6
#269530000000
1!
1%
1-
12
#269540000000
0!
0%
b101 *
0-
02
b101 6
#269550000000
1!
1%
1-
12
#269560000000
0!
0%
b110 *
0-
02
b110 6
#269570000000
1!
1%
1-
12
#269580000000
0!
0%
b111 *
0-
02
b111 6
#269590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#269600000000
0!
0%
b0 *
0-
02
b0 6
#269610000000
1!
1%
1-
12
#269620000000
0!
0%
b1 *
0-
02
b1 6
#269630000000
1!
1%
1-
12
#269640000000
0!
0%
b10 *
0-
02
b10 6
#269650000000
1!
1%
1-
12
#269660000000
0!
0%
b11 *
0-
02
b11 6
#269670000000
1!
1%
1-
12
15
#269680000000
0!
0%
b100 *
0-
02
b100 6
#269690000000
1!
1%
1-
12
#269700000000
0!
0%
b101 *
0-
02
b101 6
#269710000000
1!
1%
1-
12
#269720000000
0!
0%
b110 *
0-
02
b110 6
#269730000000
1!
1%
1-
12
#269740000000
0!
0%
b111 *
0-
02
b111 6
#269750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#269760000000
0!
0%
b0 *
0-
02
b0 6
#269770000000
1!
1%
1-
12
#269780000000
0!
0%
b1 *
0-
02
b1 6
#269790000000
1!
1%
1-
12
#269800000000
0!
0%
b10 *
0-
02
b10 6
#269810000000
1!
1%
1-
12
#269820000000
0!
0%
b11 *
0-
02
b11 6
#269830000000
1!
1%
1-
12
15
#269840000000
0!
0%
b100 *
0-
02
b100 6
#269850000000
1!
1%
1-
12
#269860000000
0!
0%
b101 *
0-
02
b101 6
#269870000000
1!
1%
1-
12
#269880000000
0!
0%
b110 *
0-
02
b110 6
#269890000000
1!
1%
1-
12
#269900000000
0!
0%
b111 *
0-
02
b111 6
#269910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#269920000000
0!
0%
b0 *
0-
02
b0 6
#269930000000
1!
1%
1-
12
#269940000000
0!
0%
b1 *
0-
02
b1 6
#269950000000
1!
1%
1-
12
#269960000000
0!
0%
b10 *
0-
02
b10 6
#269970000000
1!
1%
1-
12
#269980000000
0!
0%
b11 *
0-
02
b11 6
#269990000000
1!
1%
1-
12
15
#270000000000
0!
0%
b100 *
0-
02
b100 6
#270010000000
1!
1%
1-
12
#270020000000
0!
0%
b101 *
0-
02
b101 6
#270030000000
1!
1%
1-
12
#270040000000
0!
0%
b110 *
0-
02
b110 6
#270050000000
1!
1%
1-
12
#270060000000
0!
0%
b111 *
0-
02
b111 6
#270070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#270080000000
0!
0%
b0 *
0-
02
b0 6
#270090000000
1!
1%
1-
12
#270100000000
0!
0%
b1 *
0-
02
b1 6
#270110000000
1!
1%
1-
12
#270120000000
0!
0%
b10 *
0-
02
b10 6
#270130000000
1!
1%
1-
12
#270140000000
0!
0%
b11 *
0-
02
b11 6
#270150000000
1!
1%
1-
12
15
#270160000000
0!
0%
b100 *
0-
02
b100 6
#270170000000
1!
1%
1-
12
#270180000000
0!
0%
b101 *
0-
02
b101 6
#270190000000
1!
1%
1-
12
#270200000000
0!
0%
b110 *
0-
02
b110 6
#270210000000
1!
1%
1-
12
#270220000000
0!
0%
b111 *
0-
02
b111 6
#270230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#270240000000
0!
0%
b0 *
0-
02
b0 6
#270250000000
1!
1%
1-
12
#270260000000
0!
0%
b1 *
0-
02
b1 6
#270270000000
1!
1%
1-
12
#270280000000
0!
0%
b10 *
0-
02
b10 6
#270290000000
1!
1%
1-
12
#270300000000
0!
0%
b11 *
0-
02
b11 6
#270310000000
1!
1%
1-
12
15
#270320000000
0!
0%
b100 *
0-
02
b100 6
#270330000000
1!
1%
1-
12
#270340000000
0!
0%
b101 *
0-
02
b101 6
#270350000000
1!
1%
1-
12
#270360000000
0!
0%
b110 *
0-
02
b110 6
#270370000000
1!
1%
1-
12
#270380000000
0!
0%
b111 *
0-
02
b111 6
#270390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#270400000000
0!
0%
b0 *
0-
02
b0 6
#270410000000
1!
1%
1-
12
#270420000000
0!
0%
b1 *
0-
02
b1 6
#270430000000
1!
1%
1-
12
#270440000000
0!
0%
b10 *
0-
02
b10 6
#270450000000
1!
1%
1-
12
#270460000000
0!
0%
b11 *
0-
02
b11 6
#270470000000
1!
1%
1-
12
15
#270480000000
0!
0%
b100 *
0-
02
b100 6
#270490000000
1!
1%
1-
12
#270500000000
0!
0%
b101 *
0-
02
b101 6
#270510000000
1!
1%
1-
12
#270520000000
0!
0%
b110 *
0-
02
b110 6
#270530000000
1!
1%
1-
12
#270540000000
0!
0%
b111 *
0-
02
b111 6
#270550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#270560000000
0!
0%
b0 *
0-
02
b0 6
#270570000000
1!
1%
1-
12
#270580000000
0!
0%
b1 *
0-
02
b1 6
#270590000000
1!
1%
1-
12
#270600000000
0!
0%
b10 *
0-
02
b10 6
#270610000000
1!
1%
1-
12
#270620000000
0!
0%
b11 *
0-
02
b11 6
#270630000000
1!
1%
1-
12
15
#270640000000
0!
0%
b100 *
0-
02
b100 6
#270650000000
1!
1%
1-
12
#270660000000
0!
0%
b101 *
0-
02
b101 6
#270670000000
1!
1%
1-
12
#270680000000
0!
0%
b110 *
0-
02
b110 6
#270690000000
1!
1%
1-
12
#270700000000
0!
0%
b111 *
0-
02
b111 6
#270710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#270720000000
0!
0%
b0 *
0-
02
b0 6
#270730000000
1!
1%
1-
12
#270740000000
0!
0%
b1 *
0-
02
b1 6
#270750000000
1!
1%
1-
12
#270760000000
0!
0%
b10 *
0-
02
b10 6
#270770000000
1!
1%
1-
12
#270780000000
0!
0%
b11 *
0-
02
b11 6
#270790000000
1!
1%
1-
12
15
#270800000000
0!
0%
b100 *
0-
02
b100 6
#270810000000
1!
1%
1-
12
#270820000000
0!
0%
b101 *
0-
02
b101 6
#270830000000
1!
1%
1-
12
#270840000000
0!
0%
b110 *
0-
02
b110 6
#270850000000
1!
1%
1-
12
#270860000000
0!
0%
b111 *
0-
02
b111 6
#270870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#270880000000
0!
0%
b0 *
0-
02
b0 6
#270890000000
1!
1%
1-
12
#270900000000
0!
0%
b1 *
0-
02
b1 6
#270910000000
1!
1%
1-
12
#270920000000
0!
0%
b10 *
0-
02
b10 6
#270930000000
1!
1%
1-
12
#270940000000
0!
0%
b11 *
0-
02
b11 6
#270950000000
1!
1%
1-
12
15
#270960000000
0!
0%
b100 *
0-
02
b100 6
#270970000000
1!
1%
1-
12
#270980000000
0!
0%
b101 *
0-
02
b101 6
#270990000000
1!
1%
1-
12
#271000000000
0!
0%
b110 *
0-
02
b110 6
#271010000000
1!
1%
1-
12
#271020000000
0!
0%
b111 *
0-
02
b111 6
#271030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#271040000000
0!
0%
b0 *
0-
02
b0 6
#271050000000
1!
1%
1-
12
#271060000000
0!
0%
b1 *
0-
02
b1 6
#271070000000
1!
1%
1-
12
#271080000000
0!
0%
b10 *
0-
02
b10 6
#271090000000
1!
1%
1-
12
#271100000000
0!
0%
b11 *
0-
02
b11 6
#271110000000
1!
1%
1-
12
15
#271120000000
0!
0%
b100 *
0-
02
b100 6
#271130000000
1!
1%
1-
12
#271140000000
0!
0%
b101 *
0-
02
b101 6
#271150000000
1!
1%
1-
12
#271160000000
0!
0%
b110 *
0-
02
b110 6
#271170000000
1!
1%
1-
12
#271180000000
0!
0%
b111 *
0-
02
b111 6
#271190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#271200000000
0!
0%
b0 *
0-
02
b0 6
#271210000000
1!
1%
1-
12
#271220000000
0!
0%
b1 *
0-
02
b1 6
#271230000000
1!
1%
1-
12
#271240000000
0!
0%
b10 *
0-
02
b10 6
#271250000000
1!
1%
1-
12
#271260000000
0!
0%
b11 *
0-
02
b11 6
#271270000000
1!
1%
1-
12
15
#271280000000
0!
0%
b100 *
0-
02
b100 6
#271290000000
1!
1%
1-
12
#271300000000
0!
0%
b101 *
0-
02
b101 6
#271310000000
1!
1%
1-
12
#271320000000
0!
0%
b110 *
0-
02
b110 6
#271330000000
1!
1%
1-
12
#271340000000
0!
0%
b111 *
0-
02
b111 6
#271350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#271360000000
0!
0%
b0 *
0-
02
b0 6
#271370000000
1!
1%
1-
12
#271380000000
0!
0%
b1 *
0-
02
b1 6
#271390000000
1!
1%
1-
12
#271400000000
0!
0%
b10 *
0-
02
b10 6
#271410000000
1!
1%
1-
12
#271420000000
0!
0%
b11 *
0-
02
b11 6
#271430000000
1!
1%
1-
12
15
#271440000000
0!
0%
b100 *
0-
02
b100 6
#271450000000
1!
1%
1-
12
#271460000000
0!
0%
b101 *
0-
02
b101 6
#271470000000
1!
1%
1-
12
#271480000000
0!
0%
b110 *
0-
02
b110 6
#271490000000
1!
1%
1-
12
#271500000000
0!
0%
b111 *
0-
02
b111 6
#271510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#271520000000
0!
0%
b0 *
0-
02
b0 6
#271530000000
1!
1%
1-
12
#271540000000
0!
0%
b1 *
0-
02
b1 6
#271550000000
1!
1%
1-
12
#271560000000
0!
0%
b10 *
0-
02
b10 6
#271570000000
1!
1%
1-
12
#271580000000
0!
0%
b11 *
0-
02
b11 6
#271590000000
1!
1%
1-
12
15
#271600000000
0!
0%
b100 *
0-
02
b100 6
#271610000000
1!
1%
1-
12
#271620000000
0!
0%
b101 *
0-
02
b101 6
#271630000000
1!
1%
1-
12
#271640000000
0!
0%
b110 *
0-
02
b110 6
#271650000000
1!
1%
1-
12
#271660000000
0!
0%
b111 *
0-
02
b111 6
#271670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#271680000000
0!
0%
b0 *
0-
02
b0 6
#271690000000
1!
1%
1-
12
#271700000000
0!
0%
b1 *
0-
02
b1 6
#271710000000
1!
1%
1-
12
#271720000000
0!
0%
b10 *
0-
02
b10 6
#271730000000
1!
1%
1-
12
#271740000000
0!
0%
b11 *
0-
02
b11 6
#271750000000
1!
1%
1-
12
15
#271760000000
0!
0%
b100 *
0-
02
b100 6
#271770000000
1!
1%
1-
12
#271780000000
0!
0%
b101 *
0-
02
b101 6
#271790000000
1!
1%
1-
12
#271800000000
0!
0%
b110 *
0-
02
b110 6
#271810000000
1!
1%
1-
12
#271820000000
0!
0%
b111 *
0-
02
b111 6
#271830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#271840000000
0!
0%
b0 *
0-
02
b0 6
#271850000000
1!
1%
1-
12
#271860000000
0!
0%
b1 *
0-
02
b1 6
#271870000000
1!
1%
1-
12
#271880000000
0!
0%
b10 *
0-
02
b10 6
#271890000000
1!
1%
1-
12
#271900000000
0!
0%
b11 *
0-
02
b11 6
#271910000000
1!
1%
1-
12
15
#271920000000
0!
0%
b100 *
0-
02
b100 6
#271930000000
1!
1%
1-
12
#271940000000
0!
0%
b101 *
0-
02
b101 6
#271950000000
1!
1%
1-
12
#271960000000
0!
0%
b110 *
0-
02
b110 6
#271970000000
1!
1%
1-
12
#271980000000
0!
0%
b111 *
0-
02
b111 6
#271990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#272000000000
0!
0%
b0 *
0-
02
b0 6
#272010000000
1!
1%
1-
12
#272020000000
0!
0%
b1 *
0-
02
b1 6
#272030000000
1!
1%
1-
12
#272040000000
0!
0%
b10 *
0-
02
b10 6
#272050000000
1!
1%
1-
12
#272060000000
0!
0%
b11 *
0-
02
b11 6
#272070000000
1!
1%
1-
12
15
#272080000000
0!
0%
b100 *
0-
02
b100 6
#272090000000
1!
1%
1-
12
#272100000000
0!
0%
b101 *
0-
02
b101 6
#272110000000
1!
1%
1-
12
#272120000000
0!
0%
b110 *
0-
02
b110 6
#272130000000
1!
1%
1-
12
#272140000000
0!
0%
b111 *
0-
02
b111 6
#272150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#272160000000
0!
0%
b0 *
0-
02
b0 6
#272170000000
1!
1%
1-
12
#272180000000
0!
0%
b1 *
0-
02
b1 6
#272190000000
1!
1%
1-
12
#272200000000
0!
0%
b10 *
0-
02
b10 6
#272210000000
1!
1%
1-
12
#272220000000
0!
0%
b11 *
0-
02
b11 6
#272230000000
1!
1%
1-
12
15
#272240000000
0!
0%
b100 *
0-
02
b100 6
#272250000000
1!
1%
1-
12
#272260000000
0!
0%
b101 *
0-
02
b101 6
#272270000000
1!
1%
1-
12
#272280000000
0!
0%
b110 *
0-
02
b110 6
#272290000000
1!
1%
1-
12
#272300000000
0!
0%
b111 *
0-
02
b111 6
#272310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#272320000000
0!
0%
b0 *
0-
02
b0 6
#272330000000
1!
1%
1-
12
#272340000000
0!
0%
b1 *
0-
02
b1 6
#272350000000
1!
1%
1-
12
#272360000000
0!
0%
b10 *
0-
02
b10 6
#272370000000
1!
1%
1-
12
#272380000000
0!
0%
b11 *
0-
02
b11 6
#272390000000
1!
1%
1-
12
15
#272400000000
0!
0%
b100 *
0-
02
b100 6
#272410000000
1!
1%
1-
12
#272420000000
0!
0%
b101 *
0-
02
b101 6
#272430000000
1!
1%
1-
12
#272440000000
0!
0%
b110 *
0-
02
b110 6
#272450000000
1!
1%
1-
12
#272460000000
0!
0%
b111 *
0-
02
b111 6
#272470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#272480000000
0!
0%
b0 *
0-
02
b0 6
#272490000000
1!
1%
1-
12
#272500000000
0!
0%
b1 *
0-
02
b1 6
#272510000000
1!
1%
1-
12
#272520000000
0!
0%
b10 *
0-
02
b10 6
#272530000000
1!
1%
1-
12
#272540000000
0!
0%
b11 *
0-
02
b11 6
#272550000000
1!
1%
1-
12
15
#272560000000
0!
0%
b100 *
0-
02
b100 6
#272570000000
1!
1%
1-
12
#272580000000
0!
0%
b101 *
0-
02
b101 6
#272590000000
1!
1%
1-
12
#272600000000
0!
0%
b110 *
0-
02
b110 6
#272610000000
1!
1%
1-
12
#272620000000
0!
0%
b111 *
0-
02
b111 6
#272630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#272640000000
0!
0%
b0 *
0-
02
b0 6
#272650000000
1!
1%
1-
12
#272660000000
0!
0%
b1 *
0-
02
b1 6
#272670000000
1!
1%
1-
12
#272680000000
0!
0%
b10 *
0-
02
b10 6
#272690000000
1!
1%
1-
12
#272700000000
0!
0%
b11 *
0-
02
b11 6
#272710000000
1!
1%
1-
12
15
#272720000000
0!
0%
b100 *
0-
02
b100 6
#272730000000
1!
1%
1-
12
#272740000000
0!
0%
b101 *
0-
02
b101 6
#272750000000
1!
1%
1-
12
#272760000000
0!
0%
b110 *
0-
02
b110 6
#272770000000
1!
1%
1-
12
#272780000000
0!
0%
b111 *
0-
02
b111 6
#272790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#272800000000
0!
0%
b0 *
0-
02
b0 6
#272810000000
1!
1%
1-
12
#272820000000
0!
0%
b1 *
0-
02
b1 6
#272830000000
1!
1%
1-
12
#272840000000
0!
0%
b10 *
0-
02
b10 6
#272850000000
1!
1%
1-
12
#272860000000
0!
0%
b11 *
0-
02
b11 6
#272870000000
1!
1%
1-
12
15
#272880000000
0!
0%
b100 *
0-
02
b100 6
#272890000000
1!
1%
1-
12
#272900000000
0!
0%
b101 *
0-
02
b101 6
#272910000000
1!
1%
1-
12
#272920000000
0!
0%
b110 *
0-
02
b110 6
#272930000000
1!
1%
1-
12
#272940000000
0!
0%
b111 *
0-
02
b111 6
#272950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#272960000000
0!
0%
b0 *
0-
02
b0 6
#272970000000
1!
1%
1-
12
#272980000000
0!
0%
b1 *
0-
02
b1 6
#272990000000
1!
1%
1-
12
#273000000000
0!
0%
b10 *
0-
02
b10 6
#273010000000
1!
1%
1-
12
#273020000000
0!
0%
b11 *
0-
02
b11 6
#273030000000
1!
1%
1-
12
15
#273040000000
0!
0%
b100 *
0-
02
b100 6
#273050000000
1!
1%
1-
12
#273060000000
0!
0%
b101 *
0-
02
b101 6
#273070000000
1!
1%
1-
12
#273080000000
0!
0%
b110 *
0-
02
b110 6
#273090000000
1!
1%
1-
12
#273100000000
0!
0%
b111 *
0-
02
b111 6
#273110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#273120000000
0!
0%
b0 *
0-
02
b0 6
#273130000000
1!
1%
1-
12
#273140000000
0!
0%
b1 *
0-
02
b1 6
#273150000000
1!
1%
1-
12
#273160000000
0!
0%
b10 *
0-
02
b10 6
#273170000000
1!
1%
1-
12
#273180000000
0!
0%
b11 *
0-
02
b11 6
#273190000000
1!
1%
1-
12
15
#273200000000
0!
0%
b100 *
0-
02
b100 6
#273210000000
1!
1%
1-
12
#273220000000
0!
0%
b101 *
0-
02
b101 6
#273230000000
1!
1%
1-
12
#273240000000
0!
0%
b110 *
0-
02
b110 6
#273250000000
1!
1%
1-
12
#273260000000
0!
0%
b111 *
0-
02
b111 6
#273270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#273280000000
0!
0%
b0 *
0-
02
b0 6
#273290000000
1!
1%
1-
12
#273300000000
0!
0%
b1 *
0-
02
b1 6
#273310000000
1!
1%
1-
12
#273320000000
0!
0%
b10 *
0-
02
b10 6
#273330000000
1!
1%
1-
12
#273340000000
0!
0%
b11 *
0-
02
b11 6
#273350000000
1!
1%
1-
12
15
#273360000000
0!
0%
b100 *
0-
02
b100 6
#273370000000
1!
1%
1-
12
#273380000000
0!
0%
b101 *
0-
02
b101 6
#273390000000
1!
1%
1-
12
#273400000000
0!
0%
b110 *
0-
02
b110 6
#273410000000
1!
1%
1-
12
#273420000000
0!
0%
b111 *
0-
02
b111 6
#273430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#273440000000
0!
0%
b0 *
0-
02
b0 6
#273450000000
1!
1%
1-
12
#273460000000
0!
0%
b1 *
0-
02
b1 6
#273470000000
1!
1%
1-
12
#273480000000
0!
0%
b10 *
0-
02
b10 6
#273490000000
1!
1%
1-
12
#273500000000
0!
0%
b11 *
0-
02
b11 6
#273510000000
1!
1%
1-
12
15
#273520000000
0!
0%
b100 *
0-
02
b100 6
#273530000000
1!
1%
1-
12
#273540000000
0!
0%
b101 *
0-
02
b101 6
#273550000000
1!
1%
1-
12
#273560000000
0!
0%
b110 *
0-
02
b110 6
#273570000000
1!
1%
1-
12
#273580000000
0!
0%
b111 *
0-
02
b111 6
#273590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#273600000000
0!
0%
b0 *
0-
02
b0 6
#273610000000
1!
1%
1-
12
#273620000000
0!
0%
b1 *
0-
02
b1 6
#273630000000
1!
1%
1-
12
#273640000000
0!
0%
b10 *
0-
02
b10 6
#273650000000
1!
1%
1-
12
#273660000000
0!
0%
b11 *
0-
02
b11 6
#273670000000
1!
1%
1-
12
15
#273680000000
0!
0%
b100 *
0-
02
b100 6
#273690000000
1!
1%
1-
12
#273700000000
0!
0%
b101 *
0-
02
b101 6
#273710000000
1!
1%
1-
12
#273720000000
0!
0%
b110 *
0-
02
b110 6
#273730000000
1!
1%
1-
12
#273740000000
0!
0%
b111 *
0-
02
b111 6
#273750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#273760000000
0!
0%
b0 *
0-
02
b0 6
#273770000000
1!
1%
1-
12
#273780000000
0!
0%
b1 *
0-
02
b1 6
#273790000000
1!
1%
1-
12
#273800000000
0!
0%
b10 *
0-
02
b10 6
#273810000000
1!
1%
1-
12
#273820000000
0!
0%
b11 *
0-
02
b11 6
#273830000000
1!
1%
1-
12
15
#273840000000
0!
0%
b100 *
0-
02
b100 6
#273850000000
1!
1%
1-
12
#273860000000
0!
0%
b101 *
0-
02
b101 6
#273870000000
1!
1%
1-
12
#273880000000
0!
0%
b110 *
0-
02
b110 6
#273890000000
1!
1%
1-
12
#273900000000
0!
0%
b111 *
0-
02
b111 6
#273910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#273920000000
0!
0%
b0 *
0-
02
b0 6
#273930000000
1!
1%
1-
12
#273940000000
0!
0%
b1 *
0-
02
b1 6
#273950000000
1!
1%
1-
12
#273960000000
0!
0%
b10 *
0-
02
b10 6
#273970000000
1!
1%
1-
12
#273980000000
0!
0%
b11 *
0-
02
b11 6
#273990000000
1!
1%
1-
12
15
#274000000000
0!
0%
b100 *
0-
02
b100 6
#274010000000
1!
1%
1-
12
#274020000000
0!
0%
b101 *
0-
02
b101 6
#274030000000
1!
1%
1-
12
#274040000000
0!
0%
b110 *
0-
02
b110 6
#274050000000
1!
1%
1-
12
#274060000000
0!
0%
b111 *
0-
02
b111 6
#274070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#274080000000
0!
0%
b0 *
0-
02
b0 6
#274090000000
1!
1%
1-
12
#274100000000
0!
0%
b1 *
0-
02
b1 6
#274110000000
1!
1%
1-
12
#274120000000
0!
0%
b10 *
0-
02
b10 6
#274130000000
1!
1%
1-
12
#274140000000
0!
0%
b11 *
0-
02
b11 6
#274150000000
1!
1%
1-
12
15
#274160000000
0!
0%
b100 *
0-
02
b100 6
#274170000000
1!
1%
1-
12
#274180000000
0!
0%
b101 *
0-
02
b101 6
#274190000000
1!
1%
1-
12
#274200000000
0!
0%
b110 *
0-
02
b110 6
#274210000000
1!
1%
1-
12
#274220000000
0!
0%
b111 *
0-
02
b111 6
#274230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#274240000000
0!
0%
b0 *
0-
02
b0 6
#274250000000
1!
1%
1-
12
#274260000000
0!
0%
b1 *
0-
02
b1 6
#274270000000
1!
1%
1-
12
#274280000000
0!
0%
b10 *
0-
02
b10 6
#274290000000
1!
1%
1-
12
#274300000000
0!
0%
b11 *
0-
02
b11 6
#274310000000
1!
1%
1-
12
15
#274320000000
0!
0%
b100 *
0-
02
b100 6
#274330000000
1!
1%
1-
12
#274340000000
0!
0%
b101 *
0-
02
b101 6
#274350000000
1!
1%
1-
12
#274360000000
0!
0%
b110 *
0-
02
b110 6
#274370000000
1!
1%
1-
12
#274380000000
0!
0%
b111 *
0-
02
b111 6
#274390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#274400000000
0!
0%
b0 *
0-
02
b0 6
#274410000000
1!
1%
1-
12
#274420000000
0!
0%
b1 *
0-
02
b1 6
#274430000000
1!
1%
1-
12
#274440000000
0!
0%
b10 *
0-
02
b10 6
#274450000000
1!
1%
1-
12
#274460000000
0!
0%
b11 *
0-
02
b11 6
#274470000000
1!
1%
1-
12
15
#274480000000
0!
0%
b100 *
0-
02
b100 6
#274490000000
1!
1%
1-
12
#274500000000
0!
0%
b101 *
0-
02
b101 6
#274510000000
1!
1%
1-
12
#274520000000
0!
0%
b110 *
0-
02
b110 6
#274530000000
1!
1%
1-
12
#274540000000
0!
0%
b111 *
0-
02
b111 6
#274550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#274560000000
0!
0%
b0 *
0-
02
b0 6
#274570000000
1!
1%
1-
12
#274580000000
0!
0%
b1 *
0-
02
b1 6
#274590000000
1!
1%
1-
12
#274600000000
0!
0%
b10 *
0-
02
b10 6
#274610000000
1!
1%
1-
12
#274620000000
0!
0%
b11 *
0-
02
b11 6
#274630000000
1!
1%
1-
12
15
#274640000000
0!
0%
b100 *
0-
02
b100 6
#274650000000
1!
1%
1-
12
#274660000000
0!
0%
b101 *
0-
02
b101 6
#274670000000
1!
1%
1-
12
#274680000000
0!
0%
b110 *
0-
02
b110 6
#274690000000
1!
1%
1-
12
#274700000000
0!
0%
b111 *
0-
02
b111 6
#274710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#274720000000
0!
0%
b0 *
0-
02
b0 6
#274730000000
1!
1%
1-
12
#274740000000
0!
0%
b1 *
0-
02
b1 6
#274750000000
1!
1%
1-
12
#274760000000
0!
0%
b10 *
0-
02
b10 6
#274770000000
1!
1%
1-
12
#274780000000
0!
0%
b11 *
0-
02
b11 6
#274790000000
1!
1%
1-
12
15
#274800000000
0!
0%
b100 *
0-
02
b100 6
#274810000000
1!
1%
1-
12
#274820000000
0!
0%
b101 *
0-
02
b101 6
#274830000000
1!
1%
1-
12
#274840000000
0!
0%
b110 *
0-
02
b110 6
#274850000000
1!
1%
1-
12
#274860000000
0!
0%
b111 *
0-
02
b111 6
#274870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#274880000000
0!
0%
b0 *
0-
02
b0 6
#274890000000
1!
1%
1-
12
#274900000000
0!
0%
b1 *
0-
02
b1 6
#274910000000
1!
1%
1-
12
#274920000000
0!
0%
b10 *
0-
02
b10 6
#274930000000
1!
1%
1-
12
#274940000000
0!
0%
b11 *
0-
02
b11 6
#274950000000
1!
1%
1-
12
15
#274960000000
0!
0%
b100 *
0-
02
b100 6
#274970000000
1!
1%
1-
12
#274980000000
0!
0%
b101 *
0-
02
b101 6
#274990000000
1!
1%
1-
12
#275000000000
0!
0%
b110 *
0-
02
b110 6
#275010000000
1!
1%
1-
12
#275020000000
0!
0%
b111 *
0-
02
b111 6
#275030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#275040000000
0!
0%
b0 *
0-
02
b0 6
#275050000000
1!
1%
1-
12
#275060000000
0!
0%
b1 *
0-
02
b1 6
#275070000000
1!
1%
1-
12
#275080000000
0!
0%
b10 *
0-
02
b10 6
#275090000000
1!
1%
1-
12
#275100000000
0!
0%
b11 *
0-
02
b11 6
#275110000000
1!
1%
1-
12
15
#275120000000
0!
0%
b100 *
0-
02
b100 6
#275130000000
1!
1%
1-
12
#275140000000
0!
0%
b101 *
0-
02
b101 6
#275150000000
1!
1%
1-
12
#275160000000
0!
0%
b110 *
0-
02
b110 6
#275170000000
1!
1%
1-
12
#275180000000
0!
0%
b111 *
0-
02
b111 6
#275190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#275200000000
0!
0%
b0 *
0-
02
b0 6
#275210000000
1!
1%
1-
12
#275220000000
0!
0%
b1 *
0-
02
b1 6
#275230000000
1!
1%
1-
12
#275240000000
0!
0%
b10 *
0-
02
b10 6
#275250000000
1!
1%
1-
12
#275260000000
0!
0%
b11 *
0-
02
b11 6
#275270000000
1!
1%
1-
12
15
#275280000000
0!
0%
b100 *
0-
02
b100 6
#275290000000
1!
1%
1-
12
#275300000000
0!
0%
b101 *
0-
02
b101 6
#275310000000
1!
1%
1-
12
#275320000000
0!
0%
b110 *
0-
02
b110 6
#275330000000
1!
1%
1-
12
#275340000000
0!
0%
b111 *
0-
02
b111 6
#275350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#275360000000
0!
0%
b0 *
0-
02
b0 6
#275370000000
1!
1%
1-
12
#275380000000
0!
0%
b1 *
0-
02
b1 6
#275390000000
1!
1%
1-
12
#275400000000
0!
0%
b10 *
0-
02
b10 6
#275410000000
1!
1%
1-
12
#275420000000
0!
0%
b11 *
0-
02
b11 6
#275430000000
1!
1%
1-
12
15
#275440000000
0!
0%
b100 *
0-
02
b100 6
#275450000000
1!
1%
1-
12
#275460000000
0!
0%
b101 *
0-
02
b101 6
#275470000000
1!
1%
1-
12
#275480000000
0!
0%
b110 *
0-
02
b110 6
#275490000000
1!
1%
1-
12
#275500000000
0!
0%
b111 *
0-
02
b111 6
#275510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#275520000000
0!
0%
b0 *
0-
02
b0 6
#275530000000
1!
1%
1-
12
#275540000000
0!
0%
b1 *
0-
02
b1 6
#275550000000
1!
1%
1-
12
#275560000000
0!
0%
b10 *
0-
02
b10 6
#275570000000
1!
1%
1-
12
#275580000000
0!
0%
b11 *
0-
02
b11 6
#275590000000
1!
1%
1-
12
15
#275600000000
0!
0%
b100 *
0-
02
b100 6
#275610000000
1!
1%
1-
12
#275620000000
0!
0%
b101 *
0-
02
b101 6
#275630000000
1!
1%
1-
12
#275640000000
0!
0%
b110 *
0-
02
b110 6
#275650000000
1!
1%
1-
12
#275660000000
0!
0%
b111 *
0-
02
b111 6
#275670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#275680000000
0!
0%
b0 *
0-
02
b0 6
#275690000000
1!
1%
1-
12
#275700000000
0!
0%
b1 *
0-
02
b1 6
#275710000000
1!
1%
1-
12
#275720000000
0!
0%
b10 *
0-
02
b10 6
#275730000000
1!
1%
1-
12
#275740000000
0!
0%
b11 *
0-
02
b11 6
#275750000000
1!
1%
1-
12
15
#275760000000
0!
0%
b100 *
0-
02
b100 6
#275770000000
1!
1%
1-
12
#275780000000
0!
0%
b101 *
0-
02
b101 6
#275790000000
1!
1%
1-
12
#275800000000
0!
0%
b110 *
0-
02
b110 6
#275810000000
1!
1%
1-
12
#275820000000
0!
0%
b111 *
0-
02
b111 6
#275830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#275840000000
0!
0%
b0 *
0-
02
b0 6
#275850000000
1!
1%
1-
12
#275860000000
0!
0%
b1 *
0-
02
b1 6
#275870000000
1!
1%
1-
12
#275880000000
0!
0%
b10 *
0-
02
b10 6
#275890000000
1!
1%
1-
12
#275900000000
0!
0%
b11 *
0-
02
b11 6
#275910000000
1!
1%
1-
12
15
#275920000000
0!
0%
b100 *
0-
02
b100 6
#275930000000
1!
1%
1-
12
#275940000000
0!
0%
b101 *
0-
02
b101 6
#275950000000
1!
1%
1-
12
#275960000000
0!
0%
b110 *
0-
02
b110 6
#275970000000
1!
1%
1-
12
#275980000000
0!
0%
b111 *
0-
02
b111 6
#275990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#276000000000
0!
0%
b0 *
0-
02
b0 6
#276010000000
1!
1%
1-
12
#276020000000
0!
0%
b1 *
0-
02
b1 6
#276030000000
1!
1%
1-
12
#276040000000
0!
0%
b10 *
0-
02
b10 6
#276050000000
1!
1%
1-
12
#276060000000
0!
0%
b11 *
0-
02
b11 6
#276070000000
1!
1%
1-
12
15
#276080000000
0!
0%
b100 *
0-
02
b100 6
#276090000000
1!
1%
1-
12
#276100000000
0!
0%
b101 *
0-
02
b101 6
#276110000000
1!
1%
1-
12
#276120000000
0!
0%
b110 *
0-
02
b110 6
#276130000000
1!
1%
1-
12
#276140000000
0!
0%
b111 *
0-
02
b111 6
#276150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#276160000000
0!
0%
b0 *
0-
02
b0 6
#276170000000
1!
1%
1-
12
#276180000000
0!
0%
b1 *
0-
02
b1 6
#276190000000
1!
1%
1-
12
#276200000000
0!
0%
b10 *
0-
02
b10 6
#276210000000
1!
1%
1-
12
#276220000000
0!
0%
b11 *
0-
02
b11 6
#276230000000
1!
1%
1-
12
15
#276240000000
0!
0%
b100 *
0-
02
b100 6
#276250000000
1!
1%
1-
12
#276260000000
0!
0%
b101 *
0-
02
b101 6
#276270000000
1!
1%
1-
12
#276280000000
0!
0%
b110 *
0-
02
b110 6
#276290000000
1!
1%
1-
12
#276300000000
0!
0%
b111 *
0-
02
b111 6
#276310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#276320000000
0!
0%
b0 *
0-
02
b0 6
#276330000000
1!
1%
1-
12
#276340000000
0!
0%
b1 *
0-
02
b1 6
#276350000000
1!
1%
1-
12
#276360000000
0!
0%
b10 *
0-
02
b10 6
#276370000000
1!
1%
1-
12
#276380000000
0!
0%
b11 *
0-
02
b11 6
#276390000000
1!
1%
1-
12
15
#276400000000
0!
0%
b100 *
0-
02
b100 6
#276410000000
1!
1%
1-
12
#276420000000
0!
0%
b101 *
0-
02
b101 6
#276430000000
1!
1%
1-
12
#276440000000
0!
0%
b110 *
0-
02
b110 6
#276450000000
1!
1%
1-
12
#276460000000
0!
0%
b111 *
0-
02
b111 6
#276470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#276480000000
0!
0%
b0 *
0-
02
b0 6
#276490000000
1!
1%
1-
12
#276500000000
0!
0%
b1 *
0-
02
b1 6
#276510000000
1!
1%
1-
12
#276520000000
0!
0%
b10 *
0-
02
b10 6
#276530000000
1!
1%
1-
12
#276540000000
0!
0%
b11 *
0-
02
b11 6
#276550000000
1!
1%
1-
12
15
#276560000000
0!
0%
b100 *
0-
02
b100 6
#276570000000
1!
1%
1-
12
#276580000000
0!
0%
b101 *
0-
02
b101 6
#276590000000
1!
1%
1-
12
#276600000000
0!
0%
b110 *
0-
02
b110 6
#276610000000
1!
1%
1-
12
#276620000000
0!
0%
b111 *
0-
02
b111 6
#276630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#276640000000
0!
0%
b0 *
0-
02
b0 6
#276650000000
1!
1%
1-
12
#276660000000
0!
0%
b1 *
0-
02
b1 6
#276670000000
1!
1%
1-
12
#276680000000
0!
0%
b10 *
0-
02
b10 6
#276690000000
1!
1%
1-
12
#276700000000
0!
0%
b11 *
0-
02
b11 6
#276710000000
1!
1%
1-
12
15
#276720000000
0!
0%
b100 *
0-
02
b100 6
#276730000000
1!
1%
1-
12
#276740000000
0!
0%
b101 *
0-
02
b101 6
#276750000000
1!
1%
1-
12
#276760000000
0!
0%
b110 *
0-
02
b110 6
#276770000000
1!
1%
1-
12
#276780000000
0!
0%
b111 *
0-
02
b111 6
#276790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#276800000000
0!
0%
b0 *
0-
02
b0 6
#276810000000
1!
1%
1-
12
#276820000000
0!
0%
b1 *
0-
02
b1 6
#276830000000
1!
1%
1-
12
#276840000000
0!
0%
b10 *
0-
02
b10 6
#276850000000
1!
1%
1-
12
#276860000000
0!
0%
b11 *
0-
02
b11 6
#276870000000
1!
1%
1-
12
15
#276880000000
0!
0%
b100 *
0-
02
b100 6
#276890000000
1!
1%
1-
12
#276900000000
0!
0%
b101 *
0-
02
b101 6
#276910000000
1!
1%
1-
12
#276920000000
0!
0%
b110 *
0-
02
b110 6
#276930000000
1!
1%
1-
12
#276940000000
0!
0%
b111 *
0-
02
b111 6
#276950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#276960000000
0!
0%
b0 *
0-
02
b0 6
#276970000000
1!
1%
1-
12
#276980000000
0!
0%
b1 *
0-
02
b1 6
#276990000000
1!
1%
1-
12
#277000000000
0!
0%
b10 *
0-
02
b10 6
#277010000000
1!
1%
1-
12
#277020000000
0!
0%
b11 *
0-
02
b11 6
#277030000000
1!
1%
1-
12
15
#277040000000
0!
0%
b100 *
0-
02
b100 6
#277050000000
1!
1%
1-
12
#277060000000
0!
0%
b101 *
0-
02
b101 6
#277070000000
1!
1%
1-
12
#277080000000
0!
0%
b110 *
0-
02
b110 6
#277090000000
1!
1%
1-
12
#277100000000
0!
0%
b111 *
0-
02
b111 6
#277110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#277120000000
0!
0%
b0 *
0-
02
b0 6
#277130000000
1!
1%
1-
12
#277140000000
0!
0%
b1 *
0-
02
b1 6
#277150000000
1!
1%
1-
12
#277160000000
0!
0%
b10 *
0-
02
b10 6
#277170000000
1!
1%
1-
12
#277180000000
0!
0%
b11 *
0-
02
b11 6
#277190000000
1!
1%
1-
12
15
#277200000000
0!
0%
b100 *
0-
02
b100 6
#277210000000
1!
1%
1-
12
#277220000000
0!
0%
b101 *
0-
02
b101 6
#277230000000
1!
1%
1-
12
#277240000000
0!
0%
b110 *
0-
02
b110 6
#277250000000
1!
1%
1-
12
#277260000000
0!
0%
b111 *
0-
02
b111 6
#277270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#277280000000
0!
0%
b0 *
0-
02
b0 6
#277290000000
1!
1%
1-
12
#277300000000
0!
0%
b1 *
0-
02
b1 6
#277310000000
1!
1%
1-
12
#277320000000
0!
0%
b10 *
0-
02
b10 6
#277330000000
1!
1%
1-
12
#277340000000
0!
0%
b11 *
0-
02
b11 6
#277350000000
1!
1%
1-
12
15
#277360000000
0!
0%
b100 *
0-
02
b100 6
#277370000000
1!
1%
1-
12
#277380000000
0!
0%
b101 *
0-
02
b101 6
#277390000000
1!
1%
1-
12
#277400000000
0!
0%
b110 *
0-
02
b110 6
#277410000000
1!
1%
1-
12
#277420000000
0!
0%
b111 *
0-
02
b111 6
#277430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#277440000000
0!
0%
b0 *
0-
02
b0 6
#277450000000
1!
1%
1-
12
#277460000000
0!
0%
b1 *
0-
02
b1 6
#277470000000
1!
1%
1-
12
#277480000000
0!
0%
b10 *
0-
02
b10 6
#277490000000
1!
1%
1-
12
#277500000000
0!
0%
b11 *
0-
02
b11 6
#277510000000
1!
1%
1-
12
15
#277520000000
0!
0%
b100 *
0-
02
b100 6
#277530000000
1!
1%
1-
12
#277540000000
0!
0%
b101 *
0-
02
b101 6
#277550000000
1!
1%
1-
12
#277560000000
0!
0%
b110 *
0-
02
b110 6
#277570000000
1!
1%
1-
12
#277580000000
0!
0%
b111 *
0-
02
b111 6
#277590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#277600000000
0!
0%
b0 *
0-
02
b0 6
#277610000000
1!
1%
1-
12
#277620000000
0!
0%
b1 *
0-
02
b1 6
#277630000000
1!
1%
1-
12
#277640000000
0!
0%
b10 *
0-
02
b10 6
#277650000000
1!
1%
1-
12
#277660000000
0!
0%
b11 *
0-
02
b11 6
#277670000000
1!
1%
1-
12
15
#277680000000
0!
0%
b100 *
0-
02
b100 6
#277690000000
1!
1%
1-
12
#277700000000
0!
0%
b101 *
0-
02
b101 6
#277710000000
1!
1%
1-
12
#277720000000
0!
0%
b110 *
0-
02
b110 6
#277730000000
1!
1%
1-
12
#277740000000
0!
0%
b111 *
0-
02
b111 6
#277750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#277760000000
0!
0%
b0 *
0-
02
b0 6
#277770000000
1!
1%
1-
12
#277780000000
0!
0%
b1 *
0-
02
b1 6
#277790000000
1!
1%
1-
12
#277800000000
0!
0%
b10 *
0-
02
b10 6
#277810000000
1!
1%
1-
12
#277820000000
0!
0%
b11 *
0-
02
b11 6
#277830000000
1!
1%
1-
12
15
#277840000000
0!
0%
b100 *
0-
02
b100 6
#277850000000
1!
1%
1-
12
#277860000000
0!
0%
b101 *
0-
02
b101 6
#277870000000
1!
1%
1-
12
#277880000000
0!
0%
b110 *
0-
02
b110 6
#277890000000
1!
1%
1-
12
#277900000000
0!
0%
b111 *
0-
02
b111 6
#277910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#277920000000
0!
0%
b0 *
0-
02
b0 6
#277930000000
1!
1%
1-
12
#277940000000
0!
0%
b1 *
0-
02
b1 6
#277950000000
1!
1%
1-
12
#277960000000
0!
0%
b10 *
0-
02
b10 6
#277970000000
1!
1%
1-
12
#277980000000
0!
0%
b11 *
0-
02
b11 6
#277990000000
1!
1%
1-
12
15
#278000000000
0!
0%
b100 *
0-
02
b100 6
#278010000000
1!
1%
1-
12
#278020000000
0!
0%
b101 *
0-
02
b101 6
#278030000000
1!
1%
1-
12
#278040000000
0!
0%
b110 *
0-
02
b110 6
#278050000000
1!
1%
1-
12
#278060000000
0!
0%
b111 *
0-
02
b111 6
#278070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#278080000000
0!
0%
b0 *
0-
02
b0 6
#278090000000
1!
1%
1-
12
#278100000000
0!
0%
b1 *
0-
02
b1 6
#278110000000
1!
1%
1-
12
#278120000000
0!
0%
b10 *
0-
02
b10 6
#278130000000
1!
1%
1-
12
#278140000000
0!
0%
b11 *
0-
02
b11 6
#278150000000
1!
1%
1-
12
15
#278160000000
0!
0%
b100 *
0-
02
b100 6
#278170000000
1!
1%
1-
12
#278180000000
0!
0%
b101 *
0-
02
b101 6
#278190000000
1!
1%
1-
12
#278200000000
0!
0%
b110 *
0-
02
b110 6
#278210000000
1!
1%
1-
12
#278220000000
0!
0%
b111 *
0-
02
b111 6
#278230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#278240000000
0!
0%
b0 *
0-
02
b0 6
#278250000000
1!
1%
1-
12
#278260000000
0!
0%
b1 *
0-
02
b1 6
#278270000000
1!
1%
1-
12
#278280000000
0!
0%
b10 *
0-
02
b10 6
#278290000000
1!
1%
1-
12
#278300000000
0!
0%
b11 *
0-
02
b11 6
#278310000000
1!
1%
1-
12
15
#278320000000
0!
0%
b100 *
0-
02
b100 6
#278330000000
1!
1%
1-
12
#278340000000
0!
0%
b101 *
0-
02
b101 6
#278350000000
1!
1%
1-
12
#278360000000
0!
0%
b110 *
0-
02
b110 6
#278370000000
1!
1%
1-
12
#278380000000
0!
0%
b111 *
0-
02
b111 6
#278390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#278400000000
0!
0%
b0 *
0-
02
b0 6
#278410000000
1!
1%
1-
12
#278420000000
0!
0%
b1 *
0-
02
b1 6
#278430000000
1!
1%
1-
12
#278440000000
0!
0%
b10 *
0-
02
b10 6
#278450000000
1!
1%
1-
12
#278460000000
0!
0%
b11 *
0-
02
b11 6
#278470000000
1!
1%
1-
12
15
#278480000000
0!
0%
b100 *
0-
02
b100 6
#278490000000
1!
1%
1-
12
#278500000000
0!
0%
b101 *
0-
02
b101 6
#278510000000
1!
1%
1-
12
#278520000000
0!
0%
b110 *
0-
02
b110 6
#278530000000
1!
1%
1-
12
#278540000000
0!
0%
b111 *
0-
02
b111 6
#278550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#278560000000
0!
0%
b0 *
0-
02
b0 6
#278570000000
1!
1%
1-
12
#278580000000
0!
0%
b1 *
0-
02
b1 6
#278590000000
1!
1%
1-
12
#278600000000
0!
0%
b10 *
0-
02
b10 6
#278610000000
1!
1%
1-
12
#278620000000
0!
0%
b11 *
0-
02
b11 6
#278630000000
1!
1%
1-
12
15
#278640000000
0!
0%
b100 *
0-
02
b100 6
#278650000000
1!
1%
1-
12
#278660000000
0!
0%
b101 *
0-
02
b101 6
#278670000000
1!
1%
1-
12
#278680000000
0!
0%
b110 *
0-
02
b110 6
#278690000000
1!
1%
1-
12
#278700000000
0!
0%
b111 *
0-
02
b111 6
#278710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#278720000000
0!
0%
b0 *
0-
02
b0 6
#278730000000
1!
1%
1-
12
#278740000000
0!
0%
b1 *
0-
02
b1 6
#278750000000
1!
1%
1-
12
#278760000000
0!
0%
b10 *
0-
02
b10 6
#278770000000
1!
1%
1-
12
#278780000000
0!
0%
b11 *
0-
02
b11 6
#278790000000
1!
1%
1-
12
15
#278800000000
0!
0%
b100 *
0-
02
b100 6
#278810000000
1!
1%
1-
12
#278820000000
0!
0%
b101 *
0-
02
b101 6
#278830000000
1!
1%
1-
12
#278840000000
0!
0%
b110 *
0-
02
b110 6
#278850000000
1!
1%
1-
12
#278860000000
0!
0%
b111 *
0-
02
b111 6
#278870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#278880000000
0!
0%
b0 *
0-
02
b0 6
#278890000000
1!
1%
1-
12
#278900000000
0!
0%
b1 *
0-
02
b1 6
#278910000000
1!
1%
1-
12
#278920000000
0!
0%
b10 *
0-
02
b10 6
#278930000000
1!
1%
1-
12
#278940000000
0!
0%
b11 *
0-
02
b11 6
#278950000000
1!
1%
1-
12
15
#278960000000
0!
0%
b100 *
0-
02
b100 6
#278970000000
1!
1%
1-
12
#278980000000
0!
0%
b101 *
0-
02
b101 6
#278990000000
1!
1%
1-
12
#279000000000
0!
0%
b110 *
0-
02
b110 6
#279010000000
1!
1%
1-
12
#279020000000
0!
0%
b111 *
0-
02
b111 6
#279030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#279040000000
0!
0%
b0 *
0-
02
b0 6
#279050000000
1!
1%
1-
12
#279060000000
0!
0%
b1 *
0-
02
b1 6
#279070000000
1!
1%
1-
12
#279080000000
0!
0%
b10 *
0-
02
b10 6
#279090000000
1!
1%
1-
12
#279100000000
0!
0%
b11 *
0-
02
b11 6
#279110000000
1!
1%
1-
12
15
#279120000000
0!
0%
b100 *
0-
02
b100 6
#279130000000
1!
1%
1-
12
#279140000000
0!
0%
b101 *
0-
02
b101 6
#279150000000
1!
1%
1-
12
#279160000000
0!
0%
b110 *
0-
02
b110 6
#279170000000
1!
1%
1-
12
#279180000000
0!
0%
b111 *
0-
02
b111 6
#279190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#279200000000
0!
0%
b0 *
0-
02
b0 6
#279210000000
1!
1%
1-
12
#279220000000
0!
0%
b1 *
0-
02
b1 6
#279230000000
1!
1%
1-
12
#279240000000
0!
0%
b10 *
0-
02
b10 6
#279250000000
1!
1%
1-
12
#279260000000
0!
0%
b11 *
0-
02
b11 6
#279270000000
1!
1%
1-
12
15
#279280000000
0!
0%
b100 *
0-
02
b100 6
#279290000000
1!
1%
1-
12
#279300000000
0!
0%
b101 *
0-
02
b101 6
#279310000000
1!
1%
1-
12
#279320000000
0!
0%
b110 *
0-
02
b110 6
#279330000000
1!
1%
1-
12
#279340000000
0!
0%
b111 *
0-
02
b111 6
#279350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#279360000000
0!
0%
b0 *
0-
02
b0 6
#279370000000
1!
1%
1-
12
#279380000000
0!
0%
b1 *
0-
02
b1 6
#279390000000
1!
1%
1-
12
#279400000000
0!
0%
b10 *
0-
02
b10 6
#279410000000
1!
1%
1-
12
#279420000000
0!
0%
b11 *
0-
02
b11 6
#279430000000
1!
1%
1-
12
15
#279440000000
0!
0%
b100 *
0-
02
b100 6
#279450000000
1!
1%
1-
12
#279460000000
0!
0%
b101 *
0-
02
b101 6
#279470000000
1!
1%
1-
12
#279480000000
0!
0%
b110 *
0-
02
b110 6
#279490000000
1!
1%
1-
12
#279500000000
0!
0%
b111 *
0-
02
b111 6
#279510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#279520000000
0!
0%
b0 *
0-
02
b0 6
#279530000000
1!
1%
1-
12
#279540000000
0!
0%
b1 *
0-
02
b1 6
#279550000000
1!
1%
1-
12
#279560000000
0!
0%
b10 *
0-
02
b10 6
#279570000000
1!
1%
1-
12
#279580000000
0!
0%
b11 *
0-
02
b11 6
#279590000000
1!
1%
1-
12
15
#279600000000
0!
0%
b100 *
0-
02
b100 6
#279610000000
1!
1%
1-
12
#279620000000
0!
0%
b101 *
0-
02
b101 6
#279630000000
1!
1%
1-
12
#279640000000
0!
0%
b110 *
0-
02
b110 6
#279650000000
1!
1%
1-
12
#279660000000
0!
0%
b111 *
0-
02
b111 6
#279670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#279680000000
0!
0%
b0 *
0-
02
b0 6
#279690000000
1!
1%
1-
12
#279700000000
0!
0%
b1 *
0-
02
b1 6
#279710000000
1!
1%
1-
12
#279720000000
0!
0%
b10 *
0-
02
b10 6
#279730000000
1!
1%
1-
12
#279740000000
0!
0%
b11 *
0-
02
b11 6
#279750000000
1!
1%
1-
12
15
#279760000000
0!
0%
b100 *
0-
02
b100 6
#279770000000
1!
1%
1-
12
#279780000000
0!
0%
b101 *
0-
02
b101 6
#279790000000
1!
1%
1-
12
#279800000000
0!
0%
b110 *
0-
02
b110 6
#279810000000
1!
1%
1-
12
#279820000000
0!
0%
b111 *
0-
02
b111 6
#279830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#279840000000
0!
0%
b0 *
0-
02
b0 6
#279850000000
1!
1%
1-
12
#279860000000
0!
0%
b1 *
0-
02
b1 6
#279870000000
1!
1%
1-
12
#279880000000
0!
0%
b10 *
0-
02
b10 6
#279890000000
1!
1%
1-
12
#279900000000
0!
0%
b11 *
0-
02
b11 6
#279910000000
1!
1%
1-
12
15
#279920000000
0!
0%
b100 *
0-
02
b100 6
#279930000000
1!
1%
1-
12
#279940000000
0!
0%
b101 *
0-
02
b101 6
#279950000000
1!
1%
1-
12
#279960000000
0!
0%
b110 *
0-
02
b110 6
#279970000000
1!
1%
1-
12
#279980000000
0!
0%
b111 *
0-
02
b111 6
#279990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#280000000000
0!
0%
b0 *
0-
02
b0 6
#280010000000
1!
1%
1-
12
#280020000000
0!
0%
b1 *
0-
02
b1 6
#280030000000
1!
1%
1-
12
#280040000000
0!
0%
b10 *
0-
02
b10 6
#280050000000
1!
1%
1-
12
#280060000000
0!
0%
b11 *
0-
02
b11 6
#280070000000
1!
1%
1-
12
15
#280080000000
0!
0%
b100 *
0-
02
b100 6
#280090000000
1!
1%
1-
12
#280100000000
0!
0%
b101 *
0-
02
b101 6
#280110000000
1!
1%
1-
12
#280120000000
0!
0%
b110 *
0-
02
b110 6
#280130000000
1!
1%
1-
12
#280140000000
0!
0%
b111 *
0-
02
b111 6
#280150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#280160000000
0!
0%
b0 *
0-
02
b0 6
#280170000000
1!
1%
1-
12
#280180000000
0!
0%
b1 *
0-
02
b1 6
#280190000000
1!
1%
1-
12
#280200000000
0!
0%
b10 *
0-
02
b10 6
#280210000000
1!
1%
1-
12
#280220000000
0!
0%
b11 *
0-
02
b11 6
#280230000000
1!
1%
1-
12
15
#280240000000
0!
0%
b100 *
0-
02
b100 6
#280250000000
1!
1%
1-
12
#280260000000
0!
0%
b101 *
0-
02
b101 6
#280270000000
1!
1%
1-
12
#280280000000
0!
0%
b110 *
0-
02
b110 6
#280290000000
1!
1%
1-
12
#280300000000
0!
0%
b111 *
0-
02
b111 6
#280310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#280320000000
0!
0%
b0 *
0-
02
b0 6
#280330000000
1!
1%
1-
12
#280340000000
0!
0%
b1 *
0-
02
b1 6
#280350000000
1!
1%
1-
12
#280360000000
0!
0%
b10 *
0-
02
b10 6
#280370000000
1!
1%
1-
12
#280380000000
0!
0%
b11 *
0-
02
b11 6
#280390000000
1!
1%
1-
12
15
#280400000000
0!
0%
b100 *
0-
02
b100 6
#280410000000
1!
1%
1-
12
#280420000000
0!
0%
b101 *
0-
02
b101 6
#280430000000
1!
1%
1-
12
#280440000000
0!
0%
b110 *
0-
02
b110 6
#280450000000
1!
1%
1-
12
#280460000000
0!
0%
b111 *
0-
02
b111 6
#280470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#280480000000
0!
0%
b0 *
0-
02
b0 6
#280490000000
1!
1%
1-
12
#280500000000
0!
0%
b1 *
0-
02
b1 6
#280510000000
1!
1%
1-
12
#280520000000
0!
0%
b10 *
0-
02
b10 6
#280530000000
1!
1%
1-
12
#280540000000
0!
0%
b11 *
0-
02
b11 6
#280550000000
1!
1%
1-
12
15
#280560000000
0!
0%
b100 *
0-
02
b100 6
#280570000000
1!
1%
1-
12
#280580000000
0!
0%
b101 *
0-
02
b101 6
#280590000000
1!
1%
1-
12
#280600000000
0!
0%
b110 *
0-
02
b110 6
#280610000000
1!
1%
1-
12
#280620000000
0!
0%
b111 *
0-
02
b111 6
#280630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#280640000000
0!
0%
b0 *
0-
02
b0 6
#280650000000
1!
1%
1-
12
#280660000000
0!
0%
b1 *
0-
02
b1 6
#280670000000
1!
1%
1-
12
#280680000000
0!
0%
b10 *
0-
02
b10 6
#280690000000
1!
1%
1-
12
#280700000000
0!
0%
b11 *
0-
02
b11 6
#280710000000
1!
1%
1-
12
15
#280720000000
0!
0%
b100 *
0-
02
b100 6
#280730000000
1!
1%
1-
12
#280740000000
0!
0%
b101 *
0-
02
b101 6
#280750000000
1!
1%
1-
12
#280760000000
0!
0%
b110 *
0-
02
b110 6
#280770000000
1!
1%
1-
12
#280780000000
0!
0%
b111 *
0-
02
b111 6
#280790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#280800000000
0!
0%
b0 *
0-
02
b0 6
#280810000000
1!
1%
1-
12
#280820000000
0!
0%
b1 *
0-
02
b1 6
#280830000000
1!
1%
1-
12
#280840000000
0!
0%
b10 *
0-
02
b10 6
#280850000000
1!
1%
1-
12
#280860000000
0!
0%
b11 *
0-
02
b11 6
#280870000000
1!
1%
1-
12
15
#280880000000
0!
0%
b100 *
0-
02
b100 6
#280890000000
1!
1%
1-
12
#280900000000
0!
0%
b101 *
0-
02
b101 6
#280910000000
1!
1%
1-
12
#280920000000
0!
0%
b110 *
0-
02
b110 6
#280930000000
1!
1%
1-
12
#280940000000
0!
0%
b111 *
0-
02
b111 6
#280950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#280960000000
0!
0%
b0 *
0-
02
b0 6
#280970000000
1!
1%
1-
12
#280980000000
0!
0%
b1 *
0-
02
b1 6
#280990000000
1!
1%
1-
12
#281000000000
0!
0%
b10 *
0-
02
b10 6
#281010000000
1!
1%
1-
12
#281020000000
0!
0%
b11 *
0-
02
b11 6
#281030000000
1!
1%
1-
12
15
#281040000000
0!
0%
b100 *
0-
02
b100 6
#281050000000
1!
1%
1-
12
#281060000000
0!
0%
b101 *
0-
02
b101 6
#281070000000
1!
1%
1-
12
#281080000000
0!
0%
b110 *
0-
02
b110 6
#281090000000
1!
1%
1-
12
#281100000000
0!
0%
b111 *
0-
02
b111 6
#281110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#281120000000
0!
0%
b0 *
0-
02
b0 6
#281130000000
1!
1%
1-
12
#281140000000
0!
0%
b1 *
0-
02
b1 6
#281150000000
1!
1%
1-
12
#281160000000
0!
0%
b10 *
0-
02
b10 6
#281170000000
1!
1%
1-
12
#281180000000
0!
0%
b11 *
0-
02
b11 6
#281190000000
1!
1%
1-
12
15
#281200000000
0!
0%
b100 *
0-
02
b100 6
#281210000000
1!
1%
1-
12
#281220000000
0!
0%
b101 *
0-
02
b101 6
#281230000000
1!
1%
1-
12
#281240000000
0!
0%
b110 *
0-
02
b110 6
#281250000000
1!
1%
1-
12
#281260000000
0!
0%
b111 *
0-
02
b111 6
#281270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#281280000000
0!
0%
b0 *
0-
02
b0 6
#281290000000
1!
1%
1-
12
#281300000000
0!
0%
b1 *
0-
02
b1 6
#281310000000
1!
1%
1-
12
#281320000000
0!
0%
b10 *
0-
02
b10 6
#281330000000
1!
1%
1-
12
#281340000000
0!
0%
b11 *
0-
02
b11 6
#281350000000
1!
1%
1-
12
15
#281360000000
0!
0%
b100 *
0-
02
b100 6
#281370000000
1!
1%
1-
12
#281380000000
0!
0%
b101 *
0-
02
b101 6
#281390000000
1!
1%
1-
12
#281400000000
0!
0%
b110 *
0-
02
b110 6
#281410000000
1!
1%
1-
12
#281420000000
0!
0%
b111 *
0-
02
b111 6
#281430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#281440000000
0!
0%
b0 *
0-
02
b0 6
#281450000000
1!
1%
1-
12
#281460000000
0!
0%
b1 *
0-
02
b1 6
#281470000000
1!
1%
1-
12
#281480000000
0!
0%
b10 *
0-
02
b10 6
#281490000000
1!
1%
1-
12
#281500000000
0!
0%
b11 *
0-
02
b11 6
#281510000000
1!
1%
1-
12
15
#281520000000
0!
0%
b100 *
0-
02
b100 6
#281530000000
1!
1%
1-
12
#281540000000
0!
0%
b101 *
0-
02
b101 6
#281550000000
1!
1%
1-
12
#281560000000
0!
0%
b110 *
0-
02
b110 6
#281570000000
1!
1%
1-
12
#281580000000
0!
0%
b111 *
0-
02
b111 6
#281590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#281600000000
0!
0%
b0 *
0-
02
b0 6
#281610000000
1!
1%
1-
12
#281620000000
0!
0%
b1 *
0-
02
b1 6
#281630000000
1!
1%
1-
12
#281640000000
0!
0%
b10 *
0-
02
b10 6
#281650000000
1!
1%
1-
12
#281660000000
0!
0%
b11 *
0-
02
b11 6
#281670000000
1!
1%
1-
12
15
#281680000000
0!
0%
b100 *
0-
02
b100 6
#281690000000
1!
1%
1-
12
#281700000000
0!
0%
b101 *
0-
02
b101 6
#281710000000
1!
1%
1-
12
#281720000000
0!
0%
b110 *
0-
02
b110 6
#281730000000
1!
1%
1-
12
#281740000000
0!
0%
b111 *
0-
02
b111 6
#281750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#281760000000
0!
0%
b0 *
0-
02
b0 6
#281770000000
1!
1%
1-
12
#281780000000
0!
0%
b1 *
0-
02
b1 6
#281790000000
1!
1%
1-
12
#281800000000
0!
0%
b10 *
0-
02
b10 6
#281810000000
1!
1%
1-
12
#281820000000
0!
0%
b11 *
0-
02
b11 6
#281830000000
1!
1%
1-
12
15
#281840000000
0!
0%
b100 *
0-
02
b100 6
#281850000000
1!
1%
1-
12
#281860000000
0!
0%
b101 *
0-
02
b101 6
#281870000000
1!
1%
1-
12
#281880000000
0!
0%
b110 *
0-
02
b110 6
#281890000000
1!
1%
1-
12
#281900000000
0!
0%
b111 *
0-
02
b111 6
#281910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#281920000000
0!
0%
b0 *
0-
02
b0 6
#281930000000
1!
1%
1-
12
#281940000000
0!
0%
b1 *
0-
02
b1 6
#281950000000
1!
1%
1-
12
#281960000000
0!
0%
b10 *
0-
02
b10 6
#281970000000
1!
1%
1-
12
#281980000000
0!
0%
b11 *
0-
02
b11 6
#281990000000
1!
1%
1-
12
15
#282000000000
0!
0%
b100 *
0-
02
b100 6
#282010000000
1!
1%
1-
12
#282020000000
0!
0%
b101 *
0-
02
b101 6
#282030000000
1!
1%
1-
12
#282040000000
0!
0%
b110 *
0-
02
b110 6
#282050000000
1!
1%
1-
12
#282060000000
0!
0%
b111 *
0-
02
b111 6
#282070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#282080000000
0!
0%
b0 *
0-
02
b0 6
#282090000000
1!
1%
1-
12
#282100000000
0!
0%
b1 *
0-
02
b1 6
#282110000000
1!
1%
1-
12
#282120000000
0!
0%
b10 *
0-
02
b10 6
#282130000000
1!
1%
1-
12
#282140000000
0!
0%
b11 *
0-
02
b11 6
#282150000000
1!
1%
1-
12
15
#282160000000
0!
0%
b100 *
0-
02
b100 6
#282170000000
1!
1%
1-
12
#282180000000
0!
0%
b101 *
0-
02
b101 6
#282190000000
1!
1%
1-
12
#282200000000
0!
0%
b110 *
0-
02
b110 6
#282210000000
1!
1%
1-
12
#282220000000
0!
0%
b111 *
0-
02
b111 6
#282230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#282240000000
0!
0%
b0 *
0-
02
b0 6
#282250000000
1!
1%
1-
12
#282260000000
0!
0%
b1 *
0-
02
b1 6
#282270000000
1!
1%
1-
12
#282280000000
0!
0%
b10 *
0-
02
b10 6
#282290000000
1!
1%
1-
12
#282300000000
0!
0%
b11 *
0-
02
b11 6
#282310000000
1!
1%
1-
12
15
#282320000000
0!
0%
b100 *
0-
02
b100 6
#282330000000
1!
1%
1-
12
#282340000000
0!
0%
b101 *
0-
02
b101 6
#282350000000
1!
1%
1-
12
#282360000000
0!
0%
b110 *
0-
02
b110 6
#282370000000
1!
1%
1-
12
#282380000000
0!
0%
b111 *
0-
02
b111 6
#282390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#282400000000
0!
0%
b0 *
0-
02
b0 6
#282410000000
1!
1%
1-
12
#282420000000
0!
0%
b1 *
0-
02
b1 6
#282430000000
1!
1%
1-
12
#282440000000
0!
0%
b10 *
0-
02
b10 6
#282450000000
1!
1%
1-
12
#282460000000
0!
0%
b11 *
0-
02
b11 6
#282470000000
1!
1%
1-
12
15
#282480000000
0!
0%
b100 *
0-
02
b100 6
#282490000000
1!
1%
1-
12
#282500000000
0!
0%
b101 *
0-
02
b101 6
#282510000000
1!
1%
1-
12
#282520000000
0!
0%
b110 *
0-
02
b110 6
#282530000000
1!
1%
1-
12
#282540000000
0!
0%
b111 *
0-
02
b111 6
#282550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#282560000000
0!
0%
b0 *
0-
02
b0 6
#282570000000
1!
1%
1-
12
#282580000000
0!
0%
b1 *
0-
02
b1 6
#282590000000
1!
1%
1-
12
#282600000000
0!
0%
b10 *
0-
02
b10 6
#282610000000
1!
1%
1-
12
#282620000000
0!
0%
b11 *
0-
02
b11 6
#282630000000
1!
1%
1-
12
15
#282640000000
0!
0%
b100 *
0-
02
b100 6
#282650000000
1!
1%
1-
12
#282660000000
0!
0%
b101 *
0-
02
b101 6
#282670000000
1!
1%
1-
12
#282680000000
0!
0%
b110 *
0-
02
b110 6
#282690000000
1!
1%
1-
12
#282700000000
0!
0%
b111 *
0-
02
b111 6
#282710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#282720000000
0!
0%
b0 *
0-
02
b0 6
#282730000000
1!
1%
1-
12
#282740000000
0!
0%
b1 *
0-
02
b1 6
#282750000000
1!
1%
1-
12
#282760000000
0!
0%
b10 *
0-
02
b10 6
#282770000000
1!
1%
1-
12
#282780000000
0!
0%
b11 *
0-
02
b11 6
#282790000000
1!
1%
1-
12
15
#282800000000
0!
0%
b100 *
0-
02
b100 6
#282810000000
1!
1%
1-
12
#282820000000
0!
0%
b101 *
0-
02
b101 6
#282830000000
1!
1%
1-
12
#282840000000
0!
0%
b110 *
0-
02
b110 6
#282850000000
1!
1%
1-
12
#282860000000
0!
0%
b111 *
0-
02
b111 6
#282870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#282880000000
0!
0%
b0 *
0-
02
b0 6
#282890000000
1!
1%
1-
12
#282900000000
0!
0%
b1 *
0-
02
b1 6
#282910000000
1!
1%
1-
12
#282920000000
0!
0%
b10 *
0-
02
b10 6
#282930000000
1!
1%
1-
12
#282940000000
0!
0%
b11 *
0-
02
b11 6
#282950000000
1!
1%
1-
12
15
#282960000000
0!
0%
b100 *
0-
02
b100 6
#282970000000
1!
1%
1-
12
#282980000000
0!
0%
b101 *
0-
02
b101 6
#282990000000
1!
1%
1-
12
#283000000000
0!
0%
b110 *
0-
02
b110 6
#283010000000
1!
1%
1-
12
#283020000000
0!
0%
b111 *
0-
02
b111 6
#283030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#283040000000
0!
0%
b0 *
0-
02
b0 6
#283050000000
1!
1%
1-
12
#283060000000
0!
0%
b1 *
0-
02
b1 6
#283070000000
1!
1%
1-
12
#283080000000
0!
0%
b10 *
0-
02
b10 6
#283090000000
1!
1%
1-
12
#283100000000
0!
0%
b11 *
0-
02
b11 6
#283110000000
1!
1%
1-
12
15
#283120000000
0!
0%
b100 *
0-
02
b100 6
#283130000000
1!
1%
1-
12
#283140000000
0!
0%
b101 *
0-
02
b101 6
#283150000000
1!
1%
1-
12
#283160000000
0!
0%
b110 *
0-
02
b110 6
#283170000000
1!
1%
1-
12
#283180000000
0!
0%
b111 *
0-
02
b111 6
#283190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#283200000000
0!
0%
b0 *
0-
02
b0 6
#283210000000
1!
1%
1-
12
#283220000000
0!
0%
b1 *
0-
02
b1 6
#283230000000
1!
1%
1-
12
#283240000000
0!
0%
b10 *
0-
02
b10 6
#283250000000
1!
1%
1-
12
#283260000000
0!
0%
b11 *
0-
02
b11 6
#283270000000
1!
1%
1-
12
15
#283280000000
0!
0%
b100 *
0-
02
b100 6
#283290000000
1!
1%
1-
12
#283300000000
0!
0%
b101 *
0-
02
b101 6
#283310000000
1!
1%
1-
12
#283320000000
0!
0%
b110 *
0-
02
b110 6
#283330000000
1!
1%
1-
12
#283340000000
0!
0%
b111 *
0-
02
b111 6
#283350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#283360000000
0!
0%
b0 *
0-
02
b0 6
#283370000000
1!
1%
1-
12
#283380000000
0!
0%
b1 *
0-
02
b1 6
#283390000000
1!
1%
1-
12
#283400000000
0!
0%
b10 *
0-
02
b10 6
#283410000000
1!
1%
1-
12
#283420000000
0!
0%
b11 *
0-
02
b11 6
#283430000000
1!
1%
1-
12
15
#283440000000
0!
0%
b100 *
0-
02
b100 6
#283450000000
1!
1%
1-
12
#283460000000
0!
0%
b101 *
0-
02
b101 6
#283470000000
1!
1%
1-
12
#283480000000
0!
0%
b110 *
0-
02
b110 6
#283490000000
1!
1%
1-
12
#283500000000
0!
0%
b111 *
0-
02
b111 6
#283510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#283520000000
0!
0%
b0 *
0-
02
b0 6
#283530000000
1!
1%
1-
12
#283540000000
0!
0%
b1 *
0-
02
b1 6
#283550000000
1!
1%
1-
12
#283560000000
0!
0%
b10 *
0-
02
b10 6
#283570000000
1!
1%
1-
12
#283580000000
0!
0%
b11 *
0-
02
b11 6
#283590000000
1!
1%
1-
12
15
#283600000000
0!
0%
b100 *
0-
02
b100 6
#283610000000
1!
1%
1-
12
#283620000000
0!
0%
b101 *
0-
02
b101 6
#283630000000
1!
1%
1-
12
#283640000000
0!
0%
b110 *
0-
02
b110 6
#283650000000
1!
1%
1-
12
#283660000000
0!
0%
b111 *
0-
02
b111 6
#283670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#283680000000
0!
0%
b0 *
0-
02
b0 6
#283690000000
1!
1%
1-
12
#283700000000
0!
0%
b1 *
0-
02
b1 6
#283710000000
1!
1%
1-
12
#283720000000
0!
0%
b10 *
0-
02
b10 6
#283730000000
1!
1%
1-
12
#283740000000
0!
0%
b11 *
0-
02
b11 6
#283750000000
1!
1%
1-
12
15
#283760000000
0!
0%
b100 *
0-
02
b100 6
#283770000000
1!
1%
1-
12
#283780000000
0!
0%
b101 *
0-
02
b101 6
#283790000000
1!
1%
1-
12
#283800000000
0!
0%
b110 *
0-
02
b110 6
#283810000000
1!
1%
1-
12
#283820000000
0!
0%
b111 *
0-
02
b111 6
#283830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#283840000000
0!
0%
b0 *
0-
02
b0 6
#283850000000
1!
1%
1-
12
#283860000000
0!
0%
b1 *
0-
02
b1 6
#283870000000
1!
1%
1-
12
#283880000000
0!
0%
b10 *
0-
02
b10 6
#283890000000
1!
1%
1-
12
#283900000000
0!
0%
b11 *
0-
02
b11 6
#283910000000
1!
1%
1-
12
15
#283920000000
0!
0%
b100 *
0-
02
b100 6
#283930000000
1!
1%
1-
12
#283940000000
0!
0%
b101 *
0-
02
b101 6
#283950000000
1!
1%
1-
12
#283960000000
0!
0%
b110 *
0-
02
b110 6
#283970000000
1!
1%
1-
12
#283980000000
0!
0%
b111 *
0-
02
b111 6
#283990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#284000000000
0!
0%
b0 *
0-
02
b0 6
#284010000000
1!
1%
1-
12
#284020000000
0!
0%
b1 *
0-
02
b1 6
#284030000000
1!
1%
1-
12
#284040000000
0!
0%
b10 *
0-
02
b10 6
#284050000000
1!
1%
1-
12
#284060000000
0!
0%
b11 *
0-
02
b11 6
#284070000000
1!
1%
1-
12
15
#284080000000
0!
0%
b100 *
0-
02
b100 6
#284090000000
1!
1%
1-
12
#284100000000
0!
0%
b101 *
0-
02
b101 6
#284110000000
1!
1%
1-
12
#284120000000
0!
0%
b110 *
0-
02
b110 6
#284130000000
1!
1%
1-
12
#284140000000
0!
0%
b111 *
0-
02
b111 6
#284150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#284160000000
0!
0%
b0 *
0-
02
b0 6
#284170000000
1!
1%
1-
12
#284180000000
0!
0%
b1 *
0-
02
b1 6
#284190000000
1!
1%
1-
12
#284200000000
0!
0%
b10 *
0-
02
b10 6
#284210000000
1!
1%
1-
12
#284220000000
0!
0%
b11 *
0-
02
b11 6
#284230000000
1!
1%
1-
12
15
#284240000000
0!
0%
b100 *
0-
02
b100 6
#284250000000
1!
1%
1-
12
#284260000000
0!
0%
b101 *
0-
02
b101 6
#284270000000
1!
1%
1-
12
#284280000000
0!
0%
b110 *
0-
02
b110 6
#284290000000
1!
1%
1-
12
#284300000000
0!
0%
b111 *
0-
02
b111 6
#284310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#284320000000
0!
0%
b0 *
0-
02
b0 6
#284330000000
1!
1%
1-
12
#284340000000
0!
0%
b1 *
0-
02
b1 6
#284350000000
1!
1%
1-
12
#284360000000
0!
0%
b10 *
0-
02
b10 6
#284370000000
1!
1%
1-
12
#284380000000
0!
0%
b11 *
0-
02
b11 6
#284390000000
1!
1%
1-
12
15
#284400000000
0!
0%
b100 *
0-
02
b100 6
#284410000000
1!
1%
1-
12
#284420000000
0!
0%
b101 *
0-
02
b101 6
#284430000000
1!
1%
1-
12
#284440000000
0!
0%
b110 *
0-
02
b110 6
#284450000000
1!
1%
1-
12
#284460000000
0!
0%
b111 *
0-
02
b111 6
#284470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#284480000000
0!
0%
b0 *
0-
02
b0 6
#284490000000
1!
1%
1-
12
#284500000000
0!
0%
b1 *
0-
02
b1 6
#284510000000
1!
1%
1-
12
#284520000000
0!
0%
b10 *
0-
02
b10 6
#284530000000
1!
1%
1-
12
#284540000000
0!
0%
b11 *
0-
02
b11 6
#284550000000
1!
1%
1-
12
15
#284560000000
0!
0%
b100 *
0-
02
b100 6
#284570000000
1!
1%
1-
12
#284580000000
0!
0%
b101 *
0-
02
b101 6
#284590000000
1!
1%
1-
12
#284600000000
0!
0%
b110 *
0-
02
b110 6
#284610000000
1!
1%
1-
12
#284620000000
0!
0%
b111 *
0-
02
b111 6
#284630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#284640000000
0!
0%
b0 *
0-
02
b0 6
#284650000000
1!
1%
1-
12
#284660000000
0!
0%
b1 *
0-
02
b1 6
#284670000000
1!
1%
1-
12
#284680000000
0!
0%
b10 *
0-
02
b10 6
#284690000000
1!
1%
1-
12
#284700000000
0!
0%
b11 *
0-
02
b11 6
#284710000000
1!
1%
1-
12
15
#284720000000
0!
0%
b100 *
0-
02
b100 6
#284730000000
1!
1%
1-
12
#284740000000
0!
0%
b101 *
0-
02
b101 6
#284750000000
1!
1%
1-
12
#284760000000
0!
0%
b110 *
0-
02
b110 6
#284770000000
1!
1%
1-
12
#284780000000
0!
0%
b111 *
0-
02
b111 6
#284790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#284800000000
0!
0%
b0 *
0-
02
b0 6
#284810000000
1!
1%
1-
12
#284820000000
0!
0%
b1 *
0-
02
b1 6
#284830000000
1!
1%
1-
12
#284840000000
0!
0%
b10 *
0-
02
b10 6
#284850000000
1!
1%
1-
12
#284860000000
0!
0%
b11 *
0-
02
b11 6
#284870000000
1!
1%
1-
12
15
#284880000000
0!
0%
b100 *
0-
02
b100 6
#284890000000
1!
1%
1-
12
#284900000000
0!
0%
b101 *
0-
02
b101 6
#284910000000
1!
1%
1-
12
#284920000000
0!
0%
b110 *
0-
02
b110 6
#284930000000
1!
1%
1-
12
#284940000000
0!
0%
b111 *
0-
02
b111 6
#284950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#284960000000
0!
0%
b0 *
0-
02
b0 6
#284970000000
1!
1%
1-
12
#284980000000
0!
0%
b1 *
0-
02
b1 6
#284990000000
1!
1%
1-
12
#285000000000
0!
0%
b10 *
0-
02
b10 6
#285010000000
1!
1%
1-
12
#285020000000
0!
0%
b11 *
0-
02
b11 6
#285030000000
1!
1%
1-
12
15
#285040000000
0!
0%
b100 *
0-
02
b100 6
#285050000000
1!
1%
1-
12
#285060000000
0!
0%
b101 *
0-
02
b101 6
#285070000000
1!
1%
1-
12
#285080000000
0!
0%
b110 *
0-
02
b110 6
#285090000000
1!
1%
1-
12
#285100000000
0!
0%
b111 *
0-
02
b111 6
#285110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#285120000000
0!
0%
b0 *
0-
02
b0 6
#285130000000
1!
1%
1-
12
#285140000000
0!
0%
b1 *
0-
02
b1 6
#285150000000
1!
1%
1-
12
#285160000000
0!
0%
b10 *
0-
02
b10 6
#285170000000
1!
1%
1-
12
#285180000000
0!
0%
b11 *
0-
02
b11 6
#285190000000
1!
1%
1-
12
15
#285200000000
0!
0%
b100 *
0-
02
b100 6
#285210000000
1!
1%
1-
12
#285220000000
0!
0%
b101 *
0-
02
b101 6
#285230000000
1!
1%
1-
12
#285240000000
0!
0%
b110 *
0-
02
b110 6
#285250000000
1!
1%
1-
12
#285260000000
0!
0%
b111 *
0-
02
b111 6
#285270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#285280000000
0!
0%
b0 *
0-
02
b0 6
#285290000000
1!
1%
1-
12
#285300000000
0!
0%
b1 *
0-
02
b1 6
#285310000000
1!
1%
1-
12
#285320000000
0!
0%
b10 *
0-
02
b10 6
#285330000000
1!
1%
1-
12
#285340000000
0!
0%
b11 *
0-
02
b11 6
#285350000000
1!
1%
1-
12
15
#285360000000
0!
0%
b100 *
0-
02
b100 6
#285370000000
1!
1%
1-
12
#285380000000
0!
0%
b101 *
0-
02
b101 6
#285390000000
1!
1%
1-
12
#285400000000
0!
0%
b110 *
0-
02
b110 6
#285410000000
1!
1%
1-
12
#285420000000
0!
0%
b111 *
0-
02
b111 6
#285430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#285440000000
0!
0%
b0 *
0-
02
b0 6
#285450000000
1!
1%
1-
12
#285460000000
0!
0%
b1 *
0-
02
b1 6
#285470000000
1!
1%
1-
12
#285480000000
0!
0%
b10 *
0-
02
b10 6
#285490000000
1!
1%
1-
12
#285500000000
0!
0%
b11 *
0-
02
b11 6
#285510000000
1!
1%
1-
12
15
#285520000000
0!
0%
b100 *
0-
02
b100 6
#285530000000
1!
1%
1-
12
#285540000000
0!
0%
b101 *
0-
02
b101 6
#285550000000
1!
1%
1-
12
#285560000000
0!
0%
b110 *
0-
02
b110 6
#285570000000
1!
1%
1-
12
#285580000000
0!
0%
b111 *
0-
02
b111 6
#285590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#285600000000
0!
0%
b0 *
0-
02
b0 6
#285610000000
1!
1%
1-
12
#285620000000
0!
0%
b1 *
0-
02
b1 6
#285630000000
1!
1%
1-
12
#285640000000
0!
0%
b10 *
0-
02
b10 6
#285650000000
1!
1%
1-
12
#285660000000
0!
0%
b11 *
0-
02
b11 6
#285670000000
1!
1%
1-
12
15
#285680000000
0!
0%
b100 *
0-
02
b100 6
#285690000000
1!
1%
1-
12
#285700000000
0!
0%
b101 *
0-
02
b101 6
#285710000000
1!
1%
1-
12
#285720000000
0!
0%
b110 *
0-
02
b110 6
#285730000000
1!
1%
1-
12
#285740000000
0!
0%
b111 *
0-
02
b111 6
#285750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#285760000000
0!
0%
b0 *
0-
02
b0 6
#285770000000
1!
1%
1-
12
#285780000000
0!
0%
b1 *
0-
02
b1 6
#285790000000
1!
1%
1-
12
#285800000000
0!
0%
b10 *
0-
02
b10 6
#285810000000
1!
1%
1-
12
#285820000000
0!
0%
b11 *
0-
02
b11 6
#285830000000
1!
1%
1-
12
15
#285840000000
0!
0%
b100 *
0-
02
b100 6
#285850000000
1!
1%
1-
12
#285860000000
0!
0%
b101 *
0-
02
b101 6
#285870000000
1!
1%
1-
12
#285880000000
0!
0%
b110 *
0-
02
b110 6
#285890000000
1!
1%
1-
12
#285900000000
0!
0%
b111 *
0-
02
b111 6
#285910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#285920000000
0!
0%
b0 *
0-
02
b0 6
#285930000000
1!
1%
1-
12
#285940000000
0!
0%
b1 *
0-
02
b1 6
#285950000000
1!
1%
1-
12
#285960000000
0!
0%
b10 *
0-
02
b10 6
#285970000000
1!
1%
1-
12
#285980000000
0!
0%
b11 *
0-
02
b11 6
#285990000000
1!
1%
1-
12
15
#286000000000
0!
0%
b100 *
0-
02
b100 6
#286010000000
1!
1%
1-
12
#286020000000
0!
0%
b101 *
0-
02
b101 6
#286030000000
1!
1%
1-
12
#286040000000
0!
0%
b110 *
0-
02
b110 6
#286050000000
1!
1%
1-
12
#286060000000
0!
0%
b111 *
0-
02
b111 6
#286070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#286080000000
0!
0%
b0 *
0-
02
b0 6
#286090000000
1!
1%
1-
12
#286100000000
0!
0%
b1 *
0-
02
b1 6
#286110000000
1!
1%
1-
12
#286120000000
0!
0%
b10 *
0-
02
b10 6
#286130000000
1!
1%
1-
12
#286140000000
0!
0%
b11 *
0-
02
b11 6
#286150000000
1!
1%
1-
12
15
#286160000000
0!
0%
b100 *
0-
02
b100 6
#286170000000
1!
1%
1-
12
#286180000000
0!
0%
b101 *
0-
02
b101 6
#286190000000
1!
1%
1-
12
#286200000000
0!
0%
b110 *
0-
02
b110 6
#286210000000
1!
1%
1-
12
#286220000000
0!
0%
b111 *
0-
02
b111 6
#286230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#286240000000
0!
0%
b0 *
0-
02
b0 6
#286250000000
1!
1%
1-
12
#286260000000
0!
0%
b1 *
0-
02
b1 6
#286270000000
1!
1%
1-
12
#286280000000
0!
0%
b10 *
0-
02
b10 6
#286290000000
1!
1%
1-
12
#286300000000
0!
0%
b11 *
0-
02
b11 6
#286310000000
1!
1%
1-
12
15
#286320000000
0!
0%
b100 *
0-
02
b100 6
#286330000000
1!
1%
1-
12
#286340000000
0!
0%
b101 *
0-
02
b101 6
#286350000000
1!
1%
1-
12
#286360000000
0!
0%
b110 *
0-
02
b110 6
#286370000000
1!
1%
1-
12
#286380000000
0!
0%
b111 *
0-
02
b111 6
#286390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#286400000000
0!
0%
b0 *
0-
02
b0 6
#286410000000
1!
1%
1-
12
#286420000000
0!
0%
b1 *
0-
02
b1 6
#286430000000
1!
1%
1-
12
#286440000000
0!
0%
b10 *
0-
02
b10 6
#286450000000
1!
1%
1-
12
#286460000000
0!
0%
b11 *
0-
02
b11 6
#286470000000
1!
1%
1-
12
15
#286480000000
0!
0%
b100 *
0-
02
b100 6
#286490000000
1!
1%
1-
12
#286500000000
0!
0%
b101 *
0-
02
b101 6
#286510000000
1!
1%
1-
12
#286520000000
0!
0%
b110 *
0-
02
b110 6
#286530000000
1!
1%
1-
12
#286540000000
0!
0%
b111 *
0-
02
b111 6
#286550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#286560000000
0!
0%
b0 *
0-
02
b0 6
#286570000000
1!
1%
1-
12
#286580000000
0!
0%
b1 *
0-
02
b1 6
#286590000000
1!
1%
1-
12
#286600000000
0!
0%
b10 *
0-
02
b10 6
#286610000000
1!
1%
1-
12
#286620000000
0!
0%
b11 *
0-
02
b11 6
#286630000000
1!
1%
1-
12
15
#286640000000
0!
0%
b100 *
0-
02
b100 6
#286650000000
1!
1%
1-
12
#286660000000
0!
0%
b101 *
0-
02
b101 6
#286670000000
1!
1%
1-
12
#286680000000
0!
0%
b110 *
0-
02
b110 6
#286690000000
1!
1%
1-
12
#286700000000
0!
0%
b111 *
0-
02
b111 6
#286710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#286720000000
0!
0%
b0 *
0-
02
b0 6
#286730000000
1!
1%
1-
12
#286740000000
0!
0%
b1 *
0-
02
b1 6
#286750000000
1!
1%
1-
12
#286760000000
0!
0%
b10 *
0-
02
b10 6
#286770000000
1!
1%
1-
12
#286780000000
0!
0%
b11 *
0-
02
b11 6
#286790000000
1!
1%
1-
12
15
#286800000000
0!
0%
b100 *
0-
02
b100 6
#286810000000
1!
1%
1-
12
#286820000000
0!
0%
b101 *
0-
02
b101 6
#286830000000
1!
1%
1-
12
#286840000000
0!
0%
b110 *
0-
02
b110 6
#286850000000
1!
1%
1-
12
#286860000000
0!
0%
b111 *
0-
02
b111 6
#286870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#286880000000
0!
0%
b0 *
0-
02
b0 6
#286890000000
1!
1%
1-
12
#286900000000
0!
0%
b1 *
0-
02
b1 6
#286910000000
1!
1%
1-
12
#286920000000
0!
0%
b10 *
0-
02
b10 6
#286930000000
1!
1%
1-
12
#286940000000
0!
0%
b11 *
0-
02
b11 6
#286950000000
1!
1%
1-
12
15
#286960000000
0!
0%
b100 *
0-
02
b100 6
#286970000000
1!
1%
1-
12
#286980000000
0!
0%
b101 *
0-
02
b101 6
#286990000000
1!
1%
1-
12
#287000000000
0!
0%
b110 *
0-
02
b110 6
#287010000000
1!
1%
1-
12
#287020000000
0!
0%
b111 *
0-
02
b111 6
#287030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#287040000000
0!
0%
b0 *
0-
02
b0 6
#287050000000
1!
1%
1-
12
#287060000000
0!
0%
b1 *
0-
02
b1 6
#287070000000
1!
1%
1-
12
#287080000000
0!
0%
b10 *
0-
02
b10 6
#287090000000
1!
1%
1-
12
#287100000000
0!
0%
b11 *
0-
02
b11 6
#287110000000
1!
1%
1-
12
15
#287120000000
0!
0%
b100 *
0-
02
b100 6
#287130000000
1!
1%
1-
12
#287140000000
0!
0%
b101 *
0-
02
b101 6
#287150000000
1!
1%
1-
12
#287160000000
0!
0%
b110 *
0-
02
b110 6
#287170000000
1!
1%
1-
12
#287180000000
0!
0%
b111 *
0-
02
b111 6
#287190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#287200000000
0!
0%
b0 *
0-
02
b0 6
#287210000000
1!
1%
1-
12
#287220000000
0!
0%
b1 *
0-
02
b1 6
#287230000000
1!
1%
1-
12
#287240000000
0!
0%
b10 *
0-
02
b10 6
#287250000000
1!
1%
1-
12
#287260000000
0!
0%
b11 *
0-
02
b11 6
#287270000000
1!
1%
1-
12
15
#287280000000
0!
0%
b100 *
0-
02
b100 6
#287290000000
1!
1%
1-
12
#287300000000
0!
0%
b101 *
0-
02
b101 6
#287310000000
1!
1%
1-
12
#287320000000
0!
0%
b110 *
0-
02
b110 6
#287330000000
1!
1%
1-
12
#287340000000
0!
0%
b111 *
0-
02
b111 6
#287350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#287360000000
0!
0%
b0 *
0-
02
b0 6
#287370000000
1!
1%
1-
12
#287380000000
0!
0%
b1 *
0-
02
b1 6
#287390000000
1!
1%
1-
12
#287400000000
0!
0%
b10 *
0-
02
b10 6
#287410000000
1!
1%
1-
12
#287420000000
0!
0%
b11 *
0-
02
b11 6
#287430000000
1!
1%
1-
12
15
#287440000000
0!
0%
b100 *
0-
02
b100 6
#287450000000
1!
1%
1-
12
#287460000000
0!
0%
b101 *
0-
02
b101 6
#287470000000
1!
1%
1-
12
#287480000000
0!
0%
b110 *
0-
02
b110 6
#287490000000
1!
1%
1-
12
#287500000000
0!
0%
b111 *
0-
02
b111 6
#287510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#287520000000
0!
0%
b0 *
0-
02
b0 6
#287530000000
1!
1%
1-
12
#287540000000
0!
0%
b1 *
0-
02
b1 6
#287550000000
1!
1%
1-
12
#287560000000
0!
0%
b10 *
0-
02
b10 6
#287570000000
1!
1%
1-
12
#287580000000
0!
0%
b11 *
0-
02
b11 6
#287590000000
1!
1%
1-
12
15
#287600000000
0!
0%
b100 *
0-
02
b100 6
#287610000000
1!
1%
1-
12
#287620000000
0!
0%
b101 *
0-
02
b101 6
#287630000000
1!
1%
1-
12
#287640000000
0!
0%
b110 *
0-
02
b110 6
#287650000000
1!
1%
1-
12
#287660000000
0!
0%
b111 *
0-
02
b111 6
#287670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#287680000000
0!
0%
b0 *
0-
02
b0 6
#287690000000
1!
1%
1-
12
#287700000000
0!
0%
b1 *
0-
02
b1 6
#287710000000
1!
1%
1-
12
#287720000000
0!
0%
b10 *
0-
02
b10 6
#287730000000
1!
1%
1-
12
#287740000000
0!
0%
b11 *
0-
02
b11 6
#287750000000
1!
1%
1-
12
15
#287760000000
0!
0%
b100 *
0-
02
b100 6
#287770000000
1!
1%
1-
12
#287780000000
0!
0%
b101 *
0-
02
b101 6
#287790000000
1!
1%
1-
12
#287800000000
0!
0%
b110 *
0-
02
b110 6
#287810000000
1!
1%
1-
12
#287820000000
0!
0%
b111 *
0-
02
b111 6
#287830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#287840000000
0!
0%
b0 *
0-
02
b0 6
#287850000000
1!
1%
1-
12
#287860000000
0!
0%
b1 *
0-
02
b1 6
#287870000000
1!
1%
1-
12
#287880000000
0!
0%
b10 *
0-
02
b10 6
#287890000000
1!
1%
1-
12
#287900000000
0!
0%
b11 *
0-
02
b11 6
#287910000000
1!
1%
1-
12
15
#287920000000
0!
0%
b100 *
0-
02
b100 6
#287930000000
1!
1%
1-
12
#287940000000
0!
0%
b101 *
0-
02
b101 6
#287950000000
1!
1%
1-
12
#287960000000
0!
0%
b110 *
0-
02
b110 6
#287970000000
1!
1%
1-
12
#287980000000
0!
0%
b111 *
0-
02
b111 6
#287990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#288000000000
0!
0%
b0 *
0-
02
b0 6
#288010000000
1!
1%
1-
12
#288020000000
0!
0%
b1 *
0-
02
b1 6
#288030000000
1!
1%
1-
12
#288040000000
0!
0%
b10 *
0-
02
b10 6
#288050000000
1!
1%
1-
12
#288060000000
0!
0%
b11 *
0-
02
b11 6
#288070000000
1!
1%
1-
12
15
#288080000000
0!
0%
b100 *
0-
02
b100 6
#288090000000
1!
1%
1-
12
#288100000000
0!
0%
b101 *
0-
02
b101 6
#288110000000
1!
1%
1-
12
#288120000000
0!
0%
b110 *
0-
02
b110 6
#288130000000
1!
1%
1-
12
#288140000000
0!
0%
b111 *
0-
02
b111 6
#288150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#288160000000
0!
0%
b0 *
0-
02
b0 6
#288170000000
1!
1%
1-
12
#288180000000
0!
0%
b1 *
0-
02
b1 6
#288190000000
1!
1%
1-
12
#288200000000
0!
0%
b10 *
0-
02
b10 6
#288210000000
1!
1%
1-
12
#288220000000
0!
0%
b11 *
0-
02
b11 6
#288230000000
1!
1%
1-
12
15
#288240000000
0!
0%
b100 *
0-
02
b100 6
#288250000000
1!
1%
1-
12
#288260000000
0!
0%
b101 *
0-
02
b101 6
#288270000000
1!
1%
1-
12
#288280000000
0!
0%
b110 *
0-
02
b110 6
#288290000000
1!
1%
1-
12
#288300000000
0!
0%
b111 *
0-
02
b111 6
#288310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#288320000000
0!
0%
b0 *
0-
02
b0 6
#288330000000
1!
1%
1-
12
#288340000000
0!
0%
b1 *
0-
02
b1 6
#288350000000
1!
1%
1-
12
#288360000000
0!
0%
b10 *
0-
02
b10 6
#288370000000
1!
1%
1-
12
#288380000000
0!
0%
b11 *
0-
02
b11 6
#288390000000
1!
1%
1-
12
15
#288400000000
0!
0%
b100 *
0-
02
b100 6
#288410000000
1!
1%
1-
12
#288420000000
0!
0%
b101 *
0-
02
b101 6
#288430000000
1!
1%
1-
12
#288440000000
0!
0%
b110 *
0-
02
b110 6
#288450000000
1!
1%
1-
12
#288460000000
0!
0%
b111 *
0-
02
b111 6
#288470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#288480000000
0!
0%
b0 *
0-
02
b0 6
#288490000000
1!
1%
1-
12
#288500000000
0!
0%
b1 *
0-
02
b1 6
#288510000000
1!
1%
1-
12
#288520000000
0!
0%
b10 *
0-
02
b10 6
#288530000000
1!
1%
1-
12
#288540000000
0!
0%
b11 *
0-
02
b11 6
#288550000000
1!
1%
1-
12
15
#288560000000
0!
0%
b100 *
0-
02
b100 6
#288570000000
1!
1%
1-
12
#288580000000
0!
0%
b101 *
0-
02
b101 6
#288590000000
1!
1%
1-
12
#288600000000
0!
0%
b110 *
0-
02
b110 6
#288610000000
1!
1%
1-
12
#288620000000
0!
0%
b111 *
0-
02
b111 6
#288630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#288640000000
0!
0%
b0 *
0-
02
b0 6
#288650000000
1!
1%
1-
12
#288660000000
0!
0%
b1 *
0-
02
b1 6
#288670000000
1!
1%
1-
12
#288680000000
0!
0%
b10 *
0-
02
b10 6
#288690000000
1!
1%
1-
12
#288700000000
0!
0%
b11 *
0-
02
b11 6
#288710000000
1!
1%
1-
12
15
#288720000000
0!
0%
b100 *
0-
02
b100 6
#288730000000
1!
1%
1-
12
#288740000000
0!
0%
b101 *
0-
02
b101 6
#288750000000
1!
1%
1-
12
#288760000000
0!
0%
b110 *
0-
02
b110 6
#288770000000
1!
1%
1-
12
#288780000000
0!
0%
b111 *
0-
02
b111 6
#288790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#288800000000
0!
0%
b0 *
0-
02
b0 6
#288810000000
1!
1%
1-
12
#288820000000
0!
0%
b1 *
0-
02
b1 6
#288830000000
1!
1%
1-
12
#288840000000
0!
0%
b10 *
0-
02
b10 6
#288850000000
1!
1%
1-
12
#288860000000
0!
0%
b11 *
0-
02
b11 6
#288870000000
1!
1%
1-
12
15
#288880000000
0!
0%
b100 *
0-
02
b100 6
#288890000000
1!
1%
1-
12
#288900000000
0!
0%
b101 *
0-
02
b101 6
#288910000000
1!
1%
1-
12
#288920000000
0!
0%
b110 *
0-
02
b110 6
#288930000000
1!
1%
1-
12
#288940000000
0!
0%
b111 *
0-
02
b111 6
#288950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#288960000000
0!
0%
b0 *
0-
02
b0 6
#288970000000
1!
1%
1-
12
#288980000000
0!
0%
b1 *
0-
02
b1 6
#288990000000
1!
1%
1-
12
#289000000000
0!
0%
b10 *
0-
02
b10 6
#289010000000
1!
1%
1-
12
#289020000000
0!
0%
b11 *
0-
02
b11 6
#289030000000
1!
1%
1-
12
15
#289040000000
0!
0%
b100 *
0-
02
b100 6
#289050000000
1!
1%
1-
12
#289060000000
0!
0%
b101 *
0-
02
b101 6
#289070000000
1!
1%
1-
12
#289080000000
0!
0%
b110 *
0-
02
b110 6
#289090000000
1!
1%
1-
12
#289100000000
0!
0%
b111 *
0-
02
b111 6
#289110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#289120000000
0!
0%
b0 *
0-
02
b0 6
#289130000000
1!
1%
1-
12
#289140000000
0!
0%
b1 *
0-
02
b1 6
#289150000000
1!
1%
1-
12
#289160000000
0!
0%
b10 *
0-
02
b10 6
#289170000000
1!
1%
1-
12
#289180000000
0!
0%
b11 *
0-
02
b11 6
#289190000000
1!
1%
1-
12
15
#289200000000
0!
0%
b100 *
0-
02
b100 6
#289210000000
1!
1%
1-
12
#289220000000
0!
0%
b101 *
0-
02
b101 6
#289230000000
1!
1%
1-
12
#289240000000
0!
0%
b110 *
0-
02
b110 6
#289250000000
1!
1%
1-
12
#289260000000
0!
0%
b111 *
0-
02
b111 6
#289270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#289280000000
0!
0%
b0 *
0-
02
b0 6
#289290000000
1!
1%
1-
12
#289300000000
0!
0%
b1 *
0-
02
b1 6
#289310000000
1!
1%
1-
12
#289320000000
0!
0%
b10 *
0-
02
b10 6
#289330000000
1!
1%
1-
12
#289340000000
0!
0%
b11 *
0-
02
b11 6
#289350000000
1!
1%
1-
12
15
#289360000000
0!
0%
b100 *
0-
02
b100 6
#289370000000
1!
1%
1-
12
#289380000000
0!
0%
b101 *
0-
02
b101 6
#289390000000
1!
1%
1-
12
#289400000000
0!
0%
b110 *
0-
02
b110 6
#289410000000
1!
1%
1-
12
#289420000000
0!
0%
b111 *
0-
02
b111 6
#289430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#289440000000
0!
0%
b0 *
0-
02
b0 6
#289450000000
1!
1%
1-
12
#289460000000
0!
0%
b1 *
0-
02
b1 6
#289470000000
1!
1%
1-
12
#289480000000
0!
0%
b10 *
0-
02
b10 6
#289490000000
1!
1%
1-
12
#289500000000
0!
0%
b11 *
0-
02
b11 6
#289510000000
1!
1%
1-
12
15
#289520000000
0!
0%
b100 *
0-
02
b100 6
#289530000000
1!
1%
1-
12
#289540000000
0!
0%
b101 *
0-
02
b101 6
#289550000000
1!
1%
1-
12
#289560000000
0!
0%
b110 *
0-
02
b110 6
#289570000000
1!
1%
1-
12
#289580000000
0!
0%
b111 *
0-
02
b111 6
#289590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#289600000000
0!
0%
b0 *
0-
02
b0 6
#289610000000
1!
1%
1-
12
#289620000000
0!
0%
b1 *
0-
02
b1 6
#289630000000
1!
1%
1-
12
#289640000000
0!
0%
b10 *
0-
02
b10 6
#289650000000
1!
1%
1-
12
#289660000000
0!
0%
b11 *
0-
02
b11 6
#289670000000
1!
1%
1-
12
15
#289680000000
0!
0%
b100 *
0-
02
b100 6
#289690000000
1!
1%
1-
12
#289700000000
0!
0%
b101 *
0-
02
b101 6
#289710000000
1!
1%
1-
12
#289720000000
0!
0%
b110 *
0-
02
b110 6
#289730000000
1!
1%
1-
12
#289740000000
0!
0%
b111 *
0-
02
b111 6
#289750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#289760000000
0!
0%
b0 *
0-
02
b0 6
#289770000000
1!
1%
1-
12
#289780000000
0!
0%
b1 *
0-
02
b1 6
#289790000000
1!
1%
1-
12
#289800000000
0!
0%
b10 *
0-
02
b10 6
#289810000000
1!
1%
1-
12
#289820000000
0!
0%
b11 *
0-
02
b11 6
#289830000000
1!
1%
1-
12
15
#289840000000
0!
0%
b100 *
0-
02
b100 6
#289850000000
1!
1%
1-
12
#289860000000
0!
0%
b101 *
0-
02
b101 6
#289870000000
1!
1%
1-
12
#289880000000
0!
0%
b110 *
0-
02
b110 6
#289890000000
1!
1%
1-
12
#289900000000
0!
0%
b111 *
0-
02
b111 6
#289910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#289920000000
0!
0%
b0 *
0-
02
b0 6
#289930000000
1!
1%
1-
12
#289940000000
0!
0%
b1 *
0-
02
b1 6
#289950000000
1!
1%
1-
12
#289960000000
0!
0%
b10 *
0-
02
b10 6
#289970000000
1!
1%
1-
12
#289980000000
0!
0%
b11 *
0-
02
b11 6
#289990000000
1!
1%
1-
12
15
#290000000000
0!
0%
b100 *
0-
02
b100 6
#290010000000
1!
1%
1-
12
#290020000000
0!
0%
b101 *
0-
02
b101 6
#290030000000
1!
1%
1-
12
#290040000000
0!
0%
b110 *
0-
02
b110 6
#290050000000
1!
1%
1-
12
#290060000000
0!
0%
b111 *
0-
02
b111 6
#290070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#290080000000
0!
0%
b0 *
0-
02
b0 6
#290090000000
1!
1%
1-
12
#290100000000
0!
0%
b1 *
0-
02
b1 6
#290110000000
1!
1%
1-
12
#290120000000
0!
0%
b10 *
0-
02
b10 6
#290130000000
1!
1%
1-
12
#290140000000
0!
0%
b11 *
0-
02
b11 6
#290150000000
1!
1%
1-
12
15
#290160000000
0!
0%
b100 *
0-
02
b100 6
#290170000000
1!
1%
1-
12
#290180000000
0!
0%
b101 *
0-
02
b101 6
#290190000000
1!
1%
1-
12
#290200000000
0!
0%
b110 *
0-
02
b110 6
#290210000000
1!
1%
1-
12
#290220000000
0!
0%
b111 *
0-
02
b111 6
#290230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#290240000000
0!
0%
b0 *
0-
02
b0 6
#290250000000
1!
1%
1-
12
#290260000000
0!
0%
b1 *
0-
02
b1 6
#290270000000
1!
1%
1-
12
#290280000000
0!
0%
b10 *
0-
02
b10 6
#290290000000
1!
1%
1-
12
#290300000000
0!
0%
b11 *
0-
02
b11 6
#290310000000
1!
1%
1-
12
15
#290320000000
0!
0%
b100 *
0-
02
b100 6
#290330000000
1!
1%
1-
12
#290340000000
0!
0%
b101 *
0-
02
b101 6
#290350000000
1!
1%
1-
12
#290360000000
0!
0%
b110 *
0-
02
b110 6
#290370000000
1!
1%
1-
12
#290380000000
0!
0%
b111 *
0-
02
b111 6
#290390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#290400000000
0!
0%
b0 *
0-
02
b0 6
#290410000000
1!
1%
1-
12
#290420000000
0!
0%
b1 *
0-
02
b1 6
#290430000000
1!
1%
1-
12
#290440000000
0!
0%
b10 *
0-
02
b10 6
#290450000000
1!
1%
1-
12
#290460000000
0!
0%
b11 *
0-
02
b11 6
#290470000000
1!
1%
1-
12
15
#290480000000
0!
0%
b100 *
0-
02
b100 6
#290490000000
1!
1%
1-
12
#290500000000
0!
0%
b101 *
0-
02
b101 6
#290510000000
1!
1%
1-
12
#290520000000
0!
0%
b110 *
0-
02
b110 6
#290530000000
1!
1%
1-
12
#290540000000
0!
0%
b111 *
0-
02
b111 6
#290550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#290560000000
0!
0%
b0 *
0-
02
b0 6
#290570000000
1!
1%
1-
12
#290580000000
0!
0%
b1 *
0-
02
b1 6
#290590000000
1!
1%
1-
12
#290600000000
0!
0%
b10 *
0-
02
b10 6
#290610000000
1!
1%
1-
12
#290620000000
0!
0%
b11 *
0-
02
b11 6
#290630000000
1!
1%
1-
12
15
#290640000000
0!
0%
b100 *
0-
02
b100 6
#290650000000
1!
1%
1-
12
#290660000000
0!
0%
b101 *
0-
02
b101 6
#290670000000
1!
1%
1-
12
#290680000000
0!
0%
b110 *
0-
02
b110 6
#290690000000
1!
1%
1-
12
#290700000000
0!
0%
b111 *
0-
02
b111 6
#290710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#290720000000
0!
0%
b0 *
0-
02
b0 6
#290730000000
1!
1%
1-
12
#290740000000
0!
0%
b1 *
0-
02
b1 6
#290750000000
1!
1%
1-
12
#290760000000
0!
0%
b10 *
0-
02
b10 6
#290770000000
1!
1%
1-
12
#290780000000
0!
0%
b11 *
0-
02
b11 6
#290790000000
1!
1%
1-
12
15
#290800000000
0!
0%
b100 *
0-
02
b100 6
#290810000000
1!
1%
1-
12
#290820000000
0!
0%
b101 *
0-
02
b101 6
#290830000000
1!
1%
1-
12
#290840000000
0!
0%
b110 *
0-
02
b110 6
#290850000000
1!
1%
1-
12
#290860000000
0!
0%
b111 *
0-
02
b111 6
#290870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#290880000000
0!
0%
b0 *
0-
02
b0 6
#290890000000
1!
1%
1-
12
#290900000000
0!
0%
b1 *
0-
02
b1 6
#290910000000
1!
1%
1-
12
#290920000000
0!
0%
b10 *
0-
02
b10 6
#290930000000
1!
1%
1-
12
#290940000000
0!
0%
b11 *
0-
02
b11 6
#290950000000
1!
1%
1-
12
15
#290960000000
0!
0%
b100 *
0-
02
b100 6
#290970000000
1!
1%
1-
12
#290980000000
0!
0%
b101 *
0-
02
b101 6
#290990000000
1!
1%
1-
12
#291000000000
0!
0%
b110 *
0-
02
b110 6
#291010000000
1!
1%
1-
12
#291020000000
0!
0%
b111 *
0-
02
b111 6
#291030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#291040000000
0!
0%
b0 *
0-
02
b0 6
#291050000000
1!
1%
1-
12
#291060000000
0!
0%
b1 *
0-
02
b1 6
#291070000000
1!
1%
1-
12
#291080000000
0!
0%
b10 *
0-
02
b10 6
#291090000000
1!
1%
1-
12
#291100000000
0!
0%
b11 *
0-
02
b11 6
#291110000000
1!
1%
1-
12
15
#291120000000
0!
0%
b100 *
0-
02
b100 6
#291130000000
1!
1%
1-
12
#291140000000
0!
0%
b101 *
0-
02
b101 6
#291150000000
1!
1%
1-
12
#291160000000
0!
0%
b110 *
0-
02
b110 6
#291170000000
1!
1%
1-
12
#291180000000
0!
0%
b111 *
0-
02
b111 6
#291190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#291200000000
0!
0%
b0 *
0-
02
b0 6
#291210000000
1!
1%
1-
12
#291220000000
0!
0%
b1 *
0-
02
b1 6
#291230000000
1!
1%
1-
12
#291240000000
0!
0%
b10 *
0-
02
b10 6
#291250000000
1!
1%
1-
12
#291260000000
0!
0%
b11 *
0-
02
b11 6
#291270000000
1!
1%
1-
12
15
#291280000000
0!
0%
b100 *
0-
02
b100 6
#291290000000
1!
1%
1-
12
#291300000000
0!
0%
b101 *
0-
02
b101 6
#291310000000
1!
1%
1-
12
#291320000000
0!
0%
b110 *
0-
02
b110 6
#291330000000
1!
1%
1-
12
#291340000000
0!
0%
b111 *
0-
02
b111 6
#291350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#291360000000
0!
0%
b0 *
0-
02
b0 6
#291370000000
1!
1%
1-
12
#291380000000
0!
0%
b1 *
0-
02
b1 6
#291390000000
1!
1%
1-
12
#291400000000
0!
0%
b10 *
0-
02
b10 6
#291410000000
1!
1%
1-
12
#291420000000
0!
0%
b11 *
0-
02
b11 6
#291430000000
1!
1%
1-
12
15
#291440000000
0!
0%
b100 *
0-
02
b100 6
#291450000000
1!
1%
1-
12
#291460000000
0!
0%
b101 *
0-
02
b101 6
#291470000000
1!
1%
1-
12
#291480000000
0!
0%
b110 *
0-
02
b110 6
#291490000000
1!
1%
1-
12
#291500000000
0!
0%
b111 *
0-
02
b111 6
#291510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#291520000000
0!
0%
b0 *
0-
02
b0 6
#291530000000
1!
1%
1-
12
#291540000000
0!
0%
b1 *
0-
02
b1 6
#291550000000
1!
1%
1-
12
#291560000000
0!
0%
b10 *
0-
02
b10 6
#291570000000
1!
1%
1-
12
#291580000000
0!
0%
b11 *
0-
02
b11 6
#291590000000
1!
1%
1-
12
15
#291600000000
0!
0%
b100 *
0-
02
b100 6
#291610000000
1!
1%
1-
12
#291620000000
0!
0%
b101 *
0-
02
b101 6
#291630000000
1!
1%
1-
12
#291640000000
0!
0%
b110 *
0-
02
b110 6
#291650000000
1!
1%
1-
12
#291660000000
0!
0%
b111 *
0-
02
b111 6
#291670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#291680000000
0!
0%
b0 *
0-
02
b0 6
#291690000000
1!
1%
1-
12
#291700000000
0!
0%
b1 *
0-
02
b1 6
#291710000000
1!
1%
1-
12
#291720000000
0!
0%
b10 *
0-
02
b10 6
#291730000000
1!
1%
1-
12
#291740000000
0!
0%
b11 *
0-
02
b11 6
#291750000000
1!
1%
1-
12
15
#291760000000
0!
0%
b100 *
0-
02
b100 6
#291770000000
1!
1%
1-
12
#291780000000
0!
0%
b101 *
0-
02
b101 6
#291790000000
1!
1%
1-
12
#291800000000
0!
0%
b110 *
0-
02
b110 6
#291810000000
1!
1%
1-
12
#291820000000
0!
0%
b111 *
0-
02
b111 6
#291830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#291840000000
0!
0%
b0 *
0-
02
b0 6
#291850000000
1!
1%
1-
12
#291860000000
0!
0%
b1 *
0-
02
b1 6
#291870000000
1!
1%
1-
12
#291880000000
0!
0%
b10 *
0-
02
b10 6
#291890000000
1!
1%
1-
12
#291900000000
0!
0%
b11 *
0-
02
b11 6
#291910000000
1!
1%
1-
12
15
#291920000000
0!
0%
b100 *
0-
02
b100 6
#291930000000
1!
1%
1-
12
#291940000000
0!
0%
b101 *
0-
02
b101 6
#291950000000
1!
1%
1-
12
#291960000000
0!
0%
b110 *
0-
02
b110 6
#291970000000
1!
1%
1-
12
#291980000000
0!
0%
b111 *
0-
02
b111 6
#291990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#292000000000
0!
0%
b0 *
0-
02
b0 6
#292010000000
1!
1%
1-
12
#292020000000
0!
0%
b1 *
0-
02
b1 6
#292030000000
1!
1%
1-
12
#292040000000
0!
0%
b10 *
0-
02
b10 6
#292050000000
1!
1%
1-
12
#292060000000
0!
0%
b11 *
0-
02
b11 6
#292070000000
1!
1%
1-
12
15
#292080000000
0!
0%
b100 *
0-
02
b100 6
#292090000000
1!
1%
1-
12
#292100000000
0!
0%
b101 *
0-
02
b101 6
#292110000000
1!
1%
1-
12
#292120000000
0!
0%
b110 *
0-
02
b110 6
#292130000000
1!
1%
1-
12
#292140000000
0!
0%
b111 *
0-
02
b111 6
#292150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#292160000000
0!
0%
b0 *
0-
02
b0 6
#292170000000
1!
1%
1-
12
#292180000000
0!
0%
b1 *
0-
02
b1 6
#292190000000
1!
1%
1-
12
#292200000000
0!
0%
b10 *
0-
02
b10 6
#292210000000
1!
1%
1-
12
#292220000000
0!
0%
b11 *
0-
02
b11 6
#292230000000
1!
1%
1-
12
15
#292240000000
0!
0%
b100 *
0-
02
b100 6
#292250000000
1!
1%
1-
12
#292260000000
0!
0%
b101 *
0-
02
b101 6
#292270000000
1!
1%
1-
12
#292280000000
0!
0%
b110 *
0-
02
b110 6
#292290000000
1!
1%
1-
12
#292300000000
0!
0%
b111 *
0-
02
b111 6
#292310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#292320000000
0!
0%
b0 *
0-
02
b0 6
#292330000000
1!
1%
1-
12
#292340000000
0!
0%
b1 *
0-
02
b1 6
#292350000000
1!
1%
1-
12
#292360000000
0!
0%
b10 *
0-
02
b10 6
#292370000000
1!
1%
1-
12
#292380000000
0!
0%
b11 *
0-
02
b11 6
#292390000000
1!
1%
1-
12
15
#292400000000
0!
0%
b100 *
0-
02
b100 6
#292410000000
1!
1%
1-
12
#292420000000
0!
0%
b101 *
0-
02
b101 6
#292430000000
1!
1%
1-
12
#292440000000
0!
0%
b110 *
0-
02
b110 6
#292450000000
1!
1%
1-
12
#292460000000
0!
0%
b111 *
0-
02
b111 6
#292470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#292480000000
0!
0%
b0 *
0-
02
b0 6
#292490000000
1!
1%
1-
12
#292500000000
0!
0%
b1 *
0-
02
b1 6
#292510000000
1!
1%
1-
12
#292520000000
0!
0%
b10 *
0-
02
b10 6
#292530000000
1!
1%
1-
12
#292540000000
0!
0%
b11 *
0-
02
b11 6
#292550000000
1!
1%
1-
12
15
#292560000000
0!
0%
b100 *
0-
02
b100 6
#292570000000
1!
1%
1-
12
#292580000000
0!
0%
b101 *
0-
02
b101 6
#292590000000
1!
1%
1-
12
#292600000000
0!
0%
b110 *
0-
02
b110 6
#292610000000
1!
1%
1-
12
#292620000000
0!
0%
b111 *
0-
02
b111 6
#292630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#292640000000
0!
0%
b0 *
0-
02
b0 6
#292650000000
1!
1%
1-
12
#292660000000
0!
0%
b1 *
0-
02
b1 6
#292670000000
1!
1%
1-
12
#292680000000
0!
0%
b10 *
0-
02
b10 6
#292690000000
1!
1%
1-
12
#292700000000
0!
0%
b11 *
0-
02
b11 6
#292710000000
1!
1%
1-
12
15
#292720000000
0!
0%
b100 *
0-
02
b100 6
#292730000000
1!
1%
1-
12
#292740000000
0!
0%
b101 *
0-
02
b101 6
#292750000000
1!
1%
1-
12
#292760000000
0!
0%
b110 *
0-
02
b110 6
#292770000000
1!
1%
1-
12
#292780000000
0!
0%
b111 *
0-
02
b111 6
#292790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#292800000000
0!
0%
b0 *
0-
02
b0 6
#292810000000
1!
1%
1-
12
#292820000000
0!
0%
b1 *
0-
02
b1 6
#292830000000
1!
1%
1-
12
#292840000000
0!
0%
b10 *
0-
02
b10 6
#292850000000
1!
1%
1-
12
#292860000000
0!
0%
b11 *
0-
02
b11 6
#292870000000
1!
1%
1-
12
15
#292880000000
0!
0%
b100 *
0-
02
b100 6
#292890000000
1!
1%
1-
12
#292900000000
0!
0%
b101 *
0-
02
b101 6
#292910000000
1!
1%
1-
12
#292920000000
0!
0%
b110 *
0-
02
b110 6
#292930000000
1!
1%
1-
12
#292940000000
0!
0%
b111 *
0-
02
b111 6
#292950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#292960000000
0!
0%
b0 *
0-
02
b0 6
#292970000000
1!
1%
1-
12
#292980000000
0!
0%
b1 *
0-
02
b1 6
#292990000000
1!
1%
1-
12
#293000000000
0!
0%
b10 *
0-
02
b10 6
#293010000000
1!
1%
1-
12
#293020000000
0!
0%
b11 *
0-
02
b11 6
#293030000000
1!
1%
1-
12
15
#293040000000
0!
0%
b100 *
0-
02
b100 6
#293050000000
1!
1%
1-
12
#293060000000
0!
0%
b101 *
0-
02
b101 6
#293070000000
1!
1%
1-
12
#293080000000
0!
0%
b110 *
0-
02
b110 6
#293090000000
1!
1%
1-
12
#293100000000
0!
0%
b111 *
0-
02
b111 6
#293110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#293120000000
0!
0%
b0 *
0-
02
b0 6
#293130000000
1!
1%
1-
12
#293140000000
0!
0%
b1 *
0-
02
b1 6
#293150000000
1!
1%
1-
12
#293160000000
0!
0%
b10 *
0-
02
b10 6
#293170000000
1!
1%
1-
12
#293180000000
0!
0%
b11 *
0-
02
b11 6
#293190000000
1!
1%
1-
12
15
#293200000000
0!
0%
b100 *
0-
02
b100 6
#293210000000
1!
1%
1-
12
#293220000000
0!
0%
b101 *
0-
02
b101 6
#293230000000
1!
1%
1-
12
#293240000000
0!
0%
b110 *
0-
02
b110 6
#293250000000
1!
1%
1-
12
#293260000000
0!
0%
b111 *
0-
02
b111 6
#293270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#293280000000
0!
0%
b0 *
0-
02
b0 6
#293290000000
1!
1%
1-
12
#293300000000
0!
0%
b1 *
0-
02
b1 6
#293310000000
1!
1%
1-
12
#293320000000
0!
0%
b10 *
0-
02
b10 6
#293330000000
1!
1%
1-
12
#293340000000
0!
0%
b11 *
0-
02
b11 6
#293350000000
1!
1%
1-
12
15
#293360000000
0!
0%
b100 *
0-
02
b100 6
#293370000000
1!
1%
1-
12
#293380000000
0!
0%
b101 *
0-
02
b101 6
#293390000000
1!
1%
1-
12
#293400000000
0!
0%
b110 *
0-
02
b110 6
#293410000000
1!
1%
1-
12
#293420000000
0!
0%
b111 *
0-
02
b111 6
#293430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#293440000000
0!
0%
b0 *
0-
02
b0 6
#293450000000
1!
1%
1-
12
#293460000000
0!
0%
b1 *
0-
02
b1 6
#293470000000
1!
1%
1-
12
#293480000000
0!
0%
b10 *
0-
02
b10 6
#293490000000
1!
1%
1-
12
#293500000000
0!
0%
b11 *
0-
02
b11 6
#293510000000
1!
1%
1-
12
15
#293520000000
0!
0%
b100 *
0-
02
b100 6
#293530000000
1!
1%
1-
12
#293540000000
0!
0%
b101 *
0-
02
b101 6
#293550000000
1!
1%
1-
12
#293560000000
0!
0%
b110 *
0-
02
b110 6
#293570000000
1!
1%
1-
12
#293580000000
0!
0%
b111 *
0-
02
b111 6
#293590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#293600000000
0!
0%
b0 *
0-
02
b0 6
#293610000000
1!
1%
1-
12
#293620000000
0!
0%
b1 *
0-
02
b1 6
#293630000000
1!
1%
1-
12
#293640000000
0!
0%
b10 *
0-
02
b10 6
#293650000000
1!
1%
1-
12
#293660000000
0!
0%
b11 *
0-
02
b11 6
#293670000000
1!
1%
1-
12
15
#293680000000
0!
0%
b100 *
0-
02
b100 6
#293690000000
1!
1%
1-
12
#293700000000
0!
0%
b101 *
0-
02
b101 6
#293710000000
1!
1%
1-
12
#293720000000
0!
0%
b110 *
0-
02
b110 6
#293730000000
1!
1%
1-
12
#293740000000
0!
0%
b111 *
0-
02
b111 6
#293750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#293760000000
0!
0%
b0 *
0-
02
b0 6
#293770000000
1!
1%
1-
12
#293780000000
0!
0%
b1 *
0-
02
b1 6
#293790000000
1!
1%
1-
12
#293800000000
0!
0%
b10 *
0-
02
b10 6
#293810000000
1!
1%
1-
12
#293820000000
0!
0%
b11 *
0-
02
b11 6
#293830000000
1!
1%
1-
12
15
#293840000000
0!
0%
b100 *
0-
02
b100 6
#293850000000
1!
1%
1-
12
#293860000000
0!
0%
b101 *
0-
02
b101 6
#293870000000
1!
1%
1-
12
#293880000000
0!
0%
b110 *
0-
02
b110 6
#293890000000
1!
1%
1-
12
#293900000000
0!
0%
b111 *
0-
02
b111 6
#293910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#293920000000
0!
0%
b0 *
0-
02
b0 6
#293930000000
1!
1%
1-
12
#293940000000
0!
0%
b1 *
0-
02
b1 6
#293950000000
1!
1%
1-
12
#293960000000
0!
0%
b10 *
0-
02
b10 6
#293970000000
1!
1%
1-
12
#293980000000
0!
0%
b11 *
0-
02
b11 6
#293990000000
1!
1%
1-
12
15
#294000000000
0!
0%
b100 *
0-
02
b100 6
#294010000000
1!
1%
1-
12
#294020000000
0!
0%
b101 *
0-
02
b101 6
#294030000000
1!
1%
1-
12
#294040000000
0!
0%
b110 *
0-
02
b110 6
#294050000000
1!
1%
1-
12
#294060000000
0!
0%
b111 *
0-
02
b111 6
#294070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#294080000000
0!
0%
b0 *
0-
02
b0 6
#294090000000
1!
1%
1-
12
#294100000000
0!
0%
b1 *
0-
02
b1 6
#294110000000
1!
1%
1-
12
#294120000000
0!
0%
b10 *
0-
02
b10 6
#294130000000
1!
1%
1-
12
#294140000000
0!
0%
b11 *
0-
02
b11 6
#294150000000
1!
1%
1-
12
15
#294160000000
0!
0%
b100 *
0-
02
b100 6
#294170000000
1!
1%
1-
12
#294180000000
0!
0%
b101 *
0-
02
b101 6
#294190000000
1!
1%
1-
12
#294200000000
0!
0%
b110 *
0-
02
b110 6
#294210000000
1!
1%
1-
12
#294220000000
0!
0%
b111 *
0-
02
b111 6
#294230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#294240000000
0!
0%
b0 *
0-
02
b0 6
#294250000000
1!
1%
1-
12
#294260000000
0!
0%
b1 *
0-
02
b1 6
#294270000000
1!
1%
1-
12
#294280000000
0!
0%
b10 *
0-
02
b10 6
#294290000000
1!
1%
1-
12
#294300000000
0!
0%
b11 *
0-
02
b11 6
#294310000000
1!
1%
1-
12
15
#294320000000
0!
0%
b100 *
0-
02
b100 6
#294330000000
1!
1%
1-
12
#294340000000
0!
0%
b101 *
0-
02
b101 6
#294350000000
1!
1%
1-
12
#294360000000
0!
0%
b110 *
0-
02
b110 6
#294370000000
1!
1%
1-
12
#294380000000
0!
0%
b111 *
0-
02
b111 6
#294390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#294400000000
0!
0%
b0 *
0-
02
b0 6
#294410000000
1!
1%
1-
12
#294420000000
0!
0%
b1 *
0-
02
b1 6
#294430000000
1!
1%
1-
12
#294440000000
0!
0%
b10 *
0-
02
b10 6
#294450000000
1!
1%
1-
12
#294460000000
0!
0%
b11 *
0-
02
b11 6
#294470000000
1!
1%
1-
12
15
#294480000000
0!
0%
b100 *
0-
02
b100 6
#294490000000
1!
1%
1-
12
#294500000000
0!
0%
b101 *
0-
02
b101 6
#294510000000
1!
1%
1-
12
#294520000000
0!
0%
b110 *
0-
02
b110 6
#294530000000
1!
1%
1-
12
#294540000000
0!
0%
b111 *
0-
02
b111 6
#294550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#294560000000
0!
0%
b0 *
0-
02
b0 6
#294570000000
1!
1%
1-
12
#294580000000
0!
0%
b1 *
0-
02
b1 6
#294590000000
1!
1%
1-
12
#294600000000
0!
0%
b10 *
0-
02
b10 6
#294610000000
1!
1%
1-
12
#294620000000
0!
0%
b11 *
0-
02
b11 6
#294630000000
1!
1%
1-
12
15
#294640000000
0!
0%
b100 *
0-
02
b100 6
#294650000000
1!
1%
1-
12
#294660000000
0!
0%
b101 *
0-
02
b101 6
#294670000000
1!
1%
1-
12
#294680000000
0!
0%
b110 *
0-
02
b110 6
#294690000000
1!
1%
1-
12
#294700000000
0!
0%
b111 *
0-
02
b111 6
#294710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#294720000000
0!
0%
b0 *
0-
02
b0 6
#294730000000
1!
1%
1-
12
#294740000000
0!
0%
b1 *
0-
02
b1 6
#294750000000
1!
1%
1-
12
#294760000000
0!
0%
b10 *
0-
02
b10 6
#294770000000
1!
1%
1-
12
#294780000000
0!
0%
b11 *
0-
02
b11 6
#294790000000
1!
1%
1-
12
15
#294800000000
0!
0%
b100 *
0-
02
b100 6
#294810000000
1!
1%
1-
12
#294820000000
0!
0%
b101 *
0-
02
b101 6
#294830000000
1!
1%
1-
12
#294840000000
0!
0%
b110 *
0-
02
b110 6
#294850000000
1!
1%
1-
12
#294860000000
0!
0%
b111 *
0-
02
b111 6
#294870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#294880000000
0!
0%
b0 *
0-
02
b0 6
#294890000000
1!
1%
1-
12
#294900000000
0!
0%
b1 *
0-
02
b1 6
#294910000000
1!
1%
1-
12
#294920000000
0!
0%
b10 *
0-
02
b10 6
#294930000000
1!
1%
1-
12
#294940000000
0!
0%
b11 *
0-
02
b11 6
#294950000000
1!
1%
1-
12
15
#294960000000
0!
0%
b100 *
0-
02
b100 6
#294970000000
1!
1%
1-
12
#294980000000
0!
0%
b101 *
0-
02
b101 6
#294990000000
1!
1%
1-
12
#295000000000
0!
0%
b110 *
0-
02
b110 6
#295010000000
1!
1%
1-
12
#295020000000
0!
0%
b111 *
0-
02
b111 6
#295030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#295040000000
0!
0%
b0 *
0-
02
b0 6
#295050000000
1!
1%
1-
12
#295060000000
0!
0%
b1 *
0-
02
b1 6
#295070000000
1!
1%
1-
12
#295080000000
0!
0%
b10 *
0-
02
b10 6
#295090000000
1!
1%
1-
12
#295100000000
0!
0%
b11 *
0-
02
b11 6
#295110000000
1!
1%
1-
12
15
#295120000000
0!
0%
b100 *
0-
02
b100 6
#295130000000
1!
1%
1-
12
#295140000000
0!
0%
b101 *
0-
02
b101 6
#295150000000
1!
1%
1-
12
#295160000000
0!
0%
b110 *
0-
02
b110 6
#295170000000
1!
1%
1-
12
#295180000000
0!
0%
b111 *
0-
02
b111 6
#295190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#295200000000
0!
0%
b0 *
0-
02
b0 6
#295210000000
1!
1%
1-
12
#295220000000
0!
0%
b1 *
0-
02
b1 6
#295230000000
1!
1%
1-
12
#295240000000
0!
0%
b10 *
0-
02
b10 6
#295250000000
1!
1%
1-
12
#295260000000
0!
0%
b11 *
0-
02
b11 6
#295270000000
1!
1%
1-
12
15
#295280000000
0!
0%
b100 *
0-
02
b100 6
#295290000000
1!
1%
1-
12
#295300000000
0!
0%
b101 *
0-
02
b101 6
#295310000000
1!
1%
1-
12
#295320000000
0!
0%
b110 *
0-
02
b110 6
#295330000000
1!
1%
1-
12
#295340000000
0!
0%
b111 *
0-
02
b111 6
#295350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#295360000000
0!
0%
b0 *
0-
02
b0 6
#295370000000
1!
1%
1-
12
#295380000000
0!
0%
b1 *
0-
02
b1 6
#295390000000
1!
1%
1-
12
#295400000000
0!
0%
b10 *
0-
02
b10 6
#295410000000
1!
1%
1-
12
#295420000000
0!
0%
b11 *
0-
02
b11 6
#295430000000
1!
1%
1-
12
15
#295440000000
0!
0%
b100 *
0-
02
b100 6
#295450000000
1!
1%
1-
12
#295460000000
0!
0%
b101 *
0-
02
b101 6
#295470000000
1!
1%
1-
12
#295480000000
0!
0%
b110 *
0-
02
b110 6
#295490000000
1!
1%
1-
12
#295500000000
0!
0%
b111 *
0-
02
b111 6
#295510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#295520000000
0!
0%
b0 *
0-
02
b0 6
#295530000000
1!
1%
1-
12
#295540000000
0!
0%
b1 *
0-
02
b1 6
#295550000000
1!
1%
1-
12
#295560000000
0!
0%
b10 *
0-
02
b10 6
#295570000000
1!
1%
1-
12
#295580000000
0!
0%
b11 *
0-
02
b11 6
#295590000000
1!
1%
1-
12
15
#295600000000
0!
0%
b100 *
0-
02
b100 6
#295610000000
1!
1%
1-
12
#295620000000
0!
0%
b101 *
0-
02
b101 6
#295630000000
1!
1%
1-
12
#295640000000
0!
0%
b110 *
0-
02
b110 6
#295650000000
1!
1%
1-
12
#295660000000
0!
0%
b111 *
0-
02
b111 6
#295670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#295680000000
0!
0%
b0 *
0-
02
b0 6
#295690000000
1!
1%
1-
12
#295700000000
0!
0%
b1 *
0-
02
b1 6
#295710000000
1!
1%
1-
12
#295720000000
0!
0%
b10 *
0-
02
b10 6
#295730000000
1!
1%
1-
12
#295740000000
0!
0%
b11 *
0-
02
b11 6
#295750000000
1!
1%
1-
12
15
#295760000000
0!
0%
b100 *
0-
02
b100 6
#295770000000
1!
1%
1-
12
#295780000000
0!
0%
b101 *
0-
02
b101 6
#295790000000
1!
1%
1-
12
#295800000000
0!
0%
b110 *
0-
02
b110 6
#295810000000
1!
1%
1-
12
#295820000000
0!
0%
b111 *
0-
02
b111 6
#295830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#295840000000
0!
0%
b0 *
0-
02
b0 6
#295850000000
1!
1%
1-
12
#295860000000
0!
0%
b1 *
0-
02
b1 6
#295870000000
1!
1%
1-
12
#295880000000
0!
0%
b10 *
0-
02
b10 6
#295890000000
1!
1%
1-
12
#295900000000
0!
0%
b11 *
0-
02
b11 6
#295910000000
1!
1%
1-
12
15
#295920000000
0!
0%
b100 *
0-
02
b100 6
#295930000000
1!
1%
1-
12
#295940000000
0!
0%
b101 *
0-
02
b101 6
#295950000000
1!
1%
1-
12
#295960000000
0!
0%
b110 *
0-
02
b110 6
#295970000000
1!
1%
1-
12
#295980000000
0!
0%
b111 *
0-
02
b111 6
#295990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#296000000000
0!
0%
b0 *
0-
02
b0 6
#296010000000
1!
1%
1-
12
#296020000000
0!
0%
b1 *
0-
02
b1 6
#296030000000
1!
1%
1-
12
#296040000000
0!
0%
b10 *
0-
02
b10 6
#296050000000
1!
1%
1-
12
#296060000000
0!
0%
b11 *
0-
02
b11 6
#296070000000
1!
1%
1-
12
15
#296080000000
0!
0%
b100 *
0-
02
b100 6
#296090000000
1!
1%
1-
12
#296100000000
0!
0%
b101 *
0-
02
b101 6
#296110000000
1!
1%
1-
12
#296120000000
0!
0%
b110 *
0-
02
b110 6
#296130000000
1!
1%
1-
12
#296140000000
0!
0%
b111 *
0-
02
b111 6
#296150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#296160000000
0!
0%
b0 *
0-
02
b0 6
#296170000000
1!
1%
1-
12
#296180000000
0!
0%
b1 *
0-
02
b1 6
#296190000000
1!
1%
1-
12
#296200000000
0!
0%
b10 *
0-
02
b10 6
#296210000000
1!
1%
1-
12
#296220000000
0!
0%
b11 *
0-
02
b11 6
#296230000000
1!
1%
1-
12
15
#296240000000
0!
0%
b100 *
0-
02
b100 6
#296250000000
1!
1%
1-
12
#296260000000
0!
0%
b101 *
0-
02
b101 6
#296270000000
1!
1%
1-
12
#296280000000
0!
0%
b110 *
0-
02
b110 6
#296290000000
1!
1%
1-
12
#296300000000
0!
0%
b111 *
0-
02
b111 6
#296310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#296320000000
0!
0%
b0 *
0-
02
b0 6
#296330000000
1!
1%
1-
12
#296340000000
0!
0%
b1 *
0-
02
b1 6
#296350000000
1!
1%
1-
12
#296360000000
0!
0%
b10 *
0-
02
b10 6
#296370000000
1!
1%
1-
12
#296380000000
0!
0%
b11 *
0-
02
b11 6
#296390000000
1!
1%
1-
12
15
#296400000000
0!
0%
b100 *
0-
02
b100 6
#296410000000
1!
1%
1-
12
#296420000000
0!
0%
b101 *
0-
02
b101 6
#296430000000
1!
1%
1-
12
#296440000000
0!
0%
b110 *
0-
02
b110 6
#296450000000
1!
1%
1-
12
#296460000000
0!
0%
b111 *
0-
02
b111 6
#296470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#296480000000
0!
0%
b0 *
0-
02
b0 6
#296490000000
1!
1%
1-
12
#296500000000
0!
0%
b1 *
0-
02
b1 6
#296510000000
1!
1%
1-
12
#296520000000
0!
0%
b10 *
0-
02
b10 6
#296530000000
1!
1%
1-
12
#296540000000
0!
0%
b11 *
0-
02
b11 6
#296550000000
1!
1%
1-
12
15
#296560000000
0!
0%
b100 *
0-
02
b100 6
#296570000000
1!
1%
1-
12
#296580000000
0!
0%
b101 *
0-
02
b101 6
#296590000000
1!
1%
1-
12
#296600000000
0!
0%
b110 *
0-
02
b110 6
#296610000000
1!
1%
1-
12
#296620000000
0!
0%
b111 *
0-
02
b111 6
#296630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#296640000000
0!
0%
b0 *
0-
02
b0 6
#296650000000
1!
1%
1-
12
#296660000000
0!
0%
b1 *
0-
02
b1 6
#296670000000
1!
1%
1-
12
#296680000000
0!
0%
b10 *
0-
02
b10 6
#296690000000
1!
1%
1-
12
#296700000000
0!
0%
b11 *
0-
02
b11 6
#296710000000
1!
1%
1-
12
15
#296720000000
0!
0%
b100 *
0-
02
b100 6
#296730000000
1!
1%
1-
12
#296740000000
0!
0%
b101 *
0-
02
b101 6
#296750000000
1!
1%
1-
12
#296760000000
0!
0%
b110 *
0-
02
b110 6
#296770000000
1!
1%
1-
12
#296780000000
0!
0%
b111 *
0-
02
b111 6
#296790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#296800000000
0!
0%
b0 *
0-
02
b0 6
#296810000000
1!
1%
1-
12
#296820000000
0!
0%
b1 *
0-
02
b1 6
#296830000000
1!
1%
1-
12
#296840000000
0!
0%
b10 *
0-
02
b10 6
#296850000000
1!
1%
1-
12
#296860000000
0!
0%
b11 *
0-
02
b11 6
#296870000000
1!
1%
1-
12
15
#296880000000
0!
0%
b100 *
0-
02
b100 6
#296890000000
1!
1%
1-
12
#296900000000
0!
0%
b101 *
0-
02
b101 6
#296910000000
1!
1%
1-
12
#296920000000
0!
0%
b110 *
0-
02
b110 6
#296930000000
1!
1%
1-
12
#296940000000
0!
0%
b111 *
0-
02
b111 6
#296950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#296960000000
0!
0%
b0 *
0-
02
b0 6
#296970000000
1!
1%
1-
12
#296980000000
0!
0%
b1 *
0-
02
b1 6
#296990000000
1!
1%
1-
12
#297000000000
0!
0%
b10 *
0-
02
b10 6
#297010000000
1!
1%
1-
12
#297020000000
0!
0%
b11 *
0-
02
b11 6
#297030000000
1!
1%
1-
12
15
#297040000000
0!
0%
b100 *
0-
02
b100 6
#297050000000
1!
1%
1-
12
#297060000000
0!
0%
b101 *
0-
02
b101 6
#297070000000
1!
1%
1-
12
#297080000000
0!
0%
b110 *
0-
02
b110 6
#297090000000
1!
1%
1-
12
#297100000000
0!
0%
b111 *
0-
02
b111 6
#297110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#297120000000
0!
0%
b0 *
0-
02
b0 6
#297130000000
1!
1%
1-
12
#297140000000
0!
0%
b1 *
0-
02
b1 6
#297150000000
1!
1%
1-
12
#297160000000
0!
0%
b10 *
0-
02
b10 6
#297170000000
1!
1%
1-
12
#297180000000
0!
0%
b11 *
0-
02
b11 6
#297190000000
1!
1%
1-
12
15
#297200000000
0!
0%
b100 *
0-
02
b100 6
#297210000000
1!
1%
1-
12
#297220000000
0!
0%
b101 *
0-
02
b101 6
#297230000000
1!
1%
1-
12
#297240000000
0!
0%
b110 *
0-
02
b110 6
#297250000000
1!
1%
1-
12
#297260000000
0!
0%
b111 *
0-
02
b111 6
#297270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#297280000000
0!
0%
b0 *
0-
02
b0 6
#297290000000
1!
1%
1-
12
#297300000000
0!
0%
b1 *
0-
02
b1 6
#297310000000
1!
1%
1-
12
#297320000000
0!
0%
b10 *
0-
02
b10 6
#297330000000
1!
1%
1-
12
#297340000000
0!
0%
b11 *
0-
02
b11 6
#297350000000
1!
1%
1-
12
15
#297360000000
0!
0%
b100 *
0-
02
b100 6
#297370000000
1!
1%
1-
12
#297380000000
0!
0%
b101 *
0-
02
b101 6
#297390000000
1!
1%
1-
12
#297400000000
0!
0%
b110 *
0-
02
b110 6
#297410000000
1!
1%
1-
12
#297420000000
0!
0%
b111 *
0-
02
b111 6
#297430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#297440000000
0!
0%
b0 *
0-
02
b0 6
#297450000000
1!
1%
1-
12
#297460000000
0!
0%
b1 *
0-
02
b1 6
#297470000000
1!
1%
1-
12
#297480000000
0!
0%
b10 *
0-
02
b10 6
#297490000000
1!
1%
1-
12
#297500000000
0!
0%
b11 *
0-
02
b11 6
#297510000000
1!
1%
1-
12
15
#297520000000
0!
0%
b100 *
0-
02
b100 6
#297530000000
1!
1%
1-
12
#297540000000
0!
0%
b101 *
0-
02
b101 6
#297550000000
1!
1%
1-
12
#297560000000
0!
0%
b110 *
0-
02
b110 6
#297570000000
1!
1%
1-
12
#297580000000
0!
0%
b111 *
0-
02
b111 6
#297590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#297600000000
0!
0%
b0 *
0-
02
b0 6
#297610000000
1!
1%
1-
12
#297620000000
0!
0%
b1 *
0-
02
b1 6
#297630000000
1!
1%
1-
12
#297640000000
0!
0%
b10 *
0-
02
b10 6
#297650000000
1!
1%
1-
12
#297660000000
0!
0%
b11 *
0-
02
b11 6
#297670000000
1!
1%
1-
12
15
#297680000000
0!
0%
b100 *
0-
02
b100 6
#297690000000
1!
1%
1-
12
#297700000000
0!
0%
b101 *
0-
02
b101 6
#297710000000
1!
1%
1-
12
#297720000000
0!
0%
b110 *
0-
02
b110 6
#297730000000
1!
1%
1-
12
#297740000000
0!
0%
b111 *
0-
02
b111 6
#297750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#297760000000
0!
0%
b0 *
0-
02
b0 6
#297770000000
1!
1%
1-
12
#297780000000
0!
0%
b1 *
0-
02
b1 6
#297790000000
1!
1%
1-
12
#297800000000
0!
0%
b10 *
0-
02
b10 6
#297810000000
1!
1%
1-
12
#297820000000
0!
0%
b11 *
0-
02
b11 6
#297830000000
1!
1%
1-
12
15
#297840000000
0!
0%
b100 *
0-
02
b100 6
#297850000000
1!
1%
1-
12
#297860000000
0!
0%
b101 *
0-
02
b101 6
#297870000000
1!
1%
1-
12
#297880000000
0!
0%
b110 *
0-
02
b110 6
#297890000000
1!
1%
1-
12
#297900000000
0!
0%
b111 *
0-
02
b111 6
#297910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#297920000000
0!
0%
b0 *
0-
02
b0 6
#297930000000
1!
1%
1-
12
#297940000000
0!
0%
b1 *
0-
02
b1 6
#297950000000
1!
1%
1-
12
#297960000000
0!
0%
b10 *
0-
02
b10 6
#297970000000
1!
1%
1-
12
#297980000000
0!
0%
b11 *
0-
02
b11 6
#297990000000
1!
1%
1-
12
15
#298000000000
0!
0%
b100 *
0-
02
b100 6
#298010000000
1!
1%
1-
12
#298020000000
0!
0%
b101 *
0-
02
b101 6
#298030000000
1!
1%
1-
12
#298040000000
0!
0%
b110 *
0-
02
b110 6
#298050000000
1!
1%
1-
12
#298060000000
0!
0%
b111 *
0-
02
b111 6
#298070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#298080000000
0!
0%
b0 *
0-
02
b0 6
#298090000000
1!
1%
1-
12
#298100000000
0!
0%
b1 *
0-
02
b1 6
#298110000000
1!
1%
1-
12
#298120000000
0!
0%
b10 *
0-
02
b10 6
#298130000000
1!
1%
1-
12
#298140000000
0!
0%
b11 *
0-
02
b11 6
#298150000000
1!
1%
1-
12
15
#298160000000
0!
0%
b100 *
0-
02
b100 6
#298170000000
1!
1%
1-
12
#298180000000
0!
0%
b101 *
0-
02
b101 6
#298190000000
1!
1%
1-
12
#298200000000
0!
0%
b110 *
0-
02
b110 6
#298210000000
1!
1%
1-
12
#298220000000
0!
0%
b111 *
0-
02
b111 6
#298230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#298240000000
0!
0%
b0 *
0-
02
b0 6
#298250000000
1!
1%
1-
12
#298260000000
0!
0%
b1 *
0-
02
b1 6
#298270000000
1!
1%
1-
12
#298280000000
0!
0%
b10 *
0-
02
b10 6
#298290000000
1!
1%
1-
12
#298300000000
0!
0%
b11 *
0-
02
b11 6
#298310000000
1!
1%
1-
12
15
#298320000000
0!
0%
b100 *
0-
02
b100 6
#298330000000
1!
1%
1-
12
#298340000000
0!
0%
b101 *
0-
02
b101 6
#298350000000
1!
1%
1-
12
#298360000000
0!
0%
b110 *
0-
02
b110 6
#298370000000
1!
1%
1-
12
#298380000000
0!
0%
b111 *
0-
02
b111 6
#298390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#298400000000
0!
0%
b0 *
0-
02
b0 6
#298410000000
1!
1%
1-
12
#298420000000
0!
0%
b1 *
0-
02
b1 6
#298430000000
1!
1%
1-
12
#298440000000
0!
0%
b10 *
0-
02
b10 6
#298450000000
1!
1%
1-
12
#298460000000
0!
0%
b11 *
0-
02
b11 6
#298470000000
1!
1%
1-
12
15
#298480000000
0!
0%
b100 *
0-
02
b100 6
#298490000000
1!
1%
1-
12
#298500000000
0!
0%
b101 *
0-
02
b101 6
#298510000000
1!
1%
1-
12
#298520000000
0!
0%
b110 *
0-
02
b110 6
#298530000000
1!
1%
1-
12
#298540000000
0!
0%
b111 *
0-
02
b111 6
#298550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#298560000000
0!
0%
b0 *
0-
02
b0 6
#298570000000
1!
1%
1-
12
#298580000000
0!
0%
b1 *
0-
02
b1 6
#298590000000
1!
1%
1-
12
#298600000000
0!
0%
b10 *
0-
02
b10 6
#298610000000
1!
1%
1-
12
#298620000000
0!
0%
b11 *
0-
02
b11 6
#298630000000
1!
1%
1-
12
15
#298640000000
0!
0%
b100 *
0-
02
b100 6
#298650000000
1!
1%
1-
12
#298660000000
0!
0%
b101 *
0-
02
b101 6
#298670000000
1!
1%
1-
12
#298680000000
0!
0%
b110 *
0-
02
b110 6
#298690000000
1!
1%
1-
12
#298700000000
0!
0%
b111 *
0-
02
b111 6
#298710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#298720000000
0!
0%
b0 *
0-
02
b0 6
#298730000000
1!
1%
1-
12
#298740000000
0!
0%
b1 *
0-
02
b1 6
#298750000000
1!
1%
1-
12
#298760000000
0!
0%
b10 *
0-
02
b10 6
#298770000000
1!
1%
1-
12
#298780000000
0!
0%
b11 *
0-
02
b11 6
#298790000000
1!
1%
1-
12
15
#298800000000
0!
0%
b100 *
0-
02
b100 6
#298810000000
1!
1%
1-
12
#298820000000
0!
0%
b101 *
0-
02
b101 6
#298830000000
1!
1%
1-
12
#298840000000
0!
0%
b110 *
0-
02
b110 6
#298850000000
1!
1%
1-
12
#298860000000
0!
0%
b111 *
0-
02
b111 6
#298870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#298880000000
0!
0%
b0 *
0-
02
b0 6
#298890000000
1!
1%
1-
12
#298900000000
0!
0%
b1 *
0-
02
b1 6
#298910000000
1!
1%
1-
12
#298920000000
0!
0%
b10 *
0-
02
b10 6
#298930000000
1!
1%
1-
12
#298940000000
0!
0%
b11 *
0-
02
b11 6
#298950000000
1!
1%
1-
12
15
#298960000000
0!
0%
b100 *
0-
02
b100 6
#298970000000
1!
1%
1-
12
#298980000000
0!
0%
b101 *
0-
02
b101 6
#298990000000
1!
1%
1-
12
#299000000000
0!
0%
b110 *
0-
02
b110 6
#299010000000
1!
1%
1-
12
#299020000000
0!
0%
b111 *
0-
02
b111 6
#299030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#299040000000
0!
0%
b0 *
0-
02
b0 6
#299050000000
1!
1%
1-
12
#299060000000
0!
0%
b1 *
0-
02
b1 6
#299070000000
1!
1%
1-
12
#299080000000
0!
0%
b10 *
0-
02
b10 6
#299090000000
1!
1%
1-
12
#299100000000
0!
0%
b11 *
0-
02
b11 6
#299110000000
1!
1%
1-
12
15
#299120000000
0!
0%
b100 *
0-
02
b100 6
#299130000000
1!
1%
1-
12
#299140000000
0!
0%
b101 *
0-
02
b101 6
#299150000000
1!
1%
1-
12
#299160000000
0!
0%
b110 *
0-
02
b110 6
#299170000000
1!
1%
1-
12
#299180000000
0!
0%
b111 *
0-
02
b111 6
#299190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#299200000000
0!
0%
b0 *
0-
02
b0 6
#299210000000
1!
1%
1-
12
#299220000000
0!
0%
b1 *
0-
02
b1 6
#299230000000
1!
1%
1-
12
#299240000000
0!
0%
b10 *
0-
02
b10 6
#299250000000
1!
1%
1-
12
#299260000000
0!
0%
b11 *
0-
02
b11 6
#299270000000
1!
1%
1-
12
15
#299280000000
0!
0%
b100 *
0-
02
b100 6
#299290000000
1!
1%
1-
12
#299300000000
0!
0%
b101 *
0-
02
b101 6
#299310000000
1!
1%
1-
12
#299320000000
0!
0%
b110 *
0-
02
b110 6
#299330000000
1!
1%
1-
12
#299340000000
0!
0%
b111 *
0-
02
b111 6
#299350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#299360000000
0!
0%
b0 *
0-
02
b0 6
#299370000000
1!
1%
1-
12
#299380000000
0!
0%
b1 *
0-
02
b1 6
#299390000000
1!
1%
1-
12
#299400000000
0!
0%
b10 *
0-
02
b10 6
#299410000000
1!
1%
1-
12
#299420000000
0!
0%
b11 *
0-
02
b11 6
#299430000000
1!
1%
1-
12
15
#299440000000
0!
0%
b100 *
0-
02
b100 6
#299450000000
1!
1%
1-
12
#299460000000
0!
0%
b101 *
0-
02
b101 6
#299470000000
1!
1%
1-
12
#299480000000
0!
0%
b110 *
0-
02
b110 6
#299490000000
1!
1%
1-
12
#299500000000
0!
0%
b111 *
0-
02
b111 6
#299510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#299520000000
0!
0%
b0 *
0-
02
b0 6
#299530000000
1!
1%
1-
12
#299540000000
0!
0%
b1 *
0-
02
b1 6
#299550000000
1!
1%
1-
12
#299560000000
0!
0%
b10 *
0-
02
b10 6
#299570000000
1!
1%
1-
12
#299580000000
0!
0%
b11 *
0-
02
b11 6
#299590000000
1!
1%
1-
12
15
#299600000000
0!
0%
b100 *
0-
02
b100 6
#299610000000
1!
1%
1-
12
#299620000000
0!
0%
b101 *
0-
02
b101 6
#299630000000
1!
1%
1-
12
#299640000000
0!
0%
b110 *
0-
02
b110 6
#299650000000
1!
1%
1-
12
#299660000000
0!
0%
b111 *
0-
02
b111 6
#299670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#299680000000
0!
0%
b0 *
0-
02
b0 6
#299690000000
1!
1%
1-
12
#299700000000
0!
0%
b1 *
0-
02
b1 6
#299710000000
1!
1%
1-
12
#299720000000
0!
0%
b10 *
0-
02
b10 6
#299730000000
1!
1%
1-
12
#299740000000
0!
0%
b11 *
0-
02
b11 6
#299750000000
1!
1%
1-
12
15
#299760000000
0!
0%
b100 *
0-
02
b100 6
#299770000000
1!
1%
1-
12
#299780000000
0!
0%
b101 *
0-
02
b101 6
#299790000000
1!
1%
1-
12
#299800000000
0!
0%
b110 *
0-
02
b110 6
#299810000000
1!
1%
1-
12
#299820000000
0!
0%
b111 *
0-
02
b111 6
#299830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#299840000000
0!
0%
b0 *
0-
02
b0 6
#299850000000
1!
1%
1-
12
#299860000000
0!
0%
b1 *
0-
02
b1 6
#299870000000
1!
1%
1-
12
#299880000000
0!
0%
b10 *
0-
02
b10 6
#299890000000
1!
1%
1-
12
#299900000000
0!
0%
b11 *
0-
02
b11 6
#299910000000
1!
1%
1-
12
15
#299920000000
0!
0%
b100 *
0-
02
b100 6
#299930000000
1!
1%
1-
12
#299940000000
0!
0%
b101 *
0-
02
b101 6
#299950000000
1!
1%
1-
12
#299960000000
0!
0%
b110 *
0-
02
b110 6
#299970000000
1!
1%
1-
12
#299980000000
0!
0%
b111 *
0-
02
b111 6
#299990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#300000000000
0!
0%
b0 *
0-
02
b0 6
#300010000000
1!
1%
1-
12
#300020000000
0!
0%
b1 *
0-
02
b1 6
#300030000000
1!
1%
1-
12
#300040000000
0!
0%
b10 *
0-
02
b10 6
#300050000000
1!
1%
1-
12
#300060000000
0!
0%
b11 *
0-
02
b11 6
#300070000000
1!
1%
1-
12
15
#300080000000
0!
0%
b100 *
0-
02
b100 6
#300090000000
1!
1%
1-
12
#300100000000
0!
0%
b101 *
0-
02
b101 6
#300110000000
1!
1%
1-
12
#300120000000
0!
0%
b110 *
0-
02
b110 6
#300130000000
1!
1%
1-
12
#300140000000
0!
0%
b111 *
0-
02
b111 6
#300150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#300160000000
0!
0%
b0 *
0-
02
b0 6
#300170000000
1!
1%
1-
12
#300180000000
0!
0%
b1 *
0-
02
b1 6
#300190000000
1!
1%
1-
12
#300200000000
0!
0%
b10 *
0-
02
b10 6
#300210000000
1!
1%
1-
12
#300220000000
0!
0%
b11 *
0-
02
b11 6
#300230000000
1!
1%
1-
12
15
#300240000000
0!
0%
b100 *
0-
02
b100 6
#300250000000
1!
1%
1-
12
#300260000000
0!
0%
b101 *
0-
02
b101 6
#300270000000
1!
1%
1-
12
#300280000000
0!
0%
b110 *
0-
02
b110 6
#300290000000
1!
1%
1-
12
#300300000000
0!
0%
b111 *
0-
02
b111 6
#300310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#300320000000
0!
0%
b0 *
0-
02
b0 6
#300330000000
1!
1%
1-
12
#300340000000
0!
0%
b1 *
0-
02
b1 6
#300350000000
1!
1%
1-
12
#300360000000
0!
0%
b10 *
0-
02
b10 6
#300370000000
1!
1%
1-
12
#300380000000
0!
0%
b11 *
0-
02
b11 6
#300390000000
1!
1%
1-
12
15
#300400000000
0!
0%
b100 *
0-
02
b100 6
#300410000000
1!
1%
1-
12
#300420000000
0!
0%
b101 *
0-
02
b101 6
#300430000000
1!
1%
1-
12
#300440000000
0!
0%
b110 *
0-
02
b110 6
#300450000000
1!
1%
1-
12
#300460000000
0!
0%
b111 *
0-
02
b111 6
#300470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#300480000000
0!
0%
b0 *
0-
02
b0 6
#300490000000
1!
1%
1-
12
#300500000000
0!
0%
b1 *
0-
02
b1 6
#300510000000
1!
1%
1-
12
#300520000000
0!
0%
b10 *
0-
02
b10 6
#300530000000
1!
1%
1-
12
#300540000000
0!
0%
b11 *
0-
02
b11 6
#300550000000
1!
1%
1-
12
15
#300560000000
0!
0%
b100 *
0-
02
b100 6
#300570000000
1!
1%
1-
12
#300580000000
0!
0%
b101 *
0-
02
b101 6
#300590000000
1!
1%
1-
12
#300600000000
0!
0%
b110 *
0-
02
b110 6
#300610000000
1!
1%
1-
12
#300620000000
0!
0%
b111 *
0-
02
b111 6
#300630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#300640000000
0!
0%
b0 *
0-
02
b0 6
#300650000000
1!
1%
1-
12
#300660000000
0!
0%
b1 *
0-
02
b1 6
#300670000000
1!
1%
1-
12
#300680000000
0!
0%
b10 *
0-
02
b10 6
#300690000000
1!
1%
1-
12
#300700000000
0!
0%
b11 *
0-
02
b11 6
#300710000000
1!
1%
1-
12
15
#300720000000
0!
0%
b100 *
0-
02
b100 6
#300730000000
1!
1%
1-
12
#300740000000
0!
0%
b101 *
0-
02
b101 6
#300750000000
1!
1%
1-
12
#300760000000
0!
0%
b110 *
0-
02
b110 6
#300770000000
1!
1%
1-
12
#300780000000
0!
0%
b111 *
0-
02
b111 6
#300790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#300800000000
0!
0%
b0 *
0-
02
b0 6
#300810000000
1!
1%
1-
12
#300820000000
0!
0%
b1 *
0-
02
b1 6
#300830000000
1!
1%
1-
12
#300840000000
0!
0%
b10 *
0-
02
b10 6
#300850000000
1!
1%
1-
12
#300860000000
0!
0%
b11 *
0-
02
b11 6
#300870000000
1!
1%
1-
12
15
#300880000000
0!
0%
b100 *
0-
02
b100 6
#300890000000
1!
1%
1-
12
#300900000000
0!
0%
b101 *
0-
02
b101 6
#300910000000
1!
1%
1-
12
#300920000000
0!
0%
b110 *
0-
02
b110 6
#300930000000
1!
1%
1-
12
#300940000000
0!
0%
b111 *
0-
02
b111 6
#300950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#300960000000
0!
0%
b0 *
0-
02
b0 6
#300970000000
1!
1%
1-
12
#300980000000
0!
0%
b1 *
0-
02
b1 6
#300990000000
1!
1%
1-
12
#301000000000
0!
0%
b10 *
0-
02
b10 6
#301010000000
1!
1%
1-
12
#301020000000
0!
0%
b11 *
0-
02
b11 6
#301030000000
1!
1%
1-
12
15
#301040000000
0!
0%
b100 *
0-
02
b100 6
#301050000000
1!
1%
1-
12
#301060000000
0!
0%
b101 *
0-
02
b101 6
#301070000000
1!
1%
1-
12
#301080000000
0!
0%
b110 *
0-
02
b110 6
#301090000000
1!
1%
1-
12
#301100000000
0!
0%
b111 *
0-
02
b111 6
#301110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#301120000000
0!
0%
b0 *
0-
02
b0 6
#301130000000
1!
1%
1-
12
#301140000000
0!
0%
b1 *
0-
02
b1 6
#301150000000
1!
1%
1-
12
#301160000000
0!
0%
b10 *
0-
02
b10 6
#301170000000
1!
1%
1-
12
#301180000000
0!
0%
b11 *
0-
02
b11 6
#301190000000
1!
1%
1-
12
15
#301200000000
0!
0%
b100 *
0-
02
b100 6
#301210000000
1!
1%
1-
12
#301220000000
0!
0%
b101 *
0-
02
b101 6
#301230000000
1!
1%
1-
12
#301240000000
0!
0%
b110 *
0-
02
b110 6
#301250000000
1!
1%
1-
12
#301260000000
0!
0%
b111 *
0-
02
b111 6
#301270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#301280000000
0!
0%
b0 *
0-
02
b0 6
#301290000000
1!
1%
1-
12
#301300000000
0!
0%
b1 *
0-
02
b1 6
#301310000000
1!
1%
1-
12
#301320000000
0!
0%
b10 *
0-
02
b10 6
#301330000000
1!
1%
1-
12
#301340000000
0!
0%
b11 *
0-
02
b11 6
#301350000000
1!
1%
1-
12
15
#301360000000
0!
0%
b100 *
0-
02
b100 6
#301370000000
1!
1%
1-
12
#301380000000
0!
0%
b101 *
0-
02
b101 6
#301390000000
1!
1%
1-
12
#301400000000
0!
0%
b110 *
0-
02
b110 6
#301410000000
1!
1%
1-
12
#301420000000
0!
0%
b111 *
0-
02
b111 6
#301430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#301440000000
0!
0%
b0 *
0-
02
b0 6
#301450000000
1!
1%
1-
12
#301460000000
0!
0%
b1 *
0-
02
b1 6
#301470000000
1!
1%
1-
12
#301480000000
0!
0%
b10 *
0-
02
b10 6
#301490000000
1!
1%
1-
12
#301500000000
0!
0%
b11 *
0-
02
b11 6
#301510000000
1!
1%
1-
12
15
#301520000000
0!
0%
b100 *
0-
02
b100 6
#301530000000
1!
1%
1-
12
#301540000000
0!
0%
b101 *
0-
02
b101 6
#301550000000
1!
1%
1-
12
#301560000000
0!
0%
b110 *
0-
02
b110 6
#301570000000
1!
1%
1-
12
#301580000000
0!
0%
b111 *
0-
02
b111 6
#301590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#301600000000
0!
0%
b0 *
0-
02
b0 6
#301610000000
1!
1%
1-
12
#301620000000
0!
0%
b1 *
0-
02
b1 6
#301630000000
1!
1%
1-
12
#301640000000
0!
0%
b10 *
0-
02
b10 6
#301650000000
1!
1%
1-
12
#301660000000
0!
0%
b11 *
0-
02
b11 6
#301670000000
1!
1%
1-
12
15
#301680000000
0!
0%
b100 *
0-
02
b100 6
#301690000000
1!
1%
1-
12
#301700000000
0!
0%
b101 *
0-
02
b101 6
#301710000000
1!
1%
1-
12
#301720000000
0!
0%
b110 *
0-
02
b110 6
#301730000000
1!
1%
1-
12
#301740000000
0!
0%
b111 *
0-
02
b111 6
#301750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#301760000000
0!
0%
b0 *
0-
02
b0 6
#301770000000
1!
1%
1-
12
#301780000000
0!
0%
b1 *
0-
02
b1 6
#301790000000
1!
1%
1-
12
#301800000000
0!
0%
b10 *
0-
02
b10 6
#301810000000
1!
1%
1-
12
#301820000000
0!
0%
b11 *
0-
02
b11 6
#301830000000
1!
1%
1-
12
15
#301840000000
0!
0%
b100 *
0-
02
b100 6
#301850000000
1!
1%
1-
12
#301860000000
0!
0%
b101 *
0-
02
b101 6
#301870000000
1!
1%
1-
12
#301880000000
0!
0%
b110 *
0-
02
b110 6
#301890000000
1!
1%
1-
12
#301900000000
0!
0%
b111 *
0-
02
b111 6
#301910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#301920000000
0!
0%
b0 *
0-
02
b0 6
#301930000000
1!
1%
1-
12
#301940000000
0!
0%
b1 *
0-
02
b1 6
#301950000000
1!
1%
1-
12
#301960000000
0!
0%
b10 *
0-
02
b10 6
#301970000000
1!
1%
1-
12
#301980000000
0!
0%
b11 *
0-
02
b11 6
#301990000000
1!
1%
1-
12
15
#302000000000
0!
0%
b100 *
0-
02
b100 6
#302010000000
1!
1%
1-
12
#302020000000
0!
0%
b101 *
0-
02
b101 6
#302030000000
1!
1%
1-
12
#302040000000
0!
0%
b110 *
0-
02
b110 6
#302050000000
1!
1%
1-
12
#302060000000
0!
0%
b111 *
0-
02
b111 6
#302070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#302080000000
0!
0%
b0 *
0-
02
b0 6
#302090000000
1!
1%
1-
12
#302100000000
0!
0%
b1 *
0-
02
b1 6
#302110000000
1!
1%
1-
12
#302120000000
0!
0%
b10 *
0-
02
b10 6
#302130000000
1!
1%
1-
12
#302140000000
0!
0%
b11 *
0-
02
b11 6
#302150000000
1!
1%
1-
12
15
#302160000000
0!
0%
b100 *
0-
02
b100 6
#302170000000
1!
1%
1-
12
#302180000000
0!
0%
b101 *
0-
02
b101 6
#302190000000
1!
1%
1-
12
#302200000000
0!
0%
b110 *
0-
02
b110 6
#302210000000
1!
1%
1-
12
#302220000000
0!
0%
b111 *
0-
02
b111 6
#302230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#302240000000
0!
0%
b0 *
0-
02
b0 6
#302250000000
1!
1%
1-
12
#302260000000
0!
0%
b1 *
0-
02
b1 6
#302270000000
1!
1%
1-
12
#302280000000
0!
0%
b10 *
0-
02
b10 6
#302290000000
1!
1%
1-
12
#302300000000
0!
0%
b11 *
0-
02
b11 6
#302310000000
1!
1%
1-
12
15
#302320000000
0!
0%
b100 *
0-
02
b100 6
#302330000000
1!
1%
1-
12
#302340000000
0!
0%
b101 *
0-
02
b101 6
#302350000000
1!
1%
1-
12
#302360000000
0!
0%
b110 *
0-
02
b110 6
#302370000000
1!
1%
1-
12
#302380000000
0!
0%
b111 *
0-
02
b111 6
#302390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#302400000000
0!
0%
b0 *
0-
02
b0 6
#302410000000
1!
1%
1-
12
#302420000000
0!
0%
b1 *
0-
02
b1 6
#302430000000
1!
1%
1-
12
#302440000000
0!
0%
b10 *
0-
02
b10 6
#302450000000
1!
1%
1-
12
#302460000000
0!
0%
b11 *
0-
02
b11 6
#302470000000
1!
1%
1-
12
15
#302480000000
0!
0%
b100 *
0-
02
b100 6
#302490000000
1!
1%
1-
12
#302500000000
0!
0%
b101 *
0-
02
b101 6
#302510000000
1!
1%
1-
12
#302520000000
0!
0%
b110 *
0-
02
b110 6
#302530000000
1!
1%
1-
12
#302540000000
0!
0%
b111 *
0-
02
b111 6
#302550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#302560000000
0!
0%
b0 *
0-
02
b0 6
#302570000000
1!
1%
1-
12
#302580000000
0!
0%
b1 *
0-
02
b1 6
#302590000000
1!
1%
1-
12
#302600000000
0!
0%
b10 *
0-
02
b10 6
#302610000000
1!
1%
1-
12
#302620000000
0!
0%
b11 *
0-
02
b11 6
#302630000000
1!
1%
1-
12
15
#302640000000
0!
0%
b100 *
0-
02
b100 6
#302650000000
1!
1%
1-
12
#302660000000
0!
0%
b101 *
0-
02
b101 6
#302670000000
1!
1%
1-
12
#302680000000
0!
0%
b110 *
0-
02
b110 6
#302690000000
1!
1%
1-
12
#302700000000
0!
0%
b111 *
0-
02
b111 6
#302710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#302720000000
0!
0%
b0 *
0-
02
b0 6
#302730000000
1!
1%
1-
12
#302740000000
0!
0%
b1 *
0-
02
b1 6
#302750000000
1!
1%
1-
12
#302760000000
0!
0%
b10 *
0-
02
b10 6
#302770000000
1!
1%
1-
12
#302780000000
0!
0%
b11 *
0-
02
b11 6
#302790000000
1!
1%
1-
12
15
#302800000000
0!
0%
b100 *
0-
02
b100 6
#302810000000
1!
1%
1-
12
#302820000000
0!
0%
b101 *
0-
02
b101 6
#302830000000
1!
1%
1-
12
#302840000000
0!
0%
b110 *
0-
02
b110 6
#302850000000
1!
1%
1-
12
#302860000000
0!
0%
b111 *
0-
02
b111 6
#302870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#302880000000
0!
0%
b0 *
0-
02
b0 6
#302890000000
1!
1%
1-
12
#302900000000
0!
0%
b1 *
0-
02
b1 6
#302910000000
1!
1%
1-
12
#302920000000
0!
0%
b10 *
0-
02
b10 6
#302930000000
1!
1%
1-
12
#302940000000
0!
0%
b11 *
0-
02
b11 6
#302950000000
1!
1%
1-
12
15
#302960000000
0!
0%
b100 *
0-
02
b100 6
#302970000000
1!
1%
1-
12
#302980000000
0!
0%
b101 *
0-
02
b101 6
#302990000000
1!
1%
1-
12
#303000000000
0!
0%
b110 *
0-
02
b110 6
#303010000000
1!
1%
1-
12
#303020000000
0!
0%
b111 *
0-
02
b111 6
#303030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#303040000000
0!
0%
b0 *
0-
02
b0 6
#303050000000
1!
1%
1-
12
#303060000000
0!
0%
b1 *
0-
02
b1 6
#303070000000
1!
1%
1-
12
#303080000000
0!
0%
b10 *
0-
02
b10 6
#303090000000
1!
1%
1-
12
#303100000000
0!
0%
b11 *
0-
02
b11 6
#303110000000
1!
1%
1-
12
15
#303120000000
0!
0%
b100 *
0-
02
b100 6
#303130000000
1!
1%
1-
12
#303140000000
0!
0%
b101 *
0-
02
b101 6
#303150000000
1!
1%
1-
12
#303160000000
0!
0%
b110 *
0-
02
b110 6
#303170000000
1!
1%
1-
12
#303180000000
0!
0%
b111 *
0-
02
b111 6
#303190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#303200000000
0!
0%
b0 *
0-
02
b0 6
#303210000000
1!
1%
1-
12
#303220000000
0!
0%
b1 *
0-
02
b1 6
#303230000000
1!
1%
1-
12
#303240000000
0!
0%
b10 *
0-
02
b10 6
#303250000000
1!
1%
1-
12
#303260000000
0!
0%
b11 *
0-
02
b11 6
#303270000000
1!
1%
1-
12
15
#303280000000
0!
0%
b100 *
0-
02
b100 6
#303290000000
1!
1%
1-
12
#303300000000
0!
0%
b101 *
0-
02
b101 6
#303310000000
1!
1%
1-
12
#303320000000
0!
0%
b110 *
0-
02
b110 6
#303330000000
1!
1%
1-
12
#303340000000
0!
0%
b111 *
0-
02
b111 6
#303350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#303360000000
0!
0%
b0 *
0-
02
b0 6
#303370000000
1!
1%
1-
12
#303380000000
0!
0%
b1 *
0-
02
b1 6
#303390000000
1!
1%
1-
12
#303400000000
0!
0%
b10 *
0-
02
b10 6
#303410000000
1!
1%
1-
12
#303420000000
0!
0%
b11 *
0-
02
b11 6
#303430000000
1!
1%
1-
12
15
#303440000000
0!
0%
b100 *
0-
02
b100 6
#303450000000
1!
1%
1-
12
#303460000000
0!
0%
b101 *
0-
02
b101 6
#303470000000
1!
1%
1-
12
#303480000000
0!
0%
b110 *
0-
02
b110 6
#303490000000
1!
1%
1-
12
#303500000000
0!
0%
b111 *
0-
02
b111 6
#303510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#303520000000
0!
0%
b0 *
0-
02
b0 6
#303530000000
1!
1%
1-
12
#303540000000
0!
0%
b1 *
0-
02
b1 6
#303550000000
1!
1%
1-
12
#303560000000
0!
0%
b10 *
0-
02
b10 6
#303570000000
1!
1%
1-
12
#303580000000
0!
0%
b11 *
0-
02
b11 6
#303590000000
1!
1%
1-
12
15
#303600000000
0!
0%
b100 *
0-
02
b100 6
#303610000000
1!
1%
1-
12
#303620000000
0!
0%
b101 *
0-
02
b101 6
#303630000000
1!
1%
1-
12
#303640000000
0!
0%
b110 *
0-
02
b110 6
#303650000000
1!
1%
1-
12
#303660000000
0!
0%
b111 *
0-
02
b111 6
#303670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#303680000000
0!
0%
b0 *
0-
02
b0 6
#303690000000
1!
1%
1-
12
#303700000000
0!
0%
b1 *
0-
02
b1 6
#303710000000
1!
1%
1-
12
#303720000000
0!
0%
b10 *
0-
02
b10 6
#303730000000
1!
1%
1-
12
#303740000000
0!
0%
b11 *
0-
02
b11 6
#303750000000
1!
1%
1-
12
15
#303760000000
0!
0%
b100 *
0-
02
b100 6
#303770000000
1!
1%
1-
12
#303780000000
0!
0%
b101 *
0-
02
b101 6
#303790000000
1!
1%
1-
12
#303800000000
0!
0%
b110 *
0-
02
b110 6
#303810000000
1!
1%
1-
12
#303820000000
0!
0%
b111 *
0-
02
b111 6
#303830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#303840000000
0!
0%
b0 *
0-
02
b0 6
#303850000000
1!
1%
1-
12
#303860000000
0!
0%
b1 *
0-
02
b1 6
#303870000000
1!
1%
1-
12
#303880000000
0!
0%
b10 *
0-
02
b10 6
#303890000000
1!
1%
1-
12
#303900000000
0!
0%
b11 *
0-
02
b11 6
#303910000000
1!
1%
1-
12
15
#303920000000
0!
0%
b100 *
0-
02
b100 6
#303930000000
1!
1%
1-
12
#303940000000
0!
0%
b101 *
0-
02
b101 6
#303950000000
1!
1%
1-
12
#303960000000
0!
0%
b110 *
0-
02
b110 6
#303970000000
1!
1%
1-
12
#303980000000
0!
0%
b111 *
0-
02
b111 6
#303990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#304000000000
0!
0%
b0 *
0-
02
b0 6
#304010000000
1!
1%
1-
12
#304020000000
0!
0%
b1 *
0-
02
b1 6
#304030000000
1!
1%
1-
12
#304040000000
0!
0%
b10 *
0-
02
b10 6
#304050000000
1!
1%
1-
12
#304060000000
0!
0%
b11 *
0-
02
b11 6
#304070000000
1!
1%
1-
12
15
#304080000000
0!
0%
b100 *
0-
02
b100 6
#304090000000
1!
1%
1-
12
#304100000000
0!
0%
b101 *
0-
02
b101 6
#304110000000
1!
1%
1-
12
#304120000000
0!
0%
b110 *
0-
02
b110 6
#304130000000
1!
1%
1-
12
#304140000000
0!
0%
b111 *
0-
02
b111 6
#304150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#304160000000
0!
0%
b0 *
0-
02
b0 6
#304170000000
1!
1%
1-
12
#304180000000
0!
0%
b1 *
0-
02
b1 6
#304190000000
1!
1%
1-
12
#304200000000
0!
0%
b10 *
0-
02
b10 6
#304210000000
1!
1%
1-
12
#304220000000
0!
0%
b11 *
0-
02
b11 6
#304230000000
1!
1%
1-
12
15
#304240000000
0!
0%
b100 *
0-
02
b100 6
#304250000000
1!
1%
1-
12
#304260000000
0!
0%
b101 *
0-
02
b101 6
#304270000000
1!
1%
1-
12
#304280000000
0!
0%
b110 *
0-
02
b110 6
#304290000000
1!
1%
1-
12
#304300000000
0!
0%
b111 *
0-
02
b111 6
#304310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#304320000000
0!
0%
b0 *
0-
02
b0 6
#304330000000
1!
1%
1-
12
#304340000000
0!
0%
b1 *
0-
02
b1 6
#304350000000
1!
1%
1-
12
#304360000000
0!
0%
b10 *
0-
02
b10 6
#304370000000
1!
1%
1-
12
#304380000000
0!
0%
b11 *
0-
02
b11 6
#304390000000
1!
1%
1-
12
15
#304400000000
0!
0%
b100 *
0-
02
b100 6
#304410000000
1!
1%
1-
12
#304420000000
0!
0%
b101 *
0-
02
b101 6
#304430000000
1!
1%
1-
12
#304440000000
0!
0%
b110 *
0-
02
b110 6
#304450000000
1!
1%
1-
12
#304460000000
0!
0%
b111 *
0-
02
b111 6
#304470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#304480000000
0!
0%
b0 *
0-
02
b0 6
#304490000000
1!
1%
1-
12
#304500000000
0!
0%
b1 *
0-
02
b1 6
#304510000000
1!
1%
1-
12
#304520000000
0!
0%
b10 *
0-
02
b10 6
#304530000000
1!
1%
1-
12
#304540000000
0!
0%
b11 *
0-
02
b11 6
#304550000000
1!
1%
1-
12
15
#304560000000
0!
0%
b100 *
0-
02
b100 6
#304570000000
1!
1%
1-
12
#304580000000
0!
0%
b101 *
0-
02
b101 6
#304590000000
1!
1%
1-
12
#304600000000
0!
0%
b110 *
0-
02
b110 6
#304610000000
1!
1%
1-
12
#304620000000
0!
0%
b111 *
0-
02
b111 6
#304630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#304640000000
0!
0%
b0 *
0-
02
b0 6
#304650000000
1!
1%
1-
12
#304660000000
0!
0%
b1 *
0-
02
b1 6
#304670000000
1!
1%
1-
12
#304680000000
0!
0%
b10 *
0-
02
b10 6
#304690000000
1!
1%
1-
12
#304700000000
0!
0%
b11 *
0-
02
b11 6
#304710000000
1!
1%
1-
12
15
#304720000000
0!
0%
b100 *
0-
02
b100 6
#304730000000
1!
1%
1-
12
#304740000000
0!
0%
b101 *
0-
02
b101 6
#304750000000
1!
1%
1-
12
#304760000000
0!
0%
b110 *
0-
02
b110 6
#304770000000
1!
1%
1-
12
#304780000000
0!
0%
b111 *
0-
02
b111 6
#304790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#304800000000
0!
0%
b0 *
0-
02
b0 6
#304810000000
1!
1%
1-
12
#304820000000
0!
0%
b1 *
0-
02
b1 6
#304830000000
1!
1%
1-
12
#304840000000
0!
0%
b10 *
0-
02
b10 6
#304850000000
1!
1%
1-
12
#304860000000
0!
0%
b11 *
0-
02
b11 6
#304870000000
1!
1%
1-
12
15
#304880000000
0!
0%
b100 *
0-
02
b100 6
#304890000000
1!
1%
1-
12
#304900000000
0!
0%
b101 *
0-
02
b101 6
#304910000000
1!
1%
1-
12
#304920000000
0!
0%
b110 *
0-
02
b110 6
#304930000000
1!
1%
1-
12
#304940000000
0!
0%
b111 *
0-
02
b111 6
#304950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#304960000000
0!
0%
b0 *
0-
02
b0 6
#304970000000
1!
1%
1-
12
#304980000000
0!
0%
b1 *
0-
02
b1 6
#304990000000
1!
1%
1-
12
#305000000000
0!
0%
b10 *
0-
02
b10 6
#305010000000
1!
1%
1-
12
#305020000000
0!
0%
b11 *
0-
02
b11 6
#305030000000
1!
1%
1-
12
15
#305040000000
0!
0%
b100 *
0-
02
b100 6
#305050000000
1!
1%
1-
12
#305060000000
0!
0%
b101 *
0-
02
b101 6
#305070000000
1!
1%
1-
12
#305080000000
0!
0%
b110 *
0-
02
b110 6
#305090000000
1!
1%
1-
12
#305100000000
0!
0%
b111 *
0-
02
b111 6
#305110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#305120000000
0!
0%
b0 *
0-
02
b0 6
#305130000000
1!
1%
1-
12
#305140000000
0!
0%
b1 *
0-
02
b1 6
#305150000000
1!
1%
1-
12
#305160000000
0!
0%
b10 *
0-
02
b10 6
#305170000000
1!
1%
1-
12
#305180000000
0!
0%
b11 *
0-
02
b11 6
#305190000000
1!
1%
1-
12
15
#305200000000
0!
0%
b100 *
0-
02
b100 6
#305210000000
1!
1%
1-
12
#305220000000
0!
0%
b101 *
0-
02
b101 6
#305230000000
1!
1%
1-
12
#305240000000
0!
0%
b110 *
0-
02
b110 6
#305250000000
1!
1%
1-
12
#305260000000
0!
0%
b111 *
0-
02
b111 6
#305270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#305280000000
0!
0%
b0 *
0-
02
b0 6
#305290000000
1!
1%
1-
12
#305300000000
0!
0%
b1 *
0-
02
b1 6
#305310000000
1!
1%
1-
12
#305320000000
0!
0%
b10 *
0-
02
b10 6
#305330000000
1!
1%
1-
12
#305340000000
0!
0%
b11 *
0-
02
b11 6
#305350000000
1!
1%
1-
12
15
#305360000000
0!
0%
b100 *
0-
02
b100 6
#305370000000
1!
1%
1-
12
#305380000000
0!
0%
b101 *
0-
02
b101 6
#305390000000
1!
1%
1-
12
#305400000000
0!
0%
b110 *
0-
02
b110 6
#305410000000
1!
1%
1-
12
#305420000000
0!
0%
b111 *
0-
02
b111 6
#305430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#305440000000
0!
0%
b0 *
0-
02
b0 6
#305450000000
1!
1%
1-
12
#305460000000
0!
0%
b1 *
0-
02
b1 6
#305470000000
1!
1%
1-
12
#305480000000
0!
0%
b10 *
0-
02
b10 6
#305490000000
1!
1%
1-
12
#305500000000
0!
0%
b11 *
0-
02
b11 6
#305510000000
1!
1%
1-
12
15
#305520000000
0!
0%
b100 *
0-
02
b100 6
#305530000000
1!
1%
1-
12
#305540000000
0!
0%
b101 *
0-
02
b101 6
#305550000000
1!
1%
1-
12
#305560000000
0!
0%
b110 *
0-
02
b110 6
#305570000000
1!
1%
1-
12
#305580000000
0!
0%
b111 *
0-
02
b111 6
#305590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#305600000000
0!
0%
b0 *
0-
02
b0 6
#305610000000
1!
1%
1-
12
#305620000000
0!
0%
b1 *
0-
02
b1 6
#305630000000
1!
1%
1-
12
#305640000000
0!
0%
b10 *
0-
02
b10 6
#305650000000
1!
1%
1-
12
#305660000000
0!
0%
b11 *
0-
02
b11 6
#305670000000
1!
1%
1-
12
15
#305680000000
0!
0%
b100 *
0-
02
b100 6
#305690000000
1!
1%
1-
12
#305700000000
0!
0%
b101 *
0-
02
b101 6
#305710000000
1!
1%
1-
12
#305720000000
0!
0%
b110 *
0-
02
b110 6
#305730000000
1!
1%
1-
12
#305740000000
0!
0%
b111 *
0-
02
b111 6
#305750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#305760000000
0!
0%
b0 *
0-
02
b0 6
#305770000000
1!
1%
1-
12
#305780000000
0!
0%
b1 *
0-
02
b1 6
#305790000000
1!
1%
1-
12
#305800000000
0!
0%
b10 *
0-
02
b10 6
#305810000000
1!
1%
1-
12
#305820000000
0!
0%
b11 *
0-
02
b11 6
#305830000000
1!
1%
1-
12
15
#305840000000
0!
0%
b100 *
0-
02
b100 6
#305850000000
1!
1%
1-
12
#305860000000
0!
0%
b101 *
0-
02
b101 6
#305870000000
1!
1%
1-
12
#305880000000
0!
0%
b110 *
0-
02
b110 6
#305890000000
1!
1%
1-
12
#305900000000
0!
0%
b111 *
0-
02
b111 6
#305910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#305920000000
0!
0%
b0 *
0-
02
b0 6
#305930000000
1!
1%
1-
12
#305940000000
0!
0%
b1 *
0-
02
b1 6
#305950000000
1!
1%
1-
12
#305960000000
0!
0%
b10 *
0-
02
b10 6
#305970000000
1!
1%
1-
12
#305980000000
0!
0%
b11 *
0-
02
b11 6
#305990000000
1!
1%
1-
12
15
#306000000000
0!
0%
b100 *
0-
02
b100 6
#306010000000
1!
1%
1-
12
#306020000000
0!
0%
b101 *
0-
02
b101 6
#306030000000
1!
1%
1-
12
#306040000000
0!
0%
b110 *
0-
02
b110 6
#306050000000
1!
1%
1-
12
#306060000000
0!
0%
b111 *
0-
02
b111 6
#306070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#306080000000
0!
0%
b0 *
0-
02
b0 6
#306090000000
1!
1%
1-
12
#306100000000
0!
0%
b1 *
0-
02
b1 6
#306110000000
1!
1%
1-
12
#306120000000
0!
0%
b10 *
0-
02
b10 6
#306130000000
1!
1%
1-
12
#306140000000
0!
0%
b11 *
0-
02
b11 6
#306150000000
1!
1%
1-
12
15
#306160000000
0!
0%
b100 *
0-
02
b100 6
#306170000000
1!
1%
1-
12
#306180000000
0!
0%
b101 *
0-
02
b101 6
#306190000000
1!
1%
1-
12
#306200000000
0!
0%
b110 *
0-
02
b110 6
#306210000000
1!
1%
1-
12
#306220000000
0!
0%
b111 *
0-
02
b111 6
#306230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#306240000000
0!
0%
b0 *
0-
02
b0 6
#306250000000
1!
1%
1-
12
#306260000000
0!
0%
b1 *
0-
02
b1 6
#306270000000
1!
1%
1-
12
#306280000000
0!
0%
b10 *
0-
02
b10 6
#306290000000
1!
1%
1-
12
#306300000000
0!
0%
b11 *
0-
02
b11 6
#306310000000
1!
1%
1-
12
15
#306320000000
0!
0%
b100 *
0-
02
b100 6
#306330000000
1!
1%
1-
12
#306340000000
0!
0%
b101 *
0-
02
b101 6
#306350000000
1!
1%
1-
12
#306360000000
0!
0%
b110 *
0-
02
b110 6
#306370000000
1!
1%
1-
12
#306380000000
0!
0%
b111 *
0-
02
b111 6
#306390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#306400000000
0!
0%
b0 *
0-
02
b0 6
#306410000000
1!
1%
1-
12
#306420000000
0!
0%
b1 *
0-
02
b1 6
#306430000000
1!
1%
1-
12
#306440000000
0!
0%
b10 *
0-
02
b10 6
#306450000000
1!
1%
1-
12
#306460000000
0!
0%
b11 *
0-
02
b11 6
#306470000000
1!
1%
1-
12
15
#306480000000
0!
0%
b100 *
0-
02
b100 6
#306490000000
1!
1%
1-
12
#306500000000
0!
0%
b101 *
0-
02
b101 6
#306510000000
1!
1%
1-
12
#306520000000
0!
0%
b110 *
0-
02
b110 6
#306530000000
1!
1%
1-
12
#306540000000
0!
0%
b111 *
0-
02
b111 6
#306550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#306560000000
0!
0%
b0 *
0-
02
b0 6
#306570000000
1!
1%
1-
12
#306580000000
0!
0%
b1 *
0-
02
b1 6
#306590000000
1!
1%
1-
12
#306600000000
0!
0%
b10 *
0-
02
b10 6
#306610000000
1!
1%
1-
12
#306620000000
0!
0%
b11 *
0-
02
b11 6
#306630000000
1!
1%
1-
12
15
#306640000000
0!
0%
b100 *
0-
02
b100 6
#306650000000
1!
1%
1-
12
#306660000000
0!
0%
b101 *
0-
02
b101 6
#306670000000
1!
1%
1-
12
#306680000000
0!
0%
b110 *
0-
02
b110 6
#306690000000
1!
1%
1-
12
#306700000000
0!
0%
b111 *
0-
02
b111 6
#306710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#306720000000
0!
0%
b0 *
0-
02
b0 6
#306730000000
1!
1%
1-
12
#306740000000
0!
0%
b1 *
0-
02
b1 6
#306750000000
1!
1%
1-
12
#306760000000
0!
0%
b10 *
0-
02
b10 6
#306770000000
1!
1%
1-
12
#306780000000
0!
0%
b11 *
0-
02
b11 6
#306790000000
1!
1%
1-
12
15
#306800000000
0!
0%
b100 *
0-
02
b100 6
#306810000000
1!
1%
1-
12
#306820000000
0!
0%
b101 *
0-
02
b101 6
#306830000000
1!
1%
1-
12
#306840000000
0!
0%
b110 *
0-
02
b110 6
#306850000000
1!
1%
1-
12
#306860000000
0!
0%
b111 *
0-
02
b111 6
#306870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#306880000000
0!
0%
b0 *
0-
02
b0 6
#306890000000
1!
1%
1-
12
#306900000000
0!
0%
b1 *
0-
02
b1 6
#306910000000
1!
1%
1-
12
#306920000000
0!
0%
b10 *
0-
02
b10 6
#306930000000
1!
1%
1-
12
#306940000000
0!
0%
b11 *
0-
02
b11 6
#306950000000
1!
1%
1-
12
15
#306960000000
0!
0%
b100 *
0-
02
b100 6
#306970000000
1!
1%
1-
12
#306980000000
0!
0%
b101 *
0-
02
b101 6
#306990000000
1!
1%
1-
12
#307000000000
0!
0%
b110 *
0-
02
b110 6
#307010000000
1!
1%
1-
12
#307020000000
0!
0%
b111 *
0-
02
b111 6
#307030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#307040000000
0!
0%
b0 *
0-
02
b0 6
#307050000000
1!
1%
1-
12
#307060000000
0!
0%
b1 *
0-
02
b1 6
#307070000000
1!
1%
1-
12
#307080000000
0!
0%
b10 *
0-
02
b10 6
#307090000000
1!
1%
1-
12
#307100000000
0!
0%
b11 *
0-
02
b11 6
#307110000000
1!
1%
1-
12
15
#307120000000
0!
0%
b100 *
0-
02
b100 6
#307130000000
1!
1%
1-
12
#307140000000
0!
0%
b101 *
0-
02
b101 6
#307150000000
1!
1%
1-
12
#307160000000
0!
0%
b110 *
0-
02
b110 6
#307170000000
1!
1%
1-
12
#307180000000
0!
0%
b111 *
0-
02
b111 6
#307190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#307200000000
0!
0%
b0 *
0-
02
b0 6
#307210000000
1!
1%
1-
12
#307220000000
0!
0%
b1 *
0-
02
b1 6
#307230000000
1!
1%
1-
12
#307240000000
0!
0%
b10 *
0-
02
b10 6
#307250000000
1!
1%
1-
12
#307260000000
0!
0%
b11 *
0-
02
b11 6
#307270000000
1!
1%
1-
12
15
#307280000000
0!
0%
b100 *
0-
02
b100 6
#307290000000
1!
1%
1-
12
#307300000000
0!
0%
b101 *
0-
02
b101 6
#307310000000
1!
1%
1-
12
#307320000000
0!
0%
b110 *
0-
02
b110 6
#307330000000
1!
1%
1-
12
#307340000000
0!
0%
b111 *
0-
02
b111 6
#307350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#307360000000
0!
0%
b0 *
0-
02
b0 6
#307370000000
1!
1%
1-
12
#307380000000
0!
0%
b1 *
0-
02
b1 6
#307390000000
1!
1%
1-
12
#307400000000
0!
0%
b10 *
0-
02
b10 6
#307410000000
1!
1%
1-
12
#307420000000
0!
0%
b11 *
0-
02
b11 6
#307430000000
1!
1%
1-
12
15
#307440000000
0!
0%
b100 *
0-
02
b100 6
#307450000000
1!
1%
1-
12
#307460000000
0!
0%
b101 *
0-
02
b101 6
#307470000000
1!
1%
1-
12
#307480000000
0!
0%
b110 *
0-
02
b110 6
#307490000000
1!
1%
1-
12
#307500000000
0!
0%
b111 *
0-
02
b111 6
#307510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#307520000000
0!
0%
b0 *
0-
02
b0 6
#307530000000
1!
1%
1-
12
#307540000000
0!
0%
b1 *
0-
02
b1 6
#307550000000
1!
1%
1-
12
#307560000000
0!
0%
b10 *
0-
02
b10 6
#307570000000
1!
1%
1-
12
#307580000000
0!
0%
b11 *
0-
02
b11 6
#307590000000
1!
1%
1-
12
15
#307600000000
0!
0%
b100 *
0-
02
b100 6
#307610000000
1!
1%
1-
12
#307620000000
0!
0%
b101 *
0-
02
b101 6
#307630000000
1!
1%
1-
12
#307640000000
0!
0%
b110 *
0-
02
b110 6
#307650000000
1!
1%
1-
12
#307660000000
0!
0%
b111 *
0-
02
b111 6
#307670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#307680000000
0!
0%
b0 *
0-
02
b0 6
#307690000000
1!
1%
1-
12
#307700000000
0!
0%
b1 *
0-
02
b1 6
#307710000000
1!
1%
1-
12
#307720000000
0!
0%
b10 *
0-
02
b10 6
#307730000000
1!
1%
1-
12
#307740000000
0!
0%
b11 *
0-
02
b11 6
#307750000000
1!
1%
1-
12
15
#307760000000
0!
0%
b100 *
0-
02
b100 6
#307770000000
1!
1%
1-
12
#307780000000
0!
0%
b101 *
0-
02
b101 6
#307790000000
1!
1%
1-
12
#307800000000
0!
0%
b110 *
0-
02
b110 6
#307810000000
1!
1%
1-
12
#307820000000
0!
0%
b111 *
0-
02
b111 6
#307830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#307840000000
0!
0%
b0 *
0-
02
b0 6
#307850000000
1!
1%
1-
12
#307860000000
0!
0%
b1 *
0-
02
b1 6
#307870000000
1!
1%
1-
12
#307880000000
0!
0%
b10 *
0-
02
b10 6
#307890000000
1!
1%
1-
12
#307900000000
0!
0%
b11 *
0-
02
b11 6
#307910000000
1!
1%
1-
12
15
#307920000000
0!
0%
b100 *
0-
02
b100 6
#307930000000
1!
1%
1-
12
#307940000000
0!
0%
b101 *
0-
02
b101 6
#307950000000
1!
1%
1-
12
#307960000000
0!
0%
b110 *
0-
02
b110 6
#307970000000
1!
1%
1-
12
#307980000000
0!
0%
b111 *
0-
02
b111 6
#307990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#308000000000
0!
0%
b0 *
0-
02
b0 6
#308010000000
1!
1%
1-
12
#308020000000
0!
0%
b1 *
0-
02
b1 6
#308030000000
1!
1%
1-
12
#308040000000
0!
0%
b10 *
0-
02
b10 6
#308050000000
1!
1%
1-
12
#308060000000
0!
0%
b11 *
0-
02
b11 6
#308070000000
1!
1%
1-
12
15
#308080000000
0!
0%
b100 *
0-
02
b100 6
#308090000000
1!
1%
1-
12
#308100000000
0!
0%
b101 *
0-
02
b101 6
#308110000000
1!
1%
1-
12
#308120000000
0!
0%
b110 *
0-
02
b110 6
#308130000000
1!
1%
1-
12
#308140000000
0!
0%
b111 *
0-
02
b111 6
#308150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#308160000000
0!
0%
b0 *
0-
02
b0 6
#308170000000
1!
1%
1-
12
#308180000000
0!
0%
b1 *
0-
02
b1 6
#308190000000
1!
1%
1-
12
#308200000000
0!
0%
b10 *
0-
02
b10 6
#308210000000
1!
1%
1-
12
#308220000000
0!
0%
b11 *
0-
02
b11 6
#308230000000
1!
1%
1-
12
15
#308240000000
0!
0%
b100 *
0-
02
b100 6
#308250000000
1!
1%
1-
12
#308260000000
0!
0%
b101 *
0-
02
b101 6
#308270000000
1!
1%
1-
12
#308280000000
0!
0%
b110 *
0-
02
b110 6
#308290000000
1!
1%
1-
12
#308300000000
0!
0%
b111 *
0-
02
b111 6
#308310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#308320000000
0!
0%
b0 *
0-
02
b0 6
#308330000000
1!
1%
1-
12
#308340000000
0!
0%
b1 *
0-
02
b1 6
#308350000000
1!
1%
1-
12
#308360000000
0!
0%
b10 *
0-
02
b10 6
#308370000000
1!
1%
1-
12
#308380000000
0!
0%
b11 *
0-
02
b11 6
#308390000000
1!
1%
1-
12
15
#308400000000
0!
0%
b100 *
0-
02
b100 6
#308410000000
1!
1%
1-
12
#308420000000
0!
0%
b101 *
0-
02
b101 6
#308430000000
1!
1%
1-
12
#308440000000
0!
0%
b110 *
0-
02
b110 6
#308450000000
1!
1%
1-
12
#308460000000
0!
0%
b111 *
0-
02
b111 6
#308470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#308480000000
0!
0%
b0 *
0-
02
b0 6
#308490000000
1!
1%
1-
12
#308500000000
0!
0%
b1 *
0-
02
b1 6
#308510000000
1!
1%
1-
12
#308520000000
0!
0%
b10 *
0-
02
b10 6
#308530000000
1!
1%
1-
12
#308540000000
0!
0%
b11 *
0-
02
b11 6
#308550000000
1!
1%
1-
12
15
#308560000000
0!
0%
b100 *
0-
02
b100 6
#308570000000
1!
1%
1-
12
#308580000000
0!
0%
b101 *
0-
02
b101 6
#308590000000
1!
1%
1-
12
#308600000000
0!
0%
b110 *
0-
02
b110 6
#308610000000
1!
1%
1-
12
#308620000000
0!
0%
b111 *
0-
02
b111 6
#308630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#308640000000
0!
0%
b0 *
0-
02
b0 6
#308650000000
1!
1%
1-
12
#308660000000
0!
0%
b1 *
0-
02
b1 6
#308670000000
1!
1%
1-
12
#308680000000
0!
0%
b10 *
0-
02
b10 6
#308690000000
1!
1%
1-
12
#308700000000
0!
0%
b11 *
0-
02
b11 6
#308710000000
1!
1%
1-
12
15
#308720000000
0!
0%
b100 *
0-
02
b100 6
#308730000000
1!
1%
1-
12
#308740000000
0!
0%
b101 *
0-
02
b101 6
#308750000000
1!
1%
1-
12
#308760000000
0!
0%
b110 *
0-
02
b110 6
#308770000000
1!
1%
1-
12
#308780000000
0!
0%
b111 *
0-
02
b111 6
#308790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#308800000000
0!
0%
b0 *
0-
02
b0 6
#308810000000
1!
1%
1-
12
#308820000000
0!
0%
b1 *
0-
02
b1 6
#308830000000
1!
1%
1-
12
#308840000000
0!
0%
b10 *
0-
02
b10 6
#308850000000
1!
1%
1-
12
#308860000000
0!
0%
b11 *
0-
02
b11 6
#308870000000
1!
1%
1-
12
15
#308880000000
0!
0%
b100 *
0-
02
b100 6
#308890000000
1!
1%
1-
12
#308900000000
0!
0%
b101 *
0-
02
b101 6
#308910000000
1!
1%
1-
12
#308920000000
0!
0%
b110 *
0-
02
b110 6
#308930000000
1!
1%
1-
12
#308940000000
0!
0%
b111 *
0-
02
b111 6
#308950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#308960000000
0!
0%
b0 *
0-
02
b0 6
#308970000000
1!
1%
1-
12
#308980000000
0!
0%
b1 *
0-
02
b1 6
#308990000000
1!
1%
1-
12
#309000000000
0!
0%
b10 *
0-
02
b10 6
#309010000000
1!
1%
1-
12
#309020000000
0!
0%
b11 *
0-
02
b11 6
#309030000000
1!
1%
1-
12
15
#309040000000
0!
0%
b100 *
0-
02
b100 6
#309050000000
1!
1%
1-
12
#309060000000
0!
0%
b101 *
0-
02
b101 6
#309070000000
1!
1%
1-
12
#309080000000
0!
0%
b110 *
0-
02
b110 6
#309090000000
1!
1%
1-
12
#309100000000
0!
0%
b111 *
0-
02
b111 6
#309110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#309120000000
0!
0%
b0 *
0-
02
b0 6
#309130000000
1!
1%
1-
12
#309140000000
0!
0%
b1 *
0-
02
b1 6
#309150000000
1!
1%
1-
12
#309160000000
0!
0%
b10 *
0-
02
b10 6
#309170000000
1!
1%
1-
12
#309180000000
0!
0%
b11 *
0-
02
b11 6
#309190000000
1!
1%
1-
12
15
#309200000000
0!
0%
b100 *
0-
02
b100 6
#309210000000
1!
1%
1-
12
#309220000000
0!
0%
b101 *
0-
02
b101 6
#309230000000
1!
1%
1-
12
#309240000000
0!
0%
b110 *
0-
02
b110 6
#309250000000
1!
1%
1-
12
#309260000000
0!
0%
b111 *
0-
02
b111 6
#309270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#309280000000
0!
0%
b0 *
0-
02
b0 6
#309290000000
1!
1%
1-
12
#309300000000
0!
0%
b1 *
0-
02
b1 6
#309310000000
1!
1%
1-
12
#309320000000
0!
0%
b10 *
0-
02
b10 6
#309330000000
1!
1%
1-
12
#309340000000
0!
0%
b11 *
0-
02
b11 6
#309350000000
1!
1%
1-
12
15
#309360000000
0!
0%
b100 *
0-
02
b100 6
#309370000000
1!
1%
1-
12
#309380000000
0!
0%
b101 *
0-
02
b101 6
#309390000000
1!
1%
1-
12
#309400000000
0!
0%
b110 *
0-
02
b110 6
#309410000000
1!
1%
1-
12
#309420000000
0!
0%
b111 *
0-
02
b111 6
#309430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#309440000000
0!
0%
b0 *
0-
02
b0 6
#309450000000
1!
1%
1-
12
#309460000000
0!
0%
b1 *
0-
02
b1 6
#309470000000
1!
1%
1-
12
#309480000000
0!
0%
b10 *
0-
02
b10 6
#309490000000
1!
1%
1-
12
#309500000000
0!
0%
b11 *
0-
02
b11 6
#309510000000
1!
1%
1-
12
15
#309520000000
0!
0%
b100 *
0-
02
b100 6
#309530000000
1!
1%
1-
12
#309540000000
0!
0%
b101 *
0-
02
b101 6
#309550000000
1!
1%
1-
12
#309560000000
0!
0%
b110 *
0-
02
b110 6
#309570000000
1!
1%
1-
12
#309580000000
0!
0%
b111 *
0-
02
b111 6
#309590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#309600000000
0!
0%
b0 *
0-
02
b0 6
#309610000000
1!
1%
1-
12
#309620000000
0!
0%
b1 *
0-
02
b1 6
#309630000000
1!
1%
1-
12
#309640000000
0!
0%
b10 *
0-
02
b10 6
#309650000000
1!
1%
1-
12
#309660000000
0!
0%
b11 *
0-
02
b11 6
#309670000000
1!
1%
1-
12
15
#309680000000
0!
0%
b100 *
0-
02
b100 6
#309690000000
1!
1%
1-
12
#309700000000
0!
0%
b101 *
0-
02
b101 6
#309710000000
1!
1%
1-
12
#309720000000
0!
0%
b110 *
0-
02
b110 6
#309730000000
1!
1%
1-
12
#309740000000
0!
0%
b111 *
0-
02
b111 6
#309750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#309760000000
0!
0%
b0 *
0-
02
b0 6
#309770000000
1!
1%
1-
12
#309780000000
0!
0%
b1 *
0-
02
b1 6
#309790000000
1!
1%
1-
12
#309800000000
0!
0%
b10 *
0-
02
b10 6
#309810000000
1!
1%
1-
12
#309820000000
0!
0%
b11 *
0-
02
b11 6
#309830000000
1!
1%
1-
12
15
#309840000000
0!
0%
b100 *
0-
02
b100 6
#309850000000
1!
1%
1-
12
#309860000000
0!
0%
b101 *
0-
02
b101 6
#309870000000
1!
1%
1-
12
#309880000000
0!
0%
b110 *
0-
02
b110 6
#309890000000
1!
1%
1-
12
#309900000000
0!
0%
b111 *
0-
02
b111 6
#309910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#309920000000
0!
0%
b0 *
0-
02
b0 6
#309930000000
1!
1%
1-
12
#309940000000
0!
0%
b1 *
0-
02
b1 6
#309950000000
1!
1%
1-
12
#309960000000
0!
0%
b10 *
0-
02
b10 6
#309970000000
1!
1%
1-
12
#309980000000
0!
0%
b11 *
0-
02
b11 6
#309990000000
1!
1%
1-
12
15
#310000000000
0!
0%
b100 *
0-
02
b100 6
#310010000000
1!
1%
1-
12
#310020000000
0!
0%
b101 *
0-
02
b101 6
#310030000000
1!
1%
1-
12
#310040000000
0!
0%
b110 *
0-
02
b110 6
#310050000000
1!
1%
1-
12
#310060000000
0!
0%
b111 *
0-
02
b111 6
#310070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#310080000000
0!
0%
b0 *
0-
02
b0 6
#310090000000
1!
1%
1-
12
#310100000000
0!
0%
b1 *
0-
02
b1 6
#310110000000
1!
1%
1-
12
#310120000000
0!
0%
b10 *
0-
02
b10 6
#310130000000
1!
1%
1-
12
#310140000000
0!
0%
b11 *
0-
02
b11 6
#310150000000
1!
1%
1-
12
15
#310160000000
0!
0%
b100 *
0-
02
b100 6
#310170000000
1!
1%
1-
12
#310180000000
0!
0%
b101 *
0-
02
b101 6
#310190000000
1!
1%
1-
12
#310200000000
0!
0%
b110 *
0-
02
b110 6
#310210000000
1!
1%
1-
12
#310220000000
0!
0%
b111 *
0-
02
b111 6
#310230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#310240000000
0!
0%
b0 *
0-
02
b0 6
#310250000000
1!
1%
1-
12
#310260000000
0!
0%
b1 *
0-
02
b1 6
#310270000000
1!
1%
1-
12
#310280000000
0!
0%
b10 *
0-
02
b10 6
#310290000000
1!
1%
1-
12
#310300000000
0!
0%
b11 *
0-
02
b11 6
#310310000000
1!
1%
1-
12
15
#310320000000
0!
0%
b100 *
0-
02
b100 6
#310330000000
1!
1%
1-
12
#310340000000
0!
0%
b101 *
0-
02
b101 6
#310350000000
1!
1%
1-
12
#310360000000
0!
0%
b110 *
0-
02
b110 6
#310370000000
1!
1%
1-
12
#310380000000
0!
0%
b111 *
0-
02
b111 6
#310390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#310400000000
0!
0%
b0 *
0-
02
b0 6
#310410000000
1!
1%
1-
12
#310420000000
0!
0%
b1 *
0-
02
b1 6
#310430000000
1!
1%
1-
12
#310440000000
0!
0%
b10 *
0-
02
b10 6
#310450000000
1!
1%
1-
12
#310460000000
0!
0%
b11 *
0-
02
b11 6
#310470000000
1!
1%
1-
12
15
#310480000000
0!
0%
b100 *
0-
02
b100 6
#310490000000
1!
1%
1-
12
#310500000000
0!
0%
b101 *
0-
02
b101 6
#310510000000
1!
1%
1-
12
#310520000000
0!
0%
b110 *
0-
02
b110 6
#310530000000
1!
1%
1-
12
#310540000000
0!
0%
b111 *
0-
02
b111 6
#310550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#310560000000
0!
0%
b0 *
0-
02
b0 6
#310570000000
1!
1%
1-
12
#310580000000
0!
0%
b1 *
0-
02
b1 6
#310590000000
1!
1%
1-
12
#310600000000
0!
0%
b10 *
0-
02
b10 6
#310610000000
1!
1%
1-
12
#310620000000
0!
0%
b11 *
0-
02
b11 6
#310630000000
1!
1%
1-
12
15
#310640000000
0!
0%
b100 *
0-
02
b100 6
#310650000000
1!
1%
1-
12
#310660000000
0!
0%
b101 *
0-
02
b101 6
#310670000000
1!
1%
1-
12
#310680000000
0!
0%
b110 *
0-
02
b110 6
#310690000000
1!
1%
1-
12
#310700000000
0!
0%
b111 *
0-
02
b111 6
#310710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#310720000000
0!
0%
b0 *
0-
02
b0 6
#310730000000
1!
1%
1-
12
#310740000000
0!
0%
b1 *
0-
02
b1 6
#310750000000
1!
1%
1-
12
#310760000000
0!
0%
b10 *
0-
02
b10 6
#310770000000
1!
1%
1-
12
#310780000000
0!
0%
b11 *
0-
02
b11 6
#310790000000
1!
1%
1-
12
15
#310800000000
0!
0%
b100 *
0-
02
b100 6
#310810000000
1!
1%
1-
12
#310820000000
0!
0%
b101 *
0-
02
b101 6
#310830000000
1!
1%
1-
12
#310840000000
0!
0%
b110 *
0-
02
b110 6
#310850000000
1!
1%
1-
12
#310860000000
0!
0%
b111 *
0-
02
b111 6
#310870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#310880000000
0!
0%
b0 *
0-
02
b0 6
#310890000000
1!
1%
1-
12
#310900000000
0!
0%
b1 *
0-
02
b1 6
#310910000000
1!
1%
1-
12
#310920000000
0!
0%
b10 *
0-
02
b10 6
#310930000000
1!
1%
1-
12
#310940000000
0!
0%
b11 *
0-
02
b11 6
#310950000000
1!
1%
1-
12
15
#310960000000
0!
0%
b100 *
0-
02
b100 6
#310970000000
1!
1%
1-
12
#310980000000
0!
0%
b101 *
0-
02
b101 6
#310990000000
1!
1%
1-
12
#311000000000
0!
0%
b110 *
0-
02
b110 6
#311010000000
1!
1%
1-
12
#311020000000
0!
0%
b111 *
0-
02
b111 6
#311030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#311040000000
0!
0%
b0 *
0-
02
b0 6
#311050000000
1!
1%
1-
12
#311060000000
0!
0%
b1 *
0-
02
b1 6
#311070000000
1!
1%
1-
12
#311080000000
0!
0%
b10 *
0-
02
b10 6
#311090000000
1!
1%
1-
12
#311100000000
0!
0%
b11 *
0-
02
b11 6
#311110000000
1!
1%
1-
12
15
#311120000000
0!
0%
b100 *
0-
02
b100 6
#311130000000
1!
1%
1-
12
#311140000000
0!
0%
b101 *
0-
02
b101 6
#311150000000
1!
1%
1-
12
#311160000000
0!
0%
b110 *
0-
02
b110 6
#311170000000
1!
1%
1-
12
#311180000000
0!
0%
b111 *
0-
02
b111 6
#311190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#311200000000
0!
0%
b0 *
0-
02
b0 6
#311210000000
1!
1%
1-
12
#311220000000
0!
0%
b1 *
0-
02
b1 6
#311230000000
1!
1%
1-
12
#311240000000
0!
0%
b10 *
0-
02
b10 6
#311250000000
1!
1%
1-
12
#311260000000
0!
0%
b11 *
0-
02
b11 6
#311270000000
1!
1%
1-
12
15
#311280000000
0!
0%
b100 *
0-
02
b100 6
#311290000000
1!
1%
1-
12
#311300000000
0!
0%
b101 *
0-
02
b101 6
#311310000000
1!
1%
1-
12
#311320000000
0!
0%
b110 *
0-
02
b110 6
#311330000000
1!
1%
1-
12
#311340000000
0!
0%
b111 *
0-
02
b111 6
#311350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#311360000000
0!
0%
b0 *
0-
02
b0 6
#311370000000
1!
1%
1-
12
#311380000000
0!
0%
b1 *
0-
02
b1 6
#311390000000
1!
1%
1-
12
#311400000000
0!
0%
b10 *
0-
02
b10 6
#311410000000
1!
1%
1-
12
#311420000000
0!
0%
b11 *
0-
02
b11 6
#311430000000
1!
1%
1-
12
15
#311440000000
0!
0%
b100 *
0-
02
b100 6
#311450000000
1!
1%
1-
12
#311460000000
0!
0%
b101 *
0-
02
b101 6
#311470000000
1!
1%
1-
12
#311480000000
0!
0%
b110 *
0-
02
b110 6
#311490000000
1!
1%
1-
12
#311500000000
0!
0%
b111 *
0-
02
b111 6
#311510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#311520000000
0!
0%
b0 *
0-
02
b0 6
#311530000000
1!
1%
1-
12
#311540000000
0!
0%
b1 *
0-
02
b1 6
#311550000000
1!
1%
1-
12
#311560000000
0!
0%
b10 *
0-
02
b10 6
#311570000000
1!
1%
1-
12
#311580000000
0!
0%
b11 *
0-
02
b11 6
#311590000000
1!
1%
1-
12
15
#311600000000
0!
0%
b100 *
0-
02
b100 6
#311610000000
1!
1%
1-
12
#311620000000
0!
0%
b101 *
0-
02
b101 6
#311630000000
1!
1%
1-
12
#311640000000
0!
0%
b110 *
0-
02
b110 6
#311650000000
1!
1%
1-
12
#311660000000
0!
0%
b111 *
0-
02
b111 6
#311670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#311680000000
0!
0%
b0 *
0-
02
b0 6
#311690000000
1!
1%
1-
12
#311700000000
0!
0%
b1 *
0-
02
b1 6
#311710000000
1!
1%
1-
12
#311720000000
0!
0%
b10 *
0-
02
b10 6
#311730000000
1!
1%
1-
12
#311740000000
0!
0%
b11 *
0-
02
b11 6
#311750000000
1!
1%
1-
12
15
#311760000000
0!
0%
b100 *
0-
02
b100 6
#311770000000
1!
1%
1-
12
#311780000000
0!
0%
b101 *
0-
02
b101 6
#311790000000
1!
1%
1-
12
#311800000000
0!
0%
b110 *
0-
02
b110 6
#311810000000
1!
1%
1-
12
#311820000000
0!
0%
b111 *
0-
02
b111 6
#311830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#311840000000
0!
0%
b0 *
0-
02
b0 6
#311850000000
1!
1%
1-
12
#311860000000
0!
0%
b1 *
0-
02
b1 6
#311870000000
1!
1%
1-
12
#311880000000
0!
0%
b10 *
0-
02
b10 6
#311890000000
1!
1%
1-
12
#311900000000
0!
0%
b11 *
0-
02
b11 6
#311910000000
1!
1%
1-
12
15
#311920000000
0!
0%
b100 *
0-
02
b100 6
#311930000000
1!
1%
1-
12
#311940000000
0!
0%
b101 *
0-
02
b101 6
#311950000000
1!
1%
1-
12
#311960000000
0!
0%
b110 *
0-
02
b110 6
#311970000000
1!
1%
1-
12
#311980000000
0!
0%
b111 *
0-
02
b111 6
#311990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#312000000000
0!
0%
b0 *
0-
02
b0 6
#312010000000
1!
1%
1-
12
#312020000000
0!
0%
b1 *
0-
02
b1 6
#312030000000
1!
1%
1-
12
#312040000000
0!
0%
b10 *
0-
02
b10 6
#312050000000
1!
1%
1-
12
#312060000000
0!
0%
b11 *
0-
02
b11 6
#312070000000
1!
1%
1-
12
15
#312080000000
0!
0%
b100 *
0-
02
b100 6
#312090000000
1!
1%
1-
12
#312100000000
0!
0%
b101 *
0-
02
b101 6
#312110000000
1!
1%
1-
12
#312120000000
0!
0%
b110 *
0-
02
b110 6
#312130000000
1!
1%
1-
12
#312140000000
0!
0%
b111 *
0-
02
b111 6
#312150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#312160000000
0!
0%
b0 *
0-
02
b0 6
#312170000000
1!
1%
1-
12
#312180000000
0!
0%
b1 *
0-
02
b1 6
#312190000000
1!
1%
1-
12
#312200000000
0!
0%
b10 *
0-
02
b10 6
#312210000000
1!
1%
1-
12
#312220000000
0!
0%
b11 *
0-
02
b11 6
#312230000000
1!
1%
1-
12
15
#312240000000
0!
0%
b100 *
0-
02
b100 6
#312250000000
1!
1%
1-
12
#312260000000
0!
0%
b101 *
0-
02
b101 6
#312270000000
1!
1%
1-
12
#312280000000
0!
0%
b110 *
0-
02
b110 6
#312290000000
1!
1%
1-
12
#312300000000
0!
0%
b111 *
0-
02
b111 6
#312310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#312320000000
0!
0%
b0 *
0-
02
b0 6
#312330000000
1!
1%
1-
12
#312340000000
0!
0%
b1 *
0-
02
b1 6
#312350000000
1!
1%
1-
12
#312360000000
0!
0%
b10 *
0-
02
b10 6
#312370000000
1!
1%
1-
12
#312380000000
0!
0%
b11 *
0-
02
b11 6
#312390000000
1!
1%
1-
12
15
#312400000000
0!
0%
b100 *
0-
02
b100 6
#312410000000
1!
1%
1-
12
#312420000000
0!
0%
b101 *
0-
02
b101 6
#312430000000
1!
1%
1-
12
#312440000000
0!
0%
b110 *
0-
02
b110 6
#312450000000
1!
1%
1-
12
#312460000000
0!
0%
b111 *
0-
02
b111 6
#312470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#312480000000
0!
0%
b0 *
0-
02
b0 6
#312490000000
1!
1%
1-
12
#312500000000
0!
0%
b1 *
0-
02
b1 6
#312510000000
1!
1%
1-
12
#312520000000
0!
0%
b10 *
0-
02
b10 6
#312530000000
1!
1%
1-
12
#312540000000
0!
0%
b11 *
0-
02
b11 6
#312550000000
1!
1%
1-
12
15
#312560000000
0!
0%
b100 *
0-
02
b100 6
#312570000000
1!
1%
1-
12
#312580000000
0!
0%
b101 *
0-
02
b101 6
#312590000000
1!
1%
1-
12
#312600000000
0!
0%
b110 *
0-
02
b110 6
#312610000000
1!
1%
1-
12
#312620000000
0!
0%
b111 *
0-
02
b111 6
#312630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#312640000000
0!
0%
b0 *
0-
02
b0 6
#312650000000
1!
1%
1-
12
#312660000000
0!
0%
b1 *
0-
02
b1 6
#312670000000
1!
1%
1-
12
#312680000000
0!
0%
b10 *
0-
02
b10 6
#312690000000
1!
1%
1-
12
#312700000000
0!
0%
b11 *
0-
02
b11 6
#312710000000
1!
1%
1-
12
15
#312720000000
0!
0%
b100 *
0-
02
b100 6
#312730000000
1!
1%
1-
12
#312740000000
0!
0%
b101 *
0-
02
b101 6
#312750000000
1!
1%
1-
12
#312760000000
0!
0%
b110 *
0-
02
b110 6
#312770000000
1!
1%
1-
12
#312780000000
0!
0%
b111 *
0-
02
b111 6
#312790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#312800000000
0!
0%
b0 *
0-
02
b0 6
#312810000000
1!
1%
1-
12
#312820000000
0!
0%
b1 *
0-
02
b1 6
#312830000000
1!
1%
1-
12
#312840000000
0!
0%
b10 *
0-
02
b10 6
#312850000000
1!
1%
1-
12
#312860000000
0!
0%
b11 *
0-
02
b11 6
#312870000000
1!
1%
1-
12
15
#312880000000
0!
0%
b100 *
0-
02
b100 6
#312890000000
1!
1%
1-
12
#312900000000
0!
0%
b101 *
0-
02
b101 6
#312910000000
1!
1%
1-
12
#312920000000
0!
0%
b110 *
0-
02
b110 6
#312930000000
1!
1%
1-
12
#312940000000
0!
0%
b111 *
0-
02
b111 6
#312950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#312960000000
0!
0%
b0 *
0-
02
b0 6
#312970000000
1!
1%
1-
12
#312980000000
0!
0%
b1 *
0-
02
b1 6
#312990000000
1!
1%
1-
12
#313000000000
0!
0%
b10 *
0-
02
b10 6
#313010000000
1!
1%
1-
12
#313020000000
0!
0%
b11 *
0-
02
b11 6
#313030000000
1!
1%
1-
12
15
#313040000000
0!
0%
b100 *
0-
02
b100 6
#313050000000
1!
1%
1-
12
#313060000000
0!
0%
b101 *
0-
02
b101 6
#313070000000
1!
1%
1-
12
#313080000000
0!
0%
b110 *
0-
02
b110 6
#313090000000
1!
1%
1-
12
#313100000000
0!
0%
b111 *
0-
02
b111 6
#313110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#313120000000
0!
0%
b0 *
0-
02
b0 6
#313130000000
1!
1%
1-
12
#313140000000
0!
0%
b1 *
0-
02
b1 6
#313150000000
1!
1%
1-
12
#313160000000
0!
0%
b10 *
0-
02
b10 6
#313170000000
1!
1%
1-
12
#313180000000
0!
0%
b11 *
0-
02
b11 6
#313190000000
1!
1%
1-
12
15
#313200000000
0!
0%
b100 *
0-
02
b100 6
#313210000000
1!
1%
1-
12
#313220000000
0!
0%
b101 *
0-
02
b101 6
#313230000000
1!
1%
1-
12
#313240000000
0!
0%
b110 *
0-
02
b110 6
#313250000000
1!
1%
1-
12
#313260000000
0!
0%
b111 *
0-
02
b111 6
#313270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#313280000000
0!
0%
b0 *
0-
02
b0 6
#313290000000
1!
1%
1-
12
#313300000000
0!
0%
b1 *
0-
02
b1 6
#313310000000
1!
1%
1-
12
#313320000000
0!
0%
b10 *
0-
02
b10 6
#313330000000
1!
1%
1-
12
#313340000000
0!
0%
b11 *
0-
02
b11 6
#313350000000
1!
1%
1-
12
15
#313360000000
0!
0%
b100 *
0-
02
b100 6
#313370000000
1!
1%
1-
12
#313380000000
0!
0%
b101 *
0-
02
b101 6
#313390000000
1!
1%
1-
12
#313400000000
0!
0%
b110 *
0-
02
b110 6
#313410000000
1!
1%
1-
12
#313420000000
0!
0%
b111 *
0-
02
b111 6
#313430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#313440000000
0!
0%
b0 *
0-
02
b0 6
#313450000000
1!
1%
1-
12
#313460000000
0!
0%
b1 *
0-
02
b1 6
#313470000000
1!
1%
1-
12
#313480000000
0!
0%
b10 *
0-
02
b10 6
#313490000000
1!
1%
1-
12
#313500000000
0!
0%
b11 *
0-
02
b11 6
#313510000000
1!
1%
1-
12
15
#313520000000
0!
0%
b100 *
0-
02
b100 6
#313530000000
1!
1%
1-
12
#313540000000
0!
0%
b101 *
0-
02
b101 6
#313550000000
1!
1%
1-
12
#313560000000
0!
0%
b110 *
0-
02
b110 6
#313570000000
1!
1%
1-
12
#313580000000
0!
0%
b111 *
0-
02
b111 6
#313590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#313600000000
0!
0%
b0 *
0-
02
b0 6
#313610000000
1!
1%
1-
12
#313620000000
0!
0%
b1 *
0-
02
b1 6
#313630000000
1!
1%
1-
12
#313640000000
0!
0%
b10 *
0-
02
b10 6
#313650000000
1!
1%
1-
12
#313660000000
0!
0%
b11 *
0-
02
b11 6
#313670000000
1!
1%
1-
12
15
#313680000000
0!
0%
b100 *
0-
02
b100 6
#313690000000
1!
1%
1-
12
#313700000000
0!
0%
b101 *
0-
02
b101 6
#313710000000
1!
1%
1-
12
#313720000000
0!
0%
b110 *
0-
02
b110 6
#313730000000
1!
1%
1-
12
#313740000000
0!
0%
b111 *
0-
02
b111 6
#313750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#313760000000
0!
0%
b0 *
0-
02
b0 6
#313770000000
1!
1%
1-
12
#313780000000
0!
0%
b1 *
0-
02
b1 6
#313790000000
1!
1%
1-
12
#313800000000
0!
0%
b10 *
0-
02
b10 6
#313810000000
1!
1%
1-
12
#313820000000
0!
0%
b11 *
0-
02
b11 6
#313830000000
1!
1%
1-
12
15
#313840000000
0!
0%
b100 *
0-
02
b100 6
#313850000000
1!
1%
1-
12
#313860000000
0!
0%
b101 *
0-
02
b101 6
#313870000000
1!
1%
1-
12
#313880000000
0!
0%
b110 *
0-
02
b110 6
#313890000000
1!
1%
1-
12
#313900000000
0!
0%
b111 *
0-
02
b111 6
#313910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#313920000000
0!
0%
b0 *
0-
02
b0 6
#313930000000
1!
1%
1-
12
#313940000000
0!
0%
b1 *
0-
02
b1 6
#313950000000
1!
1%
1-
12
#313960000000
0!
0%
b10 *
0-
02
b10 6
#313970000000
1!
1%
1-
12
#313980000000
0!
0%
b11 *
0-
02
b11 6
#313990000000
1!
1%
1-
12
15
#314000000000
0!
0%
b100 *
0-
02
b100 6
#314010000000
1!
1%
1-
12
#314020000000
0!
0%
b101 *
0-
02
b101 6
#314030000000
1!
1%
1-
12
#314040000000
0!
0%
b110 *
0-
02
b110 6
#314050000000
1!
1%
1-
12
#314060000000
0!
0%
b111 *
0-
02
b111 6
#314070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#314080000000
0!
0%
b0 *
0-
02
b0 6
#314090000000
1!
1%
1-
12
#314100000000
0!
0%
b1 *
0-
02
b1 6
#314110000000
1!
1%
1-
12
#314120000000
0!
0%
b10 *
0-
02
b10 6
#314130000000
1!
1%
1-
12
#314140000000
0!
0%
b11 *
0-
02
b11 6
#314150000000
1!
1%
1-
12
15
#314160000000
0!
0%
b100 *
0-
02
b100 6
#314170000000
1!
1%
1-
12
#314180000000
0!
0%
b101 *
0-
02
b101 6
#314190000000
1!
1%
1-
12
#314200000000
0!
0%
b110 *
0-
02
b110 6
#314210000000
1!
1%
1-
12
#314220000000
0!
0%
b111 *
0-
02
b111 6
#314230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#314240000000
0!
0%
b0 *
0-
02
b0 6
#314250000000
1!
1%
1-
12
#314260000000
0!
0%
b1 *
0-
02
b1 6
#314270000000
1!
1%
1-
12
#314280000000
0!
0%
b10 *
0-
02
b10 6
#314290000000
1!
1%
1-
12
#314300000000
0!
0%
b11 *
0-
02
b11 6
#314310000000
1!
1%
1-
12
15
#314320000000
0!
0%
b100 *
0-
02
b100 6
#314330000000
1!
1%
1-
12
#314340000000
0!
0%
b101 *
0-
02
b101 6
#314350000000
1!
1%
1-
12
#314360000000
0!
0%
b110 *
0-
02
b110 6
#314370000000
1!
1%
1-
12
#314380000000
0!
0%
b111 *
0-
02
b111 6
#314390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#314400000000
0!
0%
b0 *
0-
02
b0 6
#314410000000
1!
1%
1-
12
#314420000000
0!
0%
b1 *
0-
02
b1 6
#314430000000
1!
1%
1-
12
#314440000000
0!
0%
b10 *
0-
02
b10 6
#314450000000
1!
1%
1-
12
#314460000000
0!
0%
b11 *
0-
02
b11 6
#314470000000
1!
1%
1-
12
15
#314480000000
0!
0%
b100 *
0-
02
b100 6
#314490000000
1!
1%
1-
12
#314500000000
0!
0%
b101 *
0-
02
b101 6
#314510000000
1!
1%
1-
12
#314520000000
0!
0%
b110 *
0-
02
b110 6
#314530000000
1!
1%
1-
12
#314540000000
0!
0%
b111 *
0-
02
b111 6
#314550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#314560000000
0!
0%
b0 *
0-
02
b0 6
#314570000000
1!
1%
1-
12
#314580000000
0!
0%
b1 *
0-
02
b1 6
#314590000000
1!
1%
1-
12
#314600000000
0!
0%
b10 *
0-
02
b10 6
#314610000000
1!
1%
1-
12
#314620000000
0!
0%
b11 *
0-
02
b11 6
#314630000000
1!
1%
1-
12
15
#314640000000
0!
0%
b100 *
0-
02
b100 6
#314650000000
1!
1%
1-
12
#314660000000
0!
0%
b101 *
0-
02
b101 6
#314670000000
1!
1%
1-
12
#314680000000
0!
0%
b110 *
0-
02
b110 6
#314690000000
1!
1%
1-
12
#314700000000
0!
0%
b111 *
0-
02
b111 6
#314710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#314720000000
0!
0%
b0 *
0-
02
b0 6
#314730000000
1!
1%
1-
12
#314740000000
0!
0%
b1 *
0-
02
b1 6
#314750000000
1!
1%
1-
12
#314760000000
0!
0%
b10 *
0-
02
b10 6
#314770000000
1!
1%
1-
12
#314780000000
0!
0%
b11 *
0-
02
b11 6
#314790000000
1!
1%
1-
12
15
#314800000000
0!
0%
b100 *
0-
02
b100 6
#314810000000
1!
1%
1-
12
#314820000000
0!
0%
b101 *
0-
02
b101 6
#314830000000
1!
1%
1-
12
#314840000000
0!
0%
b110 *
0-
02
b110 6
#314850000000
1!
1%
1-
12
#314860000000
0!
0%
b111 *
0-
02
b111 6
#314870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#314880000000
0!
0%
b0 *
0-
02
b0 6
#314890000000
1!
1%
1-
12
#314900000000
0!
0%
b1 *
0-
02
b1 6
#314910000000
1!
1%
1-
12
#314920000000
0!
0%
b10 *
0-
02
b10 6
#314930000000
1!
1%
1-
12
#314940000000
0!
0%
b11 *
0-
02
b11 6
#314950000000
1!
1%
1-
12
15
#314960000000
0!
0%
b100 *
0-
02
b100 6
#314970000000
1!
1%
1-
12
#314980000000
0!
0%
b101 *
0-
02
b101 6
#314990000000
1!
1%
1-
12
#315000000000
0!
0%
b110 *
0-
02
b110 6
#315010000000
1!
1%
1-
12
#315020000000
0!
0%
b111 *
0-
02
b111 6
#315030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#315040000000
0!
0%
b0 *
0-
02
b0 6
#315050000000
1!
1%
1-
12
#315060000000
0!
0%
b1 *
0-
02
b1 6
#315070000000
1!
1%
1-
12
#315080000000
0!
0%
b10 *
0-
02
b10 6
#315090000000
1!
1%
1-
12
#315100000000
0!
0%
b11 *
0-
02
b11 6
#315110000000
1!
1%
1-
12
15
#315120000000
0!
0%
b100 *
0-
02
b100 6
#315130000000
1!
1%
1-
12
#315140000000
0!
0%
b101 *
0-
02
b101 6
#315150000000
1!
1%
1-
12
#315160000000
0!
0%
b110 *
0-
02
b110 6
#315170000000
1!
1%
1-
12
#315180000000
0!
0%
b111 *
0-
02
b111 6
#315190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#315200000000
0!
0%
b0 *
0-
02
b0 6
#315210000000
1!
1%
1-
12
#315220000000
0!
0%
b1 *
0-
02
b1 6
#315230000000
1!
1%
1-
12
#315240000000
0!
0%
b10 *
0-
02
b10 6
#315250000000
1!
1%
1-
12
#315260000000
0!
0%
b11 *
0-
02
b11 6
#315270000000
1!
1%
1-
12
15
#315280000000
0!
0%
b100 *
0-
02
b100 6
#315290000000
1!
1%
1-
12
#315300000000
0!
0%
b101 *
0-
02
b101 6
#315310000000
1!
1%
1-
12
#315320000000
0!
0%
b110 *
0-
02
b110 6
#315330000000
1!
1%
1-
12
#315340000000
0!
0%
b111 *
0-
02
b111 6
#315350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#315360000000
0!
0%
b0 *
0-
02
b0 6
#315370000000
1!
1%
1-
12
#315380000000
0!
0%
b1 *
0-
02
b1 6
#315390000000
1!
1%
1-
12
#315400000000
0!
0%
b10 *
0-
02
b10 6
#315410000000
1!
1%
1-
12
#315420000000
0!
0%
b11 *
0-
02
b11 6
#315430000000
1!
1%
1-
12
15
#315440000000
0!
0%
b100 *
0-
02
b100 6
#315450000000
1!
1%
1-
12
#315460000000
0!
0%
b101 *
0-
02
b101 6
#315470000000
1!
1%
1-
12
#315480000000
0!
0%
b110 *
0-
02
b110 6
#315490000000
1!
1%
1-
12
#315500000000
0!
0%
b111 *
0-
02
b111 6
#315510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#315520000000
0!
0%
b0 *
0-
02
b0 6
#315530000000
1!
1%
1-
12
#315540000000
0!
0%
b1 *
0-
02
b1 6
#315550000000
1!
1%
1-
12
#315560000000
0!
0%
b10 *
0-
02
b10 6
#315570000000
1!
1%
1-
12
#315580000000
0!
0%
b11 *
0-
02
b11 6
#315590000000
1!
1%
1-
12
15
#315600000000
0!
0%
b100 *
0-
02
b100 6
#315610000000
1!
1%
1-
12
#315620000000
0!
0%
b101 *
0-
02
b101 6
#315630000000
1!
1%
1-
12
#315640000000
0!
0%
b110 *
0-
02
b110 6
#315650000000
1!
1%
1-
12
#315660000000
0!
0%
b111 *
0-
02
b111 6
#315670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#315680000000
0!
0%
b0 *
0-
02
b0 6
#315690000000
1!
1%
1-
12
#315700000000
0!
0%
b1 *
0-
02
b1 6
#315710000000
1!
1%
1-
12
#315720000000
0!
0%
b10 *
0-
02
b10 6
#315730000000
1!
1%
1-
12
#315740000000
0!
0%
b11 *
0-
02
b11 6
#315750000000
1!
1%
1-
12
15
#315760000000
0!
0%
b100 *
0-
02
b100 6
#315770000000
1!
1%
1-
12
#315780000000
0!
0%
b101 *
0-
02
b101 6
#315790000000
1!
1%
1-
12
#315800000000
0!
0%
b110 *
0-
02
b110 6
#315810000000
1!
1%
1-
12
#315820000000
0!
0%
b111 *
0-
02
b111 6
#315830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#315840000000
0!
0%
b0 *
0-
02
b0 6
#315850000000
1!
1%
1-
12
#315860000000
0!
0%
b1 *
0-
02
b1 6
#315870000000
1!
1%
1-
12
#315880000000
0!
0%
b10 *
0-
02
b10 6
#315890000000
1!
1%
1-
12
#315900000000
0!
0%
b11 *
0-
02
b11 6
#315910000000
1!
1%
1-
12
15
#315920000000
0!
0%
b100 *
0-
02
b100 6
#315930000000
1!
1%
1-
12
#315940000000
0!
0%
b101 *
0-
02
b101 6
#315950000000
1!
1%
1-
12
#315960000000
0!
0%
b110 *
0-
02
b110 6
#315970000000
1!
1%
1-
12
#315980000000
0!
0%
b111 *
0-
02
b111 6
#315990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#316000000000
0!
0%
b0 *
0-
02
b0 6
#316010000000
1!
1%
1-
12
#316020000000
0!
0%
b1 *
0-
02
b1 6
#316030000000
1!
1%
1-
12
#316040000000
0!
0%
b10 *
0-
02
b10 6
#316050000000
1!
1%
1-
12
#316060000000
0!
0%
b11 *
0-
02
b11 6
#316070000000
1!
1%
1-
12
15
#316080000000
0!
0%
b100 *
0-
02
b100 6
#316090000000
1!
1%
1-
12
#316100000000
0!
0%
b101 *
0-
02
b101 6
#316110000000
1!
1%
1-
12
#316120000000
0!
0%
b110 *
0-
02
b110 6
#316130000000
1!
1%
1-
12
#316140000000
0!
0%
b111 *
0-
02
b111 6
#316150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#316160000000
0!
0%
b0 *
0-
02
b0 6
#316170000000
1!
1%
1-
12
#316180000000
0!
0%
b1 *
0-
02
b1 6
#316190000000
1!
1%
1-
12
#316200000000
0!
0%
b10 *
0-
02
b10 6
#316210000000
1!
1%
1-
12
#316220000000
0!
0%
b11 *
0-
02
b11 6
#316230000000
1!
1%
1-
12
15
#316240000000
0!
0%
b100 *
0-
02
b100 6
#316250000000
1!
1%
1-
12
#316260000000
0!
0%
b101 *
0-
02
b101 6
#316270000000
1!
1%
1-
12
#316280000000
0!
0%
b110 *
0-
02
b110 6
#316290000000
1!
1%
1-
12
#316300000000
0!
0%
b111 *
0-
02
b111 6
#316310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#316320000000
0!
0%
b0 *
0-
02
b0 6
#316330000000
1!
1%
1-
12
#316340000000
0!
0%
b1 *
0-
02
b1 6
#316350000000
1!
1%
1-
12
#316360000000
0!
0%
b10 *
0-
02
b10 6
#316370000000
1!
1%
1-
12
#316380000000
0!
0%
b11 *
0-
02
b11 6
#316390000000
1!
1%
1-
12
15
#316400000000
0!
0%
b100 *
0-
02
b100 6
#316410000000
1!
1%
1-
12
#316420000000
0!
0%
b101 *
0-
02
b101 6
#316430000000
1!
1%
1-
12
#316440000000
0!
0%
b110 *
0-
02
b110 6
#316450000000
1!
1%
1-
12
#316460000000
0!
0%
b111 *
0-
02
b111 6
#316470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#316480000000
0!
0%
b0 *
0-
02
b0 6
#316490000000
1!
1%
1-
12
#316500000000
0!
0%
b1 *
0-
02
b1 6
#316510000000
1!
1%
1-
12
#316520000000
0!
0%
b10 *
0-
02
b10 6
#316530000000
1!
1%
1-
12
#316540000000
0!
0%
b11 *
0-
02
b11 6
#316550000000
1!
1%
1-
12
15
#316560000000
0!
0%
b100 *
0-
02
b100 6
#316570000000
1!
1%
1-
12
#316580000000
0!
0%
b101 *
0-
02
b101 6
#316590000000
1!
1%
1-
12
#316600000000
0!
0%
b110 *
0-
02
b110 6
#316610000000
1!
1%
1-
12
#316620000000
0!
0%
b111 *
0-
02
b111 6
#316630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#316640000000
0!
0%
b0 *
0-
02
b0 6
#316650000000
1!
1%
1-
12
#316660000000
0!
0%
b1 *
0-
02
b1 6
#316670000000
1!
1%
1-
12
#316680000000
0!
0%
b10 *
0-
02
b10 6
#316690000000
1!
1%
1-
12
#316700000000
0!
0%
b11 *
0-
02
b11 6
#316710000000
1!
1%
1-
12
15
#316720000000
0!
0%
b100 *
0-
02
b100 6
#316730000000
1!
1%
1-
12
#316740000000
0!
0%
b101 *
0-
02
b101 6
#316750000000
1!
1%
1-
12
#316760000000
0!
0%
b110 *
0-
02
b110 6
#316770000000
1!
1%
1-
12
#316780000000
0!
0%
b111 *
0-
02
b111 6
#316790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#316800000000
0!
0%
b0 *
0-
02
b0 6
#316810000000
1!
1%
1-
12
#316820000000
0!
0%
b1 *
0-
02
b1 6
#316830000000
1!
1%
1-
12
#316840000000
0!
0%
b10 *
0-
02
b10 6
#316850000000
1!
1%
1-
12
#316860000000
0!
0%
b11 *
0-
02
b11 6
#316870000000
1!
1%
1-
12
15
#316880000000
0!
0%
b100 *
0-
02
b100 6
#316890000000
1!
1%
1-
12
#316900000000
0!
0%
b101 *
0-
02
b101 6
#316910000000
1!
1%
1-
12
#316920000000
0!
0%
b110 *
0-
02
b110 6
#316930000000
1!
1%
1-
12
#316940000000
0!
0%
b111 *
0-
02
b111 6
#316950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#316960000000
0!
0%
b0 *
0-
02
b0 6
#316970000000
1!
1%
1-
12
#316980000000
0!
0%
b1 *
0-
02
b1 6
#316990000000
1!
1%
1-
12
#317000000000
0!
0%
b10 *
0-
02
b10 6
#317010000000
1!
1%
1-
12
#317020000000
0!
0%
b11 *
0-
02
b11 6
#317030000000
1!
1%
1-
12
15
#317040000000
0!
0%
b100 *
0-
02
b100 6
#317050000000
1!
1%
1-
12
#317060000000
0!
0%
b101 *
0-
02
b101 6
#317070000000
1!
1%
1-
12
#317080000000
0!
0%
b110 *
0-
02
b110 6
#317090000000
1!
1%
1-
12
#317100000000
0!
0%
b111 *
0-
02
b111 6
#317110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#317120000000
0!
0%
b0 *
0-
02
b0 6
#317130000000
1!
1%
1-
12
#317140000000
0!
0%
b1 *
0-
02
b1 6
#317150000000
1!
1%
1-
12
#317160000000
0!
0%
b10 *
0-
02
b10 6
#317170000000
1!
1%
1-
12
#317180000000
0!
0%
b11 *
0-
02
b11 6
#317190000000
1!
1%
1-
12
15
#317200000000
0!
0%
b100 *
0-
02
b100 6
#317210000000
1!
1%
1-
12
#317220000000
0!
0%
b101 *
0-
02
b101 6
#317230000000
1!
1%
1-
12
#317240000000
0!
0%
b110 *
0-
02
b110 6
#317250000000
1!
1%
1-
12
#317260000000
0!
0%
b111 *
0-
02
b111 6
#317270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#317280000000
0!
0%
b0 *
0-
02
b0 6
#317290000000
1!
1%
1-
12
#317300000000
0!
0%
b1 *
0-
02
b1 6
#317310000000
1!
1%
1-
12
#317320000000
0!
0%
b10 *
0-
02
b10 6
#317330000000
1!
1%
1-
12
#317340000000
0!
0%
b11 *
0-
02
b11 6
#317350000000
1!
1%
1-
12
15
#317360000000
0!
0%
b100 *
0-
02
b100 6
#317370000000
1!
1%
1-
12
#317380000000
0!
0%
b101 *
0-
02
b101 6
#317390000000
1!
1%
1-
12
#317400000000
0!
0%
b110 *
0-
02
b110 6
#317410000000
1!
1%
1-
12
#317420000000
0!
0%
b111 *
0-
02
b111 6
#317430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#317440000000
0!
0%
b0 *
0-
02
b0 6
#317450000000
1!
1%
1-
12
#317460000000
0!
0%
b1 *
0-
02
b1 6
#317470000000
1!
1%
1-
12
#317480000000
0!
0%
b10 *
0-
02
b10 6
#317490000000
1!
1%
1-
12
#317500000000
0!
0%
b11 *
0-
02
b11 6
#317510000000
1!
1%
1-
12
15
#317520000000
0!
0%
b100 *
0-
02
b100 6
#317530000000
1!
1%
1-
12
#317540000000
0!
0%
b101 *
0-
02
b101 6
#317550000000
1!
1%
1-
12
#317560000000
0!
0%
b110 *
0-
02
b110 6
#317570000000
1!
1%
1-
12
#317580000000
0!
0%
b111 *
0-
02
b111 6
#317590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#317600000000
0!
0%
b0 *
0-
02
b0 6
#317610000000
1!
1%
1-
12
#317620000000
0!
0%
b1 *
0-
02
b1 6
#317630000000
1!
1%
1-
12
#317640000000
0!
0%
b10 *
0-
02
b10 6
#317650000000
1!
1%
1-
12
#317660000000
0!
0%
b11 *
0-
02
b11 6
#317670000000
1!
1%
1-
12
15
#317680000000
0!
0%
b100 *
0-
02
b100 6
#317690000000
1!
1%
1-
12
#317700000000
0!
0%
b101 *
0-
02
b101 6
#317710000000
1!
1%
1-
12
#317720000000
0!
0%
b110 *
0-
02
b110 6
#317730000000
1!
1%
1-
12
#317740000000
0!
0%
b111 *
0-
02
b111 6
#317750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#317760000000
0!
0%
b0 *
0-
02
b0 6
#317770000000
1!
1%
1-
12
#317780000000
0!
0%
b1 *
0-
02
b1 6
#317790000000
1!
1%
1-
12
#317800000000
0!
0%
b10 *
0-
02
b10 6
#317810000000
1!
1%
1-
12
#317820000000
0!
0%
b11 *
0-
02
b11 6
#317830000000
1!
1%
1-
12
15
#317840000000
0!
0%
b100 *
0-
02
b100 6
#317850000000
1!
1%
1-
12
#317860000000
0!
0%
b101 *
0-
02
b101 6
#317870000000
1!
1%
1-
12
#317880000000
0!
0%
b110 *
0-
02
b110 6
#317890000000
1!
1%
1-
12
#317900000000
0!
0%
b111 *
0-
02
b111 6
#317910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#317920000000
0!
0%
b0 *
0-
02
b0 6
#317930000000
1!
1%
1-
12
#317940000000
0!
0%
b1 *
0-
02
b1 6
#317950000000
1!
1%
1-
12
#317960000000
0!
0%
b10 *
0-
02
b10 6
#317970000000
1!
1%
1-
12
#317980000000
0!
0%
b11 *
0-
02
b11 6
#317990000000
1!
1%
1-
12
15
#318000000000
0!
0%
b100 *
0-
02
b100 6
#318010000000
1!
1%
1-
12
#318020000000
0!
0%
b101 *
0-
02
b101 6
#318030000000
1!
1%
1-
12
#318040000000
0!
0%
b110 *
0-
02
b110 6
#318050000000
1!
1%
1-
12
#318060000000
0!
0%
b111 *
0-
02
b111 6
#318070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#318080000000
0!
0%
b0 *
0-
02
b0 6
#318090000000
1!
1%
1-
12
#318100000000
0!
0%
b1 *
0-
02
b1 6
#318110000000
1!
1%
1-
12
#318120000000
0!
0%
b10 *
0-
02
b10 6
#318130000000
1!
1%
1-
12
#318140000000
0!
0%
b11 *
0-
02
b11 6
#318150000000
1!
1%
1-
12
15
#318160000000
0!
0%
b100 *
0-
02
b100 6
#318170000000
1!
1%
1-
12
#318180000000
0!
0%
b101 *
0-
02
b101 6
#318190000000
1!
1%
1-
12
#318200000000
0!
0%
b110 *
0-
02
b110 6
#318210000000
1!
1%
1-
12
#318220000000
0!
0%
b111 *
0-
02
b111 6
#318230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#318240000000
0!
0%
b0 *
0-
02
b0 6
#318250000000
1!
1%
1-
12
#318260000000
0!
0%
b1 *
0-
02
b1 6
#318270000000
1!
1%
1-
12
#318280000000
0!
0%
b10 *
0-
02
b10 6
#318290000000
1!
1%
1-
12
#318300000000
0!
0%
b11 *
0-
02
b11 6
#318310000000
1!
1%
1-
12
15
#318320000000
0!
0%
b100 *
0-
02
b100 6
#318330000000
1!
1%
1-
12
#318340000000
0!
0%
b101 *
0-
02
b101 6
#318350000000
1!
1%
1-
12
#318360000000
0!
0%
b110 *
0-
02
b110 6
#318370000000
1!
1%
1-
12
#318380000000
0!
0%
b111 *
0-
02
b111 6
#318390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#318400000000
0!
0%
b0 *
0-
02
b0 6
#318410000000
1!
1%
1-
12
#318420000000
0!
0%
b1 *
0-
02
b1 6
#318430000000
1!
1%
1-
12
#318440000000
0!
0%
b10 *
0-
02
b10 6
#318450000000
1!
1%
1-
12
#318460000000
0!
0%
b11 *
0-
02
b11 6
#318470000000
1!
1%
1-
12
15
#318480000000
0!
0%
b100 *
0-
02
b100 6
#318490000000
1!
1%
1-
12
#318500000000
0!
0%
b101 *
0-
02
b101 6
#318510000000
1!
1%
1-
12
#318520000000
0!
0%
b110 *
0-
02
b110 6
#318530000000
1!
1%
1-
12
#318540000000
0!
0%
b111 *
0-
02
b111 6
#318550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#318560000000
0!
0%
b0 *
0-
02
b0 6
#318570000000
1!
1%
1-
12
#318580000000
0!
0%
b1 *
0-
02
b1 6
#318590000000
1!
1%
1-
12
#318600000000
0!
0%
b10 *
0-
02
b10 6
#318610000000
1!
1%
1-
12
#318620000000
0!
0%
b11 *
0-
02
b11 6
#318630000000
1!
1%
1-
12
15
#318640000000
0!
0%
b100 *
0-
02
b100 6
#318650000000
1!
1%
1-
12
#318660000000
0!
0%
b101 *
0-
02
b101 6
#318670000000
1!
1%
1-
12
#318680000000
0!
0%
b110 *
0-
02
b110 6
#318690000000
1!
1%
1-
12
#318700000000
0!
0%
b111 *
0-
02
b111 6
#318710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#318720000000
0!
0%
b0 *
0-
02
b0 6
#318730000000
1!
1%
1-
12
#318740000000
0!
0%
b1 *
0-
02
b1 6
#318750000000
1!
1%
1-
12
#318760000000
0!
0%
b10 *
0-
02
b10 6
#318770000000
1!
1%
1-
12
#318780000000
0!
0%
b11 *
0-
02
b11 6
#318790000000
1!
1%
1-
12
15
#318800000000
0!
0%
b100 *
0-
02
b100 6
#318810000000
1!
1%
1-
12
#318820000000
0!
0%
b101 *
0-
02
b101 6
#318830000000
1!
1%
1-
12
#318840000000
0!
0%
b110 *
0-
02
b110 6
#318850000000
1!
1%
1-
12
#318860000000
0!
0%
b111 *
0-
02
b111 6
#318870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#318880000000
0!
0%
b0 *
0-
02
b0 6
#318890000000
1!
1%
1-
12
#318900000000
0!
0%
b1 *
0-
02
b1 6
#318910000000
1!
1%
1-
12
#318920000000
0!
0%
b10 *
0-
02
b10 6
#318930000000
1!
1%
1-
12
#318940000000
0!
0%
b11 *
0-
02
b11 6
#318950000000
1!
1%
1-
12
15
#318960000000
0!
0%
b100 *
0-
02
b100 6
#318970000000
1!
1%
1-
12
#318980000000
0!
0%
b101 *
0-
02
b101 6
#318990000000
1!
1%
1-
12
#319000000000
0!
0%
b110 *
0-
02
b110 6
#319010000000
1!
1%
1-
12
#319020000000
0!
0%
b111 *
0-
02
b111 6
#319030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#319040000000
0!
0%
b0 *
0-
02
b0 6
#319050000000
1!
1%
1-
12
#319060000000
0!
0%
b1 *
0-
02
b1 6
#319070000000
1!
1%
1-
12
#319080000000
0!
0%
b10 *
0-
02
b10 6
#319090000000
1!
1%
1-
12
#319100000000
0!
0%
b11 *
0-
02
b11 6
#319110000000
1!
1%
1-
12
15
#319120000000
0!
0%
b100 *
0-
02
b100 6
#319130000000
1!
1%
1-
12
#319140000000
0!
0%
b101 *
0-
02
b101 6
#319150000000
1!
1%
1-
12
#319160000000
0!
0%
b110 *
0-
02
b110 6
#319170000000
1!
1%
1-
12
#319180000000
0!
0%
b111 *
0-
02
b111 6
#319190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#319200000000
0!
0%
b0 *
0-
02
b0 6
#319210000000
1!
1%
1-
12
#319220000000
0!
0%
b1 *
0-
02
b1 6
#319230000000
1!
1%
1-
12
#319240000000
0!
0%
b10 *
0-
02
b10 6
#319250000000
1!
1%
1-
12
#319260000000
0!
0%
b11 *
0-
02
b11 6
#319270000000
1!
1%
1-
12
15
#319280000000
0!
0%
b100 *
0-
02
b100 6
#319290000000
1!
1%
1-
12
#319300000000
0!
0%
b101 *
0-
02
b101 6
#319310000000
1!
1%
1-
12
#319320000000
0!
0%
b110 *
0-
02
b110 6
#319330000000
1!
1%
1-
12
#319340000000
0!
0%
b111 *
0-
02
b111 6
#319350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#319360000000
0!
0%
b0 *
0-
02
b0 6
#319370000000
1!
1%
1-
12
#319380000000
0!
0%
b1 *
0-
02
b1 6
#319390000000
1!
1%
1-
12
#319400000000
0!
0%
b10 *
0-
02
b10 6
#319410000000
1!
1%
1-
12
#319420000000
0!
0%
b11 *
0-
02
b11 6
#319430000000
1!
1%
1-
12
15
#319440000000
0!
0%
b100 *
0-
02
b100 6
#319450000000
1!
1%
1-
12
#319460000000
0!
0%
b101 *
0-
02
b101 6
#319470000000
1!
1%
1-
12
#319480000000
0!
0%
b110 *
0-
02
b110 6
#319490000000
1!
1%
1-
12
#319500000000
0!
0%
b111 *
0-
02
b111 6
#319510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#319520000000
0!
0%
b0 *
0-
02
b0 6
#319530000000
1!
1%
1-
12
#319540000000
0!
0%
b1 *
0-
02
b1 6
#319550000000
1!
1%
1-
12
#319560000000
0!
0%
b10 *
0-
02
b10 6
#319570000000
1!
1%
1-
12
#319580000000
0!
0%
b11 *
0-
02
b11 6
#319590000000
1!
1%
1-
12
15
#319600000000
0!
0%
b100 *
0-
02
b100 6
#319610000000
1!
1%
1-
12
#319620000000
0!
0%
b101 *
0-
02
b101 6
#319630000000
1!
1%
1-
12
#319640000000
0!
0%
b110 *
0-
02
b110 6
#319650000000
1!
1%
1-
12
#319660000000
0!
0%
b111 *
0-
02
b111 6
#319670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#319680000000
0!
0%
b0 *
0-
02
b0 6
#319690000000
1!
1%
1-
12
#319700000000
0!
0%
b1 *
0-
02
b1 6
#319710000000
1!
1%
1-
12
#319720000000
0!
0%
b10 *
0-
02
b10 6
#319730000000
1!
1%
1-
12
#319740000000
0!
0%
b11 *
0-
02
b11 6
#319750000000
1!
1%
1-
12
15
#319760000000
0!
0%
b100 *
0-
02
b100 6
#319770000000
1!
1%
1-
12
#319780000000
0!
0%
b101 *
0-
02
b101 6
#319790000000
1!
1%
1-
12
#319800000000
0!
0%
b110 *
0-
02
b110 6
#319810000000
1!
1%
1-
12
#319820000000
0!
0%
b111 *
0-
02
b111 6
#319830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#319840000000
0!
0%
b0 *
0-
02
b0 6
#319850000000
1!
1%
1-
12
#319860000000
0!
0%
b1 *
0-
02
b1 6
#319870000000
1!
1%
1-
12
#319880000000
0!
0%
b10 *
0-
02
b10 6
#319890000000
1!
1%
1-
12
#319900000000
0!
0%
b11 *
0-
02
b11 6
#319910000000
1!
1%
1-
12
15
#319920000000
0!
0%
b100 *
0-
02
b100 6
#319930000000
1!
1%
1-
12
#319940000000
0!
0%
b101 *
0-
02
b101 6
#319950000000
1!
1%
1-
12
#319960000000
0!
0%
b110 *
0-
02
b110 6
#319970000000
1!
1%
1-
12
#319980000000
0!
0%
b111 *
0-
02
b111 6
#319990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#320000000000
0!
0%
b0 *
0-
02
b0 6
#320010000000
1!
1%
1-
12
#320020000000
0!
0%
b1 *
0-
02
b1 6
#320030000000
1!
1%
1-
12
#320040000000
0!
0%
b10 *
0-
02
b10 6
#320050000000
1!
1%
1-
12
#320060000000
0!
0%
b11 *
0-
02
b11 6
#320070000000
1!
1%
1-
12
15
#320080000000
0!
0%
b100 *
0-
02
b100 6
#320090000000
1!
1%
1-
12
#320100000000
0!
0%
b101 *
0-
02
b101 6
#320110000000
1!
1%
1-
12
#320120000000
0!
0%
b110 *
0-
02
b110 6
#320130000000
1!
1%
1-
12
#320140000000
0!
0%
b111 *
0-
02
b111 6
#320150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#320160000000
0!
0%
b0 *
0-
02
b0 6
#320170000000
1!
1%
1-
12
#320180000000
0!
0%
b1 *
0-
02
b1 6
#320190000000
1!
1%
1-
12
#320200000000
0!
0%
b10 *
0-
02
b10 6
#320210000000
1!
1%
1-
12
#320220000000
0!
0%
b11 *
0-
02
b11 6
#320230000000
1!
1%
1-
12
15
#320240000000
0!
0%
b100 *
0-
02
b100 6
#320250000000
1!
1%
1-
12
#320260000000
0!
0%
b101 *
0-
02
b101 6
#320270000000
1!
1%
1-
12
#320280000000
0!
0%
b110 *
0-
02
b110 6
#320290000000
1!
1%
1-
12
#320300000000
0!
0%
b111 *
0-
02
b111 6
#320310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#320320000000
0!
0%
b0 *
0-
02
b0 6
#320330000000
1!
1%
1-
12
#320340000000
0!
0%
b1 *
0-
02
b1 6
#320350000000
1!
1%
1-
12
#320360000000
0!
0%
b10 *
0-
02
b10 6
#320370000000
1!
1%
1-
12
#320380000000
0!
0%
b11 *
0-
02
b11 6
#320390000000
1!
1%
1-
12
15
#320400000000
0!
0%
b100 *
0-
02
b100 6
#320410000000
1!
1%
1-
12
#320420000000
0!
0%
b101 *
0-
02
b101 6
#320430000000
1!
1%
1-
12
#320440000000
0!
0%
b110 *
0-
02
b110 6
#320450000000
1!
1%
1-
12
#320460000000
0!
0%
b111 *
0-
02
b111 6
#320470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#320480000000
0!
0%
b0 *
0-
02
b0 6
#320490000000
1!
1%
1-
12
#320500000000
0!
0%
b1 *
0-
02
b1 6
#320510000000
1!
1%
1-
12
#320520000000
0!
0%
b10 *
0-
02
b10 6
#320530000000
1!
1%
1-
12
#320540000000
0!
0%
b11 *
0-
02
b11 6
#320550000000
1!
1%
1-
12
15
#320560000000
0!
0%
b100 *
0-
02
b100 6
#320570000000
1!
1%
1-
12
#320580000000
0!
0%
b101 *
0-
02
b101 6
#320590000000
1!
1%
1-
12
#320600000000
0!
0%
b110 *
0-
02
b110 6
#320610000000
1!
1%
1-
12
#320620000000
0!
0%
b111 *
0-
02
b111 6
#320630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#320640000000
0!
0%
b0 *
0-
02
b0 6
#320650000000
1!
1%
1-
12
#320660000000
0!
0%
b1 *
0-
02
b1 6
#320670000000
1!
1%
1-
12
#320680000000
0!
0%
b10 *
0-
02
b10 6
#320690000000
1!
1%
1-
12
#320700000000
0!
0%
b11 *
0-
02
b11 6
#320710000000
1!
1%
1-
12
15
#320720000000
0!
0%
b100 *
0-
02
b100 6
#320730000000
1!
1%
1-
12
#320740000000
0!
0%
b101 *
0-
02
b101 6
#320750000000
1!
1%
1-
12
#320760000000
0!
0%
b110 *
0-
02
b110 6
#320770000000
1!
1%
1-
12
#320780000000
0!
0%
b111 *
0-
02
b111 6
#320790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#320800000000
0!
0%
b0 *
0-
02
b0 6
#320810000000
1!
1%
1-
12
#320820000000
0!
0%
b1 *
0-
02
b1 6
#320830000000
1!
1%
1-
12
#320840000000
0!
0%
b10 *
0-
02
b10 6
#320850000000
1!
1%
1-
12
#320860000000
0!
0%
b11 *
0-
02
b11 6
#320870000000
1!
1%
1-
12
15
#320880000000
0!
0%
b100 *
0-
02
b100 6
#320890000000
1!
1%
1-
12
#320900000000
0!
0%
b101 *
0-
02
b101 6
#320910000000
1!
1%
1-
12
#320920000000
0!
0%
b110 *
0-
02
b110 6
#320930000000
1!
1%
1-
12
#320940000000
0!
0%
b111 *
0-
02
b111 6
#320950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#320960000000
0!
0%
b0 *
0-
02
b0 6
#320970000000
1!
1%
1-
12
#320980000000
0!
0%
b1 *
0-
02
b1 6
#320990000000
1!
1%
1-
12
#321000000000
0!
0%
b10 *
0-
02
b10 6
#321010000000
1!
1%
1-
12
#321020000000
0!
0%
b11 *
0-
02
b11 6
#321030000000
1!
1%
1-
12
15
#321040000000
0!
0%
b100 *
0-
02
b100 6
#321050000000
1!
1%
1-
12
#321060000000
0!
0%
b101 *
0-
02
b101 6
#321070000000
1!
1%
1-
12
#321080000000
0!
0%
b110 *
0-
02
b110 6
#321090000000
1!
1%
1-
12
#321100000000
0!
0%
b111 *
0-
02
b111 6
#321110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#321120000000
0!
0%
b0 *
0-
02
b0 6
#321130000000
1!
1%
1-
12
#321140000000
0!
0%
b1 *
0-
02
b1 6
#321150000000
1!
1%
1-
12
#321160000000
0!
0%
b10 *
0-
02
b10 6
#321170000000
1!
1%
1-
12
#321180000000
0!
0%
b11 *
0-
02
b11 6
#321190000000
1!
1%
1-
12
15
#321200000000
0!
0%
b100 *
0-
02
b100 6
#321210000000
1!
1%
1-
12
#321220000000
0!
0%
b101 *
0-
02
b101 6
#321230000000
1!
1%
1-
12
#321240000000
0!
0%
b110 *
0-
02
b110 6
#321250000000
1!
1%
1-
12
#321260000000
0!
0%
b111 *
0-
02
b111 6
#321270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#321280000000
0!
0%
b0 *
0-
02
b0 6
#321290000000
1!
1%
1-
12
#321300000000
0!
0%
b1 *
0-
02
b1 6
#321310000000
1!
1%
1-
12
#321320000000
0!
0%
b10 *
0-
02
b10 6
#321330000000
1!
1%
1-
12
#321340000000
0!
0%
b11 *
0-
02
b11 6
#321350000000
1!
1%
1-
12
15
#321360000000
0!
0%
b100 *
0-
02
b100 6
#321370000000
1!
1%
1-
12
#321380000000
0!
0%
b101 *
0-
02
b101 6
#321390000000
1!
1%
1-
12
#321400000000
0!
0%
b110 *
0-
02
b110 6
#321410000000
1!
1%
1-
12
#321420000000
0!
0%
b111 *
0-
02
b111 6
#321430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#321440000000
0!
0%
b0 *
0-
02
b0 6
#321450000000
1!
1%
1-
12
#321460000000
0!
0%
b1 *
0-
02
b1 6
#321470000000
1!
1%
1-
12
#321480000000
0!
0%
b10 *
0-
02
b10 6
#321490000000
1!
1%
1-
12
#321500000000
0!
0%
b11 *
0-
02
b11 6
#321510000000
1!
1%
1-
12
15
#321520000000
0!
0%
b100 *
0-
02
b100 6
#321530000000
1!
1%
1-
12
#321540000000
0!
0%
b101 *
0-
02
b101 6
#321550000000
1!
1%
1-
12
#321560000000
0!
0%
b110 *
0-
02
b110 6
#321570000000
1!
1%
1-
12
#321580000000
0!
0%
b111 *
0-
02
b111 6
#321590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#321600000000
0!
0%
b0 *
0-
02
b0 6
#321610000000
1!
1%
1-
12
#321620000000
0!
0%
b1 *
0-
02
b1 6
#321630000000
1!
1%
1-
12
#321640000000
0!
0%
b10 *
0-
02
b10 6
#321650000000
1!
1%
1-
12
#321660000000
0!
0%
b11 *
0-
02
b11 6
#321670000000
1!
1%
1-
12
15
#321680000000
0!
0%
b100 *
0-
02
b100 6
#321690000000
1!
1%
1-
12
#321700000000
0!
0%
b101 *
0-
02
b101 6
#321710000000
1!
1%
1-
12
#321720000000
0!
0%
b110 *
0-
02
b110 6
#321730000000
1!
1%
1-
12
#321740000000
0!
0%
b111 *
0-
02
b111 6
#321750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#321760000000
0!
0%
b0 *
0-
02
b0 6
#321770000000
1!
1%
1-
12
#321780000000
0!
0%
b1 *
0-
02
b1 6
#321790000000
1!
1%
1-
12
#321800000000
0!
0%
b10 *
0-
02
b10 6
#321810000000
1!
1%
1-
12
#321820000000
0!
0%
b11 *
0-
02
b11 6
#321830000000
1!
1%
1-
12
15
#321840000000
0!
0%
b100 *
0-
02
b100 6
#321850000000
1!
1%
1-
12
#321860000000
0!
0%
b101 *
0-
02
b101 6
#321870000000
1!
1%
1-
12
#321880000000
0!
0%
b110 *
0-
02
b110 6
#321890000000
1!
1%
1-
12
#321900000000
0!
0%
b111 *
0-
02
b111 6
#321910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#321920000000
0!
0%
b0 *
0-
02
b0 6
#321930000000
1!
1%
1-
12
#321940000000
0!
0%
b1 *
0-
02
b1 6
#321950000000
1!
1%
1-
12
#321960000000
0!
0%
b10 *
0-
02
b10 6
#321970000000
1!
1%
1-
12
#321980000000
0!
0%
b11 *
0-
02
b11 6
#321990000000
1!
1%
1-
12
15
#322000000000
0!
0%
b100 *
0-
02
b100 6
#322010000000
1!
1%
1-
12
#322020000000
0!
0%
b101 *
0-
02
b101 6
#322030000000
1!
1%
1-
12
#322040000000
0!
0%
b110 *
0-
02
b110 6
#322050000000
1!
1%
1-
12
#322060000000
0!
0%
b111 *
0-
02
b111 6
#322070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#322080000000
0!
0%
b0 *
0-
02
b0 6
#322090000000
1!
1%
1-
12
#322100000000
0!
0%
b1 *
0-
02
b1 6
#322110000000
1!
1%
1-
12
#322120000000
0!
0%
b10 *
0-
02
b10 6
#322130000000
1!
1%
1-
12
#322140000000
0!
0%
b11 *
0-
02
b11 6
#322150000000
1!
1%
1-
12
15
#322160000000
0!
0%
b100 *
0-
02
b100 6
#322170000000
1!
1%
1-
12
#322180000000
0!
0%
b101 *
0-
02
b101 6
#322190000000
1!
1%
1-
12
#322200000000
0!
0%
b110 *
0-
02
b110 6
#322210000000
1!
1%
1-
12
#322220000000
0!
0%
b111 *
0-
02
b111 6
#322230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#322240000000
0!
0%
b0 *
0-
02
b0 6
#322250000000
1!
1%
1-
12
#322260000000
0!
0%
b1 *
0-
02
b1 6
#322270000000
1!
1%
1-
12
#322280000000
0!
0%
b10 *
0-
02
b10 6
#322290000000
1!
1%
1-
12
#322300000000
0!
0%
b11 *
0-
02
b11 6
#322310000000
1!
1%
1-
12
15
#322320000000
0!
0%
b100 *
0-
02
b100 6
#322330000000
1!
1%
1-
12
#322340000000
0!
0%
b101 *
0-
02
b101 6
#322350000000
1!
1%
1-
12
#322360000000
0!
0%
b110 *
0-
02
b110 6
#322370000000
1!
1%
1-
12
#322380000000
0!
0%
b111 *
0-
02
b111 6
#322390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#322400000000
0!
0%
b0 *
0-
02
b0 6
#322410000000
1!
1%
1-
12
#322420000000
0!
0%
b1 *
0-
02
b1 6
#322430000000
1!
1%
1-
12
#322440000000
0!
0%
b10 *
0-
02
b10 6
#322450000000
1!
1%
1-
12
#322460000000
0!
0%
b11 *
0-
02
b11 6
#322470000000
1!
1%
1-
12
15
#322480000000
0!
0%
b100 *
0-
02
b100 6
#322490000000
1!
1%
1-
12
#322500000000
0!
0%
b101 *
0-
02
b101 6
#322510000000
1!
1%
1-
12
#322520000000
0!
0%
b110 *
0-
02
b110 6
#322530000000
1!
1%
1-
12
#322540000000
0!
0%
b111 *
0-
02
b111 6
#322550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#322560000000
0!
0%
b0 *
0-
02
b0 6
#322570000000
1!
1%
1-
12
#322580000000
0!
0%
b1 *
0-
02
b1 6
#322590000000
1!
1%
1-
12
#322600000000
0!
0%
b10 *
0-
02
b10 6
#322610000000
1!
1%
1-
12
#322620000000
0!
0%
b11 *
0-
02
b11 6
#322630000000
1!
1%
1-
12
15
#322640000000
0!
0%
b100 *
0-
02
b100 6
#322650000000
1!
1%
1-
12
#322660000000
0!
0%
b101 *
0-
02
b101 6
#322670000000
1!
1%
1-
12
#322680000000
0!
0%
b110 *
0-
02
b110 6
#322690000000
1!
1%
1-
12
#322700000000
0!
0%
b111 *
0-
02
b111 6
#322710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#322720000000
0!
0%
b0 *
0-
02
b0 6
#322730000000
1!
1%
1-
12
#322740000000
0!
0%
b1 *
0-
02
b1 6
#322750000000
1!
1%
1-
12
#322760000000
0!
0%
b10 *
0-
02
b10 6
#322770000000
1!
1%
1-
12
#322780000000
0!
0%
b11 *
0-
02
b11 6
#322790000000
1!
1%
1-
12
15
#322800000000
0!
0%
b100 *
0-
02
b100 6
#322810000000
1!
1%
1-
12
#322820000000
0!
0%
b101 *
0-
02
b101 6
#322830000000
1!
1%
1-
12
#322840000000
0!
0%
b110 *
0-
02
b110 6
#322850000000
1!
1%
1-
12
#322860000000
0!
0%
b111 *
0-
02
b111 6
#322870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#322880000000
0!
0%
b0 *
0-
02
b0 6
#322890000000
1!
1%
1-
12
#322900000000
0!
0%
b1 *
0-
02
b1 6
#322910000000
1!
1%
1-
12
#322920000000
0!
0%
b10 *
0-
02
b10 6
#322930000000
1!
1%
1-
12
#322940000000
0!
0%
b11 *
0-
02
b11 6
#322950000000
1!
1%
1-
12
15
#322960000000
0!
0%
b100 *
0-
02
b100 6
#322970000000
1!
1%
1-
12
#322980000000
0!
0%
b101 *
0-
02
b101 6
#322990000000
1!
1%
1-
12
#323000000000
0!
0%
b110 *
0-
02
b110 6
#323010000000
1!
1%
1-
12
#323020000000
0!
0%
b111 *
0-
02
b111 6
#323030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#323040000000
0!
0%
b0 *
0-
02
b0 6
#323050000000
1!
1%
1-
12
#323060000000
0!
0%
b1 *
0-
02
b1 6
#323070000000
1!
1%
1-
12
#323080000000
0!
0%
b10 *
0-
02
b10 6
#323090000000
1!
1%
1-
12
#323100000000
0!
0%
b11 *
0-
02
b11 6
#323110000000
1!
1%
1-
12
15
#323120000000
0!
0%
b100 *
0-
02
b100 6
#323130000000
1!
1%
1-
12
#323140000000
0!
0%
b101 *
0-
02
b101 6
#323150000000
1!
1%
1-
12
#323160000000
0!
0%
b110 *
0-
02
b110 6
#323170000000
1!
1%
1-
12
#323180000000
0!
0%
b111 *
0-
02
b111 6
#323190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#323200000000
0!
0%
b0 *
0-
02
b0 6
#323210000000
1!
1%
1-
12
#323220000000
0!
0%
b1 *
0-
02
b1 6
#323230000000
1!
1%
1-
12
#323240000000
0!
0%
b10 *
0-
02
b10 6
#323250000000
1!
1%
1-
12
#323260000000
0!
0%
b11 *
0-
02
b11 6
#323270000000
1!
1%
1-
12
15
#323280000000
0!
0%
b100 *
0-
02
b100 6
#323290000000
1!
1%
1-
12
#323300000000
0!
0%
b101 *
0-
02
b101 6
#323310000000
1!
1%
1-
12
#323320000000
0!
0%
b110 *
0-
02
b110 6
#323330000000
1!
1%
1-
12
#323340000000
0!
0%
b111 *
0-
02
b111 6
#323350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#323360000000
0!
0%
b0 *
0-
02
b0 6
#323370000000
1!
1%
1-
12
#323380000000
0!
0%
b1 *
0-
02
b1 6
#323390000000
1!
1%
1-
12
#323400000000
0!
0%
b10 *
0-
02
b10 6
#323410000000
1!
1%
1-
12
#323420000000
0!
0%
b11 *
0-
02
b11 6
#323430000000
1!
1%
1-
12
15
#323440000000
0!
0%
b100 *
0-
02
b100 6
#323450000000
1!
1%
1-
12
#323460000000
0!
0%
b101 *
0-
02
b101 6
#323470000000
1!
1%
1-
12
#323480000000
0!
0%
b110 *
0-
02
b110 6
#323490000000
1!
1%
1-
12
#323500000000
0!
0%
b111 *
0-
02
b111 6
#323510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#323520000000
0!
0%
b0 *
0-
02
b0 6
#323530000000
1!
1%
1-
12
#323540000000
0!
0%
b1 *
0-
02
b1 6
#323550000000
1!
1%
1-
12
#323560000000
0!
0%
b10 *
0-
02
b10 6
#323570000000
1!
1%
1-
12
#323580000000
0!
0%
b11 *
0-
02
b11 6
#323590000000
1!
1%
1-
12
15
#323600000000
0!
0%
b100 *
0-
02
b100 6
#323610000000
1!
1%
1-
12
#323620000000
0!
0%
b101 *
0-
02
b101 6
#323630000000
1!
1%
1-
12
#323640000000
0!
0%
b110 *
0-
02
b110 6
#323650000000
1!
1%
1-
12
#323660000000
0!
0%
b111 *
0-
02
b111 6
#323670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#323680000000
0!
0%
b0 *
0-
02
b0 6
#323690000000
1!
1%
1-
12
#323700000000
0!
0%
b1 *
0-
02
b1 6
#323710000000
1!
1%
1-
12
#323720000000
0!
0%
b10 *
0-
02
b10 6
#323730000000
1!
1%
1-
12
#323740000000
0!
0%
b11 *
0-
02
b11 6
#323750000000
1!
1%
1-
12
15
#323760000000
0!
0%
b100 *
0-
02
b100 6
#323770000000
1!
1%
1-
12
#323780000000
0!
0%
b101 *
0-
02
b101 6
#323790000000
1!
1%
1-
12
#323800000000
0!
0%
b110 *
0-
02
b110 6
#323810000000
1!
1%
1-
12
#323820000000
0!
0%
b111 *
0-
02
b111 6
#323830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#323840000000
0!
0%
b0 *
0-
02
b0 6
#323850000000
1!
1%
1-
12
#323860000000
0!
0%
b1 *
0-
02
b1 6
#323870000000
1!
1%
1-
12
#323880000000
0!
0%
b10 *
0-
02
b10 6
#323890000000
1!
1%
1-
12
#323900000000
0!
0%
b11 *
0-
02
b11 6
#323910000000
1!
1%
1-
12
15
#323920000000
0!
0%
b100 *
0-
02
b100 6
#323930000000
1!
1%
1-
12
#323940000000
0!
0%
b101 *
0-
02
b101 6
#323950000000
1!
1%
1-
12
#323960000000
0!
0%
b110 *
0-
02
b110 6
#323970000000
1!
1%
1-
12
#323980000000
0!
0%
b111 *
0-
02
b111 6
#323990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#324000000000
0!
0%
b0 *
0-
02
b0 6
#324010000000
1!
1%
1-
12
#324020000000
0!
0%
b1 *
0-
02
b1 6
#324030000000
1!
1%
1-
12
#324040000000
0!
0%
b10 *
0-
02
b10 6
#324050000000
1!
1%
1-
12
#324060000000
0!
0%
b11 *
0-
02
b11 6
#324070000000
1!
1%
1-
12
15
#324080000000
0!
0%
b100 *
0-
02
b100 6
#324090000000
1!
1%
1-
12
#324100000000
0!
0%
b101 *
0-
02
b101 6
#324110000000
1!
1%
1-
12
#324120000000
0!
0%
b110 *
0-
02
b110 6
#324130000000
1!
1%
1-
12
#324140000000
0!
0%
b111 *
0-
02
b111 6
#324150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#324160000000
0!
0%
b0 *
0-
02
b0 6
#324170000000
1!
1%
1-
12
#324180000000
0!
0%
b1 *
0-
02
b1 6
#324190000000
1!
1%
1-
12
#324200000000
0!
0%
b10 *
0-
02
b10 6
#324210000000
1!
1%
1-
12
#324220000000
0!
0%
b11 *
0-
02
b11 6
#324230000000
1!
1%
1-
12
15
#324240000000
0!
0%
b100 *
0-
02
b100 6
#324250000000
1!
1%
1-
12
#324260000000
0!
0%
b101 *
0-
02
b101 6
#324270000000
1!
1%
1-
12
#324280000000
0!
0%
b110 *
0-
02
b110 6
#324290000000
1!
1%
1-
12
#324300000000
0!
0%
b111 *
0-
02
b111 6
#324310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#324320000000
0!
0%
b0 *
0-
02
b0 6
#324330000000
1!
1%
1-
12
#324340000000
0!
0%
b1 *
0-
02
b1 6
#324350000000
1!
1%
1-
12
#324360000000
0!
0%
b10 *
0-
02
b10 6
#324370000000
1!
1%
1-
12
#324380000000
0!
0%
b11 *
0-
02
b11 6
#324390000000
1!
1%
1-
12
15
#324400000000
0!
0%
b100 *
0-
02
b100 6
#324410000000
1!
1%
1-
12
#324420000000
0!
0%
b101 *
0-
02
b101 6
#324430000000
1!
1%
1-
12
#324440000000
0!
0%
b110 *
0-
02
b110 6
#324450000000
1!
1%
1-
12
#324460000000
0!
0%
b111 *
0-
02
b111 6
#324470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#324480000000
0!
0%
b0 *
0-
02
b0 6
#324490000000
1!
1%
1-
12
#324500000000
0!
0%
b1 *
0-
02
b1 6
#324510000000
1!
1%
1-
12
#324520000000
0!
0%
b10 *
0-
02
b10 6
#324530000000
1!
1%
1-
12
#324540000000
0!
0%
b11 *
0-
02
b11 6
#324550000000
1!
1%
1-
12
15
#324560000000
0!
0%
b100 *
0-
02
b100 6
#324570000000
1!
1%
1-
12
#324580000000
0!
0%
b101 *
0-
02
b101 6
#324590000000
1!
1%
1-
12
#324600000000
0!
0%
b110 *
0-
02
b110 6
#324610000000
1!
1%
1-
12
#324620000000
0!
0%
b111 *
0-
02
b111 6
#324630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#324640000000
0!
0%
b0 *
0-
02
b0 6
#324650000000
1!
1%
1-
12
#324660000000
0!
0%
b1 *
0-
02
b1 6
#324670000000
1!
1%
1-
12
#324680000000
0!
0%
b10 *
0-
02
b10 6
#324690000000
1!
1%
1-
12
#324700000000
0!
0%
b11 *
0-
02
b11 6
#324710000000
1!
1%
1-
12
15
#324720000000
0!
0%
b100 *
0-
02
b100 6
#324730000000
1!
1%
1-
12
#324740000000
0!
0%
b101 *
0-
02
b101 6
#324750000000
1!
1%
1-
12
#324760000000
0!
0%
b110 *
0-
02
b110 6
#324770000000
1!
1%
1-
12
#324780000000
0!
0%
b111 *
0-
02
b111 6
#324790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#324800000000
0!
0%
b0 *
0-
02
b0 6
#324810000000
1!
1%
1-
12
#324820000000
0!
0%
b1 *
0-
02
b1 6
#324830000000
1!
1%
1-
12
#324840000000
0!
0%
b10 *
0-
02
b10 6
#324850000000
1!
1%
1-
12
#324860000000
0!
0%
b11 *
0-
02
b11 6
#324870000000
1!
1%
1-
12
15
#324880000000
0!
0%
b100 *
0-
02
b100 6
#324890000000
1!
1%
1-
12
#324900000000
0!
0%
b101 *
0-
02
b101 6
#324910000000
1!
1%
1-
12
#324920000000
0!
0%
b110 *
0-
02
b110 6
#324930000000
1!
1%
1-
12
#324940000000
0!
0%
b111 *
0-
02
b111 6
#324950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#324960000000
0!
0%
b0 *
0-
02
b0 6
#324970000000
1!
1%
1-
12
#324980000000
0!
0%
b1 *
0-
02
b1 6
#324990000000
1!
1%
1-
12
#325000000000
0!
0%
b10 *
0-
02
b10 6
#325010000000
1!
1%
1-
12
#325020000000
0!
0%
b11 *
0-
02
b11 6
#325030000000
1!
1%
1-
12
15
#325040000000
0!
0%
b100 *
0-
02
b100 6
#325050000000
1!
1%
1-
12
#325060000000
0!
0%
b101 *
0-
02
b101 6
#325070000000
1!
1%
1-
12
#325080000000
0!
0%
b110 *
0-
02
b110 6
#325090000000
1!
1%
1-
12
#325100000000
0!
0%
b111 *
0-
02
b111 6
#325110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#325120000000
0!
0%
b0 *
0-
02
b0 6
#325130000000
1!
1%
1-
12
#325140000000
0!
0%
b1 *
0-
02
b1 6
#325150000000
1!
1%
1-
12
#325160000000
0!
0%
b10 *
0-
02
b10 6
#325170000000
1!
1%
1-
12
#325180000000
0!
0%
b11 *
0-
02
b11 6
#325190000000
1!
1%
1-
12
15
#325200000000
0!
0%
b100 *
0-
02
b100 6
#325210000000
1!
1%
1-
12
#325220000000
0!
0%
b101 *
0-
02
b101 6
#325230000000
1!
1%
1-
12
#325240000000
0!
0%
b110 *
0-
02
b110 6
#325250000000
1!
1%
1-
12
#325260000000
0!
0%
b111 *
0-
02
b111 6
#325270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#325280000000
0!
0%
b0 *
0-
02
b0 6
#325290000000
1!
1%
1-
12
#325300000000
0!
0%
b1 *
0-
02
b1 6
#325310000000
1!
1%
1-
12
#325320000000
0!
0%
b10 *
0-
02
b10 6
#325330000000
1!
1%
1-
12
#325340000000
0!
0%
b11 *
0-
02
b11 6
#325350000000
1!
1%
1-
12
15
#325360000000
0!
0%
b100 *
0-
02
b100 6
#325370000000
1!
1%
1-
12
#325380000000
0!
0%
b101 *
0-
02
b101 6
#325390000000
1!
1%
1-
12
#325400000000
0!
0%
b110 *
0-
02
b110 6
#325410000000
1!
1%
1-
12
#325420000000
0!
0%
b111 *
0-
02
b111 6
#325430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#325440000000
0!
0%
b0 *
0-
02
b0 6
#325450000000
1!
1%
1-
12
#325460000000
0!
0%
b1 *
0-
02
b1 6
#325470000000
1!
1%
1-
12
#325480000000
0!
0%
b10 *
0-
02
b10 6
#325490000000
1!
1%
1-
12
#325500000000
0!
0%
b11 *
0-
02
b11 6
#325510000000
1!
1%
1-
12
15
#325520000000
0!
0%
b100 *
0-
02
b100 6
#325530000000
1!
1%
1-
12
#325540000000
0!
0%
b101 *
0-
02
b101 6
#325550000000
1!
1%
1-
12
#325560000000
0!
0%
b110 *
0-
02
b110 6
#325570000000
1!
1%
1-
12
#325580000000
0!
0%
b111 *
0-
02
b111 6
#325590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#325600000000
0!
0%
b0 *
0-
02
b0 6
#325610000000
1!
1%
1-
12
#325620000000
0!
0%
b1 *
0-
02
b1 6
#325630000000
1!
1%
1-
12
#325640000000
0!
0%
b10 *
0-
02
b10 6
#325650000000
1!
1%
1-
12
#325660000000
0!
0%
b11 *
0-
02
b11 6
#325670000000
1!
1%
1-
12
15
#325680000000
0!
0%
b100 *
0-
02
b100 6
#325690000000
1!
1%
1-
12
#325700000000
0!
0%
b101 *
0-
02
b101 6
#325710000000
1!
1%
1-
12
#325720000000
0!
0%
b110 *
0-
02
b110 6
#325730000000
1!
1%
1-
12
#325740000000
0!
0%
b111 *
0-
02
b111 6
#325750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#325760000000
0!
0%
b0 *
0-
02
b0 6
#325770000000
1!
1%
1-
12
#325780000000
0!
0%
b1 *
0-
02
b1 6
#325790000000
1!
1%
1-
12
#325800000000
0!
0%
b10 *
0-
02
b10 6
#325810000000
1!
1%
1-
12
#325820000000
0!
0%
b11 *
0-
02
b11 6
#325830000000
1!
1%
1-
12
15
#325840000000
0!
0%
b100 *
0-
02
b100 6
#325850000000
1!
1%
1-
12
#325860000000
0!
0%
b101 *
0-
02
b101 6
#325870000000
1!
1%
1-
12
#325880000000
0!
0%
b110 *
0-
02
b110 6
#325890000000
1!
1%
1-
12
#325900000000
0!
0%
b111 *
0-
02
b111 6
#325910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#325920000000
0!
0%
b0 *
0-
02
b0 6
#325930000000
1!
1%
1-
12
#325940000000
0!
0%
b1 *
0-
02
b1 6
#325950000000
1!
1%
1-
12
#325960000000
0!
0%
b10 *
0-
02
b10 6
#325970000000
1!
1%
1-
12
#325980000000
0!
0%
b11 *
0-
02
b11 6
#325990000000
1!
1%
1-
12
15
#326000000000
0!
0%
b100 *
0-
02
b100 6
#326010000000
1!
1%
1-
12
#326020000000
0!
0%
b101 *
0-
02
b101 6
#326030000000
1!
1%
1-
12
#326040000000
0!
0%
b110 *
0-
02
b110 6
#326050000000
1!
1%
1-
12
#326060000000
0!
0%
b111 *
0-
02
b111 6
#326070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#326080000000
0!
0%
b0 *
0-
02
b0 6
#326090000000
1!
1%
1-
12
#326100000000
0!
0%
b1 *
0-
02
b1 6
#326110000000
1!
1%
1-
12
#326120000000
0!
0%
b10 *
0-
02
b10 6
#326130000000
1!
1%
1-
12
#326140000000
0!
0%
b11 *
0-
02
b11 6
#326150000000
1!
1%
1-
12
15
#326160000000
0!
0%
b100 *
0-
02
b100 6
#326170000000
1!
1%
1-
12
#326180000000
0!
0%
b101 *
0-
02
b101 6
#326190000000
1!
1%
1-
12
#326200000000
0!
0%
b110 *
0-
02
b110 6
#326210000000
1!
1%
1-
12
#326220000000
0!
0%
b111 *
0-
02
b111 6
#326230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#326240000000
0!
0%
b0 *
0-
02
b0 6
#326250000000
1!
1%
1-
12
#326260000000
0!
0%
b1 *
0-
02
b1 6
#326270000000
1!
1%
1-
12
#326280000000
0!
0%
b10 *
0-
02
b10 6
#326290000000
1!
1%
1-
12
#326300000000
0!
0%
b11 *
0-
02
b11 6
#326310000000
1!
1%
1-
12
15
#326320000000
0!
0%
b100 *
0-
02
b100 6
#326330000000
1!
1%
1-
12
#326340000000
0!
0%
b101 *
0-
02
b101 6
#326350000000
1!
1%
1-
12
#326360000000
0!
0%
b110 *
0-
02
b110 6
#326370000000
1!
1%
1-
12
#326380000000
0!
0%
b111 *
0-
02
b111 6
#326390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#326400000000
0!
0%
b0 *
0-
02
b0 6
#326410000000
1!
1%
1-
12
#326420000000
0!
0%
b1 *
0-
02
b1 6
#326430000000
1!
1%
1-
12
#326440000000
0!
0%
b10 *
0-
02
b10 6
#326450000000
1!
1%
1-
12
#326460000000
0!
0%
b11 *
0-
02
b11 6
#326470000000
1!
1%
1-
12
15
#326480000000
0!
0%
b100 *
0-
02
b100 6
#326490000000
1!
1%
1-
12
#326500000000
0!
0%
b101 *
0-
02
b101 6
#326510000000
1!
1%
1-
12
#326520000000
0!
0%
b110 *
0-
02
b110 6
#326530000000
1!
1%
1-
12
#326540000000
0!
0%
b111 *
0-
02
b111 6
#326550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#326560000000
0!
0%
b0 *
0-
02
b0 6
#326570000000
1!
1%
1-
12
#326580000000
0!
0%
b1 *
0-
02
b1 6
#326590000000
1!
1%
1-
12
#326600000000
0!
0%
b10 *
0-
02
b10 6
#326610000000
1!
1%
1-
12
#326620000000
0!
0%
b11 *
0-
02
b11 6
#326630000000
1!
1%
1-
12
15
#326640000000
0!
0%
b100 *
0-
02
b100 6
#326650000000
1!
1%
1-
12
#326660000000
0!
0%
b101 *
0-
02
b101 6
#326670000000
1!
1%
1-
12
#326680000000
0!
0%
b110 *
0-
02
b110 6
#326690000000
1!
1%
1-
12
#326700000000
0!
0%
b111 *
0-
02
b111 6
#326710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#326720000000
0!
0%
b0 *
0-
02
b0 6
#326730000000
1!
1%
1-
12
#326740000000
0!
0%
b1 *
0-
02
b1 6
#326750000000
1!
1%
1-
12
#326760000000
0!
0%
b10 *
0-
02
b10 6
#326770000000
1!
1%
1-
12
#326780000000
0!
0%
b11 *
0-
02
b11 6
#326790000000
1!
1%
1-
12
15
#326800000000
0!
0%
b100 *
0-
02
b100 6
#326810000000
1!
1%
1-
12
#326820000000
0!
0%
b101 *
0-
02
b101 6
#326830000000
1!
1%
1-
12
#326840000000
0!
0%
b110 *
0-
02
b110 6
#326850000000
1!
1%
1-
12
#326860000000
0!
0%
b111 *
0-
02
b111 6
#326870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#326880000000
0!
0%
b0 *
0-
02
b0 6
#326890000000
1!
1%
1-
12
#326900000000
0!
0%
b1 *
0-
02
b1 6
#326910000000
1!
1%
1-
12
#326920000000
0!
0%
b10 *
0-
02
b10 6
#326930000000
1!
1%
1-
12
#326940000000
0!
0%
b11 *
0-
02
b11 6
#326950000000
1!
1%
1-
12
15
#326960000000
0!
0%
b100 *
0-
02
b100 6
#326970000000
1!
1%
1-
12
#326980000000
0!
0%
b101 *
0-
02
b101 6
#326990000000
1!
1%
1-
12
#327000000000
0!
0%
b110 *
0-
02
b110 6
#327010000000
1!
1%
1-
12
#327020000000
0!
0%
b111 *
0-
02
b111 6
#327030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#327040000000
0!
0%
b0 *
0-
02
b0 6
#327050000000
1!
1%
1-
12
#327060000000
0!
0%
b1 *
0-
02
b1 6
#327070000000
1!
1%
1-
12
#327080000000
0!
0%
b10 *
0-
02
b10 6
#327090000000
1!
1%
1-
12
#327100000000
0!
0%
b11 *
0-
02
b11 6
#327110000000
1!
1%
1-
12
15
#327120000000
0!
0%
b100 *
0-
02
b100 6
#327130000000
1!
1%
1-
12
#327140000000
0!
0%
b101 *
0-
02
b101 6
#327150000000
1!
1%
1-
12
#327160000000
0!
0%
b110 *
0-
02
b110 6
#327170000000
1!
1%
1-
12
#327180000000
0!
0%
b111 *
0-
02
b111 6
#327190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#327200000000
0!
0%
b0 *
0-
02
b0 6
#327210000000
1!
1%
1-
12
#327220000000
0!
0%
b1 *
0-
02
b1 6
#327230000000
1!
1%
1-
12
#327240000000
0!
0%
b10 *
0-
02
b10 6
#327250000000
1!
1%
1-
12
#327260000000
0!
0%
b11 *
0-
02
b11 6
#327270000000
1!
1%
1-
12
15
#327280000000
0!
0%
b100 *
0-
02
b100 6
#327290000000
1!
1%
1-
12
#327300000000
0!
0%
b101 *
0-
02
b101 6
#327310000000
1!
1%
1-
12
#327320000000
0!
0%
b110 *
0-
02
b110 6
#327330000000
1!
1%
1-
12
#327340000000
0!
0%
b111 *
0-
02
b111 6
#327350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#327360000000
0!
0%
b0 *
0-
02
b0 6
#327370000000
1!
1%
1-
12
#327380000000
0!
0%
b1 *
0-
02
b1 6
#327390000000
1!
1%
1-
12
#327400000000
0!
0%
b10 *
0-
02
b10 6
#327410000000
1!
1%
1-
12
#327420000000
0!
0%
b11 *
0-
02
b11 6
#327430000000
1!
1%
1-
12
15
#327440000000
0!
0%
b100 *
0-
02
b100 6
#327450000000
1!
1%
1-
12
#327460000000
0!
0%
b101 *
0-
02
b101 6
#327470000000
1!
1%
1-
12
#327480000000
0!
0%
b110 *
0-
02
b110 6
#327490000000
1!
1%
1-
12
#327500000000
0!
0%
b111 *
0-
02
b111 6
#327510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#327520000000
0!
0%
b0 *
0-
02
b0 6
#327530000000
1!
1%
1-
12
#327540000000
0!
0%
b1 *
0-
02
b1 6
#327550000000
1!
1%
1-
12
#327560000000
0!
0%
b10 *
0-
02
b10 6
#327570000000
1!
1%
1-
12
#327580000000
0!
0%
b11 *
0-
02
b11 6
#327590000000
1!
1%
1-
12
15
#327600000000
0!
0%
b100 *
0-
02
b100 6
#327610000000
1!
1%
1-
12
#327620000000
0!
0%
b101 *
0-
02
b101 6
#327630000000
1!
1%
1-
12
#327640000000
0!
0%
b110 *
0-
02
b110 6
#327650000000
1!
1%
1-
12
#327660000000
0!
0%
b111 *
0-
02
b111 6
#327670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#327680000000
0!
0%
b0 *
0-
02
b0 6
#327690000000
1!
1%
1-
12
#327700000000
0!
0%
b1 *
0-
02
b1 6
#327710000000
1!
1%
1-
12
#327720000000
0!
0%
b10 *
0-
02
b10 6
#327730000000
1!
1%
1-
12
#327740000000
0!
0%
b11 *
0-
02
b11 6
#327750000000
1!
1%
1-
12
15
#327760000000
0!
0%
b100 *
0-
02
b100 6
#327770000000
1!
1%
1-
12
#327780000000
0!
0%
b101 *
0-
02
b101 6
#327790000000
1!
1%
1-
12
#327800000000
0!
0%
b110 *
0-
02
b110 6
#327810000000
1!
1%
1-
12
#327820000000
0!
0%
b111 *
0-
02
b111 6
#327830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#327840000000
0!
0%
b0 *
0-
02
b0 6
#327850000000
1!
1%
1-
12
#327860000000
0!
0%
b1 *
0-
02
b1 6
#327870000000
1!
1%
1-
12
#327880000000
0!
0%
b10 *
0-
02
b10 6
#327890000000
1!
1%
1-
12
#327900000000
0!
0%
b11 *
0-
02
b11 6
#327910000000
1!
1%
1-
12
15
#327920000000
0!
0%
b100 *
0-
02
b100 6
#327930000000
1!
1%
1-
12
#327940000000
0!
0%
b101 *
0-
02
b101 6
#327950000000
1!
1%
1-
12
#327960000000
0!
0%
b110 *
0-
02
b110 6
#327970000000
1!
1%
1-
12
#327980000000
0!
0%
b111 *
0-
02
b111 6
#327990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#328000000000
0!
0%
b0 *
0-
02
b0 6
#328010000000
1!
1%
1-
12
#328020000000
0!
0%
b1 *
0-
02
b1 6
#328030000000
1!
1%
1-
12
#328040000000
0!
0%
b10 *
0-
02
b10 6
#328050000000
1!
1%
1-
12
#328060000000
0!
0%
b11 *
0-
02
b11 6
#328070000000
1!
1%
1-
12
15
#328080000000
0!
0%
b100 *
0-
02
b100 6
#328090000000
1!
1%
1-
12
#328100000000
0!
0%
b101 *
0-
02
b101 6
#328110000000
1!
1%
1-
12
#328120000000
0!
0%
b110 *
0-
02
b110 6
#328130000000
1!
1%
1-
12
#328140000000
0!
0%
b111 *
0-
02
b111 6
#328150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#328160000000
0!
0%
b0 *
0-
02
b0 6
#328170000000
1!
1%
1-
12
#328180000000
0!
0%
b1 *
0-
02
b1 6
#328190000000
1!
1%
1-
12
#328200000000
0!
0%
b10 *
0-
02
b10 6
#328210000000
1!
1%
1-
12
#328220000000
0!
0%
b11 *
0-
02
b11 6
#328230000000
1!
1%
1-
12
15
#328240000000
0!
0%
b100 *
0-
02
b100 6
#328250000000
1!
1%
1-
12
#328260000000
0!
0%
b101 *
0-
02
b101 6
#328270000000
1!
1%
1-
12
#328280000000
0!
0%
b110 *
0-
02
b110 6
#328290000000
1!
1%
1-
12
#328300000000
0!
0%
b111 *
0-
02
b111 6
#328310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#328320000000
0!
0%
b0 *
0-
02
b0 6
#328330000000
1!
1%
1-
12
#328340000000
0!
0%
b1 *
0-
02
b1 6
#328350000000
1!
1%
1-
12
#328360000000
0!
0%
b10 *
0-
02
b10 6
#328370000000
1!
1%
1-
12
#328380000000
0!
0%
b11 *
0-
02
b11 6
#328390000000
1!
1%
1-
12
15
#328400000000
0!
0%
b100 *
0-
02
b100 6
#328410000000
1!
1%
1-
12
#328420000000
0!
0%
b101 *
0-
02
b101 6
#328430000000
1!
1%
1-
12
#328440000000
0!
0%
b110 *
0-
02
b110 6
#328450000000
1!
1%
1-
12
#328460000000
0!
0%
b111 *
0-
02
b111 6
#328470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#328480000000
0!
0%
b0 *
0-
02
b0 6
#328490000000
1!
1%
1-
12
#328500000000
0!
0%
b1 *
0-
02
b1 6
#328510000000
1!
1%
1-
12
#328520000000
0!
0%
b10 *
0-
02
b10 6
#328530000000
1!
1%
1-
12
#328540000000
0!
0%
b11 *
0-
02
b11 6
#328550000000
1!
1%
1-
12
15
#328560000000
0!
0%
b100 *
0-
02
b100 6
#328570000000
1!
1%
1-
12
#328580000000
0!
0%
b101 *
0-
02
b101 6
#328590000000
1!
1%
1-
12
#328600000000
0!
0%
b110 *
0-
02
b110 6
#328610000000
1!
1%
1-
12
#328620000000
0!
0%
b111 *
0-
02
b111 6
#328630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#328640000000
0!
0%
b0 *
0-
02
b0 6
#328650000000
1!
1%
1-
12
#328660000000
0!
0%
b1 *
0-
02
b1 6
#328670000000
1!
1%
1-
12
#328680000000
0!
0%
b10 *
0-
02
b10 6
#328690000000
1!
1%
1-
12
#328700000000
0!
0%
b11 *
0-
02
b11 6
#328710000000
1!
1%
1-
12
15
#328720000000
0!
0%
b100 *
0-
02
b100 6
#328730000000
1!
1%
1-
12
#328740000000
0!
0%
b101 *
0-
02
b101 6
#328750000000
1!
1%
1-
12
#328760000000
0!
0%
b110 *
0-
02
b110 6
#328770000000
1!
1%
1-
12
#328780000000
0!
0%
b111 *
0-
02
b111 6
#328790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#328800000000
0!
0%
b0 *
0-
02
b0 6
#328810000000
1!
1%
1-
12
#328820000000
0!
0%
b1 *
0-
02
b1 6
#328830000000
1!
1%
1-
12
#328840000000
0!
0%
b10 *
0-
02
b10 6
#328850000000
1!
1%
1-
12
#328860000000
0!
0%
b11 *
0-
02
b11 6
#328870000000
1!
1%
1-
12
15
#328880000000
0!
0%
b100 *
0-
02
b100 6
#328890000000
1!
1%
1-
12
#328900000000
0!
0%
b101 *
0-
02
b101 6
#328910000000
1!
1%
1-
12
#328920000000
0!
0%
b110 *
0-
02
b110 6
#328930000000
1!
1%
1-
12
#328940000000
0!
0%
b111 *
0-
02
b111 6
#328950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#328960000000
0!
0%
b0 *
0-
02
b0 6
#328970000000
1!
1%
1-
12
#328980000000
0!
0%
b1 *
0-
02
b1 6
#328990000000
1!
1%
1-
12
#329000000000
0!
0%
b10 *
0-
02
b10 6
#329010000000
1!
1%
1-
12
#329020000000
0!
0%
b11 *
0-
02
b11 6
#329030000000
1!
1%
1-
12
15
#329040000000
0!
0%
b100 *
0-
02
b100 6
#329050000000
1!
1%
1-
12
#329060000000
0!
0%
b101 *
0-
02
b101 6
#329070000000
1!
1%
1-
12
#329080000000
0!
0%
b110 *
0-
02
b110 6
#329090000000
1!
1%
1-
12
#329100000000
0!
0%
b111 *
0-
02
b111 6
#329110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#329120000000
0!
0%
b0 *
0-
02
b0 6
#329130000000
1!
1%
1-
12
#329140000000
0!
0%
b1 *
0-
02
b1 6
#329150000000
1!
1%
1-
12
#329160000000
0!
0%
b10 *
0-
02
b10 6
#329170000000
1!
1%
1-
12
#329180000000
0!
0%
b11 *
0-
02
b11 6
#329190000000
1!
1%
1-
12
15
#329200000000
0!
0%
b100 *
0-
02
b100 6
#329210000000
1!
1%
1-
12
#329220000000
0!
0%
b101 *
0-
02
b101 6
#329230000000
1!
1%
1-
12
#329240000000
0!
0%
b110 *
0-
02
b110 6
#329250000000
1!
1%
1-
12
#329260000000
0!
0%
b111 *
0-
02
b111 6
#329270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#329280000000
0!
0%
b0 *
0-
02
b0 6
#329290000000
1!
1%
1-
12
#329300000000
0!
0%
b1 *
0-
02
b1 6
#329310000000
1!
1%
1-
12
#329320000000
0!
0%
b10 *
0-
02
b10 6
#329330000000
1!
1%
1-
12
#329340000000
0!
0%
b11 *
0-
02
b11 6
#329350000000
1!
1%
1-
12
15
#329360000000
0!
0%
b100 *
0-
02
b100 6
#329370000000
1!
1%
1-
12
#329380000000
0!
0%
b101 *
0-
02
b101 6
#329390000000
1!
1%
1-
12
#329400000000
0!
0%
b110 *
0-
02
b110 6
#329410000000
1!
1%
1-
12
#329420000000
0!
0%
b111 *
0-
02
b111 6
#329430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#329440000000
0!
0%
b0 *
0-
02
b0 6
#329450000000
1!
1%
1-
12
#329460000000
0!
0%
b1 *
0-
02
b1 6
#329470000000
1!
1%
1-
12
#329480000000
0!
0%
b10 *
0-
02
b10 6
#329490000000
1!
1%
1-
12
#329500000000
0!
0%
b11 *
0-
02
b11 6
#329510000000
1!
1%
1-
12
15
#329520000000
0!
0%
b100 *
0-
02
b100 6
#329530000000
1!
1%
1-
12
#329540000000
0!
0%
b101 *
0-
02
b101 6
#329550000000
1!
1%
1-
12
#329560000000
0!
0%
b110 *
0-
02
b110 6
#329570000000
1!
1%
1-
12
#329580000000
0!
0%
b111 *
0-
02
b111 6
#329590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#329600000000
0!
0%
b0 *
0-
02
b0 6
#329610000000
1!
1%
1-
12
#329620000000
0!
0%
b1 *
0-
02
b1 6
#329630000000
1!
1%
1-
12
#329640000000
0!
0%
b10 *
0-
02
b10 6
#329650000000
1!
1%
1-
12
#329660000000
0!
0%
b11 *
0-
02
b11 6
#329670000000
1!
1%
1-
12
15
#329680000000
0!
0%
b100 *
0-
02
b100 6
#329690000000
1!
1%
1-
12
#329700000000
0!
0%
b101 *
0-
02
b101 6
#329710000000
1!
1%
1-
12
#329720000000
0!
0%
b110 *
0-
02
b110 6
#329730000000
1!
1%
1-
12
#329740000000
0!
0%
b111 *
0-
02
b111 6
#329750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#329760000000
0!
0%
b0 *
0-
02
b0 6
#329770000000
1!
1%
1-
12
#329780000000
0!
0%
b1 *
0-
02
b1 6
#329790000000
1!
1%
1-
12
#329800000000
0!
0%
b10 *
0-
02
b10 6
#329810000000
1!
1%
1-
12
#329820000000
0!
0%
b11 *
0-
02
b11 6
#329830000000
1!
1%
1-
12
15
#329840000000
0!
0%
b100 *
0-
02
b100 6
#329850000000
1!
1%
1-
12
#329860000000
0!
0%
b101 *
0-
02
b101 6
#329870000000
1!
1%
1-
12
#329880000000
0!
0%
b110 *
0-
02
b110 6
#329890000000
1!
1%
1-
12
#329900000000
0!
0%
b111 *
0-
02
b111 6
#329910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#329920000000
0!
0%
b0 *
0-
02
b0 6
#329930000000
1!
1%
1-
12
#329940000000
0!
0%
b1 *
0-
02
b1 6
#329950000000
1!
1%
1-
12
#329960000000
0!
0%
b10 *
0-
02
b10 6
#329970000000
1!
1%
1-
12
#329980000000
0!
0%
b11 *
0-
02
b11 6
#329990000000
1!
1%
1-
12
15
#330000000000
0!
0%
b100 *
0-
02
b100 6
#330010000000
1!
1%
1-
12
#330020000000
0!
0%
b101 *
0-
02
b101 6
#330030000000
1!
1%
1-
12
#330040000000
0!
0%
b110 *
0-
02
b110 6
#330050000000
1!
1%
1-
12
#330060000000
0!
0%
b111 *
0-
02
b111 6
#330070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#330080000000
0!
0%
b0 *
0-
02
b0 6
#330090000000
1!
1%
1-
12
#330100000000
0!
0%
b1 *
0-
02
b1 6
#330110000000
1!
1%
1-
12
#330120000000
0!
0%
b10 *
0-
02
b10 6
#330130000000
1!
1%
1-
12
#330140000000
0!
0%
b11 *
0-
02
b11 6
#330150000000
1!
1%
1-
12
15
#330160000000
0!
0%
b100 *
0-
02
b100 6
#330170000000
1!
1%
1-
12
#330180000000
0!
0%
b101 *
0-
02
b101 6
#330190000000
1!
1%
1-
12
#330200000000
0!
0%
b110 *
0-
02
b110 6
#330210000000
1!
1%
1-
12
#330220000000
0!
0%
b111 *
0-
02
b111 6
#330230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#330240000000
0!
0%
b0 *
0-
02
b0 6
#330250000000
1!
1%
1-
12
#330260000000
0!
0%
b1 *
0-
02
b1 6
#330270000000
1!
1%
1-
12
#330280000000
0!
0%
b10 *
0-
02
b10 6
#330290000000
1!
1%
1-
12
#330300000000
0!
0%
b11 *
0-
02
b11 6
#330310000000
1!
1%
1-
12
15
#330320000000
0!
0%
b100 *
0-
02
b100 6
#330330000000
1!
1%
1-
12
#330340000000
0!
0%
b101 *
0-
02
b101 6
#330350000000
1!
1%
1-
12
#330360000000
0!
0%
b110 *
0-
02
b110 6
#330370000000
1!
1%
1-
12
#330380000000
0!
0%
b111 *
0-
02
b111 6
#330390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#330400000000
0!
0%
b0 *
0-
02
b0 6
#330410000000
1!
1%
1-
12
#330420000000
0!
0%
b1 *
0-
02
b1 6
#330430000000
1!
1%
1-
12
#330440000000
0!
0%
b10 *
0-
02
b10 6
#330450000000
1!
1%
1-
12
#330460000000
0!
0%
b11 *
0-
02
b11 6
#330470000000
1!
1%
1-
12
15
#330480000000
0!
0%
b100 *
0-
02
b100 6
#330490000000
1!
1%
1-
12
#330500000000
0!
0%
b101 *
0-
02
b101 6
#330510000000
1!
1%
1-
12
#330520000000
0!
0%
b110 *
0-
02
b110 6
#330530000000
1!
1%
1-
12
#330540000000
0!
0%
b111 *
0-
02
b111 6
#330550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#330560000000
0!
0%
b0 *
0-
02
b0 6
#330570000000
1!
1%
1-
12
#330580000000
0!
0%
b1 *
0-
02
b1 6
#330590000000
1!
1%
1-
12
#330600000000
0!
0%
b10 *
0-
02
b10 6
#330610000000
1!
1%
1-
12
#330620000000
0!
0%
b11 *
0-
02
b11 6
#330630000000
1!
1%
1-
12
15
#330640000000
0!
0%
b100 *
0-
02
b100 6
#330650000000
1!
1%
1-
12
#330660000000
0!
0%
b101 *
0-
02
b101 6
#330670000000
1!
1%
1-
12
#330680000000
0!
0%
b110 *
0-
02
b110 6
#330690000000
1!
1%
1-
12
#330700000000
0!
0%
b111 *
0-
02
b111 6
#330710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#330720000000
0!
0%
b0 *
0-
02
b0 6
#330730000000
1!
1%
1-
12
#330740000000
0!
0%
b1 *
0-
02
b1 6
#330750000000
1!
1%
1-
12
#330760000000
0!
0%
b10 *
0-
02
b10 6
#330770000000
1!
1%
1-
12
#330780000000
0!
0%
b11 *
0-
02
b11 6
#330790000000
1!
1%
1-
12
15
#330800000000
0!
0%
b100 *
0-
02
b100 6
#330810000000
1!
1%
1-
12
#330820000000
0!
0%
b101 *
0-
02
b101 6
#330830000000
1!
1%
1-
12
#330840000000
0!
0%
b110 *
0-
02
b110 6
#330850000000
1!
1%
1-
12
#330860000000
0!
0%
b111 *
0-
02
b111 6
#330870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#330880000000
0!
0%
b0 *
0-
02
b0 6
#330890000000
1!
1%
1-
12
#330900000000
0!
0%
b1 *
0-
02
b1 6
#330910000000
1!
1%
1-
12
#330920000000
0!
0%
b10 *
0-
02
b10 6
#330930000000
1!
1%
1-
12
#330940000000
0!
0%
b11 *
0-
02
b11 6
#330950000000
1!
1%
1-
12
15
#330960000000
0!
0%
b100 *
0-
02
b100 6
#330970000000
1!
1%
1-
12
#330980000000
0!
0%
b101 *
0-
02
b101 6
#330990000000
1!
1%
1-
12
#331000000000
0!
0%
b110 *
0-
02
b110 6
#331010000000
1!
1%
1-
12
#331020000000
0!
0%
b111 *
0-
02
b111 6
#331030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#331040000000
0!
0%
b0 *
0-
02
b0 6
#331050000000
1!
1%
1-
12
#331060000000
0!
0%
b1 *
0-
02
b1 6
#331070000000
1!
1%
1-
12
#331080000000
0!
0%
b10 *
0-
02
b10 6
#331090000000
1!
1%
1-
12
#331100000000
0!
0%
b11 *
0-
02
b11 6
#331110000000
1!
1%
1-
12
15
#331120000000
0!
0%
b100 *
0-
02
b100 6
#331130000000
1!
1%
1-
12
#331140000000
0!
0%
b101 *
0-
02
b101 6
#331150000000
1!
1%
1-
12
#331160000000
0!
0%
b110 *
0-
02
b110 6
#331170000000
1!
1%
1-
12
#331180000000
0!
0%
b111 *
0-
02
b111 6
#331190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#331200000000
0!
0%
b0 *
0-
02
b0 6
#331210000000
1!
1%
1-
12
#331220000000
0!
0%
b1 *
0-
02
b1 6
#331230000000
1!
1%
1-
12
#331240000000
0!
0%
b10 *
0-
02
b10 6
#331250000000
1!
1%
1-
12
#331260000000
0!
0%
b11 *
0-
02
b11 6
#331270000000
1!
1%
1-
12
15
#331280000000
0!
0%
b100 *
0-
02
b100 6
#331290000000
1!
1%
1-
12
#331300000000
0!
0%
b101 *
0-
02
b101 6
#331310000000
1!
1%
1-
12
#331320000000
0!
0%
b110 *
0-
02
b110 6
#331330000000
1!
1%
1-
12
#331340000000
0!
0%
b111 *
0-
02
b111 6
#331350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#331360000000
0!
0%
b0 *
0-
02
b0 6
#331370000000
1!
1%
1-
12
#331380000000
0!
0%
b1 *
0-
02
b1 6
#331390000000
1!
1%
1-
12
#331400000000
0!
0%
b10 *
0-
02
b10 6
#331410000000
1!
1%
1-
12
#331420000000
0!
0%
b11 *
0-
02
b11 6
#331430000000
1!
1%
1-
12
15
#331440000000
0!
0%
b100 *
0-
02
b100 6
#331450000000
1!
1%
1-
12
#331460000000
0!
0%
b101 *
0-
02
b101 6
#331470000000
1!
1%
1-
12
#331480000000
0!
0%
b110 *
0-
02
b110 6
#331490000000
1!
1%
1-
12
#331500000000
0!
0%
b111 *
0-
02
b111 6
#331510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#331520000000
0!
0%
b0 *
0-
02
b0 6
#331530000000
1!
1%
1-
12
#331540000000
0!
0%
b1 *
0-
02
b1 6
#331550000000
1!
1%
1-
12
#331560000000
0!
0%
b10 *
0-
02
b10 6
#331570000000
1!
1%
1-
12
#331580000000
0!
0%
b11 *
0-
02
b11 6
#331590000000
1!
1%
1-
12
15
#331600000000
0!
0%
b100 *
0-
02
b100 6
#331610000000
1!
1%
1-
12
#331620000000
0!
0%
b101 *
0-
02
b101 6
#331630000000
1!
1%
1-
12
#331640000000
0!
0%
b110 *
0-
02
b110 6
#331650000000
1!
1%
1-
12
#331660000000
0!
0%
b111 *
0-
02
b111 6
#331670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#331680000000
0!
0%
b0 *
0-
02
b0 6
#331690000000
1!
1%
1-
12
#331700000000
0!
0%
b1 *
0-
02
b1 6
#331710000000
1!
1%
1-
12
#331720000000
0!
0%
b10 *
0-
02
b10 6
#331730000000
1!
1%
1-
12
#331740000000
0!
0%
b11 *
0-
02
b11 6
#331750000000
1!
1%
1-
12
15
#331760000000
0!
0%
b100 *
0-
02
b100 6
#331770000000
1!
1%
1-
12
#331780000000
0!
0%
b101 *
0-
02
b101 6
#331790000000
1!
1%
1-
12
#331800000000
0!
0%
b110 *
0-
02
b110 6
#331810000000
1!
1%
1-
12
#331820000000
0!
0%
b111 *
0-
02
b111 6
#331830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#331840000000
0!
0%
b0 *
0-
02
b0 6
#331850000000
1!
1%
1-
12
#331860000000
0!
0%
b1 *
0-
02
b1 6
#331870000000
1!
1%
1-
12
#331880000000
0!
0%
b10 *
0-
02
b10 6
#331890000000
1!
1%
1-
12
#331900000000
0!
0%
b11 *
0-
02
b11 6
#331910000000
1!
1%
1-
12
15
#331920000000
0!
0%
b100 *
0-
02
b100 6
#331930000000
1!
1%
1-
12
#331940000000
0!
0%
b101 *
0-
02
b101 6
#331950000000
1!
1%
1-
12
#331960000000
0!
0%
b110 *
0-
02
b110 6
#331970000000
1!
1%
1-
12
#331980000000
0!
0%
b111 *
0-
02
b111 6
#331990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#332000000000
0!
0%
b0 *
0-
02
b0 6
#332010000000
1!
1%
1-
12
#332020000000
0!
0%
b1 *
0-
02
b1 6
#332030000000
1!
1%
1-
12
#332040000000
0!
0%
b10 *
0-
02
b10 6
#332050000000
1!
1%
1-
12
#332060000000
0!
0%
b11 *
0-
02
b11 6
#332070000000
1!
1%
1-
12
15
#332080000000
0!
0%
b100 *
0-
02
b100 6
#332090000000
1!
1%
1-
12
#332100000000
0!
0%
b101 *
0-
02
b101 6
#332110000000
1!
1%
1-
12
#332120000000
0!
0%
b110 *
0-
02
b110 6
#332130000000
1!
1%
1-
12
#332140000000
0!
0%
b111 *
0-
02
b111 6
#332150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#332160000000
0!
0%
b0 *
0-
02
b0 6
#332170000000
1!
1%
1-
12
#332180000000
0!
0%
b1 *
0-
02
b1 6
#332190000000
1!
1%
1-
12
#332200000000
0!
0%
b10 *
0-
02
b10 6
#332210000000
1!
1%
1-
12
#332220000000
0!
0%
b11 *
0-
02
b11 6
#332230000000
1!
1%
1-
12
15
#332240000000
0!
0%
b100 *
0-
02
b100 6
#332250000000
1!
1%
1-
12
#332260000000
0!
0%
b101 *
0-
02
b101 6
#332270000000
1!
1%
1-
12
#332280000000
0!
0%
b110 *
0-
02
b110 6
#332290000000
1!
1%
1-
12
#332300000000
0!
0%
b111 *
0-
02
b111 6
#332310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#332320000000
0!
0%
b0 *
0-
02
b0 6
#332330000000
1!
1%
1-
12
#332340000000
0!
0%
b1 *
0-
02
b1 6
#332350000000
1!
1%
1-
12
#332360000000
0!
0%
b10 *
0-
02
b10 6
#332370000000
1!
1%
1-
12
#332380000000
0!
0%
b11 *
0-
02
b11 6
#332390000000
1!
1%
1-
12
15
#332400000000
0!
0%
b100 *
0-
02
b100 6
#332410000000
1!
1%
1-
12
#332420000000
0!
0%
b101 *
0-
02
b101 6
#332430000000
1!
1%
1-
12
#332440000000
0!
0%
b110 *
0-
02
b110 6
#332450000000
1!
1%
1-
12
#332460000000
0!
0%
b111 *
0-
02
b111 6
#332470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#332480000000
0!
0%
b0 *
0-
02
b0 6
#332490000000
1!
1%
1-
12
#332500000000
0!
0%
b1 *
0-
02
b1 6
#332510000000
1!
1%
1-
12
#332520000000
0!
0%
b10 *
0-
02
b10 6
#332530000000
1!
1%
1-
12
#332540000000
0!
0%
b11 *
0-
02
b11 6
#332550000000
1!
1%
1-
12
15
#332560000000
0!
0%
b100 *
0-
02
b100 6
#332570000000
1!
1%
1-
12
#332580000000
0!
0%
b101 *
0-
02
b101 6
#332590000000
1!
1%
1-
12
#332600000000
0!
0%
b110 *
0-
02
b110 6
#332610000000
1!
1%
1-
12
#332620000000
0!
0%
b111 *
0-
02
b111 6
#332630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#332640000000
0!
0%
b0 *
0-
02
b0 6
#332650000000
1!
1%
1-
12
#332660000000
0!
0%
b1 *
0-
02
b1 6
#332670000000
1!
1%
1-
12
#332680000000
0!
0%
b10 *
0-
02
b10 6
#332690000000
1!
1%
1-
12
#332700000000
0!
0%
b11 *
0-
02
b11 6
#332710000000
1!
1%
1-
12
15
#332720000000
0!
0%
b100 *
0-
02
b100 6
#332730000000
1!
1%
1-
12
#332740000000
0!
0%
b101 *
0-
02
b101 6
#332750000000
1!
1%
1-
12
#332760000000
0!
0%
b110 *
0-
02
b110 6
#332770000000
1!
1%
1-
12
#332780000000
0!
0%
b111 *
0-
02
b111 6
#332790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#332800000000
0!
0%
b0 *
0-
02
b0 6
#332810000000
1!
1%
1-
12
#332820000000
0!
0%
b1 *
0-
02
b1 6
#332830000000
1!
1%
1-
12
#332840000000
0!
0%
b10 *
0-
02
b10 6
#332850000000
1!
1%
1-
12
#332860000000
0!
0%
b11 *
0-
02
b11 6
#332870000000
1!
1%
1-
12
15
#332880000000
0!
0%
b100 *
0-
02
b100 6
#332890000000
1!
1%
1-
12
#332900000000
0!
0%
b101 *
0-
02
b101 6
#332910000000
1!
1%
1-
12
#332920000000
0!
0%
b110 *
0-
02
b110 6
#332930000000
1!
1%
1-
12
#332940000000
0!
0%
b111 *
0-
02
b111 6
#332950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#332960000000
0!
0%
b0 *
0-
02
b0 6
#332970000000
1!
1%
1-
12
#332980000000
0!
0%
b1 *
0-
02
b1 6
#332990000000
1!
1%
1-
12
#333000000000
0!
0%
b10 *
0-
02
b10 6
#333010000000
1!
1%
1-
12
#333020000000
0!
0%
b11 *
0-
02
b11 6
#333030000000
1!
1%
1-
12
15
#333040000000
0!
0%
b100 *
0-
02
b100 6
#333050000000
1!
1%
1-
12
#333060000000
0!
0%
b101 *
0-
02
b101 6
#333070000000
1!
1%
1-
12
#333080000000
0!
0%
b110 *
0-
02
b110 6
#333090000000
1!
1%
1-
12
#333100000000
0!
0%
b111 *
0-
02
b111 6
#333110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#333120000000
0!
0%
b0 *
0-
02
b0 6
#333130000000
1!
1%
1-
12
#333140000000
0!
0%
b1 *
0-
02
b1 6
#333150000000
1!
1%
1-
12
#333160000000
0!
0%
b10 *
0-
02
b10 6
#333170000000
1!
1%
1-
12
#333180000000
0!
0%
b11 *
0-
02
b11 6
#333190000000
1!
1%
1-
12
15
#333200000000
0!
0%
b100 *
0-
02
b100 6
#333210000000
1!
1%
1-
12
#333220000000
0!
0%
b101 *
0-
02
b101 6
#333230000000
1!
1%
1-
12
#333240000000
0!
0%
b110 *
0-
02
b110 6
#333250000000
1!
1%
1-
12
#333260000000
0!
0%
b111 *
0-
02
b111 6
#333270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#333280000000
0!
0%
b0 *
0-
02
b0 6
#333290000000
1!
1%
1-
12
#333300000000
0!
0%
b1 *
0-
02
b1 6
#333310000000
1!
1%
1-
12
#333320000000
0!
0%
b10 *
0-
02
b10 6
#333330000000
1!
1%
1-
12
#333340000000
0!
0%
b11 *
0-
02
b11 6
#333350000000
1!
1%
1-
12
15
#333360000000
0!
0%
b100 *
0-
02
b100 6
#333370000000
1!
1%
1-
12
#333380000000
0!
0%
b101 *
0-
02
b101 6
#333390000000
1!
1%
1-
12
#333400000000
0!
0%
b110 *
0-
02
b110 6
#333410000000
1!
1%
1-
12
#333420000000
0!
0%
b111 *
0-
02
b111 6
#333430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#333440000000
0!
0%
b0 *
0-
02
b0 6
#333450000000
1!
1%
1-
12
#333460000000
0!
0%
b1 *
0-
02
b1 6
#333470000000
1!
1%
1-
12
#333480000000
0!
0%
b10 *
0-
02
b10 6
#333490000000
1!
1%
1-
12
#333500000000
0!
0%
b11 *
0-
02
b11 6
#333510000000
1!
1%
1-
12
15
#333520000000
0!
0%
b100 *
0-
02
b100 6
#333530000000
1!
1%
1-
12
#333540000000
0!
0%
b101 *
0-
02
b101 6
#333550000000
1!
1%
1-
12
#333560000000
0!
0%
b110 *
0-
02
b110 6
#333570000000
1!
1%
1-
12
#333580000000
0!
0%
b111 *
0-
02
b111 6
#333590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#333600000000
0!
0%
b0 *
0-
02
b0 6
#333610000000
1!
1%
1-
12
#333620000000
0!
0%
b1 *
0-
02
b1 6
#333630000000
1!
1%
1-
12
#333640000000
0!
0%
b10 *
0-
02
b10 6
#333650000000
1!
1%
1-
12
#333660000000
0!
0%
b11 *
0-
02
b11 6
#333670000000
1!
1%
1-
12
15
#333680000000
0!
0%
b100 *
0-
02
b100 6
#333690000000
1!
1%
1-
12
#333700000000
0!
0%
b101 *
0-
02
b101 6
#333710000000
1!
1%
1-
12
#333720000000
0!
0%
b110 *
0-
02
b110 6
#333730000000
1!
1%
1-
12
#333740000000
0!
0%
b111 *
0-
02
b111 6
#333750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#333760000000
0!
0%
b0 *
0-
02
b0 6
#333770000000
1!
1%
1-
12
#333780000000
0!
0%
b1 *
0-
02
b1 6
#333790000000
1!
1%
1-
12
#333800000000
0!
0%
b10 *
0-
02
b10 6
#333810000000
1!
1%
1-
12
#333820000000
0!
0%
b11 *
0-
02
b11 6
#333830000000
1!
1%
1-
12
15
#333840000000
0!
0%
b100 *
0-
02
b100 6
#333850000000
1!
1%
1-
12
#333860000000
0!
0%
b101 *
0-
02
b101 6
#333870000000
1!
1%
1-
12
#333880000000
0!
0%
b110 *
0-
02
b110 6
#333890000000
1!
1%
1-
12
#333900000000
0!
0%
b111 *
0-
02
b111 6
#333910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#333920000000
0!
0%
b0 *
0-
02
b0 6
#333930000000
1!
1%
1-
12
#333940000000
0!
0%
b1 *
0-
02
b1 6
#333950000000
1!
1%
1-
12
#333960000000
0!
0%
b10 *
0-
02
b10 6
#333970000000
1!
1%
1-
12
#333980000000
0!
0%
b11 *
0-
02
b11 6
#333990000000
1!
1%
1-
12
15
#334000000000
0!
0%
b100 *
0-
02
b100 6
#334010000000
1!
1%
1-
12
#334020000000
0!
0%
b101 *
0-
02
b101 6
#334030000000
1!
1%
1-
12
#334040000000
0!
0%
b110 *
0-
02
b110 6
#334050000000
1!
1%
1-
12
#334060000000
0!
0%
b111 *
0-
02
b111 6
#334070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#334080000000
0!
0%
b0 *
0-
02
b0 6
#334090000000
1!
1%
1-
12
#334100000000
0!
0%
b1 *
0-
02
b1 6
#334110000000
1!
1%
1-
12
#334120000000
0!
0%
b10 *
0-
02
b10 6
#334130000000
1!
1%
1-
12
#334140000000
0!
0%
b11 *
0-
02
b11 6
#334150000000
1!
1%
1-
12
15
#334160000000
0!
0%
b100 *
0-
02
b100 6
#334170000000
1!
1%
1-
12
#334180000000
0!
0%
b101 *
0-
02
b101 6
#334190000000
1!
1%
1-
12
#334200000000
0!
0%
b110 *
0-
02
b110 6
#334210000000
1!
1%
1-
12
#334220000000
0!
0%
b111 *
0-
02
b111 6
#334230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#334240000000
0!
0%
b0 *
0-
02
b0 6
#334250000000
1!
1%
1-
12
#334260000000
0!
0%
b1 *
0-
02
b1 6
#334270000000
1!
1%
1-
12
#334280000000
0!
0%
b10 *
0-
02
b10 6
#334290000000
1!
1%
1-
12
#334300000000
0!
0%
b11 *
0-
02
b11 6
#334310000000
1!
1%
1-
12
15
#334320000000
0!
0%
b100 *
0-
02
b100 6
#334330000000
1!
1%
1-
12
#334340000000
0!
0%
b101 *
0-
02
b101 6
#334350000000
1!
1%
1-
12
#334360000000
0!
0%
b110 *
0-
02
b110 6
#334370000000
1!
1%
1-
12
#334380000000
0!
0%
b111 *
0-
02
b111 6
#334390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#334400000000
0!
0%
b0 *
0-
02
b0 6
#334410000000
1!
1%
1-
12
#334420000000
0!
0%
b1 *
0-
02
b1 6
#334430000000
1!
1%
1-
12
#334440000000
0!
0%
b10 *
0-
02
b10 6
#334450000000
1!
1%
1-
12
#334460000000
0!
0%
b11 *
0-
02
b11 6
#334470000000
1!
1%
1-
12
15
#334480000000
0!
0%
b100 *
0-
02
b100 6
#334490000000
1!
1%
1-
12
#334500000000
0!
0%
b101 *
0-
02
b101 6
#334510000000
1!
1%
1-
12
#334520000000
0!
0%
b110 *
0-
02
b110 6
#334530000000
1!
1%
1-
12
#334540000000
0!
0%
b111 *
0-
02
b111 6
#334550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#334560000000
0!
0%
b0 *
0-
02
b0 6
#334570000000
1!
1%
1-
12
#334580000000
0!
0%
b1 *
0-
02
b1 6
#334590000000
1!
1%
1-
12
#334600000000
0!
0%
b10 *
0-
02
b10 6
#334610000000
1!
1%
1-
12
#334620000000
0!
0%
b11 *
0-
02
b11 6
#334630000000
1!
1%
1-
12
15
#334640000000
0!
0%
b100 *
0-
02
b100 6
#334650000000
1!
1%
1-
12
#334660000000
0!
0%
b101 *
0-
02
b101 6
#334670000000
1!
1%
1-
12
#334680000000
0!
0%
b110 *
0-
02
b110 6
#334690000000
1!
1%
1-
12
#334700000000
0!
0%
b111 *
0-
02
b111 6
#334710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#334720000000
0!
0%
b0 *
0-
02
b0 6
#334730000000
1!
1%
1-
12
#334740000000
0!
0%
b1 *
0-
02
b1 6
#334750000000
1!
1%
1-
12
#334760000000
0!
0%
b10 *
0-
02
b10 6
#334770000000
1!
1%
1-
12
#334780000000
0!
0%
b11 *
0-
02
b11 6
#334790000000
1!
1%
1-
12
15
#334800000000
0!
0%
b100 *
0-
02
b100 6
#334810000000
1!
1%
1-
12
#334820000000
0!
0%
b101 *
0-
02
b101 6
#334830000000
1!
1%
1-
12
#334840000000
0!
0%
b110 *
0-
02
b110 6
#334850000000
1!
1%
1-
12
#334860000000
0!
0%
b111 *
0-
02
b111 6
#334870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#334880000000
0!
0%
b0 *
0-
02
b0 6
#334890000000
1!
1%
1-
12
#334900000000
0!
0%
b1 *
0-
02
b1 6
#334910000000
1!
1%
1-
12
#334920000000
0!
0%
b10 *
0-
02
b10 6
#334930000000
1!
1%
1-
12
#334940000000
0!
0%
b11 *
0-
02
b11 6
#334950000000
1!
1%
1-
12
15
#334960000000
0!
0%
b100 *
0-
02
b100 6
#334970000000
1!
1%
1-
12
#334980000000
0!
0%
b101 *
0-
02
b101 6
#334990000000
1!
1%
1-
12
#335000000000
0!
0%
b110 *
0-
02
b110 6
#335010000000
1!
1%
1-
12
#335020000000
0!
0%
b111 *
0-
02
b111 6
#335030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#335040000000
0!
0%
b0 *
0-
02
b0 6
#335050000000
1!
1%
1-
12
#335060000000
0!
0%
b1 *
0-
02
b1 6
#335070000000
1!
1%
1-
12
#335080000000
0!
0%
b10 *
0-
02
b10 6
#335090000000
1!
1%
1-
12
#335100000000
0!
0%
b11 *
0-
02
b11 6
#335110000000
1!
1%
1-
12
15
#335120000000
0!
0%
b100 *
0-
02
b100 6
#335130000000
1!
1%
1-
12
#335140000000
0!
0%
b101 *
0-
02
b101 6
#335150000000
1!
1%
1-
12
#335160000000
0!
0%
b110 *
0-
02
b110 6
#335170000000
1!
1%
1-
12
#335180000000
0!
0%
b111 *
0-
02
b111 6
#335190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#335200000000
0!
0%
b0 *
0-
02
b0 6
#335210000000
1!
1%
1-
12
#335220000000
0!
0%
b1 *
0-
02
b1 6
#335230000000
1!
1%
1-
12
#335240000000
0!
0%
b10 *
0-
02
b10 6
#335250000000
1!
1%
1-
12
#335260000000
0!
0%
b11 *
0-
02
b11 6
#335270000000
1!
1%
1-
12
15
#335280000000
0!
0%
b100 *
0-
02
b100 6
#335290000000
1!
1%
1-
12
#335300000000
0!
0%
b101 *
0-
02
b101 6
#335310000000
1!
1%
1-
12
#335320000000
0!
0%
b110 *
0-
02
b110 6
#335330000000
1!
1%
1-
12
#335340000000
0!
0%
b111 *
0-
02
b111 6
#335350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#335360000000
0!
0%
b0 *
0-
02
b0 6
#335370000000
1!
1%
1-
12
#335380000000
0!
0%
b1 *
0-
02
b1 6
#335390000000
1!
1%
1-
12
#335400000000
0!
0%
b10 *
0-
02
b10 6
#335410000000
1!
1%
1-
12
#335420000000
0!
0%
b11 *
0-
02
b11 6
#335430000000
1!
1%
1-
12
15
#335440000000
0!
0%
b100 *
0-
02
b100 6
#335450000000
1!
1%
1-
12
#335460000000
0!
0%
b101 *
0-
02
b101 6
#335470000000
1!
1%
1-
12
#335480000000
0!
0%
b110 *
0-
02
b110 6
#335490000000
1!
1%
1-
12
#335500000000
0!
0%
b111 *
0-
02
b111 6
#335510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#335520000000
0!
0%
b0 *
0-
02
b0 6
#335530000000
1!
1%
1-
12
#335540000000
0!
0%
b1 *
0-
02
b1 6
#335550000000
1!
1%
1-
12
#335560000000
0!
0%
b10 *
0-
02
b10 6
#335570000000
1!
1%
1-
12
#335580000000
0!
0%
b11 *
0-
02
b11 6
#335590000000
1!
1%
1-
12
15
#335600000000
0!
0%
b100 *
0-
02
b100 6
#335610000000
1!
1%
1-
12
#335620000000
0!
0%
b101 *
0-
02
b101 6
#335630000000
1!
1%
1-
12
#335640000000
0!
0%
b110 *
0-
02
b110 6
#335650000000
1!
1%
1-
12
#335660000000
0!
0%
b111 *
0-
02
b111 6
#335670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#335680000000
0!
0%
b0 *
0-
02
b0 6
#335690000000
1!
1%
1-
12
#335700000000
0!
0%
b1 *
0-
02
b1 6
#335710000000
1!
1%
1-
12
#335720000000
0!
0%
b10 *
0-
02
b10 6
#335730000000
1!
1%
1-
12
#335740000000
0!
0%
b11 *
0-
02
b11 6
#335750000000
1!
1%
1-
12
15
#335760000000
0!
0%
b100 *
0-
02
b100 6
#335770000000
1!
1%
1-
12
#335780000000
0!
0%
b101 *
0-
02
b101 6
#335790000000
1!
1%
1-
12
#335800000000
0!
0%
b110 *
0-
02
b110 6
#335810000000
1!
1%
1-
12
#335820000000
0!
0%
b111 *
0-
02
b111 6
#335830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#335840000000
0!
0%
b0 *
0-
02
b0 6
#335850000000
1!
1%
1-
12
#335860000000
0!
0%
b1 *
0-
02
b1 6
#335870000000
1!
1%
1-
12
#335880000000
0!
0%
b10 *
0-
02
b10 6
#335890000000
1!
1%
1-
12
#335900000000
0!
0%
b11 *
0-
02
b11 6
#335910000000
1!
1%
1-
12
15
#335920000000
0!
0%
b100 *
0-
02
b100 6
#335930000000
1!
1%
1-
12
#335940000000
0!
0%
b101 *
0-
02
b101 6
#335950000000
1!
1%
1-
12
#335960000000
0!
0%
b110 *
0-
02
b110 6
#335970000000
1!
1%
1-
12
#335980000000
0!
0%
b111 *
0-
02
b111 6
#335990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#336000000000
0!
0%
b0 *
0-
02
b0 6
#336010000000
1!
1%
1-
12
#336020000000
0!
0%
b1 *
0-
02
b1 6
#336030000000
1!
1%
1-
12
#336040000000
0!
0%
b10 *
0-
02
b10 6
#336050000000
1!
1%
1-
12
#336060000000
0!
0%
b11 *
0-
02
b11 6
#336070000000
1!
1%
1-
12
15
#336080000000
0!
0%
b100 *
0-
02
b100 6
#336090000000
1!
1%
1-
12
#336100000000
0!
0%
b101 *
0-
02
b101 6
#336110000000
1!
1%
1-
12
#336120000000
0!
0%
b110 *
0-
02
b110 6
#336130000000
1!
1%
1-
12
#336140000000
0!
0%
b111 *
0-
02
b111 6
#336150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#336160000000
0!
0%
b0 *
0-
02
b0 6
#336170000000
1!
1%
1-
12
#336180000000
0!
0%
b1 *
0-
02
b1 6
#336190000000
1!
1%
1-
12
#336200000000
0!
0%
b10 *
0-
02
b10 6
#336210000000
1!
1%
1-
12
#336220000000
0!
0%
b11 *
0-
02
b11 6
#336230000000
1!
1%
1-
12
15
#336240000000
0!
0%
b100 *
0-
02
b100 6
#336250000000
1!
1%
1-
12
#336260000000
0!
0%
b101 *
0-
02
b101 6
#336270000000
1!
1%
1-
12
#336280000000
0!
0%
b110 *
0-
02
b110 6
#336290000000
1!
1%
1-
12
#336300000000
0!
0%
b111 *
0-
02
b111 6
#336310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#336320000000
0!
0%
b0 *
0-
02
b0 6
#336330000000
1!
1%
1-
12
#336340000000
0!
0%
b1 *
0-
02
b1 6
#336350000000
1!
1%
1-
12
#336360000000
0!
0%
b10 *
0-
02
b10 6
#336370000000
1!
1%
1-
12
#336380000000
0!
0%
b11 *
0-
02
b11 6
#336390000000
1!
1%
1-
12
15
#336400000000
0!
0%
b100 *
0-
02
b100 6
#336410000000
1!
1%
1-
12
#336420000000
0!
0%
b101 *
0-
02
b101 6
#336430000000
1!
1%
1-
12
#336440000000
0!
0%
b110 *
0-
02
b110 6
#336450000000
1!
1%
1-
12
#336460000000
0!
0%
b111 *
0-
02
b111 6
#336470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#336480000000
0!
0%
b0 *
0-
02
b0 6
#336490000000
1!
1%
1-
12
#336500000000
0!
0%
b1 *
0-
02
b1 6
#336510000000
1!
1%
1-
12
#336520000000
0!
0%
b10 *
0-
02
b10 6
#336530000000
1!
1%
1-
12
#336540000000
0!
0%
b11 *
0-
02
b11 6
#336550000000
1!
1%
1-
12
15
#336560000000
0!
0%
b100 *
0-
02
b100 6
#336570000000
1!
1%
1-
12
#336580000000
0!
0%
b101 *
0-
02
b101 6
#336590000000
1!
1%
1-
12
#336600000000
0!
0%
b110 *
0-
02
b110 6
#336610000000
1!
1%
1-
12
#336620000000
0!
0%
b111 *
0-
02
b111 6
#336630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#336640000000
0!
0%
b0 *
0-
02
b0 6
#336650000000
1!
1%
1-
12
#336660000000
0!
0%
b1 *
0-
02
b1 6
#336670000000
1!
1%
1-
12
#336680000000
0!
0%
b10 *
0-
02
b10 6
#336690000000
1!
1%
1-
12
#336700000000
0!
0%
b11 *
0-
02
b11 6
#336710000000
1!
1%
1-
12
15
#336720000000
0!
0%
b100 *
0-
02
b100 6
#336730000000
1!
1%
1-
12
#336740000000
0!
0%
b101 *
0-
02
b101 6
#336750000000
1!
1%
1-
12
#336760000000
0!
0%
b110 *
0-
02
b110 6
#336770000000
1!
1%
1-
12
#336780000000
0!
0%
b111 *
0-
02
b111 6
#336790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#336800000000
0!
0%
b0 *
0-
02
b0 6
#336810000000
1!
1%
1-
12
#336820000000
0!
0%
b1 *
0-
02
b1 6
#336830000000
1!
1%
1-
12
#336840000000
0!
0%
b10 *
0-
02
b10 6
#336850000000
1!
1%
1-
12
#336860000000
0!
0%
b11 *
0-
02
b11 6
#336870000000
1!
1%
1-
12
15
#336880000000
0!
0%
b100 *
0-
02
b100 6
#336890000000
1!
1%
1-
12
#336900000000
0!
0%
b101 *
0-
02
b101 6
#336910000000
1!
1%
1-
12
#336920000000
0!
0%
b110 *
0-
02
b110 6
#336930000000
1!
1%
1-
12
#336940000000
0!
0%
b111 *
0-
02
b111 6
#336950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#336960000000
0!
0%
b0 *
0-
02
b0 6
#336970000000
1!
1%
1-
12
#336980000000
0!
0%
b1 *
0-
02
b1 6
#336990000000
1!
1%
1-
12
#337000000000
0!
0%
b10 *
0-
02
b10 6
#337010000000
1!
1%
1-
12
#337020000000
0!
0%
b11 *
0-
02
b11 6
#337030000000
1!
1%
1-
12
15
#337040000000
0!
0%
b100 *
0-
02
b100 6
#337050000000
1!
1%
1-
12
#337060000000
0!
0%
b101 *
0-
02
b101 6
#337070000000
1!
1%
1-
12
#337080000000
0!
0%
b110 *
0-
02
b110 6
#337090000000
1!
1%
1-
12
#337100000000
0!
0%
b111 *
0-
02
b111 6
#337110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#337120000000
0!
0%
b0 *
0-
02
b0 6
#337130000000
1!
1%
1-
12
#337140000000
0!
0%
b1 *
0-
02
b1 6
#337150000000
1!
1%
1-
12
#337160000000
0!
0%
b10 *
0-
02
b10 6
#337170000000
1!
1%
1-
12
#337180000000
0!
0%
b11 *
0-
02
b11 6
#337190000000
1!
1%
1-
12
15
#337200000000
0!
0%
b100 *
0-
02
b100 6
#337210000000
1!
1%
1-
12
#337220000000
0!
0%
b101 *
0-
02
b101 6
#337230000000
1!
1%
1-
12
#337240000000
0!
0%
b110 *
0-
02
b110 6
#337250000000
1!
1%
1-
12
#337260000000
0!
0%
b111 *
0-
02
b111 6
#337270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#337280000000
0!
0%
b0 *
0-
02
b0 6
#337290000000
1!
1%
1-
12
#337300000000
0!
0%
b1 *
0-
02
b1 6
#337310000000
1!
1%
1-
12
#337320000000
0!
0%
b10 *
0-
02
b10 6
#337330000000
1!
1%
1-
12
#337340000000
0!
0%
b11 *
0-
02
b11 6
#337350000000
1!
1%
1-
12
15
#337360000000
0!
0%
b100 *
0-
02
b100 6
#337370000000
1!
1%
1-
12
#337380000000
0!
0%
b101 *
0-
02
b101 6
#337390000000
1!
1%
1-
12
#337400000000
0!
0%
b110 *
0-
02
b110 6
#337410000000
1!
1%
1-
12
#337420000000
0!
0%
b111 *
0-
02
b111 6
#337430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#337440000000
0!
0%
b0 *
0-
02
b0 6
#337450000000
1!
1%
1-
12
#337460000000
0!
0%
b1 *
0-
02
b1 6
#337470000000
1!
1%
1-
12
#337480000000
0!
0%
b10 *
0-
02
b10 6
#337490000000
1!
1%
1-
12
#337500000000
0!
0%
b11 *
0-
02
b11 6
#337510000000
1!
1%
1-
12
15
#337520000000
0!
0%
b100 *
0-
02
b100 6
#337530000000
1!
1%
1-
12
#337540000000
0!
0%
b101 *
0-
02
b101 6
#337550000000
1!
1%
1-
12
#337560000000
0!
0%
b110 *
0-
02
b110 6
#337570000000
1!
1%
1-
12
#337580000000
0!
0%
b111 *
0-
02
b111 6
#337590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#337600000000
0!
0%
b0 *
0-
02
b0 6
#337610000000
1!
1%
1-
12
#337620000000
0!
0%
b1 *
0-
02
b1 6
#337630000000
1!
1%
1-
12
#337640000000
0!
0%
b10 *
0-
02
b10 6
#337650000000
1!
1%
1-
12
#337660000000
0!
0%
b11 *
0-
02
b11 6
#337670000000
1!
1%
1-
12
15
#337680000000
0!
0%
b100 *
0-
02
b100 6
#337690000000
1!
1%
1-
12
#337700000000
0!
0%
b101 *
0-
02
b101 6
#337710000000
1!
1%
1-
12
#337720000000
0!
0%
b110 *
0-
02
b110 6
#337730000000
1!
1%
1-
12
#337740000000
0!
0%
b111 *
0-
02
b111 6
#337750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#337760000000
0!
0%
b0 *
0-
02
b0 6
#337770000000
1!
1%
1-
12
#337780000000
0!
0%
b1 *
0-
02
b1 6
#337790000000
1!
1%
1-
12
#337800000000
0!
0%
b10 *
0-
02
b10 6
#337810000000
1!
1%
1-
12
#337820000000
0!
0%
b11 *
0-
02
b11 6
#337830000000
1!
1%
1-
12
15
#337840000000
0!
0%
b100 *
0-
02
b100 6
#337850000000
1!
1%
1-
12
#337860000000
0!
0%
b101 *
0-
02
b101 6
#337870000000
1!
1%
1-
12
#337880000000
0!
0%
b110 *
0-
02
b110 6
#337890000000
1!
1%
1-
12
#337900000000
0!
0%
b111 *
0-
02
b111 6
#337910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#337920000000
0!
0%
b0 *
0-
02
b0 6
#337930000000
1!
1%
1-
12
#337940000000
0!
0%
b1 *
0-
02
b1 6
#337950000000
1!
1%
1-
12
#337960000000
0!
0%
b10 *
0-
02
b10 6
#337970000000
1!
1%
1-
12
#337980000000
0!
0%
b11 *
0-
02
b11 6
#337990000000
1!
1%
1-
12
15
#338000000000
0!
0%
b100 *
0-
02
b100 6
#338010000000
1!
1%
1-
12
#338020000000
0!
0%
b101 *
0-
02
b101 6
#338030000000
1!
1%
1-
12
#338040000000
0!
0%
b110 *
0-
02
b110 6
#338050000000
1!
1%
1-
12
#338060000000
0!
0%
b111 *
0-
02
b111 6
#338070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#338080000000
0!
0%
b0 *
0-
02
b0 6
#338090000000
1!
1%
1-
12
#338100000000
0!
0%
b1 *
0-
02
b1 6
#338110000000
1!
1%
1-
12
#338120000000
0!
0%
b10 *
0-
02
b10 6
#338130000000
1!
1%
1-
12
#338140000000
0!
0%
b11 *
0-
02
b11 6
#338150000000
1!
1%
1-
12
15
#338160000000
0!
0%
b100 *
0-
02
b100 6
#338170000000
1!
1%
1-
12
#338180000000
0!
0%
b101 *
0-
02
b101 6
#338190000000
1!
1%
1-
12
#338200000000
0!
0%
b110 *
0-
02
b110 6
#338210000000
1!
1%
1-
12
#338220000000
0!
0%
b111 *
0-
02
b111 6
#338230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#338240000000
0!
0%
b0 *
0-
02
b0 6
#338250000000
1!
1%
1-
12
#338260000000
0!
0%
b1 *
0-
02
b1 6
#338270000000
1!
1%
1-
12
#338280000000
0!
0%
b10 *
0-
02
b10 6
#338290000000
1!
1%
1-
12
#338300000000
0!
0%
b11 *
0-
02
b11 6
#338310000000
1!
1%
1-
12
15
#338320000000
0!
0%
b100 *
0-
02
b100 6
#338330000000
1!
1%
1-
12
#338340000000
0!
0%
b101 *
0-
02
b101 6
#338350000000
1!
1%
1-
12
#338360000000
0!
0%
b110 *
0-
02
b110 6
#338370000000
1!
1%
1-
12
#338380000000
0!
0%
b111 *
0-
02
b111 6
#338390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#338400000000
0!
0%
b0 *
0-
02
b0 6
#338410000000
1!
1%
1-
12
#338420000000
0!
0%
b1 *
0-
02
b1 6
#338430000000
1!
1%
1-
12
#338440000000
0!
0%
b10 *
0-
02
b10 6
#338450000000
1!
1%
1-
12
#338460000000
0!
0%
b11 *
0-
02
b11 6
#338470000000
1!
1%
1-
12
15
#338480000000
0!
0%
b100 *
0-
02
b100 6
#338490000000
1!
1%
1-
12
#338500000000
0!
0%
b101 *
0-
02
b101 6
#338510000000
1!
1%
1-
12
#338520000000
0!
0%
b110 *
0-
02
b110 6
#338530000000
1!
1%
1-
12
#338540000000
0!
0%
b111 *
0-
02
b111 6
#338550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#338560000000
0!
0%
b0 *
0-
02
b0 6
#338570000000
1!
1%
1-
12
#338580000000
0!
0%
b1 *
0-
02
b1 6
#338590000000
1!
1%
1-
12
#338600000000
0!
0%
b10 *
0-
02
b10 6
#338610000000
1!
1%
1-
12
#338620000000
0!
0%
b11 *
0-
02
b11 6
#338630000000
1!
1%
1-
12
15
#338640000000
0!
0%
b100 *
0-
02
b100 6
#338650000000
1!
1%
1-
12
#338660000000
0!
0%
b101 *
0-
02
b101 6
#338670000000
1!
1%
1-
12
#338680000000
0!
0%
b110 *
0-
02
b110 6
#338690000000
1!
1%
1-
12
#338700000000
0!
0%
b111 *
0-
02
b111 6
#338710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#338720000000
0!
0%
b0 *
0-
02
b0 6
#338730000000
1!
1%
1-
12
#338740000000
0!
0%
b1 *
0-
02
b1 6
#338750000000
1!
1%
1-
12
#338760000000
0!
0%
b10 *
0-
02
b10 6
#338770000000
1!
1%
1-
12
#338780000000
0!
0%
b11 *
0-
02
b11 6
#338790000000
1!
1%
1-
12
15
#338800000000
0!
0%
b100 *
0-
02
b100 6
#338810000000
1!
1%
1-
12
#338820000000
0!
0%
b101 *
0-
02
b101 6
#338830000000
1!
1%
1-
12
#338840000000
0!
0%
b110 *
0-
02
b110 6
#338850000000
1!
1%
1-
12
#338860000000
0!
0%
b111 *
0-
02
b111 6
#338870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#338880000000
0!
0%
b0 *
0-
02
b0 6
#338890000000
1!
1%
1-
12
#338900000000
0!
0%
b1 *
0-
02
b1 6
#338910000000
1!
1%
1-
12
#338920000000
0!
0%
b10 *
0-
02
b10 6
#338930000000
1!
1%
1-
12
#338940000000
0!
0%
b11 *
0-
02
b11 6
#338950000000
1!
1%
1-
12
15
#338960000000
0!
0%
b100 *
0-
02
b100 6
#338970000000
1!
1%
1-
12
#338980000000
0!
0%
b101 *
0-
02
b101 6
#338990000000
1!
1%
1-
12
#339000000000
0!
0%
b110 *
0-
02
b110 6
#339010000000
1!
1%
1-
12
#339020000000
0!
0%
b111 *
0-
02
b111 6
#339030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#339040000000
0!
0%
b0 *
0-
02
b0 6
#339050000000
1!
1%
1-
12
#339060000000
0!
0%
b1 *
0-
02
b1 6
#339070000000
1!
1%
1-
12
#339080000000
0!
0%
b10 *
0-
02
b10 6
#339090000000
1!
1%
1-
12
#339100000000
0!
0%
b11 *
0-
02
b11 6
#339110000000
1!
1%
1-
12
15
#339120000000
0!
0%
b100 *
0-
02
b100 6
#339130000000
1!
1%
1-
12
#339140000000
0!
0%
b101 *
0-
02
b101 6
#339150000000
1!
1%
1-
12
#339160000000
0!
0%
b110 *
0-
02
b110 6
#339170000000
1!
1%
1-
12
#339180000000
0!
0%
b111 *
0-
02
b111 6
#339190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#339200000000
0!
0%
b0 *
0-
02
b0 6
#339210000000
1!
1%
1-
12
#339220000000
0!
0%
b1 *
0-
02
b1 6
#339230000000
1!
1%
1-
12
#339240000000
0!
0%
b10 *
0-
02
b10 6
#339250000000
1!
1%
1-
12
#339260000000
0!
0%
b11 *
0-
02
b11 6
#339270000000
1!
1%
1-
12
15
#339280000000
0!
0%
b100 *
0-
02
b100 6
#339290000000
1!
1%
1-
12
#339300000000
0!
0%
b101 *
0-
02
b101 6
#339310000000
1!
1%
1-
12
#339320000000
0!
0%
b110 *
0-
02
b110 6
#339330000000
1!
1%
1-
12
#339340000000
0!
0%
b111 *
0-
02
b111 6
#339350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#339360000000
0!
0%
b0 *
0-
02
b0 6
#339370000000
1!
1%
1-
12
#339380000000
0!
0%
b1 *
0-
02
b1 6
#339390000000
1!
1%
1-
12
#339400000000
0!
0%
b10 *
0-
02
b10 6
#339410000000
1!
1%
1-
12
#339420000000
0!
0%
b11 *
0-
02
b11 6
#339430000000
1!
1%
1-
12
15
#339440000000
0!
0%
b100 *
0-
02
b100 6
#339450000000
1!
1%
1-
12
#339460000000
0!
0%
b101 *
0-
02
b101 6
#339470000000
1!
1%
1-
12
#339480000000
0!
0%
b110 *
0-
02
b110 6
#339490000000
1!
1%
1-
12
#339500000000
0!
0%
b111 *
0-
02
b111 6
#339510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#339520000000
0!
0%
b0 *
0-
02
b0 6
#339530000000
1!
1%
1-
12
#339540000000
0!
0%
b1 *
0-
02
b1 6
#339550000000
1!
1%
1-
12
#339560000000
0!
0%
b10 *
0-
02
b10 6
#339570000000
1!
1%
1-
12
#339580000000
0!
0%
b11 *
0-
02
b11 6
#339590000000
1!
1%
1-
12
15
#339600000000
0!
0%
b100 *
0-
02
b100 6
#339610000000
1!
1%
1-
12
#339620000000
0!
0%
b101 *
0-
02
b101 6
#339630000000
1!
1%
1-
12
#339640000000
0!
0%
b110 *
0-
02
b110 6
#339650000000
1!
1%
1-
12
#339660000000
0!
0%
b111 *
0-
02
b111 6
#339670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#339680000000
0!
0%
b0 *
0-
02
b0 6
#339690000000
1!
1%
1-
12
#339700000000
0!
0%
b1 *
0-
02
b1 6
#339710000000
1!
1%
1-
12
#339720000000
0!
0%
b10 *
0-
02
b10 6
#339730000000
1!
1%
1-
12
#339740000000
0!
0%
b11 *
0-
02
b11 6
#339750000000
1!
1%
1-
12
15
#339760000000
0!
0%
b100 *
0-
02
b100 6
#339770000000
1!
1%
1-
12
#339780000000
0!
0%
b101 *
0-
02
b101 6
#339790000000
1!
1%
1-
12
#339800000000
0!
0%
b110 *
0-
02
b110 6
#339810000000
1!
1%
1-
12
#339820000000
0!
0%
b111 *
0-
02
b111 6
#339830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#339840000000
0!
0%
b0 *
0-
02
b0 6
#339850000000
1!
1%
1-
12
#339860000000
0!
0%
b1 *
0-
02
b1 6
#339870000000
1!
1%
1-
12
#339880000000
0!
0%
b10 *
0-
02
b10 6
#339890000000
1!
1%
1-
12
#339900000000
0!
0%
b11 *
0-
02
b11 6
#339910000000
1!
1%
1-
12
15
#339920000000
0!
0%
b100 *
0-
02
b100 6
#339930000000
1!
1%
1-
12
#339940000000
0!
0%
b101 *
0-
02
b101 6
#339950000000
1!
1%
1-
12
#339960000000
0!
0%
b110 *
0-
02
b110 6
#339970000000
1!
1%
1-
12
#339980000000
0!
0%
b111 *
0-
02
b111 6
#339990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#340000000000
0!
0%
b0 *
0-
02
b0 6
#340010000000
1!
1%
1-
12
#340020000000
0!
0%
b1 *
0-
02
b1 6
#340030000000
1!
1%
1-
12
#340040000000
0!
0%
b10 *
0-
02
b10 6
#340050000000
1!
1%
1-
12
#340060000000
0!
0%
b11 *
0-
02
b11 6
#340070000000
1!
1%
1-
12
15
#340080000000
0!
0%
b100 *
0-
02
b100 6
#340090000000
1!
1%
1-
12
#340100000000
0!
0%
b101 *
0-
02
b101 6
#340110000000
1!
1%
1-
12
#340120000000
0!
0%
b110 *
0-
02
b110 6
#340130000000
1!
1%
1-
12
#340140000000
0!
0%
b111 *
0-
02
b111 6
#340150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#340160000000
0!
0%
b0 *
0-
02
b0 6
#340170000000
1!
1%
1-
12
#340180000000
0!
0%
b1 *
0-
02
b1 6
#340190000000
1!
1%
1-
12
#340200000000
0!
0%
b10 *
0-
02
b10 6
#340210000000
1!
1%
1-
12
#340220000000
0!
0%
b11 *
0-
02
b11 6
#340230000000
1!
1%
1-
12
15
#340240000000
0!
0%
b100 *
0-
02
b100 6
#340250000000
1!
1%
1-
12
#340260000000
0!
0%
b101 *
0-
02
b101 6
#340270000000
1!
1%
1-
12
#340280000000
0!
0%
b110 *
0-
02
b110 6
#340290000000
1!
1%
1-
12
#340300000000
0!
0%
b111 *
0-
02
b111 6
#340310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#340320000000
0!
0%
b0 *
0-
02
b0 6
#340330000000
1!
1%
1-
12
#340340000000
0!
0%
b1 *
0-
02
b1 6
#340350000000
1!
1%
1-
12
#340360000000
0!
0%
b10 *
0-
02
b10 6
#340370000000
1!
1%
1-
12
#340380000000
0!
0%
b11 *
0-
02
b11 6
#340390000000
1!
1%
1-
12
15
#340400000000
0!
0%
b100 *
0-
02
b100 6
#340410000000
1!
1%
1-
12
#340420000000
0!
0%
b101 *
0-
02
b101 6
#340430000000
1!
1%
1-
12
#340440000000
0!
0%
b110 *
0-
02
b110 6
#340450000000
1!
1%
1-
12
#340460000000
0!
0%
b111 *
0-
02
b111 6
#340470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#340480000000
0!
0%
b0 *
0-
02
b0 6
#340490000000
1!
1%
1-
12
#340500000000
0!
0%
b1 *
0-
02
b1 6
#340510000000
1!
1%
1-
12
#340520000000
0!
0%
b10 *
0-
02
b10 6
#340530000000
1!
1%
1-
12
#340540000000
0!
0%
b11 *
0-
02
b11 6
#340550000000
1!
1%
1-
12
15
#340560000000
0!
0%
b100 *
0-
02
b100 6
#340570000000
1!
1%
1-
12
#340580000000
0!
0%
b101 *
0-
02
b101 6
#340590000000
1!
1%
1-
12
#340600000000
0!
0%
b110 *
0-
02
b110 6
#340610000000
1!
1%
1-
12
#340620000000
0!
0%
b111 *
0-
02
b111 6
#340630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#340640000000
0!
0%
b0 *
0-
02
b0 6
#340650000000
1!
1%
1-
12
#340660000000
0!
0%
b1 *
0-
02
b1 6
#340670000000
1!
1%
1-
12
#340680000000
0!
0%
b10 *
0-
02
b10 6
#340690000000
1!
1%
1-
12
#340700000000
0!
0%
b11 *
0-
02
b11 6
#340710000000
1!
1%
1-
12
15
#340720000000
0!
0%
b100 *
0-
02
b100 6
#340730000000
1!
1%
1-
12
#340740000000
0!
0%
b101 *
0-
02
b101 6
#340750000000
1!
1%
1-
12
#340760000000
0!
0%
b110 *
0-
02
b110 6
#340770000000
1!
1%
1-
12
#340780000000
0!
0%
b111 *
0-
02
b111 6
#340790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#340800000000
0!
0%
b0 *
0-
02
b0 6
#340810000000
1!
1%
1-
12
#340820000000
0!
0%
b1 *
0-
02
b1 6
#340830000000
1!
1%
1-
12
#340840000000
0!
0%
b10 *
0-
02
b10 6
#340850000000
1!
1%
1-
12
#340860000000
0!
0%
b11 *
0-
02
b11 6
#340870000000
1!
1%
1-
12
15
#340880000000
0!
0%
b100 *
0-
02
b100 6
#340890000000
1!
1%
1-
12
#340900000000
0!
0%
b101 *
0-
02
b101 6
#340910000000
1!
1%
1-
12
#340920000000
0!
0%
b110 *
0-
02
b110 6
#340930000000
1!
1%
1-
12
#340940000000
0!
0%
b111 *
0-
02
b111 6
#340950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#340960000000
0!
0%
b0 *
0-
02
b0 6
#340970000000
1!
1%
1-
12
#340980000000
0!
0%
b1 *
0-
02
b1 6
#340990000000
1!
1%
1-
12
#341000000000
0!
0%
b10 *
0-
02
b10 6
#341010000000
1!
1%
1-
12
#341020000000
0!
0%
b11 *
0-
02
b11 6
#341030000000
1!
1%
1-
12
15
#341040000000
0!
0%
b100 *
0-
02
b100 6
#341050000000
1!
1%
1-
12
#341060000000
0!
0%
b101 *
0-
02
b101 6
#341070000000
1!
1%
1-
12
#341080000000
0!
0%
b110 *
0-
02
b110 6
#341090000000
1!
1%
1-
12
#341100000000
0!
0%
b111 *
0-
02
b111 6
#341110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#341120000000
0!
0%
b0 *
0-
02
b0 6
#341130000000
1!
1%
1-
12
#341140000000
0!
0%
b1 *
0-
02
b1 6
#341150000000
1!
1%
1-
12
#341160000000
0!
0%
b10 *
0-
02
b10 6
#341170000000
1!
1%
1-
12
#341180000000
0!
0%
b11 *
0-
02
b11 6
#341190000000
1!
1%
1-
12
15
#341200000000
0!
0%
b100 *
0-
02
b100 6
#341210000000
1!
1%
1-
12
#341220000000
0!
0%
b101 *
0-
02
b101 6
#341230000000
1!
1%
1-
12
#341240000000
0!
0%
b110 *
0-
02
b110 6
#341250000000
1!
1%
1-
12
#341260000000
0!
0%
b111 *
0-
02
b111 6
#341270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#341280000000
0!
0%
b0 *
0-
02
b0 6
#341290000000
1!
1%
1-
12
#341300000000
0!
0%
b1 *
0-
02
b1 6
#341310000000
1!
1%
1-
12
#341320000000
0!
0%
b10 *
0-
02
b10 6
#341330000000
1!
1%
1-
12
#341340000000
0!
0%
b11 *
0-
02
b11 6
#341350000000
1!
1%
1-
12
15
#341360000000
0!
0%
b100 *
0-
02
b100 6
#341370000000
1!
1%
1-
12
#341380000000
0!
0%
b101 *
0-
02
b101 6
#341390000000
1!
1%
1-
12
#341400000000
0!
0%
b110 *
0-
02
b110 6
#341410000000
1!
1%
1-
12
#341420000000
0!
0%
b111 *
0-
02
b111 6
#341430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#341440000000
0!
0%
b0 *
0-
02
b0 6
#341450000000
1!
1%
1-
12
#341460000000
0!
0%
b1 *
0-
02
b1 6
#341470000000
1!
1%
1-
12
#341480000000
0!
0%
b10 *
0-
02
b10 6
#341490000000
1!
1%
1-
12
#341500000000
0!
0%
b11 *
0-
02
b11 6
#341510000000
1!
1%
1-
12
15
#341520000000
0!
0%
b100 *
0-
02
b100 6
#341530000000
1!
1%
1-
12
#341540000000
0!
0%
b101 *
0-
02
b101 6
#341550000000
1!
1%
1-
12
#341560000000
0!
0%
b110 *
0-
02
b110 6
#341570000000
1!
1%
1-
12
#341580000000
0!
0%
b111 *
0-
02
b111 6
#341590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#341600000000
0!
0%
b0 *
0-
02
b0 6
#341610000000
1!
1%
1-
12
#341620000000
0!
0%
b1 *
0-
02
b1 6
#341630000000
1!
1%
1-
12
#341640000000
0!
0%
b10 *
0-
02
b10 6
#341650000000
1!
1%
1-
12
#341660000000
0!
0%
b11 *
0-
02
b11 6
#341670000000
1!
1%
1-
12
15
#341680000000
0!
0%
b100 *
0-
02
b100 6
#341690000000
1!
1%
1-
12
#341700000000
0!
0%
b101 *
0-
02
b101 6
#341710000000
1!
1%
1-
12
#341720000000
0!
0%
b110 *
0-
02
b110 6
#341730000000
1!
1%
1-
12
#341740000000
0!
0%
b111 *
0-
02
b111 6
#341750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#341760000000
0!
0%
b0 *
0-
02
b0 6
#341770000000
1!
1%
1-
12
#341780000000
0!
0%
b1 *
0-
02
b1 6
#341790000000
1!
1%
1-
12
#341800000000
0!
0%
b10 *
0-
02
b10 6
#341810000000
1!
1%
1-
12
#341820000000
0!
0%
b11 *
0-
02
b11 6
#341830000000
1!
1%
1-
12
15
#341840000000
0!
0%
b100 *
0-
02
b100 6
#341850000000
1!
1%
1-
12
#341860000000
0!
0%
b101 *
0-
02
b101 6
#341870000000
1!
1%
1-
12
#341880000000
0!
0%
b110 *
0-
02
b110 6
#341890000000
1!
1%
1-
12
#341900000000
0!
0%
b111 *
0-
02
b111 6
#341910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#341920000000
0!
0%
b0 *
0-
02
b0 6
#341930000000
1!
1%
1-
12
#341940000000
0!
0%
b1 *
0-
02
b1 6
#341950000000
1!
1%
1-
12
#341960000000
0!
0%
b10 *
0-
02
b10 6
#341970000000
1!
1%
1-
12
#341980000000
0!
0%
b11 *
0-
02
b11 6
#341990000000
1!
1%
1-
12
15
#342000000000
0!
0%
b100 *
0-
02
b100 6
#342010000000
1!
1%
1-
12
#342020000000
0!
0%
b101 *
0-
02
b101 6
#342030000000
1!
1%
1-
12
#342040000000
0!
0%
b110 *
0-
02
b110 6
#342050000000
1!
1%
1-
12
#342060000000
0!
0%
b111 *
0-
02
b111 6
#342070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#342080000000
0!
0%
b0 *
0-
02
b0 6
#342090000000
1!
1%
1-
12
#342100000000
0!
0%
b1 *
0-
02
b1 6
#342110000000
1!
1%
1-
12
#342120000000
0!
0%
b10 *
0-
02
b10 6
#342130000000
1!
1%
1-
12
#342140000000
0!
0%
b11 *
0-
02
b11 6
#342150000000
1!
1%
1-
12
15
#342160000000
0!
0%
b100 *
0-
02
b100 6
#342170000000
1!
1%
1-
12
#342180000000
0!
0%
b101 *
0-
02
b101 6
#342190000000
1!
1%
1-
12
#342200000000
0!
0%
b110 *
0-
02
b110 6
#342210000000
1!
1%
1-
12
#342220000000
0!
0%
b111 *
0-
02
b111 6
#342230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#342240000000
0!
0%
b0 *
0-
02
b0 6
#342250000000
1!
1%
1-
12
#342260000000
0!
0%
b1 *
0-
02
b1 6
#342270000000
1!
1%
1-
12
#342280000000
0!
0%
b10 *
0-
02
b10 6
#342290000000
1!
1%
1-
12
#342300000000
0!
0%
b11 *
0-
02
b11 6
#342310000000
1!
1%
1-
12
15
#342320000000
0!
0%
b100 *
0-
02
b100 6
#342330000000
1!
1%
1-
12
#342340000000
0!
0%
b101 *
0-
02
b101 6
#342350000000
1!
1%
1-
12
#342360000000
0!
0%
b110 *
0-
02
b110 6
#342370000000
1!
1%
1-
12
#342380000000
0!
0%
b111 *
0-
02
b111 6
#342390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#342400000000
0!
0%
b0 *
0-
02
b0 6
#342410000000
1!
1%
1-
12
#342420000000
0!
0%
b1 *
0-
02
b1 6
#342430000000
1!
1%
1-
12
#342440000000
0!
0%
b10 *
0-
02
b10 6
#342450000000
1!
1%
1-
12
#342460000000
0!
0%
b11 *
0-
02
b11 6
#342470000000
1!
1%
1-
12
15
#342480000000
0!
0%
b100 *
0-
02
b100 6
#342490000000
1!
1%
1-
12
#342500000000
0!
0%
b101 *
0-
02
b101 6
#342510000000
1!
1%
1-
12
#342520000000
0!
0%
b110 *
0-
02
b110 6
#342530000000
1!
1%
1-
12
#342540000000
0!
0%
b111 *
0-
02
b111 6
#342550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#342560000000
0!
0%
b0 *
0-
02
b0 6
#342570000000
1!
1%
1-
12
#342580000000
0!
0%
b1 *
0-
02
b1 6
#342590000000
1!
1%
1-
12
#342600000000
0!
0%
b10 *
0-
02
b10 6
#342610000000
1!
1%
1-
12
#342620000000
0!
0%
b11 *
0-
02
b11 6
#342630000000
1!
1%
1-
12
15
#342640000000
0!
0%
b100 *
0-
02
b100 6
#342650000000
1!
1%
1-
12
#342660000000
0!
0%
b101 *
0-
02
b101 6
#342670000000
1!
1%
1-
12
#342680000000
0!
0%
b110 *
0-
02
b110 6
#342690000000
1!
1%
1-
12
#342700000000
0!
0%
b111 *
0-
02
b111 6
#342710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#342720000000
0!
0%
b0 *
0-
02
b0 6
#342730000000
1!
1%
1-
12
#342740000000
0!
0%
b1 *
0-
02
b1 6
#342750000000
1!
1%
1-
12
#342760000000
0!
0%
b10 *
0-
02
b10 6
#342770000000
1!
1%
1-
12
#342780000000
0!
0%
b11 *
0-
02
b11 6
#342790000000
1!
1%
1-
12
15
#342800000000
0!
0%
b100 *
0-
02
b100 6
#342810000000
1!
1%
1-
12
#342820000000
0!
0%
b101 *
0-
02
b101 6
#342830000000
1!
1%
1-
12
#342840000000
0!
0%
b110 *
0-
02
b110 6
#342850000000
1!
1%
1-
12
#342860000000
0!
0%
b111 *
0-
02
b111 6
#342870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#342880000000
0!
0%
b0 *
0-
02
b0 6
#342890000000
1!
1%
1-
12
#342900000000
0!
0%
b1 *
0-
02
b1 6
#342910000000
1!
1%
1-
12
#342920000000
0!
0%
b10 *
0-
02
b10 6
#342930000000
1!
1%
1-
12
#342940000000
0!
0%
b11 *
0-
02
b11 6
#342950000000
1!
1%
1-
12
15
#342960000000
0!
0%
b100 *
0-
02
b100 6
#342970000000
1!
1%
1-
12
#342980000000
0!
0%
b101 *
0-
02
b101 6
#342990000000
1!
1%
1-
12
#343000000000
0!
0%
b110 *
0-
02
b110 6
#343010000000
1!
1%
1-
12
#343020000000
0!
0%
b111 *
0-
02
b111 6
#343030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#343040000000
0!
0%
b0 *
0-
02
b0 6
#343050000000
1!
1%
1-
12
#343060000000
0!
0%
b1 *
0-
02
b1 6
#343070000000
1!
1%
1-
12
#343080000000
0!
0%
b10 *
0-
02
b10 6
#343090000000
1!
1%
1-
12
#343100000000
0!
0%
b11 *
0-
02
b11 6
#343110000000
1!
1%
1-
12
15
#343120000000
0!
0%
b100 *
0-
02
b100 6
#343130000000
1!
1%
1-
12
#343140000000
0!
0%
b101 *
0-
02
b101 6
#343150000000
1!
1%
1-
12
#343160000000
0!
0%
b110 *
0-
02
b110 6
#343170000000
1!
1%
1-
12
#343180000000
0!
0%
b111 *
0-
02
b111 6
#343190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#343200000000
0!
0%
b0 *
0-
02
b0 6
#343210000000
1!
1%
1-
12
#343220000000
0!
0%
b1 *
0-
02
b1 6
#343230000000
1!
1%
1-
12
#343240000000
0!
0%
b10 *
0-
02
b10 6
#343250000000
1!
1%
1-
12
#343260000000
0!
0%
b11 *
0-
02
b11 6
#343270000000
1!
1%
1-
12
15
#343280000000
0!
0%
b100 *
0-
02
b100 6
#343290000000
1!
1%
1-
12
#343300000000
0!
0%
b101 *
0-
02
b101 6
#343310000000
1!
1%
1-
12
#343320000000
0!
0%
b110 *
0-
02
b110 6
#343330000000
1!
1%
1-
12
#343340000000
0!
0%
b111 *
0-
02
b111 6
#343350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#343360000000
0!
0%
b0 *
0-
02
b0 6
#343370000000
1!
1%
1-
12
#343380000000
0!
0%
b1 *
0-
02
b1 6
#343390000000
1!
1%
1-
12
#343400000000
0!
0%
b10 *
0-
02
b10 6
#343410000000
1!
1%
1-
12
#343420000000
0!
0%
b11 *
0-
02
b11 6
#343430000000
1!
1%
1-
12
15
#343440000000
0!
0%
b100 *
0-
02
b100 6
#343450000000
1!
1%
1-
12
#343460000000
0!
0%
b101 *
0-
02
b101 6
#343470000000
1!
1%
1-
12
#343480000000
0!
0%
b110 *
0-
02
b110 6
#343490000000
1!
1%
1-
12
#343500000000
0!
0%
b111 *
0-
02
b111 6
#343510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#343520000000
0!
0%
b0 *
0-
02
b0 6
#343530000000
1!
1%
1-
12
#343540000000
0!
0%
b1 *
0-
02
b1 6
#343550000000
1!
1%
1-
12
#343560000000
0!
0%
b10 *
0-
02
b10 6
#343570000000
1!
1%
1-
12
#343580000000
0!
0%
b11 *
0-
02
b11 6
#343590000000
1!
1%
1-
12
15
#343600000000
0!
0%
b100 *
0-
02
b100 6
#343610000000
1!
1%
1-
12
#343620000000
0!
0%
b101 *
0-
02
b101 6
#343630000000
1!
1%
1-
12
#343640000000
0!
0%
b110 *
0-
02
b110 6
#343650000000
1!
1%
1-
12
#343660000000
0!
0%
b111 *
0-
02
b111 6
#343670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#343680000000
0!
0%
b0 *
0-
02
b0 6
#343690000000
1!
1%
1-
12
#343700000000
0!
0%
b1 *
0-
02
b1 6
#343710000000
1!
1%
1-
12
#343720000000
0!
0%
b10 *
0-
02
b10 6
#343730000000
1!
1%
1-
12
#343740000000
0!
0%
b11 *
0-
02
b11 6
#343750000000
1!
1%
1-
12
15
#343760000000
0!
0%
b100 *
0-
02
b100 6
#343770000000
1!
1%
1-
12
#343780000000
0!
0%
b101 *
0-
02
b101 6
#343790000000
1!
1%
1-
12
#343800000000
0!
0%
b110 *
0-
02
b110 6
#343810000000
1!
1%
1-
12
#343820000000
0!
0%
b111 *
0-
02
b111 6
#343830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#343840000000
0!
0%
b0 *
0-
02
b0 6
#343850000000
1!
1%
1-
12
#343860000000
0!
0%
b1 *
0-
02
b1 6
#343870000000
1!
1%
1-
12
#343880000000
0!
0%
b10 *
0-
02
b10 6
#343890000000
1!
1%
1-
12
#343900000000
0!
0%
b11 *
0-
02
b11 6
#343910000000
1!
1%
1-
12
15
#343920000000
0!
0%
b100 *
0-
02
b100 6
#343930000000
1!
1%
1-
12
#343940000000
0!
0%
b101 *
0-
02
b101 6
#343950000000
1!
1%
1-
12
#343960000000
0!
0%
b110 *
0-
02
b110 6
#343970000000
1!
1%
1-
12
#343980000000
0!
0%
b111 *
0-
02
b111 6
#343990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#344000000000
0!
0%
b0 *
0-
02
b0 6
#344010000000
1!
1%
1-
12
#344020000000
0!
0%
b1 *
0-
02
b1 6
#344030000000
1!
1%
1-
12
#344040000000
0!
0%
b10 *
0-
02
b10 6
#344050000000
1!
1%
1-
12
#344060000000
0!
0%
b11 *
0-
02
b11 6
#344070000000
1!
1%
1-
12
15
#344080000000
0!
0%
b100 *
0-
02
b100 6
#344090000000
1!
1%
1-
12
#344100000000
0!
0%
b101 *
0-
02
b101 6
#344110000000
1!
1%
1-
12
#344120000000
0!
0%
b110 *
0-
02
b110 6
#344130000000
1!
1%
1-
12
#344140000000
0!
0%
b111 *
0-
02
b111 6
#344150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#344160000000
0!
0%
b0 *
0-
02
b0 6
#344170000000
1!
1%
1-
12
#344180000000
0!
0%
b1 *
0-
02
b1 6
#344190000000
1!
1%
1-
12
#344200000000
0!
0%
b10 *
0-
02
b10 6
#344210000000
1!
1%
1-
12
#344220000000
0!
0%
b11 *
0-
02
b11 6
#344230000000
1!
1%
1-
12
15
#344240000000
0!
0%
b100 *
0-
02
b100 6
#344250000000
1!
1%
1-
12
#344260000000
0!
0%
b101 *
0-
02
b101 6
#344270000000
1!
1%
1-
12
#344280000000
0!
0%
b110 *
0-
02
b110 6
#344290000000
1!
1%
1-
12
#344300000000
0!
0%
b111 *
0-
02
b111 6
#344310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#344320000000
0!
0%
b0 *
0-
02
b0 6
#344330000000
1!
1%
1-
12
#344340000000
0!
0%
b1 *
0-
02
b1 6
#344350000000
1!
1%
1-
12
#344360000000
0!
0%
b10 *
0-
02
b10 6
#344370000000
1!
1%
1-
12
#344380000000
0!
0%
b11 *
0-
02
b11 6
#344390000000
1!
1%
1-
12
15
#344400000000
0!
0%
b100 *
0-
02
b100 6
#344410000000
1!
1%
1-
12
#344420000000
0!
0%
b101 *
0-
02
b101 6
#344430000000
1!
1%
1-
12
#344440000000
0!
0%
b110 *
0-
02
b110 6
#344450000000
1!
1%
1-
12
#344460000000
0!
0%
b111 *
0-
02
b111 6
#344470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#344480000000
0!
0%
b0 *
0-
02
b0 6
#344490000000
1!
1%
1-
12
#344500000000
0!
0%
b1 *
0-
02
b1 6
#344510000000
1!
1%
1-
12
#344520000000
0!
0%
b10 *
0-
02
b10 6
#344530000000
1!
1%
1-
12
#344540000000
0!
0%
b11 *
0-
02
b11 6
#344550000000
1!
1%
1-
12
15
#344560000000
0!
0%
b100 *
0-
02
b100 6
#344570000000
1!
1%
1-
12
#344580000000
0!
0%
b101 *
0-
02
b101 6
#344590000000
1!
1%
1-
12
#344600000000
0!
0%
b110 *
0-
02
b110 6
#344610000000
1!
1%
1-
12
#344620000000
0!
0%
b111 *
0-
02
b111 6
#344630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#344640000000
0!
0%
b0 *
0-
02
b0 6
#344650000000
1!
1%
1-
12
#344660000000
0!
0%
b1 *
0-
02
b1 6
#344670000000
1!
1%
1-
12
#344680000000
0!
0%
b10 *
0-
02
b10 6
#344690000000
1!
1%
1-
12
#344700000000
0!
0%
b11 *
0-
02
b11 6
#344710000000
1!
1%
1-
12
15
#344720000000
0!
0%
b100 *
0-
02
b100 6
#344730000000
1!
1%
1-
12
#344740000000
0!
0%
b101 *
0-
02
b101 6
#344750000000
1!
1%
1-
12
#344760000000
0!
0%
b110 *
0-
02
b110 6
#344770000000
1!
1%
1-
12
#344780000000
0!
0%
b111 *
0-
02
b111 6
#344790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#344800000000
0!
0%
b0 *
0-
02
b0 6
#344810000000
1!
1%
1-
12
#344820000000
0!
0%
b1 *
0-
02
b1 6
#344830000000
1!
1%
1-
12
#344840000000
0!
0%
b10 *
0-
02
b10 6
#344850000000
1!
1%
1-
12
#344860000000
0!
0%
b11 *
0-
02
b11 6
#344870000000
1!
1%
1-
12
15
#344880000000
0!
0%
b100 *
0-
02
b100 6
#344890000000
1!
1%
1-
12
#344900000000
0!
0%
b101 *
0-
02
b101 6
#344910000000
1!
1%
1-
12
#344920000000
0!
0%
b110 *
0-
02
b110 6
#344930000000
1!
1%
1-
12
#344940000000
0!
0%
b111 *
0-
02
b111 6
#344950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#344960000000
0!
0%
b0 *
0-
02
b0 6
#344970000000
1!
1%
1-
12
#344980000000
0!
0%
b1 *
0-
02
b1 6
#344990000000
1!
1%
1-
12
#345000000000
0!
0%
b10 *
0-
02
b10 6
#345010000000
1!
1%
1-
12
#345020000000
0!
0%
b11 *
0-
02
b11 6
#345030000000
1!
1%
1-
12
15
#345040000000
0!
0%
b100 *
0-
02
b100 6
#345050000000
1!
1%
1-
12
#345060000000
0!
0%
b101 *
0-
02
b101 6
#345070000000
1!
1%
1-
12
#345080000000
0!
0%
b110 *
0-
02
b110 6
#345090000000
1!
1%
1-
12
#345100000000
0!
0%
b111 *
0-
02
b111 6
#345110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#345120000000
0!
0%
b0 *
0-
02
b0 6
#345130000000
1!
1%
1-
12
#345140000000
0!
0%
b1 *
0-
02
b1 6
#345150000000
1!
1%
1-
12
#345160000000
0!
0%
b10 *
0-
02
b10 6
#345170000000
1!
1%
1-
12
#345180000000
0!
0%
b11 *
0-
02
b11 6
#345190000000
1!
1%
1-
12
15
#345200000000
0!
0%
b100 *
0-
02
b100 6
#345210000000
1!
1%
1-
12
#345220000000
0!
0%
b101 *
0-
02
b101 6
#345230000000
1!
1%
1-
12
#345240000000
0!
0%
b110 *
0-
02
b110 6
#345250000000
1!
1%
1-
12
#345260000000
0!
0%
b111 *
0-
02
b111 6
#345270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#345280000000
0!
0%
b0 *
0-
02
b0 6
#345290000000
1!
1%
1-
12
#345300000000
0!
0%
b1 *
0-
02
b1 6
#345310000000
1!
1%
1-
12
#345320000000
0!
0%
b10 *
0-
02
b10 6
#345330000000
1!
1%
1-
12
#345340000000
0!
0%
b11 *
0-
02
b11 6
#345350000000
1!
1%
1-
12
15
#345360000000
0!
0%
b100 *
0-
02
b100 6
#345370000000
1!
1%
1-
12
#345380000000
0!
0%
b101 *
0-
02
b101 6
#345390000000
1!
1%
1-
12
#345400000000
0!
0%
b110 *
0-
02
b110 6
#345410000000
1!
1%
1-
12
#345420000000
0!
0%
b111 *
0-
02
b111 6
#345430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#345440000000
0!
0%
b0 *
0-
02
b0 6
#345450000000
1!
1%
1-
12
#345460000000
0!
0%
b1 *
0-
02
b1 6
#345470000000
1!
1%
1-
12
#345480000000
0!
0%
b10 *
0-
02
b10 6
#345490000000
1!
1%
1-
12
#345500000000
0!
0%
b11 *
0-
02
b11 6
#345510000000
1!
1%
1-
12
15
#345520000000
0!
0%
b100 *
0-
02
b100 6
#345530000000
1!
1%
1-
12
#345540000000
0!
0%
b101 *
0-
02
b101 6
#345550000000
1!
1%
1-
12
#345560000000
0!
0%
b110 *
0-
02
b110 6
#345570000000
1!
1%
1-
12
#345580000000
0!
0%
b111 *
0-
02
b111 6
#345590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#345600000000
0!
0%
b0 *
0-
02
b0 6
#345610000000
1!
1%
1-
12
#345620000000
0!
0%
b1 *
0-
02
b1 6
#345630000000
1!
1%
1-
12
#345640000000
0!
0%
b10 *
0-
02
b10 6
#345650000000
1!
1%
1-
12
#345660000000
0!
0%
b11 *
0-
02
b11 6
#345670000000
1!
1%
1-
12
15
#345680000000
0!
0%
b100 *
0-
02
b100 6
#345690000000
1!
1%
1-
12
#345700000000
0!
0%
b101 *
0-
02
b101 6
#345710000000
1!
1%
1-
12
#345720000000
0!
0%
b110 *
0-
02
b110 6
#345730000000
1!
1%
1-
12
#345740000000
0!
0%
b111 *
0-
02
b111 6
#345750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#345760000000
0!
0%
b0 *
0-
02
b0 6
#345770000000
1!
1%
1-
12
#345780000000
0!
0%
b1 *
0-
02
b1 6
#345790000000
1!
1%
1-
12
#345800000000
0!
0%
b10 *
0-
02
b10 6
#345810000000
1!
1%
1-
12
#345820000000
0!
0%
b11 *
0-
02
b11 6
#345830000000
1!
1%
1-
12
15
#345840000000
0!
0%
b100 *
0-
02
b100 6
#345850000000
1!
1%
1-
12
#345860000000
0!
0%
b101 *
0-
02
b101 6
#345870000000
1!
1%
1-
12
#345880000000
0!
0%
b110 *
0-
02
b110 6
#345890000000
1!
1%
1-
12
#345900000000
0!
0%
b111 *
0-
02
b111 6
#345910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#345920000000
0!
0%
b0 *
0-
02
b0 6
#345930000000
1!
1%
1-
12
#345940000000
0!
0%
b1 *
0-
02
b1 6
#345950000000
1!
1%
1-
12
#345960000000
0!
0%
b10 *
0-
02
b10 6
#345970000000
1!
1%
1-
12
#345980000000
0!
0%
b11 *
0-
02
b11 6
#345990000000
1!
1%
1-
12
15
#346000000000
0!
0%
b100 *
0-
02
b100 6
#346010000000
1!
1%
1-
12
#346020000000
0!
0%
b101 *
0-
02
b101 6
#346030000000
1!
1%
1-
12
#346040000000
0!
0%
b110 *
0-
02
b110 6
#346050000000
1!
1%
1-
12
#346060000000
0!
0%
b111 *
0-
02
b111 6
#346070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#346080000000
0!
0%
b0 *
0-
02
b0 6
#346090000000
1!
1%
1-
12
#346100000000
0!
0%
b1 *
0-
02
b1 6
#346110000000
1!
1%
1-
12
#346120000000
0!
0%
b10 *
0-
02
b10 6
#346130000000
1!
1%
1-
12
#346140000000
0!
0%
b11 *
0-
02
b11 6
#346150000000
1!
1%
1-
12
15
#346160000000
0!
0%
b100 *
0-
02
b100 6
#346170000000
1!
1%
1-
12
#346180000000
0!
0%
b101 *
0-
02
b101 6
#346190000000
1!
1%
1-
12
#346200000000
0!
0%
b110 *
0-
02
b110 6
#346210000000
1!
1%
1-
12
#346220000000
0!
0%
b111 *
0-
02
b111 6
#346230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#346240000000
0!
0%
b0 *
0-
02
b0 6
#346250000000
1!
1%
1-
12
#346260000000
0!
0%
b1 *
0-
02
b1 6
#346270000000
1!
1%
1-
12
#346280000000
0!
0%
b10 *
0-
02
b10 6
#346290000000
1!
1%
1-
12
#346300000000
0!
0%
b11 *
0-
02
b11 6
#346310000000
1!
1%
1-
12
15
#346320000000
0!
0%
b100 *
0-
02
b100 6
#346330000000
1!
1%
1-
12
#346340000000
0!
0%
b101 *
0-
02
b101 6
#346350000000
1!
1%
1-
12
#346360000000
0!
0%
b110 *
0-
02
b110 6
#346370000000
1!
1%
1-
12
#346380000000
0!
0%
b111 *
0-
02
b111 6
#346390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#346400000000
0!
0%
b0 *
0-
02
b0 6
#346410000000
1!
1%
1-
12
#346420000000
0!
0%
b1 *
0-
02
b1 6
#346430000000
1!
1%
1-
12
#346440000000
0!
0%
b10 *
0-
02
b10 6
#346450000000
1!
1%
1-
12
#346460000000
0!
0%
b11 *
0-
02
b11 6
#346470000000
1!
1%
1-
12
15
#346480000000
0!
0%
b100 *
0-
02
b100 6
#346490000000
1!
1%
1-
12
#346500000000
0!
0%
b101 *
0-
02
b101 6
#346510000000
1!
1%
1-
12
#346520000000
0!
0%
b110 *
0-
02
b110 6
#346530000000
1!
1%
1-
12
#346540000000
0!
0%
b111 *
0-
02
b111 6
#346550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#346560000000
0!
0%
b0 *
0-
02
b0 6
#346570000000
1!
1%
1-
12
#346580000000
0!
0%
b1 *
0-
02
b1 6
#346590000000
1!
1%
1-
12
#346600000000
0!
0%
b10 *
0-
02
b10 6
#346610000000
1!
1%
1-
12
#346620000000
0!
0%
b11 *
0-
02
b11 6
#346630000000
1!
1%
1-
12
15
#346640000000
0!
0%
b100 *
0-
02
b100 6
#346650000000
1!
1%
1-
12
#346660000000
0!
0%
b101 *
0-
02
b101 6
#346670000000
1!
1%
1-
12
#346680000000
0!
0%
b110 *
0-
02
b110 6
#346690000000
1!
1%
1-
12
#346700000000
0!
0%
b111 *
0-
02
b111 6
#346710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#346720000000
0!
0%
b0 *
0-
02
b0 6
#346730000000
1!
1%
1-
12
#346740000000
0!
0%
b1 *
0-
02
b1 6
#346750000000
1!
1%
1-
12
#346760000000
0!
0%
b10 *
0-
02
b10 6
#346770000000
1!
1%
1-
12
#346780000000
0!
0%
b11 *
0-
02
b11 6
#346790000000
1!
1%
1-
12
15
#346800000000
0!
0%
b100 *
0-
02
b100 6
#346810000000
1!
1%
1-
12
#346820000000
0!
0%
b101 *
0-
02
b101 6
#346830000000
1!
1%
1-
12
#346840000000
0!
0%
b110 *
0-
02
b110 6
#346850000000
1!
1%
1-
12
#346860000000
0!
0%
b111 *
0-
02
b111 6
#346870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#346880000000
0!
0%
b0 *
0-
02
b0 6
#346890000000
1!
1%
1-
12
#346900000000
0!
0%
b1 *
0-
02
b1 6
#346910000000
1!
1%
1-
12
#346920000000
0!
0%
b10 *
0-
02
b10 6
#346930000000
1!
1%
1-
12
#346940000000
0!
0%
b11 *
0-
02
b11 6
#346950000000
1!
1%
1-
12
15
#346960000000
0!
0%
b100 *
0-
02
b100 6
#346970000000
1!
1%
1-
12
#346980000000
0!
0%
b101 *
0-
02
b101 6
#346990000000
1!
1%
1-
12
#347000000000
0!
0%
b110 *
0-
02
b110 6
#347010000000
1!
1%
1-
12
#347020000000
0!
0%
b111 *
0-
02
b111 6
#347030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#347040000000
0!
0%
b0 *
0-
02
b0 6
#347050000000
1!
1%
1-
12
#347060000000
0!
0%
b1 *
0-
02
b1 6
#347070000000
1!
1%
1-
12
#347080000000
0!
0%
b10 *
0-
02
b10 6
#347090000000
1!
1%
1-
12
#347100000000
0!
0%
b11 *
0-
02
b11 6
#347110000000
1!
1%
1-
12
15
#347120000000
0!
0%
b100 *
0-
02
b100 6
#347130000000
1!
1%
1-
12
#347140000000
0!
0%
b101 *
0-
02
b101 6
#347150000000
1!
1%
1-
12
#347160000000
0!
0%
b110 *
0-
02
b110 6
#347170000000
1!
1%
1-
12
#347180000000
0!
0%
b111 *
0-
02
b111 6
#347190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#347200000000
0!
0%
b0 *
0-
02
b0 6
#347210000000
1!
1%
1-
12
#347220000000
0!
0%
b1 *
0-
02
b1 6
#347230000000
1!
1%
1-
12
#347240000000
0!
0%
b10 *
0-
02
b10 6
#347250000000
1!
1%
1-
12
#347260000000
0!
0%
b11 *
0-
02
b11 6
#347270000000
1!
1%
1-
12
15
#347280000000
0!
0%
b100 *
0-
02
b100 6
#347290000000
1!
1%
1-
12
#347300000000
0!
0%
b101 *
0-
02
b101 6
#347310000000
1!
1%
1-
12
#347320000000
0!
0%
b110 *
0-
02
b110 6
#347330000000
1!
1%
1-
12
#347340000000
0!
0%
b111 *
0-
02
b111 6
#347350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#347360000000
0!
0%
b0 *
0-
02
b0 6
#347370000000
1!
1%
1-
12
#347380000000
0!
0%
b1 *
0-
02
b1 6
#347390000000
1!
1%
1-
12
#347400000000
0!
0%
b10 *
0-
02
b10 6
#347410000000
1!
1%
1-
12
#347420000000
0!
0%
b11 *
0-
02
b11 6
#347430000000
1!
1%
1-
12
15
#347440000000
0!
0%
b100 *
0-
02
b100 6
#347450000000
1!
1%
1-
12
#347460000000
0!
0%
b101 *
0-
02
b101 6
#347470000000
1!
1%
1-
12
#347480000000
0!
0%
b110 *
0-
02
b110 6
#347490000000
1!
1%
1-
12
#347500000000
0!
0%
b111 *
0-
02
b111 6
#347510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#347520000000
0!
0%
b0 *
0-
02
b0 6
#347530000000
1!
1%
1-
12
#347540000000
0!
0%
b1 *
0-
02
b1 6
#347550000000
1!
1%
1-
12
#347560000000
0!
0%
b10 *
0-
02
b10 6
#347570000000
1!
1%
1-
12
#347580000000
0!
0%
b11 *
0-
02
b11 6
#347590000000
1!
1%
1-
12
15
#347600000000
0!
0%
b100 *
0-
02
b100 6
#347610000000
1!
1%
1-
12
#347620000000
0!
0%
b101 *
0-
02
b101 6
#347630000000
1!
1%
1-
12
#347640000000
0!
0%
b110 *
0-
02
b110 6
#347650000000
1!
1%
1-
12
#347660000000
0!
0%
b111 *
0-
02
b111 6
#347670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#347680000000
0!
0%
b0 *
0-
02
b0 6
#347690000000
1!
1%
1-
12
#347700000000
0!
0%
b1 *
0-
02
b1 6
#347710000000
1!
1%
1-
12
#347720000000
0!
0%
b10 *
0-
02
b10 6
#347730000000
1!
1%
1-
12
#347740000000
0!
0%
b11 *
0-
02
b11 6
#347750000000
1!
1%
1-
12
15
#347760000000
0!
0%
b100 *
0-
02
b100 6
#347770000000
1!
1%
1-
12
#347780000000
0!
0%
b101 *
0-
02
b101 6
#347790000000
1!
1%
1-
12
#347800000000
0!
0%
b110 *
0-
02
b110 6
#347810000000
1!
1%
1-
12
#347820000000
0!
0%
b111 *
0-
02
b111 6
#347830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#347840000000
0!
0%
b0 *
0-
02
b0 6
#347850000000
1!
1%
1-
12
#347860000000
0!
0%
b1 *
0-
02
b1 6
#347870000000
1!
1%
1-
12
#347880000000
0!
0%
b10 *
0-
02
b10 6
#347890000000
1!
1%
1-
12
#347900000000
0!
0%
b11 *
0-
02
b11 6
#347910000000
1!
1%
1-
12
15
#347920000000
0!
0%
b100 *
0-
02
b100 6
#347930000000
1!
1%
1-
12
#347940000000
0!
0%
b101 *
0-
02
b101 6
#347950000000
1!
1%
1-
12
#347960000000
0!
0%
b110 *
0-
02
b110 6
#347970000000
1!
1%
1-
12
#347980000000
0!
0%
b111 *
0-
02
b111 6
#347990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#348000000000
0!
0%
b0 *
0-
02
b0 6
#348010000000
1!
1%
1-
12
#348020000000
0!
0%
b1 *
0-
02
b1 6
#348030000000
1!
1%
1-
12
#348040000000
0!
0%
b10 *
0-
02
b10 6
#348050000000
1!
1%
1-
12
#348060000000
0!
0%
b11 *
0-
02
b11 6
#348070000000
1!
1%
1-
12
15
#348080000000
0!
0%
b100 *
0-
02
b100 6
#348090000000
1!
1%
1-
12
#348100000000
0!
0%
b101 *
0-
02
b101 6
#348110000000
1!
1%
1-
12
#348120000000
0!
0%
b110 *
0-
02
b110 6
#348130000000
1!
1%
1-
12
#348140000000
0!
0%
b111 *
0-
02
b111 6
#348150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#348160000000
0!
0%
b0 *
0-
02
b0 6
#348170000000
1!
1%
1-
12
#348180000000
0!
0%
b1 *
0-
02
b1 6
#348190000000
1!
1%
1-
12
#348200000000
0!
0%
b10 *
0-
02
b10 6
#348210000000
1!
1%
1-
12
#348220000000
0!
0%
b11 *
0-
02
b11 6
#348230000000
1!
1%
1-
12
15
#348240000000
0!
0%
b100 *
0-
02
b100 6
#348250000000
1!
1%
1-
12
#348260000000
0!
0%
b101 *
0-
02
b101 6
#348270000000
1!
1%
1-
12
#348280000000
0!
0%
b110 *
0-
02
b110 6
#348290000000
1!
1%
1-
12
#348300000000
0!
0%
b111 *
0-
02
b111 6
#348310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#348320000000
0!
0%
b0 *
0-
02
b0 6
#348330000000
1!
1%
1-
12
#348340000000
0!
0%
b1 *
0-
02
b1 6
#348350000000
1!
1%
1-
12
#348360000000
0!
0%
b10 *
0-
02
b10 6
#348370000000
1!
1%
1-
12
#348380000000
0!
0%
b11 *
0-
02
b11 6
#348390000000
1!
1%
1-
12
15
#348400000000
0!
0%
b100 *
0-
02
b100 6
#348410000000
1!
1%
1-
12
#348420000000
0!
0%
b101 *
0-
02
b101 6
#348430000000
1!
1%
1-
12
#348440000000
0!
0%
b110 *
0-
02
b110 6
#348450000000
1!
1%
1-
12
#348460000000
0!
0%
b111 *
0-
02
b111 6
#348470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#348480000000
0!
0%
b0 *
0-
02
b0 6
#348490000000
1!
1%
1-
12
#348500000000
0!
0%
b1 *
0-
02
b1 6
#348510000000
1!
1%
1-
12
#348520000000
0!
0%
b10 *
0-
02
b10 6
#348530000000
1!
1%
1-
12
#348540000000
0!
0%
b11 *
0-
02
b11 6
#348550000000
1!
1%
1-
12
15
#348560000000
0!
0%
b100 *
0-
02
b100 6
#348570000000
1!
1%
1-
12
#348580000000
0!
0%
b101 *
0-
02
b101 6
#348590000000
1!
1%
1-
12
#348600000000
0!
0%
b110 *
0-
02
b110 6
#348610000000
1!
1%
1-
12
#348620000000
0!
0%
b111 *
0-
02
b111 6
#348630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#348640000000
0!
0%
b0 *
0-
02
b0 6
#348650000000
1!
1%
1-
12
#348660000000
0!
0%
b1 *
0-
02
b1 6
#348670000000
1!
1%
1-
12
#348680000000
0!
0%
b10 *
0-
02
b10 6
#348690000000
1!
1%
1-
12
#348700000000
0!
0%
b11 *
0-
02
b11 6
#348710000000
1!
1%
1-
12
15
#348720000000
0!
0%
b100 *
0-
02
b100 6
#348730000000
1!
1%
1-
12
#348740000000
0!
0%
b101 *
0-
02
b101 6
#348750000000
1!
1%
1-
12
#348760000000
0!
0%
b110 *
0-
02
b110 6
#348770000000
1!
1%
1-
12
#348780000000
0!
0%
b111 *
0-
02
b111 6
#348790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#348800000000
0!
0%
b0 *
0-
02
b0 6
#348810000000
1!
1%
1-
12
#348820000000
0!
0%
b1 *
0-
02
b1 6
#348830000000
1!
1%
1-
12
#348840000000
0!
0%
b10 *
0-
02
b10 6
#348850000000
1!
1%
1-
12
#348860000000
0!
0%
b11 *
0-
02
b11 6
#348870000000
1!
1%
1-
12
15
#348880000000
0!
0%
b100 *
0-
02
b100 6
#348890000000
1!
1%
1-
12
#348900000000
0!
0%
b101 *
0-
02
b101 6
#348910000000
1!
1%
1-
12
#348920000000
0!
0%
b110 *
0-
02
b110 6
#348930000000
1!
1%
1-
12
#348940000000
0!
0%
b111 *
0-
02
b111 6
#348950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#348960000000
0!
0%
b0 *
0-
02
b0 6
#348970000000
1!
1%
1-
12
#348980000000
0!
0%
b1 *
0-
02
b1 6
#348990000000
1!
1%
1-
12
#349000000000
0!
0%
b10 *
0-
02
b10 6
#349010000000
1!
1%
1-
12
#349020000000
0!
0%
b11 *
0-
02
b11 6
#349030000000
1!
1%
1-
12
15
#349040000000
0!
0%
b100 *
0-
02
b100 6
#349050000000
1!
1%
1-
12
#349060000000
0!
0%
b101 *
0-
02
b101 6
#349070000000
1!
1%
1-
12
#349080000000
0!
0%
b110 *
0-
02
b110 6
#349090000000
1!
1%
1-
12
#349100000000
0!
0%
b111 *
0-
02
b111 6
#349110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#349120000000
0!
0%
b0 *
0-
02
b0 6
#349130000000
1!
1%
1-
12
#349140000000
0!
0%
b1 *
0-
02
b1 6
#349150000000
1!
1%
1-
12
#349160000000
0!
0%
b10 *
0-
02
b10 6
#349170000000
1!
1%
1-
12
#349180000000
0!
0%
b11 *
0-
02
b11 6
#349190000000
1!
1%
1-
12
15
#349200000000
0!
0%
b100 *
0-
02
b100 6
#349210000000
1!
1%
1-
12
#349220000000
0!
0%
b101 *
0-
02
b101 6
#349230000000
1!
1%
1-
12
#349240000000
0!
0%
b110 *
0-
02
b110 6
#349250000000
1!
1%
1-
12
#349260000000
0!
0%
b111 *
0-
02
b111 6
#349270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#349280000000
0!
0%
b0 *
0-
02
b0 6
#349290000000
1!
1%
1-
12
#349300000000
0!
0%
b1 *
0-
02
b1 6
#349310000000
1!
1%
1-
12
#349320000000
0!
0%
b10 *
0-
02
b10 6
#349330000000
1!
1%
1-
12
#349340000000
0!
0%
b11 *
0-
02
b11 6
#349350000000
1!
1%
1-
12
15
#349360000000
0!
0%
b100 *
0-
02
b100 6
#349370000000
1!
1%
1-
12
#349380000000
0!
0%
b101 *
0-
02
b101 6
#349390000000
1!
1%
1-
12
#349400000000
0!
0%
b110 *
0-
02
b110 6
#349410000000
1!
1%
1-
12
#349420000000
0!
0%
b111 *
0-
02
b111 6
#349430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#349440000000
0!
0%
b0 *
0-
02
b0 6
#349450000000
1!
1%
1-
12
#349460000000
0!
0%
b1 *
0-
02
b1 6
#349470000000
1!
1%
1-
12
#349480000000
0!
0%
b10 *
0-
02
b10 6
#349490000000
1!
1%
1-
12
#349500000000
0!
0%
b11 *
0-
02
b11 6
#349510000000
1!
1%
1-
12
15
#349520000000
0!
0%
b100 *
0-
02
b100 6
#349530000000
1!
1%
1-
12
#349540000000
0!
0%
b101 *
0-
02
b101 6
#349550000000
1!
1%
1-
12
#349560000000
0!
0%
b110 *
0-
02
b110 6
#349570000000
1!
1%
1-
12
#349580000000
0!
0%
b111 *
0-
02
b111 6
#349590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#349600000000
0!
0%
b0 *
0-
02
b0 6
#349610000000
1!
1%
1-
12
#349620000000
0!
0%
b1 *
0-
02
b1 6
#349630000000
1!
1%
1-
12
#349640000000
0!
0%
b10 *
0-
02
b10 6
#349650000000
1!
1%
1-
12
#349660000000
0!
0%
b11 *
0-
02
b11 6
#349670000000
1!
1%
1-
12
15
#349680000000
0!
0%
b100 *
0-
02
b100 6
#349690000000
1!
1%
1-
12
#349700000000
0!
0%
b101 *
0-
02
b101 6
#349710000000
1!
1%
1-
12
#349720000000
0!
0%
b110 *
0-
02
b110 6
#349730000000
1!
1%
1-
12
#349740000000
0!
0%
b111 *
0-
02
b111 6
#349750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#349760000000
0!
0%
b0 *
0-
02
b0 6
#349770000000
1!
1%
1-
12
#349780000000
0!
0%
b1 *
0-
02
b1 6
#349790000000
1!
1%
1-
12
#349800000000
0!
0%
b10 *
0-
02
b10 6
#349810000000
1!
1%
1-
12
#349820000000
0!
0%
b11 *
0-
02
b11 6
#349830000000
1!
1%
1-
12
15
#349840000000
0!
0%
b100 *
0-
02
b100 6
#349850000000
1!
1%
1-
12
#349860000000
0!
0%
b101 *
0-
02
b101 6
#349870000000
1!
1%
1-
12
#349880000000
0!
0%
b110 *
0-
02
b110 6
#349890000000
1!
1%
1-
12
#349900000000
0!
0%
b111 *
0-
02
b111 6
#349910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#349920000000
0!
0%
b0 *
0-
02
b0 6
#349930000000
1!
1%
1-
12
#349940000000
0!
0%
b1 *
0-
02
b1 6
#349950000000
1!
1%
1-
12
#349960000000
0!
0%
b10 *
0-
02
b10 6
#349970000000
1!
1%
1-
12
#349980000000
0!
0%
b11 *
0-
02
b11 6
#349990000000
1!
1%
1-
12
15
#350000000000
0!
0%
b100 *
0-
02
b100 6
#350010000000
1!
1%
1-
12
#350020000000
0!
0%
b101 *
0-
02
b101 6
#350030000000
1!
1%
1-
12
#350040000000
0!
0%
b110 *
0-
02
b110 6
#350050000000
1!
1%
1-
12
#350060000000
0!
0%
b111 *
0-
02
b111 6
#350070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#350080000000
0!
0%
b0 *
0-
02
b0 6
#350090000000
1!
1%
1-
12
#350100000000
0!
0%
b1 *
0-
02
b1 6
#350110000000
1!
1%
1-
12
#350120000000
0!
0%
b10 *
0-
02
b10 6
#350130000000
1!
1%
1-
12
#350140000000
0!
0%
b11 *
0-
02
b11 6
#350150000000
1!
1%
1-
12
15
#350160000000
0!
0%
b100 *
0-
02
b100 6
#350170000000
1!
1%
1-
12
#350180000000
0!
0%
b101 *
0-
02
b101 6
#350190000000
1!
1%
1-
12
#350200000000
0!
0%
b110 *
0-
02
b110 6
#350210000000
1!
1%
1-
12
#350220000000
0!
0%
b111 *
0-
02
b111 6
#350230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#350240000000
0!
0%
b0 *
0-
02
b0 6
#350250000000
1!
1%
1-
12
#350260000000
0!
0%
b1 *
0-
02
b1 6
#350270000000
1!
1%
1-
12
#350280000000
0!
0%
b10 *
0-
02
b10 6
#350290000000
1!
1%
1-
12
#350300000000
0!
0%
b11 *
0-
02
b11 6
#350310000000
1!
1%
1-
12
15
#350320000000
0!
0%
b100 *
0-
02
b100 6
#350330000000
1!
1%
1-
12
#350340000000
0!
0%
b101 *
0-
02
b101 6
#350350000000
1!
1%
1-
12
#350360000000
0!
0%
b110 *
0-
02
b110 6
#350370000000
1!
1%
1-
12
#350380000000
0!
0%
b111 *
0-
02
b111 6
#350390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#350400000000
0!
0%
b0 *
0-
02
b0 6
#350410000000
1!
1%
1-
12
#350420000000
0!
0%
b1 *
0-
02
b1 6
#350430000000
1!
1%
1-
12
#350440000000
0!
0%
b10 *
0-
02
b10 6
#350450000000
1!
1%
1-
12
#350460000000
0!
0%
b11 *
0-
02
b11 6
#350470000000
1!
1%
1-
12
15
#350480000000
0!
0%
b100 *
0-
02
b100 6
#350490000000
1!
1%
1-
12
#350500000000
0!
0%
b101 *
0-
02
b101 6
#350510000000
1!
1%
1-
12
#350520000000
0!
0%
b110 *
0-
02
b110 6
#350530000000
1!
1%
1-
12
#350540000000
0!
0%
b111 *
0-
02
b111 6
#350550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#350560000000
0!
0%
b0 *
0-
02
b0 6
#350570000000
1!
1%
1-
12
#350580000000
0!
0%
b1 *
0-
02
b1 6
#350590000000
1!
1%
1-
12
#350600000000
0!
0%
b10 *
0-
02
b10 6
#350610000000
1!
1%
1-
12
#350620000000
0!
0%
b11 *
0-
02
b11 6
#350630000000
1!
1%
1-
12
15
#350640000000
0!
0%
b100 *
0-
02
b100 6
#350650000000
1!
1%
1-
12
#350660000000
0!
0%
b101 *
0-
02
b101 6
#350670000000
1!
1%
1-
12
#350680000000
0!
0%
b110 *
0-
02
b110 6
#350690000000
1!
1%
1-
12
#350700000000
0!
0%
b111 *
0-
02
b111 6
#350710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#350720000000
0!
0%
b0 *
0-
02
b0 6
#350730000000
1!
1%
1-
12
#350740000000
0!
0%
b1 *
0-
02
b1 6
#350750000000
1!
1%
1-
12
#350760000000
0!
0%
b10 *
0-
02
b10 6
#350770000000
1!
1%
1-
12
#350780000000
0!
0%
b11 *
0-
02
b11 6
#350790000000
1!
1%
1-
12
15
#350800000000
0!
0%
b100 *
0-
02
b100 6
#350810000000
1!
1%
1-
12
#350820000000
0!
0%
b101 *
0-
02
b101 6
#350830000000
1!
1%
1-
12
#350840000000
0!
0%
b110 *
0-
02
b110 6
#350850000000
1!
1%
1-
12
#350860000000
0!
0%
b111 *
0-
02
b111 6
#350870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#350880000000
0!
0%
b0 *
0-
02
b0 6
#350890000000
1!
1%
1-
12
#350900000000
0!
0%
b1 *
0-
02
b1 6
#350910000000
1!
1%
1-
12
#350920000000
0!
0%
b10 *
0-
02
b10 6
#350930000000
1!
1%
1-
12
#350940000000
0!
0%
b11 *
0-
02
b11 6
#350950000000
1!
1%
1-
12
15
#350960000000
0!
0%
b100 *
0-
02
b100 6
#350970000000
1!
1%
1-
12
#350980000000
0!
0%
b101 *
0-
02
b101 6
#350990000000
1!
1%
1-
12
#351000000000
0!
0%
b110 *
0-
02
b110 6
#351010000000
1!
1%
1-
12
#351020000000
0!
0%
b111 *
0-
02
b111 6
#351030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#351040000000
0!
0%
b0 *
0-
02
b0 6
#351050000000
1!
1%
1-
12
#351060000000
0!
0%
b1 *
0-
02
b1 6
#351070000000
1!
1%
1-
12
#351080000000
0!
0%
b10 *
0-
02
b10 6
#351090000000
1!
1%
1-
12
#351100000000
0!
0%
b11 *
0-
02
b11 6
#351110000000
1!
1%
1-
12
15
#351120000000
0!
0%
b100 *
0-
02
b100 6
#351130000000
1!
1%
1-
12
#351140000000
0!
0%
b101 *
0-
02
b101 6
#351150000000
1!
1%
1-
12
#351160000000
0!
0%
b110 *
0-
02
b110 6
#351170000000
1!
1%
1-
12
#351180000000
0!
0%
b111 *
0-
02
b111 6
#351190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#351200000000
0!
0%
b0 *
0-
02
b0 6
#351210000000
1!
1%
1-
12
#351220000000
0!
0%
b1 *
0-
02
b1 6
#351230000000
1!
1%
1-
12
#351240000000
0!
0%
b10 *
0-
02
b10 6
#351250000000
1!
1%
1-
12
#351260000000
0!
0%
b11 *
0-
02
b11 6
#351270000000
1!
1%
1-
12
15
#351280000000
0!
0%
b100 *
0-
02
b100 6
#351290000000
1!
1%
1-
12
#351300000000
0!
0%
b101 *
0-
02
b101 6
#351310000000
1!
1%
1-
12
#351320000000
0!
0%
b110 *
0-
02
b110 6
#351330000000
1!
1%
1-
12
#351340000000
0!
0%
b111 *
0-
02
b111 6
#351350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#351360000000
0!
0%
b0 *
0-
02
b0 6
#351370000000
1!
1%
1-
12
#351380000000
0!
0%
b1 *
0-
02
b1 6
#351390000000
1!
1%
1-
12
#351400000000
0!
0%
b10 *
0-
02
b10 6
#351410000000
1!
1%
1-
12
#351420000000
0!
0%
b11 *
0-
02
b11 6
#351430000000
1!
1%
1-
12
15
#351440000000
0!
0%
b100 *
0-
02
b100 6
#351450000000
1!
1%
1-
12
#351460000000
0!
0%
b101 *
0-
02
b101 6
#351470000000
1!
1%
1-
12
#351480000000
0!
0%
b110 *
0-
02
b110 6
#351490000000
1!
1%
1-
12
#351500000000
0!
0%
b111 *
0-
02
b111 6
#351510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#351520000000
0!
0%
b0 *
0-
02
b0 6
#351530000000
1!
1%
1-
12
#351540000000
0!
0%
b1 *
0-
02
b1 6
#351550000000
1!
1%
1-
12
#351560000000
0!
0%
b10 *
0-
02
b10 6
#351570000000
1!
1%
1-
12
#351580000000
0!
0%
b11 *
0-
02
b11 6
#351590000000
1!
1%
1-
12
15
#351600000000
0!
0%
b100 *
0-
02
b100 6
#351610000000
1!
1%
1-
12
#351620000000
0!
0%
b101 *
0-
02
b101 6
#351630000000
1!
1%
1-
12
#351640000000
0!
0%
b110 *
0-
02
b110 6
#351650000000
1!
1%
1-
12
#351660000000
0!
0%
b111 *
0-
02
b111 6
#351670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#351680000000
0!
0%
b0 *
0-
02
b0 6
#351690000000
1!
1%
1-
12
#351700000000
0!
0%
b1 *
0-
02
b1 6
#351710000000
1!
1%
1-
12
#351720000000
0!
0%
b10 *
0-
02
b10 6
#351730000000
1!
1%
1-
12
#351740000000
0!
0%
b11 *
0-
02
b11 6
#351750000000
1!
1%
1-
12
15
#351760000000
0!
0%
b100 *
0-
02
b100 6
#351770000000
1!
1%
1-
12
#351780000000
0!
0%
b101 *
0-
02
b101 6
#351790000000
1!
1%
1-
12
#351800000000
0!
0%
b110 *
0-
02
b110 6
#351810000000
1!
1%
1-
12
#351820000000
0!
0%
b111 *
0-
02
b111 6
#351830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#351840000000
0!
0%
b0 *
0-
02
b0 6
#351850000000
1!
1%
1-
12
#351860000000
0!
0%
b1 *
0-
02
b1 6
#351870000000
1!
1%
1-
12
#351880000000
0!
0%
b10 *
0-
02
b10 6
#351890000000
1!
1%
1-
12
#351900000000
0!
0%
b11 *
0-
02
b11 6
#351910000000
1!
1%
1-
12
15
#351920000000
0!
0%
b100 *
0-
02
b100 6
#351930000000
1!
1%
1-
12
#351940000000
0!
0%
b101 *
0-
02
b101 6
#351950000000
1!
1%
1-
12
#351960000000
0!
0%
b110 *
0-
02
b110 6
#351970000000
1!
1%
1-
12
#351980000000
0!
0%
b111 *
0-
02
b111 6
#351990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#352000000000
0!
0%
b0 *
0-
02
b0 6
#352010000000
1!
1%
1-
12
#352020000000
0!
0%
b1 *
0-
02
b1 6
#352030000000
1!
1%
1-
12
#352040000000
0!
0%
b10 *
0-
02
b10 6
#352050000000
1!
1%
1-
12
#352060000000
0!
0%
b11 *
0-
02
b11 6
#352070000000
1!
1%
1-
12
15
#352080000000
0!
0%
b100 *
0-
02
b100 6
#352090000000
1!
1%
1-
12
#352100000000
0!
0%
b101 *
0-
02
b101 6
#352110000000
1!
1%
1-
12
#352120000000
0!
0%
b110 *
0-
02
b110 6
#352130000000
1!
1%
1-
12
#352140000000
0!
0%
b111 *
0-
02
b111 6
#352150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#352160000000
0!
0%
b0 *
0-
02
b0 6
#352170000000
1!
1%
1-
12
#352180000000
0!
0%
b1 *
0-
02
b1 6
#352190000000
1!
1%
1-
12
#352200000000
0!
0%
b10 *
0-
02
b10 6
#352210000000
1!
1%
1-
12
#352220000000
0!
0%
b11 *
0-
02
b11 6
#352230000000
1!
1%
1-
12
15
#352240000000
0!
0%
b100 *
0-
02
b100 6
#352250000000
1!
1%
1-
12
#352260000000
0!
0%
b101 *
0-
02
b101 6
#352270000000
1!
1%
1-
12
#352280000000
0!
0%
b110 *
0-
02
b110 6
#352290000000
1!
1%
1-
12
#352300000000
0!
0%
b111 *
0-
02
b111 6
#352310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#352320000000
0!
0%
b0 *
0-
02
b0 6
#352330000000
1!
1%
1-
12
#352340000000
0!
0%
b1 *
0-
02
b1 6
#352350000000
1!
1%
1-
12
#352360000000
0!
0%
b10 *
0-
02
b10 6
#352370000000
1!
1%
1-
12
#352380000000
0!
0%
b11 *
0-
02
b11 6
#352390000000
1!
1%
1-
12
15
#352400000000
0!
0%
b100 *
0-
02
b100 6
#352410000000
1!
1%
1-
12
#352420000000
0!
0%
b101 *
0-
02
b101 6
#352430000000
1!
1%
1-
12
#352440000000
0!
0%
b110 *
0-
02
b110 6
#352450000000
1!
1%
1-
12
#352460000000
0!
0%
b111 *
0-
02
b111 6
#352470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#352480000000
0!
0%
b0 *
0-
02
b0 6
#352490000000
1!
1%
1-
12
#352500000000
0!
0%
b1 *
0-
02
b1 6
#352510000000
1!
1%
1-
12
#352520000000
0!
0%
b10 *
0-
02
b10 6
#352530000000
1!
1%
1-
12
#352540000000
0!
0%
b11 *
0-
02
b11 6
#352550000000
1!
1%
1-
12
15
#352560000000
0!
0%
b100 *
0-
02
b100 6
#352570000000
1!
1%
1-
12
#352580000000
0!
0%
b101 *
0-
02
b101 6
#352590000000
1!
1%
1-
12
#352600000000
0!
0%
b110 *
0-
02
b110 6
#352610000000
1!
1%
1-
12
#352620000000
0!
0%
b111 *
0-
02
b111 6
#352630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#352640000000
0!
0%
b0 *
0-
02
b0 6
#352650000000
1!
1%
1-
12
#352660000000
0!
0%
b1 *
0-
02
b1 6
#352670000000
1!
1%
1-
12
#352680000000
0!
0%
b10 *
0-
02
b10 6
#352690000000
1!
1%
1-
12
#352700000000
0!
0%
b11 *
0-
02
b11 6
#352710000000
1!
1%
1-
12
15
#352720000000
0!
0%
b100 *
0-
02
b100 6
#352730000000
1!
1%
1-
12
#352740000000
0!
0%
b101 *
0-
02
b101 6
#352750000000
1!
1%
1-
12
#352760000000
0!
0%
b110 *
0-
02
b110 6
#352770000000
1!
1%
1-
12
#352780000000
0!
0%
b111 *
0-
02
b111 6
#352790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#352800000000
0!
0%
b0 *
0-
02
b0 6
#352810000000
1!
1%
1-
12
#352820000000
0!
0%
b1 *
0-
02
b1 6
#352830000000
1!
1%
1-
12
#352840000000
0!
0%
b10 *
0-
02
b10 6
#352850000000
1!
1%
1-
12
#352860000000
0!
0%
b11 *
0-
02
b11 6
#352870000000
1!
1%
1-
12
15
#352880000000
0!
0%
b100 *
0-
02
b100 6
#352890000000
1!
1%
1-
12
#352900000000
0!
0%
b101 *
0-
02
b101 6
#352910000000
1!
1%
1-
12
#352920000000
0!
0%
b110 *
0-
02
b110 6
#352930000000
1!
1%
1-
12
#352940000000
0!
0%
b111 *
0-
02
b111 6
#352950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#352960000000
0!
0%
b0 *
0-
02
b0 6
#352970000000
1!
1%
1-
12
#352980000000
0!
0%
b1 *
0-
02
b1 6
#352990000000
1!
1%
1-
12
#353000000000
0!
0%
b10 *
0-
02
b10 6
#353010000000
1!
1%
1-
12
#353020000000
0!
0%
b11 *
0-
02
b11 6
#353030000000
1!
1%
1-
12
15
#353040000000
0!
0%
b100 *
0-
02
b100 6
#353050000000
1!
1%
1-
12
#353060000000
0!
0%
b101 *
0-
02
b101 6
#353070000000
1!
1%
1-
12
#353080000000
0!
0%
b110 *
0-
02
b110 6
#353090000000
1!
1%
1-
12
#353100000000
0!
0%
b111 *
0-
02
b111 6
#353110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#353120000000
0!
0%
b0 *
0-
02
b0 6
#353130000000
1!
1%
1-
12
#353140000000
0!
0%
b1 *
0-
02
b1 6
#353150000000
1!
1%
1-
12
#353160000000
0!
0%
b10 *
0-
02
b10 6
#353170000000
1!
1%
1-
12
#353180000000
0!
0%
b11 *
0-
02
b11 6
#353190000000
1!
1%
1-
12
15
#353200000000
0!
0%
b100 *
0-
02
b100 6
#353210000000
1!
1%
1-
12
#353220000000
0!
0%
b101 *
0-
02
b101 6
#353230000000
1!
1%
1-
12
#353240000000
0!
0%
b110 *
0-
02
b110 6
#353250000000
1!
1%
1-
12
#353260000000
0!
0%
b111 *
0-
02
b111 6
#353270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#353280000000
0!
0%
b0 *
0-
02
b0 6
#353290000000
1!
1%
1-
12
#353300000000
0!
0%
b1 *
0-
02
b1 6
#353310000000
1!
1%
1-
12
#353320000000
0!
0%
b10 *
0-
02
b10 6
#353330000000
1!
1%
1-
12
#353340000000
0!
0%
b11 *
0-
02
b11 6
#353350000000
1!
1%
1-
12
15
#353360000000
0!
0%
b100 *
0-
02
b100 6
#353370000000
1!
1%
1-
12
#353380000000
0!
0%
b101 *
0-
02
b101 6
#353390000000
1!
1%
1-
12
#353400000000
0!
0%
b110 *
0-
02
b110 6
#353410000000
1!
1%
1-
12
#353420000000
0!
0%
b111 *
0-
02
b111 6
#353430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#353440000000
0!
0%
b0 *
0-
02
b0 6
#353450000000
1!
1%
1-
12
#353460000000
0!
0%
b1 *
0-
02
b1 6
#353470000000
1!
1%
1-
12
#353480000000
0!
0%
b10 *
0-
02
b10 6
#353490000000
1!
1%
1-
12
#353500000000
0!
0%
b11 *
0-
02
b11 6
#353510000000
1!
1%
1-
12
15
#353520000000
0!
0%
b100 *
0-
02
b100 6
#353530000000
1!
1%
1-
12
#353540000000
0!
0%
b101 *
0-
02
b101 6
#353550000000
1!
1%
1-
12
#353560000000
0!
0%
b110 *
0-
02
b110 6
#353570000000
1!
1%
1-
12
#353580000000
0!
0%
b111 *
0-
02
b111 6
#353590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#353600000000
0!
0%
b0 *
0-
02
b0 6
#353610000000
1!
1%
1-
12
#353620000000
0!
0%
b1 *
0-
02
b1 6
#353630000000
1!
1%
1-
12
#353640000000
0!
0%
b10 *
0-
02
b10 6
#353650000000
1!
1%
1-
12
#353660000000
0!
0%
b11 *
0-
02
b11 6
#353670000000
1!
1%
1-
12
15
#353680000000
0!
0%
b100 *
0-
02
b100 6
#353690000000
1!
1%
1-
12
#353700000000
0!
0%
b101 *
0-
02
b101 6
#353710000000
1!
1%
1-
12
#353720000000
0!
0%
b110 *
0-
02
b110 6
#353730000000
1!
1%
1-
12
#353740000000
0!
0%
b111 *
0-
02
b111 6
#353750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#353760000000
0!
0%
b0 *
0-
02
b0 6
#353770000000
1!
1%
1-
12
#353780000000
0!
0%
b1 *
0-
02
b1 6
#353790000000
1!
1%
1-
12
#353800000000
0!
0%
b10 *
0-
02
b10 6
#353810000000
1!
1%
1-
12
#353820000000
0!
0%
b11 *
0-
02
b11 6
#353830000000
1!
1%
1-
12
15
#353840000000
0!
0%
b100 *
0-
02
b100 6
#353850000000
1!
1%
1-
12
#353860000000
0!
0%
b101 *
0-
02
b101 6
#353870000000
1!
1%
1-
12
#353880000000
0!
0%
b110 *
0-
02
b110 6
#353890000000
1!
1%
1-
12
#353900000000
0!
0%
b111 *
0-
02
b111 6
#353910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#353920000000
0!
0%
b0 *
0-
02
b0 6
#353930000000
1!
1%
1-
12
#353940000000
0!
0%
b1 *
0-
02
b1 6
#353950000000
1!
1%
1-
12
#353960000000
0!
0%
b10 *
0-
02
b10 6
#353970000000
1!
1%
1-
12
#353980000000
0!
0%
b11 *
0-
02
b11 6
#353990000000
1!
1%
1-
12
15
#354000000000
0!
0%
b100 *
0-
02
b100 6
#354010000000
1!
1%
1-
12
#354020000000
0!
0%
b101 *
0-
02
b101 6
#354030000000
1!
1%
1-
12
#354040000000
0!
0%
b110 *
0-
02
b110 6
#354050000000
1!
1%
1-
12
#354060000000
0!
0%
b111 *
0-
02
b111 6
#354070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#354080000000
0!
0%
b0 *
0-
02
b0 6
#354090000000
1!
1%
1-
12
#354100000000
0!
0%
b1 *
0-
02
b1 6
#354110000000
1!
1%
1-
12
#354120000000
0!
0%
b10 *
0-
02
b10 6
#354130000000
1!
1%
1-
12
#354140000000
0!
0%
b11 *
0-
02
b11 6
#354150000000
1!
1%
1-
12
15
#354160000000
0!
0%
b100 *
0-
02
b100 6
#354170000000
1!
1%
1-
12
#354180000000
0!
0%
b101 *
0-
02
b101 6
#354190000000
1!
1%
1-
12
#354200000000
0!
0%
b110 *
0-
02
b110 6
#354210000000
1!
1%
1-
12
#354220000000
0!
0%
b111 *
0-
02
b111 6
#354230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#354240000000
0!
0%
b0 *
0-
02
b0 6
#354250000000
1!
1%
1-
12
#354260000000
0!
0%
b1 *
0-
02
b1 6
#354270000000
1!
1%
1-
12
#354280000000
0!
0%
b10 *
0-
02
b10 6
#354290000000
1!
1%
1-
12
#354300000000
0!
0%
b11 *
0-
02
b11 6
#354310000000
1!
1%
1-
12
15
#354320000000
0!
0%
b100 *
0-
02
b100 6
#354330000000
1!
1%
1-
12
#354340000000
0!
0%
b101 *
0-
02
b101 6
#354350000000
1!
1%
1-
12
#354360000000
0!
0%
b110 *
0-
02
b110 6
#354370000000
1!
1%
1-
12
#354380000000
0!
0%
b111 *
0-
02
b111 6
#354390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#354400000000
0!
0%
b0 *
0-
02
b0 6
#354410000000
1!
1%
1-
12
#354420000000
0!
0%
b1 *
0-
02
b1 6
#354430000000
1!
1%
1-
12
#354440000000
0!
0%
b10 *
0-
02
b10 6
#354450000000
1!
1%
1-
12
#354460000000
0!
0%
b11 *
0-
02
b11 6
#354470000000
1!
1%
1-
12
15
#354480000000
0!
0%
b100 *
0-
02
b100 6
#354490000000
1!
1%
1-
12
#354500000000
0!
0%
b101 *
0-
02
b101 6
#354510000000
1!
1%
1-
12
#354520000000
0!
0%
b110 *
0-
02
b110 6
#354530000000
1!
1%
1-
12
#354540000000
0!
0%
b111 *
0-
02
b111 6
#354550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#354560000000
0!
0%
b0 *
0-
02
b0 6
#354570000000
1!
1%
1-
12
#354580000000
0!
0%
b1 *
0-
02
b1 6
#354590000000
1!
1%
1-
12
#354600000000
0!
0%
b10 *
0-
02
b10 6
#354610000000
1!
1%
1-
12
#354620000000
0!
0%
b11 *
0-
02
b11 6
#354630000000
1!
1%
1-
12
15
#354640000000
0!
0%
b100 *
0-
02
b100 6
#354650000000
1!
1%
1-
12
#354660000000
0!
0%
b101 *
0-
02
b101 6
#354670000000
1!
1%
1-
12
#354680000000
0!
0%
b110 *
0-
02
b110 6
#354690000000
1!
1%
1-
12
#354700000000
0!
0%
b111 *
0-
02
b111 6
#354710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#354720000000
0!
0%
b0 *
0-
02
b0 6
#354730000000
1!
1%
1-
12
#354740000000
0!
0%
b1 *
0-
02
b1 6
#354750000000
1!
1%
1-
12
#354760000000
0!
0%
b10 *
0-
02
b10 6
#354770000000
1!
1%
1-
12
#354780000000
0!
0%
b11 *
0-
02
b11 6
#354790000000
1!
1%
1-
12
15
#354800000000
0!
0%
b100 *
0-
02
b100 6
#354810000000
1!
1%
1-
12
#354820000000
0!
0%
b101 *
0-
02
b101 6
#354830000000
1!
1%
1-
12
#354840000000
0!
0%
b110 *
0-
02
b110 6
#354850000000
1!
1%
1-
12
#354860000000
0!
0%
b111 *
0-
02
b111 6
#354870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#354880000000
0!
0%
b0 *
0-
02
b0 6
#354890000000
1!
1%
1-
12
#354900000000
0!
0%
b1 *
0-
02
b1 6
#354910000000
1!
1%
1-
12
#354920000000
0!
0%
b10 *
0-
02
b10 6
#354930000000
1!
1%
1-
12
#354940000000
0!
0%
b11 *
0-
02
b11 6
#354950000000
1!
1%
1-
12
15
#354960000000
0!
0%
b100 *
0-
02
b100 6
#354970000000
1!
1%
1-
12
#354980000000
0!
0%
b101 *
0-
02
b101 6
#354990000000
1!
1%
1-
12
#355000000000
0!
0%
b110 *
0-
02
b110 6
#355010000000
1!
1%
1-
12
#355020000000
0!
0%
b111 *
0-
02
b111 6
#355030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#355040000000
0!
0%
b0 *
0-
02
b0 6
#355050000000
1!
1%
1-
12
#355060000000
0!
0%
b1 *
0-
02
b1 6
#355070000000
1!
1%
1-
12
#355080000000
0!
0%
b10 *
0-
02
b10 6
#355090000000
1!
1%
1-
12
#355100000000
0!
0%
b11 *
0-
02
b11 6
#355110000000
1!
1%
1-
12
15
#355120000000
0!
0%
b100 *
0-
02
b100 6
#355130000000
1!
1%
1-
12
#355140000000
0!
0%
b101 *
0-
02
b101 6
#355150000000
1!
1%
1-
12
#355160000000
0!
0%
b110 *
0-
02
b110 6
#355170000000
1!
1%
1-
12
#355180000000
0!
0%
b111 *
0-
02
b111 6
#355190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#355200000000
0!
0%
b0 *
0-
02
b0 6
#355210000000
1!
1%
1-
12
#355220000000
0!
0%
b1 *
0-
02
b1 6
#355230000000
1!
1%
1-
12
#355240000000
0!
0%
b10 *
0-
02
b10 6
#355250000000
1!
1%
1-
12
#355260000000
0!
0%
b11 *
0-
02
b11 6
#355270000000
1!
1%
1-
12
15
#355280000000
0!
0%
b100 *
0-
02
b100 6
#355290000000
1!
1%
1-
12
#355300000000
0!
0%
b101 *
0-
02
b101 6
#355310000000
1!
1%
1-
12
#355320000000
0!
0%
b110 *
0-
02
b110 6
#355330000000
1!
1%
1-
12
#355340000000
0!
0%
b111 *
0-
02
b111 6
#355350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#355360000000
0!
0%
b0 *
0-
02
b0 6
#355370000000
1!
1%
1-
12
#355380000000
0!
0%
b1 *
0-
02
b1 6
#355390000000
1!
1%
1-
12
#355400000000
0!
0%
b10 *
0-
02
b10 6
#355410000000
1!
1%
1-
12
#355420000000
0!
0%
b11 *
0-
02
b11 6
#355430000000
1!
1%
1-
12
15
#355440000000
0!
0%
b100 *
0-
02
b100 6
#355450000000
1!
1%
1-
12
#355460000000
0!
0%
b101 *
0-
02
b101 6
#355470000000
1!
1%
1-
12
#355480000000
0!
0%
b110 *
0-
02
b110 6
#355490000000
1!
1%
1-
12
#355500000000
0!
0%
b111 *
0-
02
b111 6
#355510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#355520000000
0!
0%
b0 *
0-
02
b0 6
#355530000000
1!
1%
1-
12
#355540000000
0!
0%
b1 *
0-
02
b1 6
#355550000000
1!
1%
1-
12
#355560000000
0!
0%
b10 *
0-
02
b10 6
#355570000000
1!
1%
1-
12
#355580000000
0!
0%
b11 *
0-
02
b11 6
#355590000000
1!
1%
1-
12
15
#355600000000
0!
0%
b100 *
0-
02
b100 6
#355610000000
1!
1%
1-
12
#355620000000
0!
0%
b101 *
0-
02
b101 6
#355630000000
1!
1%
1-
12
#355640000000
0!
0%
b110 *
0-
02
b110 6
#355650000000
1!
1%
1-
12
#355660000000
0!
0%
b111 *
0-
02
b111 6
#355670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#355680000000
0!
0%
b0 *
0-
02
b0 6
#355690000000
1!
1%
1-
12
#355700000000
0!
0%
b1 *
0-
02
b1 6
#355710000000
1!
1%
1-
12
#355720000000
0!
0%
b10 *
0-
02
b10 6
#355730000000
1!
1%
1-
12
#355740000000
0!
0%
b11 *
0-
02
b11 6
#355750000000
1!
1%
1-
12
15
#355760000000
0!
0%
b100 *
0-
02
b100 6
#355770000000
1!
1%
1-
12
#355780000000
0!
0%
b101 *
0-
02
b101 6
#355790000000
1!
1%
1-
12
#355800000000
0!
0%
b110 *
0-
02
b110 6
#355810000000
1!
1%
1-
12
#355820000000
0!
0%
b111 *
0-
02
b111 6
#355830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#355840000000
0!
0%
b0 *
0-
02
b0 6
#355850000000
1!
1%
1-
12
#355860000000
0!
0%
b1 *
0-
02
b1 6
#355870000000
1!
1%
1-
12
#355880000000
0!
0%
b10 *
0-
02
b10 6
#355890000000
1!
1%
1-
12
#355900000000
0!
0%
b11 *
0-
02
b11 6
#355910000000
1!
1%
1-
12
15
#355920000000
0!
0%
b100 *
0-
02
b100 6
#355930000000
1!
1%
1-
12
#355940000000
0!
0%
b101 *
0-
02
b101 6
#355950000000
1!
1%
1-
12
#355960000000
0!
0%
b110 *
0-
02
b110 6
#355970000000
1!
1%
1-
12
#355980000000
0!
0%
b111 *
0-
02
b111 6
#355990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#356000000000
0!
0%
b0 *
0-
02
b0 6
#356010000000
1!
1%
1-
12
#356020000000
0!
0%
b1 *
0-
02
b1 6
#356030000000
1!
1%
1-
12
#356040000000
0!
0%
b10 *
0-
02
b10 6
#356050000000
1!
1%
1-
12
#356060000000
0!
0%
b11 *
0-
02
b11 6
#356070000000
1!
1%
1-
12
15
#356080000000
0!
0%
b100 *
0-
02
b100 6
#356090000000
1!
1%
1-
12
#356100000000
0!
0%
b101 *
0-
02
b101 6
#356110000000
1!
1%
1-
12
#356120000000
0!
0%
b110 *
0-
02
b110 6
#356130000000
1!
1%
1-
12
#356140000000
0!
0%
b111 *
0-
02
b111 6
#356150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#356160000000
0!
0%
b0 *
0-
02
b0 6
#356170000000
1!
1%
1-
12
#356180000000
0!
0%
b1 *
0-
02
b1 6
#356190000000
1!
1%
1-
12
#356200000000
0!
0%
b10 *
0-
02
b10 6
#356210000000
1!
1%
1-
12
#356220000000
0!
0%
b11 *
0-
02
b11 6
#356230000000
1!
1%
1-
12
15
#356240000000
0!
0%
b100 *
0-
02
b100 6
#356250000000
1!
1%
1-
12
#356260000000
0!
0%
b101 *
0-
02
b101 6
#356270000000
1!
1%
1-
12
#356280000000
0!
0%
b110 *
0-
02
b110 6
#356290000000
1!
1%
1-
12
#356300000000
0!
0%
b111 *
0-
02
b111 6
#356310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#356320000000
0!
0%
b0 *
0-
02
b0 6
#356330000000
1!
1%
1-
12
#356340000000
0!
0%
b1 *
0-
02
b1 6
#356350000000
1!
1%
1-
12
#356360000000
0!
0%
b10 *
0-
02
b10 6
#356370000000
1!
1%
1-
12
#356380000000
0!
0%
b11 *
0-
02
b11 6
#356390000000
1!
1%
1-
12
15
#356400000000
0!
0%
b100 *
0-
02
b100 6
#356410000000
1!
1%
1-
12
#356420000000
0!
0%
b101 *
0-
02
b101 6
#356430000000
1!
1%
1-
12
#356440000000
0!
0%
b110 *
0-
02
b110 6
#356450000000
1!
1%
1-
12
#356460000000
0!
0%
b111 *
0-
02
b111 6
#356470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#356480000000
0!
0%
b0 *
0-
02
b0 6
#356490000000
1!
1%
1-
12
#356500000000
0!
0%
b1 *
0-
02
b1 6
#356510000000
1!
1%
1-
12
#356520000000
0!
0%
b10 *
0-
02
b10 6
#356530000000
1!
1%
1-
12
#356540000000
0!
0%
b11 *
0-
02
b11 6
#356550000000
1!
1%
1-
12
15
#356560000000
0!
0%
b100 *
0-
02
b100 6
#356570000000
1!
1%
1-
12
#356580000000
0!
0%
b101 *
0-
02
b101 6
#356590000000
1!
1%
1-
12
#356600000000
0!
0%
b110 *
0-
02
b110 6
#356610000000
1!
1%
1-
12
#356620000000
0!
0%
b111 *
0-
02
b111 6
#356630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#356640000000
0!
0%
b0 *
0-
02
b0 6
#356650000000
1!
1%
1-
12
#356660000000
0!
0%
b1 *
0-
02
b1 6
#356670000000
1!
1%
1-
12
#356680000000
0!
0%
b10 *
0-
02
b10 6
#356690000000
1!
1%
1-
12
#356700000000
0!
0%
b11 *
0-
02
b11 6
#356710000000
1!
1%
1-
12
15
#356720000000
0!
0%
b100 *
0-
02
b100 6
#356730000000
1!
1%
1-
12
#356740000000
0!
0%
b101 *
0-
02
b101 6
#356750000000
1!
1%
1-
12
#356760000000
0!
0%
b110 *
0-
02
b110 6
#356770000000
1!
1%
1-
12
#356780000000
0!
0%
b111 *
0-
02
b111 6
#356790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#356800000000
0!
0%
b0 *
0-
02
b0 6
#356810000000
1!
1%
1-
12
#356820000000
0!
0%
b1 *
0-
02
b1 6
#356830000000
1!
1%
1-
12
#356840000000
0!
0%
b10 *
0-
02
b10 6
#356850000000
1!
1%
1-
12
#356860000000
0!
0%
b11 *
0-
02
b11 6
#356870000000
1!
1%
1-
12
15
#356880000000
0!
0%
b100 *
0-
02
b100 6
#356890000000
1!
1%
1-
12
#356900000000
0!
0%
b101 *
0-
02
b101 6
#356910000000
1!
1%
1-
12
#356920000000
0!
0%
b110 *
0-
02
b110 6
#356930000000
1!
1%
1-
12
#356940000000
0!
0%
b111 *
0-
02
b111 6
#356950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#356960000000
0!
0%
b0 *
0-
02
b0 6
#356970000000
1!
1%
1-
12
#356980000000
0!
0%
b1 *
0-
02
b1 6
#356990000000
1!
1%
1-
12
#357000000000
0!
0%
b10 *
0-
02
b10 6
#357010000000
1!
1%
1-
12
#357020000000
0!
0%
b11 *
0-
02
b11 6
#357030000000
1!
1%
1-
12
15
#357040000000
0!
0%
b100 *
0-
02
b100 6
#357050000000
1!
1%
1-
12
#357060000000
0!
0%
b101 *
0-
02
b101 6
#357070000000
1!
1%
1-
12
#357080000000
0!
0%
b110 *
0-
02
b110 6
#357090000000
1!
1%
1-
12
#357100000000
0!
0%
b111 *
0-
02
b111 6
#357110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#357120000000
0!
0%
b0 *
0-
02
b0 6
#357130000000
1!
1%
1-
12
#357140000000
0!
0%
b1 *
0-
02
b1 6
#357150000000
1!
1%
1-
12
#357160000000
0!
0%
b10 *
0-
02
b10 6
#357170000000
1!
1%
1-
12
#357180000000
0!
0%
b11 *
0-
02
b11 6
#357190000000
1!
1%
1-
12
15
#357200000000
0!
0%
b100 *
0-
02
b100 6
#357210000000
1!
1%
1-
12
#357220000000
0!
0%
b101 *
0-
02
b101 6
#357230000000
1!
1%
1-
12
#357240000000
0!
0%
b110 *
0-
02
b110 6
#357250000000
1!
1%
1-
12
#357260000000
0!
0%
b111 *
0-
02
b111 6
#357270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#357280000000
0!
0%
b0 *
0-
02
b0 6
#357290000000
1!
1%
1-
12
#357300000000
0!
0%
b1 *
0-
02
b1 6
#357310000000
1!
1%
1-
12
#357320000000
0!
0%
b10 *
0-
02
b10 6
#357330000000
1!
1%
1-
12
#357340000000
0!
0%
b11 *
0-
02
b11 6
#357350000000
1!
1%
1-
12
15
#357360000000
0!
0%
b100 *
0-
02
b100 6
#357370000000
1!
1%
1-
12
#357380000000
0!
0%
b101 *
0-
02
b101 6
#357390000000
1!
1%
1-
12
#357400000000
0!
0%
b110 *
0-
02
b110 6
#357410000000
1!
1%
1-
12
#357420000000
0!
0%
b111 *
0-
02
b111 6
#357430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#357440000000
0!
0%
b0 *
0-
02
b0 6
#357450000000
1!
1%
1-
12
#357460000000
0!
0%
b1 *
0-
02
b1 6
#357470000000
1!
1%
1-
12
#357480000000
0!
0%
b10 *
0-
02
b10 6
#357490000000
1!
1%
1-
12
#357500000000
0!
0%
b11 *
0-
02
b11 6
#357510000000
1!
1%
1-
12
15
#357520000000
0!
0%
b100 *
0-
02
b100 6
#357530000000
1!
1%
1-
12
#357540000000
0!
0%
b101 *
0-
02
b101 6
#357550000000
1!
1%
1-
12
#357560000000
0!
0%
b110 *
0-
02
b110 6
#357570000000
1!
1%
1-
12
#357580000000
0!
0%
b111 *
0-
02
b111 6
#357590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#357600000000
0!
0%
b0 *
0-
02
b0 6
#357610000000
1!
1%
1-
12
#357620000000
0!
0%
b1 *
0-
02
b1 6
#357630000000
1!
1%
1-
12
#357640000000
0!
0%
b10 *
0-
02
b10 6
#357650000000
1!
1%
1-
12
#357660000000
0!
0%
b11 *
0-
02
b11 6
#357670000000
1!
1%
1-
12
15
#357680000000
0!
0%
b100 *
0-
02
b100 6
#357690000000
1!
1%
1-
12
#357700000000
0!
0%
b101 *
0-
02
b101 6
#357710000000
1!
1%
1-
12
#357720000000
0!
0%
b110 *
0-
02
b110 6
#357730000000
1!
1%
1-
12
#357740000000
0!
0%
b111 *
0-
02
b111 6
#357750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#357760000000
0!
0%
b0 *
0-
02
b0 6
#357770000000
1!
1%
1-
12
#357780000000
0!
0%
b1 *
0-
02
b1 6
#357790000000
1!
1%
1-
12
#357800000000
0!
0%
b10 *
0-
02
b10 6
#357810000000
1!
1%
1-
12
#357820000000
0!
0%
b11 *
0-
02
b11 6
#357830000000
1!
1%
1-
12
15
#357840000000
0!
0%
b100 *
0-
02
b100 6
#357850000000
1!
1%
1-
12
#357860000000
0!
0%
b101 *
0-
02
b101 6
#357870000000
1!
1%
1-
12
#357880000000
0!
0%
b110 *
0-
02
b110 6
#357890000000
1!
1%
1-
12
#357900000000
0!
0%
b111 *
0-
02
b111 6
#357910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#357920000000
0!
0%
b0 *
0-
02
b0 6
#357930000000
1!
1%
1-
12
#357940000000
0!
0%
b1 *
0-
02
b1 6
#357950000000
1!
1%
1-
12
#357960000000
0!
0%
b10 *
0-
02
b10 6
#357970000000
1!
1%
1-
12
#357980000000
0!
0%
b11 *
0-
02
b11 6
#357990000000
1!
1%
1-
12
15
#358000000000
0!
0%
b100 *
0-
02
b100 6
#358010000000
1!
1%
1-
12
#358020000000
0!
0%
b101 *
0-
02
b101 6
#358030000000
1!
1%
1-
12
#358040000000
0!
0%
b110 *
0-
02
b110 6
#358050000000
1!
1%
1-
12
#358060000000
0!
0%
b111 *
0-
02
b111 6
#358070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#358080000000
0!
0%
b0 *
0-
02
b0 6
#358090000000
1!
1%
1-
12
#358100000000
0!
0%
b1 *
0-
02
b1 6
#358110000000
1!
1%
1-
12
#358120000000
0!
0%
b10 *
0-
02
b10 6
#358130000000
1!
1%
1-
12
#358140000000
0!
0%
b11 *
0-
02
b11 6
#358150000000
1!
1%
1-
12
15
#358160000000
0!
0%
b100 *
0-
02
b100 6
#358170000000
1!
1%
1-
12
#358180000000
0!
0%
b101 *
0-
02
b101 6
#358190000000
1!
1%
1-
12
#358200000000
0!
0%
b110 *
0-
02
b110 6
#358210000000
1!
1%
1-
12
#358220000000
0!
0%
b111 *
0-
02
b111 6
#358230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#358240000000
0!
0%
b0 *
0-
02
b0 6
#358250000000
1!
1%
1-
12
#358260000000
0!
0%
b1 *
0-
02
b1 6
#358270000000
1!
1%
1-
12
#358280000000
0!
0%
b10 *
0-
02
b10 6
#358290000000
1!
1%
1-
12
#358300000000
0!
0%
b11 *
0-
02
b11 6
#358310000000
1!
1%
1-
12
15
#358320000000
0!
0%
b100 *
0-
02
b100 6
#358330000000
1!
1%
1-
12
#358340000000
0!
0%
b101 *
0-
02
b101 6
#358350000000
1!
1%
1-
12
#358360000000
0!
0%
b110 *
0-
02
b110 6
#358370000000
1!
1%
1-
12
#358380000000
0!
0%
b111 *
0-
02
b111 6
#358390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#358400000000
0!
0%
b0 *
0-
02
b0 6
#358410000000
1!
1%
1-
12
#358420000000
0!
0%
b1 *
0-
02
b1 6
#358430000000
1!
1%
1-
12
#358440000000
0!
0%
b10 *
0-
02
b10 6
#358450000000
1!
1%
1-
12
#358460000000
0!
0%
b11 *
0-
02
b11 6
#358470000000
1!
1%
1-
12
15
#358480000000
0!
0%
b100 *
0-
02
b100 6
#358490000000
1!
1%
1-
12
#358500000000
0!
0%
b101 *
0-
02
b101 6
#358510000000
1!
1%
1-
12
#358520000000
0!
0%
b110 *
0-
02
b110 6
#358530000000
1!
1%
1-
12
#358540000000
0!
0%
b111 *
0-
02
b111 6
#358550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#358560000000
0!
0%
b0 *
0-
02
b0 6
#358570000000
1!
1%
1-
12
#358580000000
0!
0%
b1 *
0-
02
b1 6
#358590000000
1!
1%
1-
12
#358600000000
0!
0%
b10 *
0-
02
b10 6
#358610000000
1!
1%
1-
12
#358620000000
0!
0%
b11 *
0-
02
b11 6
#358630000000
1!
1%
1-
12
15
#358640000000
0!
0%
b100 *
0-
02
b100 6
#358650000000
1!
1%
1-
12
#358660000000
0!
0%
b101 *
0-
02
b101 6
#358670000000
1!
1%
1-
12
#358680000000
0!
0%
b110 *
0-
02
b110 6
#358690000000
1!
1%
1-
12
#358700000000
0!
0%
b111 *
0-
02
b111 6
#358710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#358720000000
0!
0%
b0 *
0-
02
b0 6
#358730000000
1!
1%
1-
12
#358740000000
0!
0%
b1 *
0-
02
b1 6
#358750000000
1!
1%
1-
12
#358760000000
0!
0%
b10 *
0-
02
b10 6
#358770000000
1!
1%
1-
12
#358780000000
0!
0%
b11 *
0-
02
b11 6
#358790000000
1!
1%
1-
12
15
#358800000000
0!
0%
b100 *
0-
02
b100 6
#358810000000
1!
1%
1-
12
#358820000000
0!
0%
b101 *
0-
02
b101 6
#358830000000
1!
1%
1-
12
#358840000000
0!
0%
b110 *
0-
02
b110 6
#358850000000
1!
1%
1-
12
#358860000000
0!
0%
b111 *
0-
02
b111 6
#358870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#358880000000
0!
0%
b0 *
0-
02
b0 6
#358890000000
1!
1%
1-
12
#358900000000
0!
0%
b1 *
0-
02
b1 6
#358910000000
1!
1%
1-
12
#358920000000
0!
0%
b10 *
0-
02
b10 6
#358930000000
1!
1%
1-
12
#358940000000
0!
0%
b11 *
0-
02
b11 6
#358950000000
1!
1%
1-
12
15
#358960000000
0!
0%
b100 *
0-
02
b100 6
#358970000000
1!
1%
1-
12
#358980000000
0!
0%
b101 *
0-
02
b101 6
#358990000000
1!
1%
1-
12
#359000000000
0!
0%
b110 *
0-
02
b110 6
#359010000000
1!
1%
1-
12
#359020000000
0!
0%
b111 *
0-
02
b111 6
#359030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#359040000000
0!
0%
b0 *
0-
02
b0 6
#359050000000
1!
1%
1-
12
#359060000000
0!
0%
b1 *
0-
02
b1 6
#359070000000
1!
1%
1-
12
#359080000000
0!
0%
b10 *
0-
02
b10 6
#359090000000
1!
1%
1-
12
#359100000000
0!
0%
b11 *
0-
02
b11 6
#359110000000
1!
1%
1-
12
15
#359120000000
0!
0%
b100 *
0-
02
b100 6
#359130000000
1!
1%
1-
12
#359140000000
0!
0%
b101 *
0-
02
b101 6
#359150000000
1!
1%
1-
12
#359160000000
0!
0%
b110 *
0-
02
b110 6
#359170000000
1!
1%
1-
12
#359180000000
0!
0%
b111 *
0-
02
b111 6
#359190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#359200000000
0!
0%
b0 *
0-
02
b0 6
#359210000000
1!
1%
1-
12
#359220000000
0!
0%
b1 *
0-
02
b1 6
#359230000000
1!
1%
1-
12
#359240000000
0!
0%
b10 *
0-
02
b10 6
#359250000000
1!
1%
1-
12
#359260000000
0!
0%
b11 *
0-
02
b11 6
#359270000000
1!
1%
1-
12
15
#359280000000
0!
0%
b100 *
0-
02
b100 6
#359290000000
1!
1%
1-
12
#359300000000
0!
0%
b101 *
0-
02
b101 6
#359310000000
1!
1%
1-
12
#359320000000
0!
0%
b110 *
0-
02
b110 6
#359330000000
1!
1%
1-
12
#359340000000
0!
0%
b111 *
0-
02
b111 6
#359350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#359360000000
0!
0%
b0 *
0-
02
b0 6
#359370000000
1!
1%
1-
12
#359380000000
0!
0%
b1 *
0-
02
b1 6
#359390000000
1!
1%
1-
12
#359400000000
0!
0%
b10 *
0-
02
b10 6
#359410000000
1!
1%
1-
12
#359420000000
0!
0%
b11 *
0-
02
b11 6
#359430000000
1!
1%
1-
12
15
#359440000000
0!
0%
b100 *
0-
02
b100 6
#359450000000
1!
1%
1-
12
#359460000000
0!
0%
b101 *
0-
02
b101 6
#359470000000
1!
1%
1-
12
#359480000000
0!
0%
b110 *
0-
02
b110 6
#359490000000
1!
1%
1-
12
#359500000000
0!
0%
b111 *
0-
02
b111 6
#359510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#359520000000
0!
0%
b0 *
0-
02
b0 6
#359530000000
1!
1%
1-
12
#359540000000
0!
0%
b1 *
0-
02
b1 6
#359550000000
1!
1%
1-
12
#359560000000
0!
0%
b10 *
0-
02
b10 6
#359570000000
1!
1%
1-
12
#359580000000
0!
0%
b11 *
0-
02
b11 6
#359590000000
1!
1%
1-
12
15
#359600000000
0!
0%
b100 *
0-
02
b100 6
#359610000000
1!
1%
1-
12
#359620000000
0!
0%
b101 *
0-
02
b101 6
#359630000000
1!
1%
1-
12
#359640000000
0!
0%
b110 *
0-
02
b110 6
#359650000000
1!
1%
1-
12
#359660000000
0!
0%
b111 *
0-
02
b111 6
#359670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#359680000000
0!
0%
b0 *
0-
02
b0 6
#359690000000
1!
1%
1-
12
#359700000000
0!
0%
b1 *
0-
02
b1 6
#359710000000
1!
1%
1-
12
#359720000000
0!
0%
b10 *
0-
02
b10 6
#359730000000
1!
1%
1-
12
#359740000000
0!
0%
b11 *
0-
02
b11 6
#359750000000
1!
1%
1-
12
15
#359760000000
0!
0%
b100 *
0-
02
b100 6
#359770000000
1!
1%
1-
12
#359780000000
0!
0%
b101 *
0-
02
b101 6
#359790000000
1!
1%
1-
12
#359800000000
0!
0%
b110 *
0-
02
b110 6
#359810000000
1!
1%
1-
12
#359820000000
0!
0%
b111 *
0-
02
b111 6
#359830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#359840000000
0!
0%
b0 *
0-
02
b0 6
#359850000000
1!
1%
1-
12
#359860000000
0!
0%
b1 *
0-
02
b1 6
#359870000000
1!
1%
1-
12
#359880000000
0!
0%
b10 *
0-
02
b10 6
#359890000000
1!
1%
1-
12
#359900000000
0!
0%
b11 *
0-
02
b11 6
#359910000000
1!
1%
1-
12
15
#359920000000
0!
0%
b100 *
0-
02
b100 6
#359930000000
1!
1%
1-
12
#359940000000
0!
0%
b101 *
0-
02
b101 6
#359950000000
1!
1%
1-
12
#359960000000
0!
0%
b110 *
0-
02
b110 6
#359970000000
1!
1%
1-
12
#359980000000
0!
0%
b111 *
0-
02
b111 6
#359990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#360000000000
0!
0%
b0 *
0-
02
b0 6
#360010000000
1!
1%
1-
12
#360020000000
0!
0%
b1 *
0-
02
b1 6
#360030000000
1!
1%
1-
12
#360040000000
0!
0%
b10 *
0-
02
b10 6
#360050000000
1!
1%
1-
12
#360060000000
0!
0%
b11 *
0-
02
b11 6
#360070000000
1!
1%
1-
12
15
#360080000000
0!
0%
b100 *
0-
02
b100 6
#360090000000
1!
1%
1-
12
#360100000000
0!
0%
b101 *
0-
02
b101 6
#360110000000
1!
1%
1-
12
#360120000000
0!
0%
b110 *
0-
02
b110 6
#360130000000
1!
1%
1-
12
#360140000000
0!
0%
b111 *
0-
02
b111 6
#360150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#360160000000
0!
0%
b0 *
0-
02
b0 6
#360170000000
1!
1%
1-
12
#360180000000
0!
0%
b1 *
0-
02
b1 6
#360190000000
1!
1%
1-
12
#360200000000
0!
0%
b10 *
0-
02
b10 6
#360210000000
1!
1%
1-
12
#360220000000
0!
0%
b11 *
0-
02
b11 6
#360230000000
1!
1%
1-
12
15
#360240000000
0!
0%
b100 *
0-
02
b100 6
#360250000000
1!
1%
1-
12
#360260000000
0!
0%
b101 *
0-
02
b101 6
#360270000000
1!
1%
1-
12
#360280000000
0!
0%
b110 *
0-
02
b110 6
#360290000000
1!
1%
1-
12
#360300000000
0!
0%
b111 *
0-
02
b111 6
#360310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#360320000000
0!
0%
b0 *
0-
02
b0 6
#360330000000
1!
1%
1-
12
#360340000000
0!
0%
b1 *
0-
02
b1 6
#360350000000
1!
1%
1-
12
#360360000000
0!
0%
b10 *
0-
02
b10 6
#360370000000
1!
1%
1-
12
#360380000000
0!
0%
b11 *
0-
02
b11 6
#360390000000
1!
1%
1-
12
15
#360400000000
0!
0%
b100 *
0-
02
b100 6
#360410000000
1!
1%
1-
12
#360420000000
0!
0%
b101 *
0-
02
b101 6
#360430000000
1!
1%
1-
12
#360440000000
0!
0%
b110 *
0-
02
b110 6
#360450000000
1!
1%
1-
12
#360460000000
0!
0%
b111 *
0-
02
b111 6
#360470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#360480000000
0!
0%
b0 *
0-
02
b0 6
#360490000000
1!
1%
1-
12
#360500000000
0!
0%
b1 *
0-
02
b1 6
#360510000000
1!
1%
1-
12
#360520000000
0!
0%
b10 *
0-
02
b10 6
#360530000000
1!
1%
1-
12
#360540000000
0!
0%
b11 *
0-
02
b11 6
#360550000000
1!
1%
1-
12
15
#360560000000
0!
0%
b100 *
0-
02
b100 6
#360570000000
1!
1%
1-
12
#360580000000
0!
0%
b101 *
0-
02
b101 6
#360590000000
1!
1%
1-
12
#360600000000
0!
0%
b110 *
0-
02
b110 6
#360610000000
1!
1%
1-
12
#360620000000
0!
0%
b111 *
0-
02
b111 6
#360630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#360640000000
0!
0%
b0 *
0-
02
b0 6
#360650000000
1!
1%
1-
12
#360660000000
0!
0%
b1 *
0-
02
b1 6
#360670000000
1!
1%
1-
12
#360680000000
0!
0%
b10 *
0-
02
b10 6
#360690000000
1!
1%
1-
12
#360700000000
0!
0%
b11 *
0-
02
b11 6
#360710000000
1!
1%
1-
12
15
#360720000000
0!
0%
b100 *
0-
02
b100 6
#360730000000
1!
1%
1-
12
#360740000000
0!
0%
b101 *
0-
02
b101 6
#360750000000
1!
1%
1-
12
#360760000000
0!
0%
b110 *
0-
02
b110 6
#360770000000
1!
1%
1-
12
#360780000000
0!
0%
b111 *
0-
02
b111 6
#360790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#360800000000
0!
0%
b0 *
0-
02
b0 6
#360810000000
1!
1%
1-
12
#360820000000
0!
0%
b1 *
0-
02
b1 6
#360830000000
1!
1%
1-
12
#360840000000
0!
0%
b10 *
0-
02
b10 6
#360850000000
1!
1%
1-
12
#360860000000
0!
0%
b11 *
0-
02
b11 6
#360870000000
1!
1%
1-
12
15
#360880000000
0!
0%
b100 *
0-
02
b100 6
#360890000000
1!
1%
1-
12
#360900000000
0!
0%
b101 *
0-
02
b101 6
#360910000000
1!
1%
1-
12
#360920000000
0!
0%
b110 *
0-
02
b110 6
#360930000000
1!
1%
1-
12
#360940000000
0!
0%
b111 *
0-
02
b111 6
#360950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#360960000000
0!
0%
b0 *
0-
02
b0 6
#360970000000
1!
1%
1-
12
#360980000000
0!
0%
b1 *
0-
02
b1 6
#360990000000
1!
1%
1-
12
#361000000000
0!
0%
b10 *
0-
02
b10 6
#361010000000
1!
1%
1-
12
#361020000000
0!
0%
b11 *
0-
02
b11 6
#361030000000
1!
1%
1-
12
15
#361040000000
0!
0%
b100 *
0-
02
b100 6
#361050000000
1!
1%
1-
12
#361060000000
0!
0%
b101 *
0-
02
b101 6
#361070000000
1!
1%
1-
12
#361080000000
0!
0%
b110 *
0-
02
b110 6
#361090000000
1!
1%
1-
12
#361100000000
0!
0%
b111 *
0-
02
b111 6
#361110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#361120000000
0!
0%
b0 *
0-
02
b0 6
#361130000000
1!
1%
1-
12
#361140000000
0!
0%
b1 *
0-
02
b1 6
#361150000000
1!
1%
1-
12
#361160000000
0!
0%
b10 *
0-
02
b10 6
#361170000000
1!
1%
1-
12
#361180000000
0!
0%
b11 *
0-
02
b11 6
#361190000000
1!
1%
1-
12
15
#361200000000
0!
0%
b100 *
0-
02
b100 6
#361210000000
1!
1%
1-
12
#361220000000
0!
0%
b101 *
0-
02
b101 6
#361230000000
1!
1%
1-
12
#361240000000
0!
0%
b110 *
0-
02
b110 6
#361250000000
1!
1%
1-
12
#361260000000
0!
0%
b111 *
0-
02
b111 6
#361270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#361280000000
0!
0%
b0 *
0-
02
b0 6
#361290000000
1!
1%
1-
12
#361300000000
0!
0%
b1 *
0-
02
b1 6
#361310000000
1!
1%
1-
12
#361320000000
0!
0%
b10 *
0-
02
b10 6
#361330000000
1!
1%
1-
12
#361340000000
0!
0%
b11 *
0-
02
b11 6
#361350000000
1!
1%
1-
12
15
#361360000000
0!
0%
b100 *
0-
02
b100 6
#361370000000
1!
1%
1-
12
#361380000000
0!
0%
b101 *
0-
02
b101 6
#361390000000
1!
1%
1-
12
#361400000000
0!
0%
b110 *
0-
02
b110 6
#361410000000
1!
1%
1-
12
#361420000000
0!
0%
b111 *
0-
02
b111 6
#361430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#361440000000
0!
0%
b0 *
0-
02
b0 6
#361450000000
1!
1%
1-
12
#361460000000
0!
0%
b1 *
0-
02
b1 6
#361470000000
1!
1%
1-
12
#361480000000
0!
0%
b10 *
0-
02
b10 6
#361490000000
1!
1%
1-
12
#361500000000
0!
0%
b11 *
0-
02
b11 6
#361510000000
1!
1%
1-
12
15
#361520000000
0!
0%
b100 *
0-
02
b100 6
#361530000000
1!
1%
1-
12
#361540000000
0!
0%
b101 *
0-
02
b101 6
#361550000000
1!
1%
1-
12
#361560000000
0!
0%
b110 *
0-
02
b110 6
#361570000000
1!
1%
1-
12
#361580000000
0!
0%
b111 *
0-
02
b111 6
#361590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#361600000000
0!
0%
b0 *
0-
02
b0 6
#361610000000
1!
1%
1-
12
#361620000000
0!
0%
b1 *
0-
02
b1 6
#361630000000
1!
1%
1-
12
#361640000000
0!
0%
b10 *
0-
02
b10 6
#361650000000
1!
1%
1-
12
#361660000000
0!
0%
b11 *
0-
02
b11 6
#361670000000
1!
1%
1-
12
15
#361680000000
0!
0%
b100 *
0-
02
b100 6
#361690000000
1!
1%
1-
12
#361700000000
0!
0%
b101 *
0-
02
b101 6
#361710000000
1!
1%
1-
12
#361720000000
0!
0%
b110 *
0-
02
b110 6
#361730000000
1!
1%
1-
12
#361740000000
0!
0%
b111 *
0-
02
b111 6
#361750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#361760000000
0!
0%
b0 *
0-
02
b0 6
#361770000000
1!
1%
1-
12
#361780000000
0!
0%
b1 *
0-
02
b1 6
#361790000000
1!
1%
1-
12
#361800000000
0!
0%
b10 *
0-
02
b10 6
#361810000000
1!
1%
1-
12
#361820000000
0!
0%
b11 *
0-
02
b11 6
#361830000000
1!
1%
1-
12
15
#361840000000
0!
0%
b100 *
0-
02
b100 6
#361850000000
1!
1%
1-
12
#361860000000
0!
0%
b101 *
0-
02
b101 6
#361870000000
1!
1%
1-
12
#361880000000
0!
0%
b110 *
0-
02
b110 6
#361890000000
1!
1%
1-
12
#361900000000
0!
0%
b111 *
0-
02
b111 6
#361910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#361920000000
0!
0%
b0 *
0-
02
b0 6
#361930000000
1!
1%
1-
12
#361940000000
0!
0%
b1 *
0-
02
b1 6
#361950000000
1!
1%
1-
12
#361960000000
0!
0%
b10 *
0-
02
b10 6
#361970000000
1!
1%
1-
12
#361980000000
0!
0%
b11 *
0-
02
b11 6
#361990000000
1!
1%
1-
12
15
#362000000000
0!
0%
b100 *
0-
02
b100 6
#362010000000
1!
1%
1-
12
#362020000000
0!
0%
b101 *
0-
02
b101 6
#362030000000
1!
1%
1-
12
#362040000000
0!
0%
b110 *
0-
02
b110 6
#362050000000
1!
1%
1-
12
#362060000000
0!
0%
b111 *
0-
02
b111 6
#362070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#362080000000
0!
0%
b0 *
0-
02
b0 6
#362090000000
1!
1%
1-
12
#362100000000
0!
0%
b1 *
0-
02
b1 6
#362110000000
1!
1%
1-
12
#362120000000
0!
0%
b10 *
0-
02
b10 6
#362130000000
1!
1%
1-
12
#362140000000
0!
0%
b11 *
0-
02
b11 6
#362150000000
1!
1%
1-
12
15
#362160000000
0!
0%
b100 *
0-
02
b100 6
#362170000000
1!
1%
1-
12
#362180000000
0!
0%
b101 *
0-
02
b101 6
#362190000000
1!
1%
1-
12
#362200000000
0!
0%
b110 *
0-
02
b110 6
#362210000000
1!
1%
1-
12
#362220000000
0!
0%
b111 *
0-
02
b111 6
#362230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#362240000000
0!
0%
b0 *
0-
02
b0 6
#362250000000
1!
1%
1-
12
#362260000000
0!
0%
b1 *
0-
02
b1 6
#362270000000
1!
1%
1-
12
#362280000000
0!
0%
b10 *
0-
02
b10 6
#362290000000
1!
1%
1-
12
#362300000000
0!
0%
b11 *
0-
02
b11 6
#362310000000
1!
1%
1-
12
15
#362320000000
0!
0%
b100 *
0-
02
b100 6
#362330000000
1!
1%
1-
12
#362340000000
0!
0%
b101 *
0-
02
b101 6
#362350000000
1!
1%
1-
12
#362360000000
0!
0%
b110 *
0-
02
b110 6
#362370000000
1!
1%
1-
12
#362380000000
0!
0%
b111 *
0-
02
b111 6
#362390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#362400000000
0!
0%
b0 *
0-
02
b0 6
#362410000000
1!
1%
1-
12
#362420000000
0!
0%
b1 *
0-
02
b1 6
#362430000000
1!
1%
1-
12
#362440000000
0!
0%
b10 *
0-
02
b10 6
#362450000000
1!
1%
1-
12
#362460000000
0!
0%
b11 *
0-
02
b11 6
#362470000000
1!
1%
1-
12
15
#362480000000
0!
0%
b100 *
0-
02
b100 6
#362490000000
1!
1%
1-
12
#362500000000
0!
0%
b101 *
0-
02
b101 6
#362510000000
1!
1%
1-
12
#362520000000
0!
0%
b110 *
0-
02
b110 6
#362530000000
1!
1%
1-
12
#362540000000
0!
0%
b111 *
0-
02
b111 6
#362550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#362560000000
0!
0%
b0 *
0-
02
b0 6
#362570000000
1!
1%
1-
12
#362580000000
0!
0%
b1 *
0-
02
b1 6
#362590000000
1!
1%
1-
12
#362600000000
0!
0%
b10 *
0-
02
b10 6
#362610000000
1!
1%
1-
12
#362620000000
0!
0%
b11 *
0-
02
b11 6
#362630000000
1!
1%
1-
12
15
#362640000000
0!
0%
b100 *
0-
02
b100 6
#362650000000
1!
1%
1-
12
#362660000000
0!
0%
b101 *
0-
02
b101 6
#362670000000
1!
1%
1-
12
#362680000000
0!
0%
b110 *
0-
02
b110 6
#362690000000
1!
1%
1-
12
#362700000000
0!
0%
b111 *
0-
02
b111 6
#362710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#362720000000
0!
0%
b0 *
0-
02
b0 6
#362730000000
1!
1%
1-
12
#362740000000
0!
0%
b1 *
0-
02
b1 6
#362750000000
1!
1%
1-
12
#362760000000
0!
0%
b10 *
0-
02
b10 6
#362770000000
1!
1%
1-
12
#362780000000
0!
0%
b11 *
0-
02
b11 6
#362790000000
1!
1%
1-
12
15
#362800000000
0!
0%
b100 *
0-
02
b100 6
#362810000000
1!
1%
1-
12
#362820000000
0!
0%
b101 *
0-
02
b101 6
#362830000000
1!
1%
1-
12
#362840000000
0!
0%
b110 *
0-
02
b110 6
#362850000000
1!
1%
1-
12
#362860000000
0!
0%
b111 *
0-
02
b111 6
#362870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#362880000000
0!
0%
b0 *
0-
02
b0 6
#362890000000
1!
1%
1-
12
#362900000000
0!
0%
b1 *
0-
02
b1 6
#362910000000
1!
1%
1-
12
#362920000000
0!
0%
b10 *
0-
02
b10 6
#362930000000
1!
1%
1-
12
#362940000000
0!
0%
b11 *
0-
02
b11 6
#362950000000
1!
1%
1-
12
15
#362960000000
0!
0%
b100 *
0-
02
b100 6
#362970000000
1!
1%
1-
12
#362980000000
0!
0%
b101 *
0-
02
b101 6
#362990000000
1!
1%
1-
12
#363000000000
0!
0%
b110 *
0-
02
b110 6
#363010000000
1!
1%
1-
12
#363020000000
0!
0%
b111 *
0-
02
b111 6
#363030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#363040000000
0!
0%
b0 *
0-
02
b0 6
#363050000000
1!
1%
1-
12
#363060000000
0!
0%
b1 *
0-
02
b1 6
#363070000000
1!
1%
1-
12
#363080000000
0!
0%
b10 *
0-
02
b10 6
#363090000000
1!
1%
1-
12
#363100000000
0!
0%
b11 *
0-
02
b11 6
#363110000000
1!
1%
1-
12
15
#363120000000
0!
0%
b100 *
0-
02
b100 6
#363130000000
1!
1%
1-
12
#363140000000
0!
0%
b101 *
0-
02
b101 6
#363150000000
1!
1%
1-
12
#363160000000
0!
0%
b110 *
0-
02
b110 6
#363170000000
1!
1%
1-
12
#363180000000
0!
0%
b111 *
0-
02
b111 6
#363190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#363200000000
0!
0%
b0 *
0-
02
b0 6
#363210000000
1!
1%
1-
12
#363220000000
0!
0%
b1 *
0-
02
b1 6
#363230000000
1!
1%
1-
12
#363240000000
0!
0%
b10 *
0-
02
b10 6
#363250000000
1!
1%
1-
12
#363260000000
0!
0%
b11 *
0-
02
b11 6
#363270000000
1!
1%
1-
12
15
#363280000000
0!
0%
b100 *
0-
02
b100 6
#363290000000
1!
1%
1-
12
#363300000000
0!
0%
b101 *
0-
02
b101 6
#363310000000
1!
1%
1-
12
#363320000000
0!
0%
b110 *
0-
02
b110 6
#363330000000
1!
1%
1-
12
#363340000000
0!
0%
b111 *
0-
02
b111 6
#363350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#363360000000
0!
0%
b0 *
0-
02
b0 6
#363370000000
1!
1%
1-
12
#363380000000
0!
0%
b1 *
0-
02
b1 6
#363390000000
1!
1%
1-
12
#363400000000
0!
0%
b10 *
0-
02
b10 6
#363410000000
1!
1%
1-
12
#363420000000
0!
0%
b11 *
0-
02
b11 6
#363430000000
1!
1%
1-
12
15
#363440000000
0!
0%
b100 *
0-
02
b100 6
#363450000000
1!
1%
1-
12
#363460000000
0!
0%
b101 *
0-
02
b101 6
#363470000000
1!
1%
1-
12
#363480000000
0!
0%
b110 *
0-
02
b110 6
#363490000000
1!
1%
1-
12
#363500000000
0!
0%
b111 *
0-
02
b111 6
#363510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#363520000000
0!
0%
b0 *
0-
02
b0 6
#363530000000
1!
1%
1-
12
#363540000000
0!
0%
b1 *
0-
02
b1 6
#363550000000
1!
1%
1-
12
#363560000000
0!
0%
b10 *
0-
02
b10 6
#363570000000
1!
1%
1-
12
#363580000000
0!
0%
b11 *
0-
02
b11 6
#363590000000
1!
1%
1-
12
15
#363600000000
0!
0%
b100 *
0-
02
b100 6
#363610000000
1!
1%
1-
12
#363620000000
0!
0%
b101 *
0-
02
b101 6
#363630000000
1!
1%
1-
12
#363640000000
0!
0%
b110 *
0-
02
b110 6
#363650000000
1!
1%
1-
12
#363660000000
0!
0%
b111 *
0-
02
b111 6
#363670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#363680000000
0!
0%
b0 *
0-
02
b0 6
#363690000000
1!
1%
1-
12
#363700000000
0!
0%
b1 *
0-
02
b1 6
#363710000000
1!
1%
1-
12
#363720000000
0!
0%
b10 *
0-
02
b10 6
#363730000000
1!
1%
1-
12
#363740000000
0!
0%
b11 *
0-
02
b11 6
#363750000000
1!
1%
1-
12
15
#363760000000
0!
0%
b100 *
0-
02
b100 6
#363770000000
1!
1%
1-
12
#363780000000
0!
0%
b101 *
0-
02
b101 6
#363790000000
1!
1%
1-
12
#363800000000
0!
0%
b110 *
0-
02
b110 6
#363810000000
1!
1%
1-
12
#363820000000
0!
0%
b111 *
0-
02
b111 6
#363830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#363840000000
0!
0%
b0 *
0-
02
b0 6
#363850000000
1!
1%
1-
12
#363860000000
0!
0%
b1 *
0-
02
b1 6
#363870000000
1!
1%
1-
12
#363880000000
0!
0%
b10 *
0-
02
b10 6
#363890000000
1!
1%
1-
12
#363900000000
0!
0%
b11 *
0-
02
b11 6
#363910000000
1!
1%
1-
12
15
#363920000000
0!
0%
b100 *
0-
02
b100 6
#363930000000
1!
1%
1-
12
#363940000000
0!
0%
b101 *
0-
02
b101 6
#363950000000
1!
1%
1-
12
#363960000000
0!
0%
b110 *
0-
02
b110 6
#363970000000
1!
1%
1-
12
#363980000000
0!
0%
b111 *
0-
02
b111 6
#363990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#364000000000
0!
0%
b0 *
0-
02
b0 6
#364010000000
1!
1%
1-
12
#364020000000
0!
0%
b1 *
0-
02
b1 6
#364030000000
1!
1%
1-
12
#364040000000
0!
0%
b10 *
0-
02
b10 6
#364050000000
1!
1%
1-
12
#364060000000
0!
0%
b11 *
0-
02
b11 6
#364070000000
1!
1%
1-
12
15
#364080000000
0!
0%
b100 *
0-
02
b100 6
#364090000000
1!
1%
1-
12
#364100000000
0!
0%
b101 *
0-
02
b101 6
#364110000000
1!
1%
1-
12
#364120000000
0!
0%
b110 *
0-
02
b110 6
#364130000000
1!
1%
1-
12
#364140000000
0!
0%
b111 *
0-
02
b111 6
#364150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#364160000000
0!
0%
b0 *
0-
02
b0 6
#364170000000
1!
1%
1-
12
#364180000000
0!
0%
b1 *
0-
02
b1 6
#364190000000
1!
1%
1-
12
#364200000000
0!
0%
b10 *
0-
02
b10 6
#364210000000
1!
1%
1-
12
#364220000000
0!
0%
b11 *
0-
02
b11 6
#364230000000
1!
1%
1-
12
15
#364240000000
0!
0%
b100 *
0-
02
b100 6
#364250000000
1!
1%
1-
12
#364260000000
0!
0%
b101 *
0-
02
b101 6
#364270000000
1!
1%
1-
12
#364280000000
0!
0%
b110 *
0-
02
b110 6
#364290000000
1!
1%
1-
12
#364300000000
0!
0%
b111 *
0-
02
b111 6
#364310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#364320000000
0!
0%
b0 *
0-
02
b0 6
#364330000000
1!
1%
1-
12
#364340000000
0!
0%
b1 *
0-
02
b1 6
#364350000000
1!
1%
1-
12
#364360000000
0!
0%
b10 *
0-
02
b10 6
#364370000000
1!
1%
1-
12
#364380000000
0!
0%
b11 *
0-
02
b11 6
#364390000000
1!
1%
1-
12
15
#364400000000
0!
0%
b100 *
0-
02
b100 6
#364410000000
1!
1%
1-
12
#364420000000
0!
0%
b101 *
0-
02
b101 6
#364430000000
1!
1%
1-
12
#364440000000
0!
0%
b110 *
0-
02
b110 6
#364450000000
1!
1%
1-
12
#364460000000
0!
0%
b111 *
0-
02
b111 6
#364470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#364480000000
0!
0%
b0 *
0-
02
b0 6
#364490000000
1!
1%
1-
12
#364500000000
0!
0%
b1 *
0-
02
b1 6
#364510000000
1!
1%
1-
12
#364520000000
0!
0%
b10 *
0-
02
b10 6
#364530000000
1!
1%
1-
12
#364540000000
0!
0%
b11 *
0-
02
b11 6
#364550000000
1!
1%
1-
12
15
#364560000000
0!
0%
b100 *
0-
02
b100 6
#364570000000
1!
1%
1-
12
#364580000000
0!
0%
b101 *
0-
02
b101 6
#364590000000
1!
1%
1-
12
#364600000000
0!
0%
b110 *
0-
02
b110 6
#364610000000
1!
1%
1-
12
#364620000000
0!
0%
b111 *
0-
02
b111 6
#364630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#364640000000
0!
0%
b0 *
0-
02
b0 6
#364650000000
1!
1%
1-
12
#364660000000
0!
0%
b1 *
0-
02
b1 6
#364670000000
1!
1%
1-
12
#364680000000
0!
0%
b10 *
0-
02
b10 6
#364690000000
1!
1%
1-
12
#364700000000
0!
0%
b11 *
0-
02
b11 6
#364710000000
1!
1%
1-
12
15
#364720000000
0!
0%
b100 *
0-
02
b100 6
#364730000000
1!
1%
1-
12
#364740000000
0!
0%
b101 *
0-
02
b101 6
#364750000000
1!
1%
1-
12
#364760000000
0!
0%
b110 *
0-
02
b110 6
#364770000000
1!
1%
1-
12
#364780000000
0!
0%
b111 *
0-
02
b111 6
#364790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#364800000000
0!
0%
b0 *
0-
02
b0 6
#364810000000
1!
1%
1-
12
#364820000000
0!
0%
b1 *
0-
02
b1 6
#364830000000
1!
1%
1-
12
#364840000000
0!
0%
b10 *
0-
02
b10 6
#364850000000
1!
1%
1-
12
#364860000000
0!
0%
b11 *
0-
02
b11 6
#364870000000
1!
1%
1-
12
15
#364880000000
0!
0%
b100 *
0-
02
b100 6
#364890000000
1!
1%
1-
12
#364900000000
0!
0%
b101 *
0-
02
b101 6
#364910000000
1!
1%
1-
12
#364920000000
0!
0%
b110 *
0-
02
b110 6
#364930000000
1!
1%
1-
12
#364940000000
0!
0%
b111 *
0-
02
b111 6
#364950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#364960000000
0!
0%
b0 *
0-
02
b0 6
#364970000000
1!
1%
1-
12
#364980000000
0!
0%
b1 *
0-
02
b1 6
#364990000000
1!
1%
1-
12
#365000000000
0!
0%
b10 *
0-
02
b10 6
#365010000000
1!
1%
1-
12
#365020000000
0!
0%
b11 *
0-
02
b11 6
#365030000000
1!
1%
1-
12
15
#365040000000
0!
0%
b100 *
0-
02
b100 6
#365050000000
1!
1%
1-
12
#365060000000
0!
0%
b101 *
0-
02
b101 6
#365070000000
1!
1%
1-
12
#365080000000
0!
0%
b110 *
0-
02
b110 6
#365090000000
1!
1%
1-
12
#365100000000
0!
0%
b111 *
0-
02
b111 6
#365110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#365120000000
0!
0%
b0 *
0-
02
b0 6
#365130000000
1!
1%
1-
12
#365140000000
0!
0%
b1 *
0-
02
b1 6
#365150000000
1!
1%
1-
12
#365160000000
0!
0%
b10 *
0-
02
b10 6
#365170000000
1!
1%
1-
12
#365180000000
0!
0%
b11 *
0-
02
b11 6
#365190000000
1!
1%
1-
12
15
#365200000000
0!
0%
b100 *
0-
02
b100 6
#365210000000
1!
1%
1-
12
#365220000000
0!
0%
b101 *
0-
02
b101 6
#365230000000
1!
1%
1-
12
#365240000000
0!
0%
b110 *
0-
02
b110 6
#365250000000
1!
1%
1-
12
#365260000000
0!
0%
b111 *
0-
02
b111 6
#365270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#365280000000
0!
0%
b0 *
0-
02
b0 6
#365290000000
1!
1%
1-
12
#365300000000
0!
0%
b1 *
0-
02
b1 6
#365310000000
1!
1%
1-
12
#365320000000
0!
0%
b10 *
0-
02
b10 6
#365330000000
1!
1%
1-
12
#365340000000
0!
0%
b11 *
0-
02
b11 6
#365350000000
1!
1%
1-
12
15
#365360000000
0!
0%
b100 *
0-
02
b100 6
#365370000000
1!
1%
1-
12
#365380000000
0!
0%
b101 *
0-
02
b101 6
#365390000000
1!
1%
1-
12
#365400000000
0!
0%
b110 *
0-
02
b110 6
#365410000000
1!
1%
1-
12
#365420000000
0!
0%
b111 *
0-
02
b111 6
#365430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#365440000000
0!
0%
b0 *
0-
02
b0 6
#365450000000
1!
1%
1-
12
#365460000000
0!
0%
b1 *
0-
02
b1 6
#365470000000
1!
1%
1-
12
#365480000000
0!
0%
b10 *
0-
02
b10 6
#365490000000
1!
1%
1-
12
#365500000000
0!
0%
b11 *
0-
02
b11 6
#365510000000
1!
1%
1-
12
15
#365520000000
0!
0%
b100 *
0-
02
b100 6
#365530000000
1!
1%
1-
12
#365540000000
0!
0%
b101 *
0-
02
b101 6
#365550000000
1!
1%
1-
12
#365560000000
0!
0%
b110 *
0-
02
b110 6
#365570000000
1!
1%
1-
12
#365580000000
0!
0%
b111 *
0-
02
b111 6
#365590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#365600000000
0!
0%
b0 *
0-
02
b0 6
#365610000000
1!
1%
1-
12
#365620000000
0!
0%
b1 *
0-
02
b1 6
#365630000000
1!
1%
1-
12
#365640000000
0!
0%
b10 *
0-
02
b10 6
#365650000000
1!
1%
1-
12
#365660000000
0!
0%
b11 *
0-
02
b11 6
#365670000000
1!
1%
1-
12
15
#365680000000
0!
0%
b100 *
0-
02
b100 6
#365690000000
1!
1%
1-
12
#365700000000
0!
0%
b101 *
0-
02
b101 6
#365710000000
1!
1%
1-
12
#365720000000
0!
0%
b110 *
0-
02
b110 6
#365730000000
1!
1%
1-
12
#365740000000
0!
0%
b111 *
0-
02
b111 6
#365750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#365760000000
0!
0%
b0 *
0-
02
b0 6
#365770000000
1!
1%
1-
12
#365780000000
0!
0%
b1 *
0-
02
b1 6
#365790000000
1!
1%
1-
12
#365800000000
0!
0%
b10 *
0-
02
b10 6
#365810000000
1!
1%
1-
12
#365820000000
0!
0%
b11 *
0-
02
b11 6
#365830000000
1!
1%
1-
12
15
#365840000000
0!
0%
b100 *
0-
02
b100 6
#365850000000
1!
1%
1-
12
#365860000000
0!
0%
b101 *
0-
02
b101 6
#365870000000
1!
1%
1-
12
#365880000000
0!
0%
b110 *
0-
02
b110 6
#365890000000
1!
1%
1-
12
#365900000000
0!
0%
b111 *
0-
02
b111 6
#365910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#365920000000
0!
0%
b0 *
0-
02
b0 6
#365930000000
1!
1%
1-
12
#365940000000
0!
0%
b1 *
0-
02
b1 6
#365950000000
1!
1%
1-
12
#365960000000
0!
0%
b10 *
0-
02
b10 6
#365970000000
1!
1%
1-
12
#365980000000
0!
0%
b11 *
0-
02
b11 6
#365990000000
1!
1%
1-
12
15
#366000000000
0!
0%
b100 *
0-
02
b100 6
#366010000000
1!
1%
1-
12
#366020000000
0!
0%
b101 *
0-
02
b101 6
#366030000000
1!
1%
1-
12
#366040000000
0!
0%
b110 *
0-
02
b110 6
#366050000000
1!
1%
1-
12
#366060000000
0!
0%
b111 *
0-
02
b111 6
#366070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#366080000000
0!
0%
b0 *
0-
02
b0 6
#366090000000
1!
1%
1-
12
#366100000000
0!
0%
b1 *
0-
02
b1 6
#366110000000
1!
1%
1-
12
#366120000000
0!
0%
b10 *
0-
02
b10 6
#366130000000
1!
1%
1-
12
#366140000000
0!
0%
b11 *
0-
02
b11 6
#366150000000
1!
1%
1-
12
15
#366160000000
0!
0%
b100 *
0-
02
b100 6
#366170000000
1!
1%
1-
12
#366180000000
0!
0%
b101 *
0-
02
b101 6
#366190000000
1!
1%
1-
12
#366200000000
0!
0%
b110 *
0-
02
b110 6
#366210000000
1!
1%
1-
12
#366220000000
0!
0%
b111 *
0-
02
b111 6
#366230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#366240000000
0!
0%
b0 *
0-
02
b0 6
#366250000000
1!
1%
1-
12
#366260000000
0!
0%
b1 *
0-
02
b1 6
#366270000000
1!
1%
1-
12
#366280000000
0!
0%
b10 *
0-
02
b10 6
#366290000000
1!
1%
1-
12
#366300000000
0!
0%
b11 *
0-
02
b11 6
#366310000000
1!
1%
1-
12
15
#366320000000
0!
0%
b100 *
0-
02
b100 6
#366330000000
1!
1%
1-
12
#366340000000
0!
0%
b101 *
0-
02
b101 6
#366350000000
1!
1%
1-
12
#366360000000
0!
0%
b110 *
0-
02
b110 6
#366370000000
1!
1%
1-
12
#366380000000
0!
0%
b111 *
0-
02
b111 6
#366390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#366400000000
0!
0%
b0 *
0-
02
b0 6
#366410000000
1!
1%
1-
12
#366420000000
0!
0%
b1 *
0-
02
b1 6
#366430000000
1!
1%
1-
12
#366440000000
0!
0%
b10 *
0-
02
b10 6
#366450000000
1!
1%
1-
12
#366460000000
0!
0%
b11 *
0-
02
b11 6
#366470000000
1!
1%
1-
12
15
#366480000000
0!
0%
b100 *
0-
02
b100 6
#366490000000
1!
1%
1-
12
#366500000000
0!
0%
b101 *
0-
02
b101 6
#366510000000
1!
1%
1-
12
#366520000000
0!
0%
b110 *
0-
02
b110 6
#366530000000
1!
1%
1-
12
#366540000000
0!
0%
b111 *
0-
02
b111 6
#366550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#366560000000
0!
0%
b0 *
0-
02
b0 6
#366570000000
1!
1%
1-
12
#366580000000
0!
0%
b1 *
0-
02
b1 6
#366590000000
1!
1%
1-
12
#366600000000
0!
0%
b10 *
0-
02
b10 6
#366610000000
1!
1%
1-
12
#366620000000
0!
0%
b11 *
0-
02
b11 6
#366630000000
1!
1%
1-
12
15
#366640000000
0!
0%
b100 *
0-
02
b100 6
#366650000000
1!
1%
1-
12
#366660000000
0!
0%
b101 *
0-
02
b101 6
#366670000000
1!
1%
1-
12
#366680000000
0!
0%
b110 *
0-
02
b110 6
#366690000000
1!
1%
1-
12
#366700000000
0!
0%
b111 *
0-
02
b111 6
#366710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#366720000000
0!
0%
b0 *
0-
02
b0 6
#366730000000
1!
1%
1-
12
#366740000000
0!
0%
b1 *
0-
02
b1 6
#366750000000
1!
1%
1-
12
#366760000000
0!
0%
b10 *
0-
02
b10 6
#366770000000
1!
1%
1-
12
#366780000000
0!
0%
b11 *
0-
02
b11 6
#366790000000
1!
1%
1-
12
15
#366800000000
0!
0%
b100 *
0-
02
b100 6
#366810000000
1!
1%
1-
12
#366820000000
0!
0%
b101 *
0-
02
b101 6
#366830000000
1!
1%
1-
12
#366840000000
0!
0%
b110 *
0-
02
b110 6
#366850000000
1!
1%
1-
12
#366860000000
0!
0%
b111 *
0-
02
b111 6
#366870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#366880000000
0!
0%
b0 *
0-
02
b0 6
#366890000000
1!
1%
1-
12
#366900000000
0!
0%
b1 *
0-
02
b1 6
#366910000000
1!
1%
1-
12
#366920000000
0!
0%
b10 *
0-
02
b10 6
#366930000000
1!
1%
1-
12
#366940000000
0!
0%
b11 *
0-
02
b11 6
#366950000000
1!
1%
1-
12
15
#366960000000
0!
0%
b100 *
0-
02
b100 6
#366970000000
1!
1%
1-
12
#366980000000
0!
0%
b101 *
0-
02
b101 6
#366990000000
1!
1%
1-
12
#367000000000
0!
0%
b110 *
0-
02
b110 6
#367010000000
1!
1%
1-
12
#367020000000
0!
0%
b111 *
0-
02
b111 6
#367030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#367040000000
0!
0%
b0 *
0-
02
b0 6
#367050000000
1!
1%
1-
12
#367060000000
0!
0%
b1 *
0-
02
b1 6
#367070000000
1!
1%
1-
12
#367080000000
0!
0%
b10 *
0-
02
b10 6
#367090000000
1!
1%
1-
12
#367100000000
0!
0%
b11 *
0-
02
b11 6
#367110000000
1!
1%
1-
12
15
#367120000000
0!
0%
b100 *
0-
02
b100 6
#367130000000
1!
1%
1-
12
#367140000000
0!
0%
b101 *
0-
02
b101 6
#367150000000
1!
1%
1-
12
#367160000000
0!
0%
b110 *
0-
02
b110 6
#367170000000
1!
1%
1-
12
#367180000000
0!
0%
b111 *
0-
02
b111 6
#367190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#367200000000
0!
0%
b0 *
0-
02
b0 6
#367210000000
1!
1%
1-
12
#367220000000
0!
0%
b1 *
0-
02
b1 6
#367230000000
1!
1%
1-
12
#367240000000
0!
0%
b10 *
0-
02
b10 6
#367250000000
1!
1%
1-
12
#367260000000
0!
0%
b11 *
0-
02
b11 6
#367270000000
1!
1%
1-
12
15
#367280000000
0!
0%
b100 *
0-
02
b100 6
#367290000000
1!
1%
1-
12
#367300000000
0!
0%
b101 *
0-
02
b101 6
#367310000000
1!
1%
1-
12
#367320000000
0!
0%
b110 *
0-
02
b110 6
#367330000000
1!
1%
1-
12
#367340000000
0!
0%
b111 *
0-
02
b111 6
#367350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#367360000000
0!
0%
b0 *
0-
02
b0 6
#367370000000
1!
1%
1-
12
#367380000000
0!
0%
b1 *
0-
02
b1 6
#367390000000
1!
1%
1-
12
#367400000000
0!
0%
b10 *
0-
02
b10 6
#367410000000
1!
1%
1-
12
#367420000000
0!
0%
b11 *
0-
02
b11 6
#367430000000
1!
1%
1-
12
15
#367440000000
0!
0%
b100 *
0-
02
b100 6
#367450000000
1!
1%
1-
12
#367460000000
0!
0%
b101 *
0-
02
b101 6
#367470000000
1!
1%
1-
12
#367480000000
0!
0%
b110 *
0-
02
b110 6
#367490000000
1!
1%
1-
12
#367500000000
0!
0%
b111 *
0-
02
b111 6
#367510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#367520000000
0!
0%
b0 *
0-
02
b0 6
#367530000000
1!
1%
1-
12
#367540000000
0!
0%
b1 *
0-
02
b1 6
#367550000000
1!
1%
1-
12
#367560000000
0!
0%
b10 *
0-
02
b10 6
#367570000000
1!
1%
1-
12
#367580000000
0!
0%
b11 *
0-
02
b11 6
#367590000000
1!
1%
1-
12
15
#367600000000
0!
0%
b100 *
0-
02
b100 6
#367610000000
1!
1%
1-
12
#367620000000
0!
0%
b101 *
0-
02
b101 6
#367630000000
1!
1%
1-
12
#367640000000
0!
0%
b110 *
0-
02
b110 6
#367650000000
1!
1%
1-
12
#367660000000
0!
0%
b111 *
0-
02
b111 6
#367670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#367680000000
0!
0%
b0 *
0-
02
b0 6
#367690000000
1!
1%
1-
12
#367700000000
0!
0%
b1 *
0-
02
b1 6
#367710000000
1!
1%
1-
12
#367720000000
0!
0%
b10 *
0-
02
b10 6
#367730000000
1!
1%
1-
12
#367740000000
0!
0%
b11 *
0-
02
b11 6
#367750000000
1!
1%
1-
12
15
#367760000000
0!
0%
b100 *
0-
02
b100 6
#367770000000
1!
1%
1-
12
#367780000000
0!
0%
b101 *
0-
02
b101 6
#367790000000
1!
1%
1-
12
#367800000000
0!
0%
b110 *
0-
02
b110 6
#367810000000
1!
1%
1-
12
#367820000000
0!
0%
b111 *
0-
02
b111 6
#367830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#367840000000
0!
0%
b0 *
0-
02
b0 6
#367850000000
1!
1%
1-
12
#367860000000
0!
0%
b1 *
0-
02
b1 6
#367870000000
1!
1%
1-
12
#367880000000
0!
0%
b10 *
0-
02
b10 6
#367890000000
1!
1%
1-
12
#367900000000
0!
0%
b11 *
0-
02
b11 6
#367910000000
1!
1%
1-
12
15
#367920000000
0!
0%
b100 *
0-
02
b100 6
#367930000000
1!
1%
1-
12
#367940000000
0!
0%
b101 *
0-
02
b101 6
#367950000000
1!
1%
1-
12
#367960000000
0!
0%
b110 *
0-
02
b110 6
#367970000000
1!
1%
1-
12
#367980000000
0!
0%
b111 *
0-
02
b111 6
#367990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#368000000000
0!
0%
b0 *
0-
02
b0 6
#368010000000
1!
1%
1-
12
#368020000000
0!
0%
b1 *
0-
02
b1 6
#368030000000
1!
1%
1-
12
#368040000000
0!
0%
b10 *
0-
02
b10 6
#368050000000
1!
1%
1-
12
#368060000000
0!
0%
b11 *
0-
02
b11 6
#368070000000
1!
1%
1-
12
15
#368080000000
0!
0%
b100 *
0-
02
b100 6
#368090000000
1!
1%
1-
12
#368100000000
0!
0%
b101 *
0-
02
b101 6
#368110000000
1!
1%
1-
12
#368120000000
0!
0%
b110 *
0-
02
b110 6
#368130000000
1!
1%
1-
12
#368140000000
0!
0%
b111 *
0-
02
b111 6
#368150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#368160000000
0!
0%
b0 *
0-
02
b0 6
#368170000000
1!
1%
1-
12
#368180000000
0!
0%
b1 *
0-
02
b1 6
#368190000000
1!
1%
1-
12
#368200000000
0!
0%
b10 *
0-
02
b10 6
#368210000000
1!
1%
1-
12
#368220000000
0!
0%
b11 *
0-
02
b11 6
#368230000000
1!
1%
1-
12
15
#368240000000
0!
0%
b100 *
0-
02
b100 6
#368250000000
1!
1%
1-
12
#368260000000
0!
0%
b101 *
0-
02
b101 6
#368270000000
1!
1%
1-
12
#368280000000
0!
0%
b110 *
0-
02
b110 6
#368290000000
1!
1%
1-
12
#368300000000
0!
0%
b111 *
0-
02
b111 6
#368310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#368320000000
0!
0%
b0 *
0-
02
b0 6
#368330000000
1!
1%
1-
12
#368340000000
0!
0%
b1 *
0-
02
b1 6
#368350000000
1!
1%
1-
12
#368360000000
0!
0%
b10 *
0-
02
b10 6
#368370000000
1!
1%
1-
12
#368380000000
0!
0%
b11 *
0-
02
b11 6
#368390000000
1!
1%
1-
12
15
#368400000000
0!
0%
b100 *
0-
02
b100 6
#368410000000
1!
1%
1-
12
#368420000000
0!
0%
b101 *
0-
02
b101 6
#368430000000
1!
1%
1-
12
#368440000000
0!
0%
b110 *
0-
02
b110 6
#368450000000
1!
1%
1-
12
#368460000000
0!
0%
b111 *
0-
02
b111 6
#368470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#368480000000
0!
0%
b0 *
0-
02
b0 6
#368490000000
1!
1%
1-
12
#368500000000
0!
0%
b1 *
0-
02
b1 6
#368510000000
1!
1%
1-
12
#368520000000
0!
0%
b10 *
0-
02
b10 6
#368530000000
1!
1%
1-
12
#368540000000
0!
0%
b11 *
0-
02
b11 6
#368550000000
1!
1%
1-
12
15
#368560000000
0!
0%
b100 *
0-
02
b100 6
#368570000000
1!
1%
1-
12
#368580000000
0!
0%
b101 *
0-
02
b101 6
#368590000000
1!
1%
1-
12
#368600000000
0!
0%
b110 *
0-
02
b110 6
#368610000000
1!
1%
1-
12
#368620000000
0!
0%
b111 *
0-
02
b111 6
#368630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#368640000000
0!
0%
b0 *
0-
02
b0 6
#368650000000
1!
1%
1-
12
#368660000000
0!
0%
b1 *
0-
02
b1 6
#368670000000
1!
1%
1-
12
#368680000000
0!
0%
b10 *
0-
02
b10 6
#368690000000
1!
1%
1-
12
#368700000000
0!
0%
b11 *
0-
02
b11 6
#368710000000
1!
1%
1-
12
15
#368720000000
0!
0%
b100 *
0-
02
b100 6
#368730000000
1!
1%
1-
12
#368740000000
0!
0%
b101 *
0-
02
b101 6
#368750000000
1!
1%
1-
12
#368760000000
0!
0%
b110 *
0-
02
b110 6
#368770000000
1!
1%
1-
12
#368780000000
0!
0%
b111 *
0-
02
b111 6
#368790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#368800000000
0!
0%
b0 *
0-
02
b0 6
#368810000000
1!
1%
1-
12
#368820000000
0!
0%
b1 *
0-
02
b1 6
#368830000000
1!
1%
1-
12
#368840000000
0!
0%
b10 *
0-
02
b10 6
#368850000000
1!
1%
1-
12
#368860000000
0!
0%
b11 *
0-
02
b11 6
#368870000000
1!
1%
1-
12
15
#368880000000
0!
0%
b100 *
0-
02
b100 6
#368890000000
1!
1%
1-
12
#368900000000
0!
0%
b101 *
0-
02
b101 6
#368910000000
1!
1%
1-
12
#368920000000
0!
0%
b110 *
0-
02
b110 6
#368930000000
1!
1%
1-
12
#368940000000
0!
0%
b111 *
0-
02
b111 6
#368950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#368960000000
0!
0%
b0 *
0-
02
b0 6
#368970000000
1!
1%
1-
12
#368980000000
0!
0%
b1 *
0-
02
b1 6
#368990000000
1!
1%
1-
12
#369000000000
0!
0%
b10 *
0-
02
b10 6
#369010000000
1!
1%
1-
12
#369020000000
0!
0%
b11 *
0-
02
b11 6
#369030000000
1!
1%
1-
12
15
#369040000000
0!
0%
b100 *
0-
02
b100 6
#369050000000
1!
1%
1-
12
#369060000000
0!
0%
b101 *
0-
02
b101 6
#369070000000
1!
1%
1-
12
#369080000000
0!
0%
b110 *
0-
02
b110 6
#369090000000
1!
1%
1-
12
#369100000000
0!
0%
b111 *
0-
02
b111 6
#369110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#369120000000
0!
0%
b0 *
0-
02
b0 6
#369130000000
1!
1%
1-
12
#369140000000
0!
0%
b1 *
0-
02
b1 6
#369150000000
1!
1%
1-
12
#369160000000
0!
0%
b10 *
0-
02
b10 6
#369170000000
1!
1%
1-
12
#369180000000
0!
0%
b11 *
0-
02
b11 6
#369190000000
1!
1%
1-
12
15
#369200000000
0!
0%
b100 *
0-
02
b100 6
#369210000000
1!
1%
1-
12
#369220000000
0!
0%
b101 *
0-
02
b101 6
#369230000000
1!
1%
1-
12
#369240000000
0!
0%
b110 *
0-
02
b110 6
#369250000000
1!
1%
1-
12
#369260000000
0!
0%
b111 *
0-
02
b111 6
#369270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#369280000000
0!
0%
b0 *
0-
02
b0 6
#369290000000
1!
1%
1-
12
#369300000000
0!
0%
b1 *
0-
02
b1 6
#369310000000
1!
1%
1-
12
#369320000000
0!
0%
b10 *
0-
02
b10 6
#369330000000
1!
1%
1-
12
#369340000000
0!
0%
b11 *
0-
02
b11 6
#369350000000
1!
1%
1-
12
15
#369360000000
0!
0%
b100 *
0-
02
b100 6
#369370000000
1!
1%
1-
12
#369380000000
0!
0%
b101 *
0-
02
b101 6
#369390000000
1!
1%
1-
12
#369400000000
0!
0%
b110 *
0-
02
b110 6
#369410000000
1!
1%
1-
12
#369420000000
0!
0%
b111 *
0-
02
b111 6
#369430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#369440000000
0!
0%
b0 *
0-
02
b0 6
#369450000000
1!
1%
1-
12
#369460000000
0!
0%
b1 *
0-
02
b1 6
#369470000000
1!
1%
1-
12
#369480000000
0!
0%
b10 *
0-
02
b10 6
#369490000000
1!
1%
1-
12
#369500000000
0!
0%
b11 *
0-
02
b11 6
#369510000000
1!
1%
1-
12
15
#369520000000
0!
0%
b100 *
0-
02
b100 6
#369530000000
1!
1%
1-
12
#369540000000
0!
0%
b101 *
0-
02
b101 6
#369550000000
1!
1%
1-
12
#369560000000
0!
0%
b110 *
0-
02
b110 6
#369570000000
1!
1%
1-
12
#369580000000
0!
0%
b111 *
0-
02
b111 6
#369590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#369600000000
0!
0%
b0 *
0-
02
b0 6
#369610000000
1!
1%
1-
12
#369620000000
0!
0%
b1 *
0-
02
b1 6
#369630000000
1!
1%
1-
12
#369640000000
0!
0%
b10 *
0-
02
b10 6
#369650000000
1!
1%
1-
12
#369660000000
0!
0%
b11 *
0-
02
b11 6
#369670000000
1!
1%
1-
12
15
#369680000000
0!
0%
b100 *
0-
02
b100 6
#369690000000
1!
1%
1-
12
#369700000000
0!
0%
b101 *
0-
02
b101 6
#369710000000
1!
1%
1-
12
#369720000000
0!
0%
b110 *
0-
02
b110 6
#369730000000
1!
1%
1-
12
#369740000000
0!
0%
b111 *
0-
02
b111 6
#369750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#369760000000
0!
0%
b0 *
0-
02
b0 6
#369770000000
1!
1%
1-
12
#369780000000
0!
0%
b1 *
0-
02
b1 6
#369790000000
1!
1%
1-
12
#369800000000
0!
0%
b10 *
0-
02
b10 6
#369810000000
1!
1%
1-
12
#369820000000
0!
0%
b11 *
0-
02
b11 6
#369830000000
1!
1%
1-
12
15
#369840000000
0!
0%
b100 *
0-
02
b100 6
#369850000000
1!
1%
1-
12
#369860000000
0!
0%
b101 *
0-
02
b101 6
#369870000000
1!
1%
1-
12
#369880000000
0!
0%
b110 *
0-
02
b110 6
#369890000000
1!
1%
1-
12
#369900000000
0!
0%
b111 *
0-
02
b111 6
#369910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#369920000000
0!
0%
b0 *
0-
02
b0 6
#369930000000
1!
1%
1-
12
#369940000000
0!
0%
b1 *
0-
02
b1 6
#369950000000
1!
1%
1-
12
#369960000000
0!
0%
b10 *
0-
02
b10 6
#369970000000
1!
1%
1-
12
#369980000000
0!
0%
b11 *
0-
02
b11 6
#369990000000
1!
1%
1-
12
15
#370000000000
0!
0%
b100 *
0-
02
b100 6
#370010000000
1!
1%
1-
12
#370020000000
0!
0%
b101 *
0-
02
b101 6
#370030000000
1!
1%
1-
12
#370040000000
0!
0%
b110 *
0-
02
b110 6
#370050000000
1!
1%
1-
12
#370060000000
0!
0%
b111 *
0-
02
b111 6
#370070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#370080000000
0!
0%
b0 *
0-
02
b0 6
#370090000000
1!
1%
1-
12
#370100000000
0!
0%
b1 *
0-
02
b1 6
#370110000000
1!
1%
1-
12
#370120000000
0!
0%
b10 *
0-
02
b10 6
#370130000000
1!
1%
1-
12
#370140000000
0!
0%
b11 *
0-
02
b11 6
#370150000000
1!
1%
1-
12
15
#370160000000
0!
0%
b100 *
0-
02
b100 6
#370170000000
1!
1%
1-
12
#370180000000
0!
0%
b101 *
0-
02
b101 6
#370190000000
1!
1%
1-
12
#370200000000
0!
0%
b110 *
0-
02
b110 6
#370210000000
1!
1%
1-
12
#370220000000
0!
0%
b111 *
0-
02
b111 6
#370230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#370240000000
0!
0%
b0 *
0-
02
b0 6
#370250000000
1!
1%
1-
12
#370260000000
0!
0%
b1 *
0-
02
b1 6
#370270000000
1!
1%
1-
12
#370280000000
0!
0%
b10 *
0-
02
b10 6
#370290000000
1!
1%
1-
12
#370300000000
0!
0%
b11 *
0-
02
b11 6
#370310000000
1!
1%
1-
12
15
#370320000000
0!
0%
b100 *
0-
02
b100 6
#370330000000
1!
1%
1-
12
#370340000000
0!
0%
b101 *
0-
02
b101 6
#370350000000
1!
1%
1-
12
#370360000000
0!
0%
b110 *
0-
02
b110 6
#370370000000
1!
1%
1-
12
#370380000000
0!
0%
b111 *
0-
02
b111 6
#370390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#370400000000
0!
0%
b0 *
0-
02
b0 6
#370410000000
1!
1%
1-
12
#370420000000
0!
0%
b1 *
0-
02
b1 6
#370430000000
1!
1%
1-
12
#370440000000
0!
0%
b10 *
0-
02
b10 6
#370450000000
1!
1%
1-
12
#370460000000
0!
0%
b11 *
0-
02
b11 6
#370470000000
1!
1%
1-
12
15
#370480000000
0!
0%
b100 *
0-
02
b100 6
#370490000000
1!
1%
1-
12
#370500000000
0!
0%
b101 *
0-
02
b101 6
#370510000000
1!
1%
1-
12
#370520000000
0!
0%
b110 *
0-
02
b110 6
#370530000000
1!
1%
1-
12
#370540000000
0!
0%
b111 *
0-
02
b111 6
#370550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#370560000000
0!
0%
b0 *
0-
02
b0 6
#370570000000
1!
1%
1-
12
#370580000000
0!
0%
b1 *
0-
02
b1 6
#370590000000
1!
1%
1-
12
#370600000000
0!
0%
b10 *
0-
02
b10 6
#370610000000
1!
1%
1-
12
#370620000000
0!
0%
b11 *
0-
02
b11 6
#370630000000
1!
1%
1-
12
15
#370640000000
0!
0%
b100 *
0-
02
b100 6
#370650000000
1!
1%
1-
12
#370660000000
0!
0%
b101 *
0-
02
b101 6
#370670000000
1!
1%
1-
12
#370680000000
0!
0%
b110 *
0-
02
b110 6
#370690000000
1!
1%
1-
12
#370700000000
0!
0%
b111 *
0-
02
b111 6
#370710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#370720000000
0!
0%
b0 *
0-
02
b0 6
#370730000000
1!
1%
1-
12
#370740000000
0!
0%
b1 *
0-
02
b1 6
#370750000000
1!
1%
1-
12
#370760000000
0!
0%
b10 *
0-
02
b10 6
#370770000000
1!
1%
1-
12
#370780000000
0!
0%
b11 *
0-
02
b11 6
#370790000000
1!
1%
1-
12
15
#370800000000
0!
0%
b100 *
0-
02
b100 6
#370810000000
1!
1%
1-
12
#370820000000
0!
0%
b101 *
0-
02
b101 6
#370830000000
1!
1%
1-
12
#370840000000
0!
0%
b110 *
0-
02
b110 6
#370850000000
1!
1%
1-
12
#370860000000
0!
0%
b111 *
0-
02
b111 6
#370870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#370880000000
0!
0%
b0 *
0-
02
b0 6
#370890000000
1!
1%
1-
12
#370900000000
0!
0%
b1 *
0-
02
b1 6
#370910000000
1!
1%
1-
12
#370920000000
0!
0%
b10 *
0-
02
b10 6
#370930000000
1!
1%
1-
12
#370940000000
0!
0%
b11 *
0-
02
b11 6
#370950000000
1!
1%
1-
12
15
#370960000000
0!
0%
b100 *
0-
02
b100 6
#370970000000
1!
1%
1-
12
#370980000000
0!
0%
b101 *
0-
02
b101 6
#370990000000
1!
1%
1-
12
#371000000000
0!
0%
b110 *
0-
02
b110 6
#371010000000
1!
1%
1-
12
#371020000000
0!
0%
b111 *
0-
02
b111 6
#371030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#371040000000
0!
0%
b0 *
0-
02
b0 6
#371050000000
1!
1%
1-
12
#371060000000
0!
0%
b1 *
0-
02
b1 6
#371070000000
1!
1%
1-
12
#371080000000
0!
0%
b10 *
0-
02
b10 6
#371090000000
1!
1%
1-
12
#371100000000
0!
0%
b11 *
0-
02
b11 6
#371110000000
1!
1%
1-
12
15
#371120000000
0!
0%
b100 *
0-
02
b100 6
#371130000000
1!
1%
1-
12
#371140000000
0!
0%
b101 *
0-
02
b101 6
#371150000000
1!
1%
1-
12
#371160000000
0!
0%
b110 *
0-
02
b110 6
#371170000000
1!
1%
1-
12
#371180000000
0!
0%
b111 *
0-
02
b111 6
#371190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#371200000000
0!
0%
b0 *
0-
02
b0 6
#371210000000
1!
1%
1-
12
#371220000000
0!
0%
b1 *
0-
02
b1 6
#371230000000
1!
1%
1-
12
#371240000000
0!
0%
b10 *
0-
02
b10 6
#371250000000
1!
1%
1-
12
#371260000000
0!
0%
b11 *
0-
02
b11 6
#371270000000
1!
1%
1-
12
15
#371280000000
0!
0%
b100 *
0-
02
b100 6
#371290000000
1!
1%
1-
12
#371300000000
0!
0%
b101 *
0-
02
b101 6
#371310000000
1!
1%
1-
12
#371320000000
0!
0%
b110 *
0-
02
b110 6
#371330000000
1!
1%
1-
12
#371340000000
0!
0%
b111 *
0-
02
b111 6
#371350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#371360000000
0!
0%
b0 *
0-
02
b0 6
#371370000000
1!
1%
1-
12
#371380000000
0!
0%
b1 *
0-
02
b1 6
#371390000000
1!
1%
1-
12
#371400000000
0!
0%
b10 *
0-
02
b10 6
#371410000000
1!
1%
1-
12
#371420000000
0!
0%
b11 *
0-
02
b11 6
#371430000000
1!
1%
1-
12
15
#371440000000
0!
0%
b100 *
0-
02
b100 6
#371450000000
1!
1%
1-
12
#371460000000
0!
0%
b101 *
0-
02
b101 6
#371470000000
1!
1%
1-
12
#371480000000
0!
0%
b110 *
0-
02
b110 6
#371490000000
1!
1%
1-
12
#371500000000
0!
0%
b111 *
0-
02
b111 6
#371510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#371520000000
0!
0%
b0 *
0-
02
b0 6
#371530000000
1!
1%
1-
12
#371540000000
0!
0%
b1 *
0-
02
b1 6
#371550000000
1!
1%
1-
12
#371560000000
0!
0%
b10 *
0-
02
b10 6
#371570000000
1!
1%
1-
12
#371580000000
0!
0%
b11 *
0-
02
b11 6
#371590000000
1!
1%
1-
12
15
#371600000000
0!
0%
b100 *
0-
02
b100 6
#371610000000
1!
1%
1-
12
#371620000000
0!
0%
b101 *
0-
02
b101 6
#371630000000
1!
1%
1-
12
#371640000000
0!
0%
b110 *
0-
02
b110 6
#371650000000
1!
1%
1-
12
#371660000000
0!
0%
b111 *
0-
02
b111 6
#371670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#371680000000
0!
0%
b0 *
0-
02
b0 6
#371690000000
1!
1%
1-
12
#371700000000
0!
0%
b1 *
0-
02
b1 6
#371710000000
1!
1%
1-
12
#371720000000
0!
0%
b10 *
0-
02
b10 6
#371730000000
1!
1%
1-
12
#371740000000
0!
0%
b11 *
0-
02
b11 6
#371750000000
1!
1%
1-
12
15
#371760000000
0!
0%
b100 *
0-
02
b100 6
#371770000000
1!
1%
1-
12
#371780000000
0!
0%
b101 *
0-
02
b101 6
#371790000000
1!
1%
1-
12
#371800000000
0!
0%
b110 *
0-
02
b110 6
#371810000000
1!
1%
1-
12
#371820000000
0!
0%
b111 *
0-
02
b111 6
#371830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#371840000000
0!
0%
b0 *
0-
02
b0 6
#371850000000
1!
1%
1-
12
#371860000000
0!
0%
b1 *
0-
02
b1 6
#371870000000
1!
1%
1-
12
#371880000000
0!
0%
b10 *
0-
02
b10 6
#371890000000
1!
1%
1-
12
#371900000000
0!
0%
b11 *
0-
02
b11 6
#371910000000
1!
1%
1-
12
15
#371920000000
0!
0%
b100 *
0-
02
b100 6
#371930000000
1!
1%
1-
12
#371940000000
0!
0%
b101 *
0-
02
b101 6
#371950000000
1!
1%
1-
12
#371960000000
0!
0%
b110 *
0-
02
b110 6
#371970000000
1!
1%
1-
12
#371980000000
0!
0%
b111 *
0-
02
b111 6
#371990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#372000000000
0!
0%
b0 *
0-
02
b0 6
#372010000000
1!
1%
1-
12
#372020000000
0!
0%
b1 *
0-
02
b1 6
#372030000000
1!
1%
1-
12
#372040000000
0!
0%
b10 *
0-
02
b10 6
#372050000000
1!
1%
1-
12
#372060000000
0!
0%
b11 *
0-
02
b11 6
#372070000000
1!
1%
1-
12
15
#372080000000
0!
0%
b100 *
0-
02
b100 6
#372090000000
1!
1%
1-
12
#372100000000
0!
0%
b101 *
0-
02
b101 6
#372110000000
1!
1%
1-
12
#372120000000
0!
0%
b110 *
0-
02
b110 6
#372130000000
1!
1%
1-
12
#372140000000
0!
0%
b111 *
0-
02
b111 6
#372150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#372160000000
0!
0%
b0 *
0-
02
b0 6
#372170000000
1!
1%
1-
12
#372180000000
0!
0%
b1 *
0-
02
b1 6
#372190000000
1!
1%
1-
12
#372200000000
0!
0%
b10 *
0-
02
b10 6
#372210000000
1!
1%
1-
12
#372220000000
0!
0%
b11 *
0-
02
b11 6
#372230000000
1!
1%
1-
12
15
#372240000000
0!
0%
b100 *
0-
02
b100 6
#372250000000
1!
1%
1-
12
#372260000000
0!
0%
b101 *
0-
02
b101 6
#372270000000
1!
1%
1-
12
#372280000000
0!
0%
b110 *
0-
02
b110 6
#372290000000
1!
1%
1-
12
#372300000000
0!
0%
b111 *
0-
02
b111 6
#372310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#372320000000
0!
0%
b0 *
0-
02
b0 6
#372330000000
1!
1%
1-
12
#372340000000
0!
0%
b1 *
0-
02
b1 6
#372350000000
1!
1%
1-
12
#372360000000
0!
0%
b10 *
0-
02
b10 6
#372370000000
1!
1%
1-
12
#372380000000
0!
0%
b11 *
0-
02
b11 6
#372390000000
1!
1%
1-
12
15
#372400000000
0!
0%
b100 *
0-
02
b100 6
#372410000000
1!
1%
1-
12
#372420000000
0!
0%
b101 *
0-
02
b101 6
#372430000000
1!
1%
1-
12
#372440000000
0!
0%
b110 *
0-
02
b110 6
#372450000000
1!
1%
1-
12
#372460000000
0!
0%
b111 *
0-
02
b111 6
#372470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#372480000000
0!
0%
b0 *
0-
02
b0 6
#372490000000
1!
1%
1-
12
#372500000000
0!
0%
b1 *
0-
02
b1 6
#372510000000
1!
1%
1-
12
#372520000000
0!
0%
b10 *
0-
02
b10 6
#372530000000
1!
1%
1-
12
#372540000000
0!
0%
b11 *
0-
02
b11 6
#372550000000
1!
1%
1-
12
15
#372560000000
0!
0%
b100 *
0-
02
b100 6
#372570000000
1!
1%
1-
12
#372580000000
0!
0%
b101 *
0-
02
b101 6
#372590000000
1!
1%
1-
12
#372600000000
0!
0%
b110 *
0-
02
b110 6
#372610000000
1!
1%
1-
12
#372620000000
0!
0%
b111 *
0-
02
b111 6
#372630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#372640000000
0!
0%
b0 *
0-
02
b0 6
#372650000000
1!
1%
1-
12
#372660000000
0!
0%
b1 *
0-
02
b1 6
#372670000000
1!
1%
1-
12
#372680000000
0!
0%
b10 *
0-
02
b10 6
#372690000000
1!
1%
1-
12
#372700000000
0!
0%
b11 *
0-
02
b11 6
#372710000000
1!
1%
1-
12
15
#372720000000
0!
0%
b100 *
0-
02
b100 6
#372730000000
1!
1%
1-
12
#372740000000
0!
0%
b101 *
0-
02
b101 6
#372750000000
1!
1%
1-
12
#372760000000
0!
0%
b110 *
0-
02
b110 6
#372770000000
1!
1%
1-
12
#372780000000
0!
0%
b111 *
0-
02
b111 6
#372790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#372800000000
0!
0%
b0 *
0-
02
b0 6
#372810000000
1!
1%
1-
12
#372820000000
0!
0%
b1 *
0-
02
b1 6
#372830000000
1!
1%
1-
12
#372840000000
0!
0%
b10 *
0-
02
b10 6
#372850000000
1!
1%
1-
12
#372860000000
0!
0%
b11 *
0-
02
b11 6
#372870000000
1!
1%
1-
12
15
#372880000000
0!
0%
b100 *
0-
02
b100 6
#372890000000
1!
1%
1-
12
#372900000000
0!
0%
b101 *
0-
02
b101 6
#372910000000
1!
1%
1-
12
#372920000000
0!
0%
b110 *
0-
02
b110 6
#372930000000
1!
1%
1-
12
#372940000000
0!
0%
b111 *
0-
02
b111 6
#372950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#372960000000
0!
0%
b0 *
0-
02
b0 6
#372970000000
1!
1%
1-
12
#372980000000
0!
0%
b1 *
0-
02
b1 6
#372990000000
1!
1%
1-
12
#373000000000
0!
0%
b10 *
0-
02
b10 6
#373010000000
1!
1%
1-
12
#373020000000
0!
0%
b11 *
0-
02
b11 6
#373030000000
1!
1%
1-
12
15
#373040000000
0!
0%
b100 *
0-
02
b100 6
#373050000000
1!
1%
1-
12
#373060000000
0!
0%
b101 *
0-
02
b101 6
#373070000000
1!
1%
1-
12
#373080000000
0!
0%
b110 *
0-
02
b110 6
#373090000000
1!
1%
1-
12
#373100000000
0!
0%
b111 *
0-
02
b111 6
#373110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#373120000000
0!
0%
b0 *
0-
02
b0 6
#373130000000
1!
1%
1-
12
#373140000000
0!
0%
b1 *
0-
02
b1 6
#373150000000
1!
1%
1-
12
#373160000000
0!
0%
b10 *
0-
02
b10 6
#373170000000
1!
1%
1-
12
#373180000000
0!
0%
b11 *
0-
02
b11 6
#373190000000
1!
1%
1-
12
15
#373200000000
0!
0%
b100 *
0-
02
b100 6
#373210000000
1!
1%
1-
12
#373220000000
0!
0%
b101 *
0-
02
b101 6
#373230000000
1!
1%
1-
12
#373240000000
0!
0%
b110 *
0-
02
b110 6
#373250000000
1!
1%
1-
12
#373260000000
0!
0%
b111 *
0-
02
b111 6
#373270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#373280000000
0!
0%
b0 *
0-
02
b0 6
#373290000000
1!
1%
1-
12
#373300000000
0!
0%
b1 *
0-
02
b1 6
#373310000000
1!
1%
1-
12
#373320000000
0!
0%
b10 *
0-
02
b10 6
#373330000000
1!
1%
1-
12
#373340000000
0!
0%
b11 *
0-
02
b11 6
#373350000000
1!
1%
1-
12
15
#373360000000
0!
0%
b100 *
0-
02
b100 6
#373370000000
1!
1%
1-
12
#373380000000
0!
0%
b101 *
0-
02
b101 6
#373390000000
1!
1%
1-
12
#373400000000
0!
0%
b110 *
0-
02
b110 6
#373410000000
1!
1%
1-
12
#373420000000
0!
0%
b111 *
0-
02
b111 6
#373430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#373440000000
0!
0%
b0 *
0-
02
b0 6
#373450000000
1!
1%
1-
12
#373460000000
0!
0%
b1 *
0-
02
b1 6
#373470000000
1!
1%
1-
12
#373480000000
0!
0%
b10 *
0-
02
b10 6
#373490000000
1!
1%
1-
12
#373500000000
0!
0%
b11 *
0-
02
b11 6
#373510000000
1!
1%
1-
12
15
#373520000000
0!
0%
b100 *
0-
02
b100 6
#373530000000
1!
1%
1-
12
#373540000000
0!
0%
b101 *
0-
02
b101 6
#373550000000
1!
1%
1-
12
#373560000000
0!
0%
b110 *
0-
02
b110 6
#373570000000
1!
1%
1-
12
#373580000000
0!
0%
b111 *
0-
02
b111 6
#373590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#373600000000
0!
0%
b0 *
0-
02
b0 6
#373610000000
1!
1%
1-
12
#373620000000
0!
0%
b1 *
0-
02
b1 6
#373630000000
1!
1%
1-
12
#373640000000
0!
0%
b10 *
0-
02
b10 6
#373650000000
1!
1%
1-
12
#373660000000
0!
0%
b11 *
0-
02
b11 6
#373670000000
1!
1%
1-
12
15
#373680000000
0!
0%
b100 *
0-
02
b100 6
#373690000000
1!
1%
1-
12
#373700000000
0!
0%
b101 *
0-
02
b101 6
#373710000000
1!
1%
1-
12
#373720000000
0!
0%
b110 *
0-
02
b110 6
#373730000000
1!
1%
1-
12
#373740000000
0!
0%
b111 *
0-
02
b111 6
#373750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#373760000000
0!
0%
b0 *
0-
02
b0 6
#373770000000
1!
1%
1-
12
#373780000000
0!
0%
b1 *
0-
02
b1 6
#373790000000
1!
1%
1-
12
#373800000000
0!
0%
b10 *
0-
02
b10 6
#373810000000
1!
1%
1-
12
#373820000000
0!
0%
b11 *
0-
02
b11 6
#373830000000
1!
1%
1-
12
15
#373840000000
0!
0%
b100 *
0-
02
b100 6
#373850000000
1!
1%
1-
12
#373860000000
0!
0%
b101 *
0-
02
b101 6
#373870000000
1!
1%
1-
12
#373880000000
0!
0%
b110 *
0-
02
b110 6
#373890000000
1!
1%
1-
12
#373900000000
0!
0%
b111 *
0-
02
b111 6
#373910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#373920000000
0!
0%
b0 *
0-
02
b0 6
#373930000000
1!
1%
1-
12
#373940000000
0!
0%
b1 *
0-
02
b1 6
#373950000000
1!
1%
1-
12
#373960000000
0!
0%
b10 *
0-
02
b10 6
#373970000000
1!
1%
1-
12
#373980000000
0!
0%
b11 *
0-
02
b11 6
#373990000000
1!
1%
1-
12
15
#374000000000
0!
0%
b100 *
0-
02
b100 6
#374010000000
1!
1%
1-
12
#374020000000
0!
0%
b101 *
0-
02
b101 6
#374030000000
1!
1%
1-
12
#374040000000
0!
0%
b110 *
0-
02
b110 6
#374050000000
1!
1%
1-
12
#374060000000
0!
0%
b111 *
0-
02
b111 6
#374070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#374080000000
0!
0%
b0 *
0-
02
b0 6
#374090000000
1!
1%
1-
12
#374100000000
0!
0%
b1 *
0-
02
b1 6
#374110000000
1!
1%
1-
12
#374120000000
0!
0%
b10 *
0-
02
b10 6
#374130000000
1!
1%
1-
12
#374140000000
0!
0%
b11 *
0-
02
b11 6
#374150000000
1!
1%
1-
12
15
#374160000000
0!
0%
b100 *
0-
02
b100 6
#374170000000
1!
1%
1-
12
#374180000000
0!
0%
b101 *
0-
02
b101 6
#374190000000
1!
1%
1-
12
#374200000000
0!
0%
b110 *
0-
02
b110 6
#374210000000
1!
1%
1-
12
#374220000000
0!
0%
b111 *
0-
02
b111 6
#374230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#374240000000
0!
0%
b0 *
0-
02
b0 6
#374250000000
1!
1%
1-
12
#374260000000
0!
0%
b1 *
0-
02
b1 6
#374270000000
1!
1%
1-
12
#374280000000
0!
0%
b10 *
0-
02
b10 6
#374290000000
1!
1%
1-
12
#374300000000
0!
0%
b11 *
0-
02
b11 6
#374310000000
1!
1%
1-
12
15
#374320000000
0!
0%
b100 *
0-
02
b100 6
#374330000000
1!
1%
1-
12
#374340000000
0!
0%
b101 *
0-
02
b101 6
#374350000000
1!
1%
1-
12
#374360000000
0!
0%
b110 *
0-
02
b110 6
#374370000000
1!
1%
1-
12
#374380000000
0!
0%
b111 *
0-
02
b111 6
#374390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#374400000000
0!
0%
b0 *
0-
02
b0 6
#374410000000
1!
1%
1-
12
#374420000000
0!
0%
b1 *
0-
02
b1 6
#374430000000
1!
1%
1-
12
#374440000000
0!
0%
b10 *
0-
02
b10 6
#374450000000
1!
1%
1-
12
#374460000000
0!
0%
b11 *
0-
02
b11 6
#374470000000
1!
1%
1-
12
15
#374480000000
0!
0%
b100 *
0-
02
b100 6
#374490000000
1!
1%
1-
12
#374500000000
0!
0%
b101 *
0-
02
b101 6
#374510000000
1!
1%
1-
12
#374520000000
0!
0%
b110 *
0-
02
b110 6
#374530000000
1!
1%
1-
12
#374540000000
0!
0%
b111 *
0-
02
b111 6
#374550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#374560000000
0!
0%
b0 *
0-
02
b0 6
#374570000000
1!
1%
1-
12
#374580000000
0!
0%
b1 *
0-
02
b1 6
#374590000000
1!
1%
1-
12
#374600000000
0!
0%
b10 *
0-
02
b10 6
#374610000000
1!
1%
1-
12
#374620000000
0!
0%
b11 *
0-
02
b11 6
#374630000000
1!
1%
1-
12
15
#374640000000
0!
0%
b100 *
0-
02
b100 6
#374650000000
1!
1%
1-
12
#374660000000
0!
0%
b101 *
0-
02
b101 6
#374670000000
1!
1%
1-
12
#374680000000
0!
0%
b110 *
0-
02
b110 6
#374690000000
1!
1%
1-
12
#374700000000
0!
0%
b111 *
0-
02
b111 6
#374710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#374720000000
0!
0%
b0 *
0-
02
b0 6
#374730000000
1!
1%
1-
12
#374740000000
0!
0%
b1 *
0-
02
b1 6
#374750000000
1!
1%
1-
12
#374760000000
0!
0%
b10 *
0-
02
b10 6
#374770000000
1!
1%
1-
12
#374780000000
0!
0%
b11 *
0-
02
b11 6
#374790000000
1!
1%
1-
12
15
#374800000000
0!
0%
b100 *
0-
02
b100 6
#374810000000
1!
1%
1-
12
#374820000000
0!
0%
b101 *
0-
02
b101 6
#374830000000
1!
1%
1-
12
#374840000000
0!
0%
b110 *
0-
02
b110 6
#374850000000
1!
1%
1-
12
#374860000000
0!
0%
b111 *
0-
02
b111 6
#374870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#374880000000
0!
0%
b0 *
0-
02
b0 6
#374890000000
1!
1%
1-
12
#374900000000
0!
0%
b1 *
0-
02
b1 6
#374910000000
1!
1%
1-
12
#374920000000
0!
0%
b10 *
0-
02
b10 6
#374930000000
1!
1%
1-
12
#374940000000
0!
0%
b11 *
0-
02
b11 6
#374950000000
1!
1%
1-
12
15
#374960000000
0!
0%
b100 *
0-
02
b100 6
#374970000000
1!
1%
1-
12
#374980000000
0!
0%
b101 *
0-
02
b101 6
#374990000000
1!
1%
1-
12
#375000000000
0!
0%
b110 *
0-
02
b110 6
#375010000000
1!
1%
1-
12
#375020000000
0!
0%
b111 *
0-
02
b111 6
#375030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#375040000000
0!
0%
b0 *
0-
02
b0 6
#375050000000
1!
1%
1-
12
#375060000000
0!
0%
b1 *
0-
02
b1 6
#375070000000
1!
1%
1-
12
#375080000000
0!
0%
b10 *
0-
02
b10 6
#375090000000
1!
1%
1-
12
#375100000000
0!
0%
b11 *
0-
02
b11 6
#375110000000
1!
1%
1-
12
15
#375120000000
0!
0%
b100 *
0-
02
b100 6
#375130000000
1!
1%
1-
12
#375140000000
0!
0%
b101 *
0-
02
b101 6
#375150000000
1!
1%
1-
12
#375160000000
0!
0%
b110 *
0-
02
b110 6
#375170000000
1!
1%
1-
12
#375180000000
0!
0%
b111 *
0-
02
b111 6
#375190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#375200000000
0!
0%
b0 *
0-
02
b0 6
#375210000000
1!
1%
1-
12
#375220000000
0!
0%
b1 *
0-
02
b1 6
#375230000000
1!
1%
1-
12
#375240000000
0!
0%
b10 *
0-
02
b10 6
#375250000000
1!
1%
1-
12
#375260000000
0!
0%
b11 *
0-
02
b11 6
#375270000000
1!
1%
1-
12
15
#375280000000
0!
0%
b100 *
0-
02
b100 6
#375290000000
1!
1%
1-
12
#375300000000
0!
0%
b101 *
0-
02
b101 6
#375310000000
1!
1%
1-
12
#375320000000
0!
0%
b110 *
0-
02
b110 6
#375330000000
1!
1%
1-
12
#375340000000
0!
0%
b111 *
0-
02
b111 6
#375350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#375360000000
0!
0%
b0 *
0-
02
b0 6
#375370000000
1!
1%
1-
12
#375380000000
0!
0%
b1 *
0-
02
b1 6
#375390000000
1!
1%
1-
12
#375400000000
0!
0%
b10 *
0-
02
b10 6
#375410000000
1!
1%
1-
12
#375420000000
0!
0%
b11 *
0-
02
b11 6
#375430000000
1!
1%
1-
12
15
#375440000000
0!
0%
b100 *
0-
02
b100 6
#375450000000
1!
1%
1-
12
#375460000000
0!
0%
b101 *
0-
02
b101 6
#375470000000
1!
1%
1-
12
#375480000000
0!
0%
b110 *
0-
02
b110 6
#375490000000
1!
1%
1-
12
#375500000000
0!
0%
b111 *
0-
02
b111 6
#375510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#375520000000
0!
0%
b0 *
0-
02
b0 6
#375530000000
1!
1%
1-
12
#375540000000
0!
0%
b1 *
0-
02
b1 6
#375550000000
1!
1%
1-
12
#375560000000
0!
0%
b10 *
0-
02
b10 6
#375570000000
1!
1%
1-
12
#375580000000
0!
0%
b11 *
0-
02
b11 6
#375590000000
1!
1%
1-
12
15
#375600000000
0!
0%
b100 *
0-
02
b100 6
#375610000000
1!
1%
1-
12
#375620000000
0!
0%
b101 *
0-
02
b101 6
#375630000000
1!
1%
1-
12
#375640000000
0!
0%
b110 *
0-
02
b110 6
#375650000000
1!
1%
1-
12
#375660000000
0!
0%
b111 *
0-
02
b111 6
#375670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#375680000000
0!
0%
b0 *
0-
02
b0 6
#375690000000
1!
1%
1-
12
#375700000000
0!
0%
b1 *
0-
02
b1 6
#375710000000
1!
1%
1-
12
#375720000000
0!
0%
b10 *
0-
02
b10 6
#375730000000
1!
1%
1-
12
#375740000000
0!
0%
b11 *
0-
02
b11 6
#375750000000
1!
1%
1-
12
15
#375760000000
0!
0%
b100 *
0-
02
b100 6
#375770000000
1!
1%
1-
12
#375780000000
0!
0%
b101 *
0-
02
b101 6
#375790000000
1!
1%
1-
12
#375800000000
0!
0%
b110 *
0-
02
b110 6
#375810000000
1!
1%
1-
12
#375820000000
0!
0%
b111 *
0-
02
b111 6
#375830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#375840000000
0!
0%
b0 *
0-
02
b0 6
#375850000000
1!
1%
1-
12
#375860000000
0!
0%
b1 *
0-
02
b1 6
#375870000000
1!
1%
1-
12
#375880000000
0!
0%
b10 *
0-
02
b10 6
#375890000000
1!
1%
1-
12
#375900000000
0!
0%
b11 *
0-
02
b11 6
#375910000000
1!
1%
1-
12
15
#375920000000
0!
0%
b100 *
0-
02
b100 6
#375930000000
1!
1%
1-
12
#375940000000
0!
0%
b101 *
0-
02
b101 6
#375950000000
1!
1%
1-
12
#375960000000
0!
0%
b110 *
0-
02
b110 6
#375970000000
1!
1%
1-
12
#375980000000
0!
0%
b111 *
0-
02
b111 6
#375990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#376000000000
0!
0%
b0 *
0-
02
b0 6
#376010000000
1!
1%
1-
12
#376020000000
0!
0%
b1 *
0-
02
b1 6
#376030000000
1!
1%
1-
12
#376040000000
0!
0%
b10 *
0-
02
b10 6
#376050000000
1!
1%
1-
12
#376060000000
0!
0%
b11 *
0-
02
b11 6
#376070000000
1!
1%
1-
12
15
#376080000000
0!
0%
b100 *
0-
02
b100 6
#376090000000
1!
1%
1-
12
#376100000000
0!
0%
b101 *
0-
02
b101 6
#376110000000
1!
1%
1-
12
#376120000000
0!
0%
b110 *
0-
02
b110 6
#376130000000
1!
1%
1-
12
#376140000000
0!
0%
b111 *
0-
02
b111 6
#376150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#376160000000
0!
0%
b0 *
0-
02
b0 6
#376170000000
1!
1%
1-
12
#376180000000
0!
0%
b1 *
0-
02
b1 6
#376190000000
1!
1%
1-
12
#376200000000
0!
0%
b10 *
0-
02
b10 6
#376210000000
1!
1%
1-
12
#376220000000
0!
0%
b11 *
0-
02
b11 6
#376230000000
1!
1%
1-
12
15
#376240000000
0!
0%
b100 *
0-
02
b100 6
#376250000000
1!
1%
1-
12
#376260000000
0!
0%
b101 *
0-
02
b101 6
#376270000000
1!
1%
1-
12
#376280000000
0!
0%
b110 *
0-
02
b110 6
#376290000000
1!
1%
1-
12
#376300000000
0!
0%
b111 *
0-
02
b111 6
#376310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#376320000000
0!
0%
b0 *
0-
02
b0 6
#376330000000
1!
1%
1-
12
#376340000000
0!
0%
b1 *
0-
02
b1 6
#376350000000
1!
1%
1-
12
#376360000000
0!
0%
b10 *
0-
02
b10 6
#376370000000
1!
1%
1-
12
#376380000000
0!
0%
b11 *
0-
02
b11 6
#376390000000
1!
1%
1-
12
15
#376400000000
0!
0%
b100 *
0-
02
b100 6
#376410000000
1!
1%
1-
12
#376420000000
0!
0%
b101 *
0-
02
b101 6
#376430000000
1!
1%
1-
12
#376440000000
0!
0%
b110 *
0-
02
b110 6
#376450000000
1!
1%
1-
12
#376460000000
0!
0%
b111 *
0-
02
b111 6
#376470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#376480000000
0!
0%
b0 *
0-
02
b0 6
#376490000000
1!
1%
1-
12
#376500000000
0!
0%
b1 *
0-
02
b1 6
#376510000000
1!
1%
1-
12
#376520000000
0!
0%
b10 *
0-
02
b10 6
#376530000000
1!
1%
1-
12
#376540000000
0!
0%
b11 *
0-
02
b11 6
#376550000000
1!
1%
1-
12
15
#376560000000
0!
0%
b100 *
0-
02
b100 6
#376570000000
1!
1%
1-
12
#376580000000
0!
0%
b101 *
0-
02
b101 6
#376590000000
1!
1%
1-
12
#376600000000
0!
0%
b110 *
0-
02
b110 6
#376610000000
1!
1%
1-
12
#376620000000
0!
0%
b111 *
0-
02
b111 6
#376630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#376640000000
0!
0%
b0 *
0-
02
b0 6
#376650000000
1!
1%
1-
12
#376660000000
0!
0%
b1 *
0-
02
b1 6
#376670000000
1!
1%
1-
12
#376680000000
0!
0%
b10 *
0-
02
b10 6
#376690000000
1!
1%
1-
12
#376700000000
0!
0%
b11 *
0-
02
b11 6
#376710000000
1!
1%
1-
12
15
#376720000000
0!
0%
b100 *
0-
02
b100 6
#376730000000
1!
1%
1-
12
#376740000000
0!
0%
b101 *
0-
02
b101 6
#376750000000
1!
1%
1-
12
#376760000000
0!
0%
b110 *
0-
02
b110 6
#376770000000
1!
1%
1-
12
#376780000000
0!
0%
b111 *
0-
02
b111 6
#376790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#376800000000
0!
0%
b0 *
0-
02
b0 6
#376810000000
1!
1%
1-
12
#376820000000
0!
0%
b1 *
0-
02
b1 6
#376830000000
1!
1%
1-
12
#376840000000
0!
0%
b10 *
0-
02
b10 6
#376850000000
1!
1%
1-
12
#376860000000
0!
0%
b11 *
0-
02
b11 6
#376870000000
1!
1%
1-
12
15
#376880000000
0!
0%
b100 *
0-
02
b100 6
#376890000000
1!
1%
1-
12
#376900000000
0!
0%
b101 *
0-
02
b101 6
#376910000000
1!
1%
1-
12
#376920000000
0!
0%
b110 *
0-
02
b110 6
#376930000000
1!
1%
1-
12
#376940000000
0!
0%
b111 *
0-
02
b111 6
#376950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#376960000000
0!
0%
b0 *
0-
02
b0 6
#376970000000
1!
1%
1-
12
#376980000000
0!
0%
b1 *
0-
02
b1 6
#376990000000
1!
1%
1-
12
#377000000000
0!
0%
b10 *
0-
02
b10 6
#377010000000
1!
1%
1-
12
#377020000000
0!
0%
b11 *
0-
02
b11 6
#377030000000
1!
1%
1-
12
15
#377040000000
0!
0%
b100 *
0-
02
b100 6
#377050000000
1!
1%
1-
12
#377060000000
0!
0%
b101 *
0-
02
b101 6
#377070000000
1!
1%
1-
12
#377080000000
0!
0%
b110 *
0-
02
b110 6
#377090000000
1!
1%
1-
12
#377100000000
0!
0%
b111 *
0-
02
b111 6
#377110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#377120000000
0!
0%
b0 *
0-
02
b0 6
#377130000000
1!
1%
1-
12
#377140000000
0!
0%
b1 *
0-
02
b1 6
#377150000000
1!
1%
1-
12
#377160000000
0!
0%
b10 *
0-
02
b10 6
#377170000000
1!
1%
1-
12
#377180000000
0!
0%
b11 *
0-
02
b11 6
#377190000000
1!
1%
1-
12
15
#377200000000
0!
0%
b100 *
0-
02
b100 6
#377210000000
1!
1%
1-
12
#377220000000
0!
0%
b101 *
0-
02
b101 6
#377230000000
1!
1%
1-
12
#377240000000
0!
0%
b110 *
0-
02
b110 6
#377250000000
1!
1%
1-
12
#377260000000
0!
0%
b111 *
0-
02
b111 6
#377270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#377280000000
0!
0%
b0 *
0-
02
b0 6
#377290000000
1!
1%
1-
12
#377300000000
0!
0%
b1 *
0-
02
b1 6
#377310000000
1!
1%
1-
12
#377320000000
0!
0%
b10 *
0-
02
b10 6
#377330000000
1!
1%
1-
12
#377340000000
0!
0%
b11 *
0-
02
b11 6
#377350000000
1!
1%
1-
12
15
#377360000000
0!
0%
b100 *
0-
02
b100 6
#377370000000
1!
1%
1-
12
#377380000000
0!
0%
b101 *
0-
02
b101 6
#377390000000
1!
1%
1-
12
#377400000000
0!
0%
b110 *
0-
02
b110 6
#377410000000
1!
1%
1-
12
#377420000000
0!
0%
b111 *
0-
02
b111 6
#377430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#377440000000
0!
0%
b0 *
0-
02
b0 6
#377450000000
1!
1%
1-
12
#377460000000
0!
0%
b1 *
0-
02
b1 6
#377470000000
1!
1%
1-
12
#377480000000
0!
0%
b10 *
0-
02
b10 6
#377490000000
1!
1%
1-
12
#377500000000
0!
0%
b11 *
0-
02
b11 6
#377510000000
1!
1%
1-
12
15
#377520000000
0!
0%
b100 *
0-
02
b100 6
#377530000000
1!
1%
1-
12
#377540000000
0!
0%
b101 *
0-
02
b101 6
#377550000000
1!
1%
1-
12
#377560000000
0!
0%
b110 *
0-
02
b110 6
#377570000000
1!
1%
1-
12
#377580000000
0!
0%
b111 *
0-
02
b111 6
#377590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#377600000000
0!
0%
b0 *
0-
02
b0 6
#377610000000
1!
1%
1-
12
#377620000000
0!
0%
b1 *
0-
02
b1 6
#377630000000
1!
1%
1-
12
#377640000000
0!
0%
b10 *
0-
02
b10 6
#377650000000
1!
1%
1-
12
#377660000000
0!
0%
b11 *
0-
02
b11 6
#377670000000
1!
1%
1-
12
15
#377680000000
0!
0%
b100 *
0-
02
b100 6
#377690000000
1!
1%
1-
12
#377700000000
0!
0%
b101 *
0-
02
b101 6
#377710000000
1!
1%
1-
12
#377720000000
0!
0%
b110 *
0-
02
b110 6
#377730000000
1!
1%
1-
12
#377740000000
0!
0%
b111 *
0-
02
b111 6
#377750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#377760000000
0!
0%
b0 *
0-
02
b0 6
#377770000000
1!
1%
1-
12
#377780000000
0!
0%
b1 *
0-
02
b1 6
#377790000000
1!
1%
1-
12
#377800000000
0!
0%
b10 *
0-
02
b10 6
#377810000000
1!
1%
1-
12
#377820000000
0!
0%
b11 *
0-
02
b11 6
#377830000000
1!
1%
1-
12
15
#377840000000
0!
0%
b100 *
0-
02
b100 6
#377850000000
1!
1%
1-
12
#377860000000
0!
0%
b101 *
0-
02
b101 6
#377870000000
1!
1%
1-
12
#377880000000
0!
0%
b110 *
0-
02
b110 6
#377890000000
1!
1%
1-
12
#377900000000
0!
0%
b111 *
0-
02
b111 6
#377910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#377920000000
0!
0%
b0 *
0-
02
b0 6
#377930000000
1!
1%
1-
12
#377940000000
0!
0%
b1 *
0-
02
b1 6
#377950000000
1!
1%
1-
12
#377960000000
0!
0%
b10 *
0-
02
b10 6
#377970000000
1!
1%
1-
12
#377980000000
0!
0%
b11 *
0-
02
b11 6
#377990000000
1!
1%
1-
12
15
#378000000000
0!
0%
b100 *
0-
02
b100 6
#378010000000
1!
1%
1-
12
#378020000000
0!
0%
b101 *
0-
02
b101 6
#378030000000
1!
1%
1-
12
#378040000000
0!
0%
b110 *
0-
02
b110 6
#378050000000
1!
1%
1-
12
#378060000000
0!
0%
b111 *
0-
02
b111 6
#378070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#378080000000
0!
0%
b0 *
0-
02
b0 6
#378090000000
1!
1%
1-
12
#378100000000
0!
0%
b1 *
0-
02
b1 6
#378110000000
1!
1%
1-
12
#378120000000
0!
0%
b10 *
0-
02
b10 6
#378130000000
1!
1%
1-
12
#378140000000
0!
0%
b11 *
0-
02
b11 6
#378150000000
1!
1%
1-
12
15
#378160000000
0!
0%
b100 *
0-
02
b100 6
#378170000000
1!
1%
1-
12
#378180000000
0!
0%
b101 *
0-
02
b101 6
#378190000000
1!
1%
1-
12
#378200000000
0!
0%
b110 *
0-
02
b110 6
#378210000000
1!
1%
1-
12
#378220000000
0!
0%
b111 *
0-
02
b111 6
#378230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#378240000000
0!
0%
b0 *
0-
02
b0 6
#378250000000
1!
1%
1-
12
#378260000000
0!
0%
b1 *
0-
02
b1 6
#378270000000
1!
1%
1-
12
#378280000000
0!
0%
b10 *
0-
02
b10 6
#378290000000
1!
1%
1-
12
#378300000000
0!
0%
b11 *
0-
02
b11 6
#378310000000
1!
1%
1-
12
15
#378320000000
0!
0%
b100 *
0-
02
b100 6
#378330000000
1!
1%
1-
12
#378340000000
0!
0%
b101 *
0-
02
b101 6
#378350000000
1!
1%
1-
12
#378360000000
0!
0%
b110 *
0-
02
b110 6
#378370000000
1!
1%
1-
12
#378380000000
0!
0%
b111 *
0-
02
b111 6
#378390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#378400000000
0!
0%
b0 *
0-
02
b0 6
#378410000000
1!
1%
1-
12
#378420000000
0!
0%
b1 *
0-
02
b1 6
#378430000000
1!
1%
1-
12
#378440000000
0!
0%
b10 *
0-
02
b10 6
#378450000000
1!
1%
1-
12
#378460000000
0!
0%
b11 *
0-
02
b11 6
#378470000000
1!
1%
1-
12
15
#378480000000
0!
0%
b100 *
0-
02
b100 6
#378490000000
1!
1%
1-
12
#378500000000
0!
0%
b101 *
0-
02
b101 6
#378510000000
1!
1%
1-
12
#378520000000
0!
0%
b110 *
0-
02
b110 6
#378530000000
1!
1%
1-
12
#378540000000
0!
0%
b111 *
0-
02
b111 6
#378550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#378560000000
0!
0%
b0 *
0-
02
b0 6
#378570000000
1!
1%
1-
12
#378580000000
0!
0%
b1 *
0-
02
b1 6
#378590000000
1!
1%
1-
12
#378600000000
0!
0%
b10 *
0-
02
b10 6
#378610000000
1!
1%
1-
12
#378620000000
0!
0%
b11 *
0-
02
b11 6
#378630000000
1!
1%
1-
12
15
#378640000000
0!
0%
b100 *
0-
02
b100 6
#378650000000
1!
1%
1-
12
#378660000000
0!
0%
b101 *
0-
02
b101 6
#378670000000
1!
1%
1-
12
#378680000000
0!
0%
b110 *
0-
02
b110 6
#378690000000
1!
1%
1-
12
#378700000000
0!
0%
b111 *
0-
02
b111 6
#378710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#378720000000
0!
0%
b0 *
0-
02
b0 6
#378730000000
1!
1%
1-
12
#378740000000
0!
0%
b1 *
0-
02
b1 6
#378750000000
1!
1%
1-
12
#378760000000
0!
0%
b10 *
0-
02
b10 6
#378770000000
1!
1%
1-
12
#378780000000
0!
0%
b11 *
0-
02
b11 6
#378790000000
1!
1%
1-
12
15
#378800000000
0!
0%
b100 *
0-
02
b100 6
#378810000000
1!
1%
1-
12
#378820000000
0!
0%
b101 *
0-
02
b101 6
#378830000000
1!
1%
1-
12
#378840000000
0!
0%
b110 *
0-
02
b110 6
#378850000000
1!
1%
1-
12
#378860000000
0!
0%
b111 *
0-
02
b111 6
#378870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#378880000000
0!
0%
b0 *
0-
02
b0 6
#378890000000
1!
1%
1-
12
#378900000000
0!
0%
b1 *
0-
02
b1 6
#378910000000
1!
1%
1-
12
#378920000000
0!
0%
b10 *
0-
02
b10 6
#378930000000
1!
1%
1-
12
#378940000000
0!
0%
b11 *
0-
02
b11 6
#378950000000
1!
1%
1-
12
15
#378960000000
0!
0%
b100 *
0-
02
b100 6
#378970000000
1!
1%
1-
12
#378980000000
0!
0%
b101 *
0-
02
b101 6
#378990000000
1!
1%
1-
12
#379000000000
0!
0%
b110 *
0-
02
b110 6
#379010000000
1!
1%
1-
12
#379020000000
0!
0%
b111 *
0-
02
b111 6
#379030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#379040000000
0!
0%
b0 *
0-
02
b0 6
#379050000000
1!
1%
1-
12
#379060000000
0!
0%
b1 *
0-
02
b1 6
#379070000000
1!
1%
1-
12
#379080000000
0!
0%
b10 *
0-
02
b10 6
#379090000000
1!
1%
1-
12
#379100000000
0!
0%
b11 *
0-
02
b11 6
#379110000000
1!
1%
1-
12
15
#379120000000
0!
0%
b100 *
0-
02
b100 6
#379130000000
1!
1%
1-
12
#379140000000
0!
0%
b101 *
0-
02
b101 6
#379150000000
1!
1%
1-
12
#379160000000
0!
0%
b110 *
0-
02
b110 6
#379170000000
1!
1%
1-
12
#379180000000
0!
0%
b111 *
0-
02
b111 6
#379190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#379200000000
0!
0%
b0 *
0-
02
b0 6
#379210000000
1!
1%
1-
12
#379220000000
0!
0%
b1 *
0-
02
b1 6
#379230000000
1!
1%
1-
12
#379240000000
0!
0%
b10 *
0-
02
b10 6
#379250000000
1!
1%
1-
12
#379260000000
0!
0%
b11 *
0-
02
b11 6
#379270000000
1!
1%
1-
12
15
#379280000000
0!
0%
b100 *
0-
02
b100 6
#379290000000
1!
1%
1-
12
#379300000000
0!
0%
b101 *
0-
02
b101 6
#379310000000
1!
1%
1-
12
#379320000000
0!
0%
b110 *
0-
02
b110 6
#379330000000
1!
1%
1-
12
#379340000000
0!
0%
b111 *
0-
02
b111 6
#379350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#379360000000
0!
0%
b0 *
0-
02
b0 6
#379370000000
1!
1%
1-
12
#379380000000
0!
0%
b1 *
0-
02
b1 6
#379390000000
1!
1%
1-
12
#379400000000
0!
0%
b10 *
0-
02
b10 6
#379410000000
1!
1%
1-
12
#379420000000
0!
0%
b11 *
0-
02
b11 6
#379430000000
1!
1%
1-
12
15
#379440000000
0!
0%
b100 *
0-
02
b100 6
#379450000000
1!
1%
1-
12
#379460000000
0!
0%
b101 *
0-
02
b101 6
#379470000000
1!
1%
1-
12
#379480000000
0!
0%
b110 *
0-
02
b110 6
#379490000000
1!
1%
1-
12
#379500000000
0!
0%
b111 *
0-
02
b111 6
#379510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#379520000000
0!
0%
b0 *
0-
02
b0 6
#379530000000
1!
1%
1-
12
#379540000000
0!
0%
b1 *
0-
02
b1 6
#379550000000
1!
1%
1-
12
#379560000000
0!
0%
b10 *
0-
02
b10 6
#379570000000
1!
1%
1-
12
#379580000000
0!
0%
b11 *
0-
02
b11 6
#379590000000
1!
1%
1-
12
15
#379600000000
0!
0%
b100 *
0-
02
b100 6
#379610000000
1!
1%
1-
12
#379620000000
0!
0%
b101 *
0-
02
b101 6
#379630000000
1!
1%
1-
12
#379640000000
0!
0%
b110 *
0-
02
b110 6
#379650000000
1!
1%
1-
12
#379660000000
0!
0%
b111 *
0-
02
b111 6
#379670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#379680000000
0!
0%
b0 *
0-
02
b0 6
#379690000000
1!
1%
1-
12
#379700000000
0!
0%
b1 *
0-
02
b1 6
#379710000000
1!
1%
1-
12
#379720000000
0!
0%
b10 *
0-
02
b10 6
#379730000000
1!
1%
1-
12
#379740000000
0!
0%
b11 *
0-
02
b11 6
#379750000000
1!
1%
1-
12
15
#379760000000
0!
0%
b100 *
0-
02
b100 6
#379770000000
1!
1%
1-
12
#379780000000
0!
0%
b101 *
0-
02
b101 6
#379790000000
1!
1%
1-
12
#379800000000
0!
0%
b110 *
0-
02
b110 6
#379810000000
1!
1%
1-
12
#379820000000
0!
0%
b111 *
0-
02
b111 6
#379830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#379840000000
0!
0%
b0 *
0-
02
b0 6
#379850000000
1!
1%
1-
12
#379860000000
0!
0%
b1 *
0-
02
b1 6
#379870000000
1!
1%
1-
12
#379880000000
0!
0%
b10 *
0-
02
b10 6
#379890000000
1!
1%
1-
12
#379900000000
0!
0%
b11 *
0-
02
b11 6
#379910000000
1!
1%
1-
12
15
#379920000000
0!
0%
b100 *
0-
02
b100 6
#379930000000
1!
1%
1-
12
#379940000000
0!
0%
b101 *
0-
02
b101 6
#379950000000
1!
1%
1-
12
#379960000000
0!
0%
b110 *
0-
02
b110 6
#379970000000
1!
1%
1-
12
#379980000000
0!
0%
b111 *
0-
02
b111 6
#379990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#380000000000
0!
0%
b0 *
0-
02
b0 6
#380010000000
1!
1%
1-
12
#380020000000
0!
0%
b1 *
0-
02
b1 6
#380030000000
1!
1%
1-
12
#380040000000
0!
0%
b10 *
0-
02
b10 6
#380050000000
1!
1%
1-
12
#380060000000
0!
0%
b11 *
0-
02
b11 6
#380070000000
1!
1%
1-
12
15
#380080000000
0!
0%
b100 *
0-
02
b100 6
#380090000000
1!
1%
1-
12
#380100000000
0!
0%
b101 *
0-
02
b101 6
#380110000000
1!
1%
1-
12
#380120000000
0!
0%
b110 *
0-
02
b110 6
#380130000000
1!
1%
1-
12
#380140000000
0!
0%
b111 *
0-
02
b111 6
#380150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#380160000000
0!
0%
b0 *
0-
02
b0 6
#380170000000
1!
1%
1-
12
#380180000000
0!
0%
b1 *
0-
02
b1 6
#380190000000
1!
1%
1-
12
#380200000000
0!
0%
b10 *
0-
02
b10 6
#380210000000
1!
1%
1-
12
#380220000000
0!
0%
b11 *
0-
02
b11 6
#380230000000
1!
1%
1-
12
15
#380240000000
0!
0%
b100 *
0-
02
b100 6
#380250000000
1!
1%
1-
12
#380260000000
0!
0%
b101 *
0-
02
b101 6
#380270000000
1!
1%
1-
12
#380280000000
0!
0%
b110 *
0-
02
b110 6
#380290000000
1!
1%
1-
12
#380300000000
0!
0%
b111 *
0-
02
b111 6
#380310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#380320000000
0!
0%
b0 *
0-
02
b0 6
#380330000000
1!
1%
1-
12
#380340000000
0!
0%
b1 *
0-
02
b1 6
#380350000000
1!
1%
1-
12
#380360000000
0!
0%
b10 *
0-
02
b10 6
#380370000000
1!
1%
1-
12
#380380000000
0!
0%
b11 *
0-
02
b11 6
#380390000000
1!
1%
1-
12
15
#380400000000
0!
0%
b100 *
0-
02
b100 6
#380410000000
1!
1%
1-
12
#380420000000
0!
0%
b101 *
0-
02
b101 6
#380430000000
1!
1%
1-
12
#380440000000
0!
0%
b110 *
0-
02
b110 6
#380450000000
1!
1%
1-
12
#380460000000
0!
0%
b111 *
0-
02
b111 6
#380470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#380480000000
0!
0%
b0 *
0-
02
b0 6
#380490000000
1!
1%
1-
12
#380500000000
0!
0%
b1 *
0-
02
b1 6
#380510000000
1!
1%
1-
12
#380520000000
0!
0%
b10 *
0-
02
b10 6
#380530000000
1!
1%
1-
12
#380540000000
0!
0%
b11 *
0-
02
b11 6
#380550000000
1!
1%
1-
12
15
#380560000000
0!
0%
b100 *
0-
02
b100 6
#380570000000
1!
1%
1-
12
#380580000000
0!
0%
b101 *
0-
02
b101 6
#380590000000
1!
1%
1-
12
#380600000000
0!
0%
b110 *
0-
02
b110 6
#380610000000
1!
1%
1-
12
#380620000000
0!
0%
b111 *
0-
02
b111 6
#380630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#380640000000
0!
0%
b0 *
0-
02
b0 6
#380650000000
1!
1%
1-
12
#380660000000
0!
0%
b1 *
0-
02
b1 6
#380670000000
1!
1%
1-
12
#380680000000
0!
0%
b10 *
0-
02
b10 6
#380690000000
1!
1%
1-
12
#380700000000
0!
0%
b11 *
0-
02
b11 6
#380710000000
1!
1%
1-
12
15
#380720000000
0!
0%
b100 *
0-
02
b100 6
#380730000000
1!
1%
1-
12
#380740000000
0!
0%
b101 *
0-
02
b101 6
#380750000000
1!
1%
1-
12
#380760000000
0!
0%
b110 *
0-
02
b110 6
#380770000000
1!
1%
1-
12
#380780000000
0!
0%
b111 *
0-
02
b111 6
#380790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#380800000000
0!
0%
b0 *
0-
02
b0 6
#380810000000
1!
1%
1-
12
#380820000000
0!
0%
b1 *
0-
02
b1 6
#380830000000
1!
1%
1-
12
#380840000000
0!
0%
b10 *
0-
02
b10 6
#380850000000
1!
1%
1-
12
#380860000000
0!
0%
b11 *
0-
02
b11 6
#380870000000
1!
1%
1-
12
15
#380880000000
0!
0%
b100 *
0-
02
b100 6
#380890000000
1!
1%
1-
12
#380900000000
0!
0%
b101 *
0-
02
b101 6
#380910000000
1!
1%
1-
12
#380920000000
0!
0%
b110 *
0-
02
b110 6
#380930000000
1!
1%
1-
12
#380940000000
0!
0%
b111 *
0-
02
b111 6
#380950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#380960000000
0!
0%
b0 *
0-
02
b0 6
#380970000000
1!
1%
1-
12
#380980000000
0!
0%
b1 *
0-
02
b1 6
#380990000000
1!
1%
1-
12
#381000000000
0!
0%
b10 *
0-
02
b10 6
#381010000000
1!
1%
1-
12
#381020000000
0!
0%
b11 *
0-
02
b11 6
#381030000000
1!
1%
1-
12
15
#381040000000
0!
0%
b100 *
0-
02
b100 6
#381050000000
1!
1%
1-
12
#381060000000
0!
0%
b101 *
0-
02
b101 6
#381070000000
1!
1%
1-
12
#381080000000
0!
0%
b110 *
0-
02
b110 6
#381090000000
1!
1%
1-
12
#381100000000
0!
0%
b111 *
0-
02
b111 6
#381110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#381120000000
0!
0%
b0 *
0-
02
b0 6
#381130000000
1!
1%
1-
12
#381140000000
0!
0%
b1 *
0-
02
b1 6
#381150000000
1!
1%
1-
12
#381160000000
0!
0%
b10 *
0-
02
b10 6
#381170000000
1!
1%
1-
12
#381180000000
0!
0%
b11 *
0-
02
b11 6
#381190000000
1!
1%
1-
12
15
#381200000000
0!
0%
b100 *
0-
02
b100 6
#381210000000
1!
1%
1-
12
#381220000000
0!
0%
b101 *
0-
02
b101 6
#381230000000
1!
1%
1-
12
#381240000000
0!
0%
b110 *
0-
02
b110 6
#381250000000
1!
1%
1-
12
#381260000000
0!
0%
b111 *
0-
02
b111 6
#381270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#381280000000
0!
0%
b0 *
0-
02
b0 6
#381290000000
1!
1%
1-
12
#381300000000
0!
0%
b1 *
0-
02
b1 6
#381310000000
1!
1%
1-
12
#381320000000
0!
0%
b10 *
0-
02
b10 6
#381330000000
1!
1%
1-
12
#381340000000
0!
0%
b11 *
0-
02
b11 6
#381350000000
1!
1%
1-
12
15
#381360000000
0!
0%
b100 *
0-
02
b100 6
#381370000000
1!
1%
1-
12
#381380000000
0!
0%
b101 *
0-
02
b101 6
#381390000000
1!
1%
1-
12
#381400000000
0!
0%
b110 *
0-
02
b110 6
#381410000000
1!
1%
1-
12
#381420000000
0!
0%
b111 *
0-
02
b111 6
#381430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#381440000000
0!
0%
b0 *
0-
02
b0 6
#381450000000
1!
1%
1-
12
#381460000000
0!
0%
b1 *
0-
02
b1 6
#381470000000
1!
1%
1-
12
#381480000000
0!
0%
b10 *
0-
02
b10 6
#381490000000
1!
1%
1-
12
#381500000000
0!
0%
b11 *
0-
02
b11 6
#381510000000
1!
1%
1-
12
15
#381520000000
0!
0%
b100 *
0-
02
b100 6
#381530000000
1!
1%
1-
12
#381540000000
0!
0%
b101 *
0-
02
b101 6
#381550000000
1!
1%
1-
12
#381560000000
0!
0%
b110 *
0-
02
b110 6
#381570000000
1!
1%
1-
12
#381580000000
0!
0%
b111 *
0-
02
b111 6
#381590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#381600000000
0!
0%
b0 *
0-
02
b0 6
#381610000000
1!
1%
1-
12
#381620000000
0!
0%
b1 *
0-
02
b1 6
#381630000000
1!
1%
1-
12
#381640000000
0!
0%
b10 *
0-
02
b10 6
#381650000000
1!
1%
1-
12
#381660000000
0!
0%
b11 *
0-
02
b11 6
#381670000000
1!
1%
1-
12
15
#381680000000
0!
0%
b100 *
0-
02
b100 6
#381690000000
1!
1%
1-
12
#381700000000
0!
0%
b101 *
0-
02
b101 6
#381710000000
1!
1%
1-
12
#381720000000
0!
0%
b110 *
0-
02
b110 6
#381730000000
1!
1%
1-
12
#381740000000
0!
0%
b111 *
0-
02
b111 6
#381750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#381760000000
0!
0%
b0 *
0-
02
b0 6
#381770000000
1!
1%
1-
12
#381780000000
0!
0%
b1 *
0-
02
b1 6
#381790000000
1!
1%
1-
12
#381800000000
0!
0%
b10 *
0-
02
b10 6
#381810000000
1!
1%
1-
12
#381820000000
0!
0%
b11 *
0-
02
b11 6
#381830000000
1!
1%
1-
12
15
#381840000000
0!
0%
b100 *
0-
02
b100 6
#381850000000
1!
1%
1-
12
#381860000000
0!
0%
b101 *
0-
02
b101 6
#381870000000
1!
1%
1-
12
#381880000000
0!
0%
b110 *
0-
02
b110 6
#381890000000
1!
1%
1-
12
#381900000000
0!
0%
b111 *
0-
02
b111 6
#381910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#381920000000
0!
0%
b0 *
0-
02
b0 6
#381930000000
1!
1%
1-
12
#381940000000
0!
0%
b1 *
0-
02
b1 6
#381950000000
1!
1%
1-
12
#381960000000
0!
0%
b10 *
0-
02
b10 6
#381970000000
1!
1%
1-
12
#381980000000
0!
0%
b11 *
0-
02
b11 6
#381990000000
1!
1%
1-
12
15
#382000000000
0!
0%
b100 *
0-
02
b100 6
#382010000000
1!
1%
1-
12
#382020000000
0!
0%
b101 *
0-
02
b101 6
#382030000000
1!
1%
1-
12
#382040000000
0!
0%
b110 *
0-
02
b110 6
#382050000000
1!
1%
1-
12
#382060000000
0!
0%
b111 *
0-
02
b111 6
#382070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#382080000000
0!
0%
b0 *
0-
02
b0 6
#382090000000
1!
1%
1-
12
#382100000000
0!
0%
b1 *
0-
02
b1 6
#382110000000
1!
1%
1-
12
#382120000000
0!
0%
b10 *
0-
02
b10 6
#382130000000
1!
1%
1-
12
#382140000000
0!
0%
b11 *
0-
02
b11 6
#382150000000
1!
1%
1-
12
15
#382160000000
0!
0%
b100 *
0-
02
b100 6
#382170000000
1!
1%
1-
12
#382180000000
0!
0%
b101 *
0-
02
b101 6
#382190000000
1!
1%
1-
12
#382200000000
0!
0%
b110 *
0-
02
b110 6
#382210000000
1!
1%
1-
12
#382220000000
0!
0%
b111 *
0-
02
b111 6
#382230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#382240000000
0!
0%
b0 *
0-
02
b0 6
#382250000000
1!
1%
1-
12
#382260000000
0!
0%
b1 *
0-
02
b1 6
#382270000000
1!
1%
1-
12
#382280000000
0!
0%
b10 *
0-
02
b10 6
#382290000000
1!
1%
1-
12
#382300000000
0!
0%
b11 *
0-
02
b11 6
#382310000000
1!
1%
1-
12
15
#382320000000
0!
0%
b100 *
0-
02
b100 6
#382330000000
1!
1%
1-
12
#382340000000
0!
0%
b101 *
0-
02
b101 6
#382350000000
1!
1%
1-
12
#382360000000
0!
0%
b110 *
0-
02
b110 6
#382370000000
1!
1%
1-
12
#382380000000
0!
0%
b111 *
0-
02
b111 6
#382390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#382400000000
0!
0%
b0 *
0-
02
b0 6
#382410000000
1!
1%
1-
12
#382420000000
0!
0%
b1 *
0-
02
b1 6
#382430000000
1!
1%
1-
12
#382440000000
0!
0%
b10 *
0-
02
b10 6
#382450000000
1!
1%
1-
12
#382460000000
0!
0%
b11 *
0-
02
b11 6
#382470000000
1!
1%
1-
12
15
#382480000000
0!
0%
b100 *
0-
02
b100 6
#382490000000
1!
1%
1-
12
#382500000000
0!
0%
b101 *
0-
02
b101 6
#382510000000
1!
1%
1-
12
#382520000000
0!
0%
b110 *
0-
02
b110 6
#382530000000
1!
1%
1-
12
#382540000000
0!
0%
b111 *
0-
02
b111 6
#382550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#382560000000
0!
0%
b0 *
0-
02
b0 6
#382570000000
1!
1%
1-
12
#382580000000
0!
0%
b1 *
0-
02
b1 6
#382590000000
1!
1%
1-
12
#382600000000
0!
0%
b10 *
0-
02
b10 6
#382610000000
1!
1%
1-
12
#382620000000
0!
0%
b11 *
0-
02
b11 6
#382630000000
1!
1%
1-
12
15
#382640000000
0!
0%
b100 *
0-
02
b100 6
#382650000000
1!
1%
1-
12
#382660000000
0!
0%
b101 *
0-
02
b101 6
#382670000000
1!
1%
1-
12
#382680000000
0!
0%
b110 *
0-
02
b110 6
#382690000000
1!
1%
1-
12
#382700000000
0!
0%
b111 *
0-
02
b111 6
#382710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#382720000000
0!
0%
b0 *
0-
02
b0 6
#382730000000
1!
1%
1-
12
#382740000000
0!
0%
b1 *
0-
02
b1 6
#382750000000
1!
1%
1-
12
#382760000000
0!
0%
b10 *
0-
02
b10 6
#382770000000
1!
1%
1-
12
#382780000000
0!
0%
b11 *
0-
02
b11 6
#382790000000
1!
1%
1-
12
15
#382800000000
0!
0%
b100 *
0-
02
b100 6
#382810000000
1!
1%
1-
12
#382820000000
0!
0%
b101 *
0-
02
b101 6
#382830000000
1!
1%
1-
12
#382840000000
0!
0%
b110 *
0-
02
b110 6
#382850000000
1!
1%
1-
12
#382860000000
0!
0%
b111 *
0-
02
b111 6
#382870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#382880000000
0!
0%
b0 *
0-
02
b0 6
#382890000000
1!
1%
1-
12
#382900000000
0!
0%
b1 *
0-
02
b1 6
#382910000000
1!
1%
1-
12
#382920000000
0!
0%
b10 *
0-
02
b10 6
#382930000000
1!
1%
1-
12
#382940000000
0!
0%
b11 *
0-
02
b11 6
#382950000000
1!
1%
1-
12
15
#382960000000
0!
0%
b100 *
0-
02
b100 6
#382970000000
1!
1%
1-
12
#382980000000
0!
0%
b101 *
0-
02
b101 6
#382990000000
1!
1%
1-
12
#383000000000
0!
0%
b110 *
0-
02
b110 6
#383010000000
1!
1%
1-
12
#383020000000
0!
0%
b111 *
0-
02
b111 6
#383030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#383040000000
0!
0%
b0 *
0-
02
b0 6
#383050000000
1!
1%
1-
12
#383060000000
0!
0%
b1 *
0-
02
b1 6
#383070000000
1!
1%
1-
12
#383080000000
0!
0%
b10 *
0-
02
b10 6
#383090000000
1!
1%
1-
12
#383100000000
0!
0%
b11 *
0-
02
b11 6
#383110000000
1!
1%
1-
12
15
#383120000000
0!
0%
b100 *
0-
02
b100 6
#383130000000
1!
1%
1-
12
#383140000000
0!
0%
b101 *
0-
02
b101 6
#383150000000
1!
1%
1-
12
#383160000000
0!
0%
b110 *
0-
02
b110 6
#383170000000
1!
1%
1-
12
#383180000000
0!
0%
b111 *
0-
02
b111 6
#383190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#383200000000
0!
0%
b0 *
0-
02
b0 6
#383210000000
1!
1%
1-
12
#383220000000
0!
0%
b1 *
0-
02
b1 6
#383230000000
1!
1%
1-
12
#383240000000
0!
0%
b10 *
0-
02
b10 6
#383250000000
1!
1%
1-
12
#383260000000
0!
0%
b11 *
0-
02
b11 6
#383270000000
1!
1%
1-
12
15
#383280000000
0!
0%
b100 *
0-
02
b100 6
#383290000000
1!
1%
1-
12
#383300000000
0!
0%
b101 *
0-
02
b101 6
#383310000000
1!
1%
1-
12
#383320000000
0!
0%
b110 *
0-
02
b110 6
#383330000000
1!
1%
1-
12
#383340000000
0!
0%
b111 *
0-
02
b111 6
#383350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#383360000000
0!
0%
b0 *
0-
02
b0 6
#383370000000
1!
1%
1-
12
#383380000000
0!
0%
b1 *
0-
02
b1 6
#383390000000
1!
1%
1-
12
#383400000000
0!
0%
b10 *
0-
02
b10 6
#383410000000
1!
1%
1-
12
#383420000000
0!
0%
b11 *
0-
02
b11 6
#383430000000
1!
1%
1-
12
15
#383440000000
0!
0%
b100 *
0-
02
b100 6
#383450000000
1!
1%
1-
12
#383460000000
0!
0%
b101 *
0-
02
b101 6
#383470000000
1!
1%
1-
12
#383480000000
0!
0%
b110 *
0-
02
b110 6
#383490000000
1!
1%
1-
12
#383500000000
0!
0%
b111 *
0-
02
b111 6
#383510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#383520000000
0!
0%
b0 *
0-
02
b0 6
#383530000000
1!
1%
1-
12
#383540000000
0!
0%
b1 *
0-
02
b1 6
#383550000000
1!
1%
1-
12
#383560000000
0!
0%
b10 *
0-
02
b10 6
#383570000000
1!
1%
1-
12
#383580000000
0!
0%
b11 *
0-
02
b11 6
#383590000000
1!
1%
1-
12
15
#383600000000
0!
0%
b100 *
0-
02
b100 6
#383610000000
1!
1%
1-
12
#383620000000
0!
0%
b101 *
0-
02
b101 6
#383630000000
1!
1%
1-
12
#383640000000
0!
0%
b110 *
0-
02
b110 6
#383650000000
1!
1%
1-
12
#383660000000
0!
0%
b111 *
0-
02
b111 6
#383670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#383680000000
0!
0%
b0 *
0-
02
b0 6
#383690000000
1!
1%
1-
12
#383700000000
0!
0%
b1 *
0-
02
b1 6
#383710000000
1!
1%
1-
12
#383720000000
0!
0%
b10 *
0-
02
b10 6
#383730000000
1!
1%
1-
12
#383740000000
0!
0%
b11 *
0-
02
b11 6
#383750000000
1!
1%
1-
12
15
#383760000000
0!
0%
b100 *
0-
02
b100 6
#383770000000
1!
1%
1-
12
#383780000000
0!
0%
b101 *
0-
02
b101 6
#383790000000
1!
1%
1-
12
#383800000000
0!
0%
b110 *
0-
02
b110 6
#383810000000
1!
1%
1-
12
#383820000000
0!
0%
b111 *
0-
02
b111 6
#383830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#383840000000
0!
0%
b0 *
0-
02
b0 6
#383850000000
1!
1%
1-
12
#383860000000
0!
0%
b1 *
0-
02
b1 6
#383870000000
1!
1%
1-
12
#383880000000
0!
0%
b10 *
0-
02
b10 6
#383890000000
1!
1%
1-
12
#383900000000
0!
0%
b11 *
0-
02
b11 6
#383910000000
1!
1%
1-
12
15
#383920000000
0!
0%
b100 *
0-
02
b100 6
#383930000000
1!
1%
1-
12
#383940000000
0!
0%
b101 *
0-
02
b101 6
#383950000000
1!
1%
1-
12
#383960000000
0!
0%
b110 *
0-
02
b110 6
#383970000000
1!
1%
1-
12
#383980000000
0!
0%
b111 *
0-
02
b111 6
#383990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#384000000000
0!
0%
b0 *
0-
02
b0 6
#384010000000
1!
1%
1-
12
#384020000000
0!
0%
b1 *
0-
02
b1 6
#384030000000
1!
1%
1-
12
#384040000000
0!
0%
b10 *
0-
02
b10 6
#384050000000
1!
1%
1-
12
#384060000000
0!
0%
b11 *
0-
02
b11 6
#384070000000
1!
1%
1-
12
15
#384080000000
0!
0%
b100 *
0-
02
b100 6
#384090000000
1!
1%
1-
12
#384100000000
0!
0%
b101 *
0-
02
b101 6
#384110000000
1!
1%
1-
12
#384120000000
0!
0%
b110 *
0-
02
b110 6
#384130000000
1!
1%
1-
12
#384140000000
0!
0%
b111 *
0-
02
b111 6
#384150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#384160000000
0!
0%
b0 *
0-
02
b0 6
#384170000000
1!
1%
1-
12
#384180000000
0!
0%
b1 *
0-
02
b1 6
#384190000000
1!
1%
1-
12
#384200000000
0!
0%
b10 *
0-
02
b10 6
#384210000000
1!
1%
1-
12
#384220000000
0!
0%
b11 *
0-
02
b11 6
#384230000000
1!
1%
1-
12
15
#384240000000
0!
0%
b100 *
0-
02
b100 6
#384250000000
1!
1%
1-
12
#384260000000
0!
0%
b101 *
0-
02
b101 6
#384270000000
1!
1%
1-
12
#384280000000
0!
0%
b110 *
0-
02
b110 6
#384290000000
1!
1%
1-
12
#384300000000
0!
0%
b111 *
0-
02
b111 6
#384310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#384320000000
0!
0%
b0 *
0-
02
b0 6
#384330000000
1!
1%
1-
12
#384340000000
0!
0%
b1 *
0-
02
b1 6
#384350000000
1!
1%
1-
12
#384360000000
0!
0%
b10 *
0-
02
b10 6
#384370000000
1!
1%
1-
12
#384380000000
0!
0%
b11 *
0-
02
b11 6
#384390000000
1!
1%
1-
12
15
#384400000000
0!
0%
b100 *
0-
02
b100 6
#384410000000
1!
1%
1-
12
#384420000000
0!
0%
b101 *
0-
02
b101 6
#384430000000
1!
1%
1-
12
#384440000000
0!
0%
b110 *
0-
02
b110 6
#384450000000
1!
1%
1-
12
#384460000000
0!
0%
b111 *
0-
02
b111 6
#384470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#384480000000
0!
0%
b0 *
0-
02
b0 6
#384490000000
1!
1%
1-
12
#384500000000
0!
0%
b1 *
0-
02
b1 6
#384510000000
1!
1%
1-
12
#384520000000
0!
0%
b10 *
0-
02
b10 6
#384530000000
1!
1%
1-
12
#384540000000
0!
0%
b11 *
0-
02
b11 6
#384550000000
1!
1%
1-
12
15
#384560000000
0!
0%
b100 *
0-
02
b100 6
#384570000000
1!
1%
1-
12
#384580000000
0!
0%
b101 *
0-
02
b101 6
#384590000000
1!
1%
1-
12
#384600000000
0!
0%
b110 *
0-
02
b110 6
#384610000000
1!
1%
1-
12
#384620000000
0!
0%
b111 *
0-
02
b111 6
#384630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#384640000000
0!
0%
b0 *
0-
02
b0 6
#384650000000
1!
1%
1-
12
#384660000000
0!
0%
b1 *
0-
02
b1 6
#384670000000
1!
1%
1-
12
#384680000000
0!
0%
b10 *
0-
02
b10 6
#384690000000
1!
1%
1-
12
#384700000000
0!
0%
b11 *
0-
02
b11 6
#384710000000
1!
1%
1-
12
15
#384720000000
0!
0%
b100 *
0-
02
b100 6
#384730000000
1!
1%
1-
12
#384740000000
0!
0%
b101 *
0-
02
b101 6
#384750000000
1!
1%
1-
12
#384760000000
0!
0%
b110 *
0-
02
b110 6
#384770000000
1!
1%
1-
12
#384780000000
0!
0%
b111 *
0-
02
b111 6
#384790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#384800000000
0!
0%
b0 *
0-
02
b0 6
#384810000000
1!
1%
1-
12
#384820000000
0!
0%
b1 *
0-
02
b1 6
#384830000000
1!
1%
1-
12
#384840000000
0!
0%
b10 *
0-
02
b10 6
#384850000000
1!
1%
1-
12
#384860000000
0!
0%
b11 *
0-
02
b11 6
#384870000000
1!
1%
1-
12
15
#384880000000
0!
0%
b100 *
0-
02
b100 6
#384890000000
1!
1%
1-
12
#384900000000
0!
0%
b101 *
0-
02
b101 6
#384910000000
1!
1%
1-
12
#384920000000
0!
0%
b110 *
0-
02
b110 6
#384930000000
1!
1%
1-
12
#384940000000
0!
0%
b111 *
0-
02
b111 6
#384950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#384960000000
0!
0%
b0 *
0-
02
b0 6
#384970000000
1!
1%
1-
12
#384980000000
0!
0%
b1 *
0-
02
b1 6
#384990000000
1!
1%
1-
12
#385000000000
0!
0%
b10 *
0-
02
b10 6
#385010000000
1!
1%
1-
12
#385020000000
0!
0%
b11 *
0-
02
b11 6
#385030000000
1!
1%
1-
12
15
#385040000000
0!
0%
b100 *
0-
02
b100 6
#385050000000
1!
1%
1-
12
#385060000000
0!
0%
b101 *
0-
02
b101 6
#385070000000
1!
1%
1-
12
#385080000000
0!
0%
b110 *
0-
02
b110 6
#385090000000
1!
1%
1-
12
#385100000000
0!
0%
b111 *
0-
02
b111 6
#385110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#385120000000
0!
0%
b0 *
0-
02
b0 6
#385130000000
1!
1%
1-
12
#385140000000
0!
0%
b1 *
0-
02
b1 6
#385150000000
1!
1%
1-
12
#385160000000
0!
0%
b10 *
0-
02
b10 6
#385170000000
1!
1%
1-
12
#385180000000
0!
0%
b11 *
0-
02
b11 6
#385190000000
1!
1%
1-
12
15
#385200000000
0!
0%
b100 *
0-
02
b100 6
#385210000000
1!
1%
1-
12
#385220000000
0!
0%
b101 *
0-
02
b101 6
#385230000000
1!
1%
1-
12
#385240000000
0!
0%
b110 *
0-
02
b110 6
#385250000000
1!
1%
1-
12
#385260000000
0!
0%
b111 *
0-
02
b111 6
#385270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#385280000000
0!
0%
b0 *
0-
02
b0 6
#385290000000
1!
1%
1-
12
#385300000000
0!
0%
b1 *
0-
02
b1 6
#385310000000
1!
1%
1-
12
#385320000000
0!
0%
b10 *
0-
02
b10 6
#385330000000
1!
1%
1-
12
#385340000000
0!
0%
b11 *
0-
02
b11 6
#385350000000
1!
1%
1-
12
15
#385360000000
0!
0%
b100 *
0-
02
b100 6
#385370000000
1!
1%
1-
12
#385380000000
0!
0%
b101 *
0-
02
b101 6
#385390000000
1!
1%
1-
12
#385400000000
0!
0%
b110 *
0-
02
b110 6
#385410000000
1!
1%
1-
12
#385420000000
0!
0%
b111 *
0-
02
b111 6
#385430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#385440000000
0!
0%
b0 *
0-
02
b0 6
#385450000000
1!
1%
1-
12
#385460000000
0!
0%
b1 *
0-
02
b1 6
#385470000000
1!
1%
1-
12
#385480000000
0!
0%
b10 *
0-
02
b10 6
#385490000000
1!
1%
1-
12
#385500000000
0!
0%
b11 *
0-
02
b11 6
#385510000000
1!
1%
1-
12
15
#385520000000
0!
0%
b100 *
0-
02
b100 6
#385530000000
1!
1%
1-
12
#385540000000
0!
0%
b101 *
0-
02
b101 6
#385550000000
1!
1%
1-
12
#385560000000
0!
0%
b110 *
0-
02
b110 6
#385570000000
1!
1%
1-
12
#385580000000
0!
0%
b111 *
0-
02
b111 6
#385590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#385600000000
0!
0%
b0 *
0-
02
b0 6
#385610000000
1!
1%
1-
12
#385620000000
0!
0%
b1 *
0-
02
b1 6
#385630000000
1!
1%
1-
12
#385640000000
0!
0%
b10 *
0-
02
b10 6
#385650000000
1!
1%
1-
12
#385660000000
0!
0%
b11 *
0-
02
b11 6
#385670000000
1!
1%
1-
12
15
#385680000000
0!
0%
b100 *
0-
02
b100 6
#385690000000
1!
1%
1-
12
#385700000000
0!
0%
b101 *
0-
02
b101 6
#385710000000
1!
1%
1-
12
#385720000000
0!
0%
b110 *
0-
02
b110 6
#385730000000
1!
1%
1-
12
#385740000000
0!
0%
b111 *
0-
02
b111 6
#385750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#385760000000
0!
0%
b0 *
0-
02
b0 6
#385770000000
1!
1%
1-
12
#385780000000
0!
0%
b1 *
0-
02
b1 6
#385790000000
1!
1%
1-
12
#385800000000
0!
0%
b10 *
0-
02
b10 6
#385810000000
1!
1%
1-
12
#385820000000
0!
0%
b11 *
0-
02
b11 6
#385830000000
1!
1%
1-
12
15
#385840000000
0!
0%
b100 *
0-
02
b100 6
#385850000000
1!
1%
1-
12
#385860000000
0!
0%
b101 *
0-
02
b101 6
#385870000000
1!
1%
1-
12
#385880000000
0!
0%
b110 *
0-
02
b110 6
#385890000000
1!
1%
1-
12
#385900000000
0!
0%
b111 *
0-
02
b111 6
#385910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#385920000000
0!
0%
b0 *
0-
02
b0 6
#385930000000
1!
1%
1-
12
#385940000000
0!
0%
b1 *
0-
02
b1 6
#385950000000
1!
1%
1-
12
#385960000000
0!
0%
b10 *
0-
02
b10 6
#385970000000
1!
1%
1-
12
#385980000000
0!
0%
b11 *
0-
02
b11 6
#385990000000
1!
1%
1-
12
15
#386000000000
0!
0%
b100 *
0-
02
b100 6
#386010000000
1!
1%
1-
12
#386020000000
0!
0%
b101 *
0-
02
b101 6
#386030000000
1!
1%
1-
12
#386040000000
0!
0%
b110 *
0-
02
b110 6
#386050000000
1!
1%
1-
12
#386060000000
0!
0%
b111 *
0-
02
b111 6
#386070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#386080000000
0!
0%
b0 *
0-
02
b0 6
#386090000000
1!
1%
1-
12
#386100000000
0!
0%
b1 *
0-
02
b1 6
#386110000000
1!
1%
1-
12
#386120000000
0!
0%
b10 *
0-
02
b10 6
#386130000000
1!
1%
1-
12
#386140000000
0!
0%
b11 *
0-
02
b11 6
#386150000000
1!
1%
1-
12
15
#386160000000
0!
0%
b100 *
0-
02
b100 6
#386170000000
1!
1%
1-
12
#386180000000
0!
0%
b101 *
0-
02
b101 6
#386190000000
1!
1%
1-
12
#386200000000
0!
0%
b110 *
0-
02
b110 6
#386210000000
1!
1%
1-
12
#386220000000
0!
0%
b111 *
0-
02
b111 6
#386230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#386240000000
0!
0%
b0 *
0-
02
b0 6
#386250000000
1!
1%
1-
12
#386260000000
0!
0%
b1 *
0-
02
b1 6
#386270000000
1!
1%
1-
12
#386280000000
0!
0%
b10 *
0-
02
b10 6
#386290000000
1!
1%
1-
12
#386300000000
0!
0%
b11 *
0-
02
b11 6
#386310000000
1!
1%
1-
12
15
#386320000000
0!
0%
b100 *
0-
02
b100 6
#386330000000
1!
1%
1-
12
#386340000000
0!
0%
b101 *
0-
02
b101 6
#386350000000
1!
1%
1-
12
#386360000000
0!
0%
b110 *
0-
02
b110 6
#386370000000
1!
1%
1-
12
#386380000000
0!
0%
b111 *
0-
02
b111 6
#386390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#386400000000
0!
0%
b0 *
0-
02
b0 6
#386410000000
1!
1%
1-
12
#386420000000
0!
0%
b1 *
0-
02
b1 6
#386430000000
1!
1%
1-
12
#386440000000
0!
0%
b10 *
0-
02
b10 6
#386450000000
1!
1%
1-
12
#386460000000
0!
0%
b11 *
0-
02
b11 6
#386470000000
1!
1%
1-
12
15
#386480000000
0!
0%
b100 *
0-
02
b100 6
#386490000000
1!
1%
1-
12
#386500000000
0!
0%
b101 *
0-
02
b101 6
#386510000000
1!
1%
1-
12
#386520000000
0!
0%
b110 *
0-
02
b110 6
#386530000000
1!
1%
1-
12
#386540000000
0!
0%
b111 *
0-
02
b111 6
#386550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#386560000000
0!
0%
b0 *
0-
02
b0 6
#386570000000
1!
1%
1-
12
#386580000000
0!
0%
b1 *
0-
02
b1 6
#386590000000
1!
1%
1-
12
#386600000000
0!
0%
b10 *
0-
02
b10 6
#386610000000
1!
1%
1-
12
#386620000000
0!
0%
b11 *
0-
02
b11 6
#386630000000
1!
1%
1-
12
15
#386640000000
0!
0%
b100 *
0-
02
b100 6
#386650000000
1!
1%
1-
12
#386660000000
0!
0%
b101 *
0-
02
b101 6
#386670000000
1!
1%
1-
12
#386680000000
0!
0%
b110 *
0-
02
b110 6
#386690000000
1!
1%
1-
12
#386700000000
0!
0%
b111 *
0-
02
b111 6
#386710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#386720000000
0!
0%
b0 *
0-
02
b0 6
#386730000000
1!
1%
1-
12
#386740000000
0!
0%
b1 *
0-
02
b1 6
#386750000000
1!
1%
1-
12
#386760000000
0!
0%
b10 *
0-
02
b10 6
#386770000000
1!
1%
1-
12
#386780000000
0!
0%
b11 *
0-
02
b11 6
#386790000000
1!
1%
1-
12
15
#386800000000
0!
0%
b100 *
0-
02
b100 6
#386810000000
1!
1%
1-
12
#386820000000
0!
0%
b101 *
0-
02
b101 6
#386830000000
1!
1%
1-
12
#386840000000
0!
0%
b110 *
0-
02
b110 6
#386850000000
1!
1%
1-
12
#386860000000
0!
0%
b111 *
0-
02
b111 6
#386870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#386880000000
0!
0%
b0 *
0-
02
b0 6
#386890000000
1!
1%
1-
12
#386900000000
0!
0%
b1 *
0-
02
b1 6
#386910000000
1!
1%
1-
12
#386920000000
0!
0%
b10 *
0-
02
b10 6
#386930000000
1!
1%
1-
12
#386940000000
0!
0%
b11 *
0-
02
b11 6
#386950000000
1!
1%
1-
12
15
#386960000000
0!
0%
b100 *
0-
02
b100 6
#386970000000
1!
1%
1-
12
#386980000000
0!
0%
b101 *
0-
02
b101 6
#386990000000
1!
1%
1-
12
#387000000000
0!
0%
b110 *
0-
02
b110 6
#387010000000
1!
1%
1-
12
#387020000000
0!
0%
b111 *
0-
02
b111 6
#387030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#387040000000
0!
0%
b0 *
0-
02
b0 6
#387050000000
1!
1%
1-
12
#387060000000
0!
0%
b1 *
0-
02
b1 6
#387070000000
1!
1%
1-
12
#387080000000
0!
0%
b10 *
0-
02
b10 6
#387090000000
1!
1%
1-
12
#387100000000
0!
0%
b11 *
0-
02
b11 6
#387110000000
1!
1%
1-
12
15
#387120000000
0!
0%
b100 *
0-
02
b100 6
#387130000000
1!
1%
1-
12
#387140000000
0!
0%
b101 *
0-
02
b101 6
#387150000000
1!
1%
1-
12
#387160000000
0!
0%
b110 *
0-
02
b110 6
#387170000000
1!
1%
1-
12
#387180000000
0!
0%
b111 *
0-
02
b111 6
#387190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#387200000000
0!
0%
b0 *
0-
02
b0 6
#387210000000
1!
1%
1-
12
#387220000000
0!
0%
b1 *
0-
02
b1 6
#387230000000
1!
1%
1-
12
#387240000000
0!
0%
b10 *
0-
02
b10 6
#387250000000
1!
1%
1-
12
#387260000000
0!
0%
b11 *
0-
02
b11 6
#387270000000
1!
1%
1-
12
15
#387280000000
0!
0%
b100 *
0-
02
b100 6
#387290000000
1!
1%
1-
12
#387300000000
0!
0%
b101 *
0-
02
b101 6
#387310000000
1!
1%
1-
12
#387320000000
0!
0%
b110 *
0-
02
b110 6
#387330000000
1!
1%
1-
12
#387340000000
0!
0%
b111 *
0-
02
b111 6
#387350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#387360000000
0!
0%
b0 *
0-
02
b0 6
#387370000000
1!
1%
1-
12
#387380000000
0!
0%
b1 *
0-
02
b1 6
#387390000000
1!
1%
1-
12
#387400000000
0!
0%
b10 *
0-
02
b10 6
#387410000000
1!
1%
1-
12
#387420000000
0!
0%
b11 *
0-
02
b11 6
#387430000000
1!
1%
1-
12
15
#387440000000
0!
0%
b100 *
0-
02
b100 6
#387450000000
1!
1%
1-
12
#387460000000
0!
0%
b101 *
0-
02
b101 6
#387470000000
1!
1%
1-
12
#387480000000
0!
0%
b110 *
0-
02
b110 6
#387490000000
1!
1%
1-
12
#387500000000
0!
0%
b111 *
0-
02
b111 6
#387510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#387520000000
0!
0%
b0 *
0-
02
b0 6
#387530000000
1!
1%
1-
12
#387540000000
0!
0%
b1 *
0-
02
b1 6
#387550000000
1!
1%
1-
12
#387560000000
0!
0%
b10 *
0-
02
b10 6
#387570000000
1!
1%
1-
12
#387580000000
0!
0%
b11 *
0-
02
b11 6
#387590000000
1!
1%
1-
12
15
#387600000000
0!
0%
b100 *
0-
02
b100 6
#387610000000
1!
1%
1-
12
#387620000000
0!
0%
b101 *
0-
02
b101 6
#387630000000
1!
1%
1-
12
#387640000000
0!
0%
b110 *
0-
02
b110 6
#387650000000
1!
1%
1-
12
#387660000000
0!
0%
b111 *
0-
02
b111 6
#387670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#387680000000
0!
0%
b0 *
0-
02
b0 6
#387690000000
1!
1%
1-
12
#387700000000
0!
0%
b1 *
0-
02
b1 6
#387710000000
1!
1%
1-
12
#387720000000
0!
0%
b10 *
0-
02
b10 6
#387730000000
1!
1%
1-
12
#387740000000
0!
0%
b11 *
0-
02
b11 6
#387750000000
1!
1%
1-
12
15
#387760000000
0!
0%
b100 *
0-
02
b100 6
#387770000000
1!
1%
1-
12
#387780000000
0!
0%
b101 *
0-
02
b101 6
#387790000000
1!
1%
1-
12
#387800000000
0!
0%
b110 *
0-
02
b110 6
#387810000000
1!
1%
1-
12
#387820000000
0!
0%
b111 *
0-
02
b111 6
#387830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#387840000000
0!
0%
b0 *
0-
02
b0 6
#387850000000
1!
1%
1-
12
#387860000000
0!
0%
b1 *
0-
02
b1 6
#387870000000
1!
1%
1-
12
#387880000000
0!
0%
b10 *
0-
02
b10 6
#387890000000
1!
1%
1-
12
#387900000000
0!
0%
b11 *
0-
02
b11 6
#387910000000
1!
1%
1-
12
15
#387920000000
0!
0%
b100 *
0-
02
b100 6
#387930000000
1!
1%
1-
12
#387940000000
0!
0%
b101 *
0-
02
b101 6
#387950000000
1!
1%
1-
12
#387960000000
0!
0%
b110 *
0-
02
b110 6
#387970000000
1!
1%
1-
12
#387980000000
0!
0%
b111 *
0-
02
b111 6
#387990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#388000000000
0!
0%
b0 *
0-
02
b0 6
#388010000000
1!
1%
1-
12
#388020000000
0!
0%
b1 *
0-
02
b1 6
#388030000000
1!
1%
1-
12
#388040000000
0!
0%
b10 *
0-
02
b10 6
#388050000000
1!
1%
1-
12
#388060000000
0!
0%
b11 *
0-
02
b11 6
#388070000000
1!
1%
1-
12
15
#388080000000
0!
0%
b100 *
0-
02
b100 6
#388090000000
1!
1%
1-
12
#388100000000
0!
0%
b101 *
0-
02
b101 6
#388110000000
1!
1%
1-
12
#388120000000
0!
0%
b110 *
0-
02
b110 6
#388130000000
1!
1%
1-
12
#388140000000
0!
0%
b111 *
0-
02
b111 6
#388150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#388160000000
0!
0%
b0 *
0-
02
b0 6
#388170000000
1!
1%
1-
12
#388180000000
0!
0%
b1 *
0-
02
b1 6
#388190000000
1!
1%
1-
12
#388200000000
0!
0%
b10 *
0-
02
b10 6
#388210000000
1!
1%
1-
12
#388220000000
0!
0%
b11 *
0-
02
b11 6
#388230000000
1!
1%
1-
12
15
#388240000000
0!
0%
b100 *
0-
02
b100 6
#388250000000
1!
1%
1-
12
#388260000000
0!
0%
b101 *
0-
02
b101 6
#388270000000
1!
1%
1-
12
#388280000000
0!
0%
b110 *
0-
02
b110 6
#388290000000
1!
1%
1-
12
#388300000000
0!
0%
b111 *
0-
02
b111 6
#388310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#388320000000
0!
0%
b0 *
0-
02
b0 6
#388330000000
1!
1%
1-
12
#388340000000
0!
0%
b1 *
0-
02
b1 6
#388350000000
1!
1%
1-
12
#388360000000
0!
0%
b10 *
0-
02
b10 6
#388370000000
1!
1%
1-
12
#388380000000
0!
0%
b11 *
0-
02
b11 6
#388390000000
1!
1%
1-
12
15
#388400000000
0!
0%
b100 *
0-
02
b100 6
#388410000000
1!
1%
1-
12
#388420000000
0!
0%
b101 *
0-
02
b101 6
#388430000000
1!
1%
1-
12
#388440000000
0!
0%
b110 *
0-
02
b110 6
#388450000000
1!
1%
1-
12
#388460000000
0!
0%
b111 *
0-
02
b111 6
#388470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#388480000000
0!
0%
b0 *
0-
02
b0 6
#388490000000
1!
1%
1-
12
#388500000000
0!
0%
b1 *
0-
02
b1 6
#388510000000
1!
1%
1-
12
#388520000000
0!
0%
b10 *
0-
02
b10 6
#388530000000
1!
1%
1-
12
#388540000000
0!
0%
b11 *
0-
02
b11 6
#388550000000
1!
1%
1-
12
15
#388560000000
0!
0%
b100 *
0-
02
b100 6
#388570000000
1!
1%
1-
12
#388580000000
0!
0%
b101 *
0-
02
b101 6
#388590000000
1!
1%
1-
12
#388600000000
0!
0%
b110 *
0-
02
b110 6
#388610000000
1!
1%
1-
12
#388620000000
0!
0%
b111 *
0-
02
b111 6
#388630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#388640000000
0!
0%
b0 *
0-
02
b0 6
#388650000000
1!
1%
1-
12
#388660000000
0!
0%
b1 *
0-
02
b1 6
#388670000000
1!
1%
1-
12
#388680000000
0!
0%
b10 *
0-
02
b10 6
#388690000000
1!
1%
1-
12
#388700000000
0!
0%
b11 *
0-
02
b11 6
#388710000000
1!
1%
1-
12
15
#388720000000
0!
0%
b100 *
0-
02
b100 6
#388730000000
1!
1%
1-
12
#388740000000
0!
0%
b101 *
0-
02
b101 6
#388750000000
1!
1%
1-
12
#388760000000
0!
0%
b110 *
0-
02
b110 6
#388770000000
1!
1%
1-
12
#388780000000
0!
0%
b111 *
0-
02
b111 6
#388790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#388800000000
0!
0%
b0 *
0-
02
b0 6
#388810000000
1!
1%
1-
12
#388820000000
0!
0%
b1 *
0-
02
b1 6
#388830000000
1!
1%
1-
12
#388840000000
0!
0%
b10 *
0-
02
b10 6
#388850000000
1!
1%
1-
12
#388860000000
0!
0%
b11 *
0-
02
b11 6
#388870000000
1!
1%
1-
12
15
#388880000000
0!
0%
b100 *
0-
02
b100 6
#388890000000
1!
1%
1-
12
#388900000000
0!
0%
b101 *
0-
02
b101 6
#388910000000
1!
1%
1-
12
#388920000000
0!
0%
b110 *
0-
02
b110 6
#388930000000
1!
1%
1-
12
#388940000000
0!
0%
b111 *
0-
02
b111 6
#388950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#388960000000
0!
0%
b0 *
0-
02
b0 6
#388970000000
1!
1%
1-
12
#388980000000
0!
0%
b1 *
0-
02
b1 6
#388990000000
1!
1%
1-
12
#389000000000
0!
0%
b10 *
0-
02
b10 6
#389010000000
1!
1%
1-
12
#389020000000
0!
0%
b11 *
0-
02
b11 6
#389030000000
1!
1%
1-
12
15
#389040000000
0!
0%
b100 *
0-
02
b100 6
#389050000000
1!
1%
1-
12
#389060000000
0!
0%
b101 *
0-
02
b101 6
#389070000000
1!
1%
1-
12
#389080000000
0!
0%
b110 *
0-
02
b110 6
#389090000000
1!
1%
1-
12
#389100000000
0!
0%
b111 *
0-
02
b111 6
#389110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#389120000000
0!
0%
b0 *
0-
02
b0 6
#389130000000
1!
1%
1-
12
#389140000000
0!
0%
b1 *
0-
02
b1 6
#389150000000
1!
1%
1-
12
#389160000000
0!
0%
b10 *
0-
02
b10 6
#389170000000
1!
1%
1-
12
#389180000000
0!
0%
b11 *
0-
02
b11 6
#389190000000
1!
1%
1-
12
15
#389200000000
0!
0%
b100 *
0-
02
b100 6
#389210000000
1!
1%
1-
12
#389220000000
0!
0%
b101 *
0-
02
b101 6
#389230000000
1!
1%
1-
12
#389240000000
0!
0%
b110 *
0-
02
b110 6
#389250000000
1!
1%
1-
12
#389260000000
0!
0%
b111 *
0-
02
b111 6
#389270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#389280000000
0!
0%
b0 *
0-
02
b0 6
#389290000000
1!
1%
1-
12
#389300000000
0!
0%
b1 *
0-
02
b1 6
#389310000000
1!
1%
1-
12
#389320000000
0!
0%
b10 *
0-
02
b10 6
#389330000000
1!
1%
1-
12
#389340000000
0!
0%
b11 *
0-
02
b11 6
#389350000000
1!
1%
1-
12
15
#389360000000
0!
0%
b100 *
0-
02
b100 6
#389370000000
1!
1%
1-
12
#389380000000
0!
0%
b101 *
0-
02
b101 6
#389390000000
1!
1%
1-
12
#389400000000
0!
0%
b110 *
0-
02
b110 6
#389410000000
1!
1%
1-
12
#389420000000
0!
0%
b111 *
0-
02
b111 6
#389430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#389440000000
0!
0%
b0 *
0-
02
b0 6
#389450000000
1!
1%
1-
12
#389460000000
0!
0%
b1 *
0-
02
b1 6
#389470000000
1!
1%
1-
12
#389480000000
0!
0%
b10 *
0-
02
b10 6
#389490000000
1!
1%
1-
12
#389500000000
0!
0%
b11 *
0-
02
b11 6
#389510000000
1!
1%
1-
12
15
#389520000000
0!
0%
b100 *
0-
02
b100 6
#389530000000
1!
1%
1-
12
#389540000000
0!
0%
b101 *
0-
02
b101 6
#389550000000
1!
1%
1-
12
#389560000000
0!
0%
b110 *
0-
02
b110 6
#389570000000
1!
1%
1-
12
#389580000000
0!
0%
b111 *
0-
02
b111 6
#389590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#389600000000
0!
0%
b0 *
0-
02
b0 6
#389610000000
1!
1%
1-
12
#389620000000
0!
0%
b1 *
0-
02
b1 6
#389630000000
1!
1%
1-
12
#389640000000
0!
0%
b10 *
0-
02
b10 6
#389650000000
1!
1%
1-
12
#389660000000
0!
0%
b11 *
0-
02
b11 6
#389670000000
1!
1%
1-
12
15
#389680000000
0!
0%
b100 *
0-
02
b100 6
#389690000000
1!
1%
1-
12
#389700000000
0!
0%
b101 *
0-
02
b101 6
#389710000000
1!
1%
1-
12
#389720000000
0!
0%
b110 *
0-
02
b110 6
#389730000000
1!
1%
1-
12
#389740000000
0!
0%
b111 *
0-
02
b111 6
#389750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#389760000000
0!
0%
b0 *
0-
02
b0 6
#389770000000
1!
1%
1-
12
#389780000000
0!
0%
b1 *
0-
02
b1 6
#389790000000
1!
1%
1-
12
#389800000000
0!
0%
b10 *
0-
02
b10 6
#389810000000
1!
1%
1-
12
#389820000000
0!
0%
b11 *
0-
02
b11 6
#389830000000
1!
1%
1-
12
15
#389840000000
0!
0%
b100 *
0-
02
b100 6
#389850000000
1!
1%
1-
12
#389860000000
0!
0%
b101 *
0-
02
b101 6
#389870000000
1!
1%
1-
12
#389880000000
0!
0%
b110 *
0-
02
b110 6
#389890000000
1!
1%
1-
12
#389900000000
0!
0%
b111 *
0-
02
b111 6
#389910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#389920000000
0!
0%
b0 *
0-
02
b0 6
#389930000000
1!
1%
1-
12
#389940000000
0!
0%
b1 *
0-
02
b1 6
#389950000000
1!
1%
1-
12
#389960000000
0!
0%
b10 *
0-
02
b10 6
#389970000000
1!
1%
1-
12
#389980000000
0!
0%
b11 *
0-
02
b11 6
#389990000000
1!
1%
1-
12
15
#390000000000
0!
0%
b100 *
0-
02
b100 6
#390010000000
1!
1%
1-
12
#390020000000
0!
0%
b101 *
0-
02
b101 6
#390030000000
1!
1%
1-
12
#390040000000
0!
0%
b110 *
0-
02
b110 6
#390050000000
1!
1%
1-
12
#390060000000
0!
0%
b111 *
0-
02
b111 6
#390070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#390080000000
0!
0%
b0 *
0-
02
b0 6
#390090000000
1!
1%
1-
12
#390100000000
0!
0%
b1 *
0-
02
b1 6
#390110000000
1!
1%
1-
12
#390120000000
0!
0%
b10 *
0-
02
b10 6
#390130000000
1!
1%
1-
12
#390140000000
0!
0%
b11 *
0-
02
b11 6
#390150000000
1!
1%
1-
12
15
#390160000000
0!
0%
b100 *
0-
02
b100 6
#390170000000
1!
1%
1-
12
#390180000000
0!
0%
b101 *
0-
02
b101 6
#390190000000
1!
1%
1-
12
#390200000000
0!
0%
b110 *
0-
02
b110 6
#390210000000
1!
1%
1-
12
#390220000000
0!
0%
b111 *
0-
02
b111 6
#390230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#390240000000
0!
0%
b0 *
0-
02
b0 6
#390250000000
1!
1%
1-
12
#390260000000
0!
0%
b1 *
0-
02
b1 6
#390270000000
1!
1%
1-
12
#390280000000
0!
0%
b10 *
0-
02
b10 6
#390290000000
1!
1%
1-
12
#390300000000
0!
0%
b11 *
0-
02
b11 6
#390310000000
1!
1%
1-
12
15
#390320000000
0!
0%
b100 *
0-
02
b100 6
#390330000000
1!
1%
1-
12
#390340000000
0!
0%
b101 *
0-
02
b101 6
#390350000000
1!
1%
1-
12
#390360000000
0!
0%
b110 *
0-
02
b110 6
#390370000000
1!
1%
1-
12
#390380000000
0!
0%
b111 *
0-
02
b111 6
#390390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#390400000000
0!
0%
b0 *
0-
02
b0 6
#390410000000
1!
1%
1-
12
#390420000000
0!
0%
b1 *
0-
02
b1 6
#390430000000
1!
1%
1-
12
#390440000000
0!
0%
b10 *
0-
02
b10 6
#390450000000
1!
1%
1-
12
#390460000000
0!
0%
b11 *
0-
02
b11 6
#390470000000
1!
1%
1-
12
15
#390480000000
0!
0%
b100 *
0-
02
b100 6
#390490000000
1!
1%
1-
12
#390500000000
0!
0%
b101 *
0-
02
b101 6
#390510000000
1!
1%
1-
12
#390520000000
0!
0%
b110 *
0-
02
b110 6
#390530000000
1!
1%
1-
12
#390540000000
0!
0%
b111 *
0-
02
b111 6
#390550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#390560000000
0!
0%
b0 *
0-
02
b0 6
#390570000000
1!
1%
1-
12
#390580000000
0!
0%
b1 *
0-
02
b1 6
#390590000000
1!
1%
1-
12
#390600000000
0!
0%
b10 *
0-
02
b10 6
#390610000000
1!
1%
1-
12
#390620000000
0!
0%
b11 *
0-
02
b11 6
#390630000000
1!
1%
1-
12
15
#390640000000
0!
0%
b100 *
0-
02
b100 6
#390650000000
1!
1%
1-
12
#390660000000
0!
0%
b101 *
0-
02
b101 6
#390670000000
1!
1%
1-
12
#390680000000
0!
0%
b110 *
0-
02
b110 6
#390690000000
1!
1%
1-
12
#390700000000
0!
0%
b111 *
0-
02
b111 6
#390710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#390720000000
0!
0%
b0 *
0-
02
b0 6
#390730000000
1!
1%
1-
12
#390740000000
0!
0%
b1 *
0-
02
b1 6
#390750000000
1!
1%
1-
12
#390760000000
0!
0%
b10 *
0-
02
b10 6
#390770000000
1!
1%
1-
12
#390780000000
0!
0%
b11 *
0-
02
b11 6
#390790000000
1!
1%
1-
12
15
#390800000000
0!
0%
b100 *
0-
02
b100 6
#390810000000
1!
1%
1-
12
#390820000000
0!
0%
b101 *
0-
02
b101 6
#390830000000
1!
1%
1-
12
#390840000000
0!
0%
b110 *
0-
02
b110 6
#390850000000
1!
1%
1-
12
#390860000000
0!
0%
b111 *
0-
02
b111 6
#390870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#390880000000
0!
0%
b0 *
0-
02
b0 6
#390890000000
1!
1%
1-
12
#390900000000
0!
0%
b1 *
0-
02
b1 6
#390910000000
1!
1%
1-
12
#390920000000
0!
0%
b10 *
0-
02
b10 6
#390930000000
1!
1%
1-
12
#390940000000
0!
0%
b11 *
0-
02
b11 6
#390950000000
1!
1%
1-
12
15
#390960000000
0!
0%
b100 *
0-
02
b100 6
#390970000000
1!
1%
1-
12
#390980000000
0!
0%
b101 *
0-
02
b101 6
#390990000000
1!
1%
1-
12
#391000000000
0!
0%
b110 *
0-
02
b110 6
#391010000000
1!
1%
1-
12
#391020000000
0!
0%
b111 *
0-
02
b111 6
#391030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#391040000000
0!
0%
b0 *
0-
02
b0 6
#391050000000
1!
1%
1-
12
#391060000000
0!
0%
b1 *
0-
02
b1 6
#391070000000
1!
1%
1-
12
#391080000000
0!
0%
b10 *
0-
02
b10 6
#391090000000
1!
1%
1-
12
#391100000000
0!
0%
b11 *
0-
02
b11 6
#391110000000
1!
1%
1-
12
15
#391120000000
0!
0%
b100 *
0-
02
b100 6
#391130000000
1!
1%
1-
12
#391140000000
0!
0%
b101 *
0-
02
b101 6
#391150000000
1!
1%
1-
12
#391160000000
0!
0%
b110 *
0-
02
b110 6
#391170000000
1!
1%
1-
12
#391180000000
0!
0%
b111 *
0-
02
b111 6
#391190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#391200000000
0!
0%
b0 *
0-
02
b0 6
#391210000000
1!
1%
1-
12
#391220000000
0!
0%
b1 *
0-
02
b1 6
#391230000000
1!
1%
1-
12
#391240000000
0!
0%
b10 *
0-
02
b10 6
#391250000000
1!
1%
1-
12
#391260000000
0!
0%
b11 *
0-
02
b11 6
#391270000000
1!
1%
1-
12
15
#391280000000
0!
0%
b100 *
0-
02
b100 6
#391290000000
1!
1%
1-
12
#391300000000
0!
0%
b101 *
0-
02
b101 6
#391310000000
1!
1%
1-
12
#391320000000
0!
0%
b110 *
0-
02
b110 6
#391330000000
1!
1%
1-
12
#391340000000
0!
0%
b111 *
0-
02
b111 6
#391350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#391360000000
0!
0%
b0 *
0-
02
b0 6
#391370000000
1!
1%
1-
12
#391380000000
0!
0%
b1 *
0-
02
b1 6
#391390000000
1!
1%
1-
12
#391400000000
0!
0%
b10 *
0-
02
b10 6
#391410000000
1!
1%
1-
12
#391420000000
0!
0%
b11 *
0-
02
b11 6
#391430000000
1!
1%
1-
12
15
#391440000000
0!
0%
b100 *
0-
02
b100 6
#391450000000
1!
1%
1-
12
#391460000000
0!
0%
b101 *
0-
02
b101 6
#391470000000
1!
1%
1-
12
#391480000000
0!
0%
b110 *
0-
02
b110 6
#391490000000
1!
1%
1-
12
#391500000000
0!
0%
b111 *
0-
02
b111 6
#391510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#391520000000
0!
0%
b0 *
0-
02
b0 6
#391530000000
1!
1%
1-
12
#391540000000
0!
0%
b1 *
0-
02
b1 6
#391550000000
1!
1%
1-
12
#391560000000
0!
0%
b10 *
0-
02
b10 6
#391570000000
1!
1%
1-
12
#391580000000
0!
0%
b11 *
0-
02
b11 6
#391590000000
1!
1%
1-
12
15
#391600000000
0!
0%
b100 *
0-
02
b100 6
#391610000000
1!
1%
1-
12
#391620000000
0!
0%
b101 *
0-
02
b101 6
#391630000000
1!
1%
1-
12
#391640000000
0!
0%
b110 *
0-
02
b110 6
#391650000000
1!
1%
1-
12
#391660000000
0!
0%
b111 *
0-
02
b111 6
#391670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#391680000000
0!
0%
b0 *
0-
02
b0 6
#391690000000
1!
1%
1-
12
#391700000000
0!
0%
b1 *
0-
02
b1 6
#391710000000
1!
1%
1-
12
#391720000000
0!
0%
b10 *
0-
02
b10 6
#391730000000
1!
1%
1-
12
#391740000000
0!
0%
b11 *
0-
02
b11 6
#391750000000
1!
1%
1-
12
15
#391760000000
0!
0%
b100 *
0-
02
b100 6
#391770000000
1!
1%
1-
12
#391780000000
0!
0%
b101 *
0-
02
b101 6
#391790000000
1!
1%
1-
12
#391800000000
0!
0%
b110 *
0-
02
b110 6
#391810000000
1!
1%
1-
12
#391820000000
0!
0%
b111 *
0-
02
b111 6
#391830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#391840000000
0!
0%
b0 *
0-
02
b0 6
#391850000000
1!
1%
1-
12
#391860000000
0!
0%
b1 *
0-
02
b1 6
#391870000000
1!
1%
1-
12
#391880000000
0!
0%
b10 *
0-
02
b10 6
#391890000000
1!
1%
1-
12
#391900000000
0!
0%
b11 *
0-
02
b11 6
#391910000000
1!
1%
1-
12
15
#391920000000
0!
0%
b100 *
0-
02
b100 6
#391930000000
1!
1%
1-
12
#391940000000
0!
0%
b101 *
0-
02
b101 6
#391950000000
1!
1%
1-
12
#391960000000
0!
0%
b110 *
0-
02
b110 6
#391970000000
1!
1%
1-
12
#391980000000
0!
0%
b111 *
0-
02
b111 6
#391990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#392000000000
0!
0%
b0 *
0-
02
b0 6
#392010000000
1!
1%
1-
12
#392020000000
0!
0%
b1 *
0-
02
b1 6
#392030000000
1!
1%
1-
12
#392040000000
0!
0%
b10 *
0-
02
b10 6
#392050000000
1!
1%
1-
12
#392060000000
0!
0%
b11 *
0-
02
b11 6
#392070000000
1!
1%
1-
12
15
#392080000000
0!
0%
b100 *
0-
02
b100 6
#392090000000
1!
1%
1-
12
#392100000000
0!
0%
b101 *
0-
02
b101 6
#392110000000
1!
1%
1-
12
#392120000000
0!
0%
b110 *
0-
02
b110 6
#392130000000
1!
1%
1-
12
#392140000000
0!
0%
b111 *
0-
02
b111 6
#392150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#392160000000
0!
0%
b0 *
0-
02
b0 6
#392170000000
1!
1%
1-
12
#392180000000
0!
0%
b1 *
0-
02
b1 6
#392190000000
1!
1%
1-
12
#392200000000
0!
0%
b10 *
0-
02
b10 6
#392210000000
1!
1%
1-
12
#392220000000
0!
0%
b11 *
0-
02
b11 6
#392230000000
1!
1%
1-
12
15
#392240000000
0!
0%
b100 *
0-
02
b100 6
#392250000000
1!
1%
1-
12
#392260000000
0!
0%
b101 *
0-
02
b101 6
#392270000000
1!
1%
1-
12
#392280000000
0!
0%
b110 *
0-
02
b110 6
#392290000000
1!
1%
1-
12
#392300000000
0!
0%
b111 *
0-
02
b111 6
#392310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#392320000000
0!
0%
b0 *
0-
02
b0 6
#392330000000
1!
1%
1-
12
#392340000000
0!
0%
b1 *
0-
02
b1 6
#392350000000
1!
1%
1-
12
#392360000000
0!
0%
b10 *
0-
02
b10 6
#392370000000
1!
1%
1-
12
#392380000000
0!
0%
b11 *
0-
02
b11 6
#392390000000
1!
1%
1-
12
15
#392400000000
0!
0%
b100 *
0-
02
b100 6
#392410000000
1!
1%
1-
12
#392420000000
0!
0%
b101 *
0-
02
b101 6
#392430000000
1!
1%
1-
12
#392440000000
0!
0%
b110 *
0-
02
b110 6
#392450000000
1!
1%
1-
12
#392460000000
0!
0%
b111 *
0-
02
b111 6
#392470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#392480000000
0!
0%
b0 *
0-
02
b0 6
#392490000000
1!
1%
1-
12
#392500000000
0!
0%
b1 *
0-
02
b1 6
#392510000000
1!
1%
1-
12
#392520000000
0!
0%
b10 *
0-
02
b10 6
#392530000000
1!
1%
1-
12
#392540000000
0!
0%
b11 *
0-
02
b11 6
#392550000000
1!
1%
1-
12
15
#392560000000
0!
0%
b100 *
0-
02
b100 6
#392570000000
1!
1%
1-
12
#392580000000
0!
0%
b101 *
0-
02
b101 6
#392590000000
1!
1%
1-
12
#392600000000
0!
0%
b110 *
0-
02
b110 6
#392610000000
1!
1%
1-
12
#392620000000
0!
0%
b111 *
0-
02
b111 6
#392630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#392640000000
0!
0%
b0 *
0-
02
b0 6
#392650000000
1!
1%
1-
12
#392660000000
0!
0%
b1 *
0-
02
b1 6
#392670000000
1!
1%
1-
12
#392680000000
0!
0%
b10 *
0-
02
b10 6
#392690000000
1!
1%
1-
12
#392700000000
0!
0%
b11 *
0-
02
b11 6
#392710000000
1!
1%
1-
12
15
#392720000000
0!
0%
b100 *
0-
02
b100 6
#392730000000
1!
1%
1-
12
#392740000000
0!
0%
b101 *
0-
02
b101 6
#392750000000
1!
1%
1-
12
#392760000000
0!
0%
b110 *
0-
02
b110 6
#392770000000
1!
1%
1-
12
#392780000000
0!
0%
b111 *
0-
02
b111 6
#392790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#392800000000
0!
0%
b0 *
0-
02
b0 6
#392810000000
1!
1%
1-
12
#392820000000
0!
0%
b1 *
0-
02
b1 6
#392830000000
1!
1%
1-
12
#392840000000
0!
0%
b10 *
0-
02
b10 6
#392850000000
1!
1%
1-
12
#392860000000
0!
0%
b11 *
0-
02
b11 6
#392870000000
1!
1%
1-
12
15
#392880000000
0!
0%
b100 *
0-
02
b100 6
#392890000000
1!
1%
1-
12
#392900000000
0!
0%
b101 *
0-
02
b101 6
#392910000000
1!
1%
1-
12
#392920000000
0!
0%
b110 *
0-
02
b110 6
#392930000000
1!
1%
1-
12
#392940000000
0!
0%
b111 *
0-
02
b111 6
#392950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#392960000000
0!
0%
b0 *
0-
02
b0 6
#392970000000
1!
1%
1-
12
#392980000000
0!
0%
b1 *
0-
02
b1 6
#392990000000
1!
1%
1-
12
#393000000000
0!
0%
b10 *
0-
02
b10 6
#393010000000
1!
1%
1-
12
#393020000000
0!
0%
b11 *
0-
02
b11 6
#393030000000
1!
1%
1-
12
15
#393040000000
0!
0%
b100 *
0-
02
b100 6
#393050000000
1!
1%
1-
12
#393060000000
0!
0%
b101 *
0-
02
b101 6
#393070000000
1!
1%
1-
12
#393080000000
0!
0%
b110 *
0-
02
b110 6
#393090000000
1!
1%
1-
12
#393100000000
0!
0%
b111 *
0-
02
b111 6
#393110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#393120000000
0!
0%
b0 *
0-
02
b0 6
#393130000000
1!
1%
1-
12
#393140000000
0!
0%
b1 *
0-
02
b1 6
#393150000000
1!
1%
1-
12
#393160000000
0!
0%
b10 *
0-
02
b10 6
#393170000000
1!
1%
1-
12
#393180000000
0!
0%
b11 *
0-
02
b11 6
#393190000000
1!
1%
1-
12
15
#393200000000
0!
0%
b100 *
0-
02
b100 6
#393210000000
1!
1%
1-
12
#393220000000
0!
0%
b101 *
0-
02
b101 6
#393230000000
1!
1%
1-
12
#393240000000
0!
0%
b110 *
0-
02
b110 6
#393250000000
1!
1%
1-
12
#393260000000
0!
0%
b111 *
0-
02
b111 6
#393270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#393280000000
0!
0%
b0 *
0-
02
b0 6
#393290000000
1!
1%
1-
12
#393300000000
0!
0%
b1 *
0-
02
b1 6
#393310000000
1!
1%
1-
12
#393320000000
0!
0%
b10 *
0-
02
b10 6
#393330000000
1!
1%
1-
12
#393340000000
0!
0%
b11 *
0-
02
b11 6
#393350000000
1!
1%
1-
12
15
#393360000000
0!
0%
b100 *
0-
02
b100 6
#393370000000
1!
1%
1-
12
#393380000000
0!
0%
b101 *
0-
02
b101 6
#393390000000
1!
1%
1-
12
#393400000000
0!
0%
b110 *
0-
02
b110 6
#393410000000
1!
1%
1-
12
#393420000000
0!
0%
b111 *
0-
02
b111 6
#393430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#393440000000
0!
0%
b0 *
0-
02
b0 6
#393450000000
1!
1%
1-
12
#393460000000
0!
0%
b1 *
0-
02
b1 6
#393470000000
1!
1%
1-
12
#393480000000
0!
0%
b10 *
0-
02
b10 6
#393490000000
1!
1%
1-
12
#393500000000
0!
0%
b11 *
0-
02
b11 6
#393510000000
1!
1%
1-
12
15
#393520000000
0!
0%
b100 *
0-
02
b100 6
#393530000000
1!
1%
1-
12
#393540000000
0!
0%
b101 *
0-
02
b101 6
#393550000000
1!
1%
1-
12
#393560000000
0!
0%
b110 *
0-
02
b110 6
#393570000000
1!
1%
1-
12
#393580000000
0!
0%
b111 *
0-
02
b111 6
#393590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#393600000000
0!
0%
b0 *
0-
02
b0 6
#393610000000
1!
1%
1-
12
#393620000000
0!
0%
b1 *
0-
02
b1 6
#393630000000
1!
1%
1-
12
#393640000000
0!
0%
b10 *
0-
02
b10 6
#393650000000
1!
1%
1-
12
#393660000000
0!
0%
b11 *
0-
02
b11 6
#393670000000
1!
1%
1-
12
15
#393680000000
0!
0%
b100 *
0-
02
b100 6
#393690000000
1!
1%
1-
12
#393700000000
0!
0%
b101 *
0-
02
b101 6
#393710000000
1!
1%
1-
12
#393720000000
0!
0%
b110 *
0-
02
b110 6
#393730000000
1!
1%
1-
12
#393740000000
0!
0%
b111 *
0-
02
b111 6
#393750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#393760000000
0!
0%
b0 *
0-
02
b0 6
#393770000000
1!
1%
1-
12
#393780000000
0!
0%
b1 *
0-
02
b1 6
#393790000000
1!
1%
1-
12
#393800000000
0!
0%
b10 *
0-
02
b10 6
#393810000000
1!
1%
1-
12
#393820000000
0!
0%
b11 *
0-
02
b11 6
#393830000000
1!
1%
1-
12
15
#393840000000
0!
0%
b100 *
0-
02
b100 6
#393850000000
1!
1%
1-
12
#393860000000
0!
0%
b101 *
0-
02
b101 6
#393870000000
1!
1%
1-
12
#393880000000
0!
0%
b110 *
0-
02
b110 6
#393890000000
1!
1%
1-
12
#393900000000
0!
0%
b111 *
0-
02
b111 6
#393910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#393920000000
0!
0%
b0 *
0-
02
b0 6
#393930000000
1!
1%
1-
12
#393940000000
0!
0%
b1 *
0-
02
b1 6
#393950000000
1!
1%
1-
12
#393960000000
0!
0%
b10 *
0-
02
b10 6
#393970000000
1!
1%
1-
12
#393980000000
0!
0%
b11 *
0-
02
b11 6
#393990000000
1!
1%
1-
12
15
#394000000000
0!
0%
b100 *
0-
02
b100 6
#394010000000
1!
1%
1-
12
#394020000000
0!
0%
b101 *
0-
02
b101 6
#394030000000
1!
1%
1-
12
#394040000000
0!
0%
b110 *
0-
02
b110 6
#394050000000
1!
1%
1-
12
#394060000000
0!
0%
b111 *
0-
02
b111 6
#394070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#394080000000
0!
0%
b0 *
0-
02
b0 6
#394090000000
1!
1%
1-
12
#394100000000
0!
0%
b1 *
0-
02
b1 6
#394110000000
1!
1%
1-
12
#394120000000
0!
0%
b10 *
0-
02
b10 6
#394130000000
1!
1%
1-
12
#394140000000
0!
0%
b11 *
0-
02
b11 6
#394150000000
1!
1%
1-
12
15
#394160000000
0!
0%
b100 *
0-
02
b100 6
#394170000000
1!
1%
1-
12
#394180000000
0!
0%
b101 *
0-
02
b101 6
#394190000000
1!
1%
1-
12
#394200000000
0!
0%
b110 *
0-
02
b110 6
#394210000000
1!
1%
1-
12
#394220000000
0!
0%
b111 *
0-
02
b111 6
#394230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#394240000000
0!
0%
b0 *
0-
02
b0 6
#394250000000
1!
1%
1-
12
#394260000000
0!
0%
b1 *
0-
02
b1 6
#394270000000
1!
1%
1-
12
#394280000000
0!
0%
b10 *
0-
02
b10 6
#394290000000
1!
1%
1-
12
#394300000000
0!
0%
b11 *
0-
02
b11 6
#394310000000
1!
1%
1-
12
15
#394320000000
0!
0%
b100 *
0-
02
b100 6
#394330000000
1!
1%
1-
12
#394340000000
0!
0%
b101 *
0-
02
b101 6
#394350000000
1!
1%
1-
12
#394360000000
0!
0%
b110 *
0-
02
b110 6
#394370000000
1!
1%
1-
12
#394380000000
0!
0%
b111 *
0-
02
b111 6
#394390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#394400000000
0!
0%
b0 *
0-
02
b0 6
#394410000000
1!
1%
1-
12
#394420000000
0!
0%
b1 *
0-
02
b1 6
#394430000000
1!
1%
1-
12
#394440000000
0!
0%
b10 *
0-
02
b10 6
#394450000000
1!
1%
1-
12
#394460000000
0!
0%
b11 *
0-
02
b11 6
#394470000000
1!
1%
1-
12
15
#394480000000
0!
0%
b100 *
0-
02
b100 6
#394490000000
1!
1%
1-
12
#394500000000
0!
0%
b101 *
0-
02
b101 6
#394510000000
1!
1%
1-
12
#394520000000
0!
0%
b110 *
0-
02
b110 6
#394530000000
1!
1%
1-
12
#394540000000
0!
0%
b111 *
0-
02
b111 6
#394550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#394560000000
0!
0%
b0 *
0-
02
b0 6
#394570000000
1!
1%
1-
12
#394580000000
0!
0%
b1 *
0-
02
b1 6
#394590000000
1!
1%
1-
12
#394600000000
0!
0%
b10 *
0-
02
b10 6
#394610000000
1!
1%
1-
12
#394620000000
0!
0%
b11 *
0-
02
b11 6
#394630000000
1!
1%
1-
12
15
#394640000000
0!
0%
b100 *
0-
02
b100 6
#394650000000
1!
1%
1-
12
#394660000000
0!
0%
b101 *
0-
02
b101 6
#394670000000
1!
1%
1-
12
#394680000000
0!
0%
b110 *
0-
02
b110 6
#394690000000
1!
1%
1-
12
#394700000000
0!
0%
b111 *
0-
02
b111 6
#394710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#394720000000
0!
0%
b0 *
0-
02
b0 6
#394730000000
1!
1%
1-
12
#394740000000
0!
0%
b1 *
0-
02
b1 6
#394750000000
1!
1%
1-
12
#394760000000
0!
0%
b10 *
0-
02
b10 6
#394770000000
1!
1%
1-
12
#394780000000
0!
0%
b11 *
0-
02
b11 6
#394790000000
1!
1%
1-
12
15
#394800000000
0!
0%
b100 *
0-
02
b100 6
#394810000000
1!
1%
1-
12
#394820000000
0!
0%
b101 *
0-
02
b101 6
#394830000000
1!
1%
1-
12
#394840000000
0!
0%
b110 *
0-
02
b110 6
#394850000000
1!
1%
1-
12
#394860000000
0!
0%
b111 *
0-
02
b111 6
#394870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#394880000000
0!
0%
b0 *
0-
02
b0 6
#394890000000
1!
1%
1-
12
#394900000000
0!
0%
b1 *
0-
02
b1 6
#394910000000
1!
1%
1-
12
#394920000000
0!
0%
b10 *
0-
02
b10 6
#394930000000
1!
1%
1-
12
#394940000000
0!
0%
b11 *
0-
02
b11 6
#394950000000
1!
1%
1-
12
15
#394960000000
0!
0%
b100 *
0-
02
b100 6
#394970000000
1!
1%
1-
12
#394980000000
0!
0%
b101 *
0-
02
b101 6
#394990000000
1!
1%
1-
12
#395000000000
0!
0%
b110 *
0-
02
b110 6
#395010000000
1!
1%
1-
12
#395020000000
0!
0%
b111 *
0-
02
b111 6
#395030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#395040000000
0!
0%
b0 *
0-
02
b0 6
#395050000000
1!
1%
1-
12
#395060000000
0!
0%
b1 *
0-
02
b1 6
#395070000000
1!
1%
1-
12
#395080000000
0!
0%
b10 *
0-
02
b10 6
#395090000000
1!
1%
1-
12
#395100000000
0!
0%
b11 *
0-
02
b11 6
#395110000000
1!
1%
1-
12
15
#395120000000
0!
0%
b100 *
0-
02
b100 6
#395130000000
1!
1%
1-
12
#395140000000
0!
0%
b101 *
0-
02
b101 6
#395150000000
1!
1%
1-
12
#395160000000
0!
0%
b110 *
0-
02
b110 6
#395170000000
1!
1%
1-
12
#395180000000
0!
0%
b111 *
0-
02
b111 6
#395190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#395200000000
0!
0%
b0 *
0-
02
b0 6
#395210000000
1!
1%
1-
12
#395220000000
0!
0%
b1 *
0-
02
b1 6
#395230000000
1!
1%
1-
12
#395240000000
0!
0%
b10 *
0-
02
b10 6
#395250000000
1!
1%
1-
12
#395260000000
0!
0%
b11 *
0-
02
b11 6
#395270000000
1!
1%
1-
12
15
#395280000000
0!
0%
b100 *
0-
02
b100 6
#395290000000
1!
1%
1-
12
#395300000000
0!
0%
b101 *
0-
02
b101 6
#395310000000
1!
1%
1-
12
#395320000000
0!
0%
b110 *
0-
02
b110 6
#395330000000
1!
1%
1-
12
#395340000000
0!
0%
b111 *
0-
02
b111 6
#395350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#395360000000
0!
0%
b0 *
0-
02
b0 6
#395370000000
1!
1%
1-
12
#395380000000
0!
0%
b1 *
0-
02
b1 6
#395390000000
1!
1%
1-
12
#395400000000
0!
0%
b10 *
0-
02
b10 6
#395410000000
1!
1%
1-
12
#395420000000
0!
0%
b11 *
0-
02
b11 6
#395430000000
1!
1%
1-
12
15
#395440000000
0!
0%
b100 *
0-
02
b100 6
#395450000000
1!
1%
1-
12
#395460000000
0!
0%
b101 *
0-
02
b101 6
#395470000000
1!
1%
1-
12
#395480000000
0!
0%
b110 *
0-
02
b110 6
#395490000000
1!
1%
1-
12
#395500000000
0!
0%
b111 *
0-
02
b111 6
#395510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#395520000000
0!
0%
b0 *
0-
02
b0 6
#395530000000
1!
1%
1-
12
#395540000000
0!
0%
b1 *
0-
02
b1 6
#395550000000
1!
1%
1-
12
#395560000000
0!
0%
b10 *
0-
02
b10 6
#395570000000
1!
1%
1-
12
#395580000000
0!
0%
b11 *
0-
02
b11 6
#395590000000
1!
1%
1-
12
15
#395600000000
0!
0%
b100 *
0-
02
b100 6
#395610000000
1!
1%
1-
12
#395620000000
0!
0%
b101 *
0-
02
b101 6
#395630000000
1!
1%
1-
12
#395640000000
0!
0%
b110 *
0-
02
b110 6
#395650000000
1!
1%
1-
12
#395660000000
0!
0%
b111 *
0-
02
b111 6
#395670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#395680000000
0!
0%
b0 *
0-
02
b0 6
#395690000000
1!
1%
1-
12
#395700000000
0!
0%
b1 *
0-
02
b1 6
#395710000000
1!
1%
1-
12
#395720000000
0!
0%
b10 *
0-
02
b10 6
#395730000000
1!
1%
1-
12
#395740000000
0!
0%
b11 *
0-
02
b11 6
#395750000000
1!
1%
1-
12
15
#395760000000
0!
0%
b100 *
0-
02
b100 6
#395770000000
1!
1%
1-
12
#395780000000
0!
0%
b101 *
0-
02
b101 6
#395790000000
1!
1%
1-
12
#395800000000
0!
0%
b110 *
0-
02
b110 6
#395810000000
1!
1%
1-
12
#395820000000
0!
0%
b111 *
0-
02
b111 6
#395830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#395840000000
0!
0%
b0 *
0-
02
b0 6
#395850000000
1!
1%
1-
12
#395860000000
0!
0%
b1 *
0-
02
b1 6
#395870000000
1!
1%
1-
12
#395880000000
0!
0%
b10 *
0-
02
b10 6
#395890000000
1!
1%
1-
12
#395900000000
0!
0%
b11 *
0-
02
b11 6
#395910000000
1!
1%
1-
12
15
#395920000000
0!
0%
b100 *
0-
02
b100 6
#395930000000
1!
1%
1-
12
#395940000000
0!
0%
b101 *
0-
02
b101 6
#395950000000
1!
1%
1-
12
#395960000000
0!
0%
b110 *
0-
02
b110 6
#395970000000
1!
1%
1-
12
#395980000000
0!
0%
b111 *
0-
02
b111 6
#395990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#396000000000
0!
0%
b0 *
0-
02
b0 6
#396010000000
1!
1%
1-
12
#396020000000
0!
0%
b1 *
0-
02
b1 6
#396030000000
1!
1%
1-
12
#396040000000
0!
0%
b10 *
0-
02
b10 6
#396050000000
1!
1%
1-
12
#396060000000
0!
0%
b11 *
0-
02
b11 6
#396070000000
1!
1%
1-
12
15
#396080000000
0!
0%
b100 *
0-
02
b100 6
#396090000000
1!
1%
1-
12
#396100000000
0!
0%
b101 *
0-
02
b101 6
#396110000000
1!
1%
1-
12
#396120000000
0!
0%
b110 *
0-
02
b110 6
#396130000000
1!
1%
1-
12
#396140000000
0!
0%
b111 *
0-
02
b111 6
#396150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#396160000000
0!
0%
b0 *
0-
02
b0 6
#396170000000
1!
1%
1-
12
#396180000000
0!
0%
b1 *
0-
02
b1 6
#396190000000
1!
1%
1-
12
#396200000000
0!
0%
b10 *
0-
02
b10 6
#396210000000
1!
1%
1-
12
#396220000000
0!
0%
b11 *
0-
02
b11 6
#396230000000
1!
1%
1-
12
15
#396240000000
0!
0%
b100 *
0-
02
b100 6
#396250000000
1!
1%
1-
12
#396260000000
0!
0%
b101 *
0-
02
b101 6
#396270000000
1!
1%
1-
12
#396280000000
0!
0%
b110 *
0-
02
b110 6
#396290000000
1!
1%
1-
12
#396300000000
0!
0%
b111 *
0-
02
b111 6
#396310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#396320000000
0!
0%
b0 *
0-
02
b0 6
#396330000000
1!
1%
1-
12
#396340000000
0!
0%
b1 *
0-
02
b1 6
#396350000000
1!
1%
1-
12
#396360000000
0!
0%
b10 *
0-
02
b10 6
#396370000000
1!
1%
1-
12
#396380000000
0!
0%
b11 *
0-
02
b11 6
#396390000000
1!
1%
1-
12
15
#396400000000
0!
0%
b100 *
0-
02
b100 6
#396410000000
1!
1%
1-
12
#396420000000
0!
0%
b101 *
0-
02
b101 6
#396430000000
1!
1%
1-
12
#396440000000
0!
0%
b110 *
0-
02
b110 6
#396450000000
1!
1%
1-
12
#396460000000
0!
0%
b111 *
0-
02
b111 6
#396470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#396480000000
0!
0%
b0 *
0-
02
b0 6
#396490000000
1!
1%
1-
12
#396500000000
0!
0%
b1 *
0-
02
b1 6
#396510000000
1!
1%
1-
12
#396520000000
0!
0%
b10 *
0-
02
b10 6
#396530000000
1!
1%
1-
12
#396540000000
0!
0%
b11 *
0-
02
b11 6
#396550000000
1!
1%
1-
12
15
#396560000000
0!
0%
b100 *
0-
02
b100 6
#396570000000
1!
1%
1-
12
#396580000000
0!
0%
b101 *
0-
02
b101 6
#396590000000
1!
1%
1-
12
#396600000000
0!
0%
b110 *
0-
02
b110 6
#396610000000
1!
1%
1-
12
#396620000000
0!
0%
b111 *
0-
02
b111 6
#396630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#396640000000
0!
0%
b0 *
0-
02
b0 6
#396650000000
1!
1%
1-
12
#396660000000
0!
0%
b1 *
0-
02
b1 6
#396670000000
1!
1%
1-
12
#396680000000
0!
0%
b10 *
0-
02
b10 6
#396690000000
1!
1%
1-
12
#396700000000
0!
0%
b11 *
0-
02
b11 6
#396710000000
1!
1%
1-
12
15
#396720000000
0!
0%
b100 *
0-
02
b100 6
#396730000000
1!
1%
1-
12
#396740000000
0!
0%
b101 *
0-
02
b101 6
#396750000000
1!
1%
1-
12
#396760000000
0!
0%
b110 *
0-
02
b110 6
#396770000000
1!
1%
1-
12
#396780000000
0!
0%
b111 *
0-
02
b111 6
#396790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#396800000000
0!
0%
b0 *
0-
02
b0 6
#396810000000
1!
1%
1-
12
#396820000000
0!
0%
b1 *
0-
02
b1 6
#396830000000
1!
1%
1-
12
#396840000000
0!
0%
b10 *
0-
02
b10 6
#396850000000
1!
1%
1-
12
#396860000000
0!
0%
b11 *
0-
02
b11 6
#396870000000
1!
1%
1-
12
15
#396880000000
0!
0%
b100 *
0-
02
b100 6
#396890000000
1!
1%
1-
12
#396900000000
0!
0%
b101 *
0-
02
b101 6
#396910000000
1!
1%
1-
12
#396920000000
0!
0%
b110 *
0-
02
b110 6
#396930000000
1!
1%
1-
12
#396940000000
0!
0%
b111 *
0-
02
b111 6
#396950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#396960000000
0!
0%
b0 *
0-
02
b0 6
#396970000000
1!
1%
1-
12
#396980000000
0!
0%
b1 *
0-
02
b1 6
#396990000000
1!
1%
1-
12
#397000000000
0!
0%
b10 *
0-
02
b10 6
#397010000000
1!
1%
1-
12
#397020000000
0!
0%
b11 *
0-
02
b11 6
#397030000000
1!
1%
1-
12
15
#397040000000
0!
0%
b100 *
0-
02
b100 6
#397050000000
1!
1%
1-
12
#397060000000
0!
0%
b101 *
0-
02
b101 6
#397070000000
1!
1%
1-
12
#397080000000
0!
0%
b110 *
0-
02
b110 6
#397090000000
1!
1%
1-
12
#397100000000
0!
0%
b111 *
0-
02
b111 6
#397110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#397120000000
0!
0%
b0 *
0-
02
b0 6
#397130000000
1!
1%
1-
12
#397140000000
0!
0%
b1 *
0-
02
b1 6
#397150000000
1!
1%
1-
12
#397160000000
0!
0%
b10 *
0-
02
b10 6
#397170000000
1!
1%
1-
12
#397180000000
0!
0%
b11 *
0-
02
b11 6
#397190000000
1!
1%
1-
12
15
#397200000000
0!
0%
b100 *
0-
02
b100 6
#397210000000
1!
1%
1-
12
#397220000000
0!
0%
b101 *
0-
02
b101 6
#397230000000
1!
1%
1-
12
#397240000000
0!
0%
b110 *
0-
02
b110 6
#397250000000
1!
1%
1-
12
#397260000000
0!
0%
b111 *
0-
02
b111 6
#397270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#397280000000
0!
0%
b0 *
0-
02
b0 6
#397290000000
1!
1%
1-
12
#397300000000
0!
0%
b1 *
0-
02
b1 6
#397310000000
1!
1%
1-
12
#397320000000
0!
0%
b10 *
0-
02
b10 6
#397330000000
1!
1%
1-
12
#397340000000
0!
0%
b11 *
0-
02
b11 6
#397350000000
1!
1%
1-
12
15
#397360000000
0!
0%
b100 *
0-
02
b100 6
#397370000000
1!
1%
1-
12
#397380000000
0!
0%
b101 *
0-
02
b101 6
#397390000000
1!
1%
1-
12
#397400000000
0!
0%
b110 *
0-
02
b110 6
#397410000000
1!
1%
1-
12
#397420000000
0!
0%
b111 *
0-
02
b111 6
#397430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#397440000000
0!
0%
b0 *
0-
02
b0 6
#397450000000
1!
1%
1-
12
#397460000000
0!
0%
b1 *
0-
02
b1 6
#397470000000
1!
1%
1-
12
#397480000000
0!
0%
b10 *
0-
02
b10 6
#397490000000
1!
1%
1-
12
#397500000000
0!
0%
b11 *
0-
02
b11 6
#397510000000
1!
1%
1-
12
15
#397520000000
0!
0%
b100 *
0-
02
b100 6
#397530000000
1!
1%
1-
12
#397540000000
0!
0%
b101 *
0-
02
b101 6
#397550000000
1!
1%
1-
12
#397560000000
0!
0%
b110 *
0-
02
b110 6
#397570000000
1!
1%
1-
12
#397580000000
0!
0%
b111 *
0-
02
b111 6
#397590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#397600000000
0!
0%
b0 *
0-
02
b0 6
#397610000000
1!
1%
1-
12
#397620000000
0!
0%
b1 *
0-
02
b1 6
#397630000000
1!
1%
1-
12
#397640000000
0!
0%
b10 *
0-
02
b10 6
#397650000000
1!
1%
1-
12
#397660000000
0!
0%
b11 *
0-
02
b11 6
#397670000000
1!
1%
1-
12
15
#397680000000
0!
0%
b100 *
0-
02
b100 6
#397690000000
1!
1%
1-
12
#397700000000
0!
0%
b101 *
0-
02
b101 6
#397710000000
1!
1%
1-
12
#397720000000
0!
0%
b110 *
0-
02
b110 6
#397730000000
1!
1%
1-
12
#397740000000
0!
0%
b111 *
0-
02
b111 6
#397750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#397760000000
0!
0%
b0 *
0-
02
b0 6
#397770000000
1!
1%
1-
12
#397780000000
0!
0%
b1 *
0-
02
b1 6
#397790000000
1!
1%
1-
12
#397800000000
0!
0%
b10 *
0-
02
b10 6
#397810000000
1!
1%
1-
12
#397820000000
0!
0%
b11 *
0-
02
b11 6
#397830000000
1!
1%
1-
12
15
#397840000000
0!
0%
b100 *
0-
02
b100 6
#397850000000
1!
1%
1-
12
#397860000000
0!
0%
b101 *
0-
02
b101 6
#397870000000
1!
1%
1-
12
#397880000000
0!
0%
b110 *
0-
02
b110 6
#397890000000
1!
1%
1-
12
#397900000000
0!
0%
b111 *
0-
02
b111 6
#397910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#397920000000
0!
0%
b0 *
0-
02
b0 6
#397930000000
1!
1%
1-
12
#397940000000
0!
0%
b1 *
0-
02
b1 6
#397950000000
1!
1%
1-
12
#397960000000
0!
0%
b10 *
0-
02
b10 6
#397970000000
1!
1%
1-
12
#397980000000
0!
0%
b11 *
0-
02
b11 6
#397990000000
1!
1%
1-
12
15
#398000000000
0!
0%
b100 *
0-
02
b100 6
#398010000000
1!
1%
1-
12
#398020000000
0!
0%
b101 *
0-
02
b101 6
#398030000000
1!
1%
1-
12
#398040000000
0!
0%
b110 *
0-
02
b110 6
#398050000000
1!
1%
1-
12
#398060000000
0!
0%
b111 *
0-
02
b111 6
#398070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#398080000000
0!
0%
b0 *
0-
02
b0 6
#398090000000
1!
1%
1-
12
#398100000000
0!
0%
b1 *
0-
02
b1 6
#398110000000
1!
1%
1-
12
#398120000000
0!
0%
b10 *
0-
02
b10 6
#398130000000
1!
1%
1-
12
#398140000000
0!
0%
b11 *
0-
02
b11 6
#398150000000
1!
1%
1-
12
15
#398160000000
0!
0%
b100 *
0-
02
b100 6
#398170000000
1!
1%
1-
12
#398180000000
0!
0%
b101 *
0-
02
b101 6
#398190000000
1!
1%
1-
12
#398200000000
0!
0%
b110 *
0-
02
b110 6
#398210000000
1!
1%
1-
12
#398220000000
0!
0%
b111 *
0-
02
b111 6
#398230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#398240000000
0!
0%
b0 *
0-
02
b0 6
#398250000000
1!
1%
1-
12
#398260000000
0!
0%
b1 *
0-
02
b1 6
#398270000000
1!
1%
1-
12
#398280000000
0!
0%
b10 *
0-
02
b10 6
#398290000000
1!
1%
1-
12
#398300000000
0!
0%
b11 *
0-
02
b11 6
#398310000000
1!
1%
1-
12
15
#398320000000
0!
0%
b100 *
0-
02
b100 6
#398330000000
1!
1%
1-
12
#398340000000
0!
0%
b101 *
0-
02
b101 6
#398350000000
1!
1%
1-
12
#398360000000
0!
0%
b110 *
0-
02
b110 6
#398370000000
1!
1%
1-
12
#398380000000
0!
0%
b111 *
0-
02
b111 6
#398390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#398400000000
0!
0%
b0 *
0-
02
b0 6
#398410000000
1!
1%
1-
12
#398420000000
0!
0%
b1 *
0-
02
b1 6
#398430000000
1!
1%
1-
12
#398440000000
0!
0%
b10 *
0-
02
b10 6
#398450000000
1!
1%
1-
12
#398460000000
0!
0%
b11 *
0-
02
b11 6
#398470000000
1!
1%
1-
12
15
#398480000000
0!
0%
b100 *
0-
02
b100 6
#398490000000
1!
1%
1-
12
#398500000000
0!
0%
b101 *
0-
02
b101 6
#398510000000
1!
1%
1-
12
#398520000000
0!
0%
b110 *
0-
02
b110 6
#398530000000
1!
1%
1-
12
#398540000000
0!
0%
b111 *
0-
02
b111 6
#398550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#398560000000
0!
0%
b0 *
0-
02
b0 6
#398570000000
1!
1%
1-
12
#398580000000
0!
0%
b1 *
0-
02
b1 6
#398590000000
1!
1%
1-
12
#398600000000
0!
0%
b10 *
0-
02
b10 6
#398610000000
1!
1%
1-
12
#398620000000
0!
0%
b11 *
0-
02
b11 6
#398630000000
1!
1%
1-
12
15
#398640000000
0!
0%
b100 *
0-
02
b100 6
#398650000000
1!
1%
1-
12
#398660000000
0!
0%
b101 *
0-
02
b101 6
#398670000000
1!
1%
1-
12
#398680000000
0!
0%
b110 *
0-
02
b110 6
#398690000000
1!
1%
1-
12
#398700000000
0!
0%
b111 *
0-
02
b111 6
#398710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#398720000000
0!
0%
b0 *
0-
02
b0 6
#398730000000
1!
1%
1-
12
#398740000000
0!
0%
b1 *
0-
02
b1 6
#398750000000
1!
1%
1-
12
#398760000000
0!
0%
b10 *
0-
02
b10 6
#398770000000
1!
1%
1-
12
#398780000000
0!
0%
b11 *
0-
02
b11 6
#398790000000
1!
1%
1-
12
15
#398800000000
0!
0%
b100 *
0-
02
b100 6
#398810000000
1!
1%
1-
12
#398820000000
0!
0%
b101 *
0-
02
b101 6
#398830000000
1!
1%
1-
12
#398840000000
0!
0%
b110 *
0-
02
b110 6
#398850000000
1!
1%
1-
12
#398860000000
0!
0%
b111 *
0-
02
b111 6
#398870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#398880000000
0!
0%
b0 *
0-
02
b0 6
#398890000000
1!
1%
1-
12
#398900000000
0!
0%
b1 *
0-
02
b1 6
#398910000000
1!
1%
1-
12
#398920000000
0!
0%
b10 *
0-
02
b10 6
#398930000000
1!
1%
1-
12
#398940000000
0!
0%
b11 *
0-
02
b11 6
#398950000000
1!
1%
1-
12
15
#398960000000
0!
0%
b100 *
0-
02
b100 6
#398970000000
1!
1%
1-
12
#398980000000
0!
0%
b101 *
0-
02
b101 6
#398990000000
1!
1%
1-
12
#399000000000
0!
0%
b110 *
0-
02
b110 6
#399010000000
1!
1%
1-
12
#399020000000
0!
0%
b111 *
0-
02
b111 6
#399030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#399040000000
0!
0%
b0 *
0-
02
b0 6
#399050000000
1!
1%
1-
12
#399060000000
0!
0%
b1 *
0-
02
b1 6
#399070000000
1!
1%
1-
12
#399080000000
0!
0%
b10 *
0-
02
b10 6
#399090000000
1!
1%
1-
12
#399100000000
0!
0%
b11 *
0-
02
b11 6
#399110000000
1!
1%
1-
12
15
#399120000000
0!
0%
b100 *
0-
02
b100 6
#399130000000
1!
1%
1-
12
#399140000000
0!
0%
b101 *
0-
02
b101 6
#399150000000
1!
1%
1-
12
#399160000000
0!
0%
b110 *
0-
02
b110 6
#399170000000
1!
1%
1-
12
#399180000000
0!
0%
b111 *
0-
02
b111 6
#399190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#399200000000
0!
0%
b0 *
0-
02
b0 6
#399210000000
1!
1%
1-
12
#399220000000
0!
0%
b1 *
0-
02
b1 6
#399230000000
1!
1%
1-
12
#399240000000
0!
0%
b10 *
0-
02
b10 6
#399250000000
1!
1%
1-
12
#399260000000
0!
0%
b11 *
0-
02
b11 6
#399270000000
1!
1%
1-
12
15
#399280000000
0!
0%
b100 *
0-
02
b100 6
#399290000000
1!
1%
1-
12
#399300000000
0!
0%
b101 *
0-
02
b101 6
#399310000000
1!
1%
1-
12
#399320000000
0!
0%
b110 *
0-
02
b110 6
#399330000000
1!
1%
1-
12
#399340000000
0!
0%
b111 *
0-
02
b111 6
#399350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#399360000000
0!
0%
b0 *
0-
02
b0 6
#399370000000
1!
1%
1-
12
#399380000000
0!
0%
b1 *
0-
02
b1 6
#399390000000
1!
1%
1-
12
#399400000000
0!
0%
b10 *
0-
02
b10 6
#399410000000
1!
1%
1-
12
#399420000000
0!
0%
b11 *
0-
02
b11 6
#399430000000
1!
1%
1-
12
15
#399440000000
0!
0%
b100 *
0-
02
b100 6
#399450000000
1!
1%
1-
12
#399460000000
0!
0%
b101 *
0-
02
b101 6
#399470000000
1!
1%
1-
12
#399480000000
0!
0%
b110 *
0-
02
b110 6
#399490000000
1!
1%
1-
12
#399500000000
0!
0%
b111 *
0-
02
b111 6
#399510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#399520000000
0!
0%
b0 *
0-
02
b0 6
#399530000000
1!
1%
1-
12
#399540000000
0!
0%
b1 *
0-
02
b1 6
#399550000000
1!
1%
1-
12
#399560000000
0!
0%
b10 *
0-
02
b10 6
#399570000000
1!
1%
1-
12
#399580000000
0!
0%
b11 *
0-
02
b11 6
#399590000000
1!
1%
1-
12
15
#399600000000
0!
0%
b100 *
0-
02
b100 6
#399610000000
1!
1%
1-
12
#399620000000
0!
0%
b101 *
0-
02
b101 6
#399630000000
1!
1%
1-
12
#399640000000
0!
0%
b110 *
0-
02
b110 6
#399650000000
1!
1%
1-
12
#399660000000
0!
0%
b111 *
0-
02
b111 6
#399670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#399680000000
0!
0%
b0 *
0-
02
b0 6
#399690000000
1!
1%
1-
12
#399700000000
0!
0%
b1 *
0-
02
b1 6
#399710000000
1!
1%
1-
12
#399720000000
0!
0%
b10 *
0-
02
b10 6
#399730000000
1!
1%
1-
12
#399740000000
0!
0%
b11 *
0-
02
b11 6
#399750000000
1!
1%
1-
12
15
#399760000000
0!
0%
b100 *
0-
02
b100 6
#399770000000
1!
1%
1-
12
#399780000000
0!
0%
b101 *
0-
02
b101 6
#399790000000
1!
1%
1-
12
#399800000000
0!
0%
b110 *
0-
02
b110 6
#399810000000
1!
1%
1-
12
#399820000000
0!
0%
b111 *
0-
02
b111 6
#399830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#399840000000
0!
0%
b0 *
0-
02
b0 6
#399850000000
1!
1%
1-
12
#399860000000
0!
0%
b1 *
0-
02
b1 6
#399870000000
1!
1%
1-
12
#399880000000
0!
0%
b10 *
0-
02
b10 6
#399890000000
1!
1%
1-
12
#399900000000
0!
0%
b11 *
0-
02
b11 6
#399910000000
1!
1%
1-
12
15
#399920000000
0!
0%
b100 *
0-
02
b100 6
#399930000000
1!
1%
1-
12
#399940000000
0!
0%
b101 *
0-
02
b101 6
#399950000000
1!
1%
1-
12
#399960000000
0!
0%
b110 *
0-
02
b110 6
#399970000000
1!
1%
1-
12
#399980000000
0!
0%
b111 *
0-
02
b111 6
#399990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#400000000000
0!
0%
b0 *
0-
02
b0 6
#400010000000
1!
1%
1-
12
#400020000000
0!
0%
b1 *
0-
02
b1 6
#400030000000
1!
1%
1-
12
#400040000000
0!
0%
b10 *
0-
02
b10 6
#400050000000
1!
1%
1-
12
#400060000000
0!
0%
b11 *
0-
02
b11 6
#400070000000
1!
1%
1-
12
15
#400080000000
0!
0%
b100 *
0-
02
b100 6
#400090000000
1!
1%
1-
12
#400100000000
0!
0%
b101 *
0-
02
b101 6
#400110000000
1!
1%
1-
12
#400120000000
0!
0%
b110 *
0-
02
b110 6
#400130000000
1!
1%
1-
12
#400140000000
0!
0%
b111 *
0-
02
b111 6
#400150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#400160000000
0!
0%
b0 *
0-
02
b0 6
#400170000000
1!
1%
1-
12
#400180000000
0!
0%
b1 *
0-
02
b1 6
#400190000000
1!
1%
1-
12
#400200000000
0!
0%
b10 *
0-
02
b10 6
#400210000000
1!
1%
1-
12
#400220000000
0!
0%
b11 *
0-
02
b11 6
#400230000000
1!
1%
1-
12
15
#400240000000
0!
0%
b100 *
0-
02
b100 6
#400250000000
1!
1%
1-
12
#400260000000
0!
0%
b101 *
0-
02
b101 6
#400270000000
1!
1%
1-
12
#400280000000
0!
0%
b110 *
0-
02
b110 6
#400290000000
1!
1%
1-
12
#400300000000
0!
0%
b111 *
0-
02
b111 6
#400310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#400320000000
0!
0%
b0 *
0-
02
b0 6
#400330000000
1!
1%
1-
12
#400340000000
0!
0%
b1 *
0-
02
b1 6
#400350000000
1!
1%
1-
12
#400360000000
0!
0%
b10 *
0-
02
b10 6
#400370000000
1!
1%
1-
12
#400380000000
0!
0%
b11 *
0-
02
b11 6
#400390000000
1!
1%
1-
12
15
#400400000000
0!
0%
b100 *
0-
02
b100 6
#400410000000
1!
1%
1-
12
#400420000000
0!
0%
b101 *
0-
02
b101 6
#400430000000
1!
1%
1-
12
#400440000000
0!
0%
b110 *
0-
02
b110 6
#400450000000
1!
1%
1-
12
#400460000000
0!
0%
b111 *
0-
02
b111 6
#400470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#400480000000
0!
0%
b0 *
0-
02
b0 6
#400490000000
1!
1%
1-
12
#400500000000
0!
0%
b1 *
0-
02
b1 6
#400510000000
1!
1%
1-
12
#400520000000
0!
0%
b10 *
0-
02
b10 6
#400530000000
1!
1%
1-
12
#400540000000
0!
0%
b11 *
0-
02
b11 6
#400550000000
1!
1%
1-
12
15
#400560000000
0!
0%
b100 *
0-
02
b100 6
#400570000000
1!
1%
1-
12
#400580000000
0!
0%
b101 *
0-
02
b101 6
#400590000000
1!
1%
1-
12
#400600000000
0!
0%
b110 *
0-
02
b110 6
#400610000000
1!
1%
1-
12
#400620000000
0!
0%
b111 *
0-
02
b111 6
#400630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#400640000000
0!
0%
b0 *
0-
02
b0 6
#400650000000
1!
1%
1-
12
#400660000000
0!
0%
b1 *
0-
02
b1 6
#400670000000
1!
1%
1-
12
#400680000000
0!
0%
b10 *
0-
02
b10 6
#400690000000
1!
1%
1-
12
#400700000000
0!
0%
b11 *
0-
02
b11 6
#400710000000
1!
1%
1-
12
15
#400720000000
0!
0%
b100 *
0-
02
b100 6
#400730000000
1!
1%
1-
12
#400740000000
0!
0%
b101 *
0-
02
b101 6
#400750000000
1!
1%
1-
12
#400760000000
0!
0%
b110 *
0-
02
b110 6
#400770000000
1!
1%
1-
12
#400780000000
0!
0%
b111 *
0-
02
b111 6
#400790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#400800000000
0!
0%
b0 *
0-
02
b0 6
#400810000000
1!
1%
1-
12
#400820000000
0!
0%
b1 *
0-
02
b1 6
#400830000000
1!
1%
1-
12
#400840000000
0!
0%
b10 *
0-
02
b10 6
#400850000000
1!
1%
1-
12
#400860000000
0!
0%
b11 *
0-
02
b11 6
#400870000000
1!
1%
1-
12
15
#400880000000
0!
0%
b100 *
0-
02
b100 6
#400890000000
1!
1%
1-
12
#400900000000
0!
0%
b101 *
0-
02
b101 6
#400910000000
1!
1%
1-
12
#400920000000
0!
0%
b110 *
0-
02
b110 6
#400930000000
1!
1%
1-
12
#400940000000
0!
0%
b111 *
0-
02
b111 6
#400950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#400960000000
0!
0%
b0 *
0-
02
b0 6
#400970000000
1!
1%
1-
12
#400980000000
0!
0%
b1 *
0-
02
b1 6
#400990000000
1!
1%
1-
12
#401000000000
0!
0%
b10 *
0-
02
b10 6
#401010000000
1!
1%
1-
12
#401020000000
0!
0%
b11 *
0-
02
b11 6
#401030000000
1!
1%
1-
12
15
#401040000000
0!
0%
b100 *
0-
02
b100 6
#401050000000
1!
1%
1-
12
#401060000000
0!
0%
b101 *
0-
02
b101 6
#401070000000
1!
1%
1-
12
#401080000000
0!
0%
b110 *
0-
02
b110 6
#401090000000
1!
1%
1-
12
#401100000000
0!
0%
b111 *
0-
02
b111 6
#401110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#401120000000
0!
0%
b0 *
0-
02
b0 6
#401130000000
1!
1%
1-
12
#401140000000
0!
0%
b1 *
0-
02
b1 6
#401150000000
1!
1%
1-
12
#401160000000
0!
0%
b10 *
0-
02
b10 6
#401170000000
1!
1%
1-
12
#401180000000
0!
0%
b11 *
0-
02
b11 6
#401190000000
1!
1%
1-
12
15
#401200000000
0!
0%
b100 *
0-
02
b100 6
#401210000000
1!
1%
1-
12
#401220000000
0!
0%
b101 *
0-
02
b101 6
#401230000000
1!
1%
1-
12
#401240000000
0!
0%
b110 *
0-
02
b110 6
#401250000000
1!
1%
1-
12
#401260000000
0!
0%
b111 *
0-
02
b111 6
#401270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#401280000000
0!
0%
b0 *
0-
02
b0 6
#401290000000
1!
1%
1-
12
#401300000000
0!
0%
b1 *
0-
02
b1 6
#401310000000
1!
1%
1-
12
#401320000000
0!
0%
b10 *
0-
02
b10 6
#401330000000
1!
1%
1-
12
#401340000000
0!
0%
b11 *
0-
02
b11 6
#401350000000
1!
1%
1-
12
15
#401360000000
0!
0%
b100 *
0-
02
b100 6
#401370000000
1!
1%
1-
12
#401380000000
0!
0%
b101 *
0-
02
b101 6
#401390000000
1!
1%
1-
12
#401400000000
0!
0%
b110 *
0-
02
b110 6
#401410000000
1!
1%
1-
12
#401420000000
0!
0%
b111 *
0-
02
b111 6
#401430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#401440000000
0!
0%
b0 *
0-
02
b0 6
#401450000000
1!
1%
1-
12
#401460000000
0!
0%
b1 *
0-
02
b1 6
#401470000000
1!
1%
1-
12
#401480000000
0!
0%
b10 *
0-
02
b10 6
#401490000000
1!
1%
1-
12
#401500000000
0!
0%
b11 *
0-
02
b11 6
#401510000000
1!
1%
1-
12
15
#401520000000
0!
0%
b100 *
0-
02
b100 6
#401530000000
1!
1%
1-
12
#401540000000
0!
0%
b101 *
0-
02
b101 6
#401550000000
1!
1%
1-
12
#401560000000
0!
0%
b110 *
0-
02
b110 6
#401570000000
1!
1%
1-
12
#401580000000
0!
0%
b111 *
0-
02
b111 6
#401590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#401600000000
0!
0%
b0 *
0-
02
b0 6
#401610000000
1!
1%
1-
12
#401620000000
0!
0%
b1 *
0-
02
b1 6
#401630000000
1!
1%
1-
12
#401640000000
0!
0%
b10 *
0-
02
b10 6
#401650000000
1!
1%
1-
12
#401660000000
0!
0%
b11 *
0-
02
b11 6
#401670000000
1!
1%
1-
12
15
#401680000000
0!
0%
b100 *
0-
02
b100 6
#401690000000
1!
1%
1-
12
#401700000000
0!
0%
b101 *
0-
02
b101 6
#401710000000
1!
1%
1-
12
#401720000000
0!
0%
b110 *
0-
02
b110 6
#401730000000
1!
1%
1-
12
#401740000000
0!
0%
b111 *
0-
02
b111 6
#401750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#401760000000
0!
0%
b0 *
0-
02
b0 6
#401770000000
1!
1%
1-
12
#401780000000
0!
0%
b1 *
0-
02
b1 6
#401790000000
1!
1%
1-
12
#401800000000
0!
0%
b10 *
0-
02
b10 6
#401810000000
1!
1%
1-
12
#401820000000
0!
0%
b11 *
0-
02
b11 6
#401830000000
1!
1%
1-
12
15
#401840000000
0!
0%
b100 *
0-
02
b100 6
#401850000000
1!
1%
1-
12
#401860000000
0!
0%
b101 *
0-
02
b101 6
#401870000000
1!
1%
1-
12
#401880000000
0!
0%
b110 *
0-
02
b110 6
#401890000000
1!
1%
1-
12
#401900000000
0!
0%
b111 *
0-
02
b111 6
#401910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#401920000000
0!
0%
b0 *
0-
02
b0 6
#401930000000
1!
1%
1-
12
#401940000000
0!
0%
b1 *
0-
02
b1 6
#401950000000
1!
1%
1-
12
#401960000000
0!
0%
b10 *
0-
02
b10 6
#401970000000
1!
1%
1-
12
#401980000000
0!
0%
b11 *
0-
02
b11 6
#401990000000
1!
1%
1-
12
15
#402000000000
0!
0%
b100 *
0-
02
b100 6
#402010000000
1!
1%
1-
12
#402020000000
0!
0%
b101 *
0-
02
b101 6
#402030000000
1!
1%
1-
12
#402040000000
0!
0%
b110 *
0-
02
b110 6
#402050000000
1!
1%
1-
12
#402060000000
0!
0%
b111 *
0-
02
b111 6
#402070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#402080000000
0!
0%
b0 *
0-
02
b0 6
#402090000000
1!
1%
1-
12
#402100000000
0!
0%
b1 *
0-
02
b1 6
#402110000000
1!
1%
1-
12
#402120000000
0!
0%
b10 *
0-
02
b10 6
#402130000000
1!
1%
1-
12
#402140000000
0!
0%
b11 *
0-
02
b11 6
#402150000000
1!
1%
1-
12
15
#402160000000
0!
0%
b100 *
0-
02
b100 6
#402170000000
1!
1%
1-
12
#402180000000
0!
0%
b101 *
0-
02
b101 6
#402190000000
1!
1%
1-
12
#402200000000
0!
0%
b110 *
0-
02
b110 6
#402210000000
1!
1%
1-
12
#402220000000
0!
0%
b111 *
0-
02
b111 6
#402230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#402240000000
0!
0%
b0 *
0-
02
b0 6
#402250000000
1!
1%
1-
12
#402260000000
0!
0%
b1 *
0-
02
b1 6
#402270000000
1!
1%
1-
12
#402280000000
0!
0%
b10 *
0-
02
b10 6
#402290000000
1!
1%
1-
12
#402300000000
0!
0%
b11 *
0-
02
b11 6
#402310000000
1!
1%
1-
12
15
#402320000000
0!
0%
b100 *
0-
02
b100 6
#402330000000
1!
1%
1-
12
#402340000000
0!
0%
b101 *
0-
02
b101 6
#402350000000
1!
1%
1-
12
#402360000000
0!
0%
b110 *
0-
02
b110 6
#402370000000
1!
1%
1-
12
#402380000000
0!
0%
b111 *
0-
02
b111 6
#402390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#402400000000
0!
0%
b0 *
0-
02
b0 6
#402410000000
1!
1%
1-
12
#402420000000
0!
0%
b1 *
0-
02
b1 6
#402430000000
1!
1%
1-
12
#402440000000
0!
0%
b10 *
0-
02
b10 6
#402450000000
1!
1%
1-
12
#402460000000
0!
0%
b11 *
0-
02
b11 6
#402470000000
1!
1%
1-
12
15
#402480000000
0!
0%
b100 *
0-
02
b100 6
#402490000000
1!
1%
1-
12
#402500000000
0!
0%
b101 *
0-
02
b101 6
#402510000000
1!
1%
1-
12
#402520000000
0!
0%
b110 *
0-
02
b110 6
#402530000000
1!
1%
1-
12
#402540000000
0!
0%
b111 *
0-
02
b111 6
#402550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#402560000000
0!
0%
b0 *
0-
02
b0 6
#402570000000
1!
1%
1-
12
#402580000000
0!
0%
b1 *
0-
02
b1 6
#402590000000
1!
1%
1-
12
#402600000000
0!
0%
b10 *
0-
02
b10 6
#402610000000
1!
1%
1-
12
#402620000000
0!
0%
b11 *
0-
02
b11 6
#402630000000
1!
1%
1-
12
15
#402640000000
0!
0%
b100 *
0-
02
b100 6
#402650000000
1!
1%
1-
12
#402660000000
0!
0%
b101 *
0-
02
b101 6
#402670000000
1!
1%
1-
12
#402680000000
0!
0%
b110 *
0-
02
b110 6
#402690000000
1!
1%
1-
12
#402700000000
0!
0%
b111 *
0-
02
b111 6
#402710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#402720000000
0!
0%
b0 *
0-
02
b0 6
#402730000000
1!
1%
1-
12
#402740000000
0!
0%
b1 *
0-
02
b1 6
#402750000000
1!
1%
1-
12
#402760000000
0!
0%
b10 *
0-
02
b10 6
#402770000000
1!
1%
1-
12
#402780000000
0!
0%
b11 *
0-
02
b11 6
#402790000000
1!
1%
1-
12
15
#402800000000
0!
0%
b100 *
0-
02
b100 6
#402810000000
1!
1%
1-
12
#402820000000
0!
0%
b101 *
0-
02
b101 6
#402830000000
1!
1%
1-
12
#402840000000
0!
0%
b110 *
0-
02
b110 6
#402850000000
1!
1%
1-
12
#402860000000
0!
0%
b111 *
0-
02
b111 6
#402870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#402880000000
0!
0%
b0 *
0-
02
b0 6
#402890000000
1!
1%
1-
12
#402900000000
0!
0%
b1 *
0-
02
b1 6
#402910000000
1!
1%
1-
12
#402920000000
0!
0%
b10 *
0-
02
b10 6
#402930000000
1!
1%
1-
12
#402940000000
0!
0%
b11 *
0-
02
b11 6
#402950000000
1!
1%
1-
12
15
#402960000000
0!
0%
b100 *
0-
02
b100 6
#402970000000
1!
1%
1-
12
#402980000000
0!
0%
b101 *
0-
02
b101 6
#402990000000
1!
1%
1-
12
#403000000000
0!
0%
b110 *
0-
02
b110 6
#403010000000
1!
1%
1-
12
#403020000000
0!
0%
b111 *
0-
02
b111 6
#403030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#403040000000
0!
0%
b0 *
0-
02
b0 6
#403050000000
1!
1%
1-
12
#403060000000
0!
0%
b1 *
0-
02
b1 6
#403070000000
1!
1%
1-
12
#403080000000
0!
0%
b10 *
0-
02
b10 6
#403090000000
1!
1%
1-
12
#403100000000
0!
0%
b11 *
0-
02
b11 6
#403110000000
1!
1%
1-
12
15
#403120000000
0!
0%
b100 *
0-
02
b100 6
#403130000000
1!
1%
1-
12
#403140000000
0!
0%
b101 *
0-
02
b101 6
#403150000000
1!
1%
1-
12
#403160000000
0!
0%
b110 *
0-
02
b110 6
#403170000000
1!
1%
1-
12
#403180000000
0!
0%
b111 *
0-
02
b111 6
#403190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#403200000000
0!
0%
b0 *
0-
02
b0 6
#403210000000
1!
1%
1-
12
#403220000000
0!
0%
b1 *
0-
02
b1 6
#403230000000
1!
1%
1-
12
#403240000000
0!
0%
b10 *
0-
02
b10 6
#403250000000
1!
1%
1-
12
#403260000000
0!
0%
b11 *
0-
02
b11 6
#403270000000
1!
1%
1-
12
15
#403280000000
0!
0%
b100 *
0-
02
b100 6
#403290000000
1!
1%
1-
12
#403300000000
0!
0%
b101 *
0-
02
b101 6
#403310000000
1!
1%
1-
12
#403320000000
0!
0%
b110 *
0-
02
b110 6
#403330000000
1!
1%
1-
12
#403340000000
0!
0%
b111 *
0-
02
b111 6
#403350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#403360000000
0!
0%
b0 *
0-
02
b0 6
#403370000000
1!
1%
1-
12
#403380000000
0!
0%
b1 *
0-
02
b1 6
#403390000000
1!
1%
1-
12
#403400000000
0!
0%
b10 *
0-
02
b10 6
#403410000000
1!
1%
1-
12
#403420000000
0!
0%
b11 *
0-
02
b11 6
#403430000000
1!
1%
1-
12
15
#403440000000
0!
0%
b100 *
0-
02
b100 6
#403450000000
1!
1%
1-
12
#403460000000
0!
0%
b101 *
0-
02
b101 6
#403470000000
1!
1%
1-
12
#403480000000
0!
0%
b110 *
0-
02
b110 6
#403490000000
1!
1%
1-
12
#403500000000
0!
0%
b111 *
0-
02
b111 6
#403510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#403520000000
0!
0%
b0 *
0-
02
b0 6
#403530000000
1!
1%
1-
12
#403540000000
0!
0%
b1 *
0-
02
b1 6
#403550000000
1!
1%
1-
12
#403560000000
0!
0%
b10 *
0-
02
b10 6
#403570000000
1!
1%
1-
12
#403580000000
0!
0%
b11 *
0-
02
b11 6
#403590000000
1!
1%
1-
12
15
#403600000000
0!
0%
b100 *
0-
02
b100 6
#403610000000
1!
1%
1-
12
#403620000000
0!
0%
b101 *
0-
02
b101 6
#403630000000
1!
1%
1-
12
#403640000000
0!
0%
b110 *
0-
02
b110 6
#403650000000
1!
1%
1-
12
#403660000000
0!
0%
b111 *
0-
02
b111 6
#403670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#403680000000
0!
0%
b0 *
0-
02
b0 6
#403690000000
1!
1%
1-
12
#403700000000
0!
0%
b1 *
0-
02
b1 6
#403710000000
1!
1%
1-
12
#403720000000
0!
0%
b10 *
0-
02
b10 6
#403730000000
1!
1%
1-
12
#403740000000
0!
0%
b11 *
0-
02
b11 6
#403750000000
1!
1%
1-
12
15
#403760000000
0!
0%
b100 *
0-
02
b100 6
#403770000000
1!
1%
1-
12
#403780000000
0!
0%
b101 *
0-
02
b101 6
#403790000000
1!
1%
1-
12
#403800000000
0!
0%
b110 *
0-
02
b110 6
#403810000000
1!
1%
1-
12
#403820000000
0!
0%
b111 *
0-
02
b111 6
#403830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#403840000000
0!
0%
b0 *
0-
02
b0 6
#403850000000
1!
1%
1-
12
#403860000000
0!
0%
b1 *
0-
02
b1 6
#403870000000
1!
1%
1-
12
#403880000000
0!
0%
b10 *
0-
02
b10 6
#403890000000
1!
1%
1-
12
#403900000000
0!
0%
b11 *
0-
02
b11 6
#403910000000
1!
1%
1-
12
15
#403920000000
0!
0%
b100 *
0-
02
b100 6
#403930000000
1!
1%
1-
12
#403940000000
0!
0%
b101 *
0-
02
b101 6
#403950000000
1!
1%
1-
12
#403960000000
0!
0%
b110 *
0-
02
b110 6
#403970000000
1!
1%
1-
12
#403980000000
0!
0%
b111 *
0-
02
b111 6
#403990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#404000000000
0!
0%
b0 *
0-
02
b0 6
#404010000000
1!
1%
1-
12
#404020000000
0!
0%
b1 *
0-
02
b1 6
#404030000000
1!
1%
1-
12
#404040000000
0!
0%
b10 *
0-
02
b10 6
#404050000000
1!
1%
1-
12
#404060000000
0!
0%
b11 *
0-
02
b11 6
#404070000000
1!
1%
1-
12
15
#404080000000
0!
0%
b100 *
0-
02
b100 6
#404090000000
1!
1%
1-
12
#404100000000
0!
0%
b101 *
0-
02
b101 6
#404110000000
1!
1%
1-
12
#404120000000
0!
0%
b110 *
0-
02
b110 6
#404130000000
1!
1%
1-
12
#404140000000
0!
0%
b111 *
0-
02
b111 6
#404150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#404160000000
0!
0%
b0 *
0-
02
b0 6
#404170000000
1!
1%
1-
12
#404180000000
0!
0%
b1 *
0-
02
b1 6
#404190000000
1!
1%
1-
12
#404200000000
0!
0%
b10 *
0-
02
b10 6
#404210000000
1!
1%
1-
12
#404220000000
0!
0%
b11 *
0-
02
b11 6
#404230000000
1!
1%
1-
12
15
#404240000000
0!
0%
b100 *
0-
02
b100 6
#404250000000
1!
1%
1-
12
#404260000000
0!
0%
b101 *
0-
02
b101 6
#404270000000
1!
1%
1-
12
#404280000000
0!
0%
b110 *
0-
02
b110 6
#404290000000
1!
1%
1-
12
#404300000000
0!
0%
b111 *
0-
02
b111 6
#404310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#404320000000
0!
0%
b0 *
0-
02
b0 6
#404330000000
1!
1%
1-
12
#404340000000
0!
0%
b1 *
0-
02
b1 6
#404350000000
1!
1%
1-
12
#404360000000
0!
0%
b10 *
0-
02
b10 6
#404370000000
1!
1%
1-
12
#404380000000
0!
0%
b11 *
0-
02
b11 6
#404390000000
1!
1%
1-
12
15
#404400000000
0!
0%
b100 *
0-
02
b100 6
#404410000000
1!
1%
1-
12
#404420000000
0!
0%
b101 *
0-
02
b101 6
#404430000000
1!
1%
1-
12
#404440000000
0!
0%
b110 *
0-
02
b110 6
#404450000000
1!
1%
1-
12
#404460000000
0!
0%
b111 *
0-
02
b111 6
#404470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#404480000000
0!
0%
b0 *
0-
02
b0 6
#404490000000
1!
1%
1-
12
#404500000000
0!
0%
b1 *
0-
02
b1 6
#404510000000
1!
1%
1-
12
#404520000000
0!
0%
b10 *
0-
02
b10 6
#404530000000
1!
1%
1-
12
#404540000000
0!
0%
b11 *
0-
02
b11 6
#404550000000
1!
1%
1-
12
15
#404560000000
0!
0%
b100 *
0-
02
b100 6
#404570000000
1!
1%
1-
12
#404580000000
0!
0%
b101 *
0-
02
b101 6
#404590000000
1!
1%
1-
12
#404600000000
0!
0%
b110 *
0-
02
b110 6
#404610000000
1!
1%
1-
12
#404620000000
0!
0%
b111 *
0-
02
b111 6
#404630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#404640000000
0!
0%
b0 *
0-
02
b0 6
#404650000000
1!
1%
1-
12
#404660000000
0!
0%
b1 *
0-
02
b1 6
#404670000000
1!
1%
1-
12
#404680000000
0!
0%
b10 *
0-
02
b10 6
#404690000000
1!
1%
1-
12
#404700000000
0!
0%
b11 *
0-
02
b11 6
#404710000000
1!
1%
1-
12
15
#404720000000
0!
0%
b100 *
0-
02
b100 6
#404730000000
1!
1%
1-
12
#404740000000
0!
0%
b101 *
0-
02
b101 6
#404750000000
1!
1%
1-
12
#404760000000
0!
0%
b110 *
0-
02
b110 6
#404770000000
1!
1%
1-
12
#404780000000
0!
0%
b111 *
0-
02
b111 6
#404790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#404800000000
0!
0%
b0 *
0-
02
b0 6
#404810000000
1!
1%
1-
12
#404820000000
0!
0%
b1 *
0-
02
b1 6
#404830000000
1!
1%
1-
12
#404840000000
0!
0%
b10 *
0-
02
b10 6
#404850000000
1!
1%
1-
12
#404860000000
0!
0%
b11 *
0-
02
b11 6
#404870000000
1!
1%
1-
12
15
#404880000000
0!
0%
b100 *
0-
02
b100 6
#404890000000
1!
1%
1-
12
#404900000000
0!
0%
b101 *
0-
02
b101 6
#404910000000
1!
1%
1-
12
#404920000000
0!
0%
b110 *
0-
02
b110 6
#404930000000
1!
1%
1-
12
#404940000000
0!
0%
b111 *
0-
02
b111 6
#404950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#404960000000
0!
0%
b0 *
0-
02
b0 6
#404970000000
1!
1%
1-
12
#404980000000
0!
0%
b1 *
0-
02
b1 6
#404990000000
1!
1%
1-
12
#405000000000
0!
0%
b10 *
0-
02
b10 6
#405010000000
1!
1%
1-
12
#405020000000
0!
0%
b11 *
0-
02
b11 6
#405030000000
1!
1%
1-
12
15
#405040000000
0!
0%
b100 *
0-
02
b100 6
#405050000000
1!
1%
1-
12
#405060000000
0!
0%
b101 *
0-
02
b101 6
#405070000000
1!
1%
1-
12
#405080000000
0!
0%
b110 *
0-
02
b110 6
#405090000000
1!
1%
1-
12
#405100000000
0!
0%
b111 *
0-
02
b111 6
#405110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#405120000000
0!
0%
b0 *
0-
02
b0 6
#405130000000
1!
1%
1-
12
#405140000000
0!
0%
b1 *
0-
02
b1 6
#405150000000
1!
1%
1-
12
#405160000000
0!
0%
b10 *
0-
02
b10 6
#405170000000
1!
1%
1-
12
#405180000000
0!
0%
b11 *
0-
02
b11 6
#405190000000
1!
1%
1-
12
15
#405200000000
0!
0%
b100 *
0-
02
b100 6
#405210000000
1!
1%
1-
12
#405220000000
0!
0%
b101 *
0-
02
b101 6
#405230000000
1!
1%
1-
12
#405240000000
0!
0%
b110 *
0-
02
b110 6
#405250000000
1!
1%
1-
12
#405260000000
0!
0%
b111 *
0-
02
b111 6
#405270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#405280000000
0!
0%
b0 *
0-
02
b0 6
#405290000000
1!
1%
1-
12
#405300000000
0!
0%
b1 *
0-
02
b1 6
#405310000000
1!
1%
1-
12
#405320000000
0!
0%
b10 *
0-
02
b10 6
#405330000000
1!
1%
1-
12
#405340000000
0!
0%
b11 *
0-
02
b11 6
#405350000000
1!
1%
1-
12
15
#405360000000
0!
0%
b100 *
0-
02
b100 6
#405370000000
1!
1%
1-
12
#405380000000
0!
0%
b101 *
0-
02
b101 6
#405390000000
1!
1%
1-
12
#405400000000
0!
0%
b110 *
0-
02
b110 6
#405410000000
1!
1%
1-
12
#405420000000
0!
0%
b111 *
0-
02
b111 6
#405430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#405440000000
0!
0%
b0 *
0-
02
b0 6
#405450000000
1!
1%
1-
12
#405460000000
0!
0%
b1 *
0-
02
b1 6
#405470000000
1!
1%
1-
12
#405480000000
0!
0%
b10 *
0-
02
b10 6
#405490000000
1!
1%
1-
12
#405500000000
0!
0%
b11 *
0-
02
b11 6
#405510000000
1!
1%
1-
12
15
#405520000000
0!
0%
b100 *
0-
02
b100 6
#405530000000
1!
1%
1-
12
#405540000000
0!
0%
b101 *
0-
02
b101 6
#405550000000
1!
1%
1-
12
#405560000000
0!
0%
b110 *
0-
02
b110 6
#405570000000
1!
1%
1-
12
#405580000000
0!
0%
b111 *
0-
02
b111 6
#405590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#405600000000
0!
0%
b0 *
0-
02
b0 6
#405610000000
1!
1%
1-
12
#405620000000
0!
0%
b1 *
0-
02
b1 6
#405630000000
1!
1%
1-
12
#405640000000
0!
0%
b10 *
0-
02
b10 6
#405650000000
1!
1%
1-
12
#405660000000
0!
0%
b11 *
0-
02
b11 6
#405670000000
1!
1%
1-
12
15
#405680000000
0!
0%
b100 *
0-
02
b100 6
#405690000000
1!
1%
1-
12
#405700000000
0!
0%
b101 *
0-
02
b101 6
#405710000000
1!
1%
1-
12
#405720000000
0!
0%
b110 *
0-
02
b110 6
#405730000000
1!
1%
1-
12
#405740000000
0!
0%
b111 *
0-
02
b111 6
#405750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#405760000000
0!
0%
b0 *
0-
02
b0 6
#405770000000
1!
1%
1-
12
#405780000000
0!
0%
b1 *
0-
02
b1 6
#405790000000
1!
1%
1-
12
#405800000000
0!
0%
b10 *
0-
02
b10 6
#405810000000
1!
1%
1-
12
#405820000000
0!
0%
b11 *
0-
02
b11 6
#405830000000
1!
1%
1-
12
15
#405840000000
0!
0%
b100 *
0-
02
b100 6
#405850000000
1!
1%
1-
12
#405860000000
0!
0%
b101 *
0-
02
b101 6
#405870000000
1!
1%
1-
12
#405880000000
0!
0%
b110 *
0-
02
b110 6
#405890000000
1!
1%
1-
12
#405900000000
0!
0%
b111 *
0-
02
b111 6
#405910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#405920000000
0!
0%
b0 *
0-
02
b0 6
#405930000000
1!
1%
1-
12
#405940000000
0!
0%
b1 *
0-
02
b1 6
#405950000000
1!
1%
1-
12
#405960000000
0!
0%
b10 *
0-
02
b10 6
#405970000000
1!
1%
1-
12
#405980000000
0!
0%
b11 *
0-
02
b11 6
#405990000000
1!
1%
1-
12
15
#406000000000
0!
0%
b100 *
0-
02
b100 6
#406010000000
1!
1%
1-
12
#406020000000
0!
0%
b101 *
0-
02
b101 6
#406030000000
1!
1%
1-
12
#406040000000
0!
0%
b110 *
0-
02
b110 6
#406050000000
1!
1%
1-
12
#406060000000
0!
0%
b111 *
0-
02
b111 6
#406070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#406080000000
0!
0%
b0 *
0-
02
b0 6
#406090000000
1!
1%
1-
12
#406100000000
0!
0%
b1 *
0-
02
b1 6
#406110000000
1!
1%
1-
12
#406120000000
0!
0%
b10 *
0-
02
b10 6
#406130000000
1!
1%
1-
12
#406140000000
0!
0%
b11 *
0-
02
b11 6
#406150000000
1!
1%
1-
12
15
#406160000000
0!
0%
b100 *
0-
02
b100 6
#406170000000
1!
1%
1-
12
#406180000000
0!
0%
b101 *
0-
02
b101 6
#406190000000
1!
1%
1-
12
#406200000000
0!
0%
b110 *
0-
02
b110 6
#406210000000
1!
1%
1-
12
#406220000000
0!
0%
b111 *
0-
02
b111 6
#406230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#406240000000
0!
0%
b0 *
0-
02
b0 6
#406250000000
1!
1%
1-
12
#406260000000
0!
0%
b1 *
0-
02
b1 6
#406270000000
1!
1%
1-
12
#406280000000
0!
0%
b10 *
0-
02
b10 6
#406290000000
1!
1%
1-
12
#406300000000
0!
0%
b11 *
0-
02
b11 6
#406310000000
1!
1%
1-
12
15
#406320000000
0!
0%
b100 *
0-
02
b100 6
#406330000000
1!
1%
1-
12
#406340000000
0!
0%
b101 *
0-
02
b101 6
#406350000000
1!
1%
1-
12
#406360000000
0!
0%
b110 *
0-
02
b110 6
#406370000000
1!
1%
1-
12
#406380000000
0!
0%
b111 *
0-
02
b111 6
#406390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#406400000000
0!
0%
b0 *
0-
02
b0 6
#406410000000
1!
1%
1-
12
#406420000000
0!
0%
b1 *
0-
02
b1 6
#406430000000
1!
1%
1-
12
#406440000000
0!
0%
b10 *
0-
02
b10 6
#406450000000
1!
1%
1-
12
#406460000000
0!
0%
b11 *
0-
02
b11 6
#406470000000
1!
1%
1-
12
15
#406480000000
0!
0%
b100 *
0-
02
b100 6
#406490000000
1!
1%
1-
12
#406500000000
0!
0%
b101 *
0-
02
b101 6
#406510000000
1!
1%
1-
12
#406520000000
0!
0%
b110 *
0-
02
b110 6
#406530000000
1!
1%
1-
12
#406540000000
0!
0%
b111 *
0-
02
b111 6
#406550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#406560000000
0!
0%
b0 *
0-
02
b0 6
#406570000000
1!
1%
1-
12
#406580000000
0!
0%
b1 *
0-
02
b1 6
#406590000000
1!
1%
1-
12
#406600000000
0!
0%
b10 *
0-
02
b10 6
#406610000000
1!
1%
1-
12
#406620000000
0!
0%
b11 *
0-
02
b11 6
#406630000000
1!
1%
1-
12
15
#406640000000
0!
0%
b100 *
0-
02
b100 6
#406650000000
1!
1%
1-
12
#406660000000
0!
0%
b101 *
0-
02
b101 6
#406670000000
1!
1%
1-
12
#406680000000
0!
0%
b110 *
0-
02
b110 6
#406690000000
1!
1%
1-
12
#406700000000
0!
0%
b111 *
0-
02
b111 6
#406710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#406720000000
0!
0%
b0 *
0-
02
b0 6
#406730000000
1!
1%
1-
12
#406740000000
0!
0%
b1 *
0-
02
b1 6
#406750000000
1!
1%
1-
12
#406760000000
0!
0%
b10 *
0-
02
b10 6
#406770000000
1!
1%
1-
12
#406780000000
0!
0%
b11 *
0-
02
b11 6
#406790000000
1!
1%
1-
12
15
#406800000000
0!
0%
b100 *
0-
02
b100 6
#406810000000
1!
1%
1-
12
#406820000000
0!
0%
b101 *
0-
02
b101 6
#406830000000
1!
1%
1-
12
#406840000000
0!
0%
b110 *
0-
02
b110 6
#406850000000
1!
1%
1-
12
#406860000000
0!
0%
b111 *
0-
02
b111 6
#406870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#406880000000
0!
0%
b0 *
0-
02
b0 6
#406890000000
1!
1%
1-
12
#406900000000
0!
0%
b1 *
0-
02
b1 6
#406910000000
1!
1%
1-
12
#406920000000
0!
0%
b10 *
0-
02
b10 6
#406930000000
1!
1%
1-
12
#406940000000
0!
0%
b11 *
0-
02
b11 6
#406950000000
1!
1%
1-
12
15
#406960000000
0!
0%
b100 *
0-
02
b100 6
#406970000000
1!
1%
1-
12
#406980000000
0!
0%
b101 *
0-
02
b101 6
#406990000000
1!
1%
1-
12
#407000000000
0!
0%
b110 *
0-
02
b110 6
#407010000000
1!
1%
1-
12
#407020000000
0!
0%
b111 *
0-
02
b111 6
#407030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#407040000000
0!
0%
b0 *
0-
02
b0 6
#407050000000
1!
1%
1-
12
#407060000000
0!
0%
b1 *
0-
02
b1 6
#407070000000
1!
1%
1-
12
#407080000000
0!
0%
b10 *
0-
02
b10 6
#407090000000
1!
1%
1-
12
#407100000000
0!
0%
b11 *
0-
02
b11 6
#407110000000
1!
1%
1-
12
15
#407120000000
0!
0%
b100 *
0-
02
b100 6
#407130000000
1!
1%
1-
12
#407140000000
0!
0%
b101 *
0-
02
b101 6
#407150000000
1!
1%
1-
12
#407160000000
0!
0%
b110 *
0-
02
b110 6
#407170000000
1!
1%
1-
12
#407180000000
0!
0%
b111 *
0-
02
b111 6
#407190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#407200000000
0!
0%
b0 *
0-
02
b0 6
#407210000000
1!
1%
1-
12
#407220000000
0!
0%
b1 *
0-
02
b1 6
#407230000000
1!
1%
1-
12
#407240000000
0!
0%
b10 *
0-
02
b10 6
#407250000000
1!
1%
1-
12
#407260000000
0!
0%
b11 *
0-
02
b11 6
#407270000000
1!
1%
1-
12
15
#407280000000
0!
0%
b100 *
0-
02
b100 6
#407290000000
1!
1%
1-
12
#407300000000
0!
0%
b101 *
0-
02
b101 6
#407310000000
1!
1%
1-
12
#407320000000
0!
0%
b110 *
0-
02
b110 6
#407330000000
1!
1%
1-
12
#407340000000
0!
0%
b111 *
0-
02
b111 6
#407350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#407360000000
0!
0%
b0 *
0-
02
b0 6
#407370000000
1!
1%
1-
12
#407380000000
0!
0%
b1 *
0-
02
b1 6
#407390000000
1!
1%
1-
12
#407400000000
0!
0%
b10 *
0-
02
b10 6
#407410000000
1!
1%
1-
12
#407420000000
0!
0%
b11 *
0-
02
b11 6
#407430000000
1!
1%
1-
12
15
#407440000000
0!
0%
b100 *
0-
02
b100 6
#407450000000
1!
1%
1-
12
#407460000000
0!
0%
b101 *
0-
02
b101 6
#407470000000
1!
1%
1-
12
#407480000000
0!
0%
b110 *
0-
02
b110 6
#407490000000
1!
1%
1-
12
#407500000000
0!
0%
b111 *
0-
02
b111 6
#407510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#407520000000
0!
0%
b0 *
0-
02
b0 6
#407530000000
1!
1%
1-
12
#407540000000
0!
0%
b1 *
0-
02
b1 6
#407550000000
1!
1%
1-
12
#407560000000
0!
0%
b10 *
0-
02
b10 6
#407570000000
1!
1%
1-
12
#407580000000
0!
0%
b11 *
0-
02
b11 6
#407590000000
1!
1%
1-
12
15
#407600000000
0!
0%
b100 *
0-
02
b100 6
#407610000000
1!
1%
1-
12
#407620000000
0!
0%
b101 *
0-
02
b101 6
#407630000000
1!
1%
1-
12
#407640000000
0!
0%
b110 *
0-
02
b110 6
#407650000000
1!
1%
1-
12
#407660000000
0!
0%
b111 *
0-
02
b111 6
#407670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#407680000000
0!
0%
b0 *
0-
02
b0 6
#407690000000
1!
1%
1-
12
#407700000000
0!
0%
b1 *
0-
02
b1 6
#407710000000
1!
1%
1-
12
#407720000000
0!
0%
b10 *
0-
02
b10 6
#407730000000
1!
1%
1-
12
#407740000000
0!
0%
b11 *
0-
02
b11 6
#407750000000
1!
1%
1-
12
15
#407760000000
0!
0%
b100 *
0-
02
b100 6
#407770000000
1!
1%
1-
12
#407780000000
0!
0%
b101 *
0-
02
b101 6
#407790000000
1!
1%
1-
12
#407800000000
0!
0%
b110 *
0-
02
b110 6
#407810000000
1!
1%
1-
12
#407820000000
0!
0%
b111 *
0-
02
b111 6
#407830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#407840000000
0!
0%
b0 *
0-
02
b0 6
#407850000000
1!
1%
1-
12
#407860000000
0!
0%
b1 *
0-
02
b1 6
#407870000000
1!
1%
1-
12
#407880000000
0!
0%
b10 *
0-
02
b10 6
#407890000000
1!
1%
1-
12
#407900000000
0!
0%
b11 *
0-
02
b11 6
#407910000000
1!
1%
1-
12
15
#407920000000
0!
0%
b100 *
0-
02
b100 6
#407930000000
1!
1%
1-
12
#407940000000
0!
0%
b101 *
0-
02
b101 6
#407950000000
1!
1%
1-
12
#407960000000
0!
0%
b110 *
0-
02
b110 6
#407970000000
1!
1%
1-
12
#407980000000
0!
0%
b111 *
0-
02
b111 6
#407990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#408000000000
0!
0%
b0 *
0-
02
b0 6
#408010000000
1!
1%
1-
12
#408020000000
0!
0%
b1 *
0-
02
b1 6
#408030000000
1!
1%
1-
12
#408040000000
0!
0%
b10 *
0-
02
b10 6
#408050000000
1!
1%
1-
12
#408060000000
0!
0%
b11 *
0-
02
b11 6
#408070000000
1!
1%
1-
12
15
#408080000000
0!
0%
b100 *
0-
02
b100 6
#408090000000
1!
1%
1-
12
#408100000000
0!
0%
b101 *
0-
02
b101 6
#408110000000
1!
1%
1-
12
#408120000000
0!
0%
b110 *
0-
02
b110 6
#408130000000
1!
1%
1-
12
#408140000000
0!
0%
b111 *
0-
02
b111 6
#408150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#408160000000
0!
0%
b0 *
0-
02
b0 6
#408170000000
1!
1%
1-
12
#408180000000
0!
0%
b1 *
0-
02
b1 6
#408190000000
1!
1%
1-
12
#408200000000
0!
0%
b10 *
0-
02
b10 6
#408210000000
1!
1%
1-
12
#408220000000
0!
0%
b11 *
0-
02
b11 6
#408230000000
1!
1%
1-
12
15
#408240000000
0!
0%
b100 *
0-
02
b100 6
#408250000000
1!
1%
1-
12
#408260000000
0!
0%
b101 *
0-
02
b101 6
#408270000000
1!
1%
1-
12
#408280000000
0!
0%
b110 *
0-
02
b110 6
#408290000000
1!
1%
1-
12
#408300000000
0!
0%
b111 *
0-
02
b111 6
#408310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#408320000000
0!
0%
b0 *
0-
02
b0 6
#408330000000
1!
1%
1-
12
#408340000000
0!
0%
b1 *
0-
02
b1 6
#408350000000
1!
1%
1-
12
#408360000000
0!
0%
b10 *
0-
02
b10 6
#408370000000
1!
1%
1-
12
#408380000000
0!
0%
b11 *
0-
02
b11 6
#408390000000
1!
1%
1-
12
15
#408400000000
0!
0%
b100 *
0-
02
b100 6
#408410000000
1!
1%
1-
12
#408420000000
0!
0%
b101 *
0-
02
b101 6
#408430000000
1!
1%
1-
12
#408440000000
0!
0%
b110 *
0-
02
b110 6
#408450000000
1!
1%
1-
12
#408460000000
0!
0%
b111 *
0-
02
b111 6
#408470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#408480000000
0!
0%
b0 *
0-
02
b0 6
#408490000000
1!
1%
1-
12
#408500000000
0!
0%
b1 *
0-
02
b1 6
#408510000000
1!
1%
1-
12
#408520000000
0!
0%
b10 *
0-
02
b10 6
#408530000000
1!
1%
1-
12
#408540000000
0!
0%
b11 *
0-
02
b11 6
#408550000000
1!
1%
1-
12
15
#408560000000
0!
0%
b100 *
0-
02
b100 6
#408570000000
1!
1%
1-
12
#408580000000
0!
0%
b101 *
0-
02
b101 6
#408590000000
1!
1%
1-
12
#408600000000
0!
0%
b110 *
0-
02
b110 6
#408610000000
1!
1%
1-
12
#408620000000
0!
0%
b111 *
0-
02
b111 6
#408630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#408640000000
0!
0%
b0 *
0-
02
b0 6
#408650000000
1!
1%
1-
12
#408660000000
0!
0%
b1 *
0-
02
b1 6
#408670000000
1!
1%
1-
12
#408680000000
0!
0%
b10 *
0-
02
b10 6
#408690000000
1!
1%
1-
12
#408700000000
0!
0%
b11 *
0-
02
b11 6
#408710000000
1!
1%
1-
12
15
#408720000000
0!
0%
b100 *
0-
02
b100 6
#408730000000
1!
1%
1-
12
#408740000000
0!
0%
b101 *
0-
02
b101 6
#408750000000
1!
1%
1-
12
#408760000000
0!
0%
b110 *
0-
02
b110 6
#408770000000
1!
1%
1-
12
#408780000000
0!
0%
b111 *
0-
02
b111 6
#408790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#408800000000
0!
0%
b0 *
0-
02
b0 6
#408810000000
1!
1%
1-
12
#408820000000
0!
0%
b1 *
0-
02
b1 6
#408830000000
1!
1%
1-
12
#408840000000
0!
0%
b10 *
0-
02
b10 6
#408850000000
1!
1%
1-
12
#408860000000
0!
0%
b11 *
0-
02
b11 6
#408870000000
1!
1%
1-
12
15
#408880000000
0!
0%
b100 *
0-
02
b100 6
#408890000000
1!
1%
1-
12
#408900000000
0!
0%
b101 *
0-
02
b101 6
#408910000000
1!
1%
1-
12
#408920000000
0!
0%
b110 *
0-
02
b110 6
#408930000000
1!
1%
1-
12
#408940000000
0!
0%
b111 *
0-
02
b111 6
#408950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#408960000000
0!
0%
b0 *
0-
02
b0 6
#408970000000
1!
1%
1-
12
#408980000000
0!
0%
b1 *
0-
02
b1 6
#408990000000
1!
1%
1-
12
#409000000000
0!
0%
b10 *
0-
02
b10 6
#409010000000
1!
1%
1-
12
#409020000000
0!
0%
b11 *
0-
02
b11 6
#409030000000
1!
1%
1-
12
15
#409040000000
0!
0%
b100 *
0-
02
b100 6
#409050000000
1!
1%
1-
12
#409060000000
0!
0%
b101 *
0-
02
b101 6
#409070000000
1!
1%
1-
12
#409080000000
0!
0%
b110 *
0-
02
b110 6
#409090000000
1!
1%
1-
12
#409100000000
0!
0%
b111 *
0-
02
b111 6
#409110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#409120000000
0!
0%
b0 *
0-
02
b0 6
#409130000000
1!
1%
1-
12
#409140000000
0!
0%
b1 *
0-
02
b1 6
#409150000000
1!
1%
1-
12
#409160000000
0!
0%
b10 *
0-
02
b10 6
#409170000000
1!
1%
1-
12
#409180000000
0!
0%
b11 *
0-
02
b11 6
#409190000000
1!
1%
1-
12
15
#409200000000
0!
0%
b100 *
0-
02
b100 6
#409210000000
1!
1%
1-
12
#409220000000
0!
0%
b101 *
0-
02
b101 6
#409230000000
1!
1%
1-
12
#409240000000
0!
0%
b110 *
0-
02
b110 6
#409250000000
1!
1%
1-
12
#409260000000
0!
0%
b111 *
0-
02
b111 6
#409270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#409280000000
0!
0%
b0 *
0-
02
b0 6
#409290000000
1!
1%
1-
12
#409300000000
0!
0%
b1 *
0-
02
b1 6
#409310000000
1!
1%
1-
12
#409320000000
0!
0%
b10 *
0-
02
b10 6
#409330000000
1!
1%
1-
12
#409340000000
0!
0%
b11 *
0-
02
b11 6
#409350000000
1!
1%
1-
12
15
#409360000000
0!
0%
b100 *
0-
02
b100 6
#409370000000
1!
1%
1-
12
#409380000000
0!
0%
b101 *
0-
02
b101 6
#409390000000
1!
1%
1-
12
#409400000000
0!
0%
b110 *
0-
02
b110 6
#409410000000
1!
1%
1-
12
#409420000000
0!
0%
b111 *
0-
02
b111 6
#409430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#409440000000
0!
0%
b0 *
0-
02
b0 6
#409450000000
1!
1%
1-
12
#409460000000
0!
0%
b1 *
0-
02
b1 6
#409470000000
1!
1%
1-
12
#409480000000
0!
0%
b10 *
0-
02
b10 6
#409490000000
1!
1%
1-
12
#409500000000
0!
0%
b11 *
0-
02
b11 6
#409510000000
1!
1%
1-
12
15
#409520000000
0!
0%
b100 *
0-
02
b100 6
#409530000000
1!
1%
1-
12
#409540000000
0!
0%
b101 *
0-
02
b101 6
#409550000000
1!
1%
1-
12
#409560000000
0!
0%
b110 *
0-
02
b110 6
#409570000000
1!
1%
1-
12
#409580000000
0!
0%
b111 *
0-
02
b111 6
#409590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#409600000000
0!
0%
b0 *
0-
02
b0 6
#409610000000
1!
1%
1-
12
#409620000000
0!
0%
b1 *
0-
02
b1 6
#409630000000
1!
1%
1-
12
#409640000000
0!
0%
b10 *
0-
02
b10 6
#409650000000
1!
1%
1-
12
#409660000000
0!
0%
b11 *
0-
02
b11 6
#409670000000
1!
1%
1-
12
15
#409680000000
0!
0%
b100 *
0-
02
b100 6
#409690000000
1!
1%
1-
12
#409700000000
0!
0%
b101 *
0-
02
b101 6
#409710000000
1!
1%
1-
12
#409720000000
0!
0%
b110 *
0-
02
b110 6
#409730000000
1!
1%
1-
12
#409740000000
0!
0%
b111 *
0-
02
b111 6
#409750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#409760000000
0!
0%
b0 *
0-
02
b0 6
#409770000000
1!
1%
1-
12
#409780000000
0!
0%
b1 *
0-
02
b1 6
#409790000000
1!
1%
1-
12
#409800000000
0!
0%
b10 *
0-
02
b10 6
#409810000000
1!
1%
1-
12
#409820000000
0!
0%
b11 *
0-
02
b11 6
#409830000000
1!
1%
1-
12
15
#409840000000
0!
0%
b100 *
0-
02
b100 6
#409850000000
1!
1%
1-
12
#409860000000
0!
0%
b101 *
0-
02
b101 6
#409870000000
1!
1%
1-
12
#409880000000
0!
0%
b110 *
0-
02
b110 6
#409890000000
1!
1%
1-
12
#409900000000
0!
0%
b111 *
0-
02
b111 6
#409910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#409920000000
0!
0%
b0 *
0-
02
b0 6
#409930000000
1!
1%
1-
12
#409940000000
0!
0%
b1 *
0-
02
b1 6
#409950000000
1!
1%
1-
12
#409960000000
0!
0%
b10 *
0-
02
b10 6
#409970000000
1!
1%
1-
12
#409980000000
0!
0%
b11 *
0-
02
b11 6
#409990000000
1!
1%
1-
12
15
#410000000000
0!
0%
b100 *
0-
02
b100 6
#410010000000
1!
1%
1-
12
#410020000000
0!
0%
b101 *
0-
02
b101 6
#410030000000
1!
1%
1-
12
#410040000000
0!
0%
b110 *
0-
02
b110 6
#410050000000
1!
1%
1-
12
#410060000000
0!
0%
b111 *
0-
02
b111 6
#410070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#410080000000
0!
0%
b0 *
0-
02
b0 6
#410090000000
1!
1%
1-
12
#410100000000
0!
0%
b1 *
0-
02
b1 6
#410110000000
1!
1%
1-
12
#410120000000
0!
0%
b10 *
0-
02
b10 6
#410130000000
1!
1%
1-
12
#410140000000
0!
0%
b11 *
0-
02
b11 6
#410150000000
1!
1%
1-
12
15
#410160000000
0!
0%
b100 *
0-
02
b100 6
#410170000000
1!
1%
1-
12
#410180000000
0!
0%
b101 *
0-
02
b101 6
#410190000000
1!
1%
1-
12
#410200000000
0!
0%
b110 *
0-
02
b110 6
#410210000000
1!
1%
1-
12
#410220000000
0!
0%
b111 *
0-
02
b111 6
#410230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#410240000000
0!
0%
b0 *
0-
02
b0 6
#410250000000
1!
1%
1-
12
#410260000000
0!
0%
b1 *
0-
02
b1 6
#410270000000
1!
1%
1-
12
#410280000000
0!
0%
b10 *
0-
02
b10 6
#410290000000
1!
1%
1-
12
#410300000000
0!
0%
b11 *
0-
02
b11 6
#410310000000
1!
1%
1-
12
15
#410320000000
0!
0%
b100 *
0-
02
b100 6
#410330000000
1!
1%
1-
12
#410340000000
0!
0%
b101 *
0-
02
b101 6
#410350000000
1!
1%
1-
12
#410360000000
0!
0%
b110 *
0-
02
b110 6
#410370000000
1!
1%
1-
12
#410380000000
0!
0%
b111 *
0-
02
b111 6
#410390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#410400000000
0!
0%
b0 *
0-
02
b0 6
#410410000000
1!
1%
1-
12
#410420000000
0!
0%
b1 *
0-
02
b1 6
#410430000000
1!
1%
1-
12
#410440000000
0!
0%
b10 *
0-
02
b10 6
#410450000000
1!
1%
1-
12
#410460000000
0!
0%
b11 *
0-
02
b11 6
#410470000000
1!
1%
1-
12
15
#410480000000
0!
0%
b100 *
0-
02
b100 6
#410490000000
1!
1%
1-
12
#410500000000
0!
0%
b101 *
0-
02
b101 6
#410510000000
1!
1%
1-
12
#410520000000
0!
0%
b110 *
0-
02
b110 6
#410530000000
1!
1%
1-
12
#410540000000
0!
0%
b111 *
0-
02
b111 6
#410550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#410560000000
0!
0%
b0 *
0-
02
b0 6
#410570000000
1!
1%
1-
12
#410580000000
0!
0%
b1 *
0-
02
b1 6
#410590000000
1!
1%
1-
12
#410600000000
0!
0%
b10 *
0-
02
b10 6
#410610000000
1!
1%
1-
12
#410620000000
0!
0%
b11 *
0-
02
b11 6
#410630000000
1!
1%
1-
12
15
#410640000000
0!
0%
b100 *
0-
02
b100 6
#410650000000
1!
1%
1-
12
#410660000000
0!
0%
b101 *
0-
02
b101 6
#410670000000
1!
1%
1-
12
#410680000000
0!
0%
b110 *
0-
02
b110 6
#410690000000
1!
1%
1-
12
#410700000000
0!
0%
b111 *
0-
02
b111 6
#410710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#410720000000
0!
0%
b0 *
0-
02
b0 6
#410730000000
1!
1%
1-
12
#410740000000
0!
0%
b1 *
0-
02
b1 6
#410750000000
1!
1%
1-
12
#410760000000
0!
0%
b10 *
0-
02
b10 6
#410770000000
1!
1%
1-
12
#410780000000
0!
0%
b11 *
0-
02
b11 6
#410790000000
1!
1%
1-
12
15
#410800000000
0!
0%
b100 *
0-
02
b100 6
#410810000000
1!
1%
1-
12
#410820000000
0!
0%
b101 *
0-
02
b101 6
#410830000000
1!
1%
1-
12
#410840000000
0!
0%
b110 *
0-
02
b110 6
#410850000000
1!
1%
1-
12
#410860000000
0!
0%
b111 *
0-
02
b111 6
#410870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#410880000000
0!
0%
b0 *
0-
02
b0 6
#410890000000
1!
1%
1-
12
#410900000000
0!
0%
b1 *
0-
02
b1 6
#410910000000
1!
1%
1-
12
#410920000000
0!
0%
b10 *
0-
02
b10 6
#410930000000
1!
1%
1-
12
#410940000000
0!
0%
b11 *
0-
02
b11 6
#410950000000
1!
1%
1-
12
15
#410960000000
0!
0%
b100 *
0-
02
b100 6
#410970000000
1!
1%
1-
12
#410980000000
0!
0%
b101 *
0-
02
b101 6
#410990000000
1!
1%
1-
12
#411000000000
0!
0%
b110 *
0-
02
b110 6
#411010000000
1!
1%
1-
12
#411020000000
0!
0%
b111 *
0-
02
b111 6
#411030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#411040000000
0!
0%
b0 *
0-
02
b0 6
#411050000000
1!
1%
1-
12
#411060000000
0!
0%
b1 *
0-
02
b1 6
#411070000000
1!
1%
1-
12
#411080000000
0!
0%
b10 *
0-
02
b10 6
#411090000000
1!
1%
1-
12
#411100000000
0!
0%
b11 *
0-
02
b11 6
#411110000000
1!
1%
1-
12
15
#411120000000
0!
0%
b100 *
0-
02
b100 6
#411130000000
1!
1%
1-
12
#411140000000
0!
0%
b101 *
0-
02
b101 6
#411150000000
1!
1%
1-
12
#411160000000
0!
0%
b110 *
0-
02
b110 6
#411170000000
1!
1%
1-
12
#411180000000
0!
0%
b111 *
0-
02
b111 6
#411190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#411200000000
0!
0%
b0 *
0-
02
b0 6
#411210000000
1!
1%
1-
12
#411220000000
0!
0%
b1 *
0-
02
b1 6
#411230000000
1!
1%
1-
12
#411240000000
0!
0%
b10 *
0-
02
b10 6
#411250000000
1!
1%
1-
12
#411260000000
0!
0%
b11 *
0-
02
b11 6
#411270000000
1!
1%
1-
12
15
#411280000000
0!
0%
b100 *
0-
02
b100 6
#411290000000
1!
1%
1-
12
#411300000000
0!
0%
b101 *
0-
02
b101 6
#411310000000
1!
1%
1-
12
#411320000000
0!
0%
b110 *
0-
02
b110 6
#411330000000
1!
1%
1-
12
#411340000000
0!
0%
b111 *
0-
02
b111 6
#411350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#411360000000
0!
0%
b0 *
0-
02
b0 6
#411370000000
1!
1%
1-
12
#411380000000
0!
0%
b1 *
0-
02
b1 6
#411390000000
1!
1%
1-
12
#411400000000
0!
0%
b10 *
0-
02
b10 6
#411410000000
1!
1%
1-
12
#411420000000
0!
0%
b11 *
0-
02
b11 6
#411430000000
1!
1%
1-
12
15
#411440000000
0!
0%
b100 *
0-
02
b100 6
#411450000000
1!
1%
1-
12
#411460000000
0!
0%
b101 *
0-
02
b101 6
#411470000000
1!
1%
1-
12
#411480000000
0!
0%
b110 *
0-
02
b110 6
#411490000000
1!
1%
1-
12
#411500000000
0!
0%
b111 *
0-
02
b111 6
#411510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#411520000000
0!
0%
b0 *
0-
02
b0 6
#411530000000
1!
1%
1-
12
#411540000000
0!
0%
b1 *
0-
02
b1 6
#411550000000
1!
1%
1-
12
#411560000000
0!
0%
b10 *
0-
02
b10 6
#411570000000
1!
1%
1-
12
#411580000000
0!
0%
b11 *
0-
02
b11 6
#411590000000
1!
1%
1-
12
15
#411600000000
0!
0%
b100 *
0-
02
b100 6
#411610000000
1!
1%
1-
12
#411620000000
0!
0%
b101 *
0-
02
b101 6
#411630000000
1!
1%
1-
12
#411640000000
0!
0%
b110 *
0-
02
b110 6
#411650000000
1!
1%
1-
12
#411660000000
0!
0%
b111 *
0-
02
b111 6
#411670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#411680000000
0!
0%
b0 *
0-
02
b0 6
#411690000000
1!
1%
1-
12
#411700000000
0!
0%
b1 *
0-
02
b1 6
#411710000000
1!
1%
1-
12
#411720000000
0!
0%
b10 *
0-
02
b10 6
#411730000000
1!
1%
1-
12
#411740000000
0!
0%
b11 *
0-
02
b11 6
#411750000000
1!
1%
1-
12
15
#411760000000
0!
0%
b100 *
0-
02
b100 6
#411770000000
1!
1%
1-
12
#411780000000
0!
0%
b101 *
0-
02
b101 6
#411790000000
1!
1%
1-
12
#411800000000
0!
0%
b110 *
0-
02
b110 6
#411810000000
1!
1%
1-
12
#411820000000
0!
0%
b111 *
0-
02
b111 6
#411830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#411840000000
0!
0%
b0 *
0-
02
b0 6
#411850000000
1!
1%
1-
12
#411860000000
0!
0%
b1 *
0-
02
b1 6
#411870000000
1!
1%
1-
12
#411880000000
0!
0%
b10 *
0-
02
b10 6
#411890000000
1!
1%
1-
12
#411900000000
0!
0%
b11 *
0-
02
b11 6
#411910000000
1!
1%
1-
12
15
#411920000000
0!
0%
b100 *
0-
02
b100 6
#411930000000
1!
1%
1-
12
#411940000000
0!
0%
b101 *
0-
02
b101 6
#411950000000
1!
1%
1-
12
#411960000000
0!
0%
b110 *
0-
02
b110 6
#411970000000
1!
1%
1-
12
#411980000000
0!
0%
b111 *
0-
02
b111 6
#411990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#412000000000
0!
0%
b0 *
0-
02
b0 6
#412010000000
1!
1%
1-
12
#412020000000
0!
0%
b1 *
0-
02
b1 6
#412030000000
1!
1%
1-
12
#412040000000
0!
0%
b10 *
0-
02
b10 6
#412050000000
1!
1%
1-
12
#412060000000
0!
0%
b11 *
0-
02
b11 6
#412070000000
1!
1%
1-
12
15
#412080000000
0!
0%
b100 *
0-
02
b100 6
#412090000000
1!
1%
1-
12
#412100000000
0!
0%
b101 *
0-
02
b101 6
#412110000000
1!
1%
1-
12
#412120000000
0!
0%
b110 *
0-
02
b110 6
#412130000000
1!
1%
1-
12
#412140000000
0!
0%
b111 *
0-
02
b111 6
#412150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#412160000000
0!
0%
b0 *
0-
02
b0 6
#412170000000
1!
1%
1-
12
#412180000000
0!
0%
b1 *
0-
02
b1 6
#412190000000
1!
1%
1-
12
#412200000000
0!
0%
b10 *
0-
02
b10 6
#412210000000
1!
1%
1-
12
#412220000000
0!
0%
b11 *
0-
02
b11 6
#412230000000
1!
1%
1-
12
15
#412240000000
0!
0%
b100 *
0-
02
b100 6
#412250000000
1!
1%
1-
12
#412260000000
0!
0%
b101 *
0-
02
b101 6
#412270000000
1!
1%
1-
12
#412280000000
0!
0%
b110 *
0-
02
b110 6
#412290000000
1!
1%
1-
12
#412300000000
0!
0%
b111 *
0-
02
b111 6
#412310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#412320000000
0!
0%
b0 *
0-
02
b0 6
#412330000000
1!
1%
1-
12
#412340000000
0!
0%
b1 *
0-
02
b1 6
#412350000000
1!
1%
1-
12
#412360000000
0!
0%
b10 *
0-
02
b10 6
#412370000000
1!
1%
1-
12
#412380000000
0!
0%
b11 *
0-
02
b11 6
#412390000000
1!
1%
1-
12
15
#412400000000
0!
0%
b100 *
0-
02
b100 6
#412410000000
1!
1%
1-
12
#412420000000
0!
0%
b101 *
0-
02
b101 6
#412430000000
1!
1%
1-
12
#412440000000
0!
0%
b110 *
0-
02
b110 6
#412450000000
1!
1%
1-
12
#412460000000
0!
0%
b111 *
0-
02
b111 6
#412470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#412480000000
0!
0%
b0 *
0-
02
b0 6
#412490000000
1!
1%
1-
12
#412500000000
0!
0%
b1 *
0-
02
b1 6
#412510000000
1!
1%
1-
12
#412520000000
0!
0%
b10 *
0-
02
b10 6
#412530000000
1!
1%
1-
12
#412540000000
0!
0%
b11 *
0-
02
b11 6
#412550000000
1!
1%
1-
12
15
#412560000000
0!
0%
b100 *
0-
02
b100 6
#412570000000
1!
1%
1-
12
#412580000000
0!
0%
b101 *
0-
02
b101 6
#412590000000
1!
1%
1-
12
#412600000000
0!
0%
b110 *
0-
02
b110 6
#412610000000
1!
1%
1-
12
#412620000000
0!
0%
b111 *
0-
02
b111 6
#412630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#412640000000
0!
0%
b0 *
0-
02
b0 6
#412650000000
1!
1%
1-
12
#412660000000
0!
0%
b1 *
0-
02
b1 6
#412670000000
1!
1%
1-
12
#412680000000
0!
0%
b10 *
0-
02
b10 6
#412690000000
1!
1%
1-
12
#412700000000
0!
0%
b11 *
0-
02
b11 6
#412710000000
1!
1%
1-
12
15
#412720000000
0!
0%
b100 *
0-
02
b100 6
#412730000000
1!
1%
1-
12
#412740000000
0!
0%
b101 *
0-
02
b101 6
#412750000000
1!
1%
1-
12
#412760000000
0!
0%
b110 *
0-
02
b110 6
#412770000000
1!
1%
1-
12
#412780000000
0!
0%
b111 *
0-
02
b111 6
#412790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#412800000000
0!
0%
b0 *
0-
02
b0 6
#412810000000
1!
1%
1-
12
#412820000000
0!
0%
b1 *
0-
02
b1 6
#412830000000
1!
1%
1-
12
#412840000000
0!
0%
b10 *
0-
02
b10 6
#412850000000
1!
1%
1-
12
#412860000000
0!
0%
b11 *
0-
02
b11 6
#412870000000
1!
1%
1-
12
15
#412880000000
0!
0%
b100 *
0-
02
b100 6
#412890000000
1!
1%
1-
12
#412900000000
0!
0%
b101 *
0-
02
b101 6
#412910000000
1!
1%
1-
12
#412920000000
0!
0%
b110 *
0-
02
b110 6
#412930000000
1!
1%
1-
12
#412940000000
0!
0%
b111 *
0-
02
b111 6
#412950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#412960000000
0!
0%
b0 *
0-
02
b0 6
#412970000000
1!
1%
1-
12
#412980000000
0!
0%
b1 *
0-
02
b1 6
#412990000000
1!
1%
1-
12
#413000000000
0!
0%
b10 *
0-
02
b10 6
#413010000000
1!
1%
1-
12
#413020000000
0!
0%
b11 *
0-
02
b11 6
#413030000000
1!
1%
1-
12
15
#413040000000
0!
0%
b100 *
0-
02
b100 6
#413050000000
1!
1%
1-
12
#413060000000
0!
0%
b101 *
0-
02
b101 6
#413070000000
1!
1%
1-
12
#413080000000
0!
0%
b110 *
0-
02
b110 6
#413090000000
1!
1%
1-
12
#413100000000
0!
0%
b111 *
0-
02
b111 6
#413110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#413120000000
0!
0%
b0 *
0-
02
b0 6
#413130000000
1!
1%
1-
12
#413140000000
0!
0%
b1 *
0-
02
b1 6
#413150000000
1!
1%
1-
12
#413160000000
0!
0%
b10 *
0-
02
b10 6
#413170000000
1!
1%
1-
12
#413180000000
0!
0%
b11 *
0-
02
b11 6
#413190000000
1!
1%
1-
12
15
#413200000000
0!
0%
b100 *
0-
02
b100 6
#413210000000
1!
1%
1-
12
#413220000000
0!
0%
b101 *
0-
02
b101 6
#413230000000
1!
1%
1-
12
#413240000000
0!
0%
b110 *
0-
02
b110 6
#413250000000
1!
1%
1-
12
#413260000000
0!
0%
b111 *
0-
02
b111 6
#413270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#413280000000
0!
0%
b0 *
0-
02
b0 6
#413290000000
1!
1%
1-
12
#413300000000
0!
0%
b1 *
0-
02
b1 6
#413310000000
1!
1%
1-
12
#413320000000
0!
0%
b10 *
0-
02
b10 6
#413330000000
1!
1%
1-
12
#413340000000
0!
0%
b11 *
0-
02
b11 6
#413350000000
1!
1%
1-
12
15
#413360000000
0!
0%
b100 *
0-
02
b100 6
#413370000000
1!
1%
1-
12
#413380000000
0!
0%
b101 *
0-
02
b101 6
#413390000000
1!
1%
1-
12
#413400000000
0!
0%
b110 *
0-
02
b110 6
#413410000000
1!
1%
1-
12
#413420000000
0!
0%
b111 *
0-
02
b111 6
#413430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#413440000000
0!
0%
b0 *
0-
02
b0 6
#413450000000
1!
1%
1-
12
#413460000000
0!
0%
b1 *
0-
02
b1 6
#413470000000
1!
1%
1-
12
#413480000000
0!
0%
b10 *
0-
02
b10 6
#413490000000
1!
1%
1-
12
#413500000000
0!
0%
b11 *
0-
02
b11 6
#413510000000
1!
1%
1-
12
15
#413520000000
0!
0%
b100 *
0-
02
b100 6
#413530000000
1!
1%
1-
12
#413540000000
0!
0%
b101 *
0-
02
b101 6
#413550000000
1!
1%
1-
12
#413560000000
0!
0%
b110 *
0-
02
b110 6
#413570000000
1!
1%
1-
12
#413580000000
0!
0%
b111 *
0-
02
b111 6
#413590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#413600000000
0!
0%
b0 *
0-
02
b0 6
#413610000000
1!
1%
1-
12
#413620000000
0!
0%
b1 *
0-
02
b1 6
#413630000000
1!
1%
1-
12
#413640000000
0!
0%
b10 *
0-
02
b10 6
#413650000000
1!
1%
1-
12
#413660000000
0!
0%
b11 *
0-
02
b11 6
#413670000000
1!
1%
1-
12
15
#413680000000
0!
0%
b100 *
0-
02
b100 6
#413690000000
1!
1%
1-
12
#413700000000
0!
0%
b101 *
0-
02
b101 6
#413710000000
1!
1%
1-
12
#413720000000
0!
0%
b110 *
0-
02
b110 6
#413730000000
1!
1%
1-
12
#413740000000
0!
0%
b111 *
0-
02
b111 6
#413750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#413760000000
0!
0%
b0 *
0-
02
b0 6
#413770000000
1!
1%
1-
12
#413780000000
0!
0%
b1 *
0-
02
b1 6
#413790000000
1!
1%
1-
12
#413800000000
0!
0%
b10 *
0-
02
b10 6
#413810000000
1!
1%
1-
12
#413820000000
0!
0%
b11 *
0-
02
b11 6
#413830000000
1!
1%
1-
12
15
#413840000000
0!
0%
b100 *
0-
02
b100 6
#413850000000
1!
1%
1-
12
#413860000000
0!
0%
b101 *
0-
02
b101 6
#413870000000
1!
1%
1-
12
#413880000000
0!
0%
b110 *
0-
02
b110 6
#413890000000
1!
1%
1-
12
#413900000000
0!
0%
b111 *
0-
02
b111 6
#413910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#413920000000
0!
0%
b0 *
0-
02
b0 6
#413930000000
1!
1%
1-
12
#413940000000
0!
0%
b1 *
0-
02
b1 6
#413950000000
1!
1%
1-
12
#413960000000
0!
0%
b10 *
0-
02
b10 6
#413970000000
1!
1%
1-
12
#413980000000
0!
0%
b11 *
0-
02
b11 6
#413990000000
1!
1%
1-
12
15
#414000000000
0!
0%
b100 *
0-
02
b100 6
#414010000000
1!
1%
1-
12
#414020000000
0!
0%
b101 *
0-
02
b101 6
#414030000000
1!
1%
1-
12
#414040000000
0!
0%
b110 *
0-
02
b110 6
#414050000000
1!
1%
1-
12
#414060000000
0!
0%
b111 *
0-
02
b111 6
#414070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#414080000000
0!
0%
b0 *
0-
02
b0 6
#414090000000
1!
1%
1-
12
#414100000000
0!
0%
b1 *
0-
02
b1 6
#414110000000
1!
1%
1-
12
#414120000000
0!
0%
b10 *
0-
02
b10 6
#414130000000
1!
1%
1-
12
#414140000000
0!
0%
b11 *
0-
02
b11 6
#414150000000
1!
1%
1-
12
15
#414160000000
0!
0%
b100 *
0-
02
b100 6
#414170000000
1!
1%
1-
12
#414180000000
0!
0%
b101 *
0-
02
b101 6
#414190000000
1!
1%
1-
12
#414200000000
0!
0%
b110 *
0-
02
b110 6
#414210000000
1!
1%
1-
12
#414220000000
0!
0%
b111 *
0-
02
b111 6
#414230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#414240000000
0!
0%
b0 *
0-
02
b0 6
#414250000000
1!
1%
1-
12
#414260000000
0!
0%
b1 *
0-
02
b1 6
#414270000000
1!
1%
1-
12
#414280000000
0!
0%
b10 *
0-
02
b10 6
#414290000000
1!
1%
1-
12
#414300000000
0!
0%
b11 *
0-
02
b11 6
#414310000000
1!
1%
1-
12
15
#414320000000
0!
0%
b100 *
0-
02
b100 6
#414330000000
1!
1%
1-
12
#414340000000
0!
0%
b101 *
0-
02
b101 6
#414350000000
1!
1%
1-
12
#414360000000
0!
0%
b110 *
0-
02
b110 6
#414370000000
1!
1%
1-
12
#414380000000
0!
0%
b111 *
0-
02
b111 6
#414390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#414400000000
0!
0%
b0 *
0-
02
b0 6
#414410000000
1!
1%
1-
12
#414420000000
0!
0%
b1 *
0-
02
b1 6
#414430000000
1!
1%
1-
12
#414440000000
0!
0%
b10 *
0-
02
b10 6
#414450000000
1!
1%
1-
12
#414460000000
0!
0%
b11 *
0-
02
b11 6
#414470000000
1!
1%
1-
12
15
#414480000000
0!
0%
b100 *
0-
02
b100 6
#414490000000
1!
1%
1-
12
#414500000000
0!
0%
b101 *
0-
02
b101 6
#414510000000
1!
1%
1-
12
#414520000000
0!
0%
b110 *
0-
02
b110 6
#414530000000
1!
1%
1-
12
#414540000000
0!
0%
b111 *
0-
02
b111 6
#414550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#414560000000
0!
0%
b0 *
0-
02
b0 6
#414570000000
1!
1%
1-
12
#414580000000
0!
0%
b1 *
0-
02
b1 6
#414590000000
1!
1%
1-
12
#414600000000
0!
0%
b10 *
0-
02
b10 6
#414610000000
1!
1%
1-
12
#414620000000
0!
0%
b11 *
0-
02
b11 6
#414630000000
1!
1%
1-
12
15
#414640000000
0!
0%
b100 *
0-
02
b100 6
#414650000000
1!
1%
1-
12
#414660000000
0!
0%
b101 *
0-
02
b101 6
#414670000000
1!
1%
1-
12
#414680000000
0!
0%
b110 *
0-
02
b110 6
#414690000000
1!
1%
1-
12
#414700000000
0!
0%
b111 *
0-
02
b111 6
#414710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#414720000000
0!
0%
b0 *
0-
02
b0 6
#414730000000
1!
1%
1-
12
#414740000000
0!
0%
b1 *
0-
02
b1 6
#414750000000
1!
1%
1-
12
#414760000000
0!
0%
b10 *
0-
02
b10 6
#414770000000
1!
1%
1-
12
#414780000000
0!
0%
b11 *
0-
02
b11 6
#414790000000
1!
1%
1-
12
15
#414800000000
0!
0%
b100 *
0-
02
b100 6
#414810000000
1!
1%
1-
12
#414820000000
0!
0%
b101 *
0-
02
b101 6
#414830000000
1!
1%
1-
12
#414840000000
0!
0%
b110 *
0-
02
b110 6
#414850000000
1!
1%
1-
12
#414860000000
0!
0%
b111 *
0-
02
b111 6
#414870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#414880000000
0!
0%
b0 *
0-
02
b0 6
#414890000000
1!
1%
1-
12
#414900000000
0!
0%
b1 *
0-
02
b1 6
#414910000000
1!
1%
1-
12
#414920000000
0!
0%
b10 *
0-
02
b10 6
#414930000000
1!
1%
1-
12
#414940000000
0!
0%
b11 *
0-
02
b11 6
#414950000000
1!
1%
1-
12
15
#414960000000
0!
0%
b100 *
0-
02
b100 6
#414970000000
1!
1%
1-
12
#414980000000
0!
0%
b101 *
0-
02
b101 6
#414990000000
1!
1%
1-
12
#415000000000
0!
0%
b110 *
0-
02
b110 6
#415010000000
1!
1%
1-
12
#415020000000
0!
0%
b111 *
0-
02
b111 6
#415030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#415040000000
0!
0%
b0 *
0-
02
b0 6
#415050000000
1!
1%
1-
12
#415060000000
0!
0%
b1 *
0-
02
b1 6
#415070000000
1!
1%
1-
12
#415080000000
0!
0%
b10 *
0-
02
b10 6
#415090000000
1!
1%
1-
12
#415100000000
0!
0%
b11 *
0-
02
b11 6
#415110000000
1!
1%
1-
12
15
#415120000000
0!
0%
b100 *
0-
02
b100 6
#415130000000
1!
1%
1-
12
#415140000000
0!
0%
b101 *
0-
02
b101 6
#415150000000
1!
1%
1-
12
#415160000000
0!
0%
b110 *
0-
02
b110 6
#415170000000
1!
1%
1-
12
#415180000000
0!
0%
b111 *
0-
02
b111 6
#415190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#415200000000
0!
0%
b0 *
0-
02
b0 6
#415210000000
1!
1%
1-
12
#415220000000
0!
0%
b1 *
0-
02
b1 6
#415230000000
1!
1%
1-
12
#415240000000
0!
0%
b10 *
0-
02
b10 6
#415250000000
1!
1%
1-
12
#415260000000
0!
0%
b11 *
0-
02
b11 6
#415270000000
1!
1%
1-
12
15
#415280000000
0!
0%
b100 *
0-
02
b100 6
#415290000000
1!
1%
1-
12
#415300000000
0!
0%
b101 *
0-
02
b101 6
#415310000000
1!
1%
1-
12
#415320000000
0!
0%
b110 *
0-
02
b110 6
#415330000000
1!
1%
1-
12
#415340000000
0!
0%
b111 *
0-
02
b111 6
#415350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#415360000000
0!
0%
b0 *
0-
02
b0 6
#415370000000
1!
1%
1-
12
#415380000000
0!
0%
b1 *
0-
02
b1 6
#415390000000
1!
1%
1-
12
#415400000000
0!
0%
b10 *
0-
02
b10 6
#415410000000
1!
1%
1-
12
#415420000000
0!
0%
b11 *
0-
02
b11 6
#415430000000
1!
1%
1-
12
15
#415440000000
0!
0%
b100 *
0-
02
b100 6
#415450000000
1!
1%
1-
12
#415460000000
0!
0%
b101 *
0-
02
b101 6
#415470000000
1!
1%
1-
12
#415480000000
0!
0%
b110 *
0-
02
b110 6
#415490000000
1!
1%
1-
12
#415500000000
0!
0%
b111 *
0-
02
b111 6
#415510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#415520000000
0!
0%
b0 *
0-
02
b0 6
#415530000000
1!
1%
1-
12
#415540000000
0!
0%
b1 *
0-
02
b1 6
#415550000000
1!
1%
1-
12
#415560000000
0!
0%
b10 *
0-
02
b10 6
#415570000000
1!
1%
1-
12
#415580000000
0!
0%
b11 *
0-
02
b11 6
#415590000000
1!
1%
1-
12
15
#415600000000
0!
0%
b100 *
0-
02
b100 6
#415610000000
1!
1%
1-
12
#415620000000
0!
0%
b101 *
0-
02
b101 6
#415630000000
1!
1%
1-
12
#415640000000
0!
0%
b110 *
0-
02
b110 6
#415650000000
1!
1%
1-
12
#415660000000
0!
0%
b111 *
0-
02
b111 6
#415670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#415680000000
0!
0%
b0 *
0-
02
b0 6
#415690000000
1!
1%
1-
12
#415700000000
0!
0%
b1 *
0-
02
b1 6
#415710000000
1!
1%
1-
12
#415720000000
0!
0%
b10 *
0-
02
b10 6
#415730000000
1!
1%
1-
12
#415740000000
0!
0%
b11 *
0-
02
b11 6
#415750000000
1!
1%
1-
12
15
#415760000000
0!
0%
b100 *
0-
02
b100 6
#415770000000
1!
1%
1-
12
#415780000000
0!
0%
b101 *
0-
02
b101 6
#415790000000
1!
1%
1-
12
#415800000000
0!
0%
b110 *
0-
02
b110 6
#415810000000
1!
1%
1-
12
#415820000000
0!
0%
b111 *
0-
02
b111 6
#415830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#415840000000
0!
0%
b0 *
0-
02
b0 6
#415850000000
1!
1%
1-
12
#415860000000
0!
0%
b1 *
0-
02
b1 6
#415870000000
1!
1%
1-
12
#415880000000
0!
0%
b10 *
0-
02
b10 6
#415890000000
1!
1%
1-
12
#415900000000
0!
0%
b11 *
0-
02
b11 6
#415910000000
1!
1%
1-
12
15
#415920000000
0!
0%
b100 *
0-
02
b100 6
#415930000000
1!
1%
1-
12
#415940000000
0!
0%
b101 *
0-
02
b101 6
#415950000000
1!
1%
1-
12
#415960000000
0!
0%
b110 *
0-
02
b110 6
#415970000000
1!
1%
1-
12
#415980000000
0!
0%
b111 *
0-
02
b111 6
#415990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#416000000000
0!
0%
b0 *
0-
02
b0 6
#416010000000
1!
1%
1-
12
#416020000000
0!
0%
b1 *
0-
02
b1 6
#416030000000
1!
1%
1-
12
#416040000000
0!
0%
b10 *
0-
02
b10 6
#416050000000
1!
1%
1-
12
#416060000000
0!
0%
b11 *
0-
02
b11 6
#416070000000
1!
1%
1-
12
15
#416080000000
0!
0%
b100 *
0-
02
b100 6
#416090000000
1!
1%
1-
12
#416100000000
0!
0%
b101 *
0-
02
b101 6
#416110000000
1!
1%
1-
12
#416120000000
0!
0%
b110 *
0-
02
b110 6
#416130000000
1!
1%
1-
12
#416140000000
0!
0%
b111 *
0-
02
b111 6
#416150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#416160000000
0!
0%
b0 *
0-
02
b0 6
#416170000000
1!
1%
1-
12
#416180000000
0!
0%
b1 *
0-
02
b1 6
#416190000000
1!
1%
1-
12
#416200000000
0!
0%
b10 *
0-
02
b10 6
#416210000000
1!
1%
1-
12
#416220000000
0!
0%
b11 *
0-
02
b11 6
#416230000000
1!
1%
1-
12
15
#416240000000
0!
0%
b100 *
0-
02
b100 6
#416250000000
1!
1%
1-
12
#416260000000
0!
0%
b101 *
0-
02
b101 6
#416270000000
1!
1%
1-
12
#416280000000
0!
0%
b110 *
0-
02
b110 6
#416290000000
1!
1%
1-
12
#416300000000
0!
0%
b111 *
0-
02
b111 6
#416310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#416320000000
0!
0%
b0 *
0-
02
b0 6
#416330000000
1!
1%
1-
12
#416340000000
0!
0%
b1 *
0-
02
b1 6
#416350000000
1!
1%
1-
12
#416360000000
0!
0%
b10 *
0-
02
b10 6
#416370000000
1!
1%
1-
12
#416380000000
0!
0%
b11 *
0-
02
b11 6
#416390000000
1!
1%
1-
12
15
#416400000000
0!
0%
b100 *
0-
02
b100 6
#416410000000
1!
1%
1-
12
#416420000000
0!
0%
b101 *
0-
02
b101 6
#416430000000
1!
1%
1-
12
#416440000000
0!
0%
b110 *
0-
02
b110 6
#416450000000
1!
1%
1-
12
#416460000000
0!
0%
b111 *
0-
02
b111 6
#416470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#416480000000
0!
0%
b0 *
0-
02
b0 6
#416490000000
1!
1%
1-
12
#416500000000
0!
0%
b1 *
0-
02
b1 6
#416510000000
1!
1%
1-
12
#416520000000
0!
0%
b10 *
0-
02
b10 6
#416530000000
1!
1%
1-
12
#416540000000
0!
0%
b11 *
0-
02
b11 6
#416550000000
1!
1%
1-
12
15
#416560000000
0!
0%
b100 *
0-
02
b100 6
#416570000000
1!
1%
1-
12
#416580000000
0!
0%
b101 *
0-
02
b101 6
#416590000000
1!
1%
1-
12
#416600000000
0!
0%
b110 *
0-
02
b110 6
#416610000000
1!
1%
1-
12
#416620000000
0!
0%
b111 *
0-
02
b111 6
#416630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#416640000000
0!
0%
b0 *
0-
02
b0 6
#416650000000
1!
1%
1-
12
#416660000000
0!
0%
b1 *
0-
02
b1 6
#416670000000
1!
1%
1-
12
#416680000000
0!
0%
b10 *
0-
02
b10 6
#416690000000
1!
1%
1-
12
#416700000000
0!
0%
b11 *
0-
02
b11 6
#416710000000
1!
1%
1-
12
15
#416720000000
0!
0%
b100 *
0-
02
b100 6
#416730000000
1!
1%
1-
12
#416740000000
0!
0%
b101 *
0-
02
b101 6
#416750000000
1!
1%
1-
12
#416760000000
0!
0%
b110 *
0-
02
b110 6
#416770000000
1!
1%
1-
12
#416780000000
0!
0%
b111 *
0-
02
b111 6
#416790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#416800000000
0!
0%
b0 *
0-
02
b0 6
#416810000000
1!
1%
1-
12
#416820000000
0!
0%
b1 *
0-
02
b1 6
#416830000000
1!
1%
1-
12
#416840000000
0!
0%
b10 *
0-
02
b10 6
#416850000000
1!
1%
1-
12
#416860000000
0!
0%
b11 *
0-
02
b11 6
#416870000000
1!
1%
1-
12
15
#416880000000
0!
0%
b100 *
0-
02
b100 6
#416890000000
1!
1%
1-
12
#416900000000
0!
0%
b101 *
0-
02
b101 6
#416910000000
1!
1%
1-
12
#416920000000
0!
0%
b110 *
0-
02
b110 6
#416930000000
1!
1%
1-
12
#416940000000
0!
0%
b111 *
0-
02
b111 6
#416950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#416960000000
0!
0%
b0 *
0-
02
b0 6
#416970000000
1!
1%
1-
12
#416980000000
0!
0%
b1 *
0-
02
b1 6
#416990000000
1!
1%
1-
12
#417000000000
0!
0%
b10 *
0-
02
b10 6
#417010000000
1!
1%
1-
12
#417020000000
0!
0%
b11 *
0-
02
b11 6
#417030000000
1!
1%
1-
12
15
#417040000000
0!
0%
b100 *
0-
02
b100 6
#417050000000
1!
1%
1-
12
#417060000000
0!
0%
b101 *
0-
02
b101 6
#417070000000
1!
1%
1-
12
#417080000000
0!
0%
b110 *
0-
02
b110 6
#417090000000
1!
1%
1-
12
#417100000000
0!
0%
b111 *
0-
02
b111 6
#417110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#417120000000
0!
0%
b0 *
0-
02
b0 6
#417130000000
1!
1%
1-
12
#417140000000
0!
0%
b1 *
0-
02
b1 6
#417150000000
1!
1%
1-
12
#417160000000
0!
0%
b10 *
0-
02
b10 6
#417170000000
1!
1%
1-
12
#417180000000
0!
0%
b11 *
0-
02
b11 6
#417190000000
1!
1%
1-
12
15
#417200000000
0!
0%
b100 *
0-
02
b100 6
#417210000000
1!
1%
1-
12
#417220000000
0!
0%
b101 *
0-
02
b101 6
#417230000000
1!
1%
1-
12
#417240000000
0!
0%
b110 *
0-
02
b110 6
#417250000000
1!
1%
1-
12
#417260000000
0!
0%
b111 *
0-
02
b111 6
#417270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#417280000000
0!
0%
b0 *
0-
02
b0 6
#417290000000
1!
1%
1-
12
#417300000000
0!
0%
b1 *
0-
02
b1 6
#417310000000
1!
1%
1-
12
#417320000000
0!
0%
b10 *
0-
02
b10 6
#417330000000
1!
1%
1-
12
#417340000000
0!
0%
b11 *
0-
02
b11 6
#417350000000
1!
1%
1-
12
15
#417360000000
0!
0%
b100 *
0-
02
b100 6
#417370000000
1!
1%
1-
12
#417380000000
0!
0%
b101 *
0-
02
b101 6
#417390000000
1!
1%
1-
12
#417400000000
0!
0%
b110 *
0-
02
b110 6
#417410000000
1!
1%
1-
12
#417420000000
0!
0%
b111 *
0-
02
b111 6
#417430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#417440000000
0!
0%
b0 *
0-
02
b0 6
#417450000000
1!
1%
1-
12
#417460000000
0!
0%
b1 *
0-
02
b1 6
#417470000000
1!
1%
1-
12
#417480000000
0!
0%
b10 *
0-
02
b10 6
#417490000000
1!
1%
1-
12
#417500000000
0!
0%
b11 *
0-
02
b11 6
#417510000000
1!
1%
1-
12
15
#417520000000
0!
0%
b100 *
0-
02
b100 6
#417530000000
1!
1%
1-
12
#417540000000
0!
0%
b101 *
0-
02
b101 6
#417550000000
1!
1%
1-
12
#417560000000
0!
0%
b110 *
0-
02
b110 6
#417570000000
1!
1%
1-
12
#417580000000
0!
0%
b111 *
0-
02
b111 6
#417590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#417600000000
0!
0%
b0 *
0-
02
b0 6
#417610000000
1!
1%
1-
12
#417620000000
0!
0%
b1 *
0-
02
b1 6
#417630000000
1!
1%
1-
12
#417640000000
0!
0%
b10 *
0-
02
b10 6
#417650000000
1!
1%
1-
12
#417660000000
0!
0%
b11 *
0-
02
b11 6
#417670000000
1!
1%
1-
12
15
#417680000000
0!
0%
b100 *
0-
02
b100 6
#417690000000
1!
1%
1-
12
#417700000000
0!
0%
b101 *
0-
02
b101 6
#417710000000
1!
1%
1-
12
#417720000000
0!
0%
b110 *
0-
02
b110 6
#417730000000
1!
1%
1-
12
#417740000000
0!
0%
b111 *
0-
02
b111 6
#417750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#417760000000
0!
0%
b0 *
0-
02
b0 6
#417770000000
1!
1%
1-
12
#417780000000
0!
0%
b1 *
0-
02
b1 6
#417790000000
1!
1%
1-
12
#417800000000
0!
0%
b10 *
0-
02
b10 6
#417810000000
1!
1%
1-
12
#417820000000
0!
0%
b11 *
0-
02
b11 6
#417830000000
1!
1%
1-
12
15
#417840000000
0!
0%
b100 *
0-
02
b100 6
#417850000000
1!
1%
1-
12
#417860000000
0!
0%
b101 *
0-
02
b101 6
#417870000000
1!
1%
1-
12
#417880000000
0!
0%
b110 *
0-
02
b110 6
#417890000000
1!
1%
1-
12
#417900000000
0!
0%
b111 *
0-
02
b111 6
#417910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#417920000000
0!
0%
b0 *
0-
02
b0 6
#417930000000
1!
1%
1-
12
#417940000000
0!
0%
b1 *
0-
02
b1 6
#417950000000
1!
1%
1-
12
#417960000000
0!
0%
b10 *
0-
02
b10 6
#417970000000
1!
1%
1-
12
#417980000000
0!
0%
b11 *
0-
02
b11 6
#417990000000
1!
1%
1-
12
15
#418000000000
0!
0%
b100 *
0-
02
b100 6
#418010000000
1!
1%
1-
12
#418020000000
0!
0%
b101 *
0-
02
b101 6
#418030000000
1!
1%
1-
12
#418040000000
0!
0%
b110 *
0-
02
b110 6
#418050000000
1!
1%
1-
12
#418060000000
0!
0%
b111 *
0-
02
b111 6
#418070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#418080000000
0!
0%
b0 *
0-
02
b0 6
#418090000000
1!
1%
1-
12
#418100000000
0!
0%
b1 *
0-
02
b1 6
#418110000000
1!
1%
1-
12
#418120000000
0!
0%
b10 *
0-
02
b10 6
#418130000000
1!
1%
1-
12
#418140000000
0!
0%
b11 *
0-
02
b11 6
#418150000000
1!
1%
1-
12
15
#418160000000
0!
0%
b100 *
0-
02
b100 6
#418170000000
1!
1%
1-
12
#418180000000
0!
0%
b101 *
0-
02
b101 6
#418190000000
1!
1%
1-
12
#418200000000
0!
0%
b110 *
0-
02
b110 6
#418210000000
1!
1%
1-
12
#418220000000
0!
0%
b111 *
0-
02
b111 6
#418230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#418240000000
0!
0%
b0 *
0-
02
b0 6
#418250000000
1!
1%
1-
12
#418260000000
0!
0%
b1 *
0-
02
b1 6
#418270000000
1!
1%
1-
12
#418280000000
0!
0%
b10 *
0-
02
b10 6
#418290000000
1!
1%
1-
12
#418300000000
0!
0%
b11 *
0-
02
b11 6
#418310000000
1!
1%
1-
12
15
#418320000000
0!
0%
b100 *
0-
02
b100 6
#418330000000
1!
1%
1-
12
#418340000000
0!
0%
b101 *
0-
02
b101 6
#418350000000
1!
1%
1-
12
#418360000000
0!
0%
b110 *
0-
02
b110 6
#418370000000
1!
1%
1-
12
#418380000000
0!
0%
b111 *
0-
02
b111 6
#418390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#418400000000
0!
0%
b0 *
0-
02
b0 6
#418410000000
1!
1%
1-
12
#418420000000
0!
0%
b1 *
0-
02
b1 6
#418430000000
1!
1%
1-
12
#418440000000
0!
0%
b10 *
0-
02
b10 6
#418450000000
1!
1%
1-
12
#418460000000
0!
0%
b11 *
0-
02
b11 6
#418470000000
1!
1%
1-
12
15
#418480000000
0!
0%
b100 *
0-
02
b100 6
#418490000000
1!
1%
1-
12
#418500000000
0!
0%
b101 *
0-
02
b101 6
#418510000000
1!
1%
1-
12
#418520000000
0!
0%
b110 *
0-
02
b110 6
#418530000000
1!
1%
1-
12
#418540000000
0!
0%
b111 *
0-
02
b111 6
#418550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#418560000000
0!
0%
b0 *
0-
02
b0 6
#418570000000
1!
1%
1-
12
#418580000000
0!
0%
b1 *
0-
02
b1 6
#418590000000
1!
1%
1-
12
#418600000000
0!
0%
b10 *
0-
02
b10 6
#418610000000
1!
1%
1-
12
#418620000000
0!
0%
b11 *
0-
02
b11 6
#418630000000
1!
1%
1-
12
15
#418640000000
0!
0%
b100 *
0-
02
b100 6
#418650000000
1!
1%
1-
12
#418660000000
0!
0%
b101 *
0-
02
b101 6
#418670000000
1!
1%
1-
12
#418680000000
0!
0%
b110 *
0-
02
b110 6
#418690000000
1!
1%
1-
12
#418700000000
0!
0%
b111 *
0-
02
b111 6
#418710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#418720000000
0!
0%
b0 *
0-
02
b0 6
#418730000000
1!
1%
1-
12
#418740000000
0!
0%
b1 *
0-
02
b1 6
#418750000000
1!
1%
1-
12
#418760000000
0!
0%
b10 *
0-
02
b10 6
#418770000000
1!
1%
1-
12
#418780000000
0!
0%
b11 *
0-
02
b11 6
#418790000000
1!
1%
1-
12
15
#418800000000
0!
0%
b100 *
0-
02
b100 6
#418810000000
1!
1%
1-
12
#418820000000
0!
0%
b101 *
0-
02
b101 6
#418830000000
1!
1%
1-
12
#418840000000
0!
0%
b110 *
0-
02
b110 6
#418850000000
1!
1%
1-
12
#418860000000
0!
0%
b111 *
0-
02
b111 6
#418870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#418880000000
0!
0%
b0 *
0-
02
b0 6
#418890000000
1!
1%
1-
12
#418900000000
0!
0%
b1 *
0-
02
b1 6
#418910000000
1!
1%
1-
12
#418920000000
0!
0%
b10 *
0-
02
b10 6
#418930000000
1!
1%
1-
12
#418940000000
0!
0%
b11 *
0-
02
b11 6
#418950000000
1!
1%
1-
12
15
#418960000000
0!
0%
b100 *
0-
02
b100 6
#418970000000
1!
1%
1-
12
#418980000000
0!
0%
b101 *
0-
02
b101 6
#418990000000
1!
1%
1-
12
#419000000000
0!
0%
b110 *
0-
02
b110 6
#419010000000
1!
1%
1-
12
#419020000000
0!
0%
b111 *
0-
02
b111 6
#419030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#419040000000
0!
0%
b0 *
0-
02
b0 6
#419050000000
1!
1%
1-
12
#419060000000
0!
0%
b1 *
0-
02
b1 6
#419070000000
1!
1%
1-
12
#419080000000
0!
0%
b10 *
0-
02
b10 6
#419090000000
1!
1%
1-
12
#419100000000
0!
0%
b11 *
0-
02
b11 6
#419110000000
1!
1%
1-
12
15
#419120000000
0!
0%
b100 *
0-
02
b100 6
#419130000000
1!
1%
1-
12
#419140000000
0!
0%
b101 *
0-
02
b101 6
#419150000000
1!
1%
1-
12
#419160000000
0!
0%
b110 *
0-
02
b110 6
#419170000000
1!
1%
1-
12
#419180000000
0!
0%
b111 *
0-
02
b111 6
#419190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#419200000000
0!
0%
b0 *
0-
02
b0 6
#419210000000
1!
1%
1-
12
#419220000000
0!
0%
b1 *
0-
02
b1 6
#419230000000
1!
1%
1-
12
#419240000000
0!
0%
b10 *
0-
02
b10 6
#419250000000
1!
1%
1-
12
#419260000000
0!
0%
b11 *
0-
02
b11 6
#419270000000
1!
1%
1-
12
15
#419280000000
0!
0%
b100 *
0-
02
b100 6
#419290000000
1!
1%
1-
12
#419300000000
0!
0%
b101 *
0-
02
b101 6
#419310000000
1!
1%
1-
12
#419320000000
0!
0%
b110 *
0-
02
b110 6
#419330000000
1!
1%
1-
12
#419340000000
0!
0%
b111 *
0-
02
b111 6
#419350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#419360000000
0!
0%
b0 *
0-
02
b0 6
#419370000000
1!
1%
1-
12
#419380000000
0!
0%
b1 *
0-
02
b1 6
#419390000000
1!
1%
1-
12
#419400000000
0!
0%
b10 *
0-
02
b10 6
#419410000000
1!
1%
1-
12
#419420000000
0!
0%
b11 *
0-
02
b11 6
#419430000000
1!
1%
1-
12
15
#419440000000
0!
0%
b100 *
0-
02
b100 6
#419450000000
1!
1%
1-
12
#419460000000
0!
0%
b101 *
0-
02
b101 6
#419470000000
1!
1%
1-
12
#419480000000
0!
0%
b110 *
0-
02
b110 6
#419490000000
1!
1%
1-
12
#419500000000
0!
0%
b111 *
0-
02
b111 6
#419510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#419520000000
0!
0%
b0 *
0-
02
b0 6
#419530000000
1!
1%
1-
12
#419540000000
0!
0%
b1 *
0-
02
b1 6
#419550000000
1!
1%
1-
12
#419560000000
0!
0%
b10 *
0-
02
b10 6
#419570000000
1!
1%
1-
12
#419580000000
0!
0%
b11 *
0-
02
b11 6
#419590000000
1!
1%
1-
12
15
#419600000000
0!
0%
b100 *
0-
02
b100 6
#419610000000
1!
1%
1-
12
#419620000000
0!
0%
b101 *
0-
02
b101 6
#419630000000
1!
1%
1-
12
#419640000000
0!
0%
b110 *
0-
02
b110 6
#419650000000
1!
1%
1-
12
#419660000000
0!
0%
b111 *
0-
02
b111 6
#419670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#419680000000
0!
0%
b0 *
0-
02
b0 6
#419690000000
1!
1%
1-
12
#419700000000
0!
0%
b1 *
0-
02
b1 6
#419710000000
1!
1%
1-
12
#419720000000
0!
0%
b10 *
0-
02
b10 6
#419730000000
1!
1%
1-
12
#419740000000
0!
0%
b11 *
0-
02
b11 6
#419750000000
1!
1%
1-
12
15
#419760000000
0!
0%
b100 *
0-
02
b100 6
#419770000000
1!
1%
1-
12
#419780000000
0!
0%
b101 *
0-
02
b101 6
#419790000000
1!
1%
1-
12
#419800000000
0!
0%
b110 *
0-
02
b110 6
#419810000000
1!
1%
1-
12
#419820000000
0!
0%
b111 *
0-
02
b111 6
#419830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#419840000000
0!
0%
b0 *
0-
02
b0 6
#419850000000
1!
1%
1-
12
#419860000000
0!
0%
b1 *
0-
02
b1 6
#419870000000
1!
1%
1-
12
#419880000000
0!
0%
b10 *
0-
02
b10 6
#419890000000
1!
1%
1-
12
#419900000000
0!
0%
b11 *
0-
02
b11 6
#419910000000
1!
1%
1-
12
15
#419920000000
0!
0%
b100 *
0-
02
b100 6
#419930000000
1!
1%
1-
12
#419940000000
0!
0%
b101 *
0-
02
b101 6
#419950000000
1!
1%
1-
12
#419960000000
0!
0%
b110 *
0-
02
b110 6
#419970000000
1!
1%
1-
12
#419980000000
0!
0%
b111 *
0-
02
b111 6
#419990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#420000000000
0!
0%
b0 *
0-
02
b0 6
#420010000000
1!
1%
1-
12
#420020000000
0!
0%
b1 *
0-
02
b1 6
#420030000000
1!
1%
1-
12
#420040000000
0!
0%
b10 *
0-
02
b10 6
#420050000000
1!
1%
1-
12
#420060000000
0!
0%
b11 *
0-
02
b11 6
#420070000000
1!
1%
1-
12
15
#420080000000
0!
0%
b100 *
0-
02
b100 6
#420090000000
1!
1%
1-
12
#420100000000
0!
0%
b101 *
0-
02
b101 6
#420110000000
1!
1%
1-
12
#420120000000
0!
0%
b110 *
0-
02
b110 6
#420130000000
1!
1%
1-
12
#420140000000
0!
0%
b111 *
0-
02
b111 6
#420150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#420160000000
0!
0%
b0 *
0-
02
b0 6
#420170000000
1!
1%
1-
12
#420180000000
0!
0%
b1 *
0-
02
b1 6
#420190000000
1!
1%
1-
12
#420200000000
0!
0%
b10 *
0-
02
b10 6
#420210000000
1!
1%
1-
12
#420220000000
0!
0%
b11 *
0-
02
b11 6
#420230000000
1!
1%
1-
12
15
#420240000000
0!
0%
b100 *
0-
02
b100 6
#420250000000
1!
1%
1-
12
#420260000000
0!
0%
b101 *
0-
02
b101 6
#420270000000
1!
1%
1-
12
#420280000000
0!
0%
b110 *
0-
02
b110 6
#420290000000
1!
1%
1-
12
#420300000000
0!
0%
b111 *
0-
02
b111 6
#420310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#420320000000
0!
0%
b0 *
0-
02
b0 6
#420330000000
1!
1%
1-
12
#420340000000
0!
0%
b1 *
0-
02
b1 6
#420350000000
1!
1%
1-
12
#420360000000
0!
0%
b10 *
0-
02
b10 6
#420370000000
1!
1%
1-
12
#420380000000
0!
0%
b11 *
0-
02
b11 6
#420390000000
1!
1%
1-
12
15
#420400000000
0!
0%
b100 *
0-
02
b100 6
#420410000000
1!
1%
1-
12
#420420000000
0!
0%
b101 *
0-
02
b101 6
#420430000000
1!
1%
1-
12
#420440000000
0!
0%
b110 *
0-
02
b110 6
#420450000000
1!
1%
1-
12
#420460000000
0!
0%
b111 *
0-
02
b111 6
#420470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#420480000000
0!
0%
b0 *
0-
02
b0 6
#420490000000
1!
1%
1-
12
#420500000000
0!
0%
b1 *
0-
02
b1 6
#420510000000
1!
1%
1-
12
#420520000000
0!
0%
b10 *
0-
02
b10 6
#420530000000
1!
1%
1-
12
#420540000000
0!
0%
b11 *
0-
02
b11 6
#420550000000
1!
1%
1-
12
15
#420560000000
0!
0%
b100 *
0-
02
b100 6
#420570000000
1!
1%
1-
12
#420580000000
0!
0%
b101 *
0-
02
b101 6
#420590000000
1!
1%
1-
12
#420600000000
0!
0%
b110 *
0-
02
b110 6
#420610000000
1!
1%
1-
12
#420620000000
0!
0%
b111 *
0-
02
b111 6
#420630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#420640000000
0!
0%
b0 *
0-
02
b0 6
#420650000000
1!
1%
1-
12
#420660000000
0!
0%
b1 *
0-
02
b1 6
#420670000000
1!
1%
1-
12
#420680000000
0!
0%
b10 *
0-
02
b10 6
#420690000000
1!
1%
1-
12
#420700000000
0!
0%
b11 *
0-
02
b11 6
#420710000000
1!
1%
1-
12
15
#420720000000
0!
0%
b100 *
0-
02
b100 6
#420730000000
1!
1%
1-
12
#420740000000
0!
0%
b101 *
0-
02
b101 6
#420750000000
1!
1%
1-
12
#420760000000
0!
0%
b110 *
0-
02
b110 6
#420770000000
1!
1%
1-
12
#420780000000
0!
0%
b111 *
0-
02
b111 6
#420790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#420800000000
0!
0%
b0 *
0-
02
b0 6
#420810000000
1!
1%
1-
12
#420820000000
0!
0%
b1 *
0-
02
b1 6
#420830000000
1!
1%
1-
12
#420840000000
0!
0%
b10 *
0-
02
b10 6
#420850000000
1!
1%
1-
12
#420860000000
0!
0%
b11 *
0-
02
b11 6
#420870000000
1!
1%
1-
12
15
#420880000000
0!
0%
b100 *
0-
02
b100 6
#420890000000
1!
1%
1-
12
#420900000000
0!
0%
b101 *
0-
02
b101 6
#420910000000
1!
1%
1-
12
#420920000000
0!
0%
b110 *
0-
02
b110 6
#420930000000
1!
1%
1-
12
#420940000000
0!
0%
b111 *
0-
02
b111 6
#420950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#420960000000
0!
0%
b0 *
0-
02
b0 6
#420970000000
1!
1%
1-
12
#420980000000
0!
0%
b1 *
0-
02
b1 6
#420990000000
1!
1%
1-
12
#421000000000
0!
0%
b10 *
0-
02
b10 6
#421010000000
1!
1%
1-
12
#421020000000
0!
0%
b11 *
0-
02
b11 6
#421030000000
1!
1%
1-
12
15
#421040000000
0!
0%
b100 *
0-
02
b100 6
#421050000000
1!
1%
1-
12
#421060000000
0!
0%
b101 *
0-
02
b101 6
#421070000000
1!
1%
1-
12
#421080000000
0!
0%
b110 *
0-
02
b110 6
#421090000000
1!
1%
1-
12
#421100000000
0!
0%
b111 *
0-
02
b111 6
#421110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#421120000000
0!
0%
b0 *
0-
02
b0 6
#421130000000
1!
1%
1-
12
#421140000000
0!
0%
b1 *
0-
02
b1 6
#421150000000
1!
1%
1-
12
#421160000000
0!
0%
b10 *
0-
02
b10 6
#421170000000
1!
1%
1-
12
#421180000000
0!
0%
b11 *
0-
02
b11 6
#421190000000
1!
1%
1-
12
15
#421200000000
0!
0%
b100 *
0-
02
b100 6
#421210000000
1!
1%
1-
12
#421220000000
0!
0%
b101 *
0-
02
b101 6
#421230000000
1!
1%
1-
12
#421240000000
0!
0%
b110 *
0-
02
b110 6
#421250000000
1!
1%
1-
12
#421260000000
0!
0%
b111 *
0-
02
b111 6
#421270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#421280000000
0!
0%
b0 *
0-
02
b0 6
#421290000000
1!
1%
1-
12
#421300000000
0!
0%
b1 *
0-
02
b1 6
#421310000000
1!
1%
1-
12
#421320000000
0!
0%
b10 *
0-
02
b10 6
#421330000000
1!
1%
1-
12
#421340000000
0!
0%
b11 *
0-
02
b11 6
#421350000000
1!
1%
1-
12
15
#421360000000
0!
0%
b100 *
0-
02
b100 6
#421370000000
1!
1%
1-
12
#421380000000
0!
0%
b101 *
0-
02
b101 6
#421390000000
1!
1%
1-
12
#421400000000
0!
0%
b110 *
0-
02
b110 6
#421410000000
1!
1%
1-
12
#421420000000
0!
0%
b111 *
0-
02
b111 6
#421430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#421440000000
0!
0%
b0 *
0-
02
b0 6
#421450000000
1!
1%
1-
12
#421460000000
0!
0%
b1 *
0-
02
b1 6
#421470000000
1!
1%
1-
12
#421480000000
0!
0%
b10 *
0-
02
b10 6
#421490000000
1!
1%
1-
12
#421500000000
0!
0%
b11 *
0-
02
b11 6
#421510000000
1!
1%
1-
12
15
#421520000000
0!
0%
b100 *
0-
02
b100 6
#421530000000
1!
1%
1-
12
#421540000000
0!
0%
b101 *
0-
02
b101 6
#421550000000
1!
1%
1-
12
#421560000000
0!
0%
b110 *
0-
02
b110 6
#421570000000
1!
1%
1-
12
#421580000000
0!
0%
b111 *
0-
02
b111 6
#421590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#421600000000
0!
0%
b0 *
0-
02
b0 6
#421610000000
1!
1%
1-
12
#421620000000
0!
0%
b1 *
0-
02
b1 6
#421630000000
1!
1%
1-
12
#421640000000
0!
0%
b10 *
0-
02
b10 6
#421650000000
1!
1%
1-
12
#421660000000
0!
0%
b11 *
0-
02
b11 6
#421670000000
1!
1%
1-
12
15
#421680000000
0!
0%
b100 *
0-
02
b100 6
#421690000000
1!
1%
1-
12
#421700000000
0!
0%
b101 *
0-
02
b101 6
#421710000000
1!
1%
1-
12
#421720000000
0!
0%
b110 *
0-
02
b110 6
#421730000000
1!
1%
1-
12
#421740000000
0!
0%
b111 *
0-
02
b111 6
#421750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#421760000000
0!
0%
b0 *
0-
02
b0 6
#421770000000
1!
1%
1-
12
#421780000000
0!
0%
b1 *
0-
02
b1 6
#421790000000
1!
1%
1-
12
#421800000000
0!
0%
b10 *
0-
02
b10 6
#421810000000
1!
1%
1-
12
#421820000000
0!
0%
b11 *
0-
02
b11 6
#421830000000
1!
1%
1-
12
15
#421840000000
0!
0%
b100 *
0-
02
b100 6
#421850000000
1!
1%
1-
12
#421860000000
0!
0%
b101 *
0-
02
b101 6
#421870000000
1!
1%
1-
12
#421880000000
0!
0%
b110 *
0-
02
b110 6
#421890000000
1!
1%
1-
12
#421900000000
0!
0%
b111 *
0-
02
b111 6
#421910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#421920000000
0!
0%
b0 *
0-
02
b0 6
#421930000000
1!
1%
1-
12
#421940000000
0!
0%
b1 *
0-
02
b1 6
#421950000000
1!
1%
1-
12
#421960000000
0!
0%
b10 *
0-
02
b10 6
#421970000000
1!
1%
1-
12
#421980000000
0!
0%
b11 *
0-
02
b11 6
#421990000000
1!
1%
1-
12
15
#422000000000
0!
0%
b100 *
0-
02
b100 6
#422010000000
1!
1%
1-
12
#422020000000
0!
0%
b101 *
0-
02
b101 6
#422030000000
1!
1%
1-
12
#422040000000
0!
0%
b110 *
0-
02
b110 6
#422050000000
1!
1%
1-
12
#422060000000
0!
0%
b111 *
0-
02
b111 6
#422070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#422080000000
0!
0%
b0 *
0-
02
b0 6
#422090000000
1!
1%
1-
12
#422100000000
0!
0%
b1 *
0-
02
b1 6
#422110000000
1!
1%
1-
12
#422120000000
0!
0%
b10 *
0-
02
b10 6
#422130000000
1!
1%
1-
12
#422140000000
0!
0%
b11 *
0-
02
b11 6
#422150000000
1!
1%
1-
12
15
#422160000000
0!
0%
b100 *
0-
02
b100 6
#422170000000
1!
1%
1-
12
#422180000000
0!
0%
b101 *
0-
02
b101 6
#422190000000
1!
1%
1-
12
#422200000000
0!
0%
b110 *
0-
02
b110 6
#422210000000
1!
1%
1-
12
#422220000000
0!
0%
b111 *
0-
02
b111 6
#422230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#422240000000
0!
0%
b0 *
0-
02
b0 6
#422250000000
1!
1%
1-
12
#422260000000
0!
0%
b1 *
0-
02
b1 6
#422270000000
1!
1%
1-
12
#422280000000
0!
0%
b10 *
0-
02
b10 6
#422290000000
1!
1%
1-
12
#422300000000
0!
0%
b11 *
0-
02
b11 6
#422310000000
1!
1%
1-
12
15
#422320000000
0!
0%
b100 *
0-
02
b100 6
#422330000000
1!
1%
1-
12
#422340000000
0!
0%
b101 *
0-
02
b101 6
#422350000000
1!
1%
1-
12
#422360000000
0!
0%
b110 *
0-
02
b110 6
#422370000000
1!
1%
1-
12
#422380000000
0!
0%
b111 *
0-
02
b111 6
#422390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#422400000000
0!
0%
b0 *
0-
02
b0 6
#422410000000
1!
1%
1-
12
#422420000000
0!
0%
b1 *
0-
02
b1 6
#422430000000
1!
1%
1-
12
#422440000000
0!
0%
b10 *
0-
02
b10 6
#422450000000
1!
1%
1-
12
#422460000000
0!
0%
b11 *
0-
02
b11 6
#422470000000
1!
1%
1-
12
15
#422480000000
0!
0%
b100 *
0-
02
b100 6
#422490000000
1!
1%
1-
12
#422500000000
0!
0%
b101 *
0-
02
b101 6
#422510000000
1!
1%
1-
12
#422520000000
0!
0%
b110 *
0-
02
b110 6
#422530000000
1!
1%
1-
12
#422540000000
0!
0%
b111 *
0-
02
b111 6
#422550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#422560000000
0!
0%
b0 *
0-
02
b0 6
#422570000000
1!
1%
1-
12
#422580000000
0!
0%
b1 *
0-
02
b1 6
#422590000000
1!
1%
1-
12
#422600000000
0!
0%
b10 *
0-
02
b10 6
#422610000000
1!
1%
1-
12
#422620000000
0!
0%
b11 *
0-
02
b11 6
#422630000000
1!
1%
1-
12
15
#422640000000
0!
0%
b100 *
0-
02
b100 6
#422650000000
1!
1%
1-
12
#422660000000
0!
0%
b101 *
0-
02
b101 6
#422670000000
1!
1%
1-
12
#422680000000
0!
0%
b110 *
0-
02
b110 6
#422690000000
1!
1%
1-
12
#422700000000
0!
0%
b111 *
0-
02
b111 6
#422710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#422720000000
0!
0%
b0 *
0-
02
b0 6
#422730000000
1!
1%
1-
12
#422740000000
0!
0%
b1 *
0-
02
b1 6
#422750000000
1!
1%
1-
12
#422760000000
0!
0%
b10 *
0-
02
b10 6
#422770000000
1!
1%
1-
12
#422780000000
0!
0%
b11 *
0-
02
b11 6
#422790000000
1!
1%
1-
12
15
#422800000000
0!
0%
b100 *
0-
02
b100 6
#422810000000
1!
1%
1-
12
#422820000000
0!
0%
b101 *
0-
02
b101 6
#422830000000
1!
1%
1-
12
#422840000000
0!
0%
b110 *
0-
02
b110 6
#422850000000
1!
1%
1-
12
#422860000000
0!
0%
b111 *
0-
02
b111 6
#422870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#422880000000
0!
0%
b0 *
0-
02
b0 6
#422890000000
1!
1%
1-
12
#422900000000
0!
0%
b1 *
0-
02
b1 6
#422910000000
1!
1%
1-
12
#422920000000
0!
0%
b10 *
0-
02
b10 6
#422930000000
1!
1%
1-
12
#422940000000
0!
0%
b11 *
0-
02
b11 6
#422950000000
1!
1%
1-
12
15
#422960000000
0!
0%
b100 *
0-
02
b100 6
#422970000000
1!
1%
1-
12
#422980000000
0!
0%
b101 *
0-
02
b101 6
#422990000000
1!
1%
1-
12
#423000000000
0!
0%
b110 *
0-
02
b110 6
#423010000000
1!
1%
1-
12
#423020000000
0!
0%
b111 *
0-
02
b111 6
#423030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#423040000000
0!
0%
b0 *
0-
02
b0 6
#423050000000
1!
1%
1-
12
#423060000000
0!
0%
b1 *
0-
02
b1 6
#423070000000
1!
1%
1-
12
#423080000000
0!
0%
b10 *
0-
02
b10 6
#423090000000
1!
1%
1-
12
#423100000000
0!
0%
b11 *
0-
02
b11 6
#423110000000
1!
1%
1-
12
15
#423120000000
0!
0%
b100 *
0-
02
b100 6
#423130000000
1!
1%
1-
12
#423140000000
0!
0%
b101 *
0-
02
b101 6
#423150000000
1!
1%
1-
12
#423160000000
0!
0%
b110 *
0-
02
b110 6
#423170000000
1!
1%
1-
12
#423180000000
0!
0%
b111 *
0-
02
b111 6
#423190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#423200000000
0!
0%
b0 *
0-
02
b0 6
#423210000000
1!
1%
1-
12
#423220000000
0!
0%
b1 *
0-
02
b1 6
#423230000000
1!
1%
1-
12
#423240000000
0!
0%
b10 *
0-
02
b10 6
#423250000000
1!
1%
1-
12
#423260000000
0!
0%
b11 *
0-
02
b11 6
#423270000000
1!
1%
1-
12
15
#423280000000
0!
0%
b100 *
0-
02
b100 6
#423290000000
1!
1%
1-
12
#423300000000
0!
0%
b101 *
0-
02
b101 6
#423310000000
1!
1%
1-
12
#423320000000
0!
0%
b110 *
0-
02
b110 6
#423330000000
1!
1%
1-
12
#423340000000
0!
0%
b111 *
0-
02
b111 6
#423350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#423360000000
0!
0%
b0 *
0-
02
b0 6
#423370000000
1!
1%
1-
12
#423380000000
0!
0%
b1 *
0-
02
b1 6
#423390000000
1!
1%
1-
12
#423400000000
0!
0%
b10 *
0-
02
b10 6
#423410000000
1!
1%
1-
12
#423420000000
0!
0%
b11 *
0-
02
b11 6
#423430000000
1!
1%
1-
12
15
#423440000000
0!
0%
b100 *
0-
02
b100 6
#423450000000
1!
1%
1-
12
#423460000000
0!
0%
b101 *
0-
02
b101 6
#423470000000
1!
1%
1-
12
#423480000000
0!
0%
b110 *
0-
02
b110 6
#423490000000
1!
1%
1-
12
#423500000000
0!
0%
b111 *
0-
02
b111 6
#423510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#423520000000
0!
0%
b0 *
0-
02
b0 6
#423530000000
1!
1%
1-
12
#423540000000
0!
0%
b1 *
0-
02
b1 6
#423550000000
1!
1%
1-
12
#423560000000
0!
0%
b10 *
0-
02
b10 6
#423570000000
1!
1%
1-
12
#423580000000
0!
0%
b11 *
0-
02
b11 6
#423590000000
1!
1%
1-
12
15
#423600000000
0!
0%
b100 *
0-
02
b100 6
#423610000000
1!
1%
1-
12
#423620000000
0!
0%
b101 *
0-
02
b101 6
#423630000000
1!
1%
1-
12
#423640000000
0!
0%
b110 *
0-
02
b110 6
#423650000000
1!
1%
1-
12
#423660000000
0!
0%
b111 *
0-
02
b111 6
#423670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#423680000000
0!
0%
b0 *
0-
02
b0 6
#423690000000
1!
1%
1-
12
#423700000000
0!
0%
b1 *
0-
02
b1 6
#423710000000
1!
1%
1-
12
#423720000000
0!
0%
b10 *
0-
02
b10 6
#423730000000
1!
1%
1-
12
#423740000000
0!
0%
b11 *
0-
02
b11 6
#423750000000
1!
1%
1-
12
15
#423760000000
0!
0%
b100 *
0-
02
b100 6
#423770000000
1!
1%
1-
12
#423780000000
0!
0%
b101 *
0-
02
b101 6
#423790000000
1!
1%
1-
12
#423800000000
0!
0%
b110 *
0-
02
b110 6
#423810000000
1!
1%
1-
12
#423820000000
0!
0%
b111 *
0-
02
b111 6
#423830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#423840000000
0!
0%
b0 *
0-
02
b0 6
#423850000000
1!
1%
1-
12
#423860000000
0!
0%
b1 *
0-
02
b1 6
#423870000000
1!
1%
1-
12
#423880000000
0!
0%
b10 *
0-
02
b10 6
#423890000000
1!
1%
1-
12
#423900000000
0!
0%
b11 *
0-
02
b11 6
#423910000000
1!
1%
1-
12
15
#423920000000
0!
0%
b100 *
0-
02
b100 6
#423930000000
1!
1%
1-
12
#423940000000
0!
0%
b101 *
0-
02
b101 6
#423950000000
1!
1%
1-
12
#423960000000
0!
0%
b110 *
0-
02
b110 6
#423970000000
1!
1%
1-
12
#423980000000
0!
0%
b111 *
0-
02
b111 6
#423990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#424000000000
0!
0%
b0 *
0-
02
b0 6
#424010000000
1!
1%
1-
12
#424020000000
0!
0%
b1 *
0-
02
b1 6
#424030000000
1!
1%
1-
12
#424040000000
0!
0%
b10 *
0-
02
b10 6
#424050000000
1!
1%
1-
12
#424060000000
0!
0%
b11 *
0-
02
b11 6
#424070000000
1!
1%
1-
12
15
#424080000000
0!
0%
b100 *
0-
02
b100 6
#424090000000
1!
1%
1-
12
#424100000000
0!
0%
b101 *
0-
02
b101 6
#424110000000
1!
1%
1-
12
#424120000000
0!
0%
b110 *
0-
02
b110 6
#424130000000
1!
1%
1-
12
#424140000000
0!
0%
b111 *
0-
02
b111 6
#424150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#424160000000
0!
0%
b0 *
0-
02
b0 6
#424170000000
1!
1%
1-
12
#424180000000
0!
0%
b1 *
0-
02
b1 6
#424190000000
1!
1%
1-
12
#424200000000
0!
0%
b10 *
0-
02
b10 6
#424210000000
1!
1%
1-
12
#424220000000
0!
0%
b11 *
0-
02
b11 6
#424230000000
1!
1%
1-
12
15
#424240000000
0!
0%
b100 *
0-
02
b100 6
#424250000000
1!
1%
1-
12
#424260000000
0!
0%
b101 *
0-
02
b101 6
#424270000000
1!
1%
1-
12
#424280000000
0!
0%
b110 *
0-
02
b110 6
#424290000000
1!
1%
1-
12
#424300000000
0!
0%
b111 *
0-
02
b111 6
#424310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#424320000000
0!
0%
b0 *
0-
02
b0 6
#424330000000
1!
1%
1-
12
#424340000000
0!
0%
b1 *
0-
02
b1 6
#424350000000
1!
1%
1-
12
#424360000000
0!
0%
b10 *
0-
02
b10 6
#424370000000
1!
1%
1-
12
#424380000000
0!
0%
b11 *
0-
02
b11 6
#424390000000
1!
1%
1-
12
15
#424400000000
0!
0%
b100 *
0-
02
b100 6
#424410000000
1!
1%
1-
12
#424420000000
0!
0%
b101 *
0-
02
b101 6
#424430000000
1!
1%
1-
12
#424440000000
0!
0%
b110 *
0-
02
b110 6
#424450000000
1!
1%
1-
12
#424460000000
0!
0%
b111 *
0-
02
b111 6
#424470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#424480000000
0!
0%
b0 *
0-
02
b0 6
#424490000000
1!
1%
1-
12
#424500000000
0!
0%
b1 *
0-
02
b1 6
#424510000000
1!
1%
1-
12
#424520000000
0!
0%
b10 *
0-
02
b10 6
#424530000000
1!
1%
1-
12
#424540000000
0!
0%
b11 *
0-
02
b11 6
#424550000000
1!
1%
1-
12
15
#424560000000
0!
0%
b100 *
0-
02
b100 6
#424570000000
1!
1%
1-
12
#424580000000
0!
0%
b101 *
0-
02
b101 6
#424590000000
1!
1%
1-
12
#424600000000
0!
0%
b110 *
0-
02
b110 6
#424610000000
1!
1%
1-
12
#424620000000
0!
0%
b111 *
0-
02
b111 6
#424630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#424640000000
0!
0%
b0 *
0-
02
b0 6
#424650000000
1!
1%
1-
12
#424660000000
0!
0%
b1 *
0-
02
b1 6
#424670000000
1!
1%
1-
12
#424680000000
0!
0%
b10 *
0-
02
b10 6
#424690000000
1!
1%
1-
12
#424700000000
0!
0%
b11 *
0-
02
b11 6
#424710000000
1!
1%
1-
12
15
#424720000000
0!
0%
b100 *
0-
02
b100 6
#424730000000
1!
1%
1-
12
#424740000000
0!
0%
b101 *
0-
02
b101 6
#424750000000
1!
1%
1-
12
#424760000000
0!
0%
b110 *
0-
02
b110 6
#424770000000
1!
1%
1-
12
#424780000000
0!
0%
b111 *
0-
02
b111 6
#424790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#424800000000
0!
0%
b0 *
0-
02
b0 6
#424810000000
1!
1%
1-
12
#424820000000
0!
0%
b1 *
0-
02
b1 6
#424830000000
1!
1%
1-
12
#424840000000
0!
0%
b10 *
0-
02
b10 6
#424850000000
1!
1%
1-
12
#424860000000
0!
0%
b11 *
0-
02
b11 6
#424870000000
1!
1%
1-
12
15
#424880000000
0!
0%
b100 *
0-
02
b100 6
#424890000000
1!
1%
1-
12
#424900000000
0!
0%
b101 *
0-
02
b101 6
#424910000000
1!
1%
1-
12
#424920000000
0!
0%
b110 *
0-
02
b110 6
#424930000000
1!
1%
1-
12
#424940000000
0!
0%
b111 *
0-
02
b111 6
#424950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#424960000000
0!
0%
b0 *
0-
02
b0 6
#424970000000
1!
1%
1-
12
#424980000000
0!
0%
b1 *
0-
02
b1 6
#424990000000
1!
1%
1-
12
#425000000000
0!
0%
b10 *
0-
02
b10 6
#425010000000
1!
1%
1-
12
#425020000000
0!
0%
b11 *
0-
02
b11 6
#425030000000
1!
1%
1-
12
15
#425040000000
0!
0%
b100 *
0-
02
b100 6
#425050000000
1!
1%
1-
12
#425060000000
0!
0%
b101 *
0-
02
b101 6
#425070000000
1!
1%
1-
12
#425080000000
0!
0%
b110 *
0-
02
b110 6
#425090000000
1!
1%
1-
12
#425100000000
0!
0%
b111 *
0-
02
b111 6
#425110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#425120000000
0!
0%
b0 *
0-
02
b0 6
#425130000000
1!
1%
1-
12
#425140000000
0!
0%
b1 *
0-
02
b1 6
#425150000000
1!
1%
1-
12
#425160000000
0!
0%
b10 *
0-
02
b10 6
#425170000000
1!
1%
1-
12
#425180000000
0!
0%
b11 *
0-
02
b11 6
#425190000000
1!
1%
1-
12
15
#425200000000
0!
0%
b100 *
0-
02
b100 6
#425210000000
1!
1%
1-
12
#425220000000
0!
0%
b101 *
0-
02
b101 6
#425230000000
1!
1%
1-
12
#425240000000
0!
0%
b110 *
0-
02
b110 6
#425250000000
1!
1%
1-
12
#425260000000
0!
0%
b111 *
0-
02
b111 6
#425270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#425280000000
0!
0%
b0 *
0-
02
b0 6
#425290000000
1!
1%
1-
12
#425300000000
0!
0%
b1 *
0-
02
b1 6
#425310000000
1!
1%
1-
12
#425320000000
0!
0%
b10 *
0-
02
b10 6
#425330000000
1!
1%
1-
12
#425340000000
0!
0%
b11 *
0-
02
b11 6
#425350000000
1!
1%
1-
12
15
#425360000000
0!
0%
b100 *
0-
02
b100 6
#425370000000
1!
1%
1-
12
#425380000000
0!
0%
b101 *
0-
02
b101 6
#425390000000
1!
1%
1-
12
#425400000000
0!
0%
b110 *
0-
02
b110 6
#425410000000
1!
1%
1-
12
#425420000000
0!
0%
b111 *
0-
02
b111 6
#425430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#425440000000
0!
0%
b0 *
0-
02
b0 6
#425450000000
1!
1%
1-
12
#425460000000
0!
0%
b1 *
0-
02
b1 6
#425470000000
1!
1%
1-
12
#425480000000
0!
0%
b10 *
0-
02
b10 6
#425490000000
1!
1%
1-
12
#425500000000
0!
0%
b11 *
0-
02
b11 6
#425510000000
1!
1%
1-
12
15
#425520000000
0!
0%
b100 *
0-
02
b100 6
#425530000000
1!
1%
1-
12
#425540000000
0!
0%
b101 *
0-
02
b101 6
#425550000000
1!
1%
1-
12
#425560000000
0!
0%
b110 *
0-
02
b110 6
#425570000000
1!
1%
1-
12
#425580000000
0!
0%
b111 *
0-
02
b111 6
#425590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#425600000000
0!
0%
b0 *
0-
02
b0 6
#425610000000
1!
1%
1-
12
#425620000000
0!
0%
b1 *
0-
02
b1 6
#425630000000
1!
1%
1-
12
#425640000000
0!
0%
b10 *
0-
02
b10 6
#425650000000
1!
1%
1-
12
#425660000000
0!
0%
b11 *
0-
02
b11 6
#425670000000
1!
1%
1-
12
15
#425680000000
0!
0%
b100 *
0-
02
b100 6
#425690000000
1!
1%
1-
12
#425700000000
0!
0%
b101 *
0-
02
b101 6
#425710000000
1!
1%
1-
12
#425720000000
0!
0%
b110 *
0-
02
b110 6
#425730000000
1!
1%
1-
12
#425740000000
0!
0%
b111 *
0-
02
b111 6
#425750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#425760000000
0!
0%
b0 *
0-
02
b0 6
#425770000000
1!
1%
1-
12
#425780000000
0!
0%
b1 *
0-
02
b1 6
#425790000000
1!
1%
1-
12
#425800000000
0!
0%
b10 *
0-
02
b10 6
#425810000000
1!
1%
1-
12
#425820000000
0!
0%
b11 *
0-
02
b11 6
#425830000000
1!
1%
1-
12
15
#425840000000
0!
0%
b100 *
0-
02
b100 6
#425850000000
1!
1%
1-
12
#425860000000
0!
0%
b101 *
0-
02
b101 6
#425870000000
1!
1%
1-
12
#425880000000
0!
0%
b110 *
0-
02
b110 6
#425890000000
1!
1%
1-
12
#425900000000
0!
0%
b111 *
0-
02
b111 6
#425910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#425920000000
0!
0%
b0 *
0-
02
b0 6
#425930000000
1!
1%
1-
12
#425940000000
0!
0%
b1 *
0-
02
b1 6
#425950000000
1!
1%
1-
12
#425960000000
0!
0%
b10 *
0-
02
b10 6
#425970000000
1!
1%
1-
12
#425980000000
0!
0%
b11 *
0-
02
b11 6
#425990000000
1!
1%
1-
12
15
#426000000000
0!
0%
b100 *
0-
02
b100 6
#426010000000
1!
1%
1-
12
#426020000000
0!
0%
b101 *
0-
02
b101 6
#426030000000
1!
1%
1-
12
#426040000000
0!
0%
b110 *
0-
02
b110 6
#426050000000
1!
1%
1-
12
#426060000000
0!
0%
b111 *
0-
02
b111 6
#426070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#426080000000
0!
0%
b0 *
0-
02
b0 6
#426090000000
1!
1%
1-
12
#426100000000
0!
0%
b1 *
0-
02
b1 6
#426110000000
1!
1%
1-
12
#426120000000
0!
0%
b10 *
0-
02
b10 6
#426130000000
1!
1%
1-
12
#426140000000
0!
0%
b11 *
0-
02
b11 6
#426150000000
1!
1%
1-
12
15
#426160000000
0!
0%
b100 *
0-
02
b100 6
#426170000000
1!
1%
1-
12
#426180000000
0!
0%
b101 *
0-
02
b101 6
#426190000000
1!
1%
1-
12
#426200000000
0!
0%
b110 *
0-
02
b110 6
#426210000000
1!
1%
1-
12
#426220000000
0!
0%
b111 *
0-
02
b111 6
#426230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#426240000000
0!
0%
b0 *
0-
02
b0 6
#426250000000
1!
1%
1-
12
#426260000000
0!
0%
b1 *
0-
02
b1 6
#426270000000
1!
1%
1-
12
#426280000000
0!
0%
b10 *
0-
02
b10 6
#426290000000
1!
1%
1-
12
#426300000000
0!
0%
b11 *
0-
02
b11 6
#426310000000
1!
1%
1-
12
15
#426320000000
0!
0%
b100 *
0-
02
b100 6
#426330000000
1!
1%
1-
12
#426340000000
0!
0%
b101 *
0-
02
b101 6
#426350000000
1!
1%
1-
12
#426360000000
0!
0%
b110 *
0-
02
b110 6
#426370000000
1!
1%
1-
12
#426380000000
0!
0%
b111 *
0-
02
b111 6
#426390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#426400000000
0!
0%
b0 *
0-
02
b0 6
#426410000000
1!
1%
1-
12
#426420000000
0!
0%
b1 *
0-
02
b1 6
#426430000000
1!
1%
1-
12
#426440000000
0!
0%
b10 *
0-
02
b10 6
#426450000000
1!
1%
1-
12
#426460000000
0!
0%
b11 *
0-
02
b11 6
#426470000000
1!
1%
1-
12
15
#426480000000
0!
0%
b100 *
0-
02
b100 6
#426490000000
1!
1%
1-
12
#426500000000
0!
0%
b101 *
0-
02
b101 6
#426510000000
1!
1%
1-
12
#426520000000
0!
0%
b110 *
0-
02
b110 6
#426530000000
1!
1%
1-
12
#426540000000
0!
0%
b111 *
0-
02
b111 6
#426550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#426560000000
0!
0%
b0 *
0-
02
b0 6
#426570000000
1!
1%
1-
12
#426580000000
0!
0%
b1 *
0-
02
b1 6
#426590000000
1!
1%
1-
12
#426600000000
0!
0%
b10 *
0-
02
b10 6
#426610000000
1!
1%
1-
12
#426620000000
0!
0%
b11 *
0-
02
b11 6
#426630000000
1!
1%
1-
12
15
#426640000000
0!
0%
b100 *
0-
02
b100 6
#426650000000
1!
1%
1-
12
#426660000000
0!
0%
b101 *
0-
02
b101 6
#426670000000
1!
1%
1-
12
#426680000000
0!
0%
b110 *
0-
02
b110 6
#426690000000
1!
1%
1-
12
#426700000000
0!
0%
b111 *
0-
02
b111 6
#426710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#426720000000
0!
0%
b0 *
0-
02
b0 6
#426730000000
1!
1%
1-
12
#426740000000
0!
0%
b1 *
0-
02
b1 6
#426750000000
1!
1%
1-
12
#426760000000
0!
0%
b10 *
0-
02
b10 6
#426770000000
1!
1%
1-
12
#426780000000
0!
0%
b11 *
0-
02
b11 6
#426790000000
1!
1%
1-
12
15
#426800000000
0!
0%
b100 *
0-
02
b100 6
#426810000000
1!
1%
1-
12
#426820000000
0!
0%
b101 *
0-
02
b101 6
#426830000000
1!
1%
1-
12
#426840000000
0!
0%
b110 *
0-
02
b110 6
#426850000000
1!
1%
1-
12
#426860000000
0!
0%
b111 *
0-
02
b111 6
#426870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#426880000000
0!
0%
b0 *
0-
02
b0 6
#426890000000
1!
1%
1-
12
#426900000000
0!
0%
b1 *
0-
02
b1 6
#426910000000
1!
1%
1-
12
#426920000000
0!
0%
b10 *
0-
02
b10 6
#426930000000
1!
1%
1-
12
#426940000000
0!
0%
b11 *
0-
02
b11 6
#426950000000
1!
1%
1-
12
15
#426960000000
0!
0%
b100 *
0-
02
b100 6
#426970000000
1!
1%
1-
12
#426980000000
0!
0%
b101 *
0-
02
b101 6
#426990000000
1!
1%
1-
12
#427000000000
0!
0%
b110 *
0-
02
b110 6
#427010000000
1!
1%
1-
12
#427020000000
0!
0%
b111 *
0-
02
b111 6
#427030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#427040000000
0!
0%
b0 *
0-
02
b0 6
#427050000000
1!
1%
1-
12
#427060000000
0!
0%
b1 *
0-
02
b1 6
#427070000000
1!
1%
1-
12
#427080000000
0!
0%
b10 *
0-
02
b10 6
#427090000000
1!
1%
1-
12
#427100000000
0!
0%
b11 *
0-
02
b11 6
#427110000000
1!
1%
1-
12
15
#427120000000
0!
0%
b100 *
0-
02
b100 6
#427130000000
1!
1%
1-
12
#427140000000
0!
0%
b101 *
0-
02
b101 6
#427150000000
1!
1%
1-
12
#427160000000
0!
0%
b110 *
0-
02
b110 6
#427170000000
1!
1%
1-
12
#427180000000
0!
0%
b111 *
0-
02
b111 6
#427190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#427200000000
0!
0%
b0 *
0-
02
b0 6
#427210000000
1!
1%
1-
12
#427220000000
0!
0%
b1 *
0-
02
b1 6
#427230000000
1!
1%
1-
12
#427240000000
0!
0%
b10 *
0-
02
b10 6
#427250000000
1!
1%
1-
12
#427260000000
0!
0%
b11 *
0-
02
b11 6
#427270000000
1!
1%
1-
12
15
#427280000000
0!
0%
b100 *
0-
02
b100 6
#427290000000
1!
1%
1-
12
#427300000000
0!
0%
b101 *
0-
02
b101 6
#427310000000
1!
1%
1-
12
#427320000000
0!
0%
b110 *
0-
02
b110 6
#427330000000
1!
1%
1-
12
#427340000000
0!
0%
b111 *
0-
02
b111 6
#427350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#427360000000
0!
0%
b0 *
0-
02
b0 6
#427370000000
1!
1%
1-
12
#427380000000
0!
0%
b1 *
0-
02
b1 6
#427390000000
1!
1%
1-
12
#427400000000
0!
0%
b10 *
0-
02
b10 6
#427410000000
1!
1%
1-
12
#427420000000
0!
0%
b11 *
0-
02
b11 6
#427430000000
1!
1%
1-
12
15
#427440000000
0!
0%
b100 *
0-
02
b100 6
#427450000000
1!
1%
1-
12
#427460000000
0!
0%
b101 *
0-
02
b101 6
#427470000000
1!
1%
1-
12
#427480000000
0!
0%
b110 *
0-
02
b110 6
#427490000000
1!
1%
1-
12
#427500000000
0!
0%
b111 *
0-
02
b111 6
#427510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#427520000000
0!
0%
b0 *
0-
02
b0 6
#427530000000
1!
1%
1-
12
#427540000000
0!
0%
b1 *
0-
02
b1 6
#427550000000
1!
1%
1-
12
#427560000000
0!
0%
b10 *
0-
02
b10 6
#427570000000
1!
1%
1-
12
#427580000000
0!
0%
b11 *
0-
02
b11 6
#427590000000
1!
1%
1-
12
15
#427600000000
0!
0%
b100 *
0-
02
b100 6
#427610000000
1!
1%
1-
12
#427620000000
0!
0%
b101 *
0-
02
b101 6
#427630000000
1!
1%
1-
12
#427640000000
0!
0%
b110 *
0-
02
b110 6
#427650000000
1!
1%
1-
12
#427660000000
0!
0%
b111 *
0-
02
b111 6
#427670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#427680000000
0!
0%
b0 *
0-
02
b0 6
#427690000000
1!
1%
1-
12
#427700000000
0!
0%
b1 *
0-
02
b1 6
#427710000000
1!
1%
1-
12
#427720000000
0!
0%
b10 *
0-
02
b10 6
#427730000000
1!
1%
1-
12
#427740000000
0!
0%
b11 *
0-
02
b11 6
#427750000000
1!
1%
1-
12
15
#427760000000
0!
0%
b100 *
0-
02
b100 6
#427770000000
1!
1%
1-
12
#427780000000
0!
0%
b101 *
0-
02
b101 6
#427790000000
1!
1%
1-
12
#427800000000
0!
0%
b110 *
0-
02
b110 6
#427810000000
1!
1%
1-
12
#427820000000
0!
0%
b111 *
0-
02
b111 6
#427830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#427840000000
0!
0%
b0 *
0-
02
b0 6
#427850000000
1!
1%
1-
12
#427860000000
0!
0%
b1 *
0-
02
b1 6
#427870000000
1!
1%
1-
12
#427880000000
0!
0%
b10 *
0-
02
b10 6
#427890000000
1!
1%
1-
12
#427900000000
0!
0%
b11 *
0-
02
b11 6
#427910000000
1!
1%
1-
12
15
#427920000000
0!
0%
b100 *
0-
02
b100 6
#427930000000
1!
1%
1-
12
#427940000000
0!
0%
b101 *
0-
02
b101 6
#427950000000
1!
1%
1-
12
#427960000000
0!
0%
b110 *
0-
02
b110 6
#427970000000
1!
1%
1-
12
#427980000000
0!
0%
b111 *
0-
02
b111 6
#427990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#428000000000
0!
0%
b0 *
0-
02
b0 6
#428010000000
1!
1%
1-
12
#428020000000
0!
0%
b1 *
0-
02
b1 6
#428030000000
1!
1%
1-
12
#428040000000
0!
0%
b10 *
0-
02
b10 6
#428050000000
1!
1%
1-
12
#428060000000
0!
0%
b11 *
0-
02
b11 6
#428070000000
1!
1%
1-
12
15
#428080000000
0!
0%
b100 *
0-
02
b100 6
#428090000000
1!
1%
1-
12
#428100000000
0!
0%
b101 *
0-
02
b101 6
#428110000000
1!
1%
1-
12
#428120000000
0!
0%
b110 *
0-
02
b110 6
#428130000000
1!
1%
1-
12
#428140000000
0!
0%
b111 *
0-
02
b111 6
#428150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#428160000000
0!
0%
b0 *
0-
02
b0 6
#428170000000
1!
1%
1-
12
#428180000000
0!
0%
b1 *
0-
02
b1 6
#428190000000
1!
1%
1-
12
#428200000000
0!
0%
b10 *
0-
02
b10 6
#428210000000
1!
1%
1-
12
#428220000000
0!
0%
b11 *
0-
02
b11 6
#428230000000
1!
1%
1-
12
15
#428240000000
0!
0%
b100 *
0-
02
b100 6
#428250000000
1!
1%
1-
12
#428260000000
0!
0%
b101 *
0-
02
b101 6
#428270000000
1!
1%
1-
12
#428280000000
0!
0%
b110 *
0-
02
b110 6
#428290000000
1!
1%
1-
12
#428300000000
0!
0%
b111 *
0-
02
b111 6
#428310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#428320000000
0!
0%
b0 *
0-
02
b0 6
#428330000000
1!
1%
1-
12
#428340000000
0!
0%
b1 *
0-
02
b1 6
#428350000000
1!
1%
1-
12
#428360000000
0!
0%
b10 *
0-
02
b10 6
#428370000000
1!
1%
1-
12
#428380000000
0!
0%
b11 *
0-
02
b11 6
#428390000000
1!
1%
1-
12
15
#428400000000
0!
0%
b100 *
0-
02
b100 6
#428410000000
1!
1%
1-
12
#428420000000
0!
0%
b101 *
0-
02
b101 6
#428430000000
1!
1%
1-
12
#428440000000
0!
0%
b110 *
0-
02
b110 6
#428450000000
1!
1%
1-
12
#428460000000
0!
0%
b111 *
0-
02
b111 6
#428470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#428480000000
0!
0%
b0 *
0-
02
b0 6
#428490000000
1!
1%
1-
12
#428500000000
0!
0%
b1 *
0-
02
b1 6
#428510000000
1!
1%
1-
12
#428520000000
0!
0%
b10 *
0-
02
b10 6
#428530000000
1!
1%
1-
12
#428540000000
0!
0%
b11 *
0-
02
b11 6
#428550000000
1!
1%
1-
12
15
#428560000000
0!
0%
b100 *
0-
02
b100 6
#428570000000
1!
1%
1-
12
#428580000000
0!
0%
b101 *
0-
02
b101 6
#428590000000
1!
1%
1-
12
#428600000000
0!
0%
b110 *
0-
02
b110 6
#428610000000
1!
1%
1-
12
#428620000000
0!
0%
b111 *
0-
02
b111 6
#428630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#428640000000
0!
0%
b0 *
0-
02
b0 6
#428650000000
1!
1%
1-
12
#428660000000
0!
0%
b1 *
0-
02
b1 6
#428670000000
1!
1%
1-
12
#428680000000
0!
0%
b10 *
0-
02
b10 6
#428690000000
1!
1%
1-
12
#428700000000
0!
0%
b11 *
0-
02
b11 6
#428710000000
1!
1%
1-
12
15
#428720000000
0!
0%
b100 *
0-
02
b100 6
#428730000000
1!
1%
1-
12
#428740000000
0!
0%
b101 *
0-
02
b101 6
#428750000000
1!
1%
1-
12
#428760000000
0!
0%
b110 *
0-
02
b110 6
#428770000000
1!
1%
1-
12
#428780000000
0!
0%
b111 *
0-
02
b111 6
#428790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#428800000000
0!
0%
b0 *
0-
02
b0 6
#428810000000
1!
1%
1-
12
#428820000000
0!
0%
b1 *
0-
02
b1 6
#428830000000
1!
1%
1-
12
#428840000000
0!
0%
b10 *
0-
02
b10 6
#428850000000
1!
1%
1-
12
#428860000000
0!
0%
b11 *
0-
02
b11 6
#428870000000
1!
1%
1-
12
15
#428880000000
0!
0%
b100 *
0-
02
b100 6
#428890000000
1!
1%
1-
12
#428900000000
0!
0%
b101 *
0-
02
b101 6
#428910000000
1!
1%
1-
12
#428920000000
0!
0%
b110 *
0-
02
b110 6
#428930000000
1!
1%
1-
12
#428940000000
0!
0%
b111 *
0-
02
b111 6
#428950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#428960000000
0!
0%
b0 *
0-
02
b0 6
#428970000000
1!
1%
1-
12
#428980000000
0!
0%
b1 *
0-
02
b1 6
#428990000000
1!
1%
1-
12
#429000000000
0!
0%
b10 *
0-
02
b10 6
#429010000000
1!
1%
1-
12
#429020000000
0!
0%
b11 *
0-
02
b11 6
#429030000000
1!
1%
1-
12
15
#429040000000
0!
0%
b100 *
0-
02
b100 6
#429050000000
1!
1%
1-
12
#429060000000
0!
0%
b101 *
0-
02
b101 6
#429070000000
1!
1%
1-
12
#429080000000
0!
0%
b110 *
0-
02
b110 6
#429090000000
1!
1%
1-
12
#429100000000
0!
0%
b111 *
0-
02
b111 6
#429110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#429120000000
0!
0%
b0 *
0-
02
b0 6
#429130000000
1!
1%
1-
12
#429140000000
0!
0%
b1 *
0-
02
b1 6
#429150000000
1!
1%
1-
12
#429160000000
0!
0%
b10 *
0-
02
b10 6
#429170000000
1!
1%
1-
12
#429180000000
0!
0%
b11 *
0-
02
b11 6
#429190000000
1!
1%
1-
12
15
#429200000000
0!
0%
b100 *
0-
02
b100 6
#429210000000
1!
1%
1-
12
#429220000000
0!
0%
b101 *
0-
02
b101 6
#429230000000
1!
1%
1-
12
#429240000000
0!
0%
b110 *
0-
02
b110 6
#429250000000
1!
1%
1-
12
#429260000000
0!
0%
b111 *
0-
02
b111 6
#429270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#429280000000
0!
0%
b0 *
0-
02
b0 6
#429290000000
1!
1%
1-
12
#429300000000
0!
0%
b1 *
0-
02
b1 6
#429310000000
1!
1%
1-
12
#429320000000
0!
0%
b10 *
0-
02
b10 6
#429330000000
1!
1%
1-
12
#429340000000
0!
0%
b11 *
0-
02
b11 6
#429350000000
1!
1%
1-
12
15
#429360000000
0!
0%
b100 *
0-
02
b100 6
#429370000000
1!
1%
1-
12
#429380000000
0!
0%
b101 *
0-
02
b101 6
#429390000000
1!
1%
1-
12
#429400000000
0!
0%
b110 *
0-
02
b110 6
#429410000000
1!
1%
1-
12
#429420000000
0!
0%
b111 *
0-
02
b111 6
#429430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#429440000000
0!
0%
b0 *
0-
02
b0 6
#429450000000
1!
1%
1-
12
#429460000000
0!
0%
b1 *
0-
02
b1 6
#429470000000
1!
1%
1-
12
#429480000000
0!
0%
b10 *
0-
02
b10 6
#429490000000
1!
1%
1-
12
#429500000000
0!
0%
b11 *
0-
02
b11 6
#429510000000
1!
1%
1-
12
15
#429520000000
0!
0%
b100 *
0-
02
b100 6
#429530000000
1!
1%
1-
12
#429540000000
0!
0%
b101 *
0-
02
b101 6
#429550000000
1!
1%
1-
12
#429560000000
0!
0%
b110 *
0-
02
b110 6
#429570000000
1!
1%
1-
12
#429580000000
0!
0%
b111 *
0-
02
b111 6
#429590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#429600000000
0!
0%
b0 *
0-
02
b0 6
#429610000000
1!
1%
1-
12
#429620000000
0!
0%
b1 *
0-
02
b1 6
#429630000000
1!
1%
1-
12
#429640000000
0!
0%
b10 *
0-
02
b10 6
#429650000000
1!
1%
1-
12
#429660000000
0!
0%
b11 *
0-
02
b11 6
#429670000000
1!
1%
1-
12
15
#429680000000
0!
0%
b100 *
0-
02
b100 6
#429690000000
1!
1%
1-
12
#429700000000
0!
0%
b101 *
0-
02
b101 6
#429710000000
1!
1%
1-
12
#429720000000
0!
0%
b110 *
0-
02
b110 6
#429730000000
1!
1%
1-
12
#429740000000
0!
0%
b111 *
0-
02
b111 6
#429750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#429760000000
0!
0%
b0 *
0-
02
b0 6
#429770000000
1!
1%
1-
12
#429780000000
0!
0%
b1 *
0-
02
b1 6
#429790000000
1!
1%
1-
12
#429800000000
0!
0%
b10 *
0-
02
b10 6
#429810000000
1!
1%
1-
12
#429820000000
0!
0%
b11 *
0-
02
b11 6
#429830000000
1!
1%
1-
12
15
#429840000000
0!
0%
b100 *
0-
02
b100 6
#429850000000
1!
1%
1-
12
#429860000000
0!
0%
b101 *
0-
02
b101 6
#429870000000
1!
1%
1-
12
#429880000000
0!
0%
b110 *
0-
02
b110 6
#429890000000
1!
1%
1-
12
#429900000000
0!
0%
b111 *
0-
02
b111 6
#429910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#429920000000
0!
0%
b0 *
0-
02
b0 6
#429930000000
1!
1%
1-
12
#429940000000
0!
0%
b1 *
0-
02
b1 6
#429950000000
1!
1%
1-
12
#429960000000
0!
0%
b10 *
0-
02
b10 6
#429970000000
1!
1%
1-
12
#429980000000
0!
0%
b11 *
0-
02
b11 6
#429990000000
1!
1%
1-
12
15
#430000000000
0!
0%
b100 *
0-
02
b100 6
#430010000000
1!
1%
1-
12
#430020000000
0!
0%
b101 *
0-
02
b101 6
#430030000000
1!
1%
1-
12
#430040000000
0!
0%
b110 *
0-
02
b110 6
#430050000000
1!
1%
1-
12
#430060000000
0!
0%
b111 *
0-
02
b111 6
#430070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#430080000000
0!
0%
b0 *
0-
02
b0 6
#430090000000
1!
1%
1-
12
#430100000000
0!
0%
b1 *
0-
02
b1 6
#430110000000
1!
1%
1-
12
#430120000000
0!
0%
b10 *
0-
02
b10 6
#430130000000
1!
1%
1-
12
#430140000000
0!
0%
b11 *
0-
02
b11 6
#430150000000
1!
1%
1-
12
15
#430160000000
0!
0%
b100 *
0-
02
b100 6
#430170000000
1!
1%
1-
12
#430180000000
0!
0%
b101 *
0-
02
b101 6
#430190000000
1!
1%
1-
12
#430200000000
0!
0%
b110 *
0-
02
b110 6
#430210000000
1!
1%
1-
12
#430220000000
0!
0%
b111 *
0-
02
b111 6
#430230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#430240000000
0!
0%
b0 *
0-
02
b0 6
#430250000000
1!
1%
1-
12
#430260000000
0!
0%
b1 *
0-
02
b1 6
#430270000000
1!
1%
1-
12
#430280000000
0!
0%
b10 *
0-
02
b10 6
#430290000000
1!
1%
1-
12
#430300000000
0!
0%
b11 *
0-
02
b11 6
#430310000000
1!
1%
1-
12
15
#430320000000
0!
0%
b100 *
0-
02
b100 6
#430330000000
1!
1%
1-
12
#430340000000
0!
0%
b101 *
0-
02
b101 6
#430350000000
1!
1%
1-
12
#430360000000
0!
0%
b110 *
0-
02
b110 6
#430370000000
1!
1%
1-
12
#430380000000
0!
0%
b111 *
0-
02
b111 6
#430390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#430400000000
0!
0%
b0 *
0-
02
b0 6
#430410000000
1!
1%
1-
12
#430420000000
0!
0%
b1 *
0-
02
b1 6
#430430000000
1!
1%
1-
12
#430440000000
0!
0%
b10 *
0-
02
b10 6
#430450000000
1!
1%
1-
12
#430460000000
0!
0%
b11 *
0-
02
b11 6
#430470000000
1!
1%
1-
12
15
#430480000000
0!
0%
b100 *
0-
02
b100 6
#430490000000
1!
1%
1-
12
#430500000000
0!
0%
b101 *
0-
02
b101 6
#430510000000
1!
1%
1-
12
#430520000000
0!
0%
b110 *
0-
02
b110 6
#430530000000
1!
1%
1-
12
#430540000000
0!
0%
b111 *
0-
02
b111 6
#430550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#430560000000
0!
0%
b0 *
0-
02
b0 6
#430570000000
1!
1%
1-
12
#430580000000
0!
0%
b1 *
0-
02
b1 6
#430590000000
1!
1%
1-
12
#430600000000
0!
0%
b10 *
0-
02
b10 6
#430610000000
1!
1%
1-
12
#430620000000
0!
0%
b11 *
0-
02
b11 6
#430630000000
1!
1%
1-
12
15
#430640000000
0!
0%
b100 *
0-
02
b100 6
#430650000000
1!
1%
1-
12
#430660000000
0!
0%
b101 *
0-
02
b101 6
#430670000000
1!
1%
1-
12
#430680000000
0!
0%
b110 *
0-
02
b110 6
#430690000000
1!
1%
1-
12
#430700000000
0!
0%
b111 *
0-
02
b111 6
#430710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#430720000000
0!
0%
b0 *
0-
02
b0 6
#430730000000
1!
1%
1-
12
#430740000000
0!
0%
b1 *
0-
02
b1 6
#430750000000
1!
1%
1-
12
#430760000000
0!
0%
b10 *
0-
02
b10 6
#430770000000
1!
1%
1-
12
#430780000000
0!
0%
b11 *
0-
02
b11 6
#430790000000
1!
1%
1-
12
15
#430800000000
0!
0%
b100 *
0-
02
b100 6
#430810000000
1!
1%
1-
12
#430820000000
0!
0%
b101 *
0-
02
b101 6
#430830000000
1!
1%
1-
12
#430840000000
0!
0%
b110 *
0-
02
b110 6
#430850000000
1!
1%
1-
12
#430860000000
0!
0%
b111 *
0-
02
b111 6
#430870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#430880000000
0!
0%
b0 *
0-
02
b0 6
#430890000000
1!
1%
1-
12
#430900000000
0!
0%
b1 *
0-
02
b1 6
#430910000000
1!
1%
1-
12
#430920000000
0!
0%
b10 *
0-
02
b10 6
#430930000000
1!
1%
1-
12
#430940000000
0!
0%
b11 *
0-
02
b11 6
#430950000000
1!
1%
1-
12
15
#430960000000
0!
0%
b100 *
0-
02
b100 6
#430970000000
1!
1%
1-
12
#430980000000
0!
0%
b101 *
0-
02
b101 6
#430990000000
1!
1%
1-
12
#431000000000
0!
0%
b110 *
0-
02
b110 6
#431010000000
1!
1%
1-
12
#431020000000
0!
0%
b111 *
0-
02
b111 6
#431030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#431040000000
0!
0%
b0 *
0-
02
b0 6
#431050000000
1!
1%
1-
12
#431060000000
0!
0%
b1 *
0-
02
b1 6
#431070000000
1!
1%
1-
12
#431080000000
0!
0%
b10 *
0-
02
b10 6
#431090000000
1!
1%
1-
12
#431100000000
0!
0%
b11 *
0-
02
b11 6
#431110000000
1!
1%
1-
12
15
#431120000000
0!
0%
b100 *
0-
02
b100 6
#431130000000
1!
1%
1-
12
#431140000000
0!
0%
b101 *
0-
02
b101 6
#431150000000
1!
1%
1-
12
#431160000000
0!
0%
b110 *
0-
02
b110 6
#431170000000
1!
1%
1-
12
#431180000000
0!
0%
b111 *
0-
02
b111 6
#431190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#431200000000
0!
0%
b0 *
0-
02
b0 6
#431210000000
1!
1%
1-
12
#431220000000
0!
0%
b1 *
0-
02
b1 6
#431230000000
1!
1%
1-
12
#431240000000
0!
0%
b10 *
0-
02
b10 6
#431250000000
1!
1%
1-
12
#431260000000
0!
0%
b11 *
0-
02
b11 6
#431270000000
1!
1%
1-
12
15
#431280000000
0!
0%
b100 *
0-
02
b100 6
#431290000000
1!
1%
1-
12
#431300000000
0!
0%
b101 *
0-
02
b101 6
#431310000000
1!
1%
1-
12
#431320000000
0!
0%
b110 *
0-
02
b110 6
#431330000000
1!
1%
1-
12
#431340000000
0!
0%
b111 *
0-
02
b111 6
#431350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#431360000000
0!
0%
b0 *
0-
02
b0 6
#431370000000
1!
1%
1-
12
#431380000000
0!
0%
b1 *
0-
02
b1 6
#431390000000
1!
1%
1-
12
#431400000000
0!
0%
b10 *
0-
02
b10 6
#431410000000
1!
1%
1-
12
#431420000000
0!
0%
b11 *
0-
02
b11 6
#431430000000
1!
1%
1-
12
15
#431440000000
0!
0%
b100 *
0-
02
b100 6
#431450000000
1!
1%
1-
12
#431460000000
0!
0%
b101 *
0-
02
b101 6
#431470000000
1!
1%
1-
12
#431480000000
0!
0%
b110 *
0-
02
b110 6
#431490000000
1!
1%
1-
12
#431500000000
0!
0%
b111 *
0-
02
b111 6
#431510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#431520000000
0!
0%
b0 *
0-
02
b0 6
#431530000000
1!
1%
1-
12
#431540000000
0!
0%
b1 *
0-
02
b1 6
#431550000000
1!
1%
1-
12
#431560000000
0!
0%
b10 *
0-
02
b10 6
#431570000000
1!
1%
1-
12
#431580000000
0!
0%
b11 *
0-
02
b11 6
#431590000000
1!
1%
1-
12
15
#431600000000
0!
0%
b100 *
0-
02
b100 6
#431610000000
1!
1%
1-
12
#431620000000
0!
0%
b101 *
0-
02
b101 6
#431630000000
1!
1%
1-
12
#431640000000
0!
0%
b110 *
0-
02
b110 6
#431650000000
1!
1%
1-
12
#431660000000
0!
0%
b111 *
0-
02
b111 6
#431670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#431680000000
0!
0%
b0 *
0-
02
b0 6
#431690000000
1!
1%
1-
12
#431700000000
0!
0%
b1 *
0-
02
b1 6
#431710000000
1!
1%
1-
12
#431720000000
0!
0%
b10 *
0-
02
b10 6
#431730000000
1!
1%
1-
12
#431740000000
0!
0%
b11 *
0-
02
b11 6
#431750000000
1!
1%
1-
12
15
#431760000000
0!
0%
b100 *
0-
02
b100 6
#431770000000
1!
1%
1-
12
#431780000000
0!
0%
b101 *
0-
02
b101 6
#431790000000
1!
1%
1-
12
#431800000000
0!
0%
b110 *
0-
02
b110 6
#431810000000
1!
1%
1-
12
#431820000000
0!
0%
b111 *
0-
02
b111 6
#431830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#431840000000
0!
0%
b0 *
0-
02
b0 6
#431850000000
1!
1%
1-
12
#431860000000
0!
0%
b1 *
0-
02
b1 6
#431870000000
1!
1%
1-
12
#431880000000
0!
0%
b10 *
0-
02
b10 6
#431890000000
1!
1%
1-
12
#431900000000
0!
0%
b11 *
0-
02
b11 6
#431910000000
1!
1%
1-
12
15
#431920000000
0!
0%
b100 *
0-
02
b100 6
#431930000000
1!
1%
1-
12
#431940000000
0!
0%
b101 *
0-
02
b101 6
#431950000000
1!
1%
1-
12
#431960000000
0!
0%
b110 *
0-
02
b110 6
#431970000000
1!
1%
1-
12
#431980000000
0!
0%
b111 *
0-
02
b111 6
#431990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#432000000000
0!
0%
b0 *
0-
02
b0 6
#432010000000
1!
1%
1-
12
#432020000000
0!
0%
b1 *
0-
02
b1 6
#432030000000
1!
1%
1-
12
#432040000000
0!
0%
b10 *
0-
02
b10 6
#432050000000
1!
1%
1-
12
#432060000000
0!
0%
b11 *
0-
02
b11 6
#432070000000
1!
1%
1-
12
15
#432080000000
0!
0%
b100 *
0-
02
b100 6
#432090000000
1!
1%
1-
12
#432100000000
0!
0%
b101 *
0-
02
b101 6
#432110000000
1!
1%
1-
12
#432120000000
0!
0%
b110 *
0-
02
b110 6
#432130000000
1!
1%
1-
12
#432140000000
0!
0%
b111 *
0-
02
b111 6
#432150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#432160000000
0!
0%
b0 *
0-
02
b0 6
#432170000000
1!
1%
1-
12
#432180000000
0!
0%
b1 *
0-
02
b1 6
#432190000000
1!
1%
1-
12
#432200000000
0!
0%
b10 *
0-
02
b10 6
#432210000000
1!
1%
1-
12
#432220000000
0!
0%
b11 *
0-
02
b11 6
#432230000000
1!
1%
1-
12
15
#432240000000
0!
0%
b100 *
0-
02
b100 6
#432250000000
1!
1%
1-
12
#432260000000
0!
0%
b101 *
0-
02
b101 6
#432270000000
1!
1%
1-
12
#432280000000
0!
0%
b110 *
0-
02
b110 6
#432290000000
1!
1%
1-
12
#432300000000
0!
0%
b111 *
0-
02
b111 6
#432310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#432320000000
0!
0%
b0 *
0-
02
b0 6
#432330000000
1!
1%
1-
12
#432340000000
0!
0%
b1 *
0-
02
b1 6
#432350000000
1!
1%
1-
12
#432360000000
0!
0%
b10 *
0-
02
b10 6
#432370000000
1!
1%
1-
12
#432380000000
0!
0%
b11 *
0-
02
b11 6
#432390000000
1!
1%
1-
12
15
#432400000000
0!
0%
b100 *
0-
02
b100 6
#432410000000
1!
1%
1-
12
#432420000000
0!
0%
b101 *
0-
02
b101 6
#432430000000
1!
1%
1-
12
#432440000000
0!
0%
b110 *
0-
02
b110 6
#432450000000
1!
1%
1-
12
#432460000000
0!
0%
b111 *
0-
02
b111 6
#432470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#432480000000
0!
0%
b0 *
0-
02
b0 6
#432490000000
1!
1%
1-
12
#432500000000
0!
0%
b1 *
0-
02
b1 6
#432510000000
1!
1%
1-
12
#432520000000
0!
0%
b10 *
0-
02
b10 6
#432530000000
1!
1%
1-
12
#432540000000
0!
0%
b11 *
0-
02
b11 6
#432550000000
1!
1%
1-
12
15
#432560000000
0!
0%
b100 *
0-
02
b100 6
#432570000000
1!
1%
1-
12
#432580000000
0!
0%
b101 *
0-
02
b101 6
#432590000000
1!
1%
1-
12
#432600000000
0!
0%
b110 *
0-
02
b110 6
#432610000000
1!
1%
1-
12
#432620000000
0!
0%
b111 *
0-
02
b111 6
#432630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#432640000000
0!
0%
b0 *
0-
02
b0 6
#432650000000
1!
1%
1-
12
#432660000000
0!
0%
b1 *
0-
02
b1 6
#432670000000
1!
1%
1-
12
#432680000000
0!
0%
b10 *
0-
02
b10 6
#432690000000
1!
1%
1-
12
#432700000000
0!
0%
b11 *
0-
02
b11 6
#432710000000
1!
1%
1-
12
15
#432720000000
0!
0%
b100 *
0-
02
b100 6
#432730000000
1!
1%
1-
12
#432740000000
0!
0%
b101 *
0-
02
b101 6
#432750000000
1!
1%
1-
12
#432760000000
0!
0%
b110 *
0-
02
b110 6
#432770000000
1!
1%
1-
12
#432780000000
0!
0%
b111 *
0-
02
b111 6
#432790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#432800000000
0!
0%
b0 *
0-
02
b0 6
#432810000000
1!
1%
1-
12
#432820000000
0!
0%
b1 *
0-
02
b1 6
#432830000000
1!
1%
1-
12
#432840000000
0!
0%
b10 *
0-
02
b10 6
#432850000000
1!
1%
1-
12
#432860000000
0!
0%
b11 *
0-
02
b11 6
#432870000000
1!
1%
1-
12
15
#432880000000
0!
0%
b100 *
0-
02
b100 6
#432890000000
1!
1%
1-
12
#432900000000
0!
0%
b101 *
0-
02
b101 6
#432910000000
1!
1%
1-
12
#432920000000
0!
0%
b110 *
0-
02
b110 6
#432930000000
1!
1%
1-
12
#432940000000
0!
0%
b111 *
0-
02
b111 6
#432950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#432960000000
0!
0%
b0 *
0-
02
b0 6
#432970000000
1!
1%
1-
12
#432980000000
0!
0%
b1 *
0-
02
b1 6
#432990000000
1!
1%
1-
12
#433000000000
0!
0%
b10 *
0-
02
b10 6
#433010000000
1!
1%
1-
12
#433020000000
0!
0%
b11 *
0-
02
b11 6
#433030000000
1!
1%
1-
12
15
#433040000000
0!
0%
b100 *
0-
02
b100 6
#433050000000
1!
1%
1-
12
#433060000000
0!
0%
b101 *
0-
02
b101 6
#433070000000
1!
1%
1-
12
#433080000000
0!
0%
b110 *
0-
02
b110 6
#433090000000
1!
1%
1-
12
#433100000000
0!
0%
b111 *
0-
02
b111 6
#433110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#433120000000
0!
0%
b0 *
0-
02
b0 6
#433130000000
1!
1%
1-
12
#433140000000
0!
0%
b1 *
0-
02
b1 6
#433150000000
1!
1%
1-
12
#433160000000
0!
0%
b10 *
0-
02
b10 6
#433170000000
1!
1%
1-
12
#433180000000
0!
0%
b11 *
0-
02
b11 6
#433190000000
1!
1%
1-
12
15
#433200000000
0!
0%
b100 *
0-
02
b100 6
#433210000000
1!
1%
1-
12
#433220000000
0!
0%
b101 *
0-
02
b101 6
#433230000000
1!
1%
1-
12
#433240000000
0!
0%
b110 *
0-
02
b110 6
#433250000000
1!
1%
1-
12
#433260000000
0!
0%
b111 *
0-
02
b111 6
#433270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#433280000000
0!
0%
b0 *
0-
02
b0 6
#433290000000
1!
1%
1-
12
#433300000000
0!
0%
b1 *
0-
02
b1 6
#433310000000
1!
1%
1-
12
#433320000000
0!
0%
b10 *
0-
02
b10 6
#433330000000
1!
1%
1-
12
#433340000000
0!
0%
b11 *
0-
02
b11 6
#433350000000
1!
1%
1-
12
15
#433360000000
0!
0%
b100 *
0-
02
b100 6
#433370000000
1!
1%
1-
12
#433380000000
0!
0%
b101 *
0-
02
b101 6
#433390000000
1!
1%
1-
12
#433400000000
0!
0%
b110 *
0-
02
b110 6
#433410000000
1!
1%
1-
12
#433420000000
0!
0%
b111 *
0-
02
b111 6
#433430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#433440000000
0!
0%
b0 *
0-
02
b0 6
#433450000000
1!
1%
1-
12
#433460000000
0!
0%
b1 *
0-
02
b1 6
#433470000000
1!
1%
1-
12
#433480000000
0!
0%
b10 *
0-
02
b10 6
#433490000000
1!
1%
1-
12
#433500000000
0!
0%
b11 *
0-
02
b11 6
#433510000000
1!
1%
1-
12
15
#433520000000
0!
0%
b100 *
0-
02
b100 6
#433530000000
1!
1%
1-
12
#433540000000
0!
0%
b101 *
0-
02
b101 6
#433550000000
1!
1%
1-
12
#433560000000
0!
0%
b110 *
0-
02
b110 6
#433570000000
1!
1%
1-
12
#433580000000
0!
0%
b111 *
0-
02
b111 6
#433590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#433600000000
0!
0%
b0 *
0-
02
b0 6
#433610000000
1!
1%
1-
12
#433620000000
0!
0%
b1 *
0-
02
b1 6
#433630000000
1!
1%
1-
12
#433640000000
0!
0%
b10 *
0-
02
b10 6
#433650000000
1!
1%
1-
12
#433660000000
0!
0%
b11 *
0-
02
b11 6
#433670000000
1!
1%
1-
12
15
#433680000000
0!
0%
b100 *
0-
02
b100 6
#433690000000
1!
1%
1-
12
#433700000000
0!
0%
b101 *
0-
02
b101 6
#433710000000
1!
1%
1-
12
#433720000000
0!
0%
b110 *
0-
02
b110 6
#433730000000
1!
1%
1-
12
#433740000000
0!
0%
b111 *
0-
02
b111 6
#433750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#433760000000
0!
0%
b0 *
0-
02
b0 6
#433770000000
1!
1%
1-
12
#433780000000
0!
0%
b1 *
0-
02
b1 6
#433790000000
1!
1%
1-
12
#433800000000
0!
0%
b10 *
0-
02
b10 6
#433810000000
1!
1%
1-
12
#433820000000
0!
0%
b11 *
0-
02
b11 6
#433830000000
1!
1%
1-
12
15
#433840000000
0!
0%
b100 *
0-
02
b100 6
#433850000000
1!
1%
1-
12
#433860000000
0!
0%
b101 *
0-
02
b101 6
#433870000000
1!
1%
1-
12
#433880000000
0!
0%
b110 *
0-
02
b110 6
#433890000000
1!
1%
1-
12
#433900000000
0!
0%
b111 *
0-
02
b111 6
#433910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#433920000000
0!
0%
b0 *
0-
02
b0 6
#433930000000
1!
1%
1-
12
#433940000000
0!
0%
b1 *
0-
02
b1 6
#433950000000
1!
1%
1-
12
#433960000000
0!
0%
b10 *
0-
02
b10 6
#433970000000
1!
1%
1-
12
#433980000000
0!
0%
b11 *
0-
02
b11 6
#433990000000
1!
1%
1-
12
15
#434000000000
0!
0%
b100 *
0-
02
b100 6
#434010000000
1!
1%
1-
12
#434020000000
0!
0%
b101 *
0-
02
b101 6
#434030000000
1!
1%
1-
12
#434040000000
0!
0%
b110 *
0-
02
b110 6
#434050000000
1!
1%
1-
12
#434060000000
0!
0%
b111 *
0-
02
b111 6
#434070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#434080000000
0!
0%
b0 *
0-
02
b0 6
#434090000000
1!
1%
1-
12
#434100000000
0!
0%
b1 *
0-
02
b1 6
#434110000000
1!
1%
1-
12
#434120000000
0!
0%
b10 *
0-
02
b10 6
#434130000000
1!
1%
1-
12
#434140000000
0!
0%
b11 *
0-
02
b11 6
#434150000000
1!
1%
1-
12
15
#434160000000
0!
0%
b100 *
0-
02
b100 6
#434170000000
1!
1%
1-
12
#434180000000
0!
0%
b101 *
0-
02
b101 6
#434190000000
1!
1%
1-
12
#434200000000
0!
0%
b110 *
0-
02
b110 6
#434210000000
1!
1%
1-
12
#434220000000
0!
0%
b111 *
0-
02
b111 6
#434230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#434240000000
0!
0%
b0 *
0-
02
b0 6
#434250000000
1!
1%
1-
12
#434260000000
0!
0%
b1 *
0-
02
b1 6
#434270000000
1!
1%
1-
12
#434280000000
0!
0%
b10 *
0-
02
b10 6
#434290000000
1!
1%
1-
12
#434300000000
0!
0%
b11 *
0-
02
b11 6
#434310000000
1!
1%
1-
12
15
#434320000000
0!
0%
b100 *
0-
02
b100 6
#434330000000
1!
1%
1-
12
#434340000000
0!
0%
b101 *
0-
02
b101 6
#434350000000
1!
1%
1-
12
#434360000000
0!
0%
b110 *
0-
02
b110 6
#434370000000
1!
1%
1-
12
#434380000000
0!
0%
b111 *
0-
02
b111 6
#434390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#434400000000
0!
0%
b0 *
0-
02
b0 6
#434410000000
1!
1%
1-
12
#434420000000
0!
0%
b1 *
0-
02
b1 6
#434430000000
1!
1%
1-
12
#434440000000
0!
0%
b10 *
0-
02
b10 6
#434450000000
1!
1%
1-
12
#434460000000
0!
0%
b11 *
0-
02
b11 6
#434470000000
1!
1%
1-
12
15
#434480000000
0!
0%
b100 *
0-
02
b100 6
#434490000000
1!
1%
1-
12
#434500000000
0!
0%
b101 *
0-
02
b101 6
#434510000000
1!
1%
1-
12
#434520000000
0!
0%
b110 *
0-
02
b110 6
#434530000000
1!
1%
1-
12
#434540000000
0!
0%
b111 *
0-
02
b111 6
#434550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#434560000000
0!
0%
b0 *
0-
02
b0 6
#434570000000
1!
1%
1-
12
#434580000000
0!
0%
b1 *
0-
02
b1 6
#434590000000
1!
1%
1-
12
#434600000000
0!
0%
b10 *
0-
02
b10 6
#434610000000
1!
1%
1-
12
#434620000000
0!
0%
b11 *
0-
02
b11 6
#434630000000
1!
1%
1-
12
15
#434640000000
0!
0%
b100 *
0-
02
b100 6
#434650000000
1!
1%
1-
12
#434660000000
0!
0%
b101 *
0-
02
b101 6
#434670000000
1!
1%
1-
12
#434680000000
0!
0%
b110 *
0-
02
b110 6
#434690000000
1!
1%
1-
12
#434700000000
0!
0%
b111 *
0-
02
b111 6
#434710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#434720000000
0!
0%
b0 *
0-
02
b0 6
#434730000000
1!
1%
1-
12
#434740000000
0!
0%
b1 *
0-
02
b1 6
#434750000000
1!
1%
1-
12
#434760000000
0!
0%
b10 *
0-
02
b10 6
#434770000000
1!
1%
1-
12
#434780000000
0!
0%
b11 *
0-
02
b11 6
#434790000000
1!
1%
1-
12
15
#434800000000
0!
0%
b100 *
0-
02
b100 6
#434810000000
1!
1%
1-
12
#434820000000
0!
0%
b101 *
0-
02
b101 6
#434830000000
1!
1%
1-
12
#434840000000
0!
0%
b110 *
0-
02
b110 6
#434850000000
1!
1%
1-
12
#434860000000
0!
0%
b111 *
0-
02
b111 6
#434870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#434880000000
0!
0%
b0 *
0-
02
b0 6
#434890000000
1!
1%
1-
12
#434900000000
0!
0%
b1 *
0-
02
b1 6
#434910000000
1!
1%
1-
12
#434920000000
0!
0%
b10 *
0-
02
b10 6
#434930000000
1!
1%
1-
12
#434940000000
0!
0%
b11 *
0-
02
b11 6
#434950000000
1!
1%
1-
12
15
#434960000000
0!
0%
b100 *
0-
02
b100 6
#434970000000
1!
1%
1-
12
#434980000000
0!
0%
b101 *
0-
02
b101 6
#434990000000
1!
1%
1-
12
#435000000000
0!
0%
b110 *
0-
02
b110 6
#435010000000
1!
1%
1-
12
#435020000000
0!
0%
b111 *
0-
02
b111 6
#435030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#435040000000
0!
0%
b0 *
0-
02
b0 6
#435050000000
1!
1%
1-
12
#435060000000
0!
0%
b1 *
0-
02
b1 6
#435070000000
1!
1%
1-
12
#435080000000
0!
0%
b10 *
0-
02
b10 6
#435090000000
1!
1%
1-
12
#435100000000
0!
0%
b11 *
0-
02
b11 6
#435110000000
1!
1%
1-
12
15
#435120000000
0!
0%
b100 *
0-
02
b100 6
#435130000000
1!
1%
1-
12
#435140000000
0!
0%
b101 *
0-
02
b101 6
#435150000000
1!
1%
1-
12
#435160000000
0!
0%
b110 *
0-
02
b110 6
#435170000000
1!
1%
1-
12
#435180000000
0!
0%
b111 *
0-
02
b111 6
#435190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#435200000000
0!
0%
b0 *
0-
02
b0 6
#435210000000
1!
1%
1-
12
#435220000000
0!
0%
b1 *
0-
02
b1 6
#435230000000
1!
1%
1-
12
#435240000000
0!
0%
b10 *
0-
02
b10 6
#435250000000
1!
1%
1-
12
#435260000000
0!
0%
b11 *
0-
02
b11 6
#435270000000
1!
1%
1-
12
15
#435280000000
0!
0%
b100 *
0-
02
b100 6
#435290000000
1!
1%
1-
12
#435300000000
0!
0%
b101 *
0-
02
b101 6
#435310000000
1!
1%
1-
12
#435320000000
0!
0%
b110 *
0-
02
b110 6
#435330000000
1!
1%
1-
12
#435340000000
0!
0%
b111 *
0-
02
b111 6
#435350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#435360000000
0!
0%
b0 *
0-
02
b0 6
#435370000000
1!
1%
1-
12
#435380000000
0!
0%
b1 *
0-
02
b1 6
#435390000000
1!
1%
1-
12
#435400000000
0!
0%
b10 *
0-
02
b10 6
#435410000000
1!
1%
1-
12
#435420000000
0!
0%
b11 *
0-
02
b11 6
#435430000000
1!
1%
1-
12
15
#435440000000
0!
0%
b100 *
0-
02
b100 6
#435450000000
1!
1%
1-
12
#435460000000
0!
0%
b101 *
0-
02
b101 6
#435470000000
1!
1%
1-
12
#435480000000
0!
0%
b110 *
0-
02
b110 6
#435490000000
1!
1%
1-
12
#435500000000
0!
0%
b111 *
0-
02
b111 6
#435510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#435520000000
0!
0%
b0 *
0-
02
b0 6
#435530000000
1!
1%
1-
12
#435540000000
0!
0%
b1 *
0-
02
b1 6
#435550000000
1!
1%
1-
12
#435560000000
0!
0%
b10 *
0-
02
b10 6
#435570000000
1!
1%
1-
12
#435580000000
0!
0%
b11 *
0-
02
b11 6
#435590000000
1!
1%
1-
12
15
#435600000000
0!
0%
b100 *
0-
02
b100 6
#435610000000
1!
1%
1-
12
#435620000000
0!
0%
b101 *
0-
02
b101 6
#435630000000
1!
1%
1-
12
#435640000000
0!
0%
b110 *
0-
02
b110 6
#435650000000
1!
1%
1-
12
#435660000000
0!
0%
b111 *
0-
02
b111 6
#435670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#435680000000
0!
0%
b0 *
0-
02
b0 6
#435690000000
1!
1%
1-
12
#435700000000
0!
0%
b1 *
0-
02
b1 6
#435710000000
1!
1%
1-
12
#435720000000
0!
0%
b10 *
0-
02
b10 6
#435730000000
1!
1%
1-
12
#435740000000
0!
0%
b11 *
0-
02
b11 6
#435750000000
1!
1%
1-
12
15
#435760000000
0!
0%
b100 *
0-
02
b100 6
#435770000000
1!
1%
1-
12
#435780000000
0!
0%
b101 *
0-
02
b101 6
#435790000000
1!
1%
1-
12
#435800000000
0!
0%
b110 *
0-
02
b110 6
#435810000000
1!
1%
1-
12
#435820000000
0!
0%
b111 *
0-
02
b111 6
#435830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#435840000000
0!
0%
b0 *
0-
02
b0 6
#435850000000
1!
1%
1-
12
#435860000000
0!
0%
b1 *
0-
02
b1 6
#435870000000
1!
1%
1-
12
#435880000000
0!
0%
b10 *
0-
02
b10 6
#435890000000
1!
1%
1-
12
#435900000000
0!
0%
b11 *
0-
02
b11 6
#435910000000
1!
1%
1-
12
15
#435920000000
0!
0%
b100 *
0-
02
b100 6
#435930000000
1!
1%
1-
12
#435940000000
0!
0%
b101 *
0-
02
b101 6
#435950000000
1!
1%
1-
12
#435960000000
0!
0%
b110 *
0-
02
b110 6
#435970000000
1!
1%
1-
12
#435980000000
0!
0%
b111 *
0-
02
b111 6
#435990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#436000000000
0!
0%
b0 *
0-
02
b0 6
#436010000000
1!
1%
1-
12
#436020000000
0!
0%
b1 *
0-
02
b1 6
#436030000000
1!
1%
1-
12
#436040000000
0!
0%
b10 *
0-
02
b10 6
#436050000000
1!
1%
1-
12
#436060000000
0!
0%
b11 *
0-
02
b11 6
#436070000000
1!
1%
1-
12
15
#436080000000
0!
0%
b100 *
0-
02
b100 6
#436090000000
1!
1%
1-
12
#436100000000
0!
0%
b101 *
0-
02
b101 6
#436110000000
1!
1%
1-
12
#436120000000
0!
0%
b110 *
0-
02
b110 6
#436130000000
1!
1%
1-
12
#436140000000
0!
0%
b111 *
0-
02
b111 6
#436150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#436160000000
0!
0%
b0 *
0-
02
b0 6
#436170000000
1!
1%
1-
12
#436180000000
0!
0%
b1 *
0-
02
b1 6
#436190000000
1!
1%
1-
12
#436200000000
0!
0%
b10 *
0-
02
b10 6
#436210000000
1!
1%
1-
12
#436220000000
0!
0%
b11 *
0-
02
b11 6
#436230000000
1!
1%
1-
12
15
#436240000000
0!
0%
b100 *
0-
02
b100 6
#436250000000
1!
1%
1-
12
#436260000000
0!
0%
b101 *
0-
02
b101 6
#436270000000
1!
1%
1-
12
#436280000000
0!
0%
b110 *
0-
02
b110 6
#436290000000
1!
1%
1-
12
#436300000000
0!
0%
b111 *
0-
02
b111 6
#436310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#436320000000
0!
0%
b0 *
0-
02
b0 6
#436330000000
1!
1%
1-
12
#436340000000
0!
0%
b1 *
0-
02
b1 6
#436350000000
1!
1%
1-
12
#436360000000
0!
0%
b10 *
0-
02
b10 6
#436370000000
1!
1%
1-
12
#436380000000
0!
0%
b11 *
0-
02
b11 6
#436390000000
1!
1%
1-
12
15
#436400000000
0!
0%
b100 *
0-
02
b100 6
#436410000000
1!
1%
1-
12
#436420000000
0!
0%
b101 *
0-
02
b101 6
#436430000000
1!
1%
1-
12
#436440000000
0!
0%
b110 *
0-
02
b110 6
#436450000000
1!
1%
1-
12
#436460000000
0!
0%
b111 *
0-
02
b111 6
#436470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#436480000000
0!
0%
b0 *
0-
02
b0 6
#436490000000
1!
1%
1-
12
#436500000000
0!
0%
b1 *
0-
02
b1 6
#436510000000
1!
1%
1-
12
#436520000000
0!
0%
b10 *
0-
02
b10 6
#436530000000
1!
1%
1-
12
#436540000000
0!
0%
b11 *
0-
02
b11 6
#436550000000
1!
1%
1-
12
15
#436560000000
0!
0%
b100 *
0-
02
b100 6
#436570000000
1!
1%
1-
12
#436580000000
0!
0%
b101 *
0-
02
b101 6
#436590000000
1!
1%
1-
12
#436600000000
0!
0%
b110 *
0-
02
b110 6
#436610000000
1!
1%
1-
12
#436620000000
0!
0%
b111 *
0-
02
b111 6
#436630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#436640000000
0!
0%
b0 *
0-
02
b0 6
#436650000000
1!
1%
1-
12
#436660000000
0!
0%
b1 *
0-
02
b1 6
#436670000000
1!
1%
1-
12
#436680000000
0!
0%
b10 *
0-
02
b10 6
#436690000000
1!
1%
1-
12
#436700000000
0!
0%
b11 *
0-
02
b11 6
#436710000000
1!
1%
1-
12
15
#436720000000
0!
0%
b100 *
0-
02
b100 6
#436730000000
1!
1%
1-
12
#436740000000
0!
0%
b101 *
0-
02
b101 6
#436750000000
1!
1%
1-
12
#436760000000
0!
0%
b110 *
0-
02
b110 6
#436770000000
1!
1%
1-
12
#436780000000
0!
0%
b111 *
0-
02
b111 6
#436790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#436800000000
0!
0%
b0 *
0-
02
b0 6
#436810000000
1!
1%
1-
12
#436820000000
0!
0%
b1 *
0-
02
b1 6
#436830000000
1!
1%
1-
12
#436840000000
0!
0%
b10 *
0-
02
b10 6
#436850000000
1!
1%
1-
12
#436860000000
0!
0%
b11 *
0-
02
b11 6
#436870000000
1!
1%
1-
12
15
#436880000000
0!
0%
b100 *
0-
02
b100 6
#436890000000
1!
1%
1-
12
#436900000000
0!
0%
b101 *
0-
02
b101 6
#436910000000
1!
1%
1-
12
#436920000000
0!
0%
b110 *
0-
02
b110 6
#436930000000
1!
1%
1-
12
#436940000000
0!
0%
b111 *
0-
02
b111 6
#436950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#436960000000
0!
0%
b0 *
0-
02
b0 6
#436970000000
1!
1%
1-
12
#436980000000
0!
0%
b1 *
0-
02
b1 6
#436990000000
1!
1%
1-
12
#437000000000
0!
0%
b10 *
0-
02
b10 6
#437010000000
1!
1%
1-
12
#437020000000
0!
0%
b11 *
0-
02
b11 6
#437030000000
1!
1%
1-
12
15
#437040000000
0!
0%
b100 *
0-
02
b100 6
#437050000000
1!
1%
1-
12
#437060000000
0!
0%
b101 *
0-
02
b101 6
#437070000000
1!
1%
1-
12
#437080000000
0!
0%
b110 *
0-
02
b110 6
#437090000000
1!
1%
1-
12
#437100000000
0!
0%
b111 *
0-
02
b111 6
#437110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#437120000000
0!
0%
b0 *
0-
02
b0 6
#437130000000
1!
1%
1-
12
#437140000000
0!
0%
b1 *
0-
02
b1 6
#437150000000
1!
1%
1-
12
#437160000000
0!
0%
b10 *
0-
02
b10 6
#437170000000
1!
1%
1-
12
#437180000000
0!
0%
b11 *
0-
02
b11 6
#437190000000
1!
1%
1-
12
15
#437200000000
0!
0%
b100 *
0-
02
b100 6
#437210000000
1!
1%
1-
12
#437220000000
0!
0%
b101 *
0-
02
b101 6
#437230000000
1!
1%
1-
12
#437240000000
0!
0%
b110 *
0-
02
b110 6
#437250000000
1!
1%
1-
12
#437260000000
0!
0%
b111 *
0-
02
b111 6
#437270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#437280000000
0!
0%
b0 *
0-
02
b0 6
#437290000000
1!
1%
1-
12
#437300000000
0!
0%
b1 *
0-
02
b1 6
#437310000000
1!
1%
1-
12
#437320000000
0!
0%
b10 *
0-
02
b10 6
#437330000000
1!
1%
1-
12
#437340000000
0!
0%
b11 *
0-
02
b11 6
#437350000000
1!
1%
1-
12
15
#437360000000
0!
0%
b100 *
0-
02
b100 6
#437370000000
1!
1%
1-
12
#437380000000
0!
0%
b101 *
0-
02
b101 6
#437390000000
1!
1%
1-
12
#437400000000
0!
0%
b110 *
0-
02
b110 6
#437410000000
1!
1%
1-
12
#437420000000
0!
0%
b111 *
0-
02
b111 6
#437430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#437440000000
0!
0%
b0 *
0-
02
b0 6
#437450000000
1!
1%
1-
12
#437460000000
0!
0%
b1 *
0-
02
b1 6
#437470000000
1!
1%
1-
12
#437480000000
0!
0%
b10 *
0-
02
b10 6
#437490000000
1!
1%
1-
12
#437500000000
0!
0%
b11 *
0-
02
b11 6
#437510000000
1!
1%
1-
12
15
#437520000000
0!
0%
b100 *
0-
02
b100 6
#437530000000
1!
1%
1-
12
#437540000000
0!
0%
b101 *
0-
02
b101 6
#437550000000
1!
1%
1-
12
#437560000000
0!
0%
b110 *
0-
02
b110 6
#437570000000
1!
1%
1-
12
#437580000000
0!
0%
b111 *
0-
02
b111 6
#437590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#437600000000
0!
0%
b0 *
0-
02
b0 6
#437610000000
1!
1%
1-
12
#437620000000
0!
0%
b1 *
0-
02
b1 6
#437630000000
1!
1%
1-
12
#437640000000
0!
0%
b10 *
0-
02
b10 6
#437650000000
1!
1%
1-
12
#437660000000
0!
0%
b11 *
0-
02
b11 6
#437670000000
1!
1%
1-
12
15
#437680000000
0!
0%
b100 *
0-
02
b100 6
#437690000000
1!
1%
1-
12
#437700000000
0!
0%
b101 *
0-
02
b101 6
#437710000000
1!
1%
1-
12
#437720000000
0!
0%
b110 *
0-
02
b110 6
#437730000000
1!
1%
1-
12
#437740000000
0!
0%
b111 *
0-
02
b111 6
#437750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#437760000000
0!
0%
b0 *
0-
02
b0 6
#437770000000
1!
1%
1-
12
#437780000000
0!
0%
b1 *
0-
02
b1 6
#437790000000
1!
1%
1-
12
#437800000000
0!
0%
b10 *
0-
02
b10 6
#437810000000
1!
1%
1-
12
#437820000000
0!
0%
b11 *
0-
02
b11 6
#437830000000
1!
1%
1-
12
15
#437840000000
0!
0%
b100 *
0-
02
b100 6
#437850000000
1!
1%
1-
12
#437860000000
0!
0%
b101 *
0-
02
b101 6
#437870000000
1!
1%
1-
12
#437880000000
0!
0%
b110 *
0-
02
b110 6
#437890000000
1!
1%
1-
12
#437900000000
0!
0%
b111 *
0-
02
b111 6
#437910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#437920000000
0!
0%
b0 *
0-
02
b0 6
#437930000000
1!
1%
1-
12
#437940000000
0!
0%
b1 *
0-
02
b1 6
#437950000000
1!
1%
1-
12
#437960000000
0!
0%
b10 *
0-
02
b10 6
#437970000000
1!
1%
1-
12
#437980000000
0!
0%
b11 *
0-
02
b11 6
#437990000000
1!
1%
1-
12
15
#438000000000
0!
0%
b100 *
0-
02
b100 6
#438010000000
1!
1%
1-
12
#438020000000
0!
0%
b101 *
0-
02
b101 6
#438030000000
1!
1%
1-
12
#438040000000
0!
0%
b110 *
0-
02
b110 6
#438050000000
1!
1%
1-
12
#438060000000
0!
0%
b111 *
0-
02
b111 6
#438070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#438080000000
0!
0%
b0 *
0-
02
b0 6
#438090000000
1!
1%
1-
12
#438100000000
0!
0%
b1 *
0-
02
b1 6
#438110000000
1!
1%
1-
12
#438120000000
0!
0%
b10 *
0-
02
b10 6
#438130000000
1!
1%
1-
12
#438140000000
0!
0%
b11 *
0-
02
b11 6
#438150000000
1!
1%
1-
12
15
#438160000000
0!
0%
b100 *
0-
02
b100 6
#438170000000
1!
1%
1-
12
#438180000000
0!
0%
b101 *
0-
02
b101 6
#438190000000
1!
1%
1-
12
#438200000000
0!
0%
b110 *
0-
02
b110 6
#438210000000
1!
1%
1-
12
#438220000000
0!
0%
b111 *
0-
02
b111 6
#438230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#438240000000
0!
0%
b0 *
0-
02
b0 6
#438250000000
1!
1%
1-
12
#438260000000
0!
0%
b1 *
0-
02
b1 6
#438270000000
1!
1%
1-
12
#438280000000
0!
0%
b10 *
0-
02
b10 6
#438290000000
1!
1%
1-
12
#438300000000
0!
0%
b11 *
0-
02
b11 6
#438310000000
1!
1%
1-
12
15
#438320000000
0!
0%
b100 *
0-
02
b100 6
#438330000000
1!
1%
1-
12
#438340000000
0!
0%
b101 *
0-
02
b101 6
#438350000000
1!
1%
1-
12
#438360000000
0!
0%
b110 *
0-
02
b110 6
#438370000000
1!
1%
1-
12
#438380000000
0!
0%
b111 *
0-
02
b111 6
#438390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#438400000000
0!
0%
b0 *
0-
02
b0 6
#438410000000
1!
1%
1-
12
#438420000000
0!
0%
b1 *
0-
02
b1 6
#438430000000
1!
1%
1-
12
#438440000000
0!
0%
b10 *
0-
02
b10 6
#438450000000
1!
1%
1-
12
#438460000000
0!
0%
b11 *
0-
02
b11 6
#438470000000
1!
1%
1-
12
15
#438480000000
0!
0%
b100 *
0-
02
b100 6
#438490000000
1!
1%
1-
12
#438500000000
0!
0%
b101 *
0-
02
b101 6
#438510000000
1!
1%
1-
12
#438520000000
0!
0%
b110 *
0-
02
b110 6
#438530000000
1!
1%
1-
12
#438540000000
0!
0%
b111 *
0-
02
b111 6
#438550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#438560000000
0!
0%
b0 *
0-
02
b0 6
#438570000000
1!
1%
1-
12
#438580000000
0!
0%
b1 *
0-
02
b1 6
#438590000000
1!
1%
1-
12
#438600000000
0!
0%
b10 *
0-
02
b10 6
#438610000000
1!
1%
1-
12
#438620000000
0!
0%
b11 *
0-
02
b11 6
#438630000000
1!
1%
1-
12
15
#438640000000
0!
0%
b100 *
0-
02
b100 6
#438650000000
1!
1%
1-
12
#438660000000
0!
0%
b101 *
0-
02
b101 6
#438670000000
1!
1%
1-
12
#438680000000
0!
0%
b110 *
0-
02
b110 6
#438690000000
1!
1%
1-
12
#438700000000
0!
0%
b111 *
0-
02
b111 6
#438710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#438720000000
0!
0%
b0 *
0-
02
b0 6
#438730000000
1!
1%
1-
12
#438740000000
0!
0%
b1 *
0-
02
b1 6
#438750000000
1!
1%
1-
12
#438760000000
0!
0%
b10 *
0-
02
b10 6
#438770000000
1!
1%
1-
12
#438780000000
0!
0%
b11 *
0-
02
b11 6
#438790000000
1!
1%
1-
12
15
#438800000000
0!
0%
b100 *
0-
02
b100 6
#438810000000
1!
1%
1-
12
#438820000000
0!
0%
b101 *
0-
02
b101 6
#438830000000
1!
1%
1-
12
#438840000000
0!
0%
b110 *
0-
02
b110 6
#438850000000
1!
1%
1-
12
#438860000000
0!
0%
b111 *
0-
02
b111 6
#438870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#438880000000
0!
0%
b0 *
0-
02
b0 6
#438890000000
1!
1%
1-
12
#438900000000
0!
0%
b1 *
0-
02
b1 6
#438910000000
1!
1%
1-
12
#438920000000
0!
0%
b10 *
0-
02
b10 6
#438930000000
1!
1%
1-
12
#438940000000
0!
0%
b11 *
0-
02
b11 6
#438950000000
1!
1%
1-
12
15
#438960000000
0!
0%
b100 *
0-
02
b100 6
#438970000000
1!
1%
1-
12
#438980000000
0!
0%
b101 *
0-
02
b101 6
#438990000000
1!
1%
1-
12
#439000000000
0!
0%
b110 *
0-
02
b110 6
#439010000000
1!
1%
1-
12
#439020000000
0!
0%
b111 *
0-
02
b111 6
#439030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#439040000000
0!
0%
b0 *
0-
02
b0 6
#439050000000
1!
1%
1-
12
#439060000000
0!
0%
b1 *
0-
02
b1 6
#439070000000
1!
1%
1-
12
#439080000000
0!
0%
b10 *
0-
02
b10 6
#439090000000
1!
1%
1-
12
#439100000000
0!
0%
b11 *
0-
02
b11 6
#439110000000
1!
1%
1-
12
15
#439120000000
0!
0%
b100 *
0-
02
b100 6
#439130000000
1!
1%
1-
12
#439140000000
0!
0%
b101 *
0-
02
b101 6
#439150000000
1!
1%
1-
12
#439160000000
0!
0%
b110 *
0-
02
b110 6
#439170000000
1!
1%
1-
12
#439180000000
0!
0%
b111 *
0-
02
b111 6
#439190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#439200000000
0!
0%
b0 *
0-
02
b0 6
#439210000000
1!
1%
1-
12
#439220000000
0!
0%
b1 *
0-
02
b1 6
#439230000000
1!
1%
1-
12
#439240000000
0!
0%
b10 *
0-
02
b10 6
#439250000000
1!
1%
1-
12
#439260000000
0!
0%
b11 *
0-
02
b11 6
#439270000000
1!
1%
1-
12
15
#439280000000
0!
0%
b100 *
0-
02
b100 6
#439290000000
1!
1%
1-
12
#439300000000
0!
0%
b101 *
0-
02
b101 6
#439310000000
1!
1%
1-
12
#439320000000
0!
0%
b110 *
0-
02
b110 6
#439330000000
1!
1%
1-
12
#439340000000
0!
0%
b111 *
0-
02
b111 6
#439350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#439360000000
0!
0%
b0 *
0-
02
b0 6
#439370000000
1!
1%
1-
12
#439380000000
0!
0%
b1 *
0-
02
b1 6
#439390000000
1!
1%
1-
12
#439400000000
0!
0%
b10 *
0-
02
b10 6
#439410000000
1!
1%
1-
12
#439420000000
0!
0%
b11 *
0-
02
b11 6
#439430000000
1!
1%
1-
12
15
#439440000000
0!
0%
b100 *
0-
02
b100 6
#439450000000
1!
1%
1-
12
#439460000000
0!
0%
b101 *
0-
02
b101 6
#439470000000
1!
1%
1-
12
#439480000000
0!
0%
b110 *
0-
02
b110 6
#439490000000
1!
1%
1-
12
#439500000000
0!
0%
b111 *
0-
02
b111 6
#439510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#439520000000
0!
0%
b0 *
0-
02
b0 6
#439530000000
1!
1%
1-
12
#439540000000
0!
0%
b1 *
0-
02
b1 6
#439550000000
1!
1%
1-
12
#439560000000
0!
0%
b10 *
0-
02
b10 6
#439570000000
1!
1%
1-
12
#439580000000
0!
0%
b11 *
0-
02
b11 6
#439590000000
1!
1%
1-
12
15
#439600000000
0!
0%
b100 *
0-
02
b100 6
#439610000000
1!
1%
1-
12
#439620000000
0!
0%
b101 *
0-
02
b101 6
#439630000000
1!
1%
1-
12
#439640000000
0!
0%
b110 *
0-
02
b110 6
#439650000000
1!
1%
1-
12
#439660000000
0!
0%
b111 *
0-
02
b111 6
#439670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#439680000000
0!
0%
b0 *
0-
02
b0 6
#439690000000
1!
1%
1-
12
#439700000000
0!
0%
b1 *
0-
02
b1 6
#439710000000
1!
1%
1-
12
#439720000000
0!
0%
b10 *
0-
02
b10 6
#439730000000
1!
1%
1-
12
#439740000000
0!
0%
b11 *
0-
02
b11 6
#439750000000
1!
1%
1-
12
15
#439760000000
0!
0%
b100 *
0-
02
b100 6
#439770000000
1!
1%
1-
12
#439780000000
0!
0%
b101 *
0-
02
b101 6
#439790000000
1!
1%
1-
12
#439800000000
0!
0%
b110 *
0-
02
b110 6
#439810000000
1!
1%
1-
12
#439820000000
0!
0%
b111 *
0-
02
b111 6
#439830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#439840000000
0!
0%
b0 *
0-
02
b0 6
#439850000000
1!
1%
1-
12
#439860000000
0!
0%
b1 *
0-
02
b1 6
#439870000000
1!
1%
1-
12
#439880000000
0!
0%
b10 *
0-
02
b10 6
#439890000000
1!
1%
1-
12
#439900000000
0!
0%
b11 *
0-
02
b11 6
#439910000000
1!
1%
1-
12
15
#439920000000
0!
0%
b100 *
0-
02
b100 6
#439930000000
1!
1%
1-
12
#439940000000
0!
0%
b101 *
0-
02
b101 6
#439950000000
1!
1%
1-
12
#439960000000
0!
0%
b110 *
0-
02
b110 6
#439970000000
1!
1%
1-
12
#439980000000
0!
0%
b111 *
0-
02
b111 6
#439990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#440000000000
0!
0%
b0 *
0-
02
b0 6
#440010000000
1!
1%
1-
12
#440020000000
0!
0%
b1 *
0-
02
b1 6
#440030000000
1!
1%
1-
12
#440040000000
0!
0%
b10 *
0-
02
b10 6
#440050000000
1!
1%
1-
12
#440060000000
0!
0%
b11 *
0-
02
b11 6
#440070000000
1!
1%
1-
12
15
#440080000000
0!
0%
b100 *
0-
02
b100 6
#440090000000
1!
1%
1-
12
#440100000000
0!
0%
b101 *
0-
02
b101 6
#440110000000
1!
1%
1-
12
#440120000000
0!
0%
b110 *
0-
02
b110 6
#440130000000
1!
1%
1-
12
#440140000000
0!
0%
b111 *
0-
02
b111 6
#440150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#440160000000
0!
0%
b0 *
0-
02
b0 6
#440170000000
1!
1%
1-
12
#440180000000
0!
0%
b1 *
0-
02
b1 6
#440190000000
1!
1%
1-
12
#440200000000
0!
0%
b10 *
0-
02
b10 6
#440210000000
1!
1%
1-
12
#440220000000
0!
0%
b11 *
0-
02
b11 6
#440230000000
1!
1%
1-
12
15
#440240000000
0!
0%
b100 *
0-
02
b100 6
#440250000000
1!
1%
1-
12
#440260000000
0!
0%
b101 *
0-
02
b101 6
#440270000000
1!
1%
1-
12
#440280000000
0!
0%
b110 *
0-
02
b110 6
#440290000000
1!
1%
1-
12
#440300000000
0!
0%
b111 *
0-
02
b111 6
#440310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#440320000000
0!
0%
b0 *
0-
02
b0 6
#440330000000
1!
1%
1-
12
#440340000000
0!
0%
b1 *
0-
02
b1 6
#440350000000
1!
1%
1-
12
#440360000000
0!
0%
b10 *
0-
02
b10 6
#440370000000
1!
1%
1-
12
#440380000000
0!
0%
b11 *
0-
02
b11 6
#440390000000
1!
1%
1-
12
15
#440400000000
0!
0%
b100 *
0-
02
b100 6
#440410000000
1!
1%
1-
12
#440420000000
0!
0%
b101 *
0-
02
b101 6
#440430000000
1!
1%
1-
12
#440440000000
0!
0%
b110 *
0-
02
b110 6
#440450000000
1!
1%
1-
12
#440460000000
0!
0%
b111 *
0-
02
b111 6
#440470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#440480000000
0!
0%
b0 *
0-
02
b0 6
#440490000000
1!
1%
1-
12
#440500000000
0!
0%
b1 *
0-
02
b1 6
#440510000000
1!
1%
1-
12
#440520000000
0!
0%
b10 *
0-
02
b10 6
#440530000000
1!
1%
1-
12
#440540000000
0!
0%
b11 *
0-
02
b11 6
#440550000000
1!
1%
1-
12
15
#440560000000
0!
0%
b100 *
0-
02
b100 6
#440570000000
1!
1%
1-
12
#440580000000
0!
0%
b101 *
0-
02
b101 6
#440590000000
1!
1%
1-
12
#440600000000
0!
0%
b110 *
0-
02
b110 6
#440610000000
1!
1%
1-
12
#440620000000
0!
0%
b111 *
0-
02
b111 6
#440630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#440640000000
0!
0%
b0 *
0-
02
b0 6
#440650000000
1!
1%
1-
12
#440660000000
0!
0%
b1 *
0-
02
b1 6
#440670000000
1!
1%
1-
12
#440680000000
0!
0%
b10 *
0-
02
b10 6
#440690000000
1!
1%
1-
12
#440700000000
0!
0%
b11 *
0-
02
b11 6
#440710000000
1!
1%
1-
12
15
#440720000000
0!
0%
b100 *
0-
02
b100 6
#440730000000
1!
1%
1-
12
#440740000000
0!
0%
b101 *
0-
02
b101 6
#440750000000
1!
1%
1-
12
#440760000000
0!
0%
b110 *
0-
02
b110 6
#440770000000
1!
1%
1-
12
#440780000000
0!
0%
b111 *
0-
02
b111 6
#440790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#440800000000
0!
0%
b0 *
0-
02
b0 6
#440810000000
1!
1%
1-
12
#440820000000
0!
0%
b1 *
0-
02
b1 6
#440830000000
1!
1%
1-
12
#440840000000
0!
0%
b10 *
0-
02
b10 6
#440850000000
1!
1%
1-
12
#440860000000
0!
0%
b11 *
0-
02
b11 6
#440870000000
1!
1%
1-
12
15
#440880000000
0!
0%
b100 *
0-
02
b100 6
#440890000000
1!
1%
1-
12
#440900000000
0!
0%
b101 *
0-
02
b101 6
#440910000000
1!
1%
1-
12
#440920000000
0!
0%
b110 *
0-
02
b110 6
#440930000000
1!
1%
1-
12
#440940000000
0!
0%
b111 *
0-
02
b111 6
#440950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#440960000000
0!
0%
b0 *
0-
02
b0 6
#440970000000
1!
1%
1-
12
#440980000000
0!
0%
b1 *
0-
02
b1 6
#440990000000
1!
1%
1-
12
#441000000000
0!
0%
b10 *
0-
02
b10 6
#441010000000
1!
1%
1-
12
#441020000000
0!
0%
b11 *
0-
02
b11 6
#441030000000
1!
1%
1-
12
15
#441040000000
0!
0%
b100 *
0-
02
b100 6
#441050000000
1!
1%
1-
12
#441060000000
0!
0%
b101 *
0-
02
b101 6
#441070000000
1!
1%
1-
12
#441080000000
0!
0%
b110 *
0-
02
b110 6
#441090000000
1!
1%
1-
12
#441100000000
0!
0%
b111 *
0-
02
b111 6
#441110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#441120000000
0!
0%
b0 *
0-
02
b0 6
#441130000000
1!
1%
1-
12
#441140000000
0!
0%
b1 *
0-
02
b1 6
#441150000000
1!
1%
1-
12
#441160000000
0!
0%
b10 *
0-
02
b10 6
#441170000000
1!
1%
1-
12
#441180000000
0!
0%
b11 *
0-
02
b11 6
#441190000000
1!
1%
1-
12
15
#441200000000
0!
0%
b100 *
0-
02
b100 6
#441210000000
1!
1%
1-
12
#441220000000
0!
0%
b101 *
0-
02
b101 6
#441230000000
1!
1%
1-
12
#441240000000
0!
0%
b110 *
0-
02
b110 6
#441250000000
1!
1%
1-
12
#441260000000
0!
0%
b111 *
0-
02
b111 6
#441270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#441280000000
0!
0%
b0 *
0-
02
b0 6
#441290000000
1!
1%
1-
12
#441300000000
0!
0%
b1 *
0-
02
b1 6
#441310000000
1!
1%
1-
12
#441320000000
0!
0%
b10 *
0-
02
b10 6
#441330000000
1!
1%
1-
12
#441340000000
0!
0%
b11 *
0-
02
b11 6
#441350000000
1!
1%
1-
12
15
#441360000000
0!
0%
b100 *
0-
02
b100 6
#441370000000
1!
1%
1-
12
#441380000000
0!
0%
b101 *
0-
02
b101 6
#441390000000
1!
1%
1-
12
#441400000000
0!
0%
b110 *
0-
02
b110 6
#441410000000
1!
1%
1-
12
#441420000000
0!
0%
b111 *
0-
02
b111 6
#441430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#441440000000
0!
0%
b0 *
0-
02
b0 6
#441450000000
1!
1%
1-
12
#441460000000
0!
0%
b1 *
0-
02
b1 6
#441470000000
1!
1%
1-
12
#441480000000
0!
0%
b10 *
0-
02
b10 6
#441490000000
1!
1%
1-
12
#441500000000
0!
0%
b11 *
0-
02
b11 6
#441510000000
1!
1%
1-
12
15
#441520000000
0!
0%
b100 *
0-
02
b100 6
#441530000000
1!
1%
1-
12
#441540000000
0!
0%
b101 *
0-
02
b101 6
#441550000000
1!
1%
1-
12
#441560000000
0!
0%
b110 *
0-
02
b110 6
#441570000000
1!
1%
1-
12
#441580000000
0!
0%
b111 *
0-
02
b111 6
#441590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#441600000000
0!
0%
b0 *
0-
02
b0 6
#441610000000
1!
1%
1-
12
#441620000000
0!
0%
b1 *
0-
02
b1 6
#441630000000
1!
1%
1-
12
#441640000000
0!
0%
b10 *
0-
02
b10 6
#441650000000
1!
1%
1-
12
#441660000000
0!
0%
b11 *
0-
02
b11 6
#441670000000
1!
1%
1-
12
15
#441680000000
0!
0%
b100 *
0-
02
b100 6
#441690000000
1!
1%
1-
12
#441700000000
0!
0%
b101 *
0-
02
b101 6
#441710000000
1!
1%
1-
12
#441720000000
0!
0%
b110 *
0-
02
b110 6
#441730000000
1!
1%
1-
12
#441740000000
0!
0%
b111 *
0-
02
b111 6
#441750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#441760000000
0!
0%
b0 *
0-
02
b0 6
#441770000000
1!
1%
1-
12
#441780000000
0!
0%
b1 *
0-
02
b1 6
#441790000000
1!
1%
1-
12
#441800000000
0!
0%
b10 *
0-
02
b10 6
#441810000000
1!
1%
1-
12
#441820000000
0!
0%
b11 *
0-
02
b11 6
#441830000000
1!
1%
1-
12
15
#441840000000
0!
0%
b100 *
0-
02
b100 6
#441850000000
1!
1%
1-
12
#441860000000
0!
0%
b101 *
0-
02
b101 6
#441870000000
1!
1%
1-
12
#441880000000
0!
0%
b110 *
0-
02
b110 6
#441890000000
1!
1%
1-
12
#441900000000
0!
0%
b111 *
0-
02
b111 6
#441910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#441920000000
0!
0%
b0 *
0-
02
b0 6
#441930000000
1!
1%
1-
12
#441940000000
0!
0%
b1 *
0-
02
b1 6
#441950000000
1!
1%
1-
12
#441960000000
0!
0%
b10 *
0-
02
b10 6
#441970000000
1!
1%
1-
12
#441980000000
0!
0%
b11 *
0-
02
b11 6
#441990000000
1!
1%
1-
12
15
#442000000000
0!
0%
b100 *
0-
02
b100 6
#442010000000
1!
1%
1-
12
#442020000000
0!
0%
b101 *
0-
02
b101 6
#442030000000
1!
1%
1-
12
#442040000000
0!
0%
b110 *
0-
02
b110 6
#442050000000
1!
1%
1-
12
#442060000000
0!
0%
b111 *
0-
02
b111 6
#442070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#442080000000
0!
0%
b0 *
0-
02
b0 6
#442090000000
1!
1%
1-
12
#442100000000
0!
0%
b1 *
0-
02
b1 6
#442110000000
1!
1%
1-
12
#442120000000
0!
0%
b10 *
0-
02
b10 6
#442130000000
1!
1%
1-
12
#442140000000
0!
0%
b11 *
0-
02
b11 6
#442150000000
1!
1%
1-
12
15
#442160000000
0!
0%
b100 *
0-
02
b100 6
#442170000000
1!
1%
1-
12
#442180000000
0!
0%
b101 *
0-
02
b101 6
#442190000000
1!
1%
1-
12
#442200000000
0!
0%
b110 *
0-
02
b110 6
#442210000000
1!
1%
1-
12
#442220000000
0!
0%
b111 *
0-
02
b111 6
#442230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#442240000000
0!
0%
b0 *
0-
02
b0 6
#442250000000
1!
1%
1-
12
#442260000000
0!
0%
b1 *
0-
02
b1 6
#442270000000
1!
1%
1-
12
#442280000000
0!
0%
b10 *
0-
02
b10 6
#442290000000
1!
1%
1-
12
#442300000000
0!
0%
b11 *
0-
02
b11 6
#442310000000
1!
1%
1-
12
15
#442320000000
0!
0%
b100 *
0-
02
b100 6
#442330000000
1!
1%
1-
12
#442340000000
0!
0%
b101 *
0-
02
b101 6
#442350000000
1!
1%
1-
12
#442360000000
0!
0%
b110 *
0-
02
b110 6
#442370000000
1!
1%
1-
12
#442380000000
0!
0%
b111 *
0-
02
b111 6
#442390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#442400000000
0!
0%
b0 *
0-
02
b0 6
#442410000000
1!
1%
1-
12
#442420000000
0!
0%
b1 *
0-
02
b1 6
#442430000000
1!
1%
1-
12
#442440000000
0!
0%
b10 *
0-
02
b10 6
#442450000000
1!
1%
1-
12
#442460000000
0!
0%
b11 *
0-
02
b11 6
#442470000000
1!
1%
1-
12
15
#442480000000
0!
0%
b100 *
0-
02
b100 6
#442490000000
1!
1%
1-
12
#442500000000
0!
0%
b101 *
0-
02
b101 6
#442510000000
1!
1%
1-
12
#442520000000
0!
0%
b110 *
0-
02
b110 6
#442530000000
1!
1%
1-
12
#442540000000
0!
0%
b111 *
0-
02
b111 6
#442550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#442560000000
0!
0%
b0 *
0-
02
b0 6
#442570000000
1!
1%
1-
12
#442580000000
0!
0%
b1 *
0-
02
b1 6
#442590000000
1!
1%
1-
12
#442600000000
0!
0%
b10 *
0-
02
b10 6
#442610000000
1!
1%
1-
12
#442620000000
0!
0%
b11 *
0-
02
b11 6
#442630000000
1!
1%
1-
12
15
#442640000000
0!
0%
b100 *
0-
02
b100 6
#442650000000
1!
1%
1-
12
#442660000000
0!
0%
b101 *
0-
02
b101 6
#442670000000
1!
1%
1-
12
#442680000000
0!
0%
b110 *
0-
02
b110 6
#442690000000
1!
1%
1-
12
#442700000000
0!
0%
b111 *
0-
02
b111 6
#442710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#442720000000
0!
0%
b0 *
0-
02
b0 6
#442730000000
1!
1%
1-
12
#442740000000
0!
0%
b1 *
0-
02
b1 6
#442750000000
1!
1%
1-
12
#442760000000
0!
0%
b10 *
0-
02
b10 6
#442770000000
1!
1%
1-
12
#442780000000
0!
0%
b11 *
0-
02
b11 6
#442790000000
1!
1%
1-
12
15
#442800000000
0!
0%
b100 *
0-
02
b100 6
#442810000000
1!
1%
1-
12
#442820000000
0!
0%
b101 *
0-
02
b101 6
#442830000000
1!
1%
1-
12
#442840000000
0!
0%
b110 *
0-
02
b110 6
#442850000000
1!
1%
1-
12
#442860000000
0!
0%
b111 *
0-
02
b111 6
#442870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#442880000000
0!
0%
b0 *
0-
02
b0 6
#442890000000
1!
1%
1-
12
#442900000000
0!
0%
b1 *
0-
02
b1 6
#442910000000
1!
1%
1-
12
#442920000000
0!
0%
b10 *
0-
02
b10 6
#442930000000
1!
1%
1-
12
#442940000000
0!
0%
b11 *
0-
02
b11 6
#442950000000
1!
1%
1-
12
15
#442960000000
0!
0%
b100 *
0-
02
b100 6
#442970000000
1!
1%
1-
12
#442980000000
0!
0%
b101 *
0-
02
b101 6
#442990000000
1!
1%
1-
12
#443000000000
0!
0%
b110 *
0-
02
b110 6
#443010000000
1!
1%
1-
12
#443020000000
0!
0%
b111 *
0-
02
b111 6
#443030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#443040000000
0!
0%
b0 *
0-
02
b0 6
#443050000000
1!
1%
1-
12
#443060000000
0!
0%
b1 *
0-
02
b1 6
#443070000000
1!
1%
1-
12
#443080000000
0!
0%
b10 *
0-
02
b10 6
#443090000000
1!
1%
1-
12
#443100000000
0!
0%
b11 *
0-
02
b11 6
#443110000000
1!
1%
1-
12
15
#443120000000
0!
0%
b100 *
0-
02
b100 6
#443130000000
1!
1%
1-
12
#443140000000
0!
0%
b101 *
0-
02
b101 6
#443150000000
1!
1%
1-
12
#443160000000
0!
0%
b110 *
0-
02
b110 6
#443170000000
1!
1%
1-
12
#443180000000
0!
0%
b111 *
0-
02
b111 6
#443190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#443200000000
0!
0%
b0 *
0-
02
b0 6
#443210000000
1!
1%
1-
12
#443220000000
0!
0%
b1 *
0-
02
b1 6
#443230000000
1!
1%
1-
12
#443240000000
0!
0%
b10 *
0-
02
b10 6
#443250000000
1!
1%
1-
12
#443260000000
0!
0%
b11 *
0-
02
b11 6
#443270000000
1!
1%
1-
12
15
#443280000000
0!
0%
b100 *
0-
02
b100 6
#443290000000
1!
1%
1-
12
#443300000000
0!
0%
b101 *
0-
02
b101 6
#443310000000
1!
1%
1-
12
#443320000000
0!
0%
b110 *
0-
02
b110 6
#443330000000
1!
1%
1-
12
#443340000000
0!
0%
b111 *
0-
02
b111 6
#443350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#443360000000
0!
0%
b0 *
0-
02
b0 6
#443370000000
1!
1%
1-
12
#443380000000
0!
0%
b1 *
0-
02
b1 6
#443390000000
1!
1%
1-
12
#443400000000
0!
0%
b10 *
0-
02
b10 6
#443410000000
1!
1%
1-
12
#443420000000
0!
0%
b11 *
0-
02
b11 6
#443430000000
1!
1%
1-
12
15
#443440000000
0!
0%
b100 *
0-
02
b100 6
#443450000000
1!
1%
1-
12
#443460000000
0!
0%
b101 *
0-
02
b101 6
#443470000000
1!
1%
1-
12
#443480000000
0!
0%
b110 *
0-
02
b110 6
#443490000000
1!
1%
1-
12
#443500000000
0!
0%
b111 *
0-
02
b111 6
#443510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#443520000000
0!
0%
b0 *
0-
02
b0 6
#443530000000
1!
1%
1-
12
#443540000000
0!
0%
b1 *
0-
02
b1 6
#443550000000
1!
1%
1-
12
#443560000000
0!
0%
b10 *
0-
02
b10 6
#443570000000
1!
1%
1-
12
#443580000000
0!
0%
b11 *
0-
02
b11 6
#443590000000
1!
1%
1-
12
15
#443600000000
0!
0%
b100 *
0-
02
b100 6
#443610000000
1!
1%
1-
12
#443620000000
0!
0%
b101 *
0-
02
b101 6
#443630000000
1!
1%
1-
12
#443640000000
0!
0%
b110 *
0-
02
b110 6
#443650000000
1!
1%
1-
12
#443660000000
0!
0%
b111 *
0-
02
b111 6
#443670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#443680000000
0!
0%
b0 *
0-
02
b0 6
#443690000000
1!
1%
1-
12
#443700000000
0!
0%
b1 *
0-
02
b1 6
#443710000000
1!
1%
1-
12
#443720000000
0!
0%
b10 *
0-
02
b10 6
#443730000000
1!
1%
1-
12
#443740000000
0!
0%
b11 *
0-
02
b11 6
#443750000000
1!
1%
1-
12
15
#443760000000
0!
0%
b100 *
0-
02
b100 6
#443770000000
1!
1%
1-
12
#443780000000
0!
0%
b101 *
0-
02
b101 6
#443790000000
1!
1%
1-
12
#443800000000
0!
0%
b110 *
0-
02
b110 6
#443810000000
1!
1%
1-
12
#443820000000
0!
0%
b111 *
0-
02
b111 6
#443830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#443840000000
0!
0%
b0 *
0-
02
b0 6
#443850000000
1!
1%
1-
12
#443860000000
0!
0%
b1 *
0-
02
b1 6
#443870000000
1!
1%
1-
12
#443880000000
0!
0%
b10 *
0-
02
b10 6
#443890000000
1!
1%
1-
12
#443900000000
0!
0%
b11 *
0-
02
b11 6
#443910000000
1!
1%
1-
12
15
#443920000000
0!
0%
b100 *
0-
02
b100 6
#443930000000
1!
1%
1-
12
#443940000000
0!
0%
b101 *
0-
02
b101 6
#443950000000
1!
1%
1-
12
#443960000000
0!
0%
b110 *
0-
02
b110 6
#443970000000
1!
1%
1-
12
#443980000000
0!
0%
b111 *
0-
02
b111 6
#443990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#444000000000
0!
0%
b0 *
0-
02
b0 6
#444010000000
1!
1%
1-
12
#444020000000
0!
0%
b1 *
0-
02
b1 6
#444030000000
1!
1%
1-
12
#444040000000
0!
0%
b10 *
0-
02
b10 6
#444050000000
1!
1%
1-
12
#444060000000
0!
0%
b11 *
0-
02
b11 6
#444070000000
1!
1%
1-
12
15
#444080000000
0!
0%
b100 *
0-
02
b100 6
#444090000000
1!
1%
1-
12
#444100000000
0!
0%
b101 *
0-
02
b101 6
#444110000000
1!
1%
1-
12
#444120000000
0!
0%
b110 *
0-
02
b110 6
#444130000000
1!
1%
1-
12
#444140000000
0!
0%
b111 *
0-
02
b111 6
#444150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#444160000000
0!
0%
b0 *
0-
02
b0 6
#444170000000
1!
1%
1-
12
#444180000000
0!
0%
b1 *
0-
02
b1 6
#444190000000
1!
1%
1-
12
#444200000000
0!
0%
b10 *
0-
02
b10 6
#444210000000
1!
1%
1-
12
#444220000000
0!
0%
b11 *
0-
02
b11 6
#444230000000
1!
1%
1-
12
15
#444240000000
0!
0%
b100 *
0-
02
b100 6
#444250000000
1!
1%
1-
12
#444260000000
0!
0%
b101 *
0-
02
b101 6
#444270000000
1!
1%
1-
12
#444280000000
0!
0%
b110 *
0-
02
b110 6
#444290000000
1!
1%
1-
12
#444300000000
0!
0%
b111 *
0-
02
b111 6
#444310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#444320000000
0!
0%
b0 *
0-
02
b0 6
#444330000000
1!
1%
1-
12
#444340000000
0!
0%
b1 *
0-
02
b1 6
#444350000000
1!
1%
1-
12
#444360000000
0!
0%
b10 *
0-
02
b10 6
#444370000000
1!
1%
1-
12
#444380000000
0!
0%
b11 *
0-
02
b11 6
#444390000000
1!
1%
1-
12
15
#444400000000
0!
0%
b100 *
0-
02
b100 6
#444410000000
1!
1%
1-
12
#444420000000
0!
0%
b101 *
0-
02
b101 6
#444430000000
1!
1%
1-
12
#444440000000
0!
0%
b110 *
0-
02
b110 6
#444450000000
1!
1%
1-
12
#444460000000
0!
0%
b111 *
0-
02
b111 6
#444470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#444480000000
0!
0%
b0 *
0-
02
b0 6
#444490000000
1!
1%
1-
12
#444500000000
0!
0%
b1 *
0-
02
b1 6
#444510000000
1!
1%
1-
12
#444520000000
0!
0%
b10 *
0-
02
b10 6
#444530000000
1!
1%
1-
12
#444540000000
0!
0%
b11 *
0-
02
b11 6
#444550000000
1!
1%
1-
12
15
#444560000000
0!
0%
b100 *
0-
02
b100 6
#444570000000
1!
1%
1-
12
#444580000000
0!
0%
b101 *
0-
02
b101 6
#444590000000
1!
1%
1-
12
#444600000000
0!
0%
b110 *
0-
02
b110 6
#444610000000
1!
1%
1-
12
#444620000000
0!
0%
b111 *
0-
02
b111 6
#444630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#444640000000
0!
0%
b0 *
0-
02
b0 6
#444650000000
1!
1%
1-
12
#444660000000
0!
0%
b1 *
0-
02
b1 6
#444670000000
1!
1%
1-
12
#444680000000
0!
0%
b10 *
0-
02
b10 6
#444690000000
1!
1%
1-
12
#444700000000
0!
0%
b11 *
0-
02
b11 6
#444710000000
1!
1%
1-
12
15
#444720000000
0!
0%
b100 *
0-
02
b100 6
#444730000000
1!
1%
1-
12
#444740000000
0!
0%
b101 *
0-
02
b101 6
#444750000000
1!
1%
1-
12
#444760000000
0!
0%
b110 *
0-
02
b110 6
#444770000000
1!
1%
1-
12
#444780000000
0!
0%
b111 *
0-
02
b111 6
#444790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#444800000000
0!
0%
b0 *
0-
02
b0 6
#444810000000
1!
1%
1-
12
#444820000000
0!
0%
b1 *
0-
02
b1 6
#444830000000
1!
1%
1-
12
#444840000000
0!
0%
b10 *
0-
02
b10 6
#444850000000
1!
1%
1-
12
#444860000000
0!
0%
b11 *
0-
02
b11 6
#444870000000
1!
1%
1-
12
15
#444880000000
0!
0%
b100 *
0-
02
b100 6
#444890000000
1!
1%
1-
12
#444900000000
0!
0%
b101 *
0-
02
b101 6
#444910000000
1!
1%
1-
12
#444920000000
0!
0%
b110 *
0-
02
b110 6
#444930000000
1!
1%
1-
12
#444940000000
0!
0%
b111 *
0-
02
b111 6
#444950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#444960000000
0!
0%
b0 *
0-
02
b0 6
#444970000000
1!
1%
1-
12
#444980000000
0!
0%
b1 *
0-
02
b1 6
#444990000000
1!
1%
1-
12
#445000000000
0!
0%
b10 *
0-
02
b10 6
#445010000000
1!
1%
1-
12
#445020000000
0!
0%
b11 *
0-
02
b11 6
#445030000000
1!
1%
1-
12
15
#445040000000
0!
0%
b100 *
0-
02
b100 6
#445050000000
1!
1%
1-
12
#445060000000
0!
0%
b101 *
0-
02
b101 6
#445070000000
1!
1%
1-
12
#445080000000
0!
0%
b110 *
0-
02
b110 6
#445090000000
1!
1%
1-
12
#445100000000
0!
0%
b111 *
0-
02
b111 6
#445110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#445120000000
0!
0%
b0 *
0-
02
b0 6
#445130000000
1!
1%
1-
12
#445140000000
0!
0%
b1 *
0-
02
b1 6
#445150000000
1!
1%
1-
12
#445160000000
0!
0%
b10 *
0-
02
b10 6
#445170000000
1!
1%
1-
12
#445180000000
0!
0%
b11 *
0-
02
b11 6
#445190000000
1!
1%
1-
12
15
#445200000000
0!
0%
b100 *
0-
02
b100 6
#445210000000
1!
1%
1-
12
#445220000000
0!
0%
b101 *
0-
02
b101 6
#445230000000
1!
1%
1-
12
#445240000000
0!
0%
b110 *
0-
02
b110 6
#445250000000
1!
1%
1-
12
#445260000000
0!
0%
b111 *
0-
02
b111 6
#445270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#445280000000
0!
0%
b0 *
0-
02
b0 6
#445290000000
1!
1%
1-
12
#445300000000
0!
0%
b1 *
0-
02
b1 6
#445310000000
1!
1%
1-
12
#445320000000
0!
0%
b10 *
0-
02
b10 6
#445330000000
1!
1%
1-
12
#445340000000
0!
0%
b11 *
0-
02
b11 6
#445350000000
1!
1%
1-
12
15
#445360000000
0!
0%
b100 *
0-
02
b100 6
#445370000000
1!
1%
1-
12
#445380000000
0!
0%
b101 *
0-
02
b101 6
#445390000000
1!
1%
1-
12
#445400000000
0!
0%
b110 *
0-
02
b110 6
#445410000000
1!
1%
1-
12
#445420000000
0!
0%
b111 *
0-
02
b111 6
#445430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#445440000000
0!
0%
b0 *
0-
02
b0 6
#445450000000
1!
1%
1-
12
#445460000000
0!
0%
b1 *
0-
02
b1 6
#445470000000
1!
1%
1-
12
#445480000000
0!
0%
b10 *
0-
02
b10 6
#445490000000
1!
1%
1-
12
#445500000000
0!
0%
b11 *
0-
02
b11 6
#445510000000
1!
1%
1-
12
15
#445520000000
0!
0%
b100 *
0-
02
b100 6
#445530000000
1!
1%
1-
12
#445540000000
0!
0%
b101 *
0-
02
b101 6
#445550000000
1!
1%
1-
12
#445560000000
0!
0%
b110 *
0-
02
b110 6
#445570000000
1!
1%
1-
12
#445580000000
0!
0%
b111 *
0-
02
b111 6
#445590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#445600000000
0!
0%
b0 *
0-
02
b0 6
#445610000000
1!
1%
1-
12
#445620000000
0!
0%
b1 *
0-
02
b1 6
#445630000000
1!
1%
1-
12
#445640000000
0!
0%
b10 *
0-
02
b10 6
#445650000000
1!
1%
1-
12
#445660000000
0!
0%
b11 *
0-
02
b11 6
#445670000000
1!
1%
1-
12
15
#445680000000
0!
0%
b100 *
0-
02
b100 6
#445690000000
1!
1%
1-
12
#445700000000
0!
0%
b101 *
0-
02
b101 6
#445710000000
1!
1%
1-
12
#445720000000
0!
0%
b110 *
0-
02
b110 6
#445730000000
1!
1%
1-
12
#445740000000
0!
0%
b111 *
0-
02
b111 6
#445750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#445760000000
0!
0%
b0 *
0-
02
b0 6
#445770000000
1!
1%
1-
12
#445780000000
0!
0%
b1 *
0-
02
b1 6
#445790000000
1!
1%
1-
12
#445800000000
0!
0%
b10 *
0-
02
b10 6
#445810000000
1!
1%
1-
12
#445820000000
0!
0%
b11 *
0-
02
b11 6
#445830000000
1!
1%
1-
12
15
#445840000000
0!
0%
b100 *
0-
02
b100 6
#445850000000
1!
1%
1-
12
#445860000000
0!
0%
b101 *
0-
02
b101 6
#445870000000
1!
1%
1-
12
#445880000000
0!
0%
b110 *
0-
02
b110 6
#445890000000
1!
1%
1-
12
#445900000000
0!
0%
b111 *
0-
02
b111 6
#445910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#445920000000
0!
0%
b0 *
0-
02
b0 6
#445930000000
1!
1%
1-
12
#445940000000
0!
0%
b1 *
0-
02
b1 6
#445950000000
1!
1%
1-
12
#445960000000
0!
0%
b10 *
0-
02
b10 6
#445970000000
1!
1%
1-
12
#445980000000
0!
0%
b11 *
0-
02
b11 6
#445990000000
1!
1%
1-
12
15
#446000000000
0!
0%
b100 *
0-
02
b100 6
#446010000000
1!
1%
1-
12
#446020000000
0!
0%
b101 *
0-
02
b101 6
#446030000000
1!
1%
1-
12
#446040000000
0!
0%
b110 *
0-
02
b110 6
#446050000000
1!
1%
1-
12
#446060000000
0!
0%
b111 *
0-
02
b111 6
#446070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#446080000000
0!
0%
b0 *
0-
02
b0 6
#446090000000
1!
1%
1-
12
#446100000000
0!
0%
b1 *
0-
02
b1 6
#446110000000
1!
1%
1-
12
#446120000000
0!
0%
b10 *
0-
02
b10 6
#446130000000
1!
1%
1-
12
#446140000000
0!
0%
b11 *
0-
02
b11 6
#446150000000
1!
1%
1-
12
15
#446160000000
0!
0%
b100 *
0-
02
b100 6
#446170000000
1!
1%
1-
12
#446180000000
0!
0%
b101 *
0-
02
b101 6
#446190000000
1!
1%
1-
12
#446200000000
0!
0%
b110 *
0-
02
b110 6
#446210000000
1!
1%
1-
12
#446220000000
0!
0%
b111 *
0-
02
b111 6
#446230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#446240000000
0!
0%
b0 *
0-
02
b0 6
#446250000000
1!
1%
1-
12
#446260000000
0!
0%
b1 *
0-
02
b1 6
#446270000000
1!
1%
1-
12
#446280000000
0!
0%
b10 *
0-
02
b10 6
#446290000000
1!
1%
1-
12
#446300000000
0!
0%
b11 *
0-
02
b11 6
#446310000000
1!
1%
1-
12
15
#446320000000
0!
0%
b100 *
0-
02
b100 6
#446330000000
1!
1%
1-
12
#446340000000
0!
0%
b101 *
0-
02
b101 6
#446350000000
1!
1%
1-
12
#446360000000
0!
0%
b110 *
0-
02
b110 6
#446370000000
1!
1%
1-
12
#446380000000
0!
0%
b111 *
0-
02
b111 6
#446390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#446400000000
0!
0%
b0 *
0-
02
b0 6
#446410000000
1!
1%
1-
12
#446420000000
0!
0%
b1 *
0-
02
b1 6
#446430000000
1!
1%
1-
12
#446440000000
0!
0%
b10 *
0-
02
b10 6
#446450000000
1!
1%
1-
12
#446460000000
0!
0%
b11 *
0-
02
b11 6
#446470000000
1!
1%
1-
12
15
#446480000000
0!
0%
b100 *
0-
02
b100 6
#446490000000
1!
1%
1-
12
#446500000000
0!
0%
b101 *
0-
02
b101 6
#446510000000
1!
1%
1-
12
#446520000000
0!
0%
b110 *
0-
02
b110 6
#446530000000
1!
1%
1-
12
#446540000000
0!
0%
b111 *
0-
02
b111 6
#446550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#446560000000
0!
0%
b0 *
0-
02
b0 6
#446570000000
1!
1%
1-
12
#446580000000
0!
0%
b1 *
0-
02
b1 6
#446590000000
1!
1%
1-
12
#446600000000
0!
0%
b10 *
0-
02
b10 6
#446610000000
1!
1%
1-
12
#446620000000
0!
0%
b11 *
0-
02
b11 6
#446630000000
1!
1%
1-
12
15
#446640000000
0!
0%
b100 *
0-
02
b100 6
#446650000000
1!
1%
1-
12
#446660000000
0!
0%
b101 *
0-
02
b101 6
#446670000000
1!
1%
1-
12
#446680000000
0!
0%
b110 *
0-
02
b110 6
#446690000000
1!
1%
1-
12
#446700000000
0!
0%
b111 *
0-
02
b111 6
#446710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#446720000000
0!
0%
b0 *
0-
02
b0 6
#446730000000
1!
1%
1-
12
#446740000000
0!
0%
b1 *
0-
02
b1 6
#446750000000
1!
1%
1-
12
#446760000000
0!
0%
b10 *
0-
02
b10 6
#446770000000
1!
1%
1-
12
#446780000000
0!
0%
b11 *
0-
02
b11 6
#446790000000
1!
1%
1-
12
15
#446800000000
0!
0%
b100 *
0-
02
b100 6
#446810000000
1!
1%
1-
12
#446820000000
0!
0%
b101 *
0-
02
b101 6
#446830000000
1!
1%
1-
12
#446840000000
0!
0%
b110 *
0-
02
b110 6
#446850000000
1!
1%
1-
12
#446860000000
0!
0%
b111 *
0-
02
b111 6
#446870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#446880000000
0!
0%
b0 *
0-
02
b0 6
#446890000000
1!
1%
1-
12
#446900000000
0!
0%
b1 *
0-
02
b1 6
#446910000000
1!
1%
1-
12
#446920000000
0!
0%
b10 *
0-
02
b10 6
#446930000000
1!
1%
1-
12
#446940000000
0!
0%
b11 *
0-
02
b11 6
#446950000000
1!
1%
1-
12
15
#446960000000
0!
0%
b100 *
0-
02
b100 6
#446970000000
1!
1%
1-
12
#446980000000
0!
0%
b101 *
0-
02
b101 6
#446990000000
1!
1%
1-
12
#447000000000
0!
0%
b110 *
0-
02
b110 6
#447010000000
1!
1%
1-
12
#447020000000
0!
0%
b111 *
0-
02
b111 6
#447030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#447040000000
0!
0%
b0 *
0-
02
b0 6
#447050000000
1!
1%
1-
12
#447060000000
0!
0%
b1 *
0-
02
b1 6
#447070000000
1!
1%
1-
12
#447080000000
0!
0%
b10 *
0-
02
b10 6
#447090000000
1!
1%
1-
12
#447100000000
0!
0%
b11 *
0-
02
b11 6
#447110000000
1!
1%
1-
12
15
#447120000000
0!
0%
b100 *
0-
02
b100 6
#447130000000
1!
1%
1-
12
#447140000000
0!
0%
b101 *
0-
02
b101 6
#447150000000
1!
1%
1-
12
#447160000000
0!
0%
b110 *
0-
02
b110 6
#447170000000
1!
1%
1-
12
#447180000000
0!
0%
b111 *
0-
02
b111 6
#447190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#447200000000
0!
0%
b0 *
0-
02
b0 6
#447210000000
1!
1%
1-
12
#447220000000
0!
0%
b1 *
0-
02
b1 6
#447230000000
1!
1%
1-
12
#447240000000
0!
0%
b10 *
0-
02
b10 6
#447250000000
1!
1%
1-
12
#447260000000
0!
0%
b11 *
0-
02
b11 6
#447270000000
1!
1%
1-
12
15
#447280000000
0!
0%
b100 *
0-
02
b100 6
#447290000000
1!
1%
1-
12
#447300000000
0!
0%
b101 *
0-
02
b101 6
#447310000000
1!
1%
1-
12
#447320000000
0!
0%
b110 *
0-
02
b110 6
#447330000000
1!
1%
1-
12
#447340000000
0!
0%
b111 *
0-
02
b111 6
#447350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#447360000000
0!
0%
b0 *
0-
02
b0 6
#447370000000
1!
1%
1-
12
#447380000000
0!
0%
b1 *
0-
02
b1 6
#447390000000
1!
1%
1-
12
#447400000000
0!
0%
b10 *
0-
02
b10 6
#447410000000
1!
1%
1-
12
#447420000000
0!
0%
b11 *
0-
02
b11 6
#447430000000
1!
1%
1-
12
15
#447440000000
0!
0%
b100 *
0-
02
b100 6
#447450000000
1!
1%
1-
12
#447460000000
0!
0%
b101 *
0-
02
b101 6
#447470000000
1!
1%
1-
12
#447480000000
0!
0%
b110 *
0-
02
b110 6
#447490000000
1!
1%
1-
12
#447500000000
0!
0%
b111 *
0-
02
b111 6
#447510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#447520000000
0!
0%
b0 *
0-
02
b0 6
#447530000000
1!
1%
1-
12
#447540000000
0!
0%
b1 *
0-
02
b1 6
#447550000000
1!
1%
1-
12
#447560000000
0!
0%
b10 *
0-
02
b10 6
#447570000000
1!
1%
1-
12
#447580000000
0!
0%
b11 *
0-
02
b11 6
#447590000000
1!
1%
1-
12
15
#447600000000
0!
0%
b100 *
0-
02
b100 6
#447610000000
1!
1%
1-
12
#447620000000
0!
0%
b101 *
0-
02
b101 6
#447630000000
1!
1%
1-
12
#447640000000
0!
0%
b110 *
0-
02
b110 6
#447650000000
1!
1%
1-
12
#447660000000
0!
0%
b111 *
0-
02
b111 6
#447670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#447680000000
0!
0%
b0 *
0-
02
b0 6
#447690000000
1!
1%
1-
12
#447700000000
0!
0%
b1 *
0-
02
b1 6
#447710000000
1!
1%
1-
12
#447720000000
0!
0%
b10 *
0-
02
b10 6
#447730000000
1!
1%
1-
12
#447740000000
0!
0%
b11 *
0-
02
b11 6
#447750000000
1!
1%
1-
12
15
#447760000000
0!
0%
b100 *
0-
02
b100 6
#447770000000
1!
1%
1-
12
#447780000000
0!
0%
b101 *
0-
02
b101 6
#447790000000
1!
1%
1-
12
#447800000000
0!
0%
b110 *
0-
02
b110 6
#447810000000
1!
1%
1-
12
#447820000000
0!
0%
b111 *
0-
02
b111 6
#447830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#447840000000
0!
0%
b0 *
0-
02
b0 6
#447850000000
1!
1%
1-
12
#447860000000
0!
0%
b1 *
0-
02
b1 6
#447870000000
1!
1%
1-
12
#447880000000
0!
0%
b10 *
0-
02
b10 6
#447890000000
1!
1%
1-
12
#447900000000
0!
0%
b11 *
0-
02
b11 6
#447910000000
1!
1%
1-
12
15
#447920000000
0!
0%
b100 *
0-
02
b100 6
#447930000000
1!
1%
1-
12
#447940000000
0!
0%
b101 *
0-
02
b101 6
#447950000000
1!
1%
1-
12
#447960000000
0!
0%
b110 *
0-
02
b110 6
#447970000000
1!
1%
1-
12
#447980000000
0!
0%
b111 *
0-
02
b111 6
#447990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#448000000000
0!
0%
b0 *
0-
02
b0 6
#448010000000
1!
1%
1-
12
#448020000000
0!
0%
b1 *
0-
02
b1 6
#448030000000
1!
1%
1-
12
#448040000000
0!
0%
b10 *
0-
02
b10 6
#448050000000
1!
1%
1-
12
#448060000000
0!
0%
b11 *
0-
02
b11 6
#448070000000
1!
1%
1-
12
15
#448080000000
0!
0%
b100 *
0-
02
b100 6
#448090000000
1!
1%
1-
12
#448100000000
0!
0%
b101 *
0-
02
b101 6
#448110000000
1!
1%
1-
12
#448120000000
0!
0%
b110 *
0-
02
b110 6
#448130000000
1!
1%
1-
12
#448140000000
0!
0%
b111 *
0-
02
b111 6
#448150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#448160000000
0!
0%
b0 *
0-
02
b0 6
#448170000000
1!
1%
1-
12
#448180000000
0!
0%
b1 *
0-
02
b1 6
#448190000000
1!
1%
1-
12
#448200000000
0!
0%
b10 *
0-
02
b10 6
#448210000000
1!
1%
1-
12
#448220000000
0!
0%
b11 *
0-
02
b11 6
#448230000000
1!
1%
1-
12
15
#448240000000
0!
0%
b100 *
0-
02
b100 6
#448250000000
1!
1%
1-
12
#448260000000
0!
0%
b101 *
0-
02
b101 6
#448270000000
1!
1%
1-
12
#448280000000
0!
0%
b110 *
0-
02
b110 6
#448290000000
1!
1%
1-
12
#448300000000
0!
0%
b111 *
0-
02
b111 6
#448310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#448320000000
0!
0%
b0 *
0-
02
b0 6
#448330000000
1!
1%
1-
12
#448340000000
0!
0%
b1 *
0-
02
b1 6
#448350000000
1!
1%
1-
12
#448360000000
0!
0%
b10 *
0-
02
b10 6
#448370000000
1!
1%
1-
12
#448380000000
0!
0%
b11 *
0-
02
b11 6
#448390000000
1!
1%
1-
12
15
#448400000000
0!
0%
b100 *
0-
02
b100 6
#448410000000
1!
1%
1-
12
#448420000000
0!
0%
b101 *
0-
02
b101 6
#448430000000
1!
1%
1-
12
#448440000000
0!
0%
b110 *
0-
02
b110 6
#448450000000
1!
1%
1-
12
#448460000000
0!
0%
b111 *
0-
02
b111 6
#448470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#448480000000
0!
0%
b0 *
0-
02
b0 6
#448490000000
1!
1%
1-
12
#448500000000
0!
0%
b1 *
0-
02
b1 6
#448510000000
1!
1%
1-
12
#448520000000
0!
0%
b10 *
0-
02
b10 6
#448530000000
1!
1%
1-
12
#448540000000
0!
0%
b11 *
0-
02
b11 6
#448550000000
1!
1%
1-
12
15
#448560000000
0!
0%
b100 *
0-
02
b100 6
#448570000000
1!
1%
1-
12
#448580000000
0!
0%
b101 *
0-
02
b101 6
#448590000000
1!
1%
1-
12
#448600000000
0!
0%
b110 *
0-
02
b110 6
#448610000000
1!
1%
1-
12
#448620000000
0!
0%
b111 *
0-
02
b111 6
#448630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#448640000000
0!
0%
b0 *
0-
02
b0 6
#448650000000
1!
1%
1-
12
#448660000000
0!
0%
b1 *
0-
02
b1 6
#448670000000
1!
1%
1-
12
#448680000000
0!
0%
b10 *
0-
02
b10 6
#448690000000
1!
1%
1-
12
#448700000000
0!
0%
b11 *
0-
02
b11 6
#448710000000
1!
1%
1-
12
15
#448720000000
0!
0%
b100 *
0-
02
b100 6
#448730000000
1!
1%
1-
12
#448740000000
0!
0%
b101 *
0-
02
b101 6
#448750000000
1!
1%
1-
12
#448760000000
0!
0%
b110 *
0-
02
b110 6
#448770000000
1!
1%
1-
12
#448780000000
0!
0%
b111 *
0-
02
b111 6
#448790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#448800000000
0!
0%
b0 *
0-
02
b0 6
#448810000000
1!
1%
1-
12
#448820000000
0!
0%
b1 *
0-
02
b1 6
#448830000000
1!
1%
1-
12
#448840000000
0!
0%
b10 *
0-
02
b10 6
#448850000000
1!
1%
1-
12
#448860000000
0!
0%
b11 *
0-
02
b11 6
#448870000000
1!
1%
1-
12
15
#448880000000
0!
0%
b100 *
0-
02
b100 6
#448890000000
1!
1%
1-
12
#448900000000
0!
0%
b101 *
0-
02
b101 6
#448910000000
1!
1%
1-
12
#448920000000
0!
0%
b110 *
0-
02
b110 6
#448930000000
1!
1%
1-
12
#448940000000
0!
0%
b111 *
0-
02
b111 6
#448950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#448960000000
0!
0%
b0 *
0-
02
b0 6
#448970000000
1!
1%
1-
12
#448980000000
0!
0%
b1 *
0-
02
b1 6
#448990000000
1!
1%
1-
12
#449000000000
0!
0%
b10 *
0-
02
b10 6
#449010000000
1!
1%
1-
12
#449020000000
0!
0%
b11 *
0-
02
b11 6
#449030000000
1!
1%
1-
12
15
#449040000000
0!
0%
b100 *
0-
02
b100 6
#449050000000
1!
1%
1-
12
#449060000000
0!
0%
b101 *
0-
02
b101 6
#449070000000
1!
1%
1-
12
#449080000000
0!
0%
b110 *
0-
02
b110 6
#449090000000
1!
1%
1-
12
#449100000000
0!
0%
b111 *
0-
02
b111 6
#449110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#449120000000
0!
0%
b0 *
0-
02
b0 6
#449130000000
1!
1%
1-
12
#449140000000
0!
0%
b1 *
0-
02
b1 6
#449150000000
1!
1%
1-
12
#449160000000
0!
0%
b10 *
0-
02
b10 6
#449170000000
1!
1%
1-
12
#449180000000
0!
0%
b11 *
0-
02
b11 6
#449190000000
1!
1%
1-
12
15
#449200000000
0!
0%
b100 *
0-
02
b100 6
#449210000000
1!
1%
1-
12
#449220000000
0!
0%
b101 *
0-
02
b101 6
#449230000000
1!
1%
1-
12
#449240000000
0!
0%
b110 *
0-
02
b110 6
#449250000000
1!
1%
1-
12
#449260000000
0!
0%
b111 *
0-
02
b111 6
#449270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#449280000000
0!
0%
b0 *
0-
02
b0 6
#449290000000
1!
1%
1-
12
#449300000000
0!
0%
b1 *
0-
02
b1 6
#449310000000
1!
1%
1-
12
#449320000000
0!
0%
b10 *
0-
02
b10 6
#449330000000
1!
1%
1-
12
#449340000000
0!
0%
b11 *
0-
02
b11 6
#449350000000
1!
1%
1-
12
15
#449360000000
0!
0%
b100 *
0-
02
b100 6
#449370000000
1!
1%
1-
12
#449380000000
0!
0%
b101 *
0-
02
b101 6
#449390000000
1!
1%
1-
12
#449400000000
0!
0%
b110 *
0-
02
b110 6
#449410000000
1!
1%
1-
12
#449420000000
0!
0%
b111 *
0-
02
b111 6
#449430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#449440000000
0!
0%
b0 *
0-
02
b0 6
#449450000000
1!
1%
1-
12
#449460000000
0!
0%
b1 *
0-
02
b1 6
#449470000000
1!
1%
1-
12
#449480000000
0!
0%
b10 *
0-
02
b10 6
#449490000000
1!
1%
1-
12
#449500000000
0!
0%
b11 *
0-
02
b11 6
#449510000000
1!
1%
1-
12
15
#449520000000
0!
0%
b100 *
0-
02
b100 6
#449530000000
1!
1%
1-
12
#449540000000
0!
0%
b101 *
0-
02
b101 6
#449550000000
1!
1%
1-
12
#449560000000
0!
0%
b110 *
0-
02
b110 6
#449570000000
1!
1%
1-
12
#449580000000
0!
0%
b111 *
0-
02
b111 6
#449590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#449600000000
0!
0%
b0 *
0-
02
b0 6
#449610000000
1!
1%
1-
12
#449620000000
0!
0%
b1 *
0-
02
b1 6
#449630000000
1!
1%
1-
12
#449640000000
0!
0%
b10 *
0-
02
b10 6
#449650000000
1!
1%
1-
12
#449660000000
0!
0%
b11 *
0-
02
b11 6
#449670000000
1!
1%
1-
12
15
#449680000000
0!
0%
b100 *
0-
02
b100 6
#449690000000
1!
1%
1-
12
#449700000000
0!
0%
b101 *
0-
02
b101 6
#449710000000
1!
1%
1-
12
#449720000000
0!
0%
b110 *
0-
02
b110 6
#449730000000
1!
1%
1-
12
#449740000000
0!
0%
b111 *
0-
02
b111 6
#449750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#449760000000
0!
0%
b0 *
0-
02
b0 6
#449770000000
1!
1%
1-
12
#449780000000
0!
0%
b1 *
0-
02
b1 6
#449790000000
1!
1%
1-
12
#449800000000
0!
0%
b10 *
0-
02
b10 6
#449810000000
1!
1%
1-
12
#449820000000
0!
0%
b11 *
0-
02
b11 6
#449830000000
1!
1%
1-
12
15
#449840000000
0!
0%
b100 *
0-
02
b100 6
#449850000000
1!
1%
1-
12
#449860000000
0!
0%
b101 *
0-
02
b101 6
#449870000000
1!
1%
1-
12
#449880000000
0!
0%
b110 *
0-
02
b110 6
#449890000000
1!
1%
1-
12
#449900000000
0!
0%
b111 *
0-
02
b111 6
#449910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#449920000000
0!
0%
b0 *
0-
02
b0 6
#449930000000
1!
1%
1-
12
#449940000000
0!
0%
b1 *
0-
02
b1 6
#449950000000
1!
1%
1-
12
#449960000000
0!
0%
b10 *
0-
02
b10 6
#449970000000
1!
1%
1-
12
#449980000000
0!
0%
b11 *
0-
02
b11 6
#449990000000
1!
1%
1-
12
15
#450000000000
0!
0%
b100 *
0-
02
b100 6
#450010000000
1!
1%
1-
12
#450020000000
0!
0%
b101 *
0-
02
b101 6
#450030000000
1!
1%
1-
12
#450040000000
0!
0%
b110 *
0-
02
b110 6
#450050000000
1!
1%
1-
12
#450060000000
0!
0%
b111 *
0-
02
b111 6
#450070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#450080000000
0!
0%
b0 *
0-
02
b0 6
#450090000000
1!
1%
1-
12
#450100000000
0!
0%
b1 *
0-
02
b1 6
#450110000000
1!
1%
1-
12
#450120000000
0!
0%
b10 *
0-
02
b10 6
#450130000000
1!
1%
1-
12
#450140000000
0!
0%
b11 *
0-
02
b11 6
#450150000000
1!
1%
1-
12
15
#450160000000
0!
0%
b100 *
0-
02
b100 6
#450170000000
1!
1%
1-
12
#450180000000
0!
0%
b101 *
0-
02
b101 6
#450190000000
1!
1%
1-
12
#450200000000
0!
0%
b110 *
0-
02
b110 6
#450210000000
1!
1%
1-
12
#450220000000
0!
0%
b111 *
0-
02
b111 6
#450230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#450240000000
0!
0%
b0 *
0-
02
b0 6
#450250000000
1!
1%
1-
12
#450260000000
0!
0%
b1 *
0-
02
b1 6
#450270000000
1!
1%
1-
12
#450280000000
0!
0%
b10 *
0-
02
b10 6
#450290000000
1!
1%
1-
12
#450300000000
0!
0%
b11 *
0-
02
b11 6
#450310000000
1!
1%
1-
12
15
#450320000000
0!
0%
b100 *
0-
02
b100 6
#450330000000
1!
1%
1-
12
#450340000000
0!
0%
b101 *
0-
02
b101 6
#450350000000
1!
1%
1-
12
#450360000000
0!
0%
b110 *
0-
02
b110 6
#450370000000
1!
1%
1-
12
#450380000000
0!
0%
b111 *
0-
02
b111 6
#450390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#450400000000
0!
0%
b0 *
0-
02
b0 6
#450410000000
1!
1%
1-
12
#450420000000
0!
0%
b1 *
0-
02
b1 6
#450430000000
1!
1%
1-
12
#450440000000
0!
0%
b10 *
0-
02
b10 6
#450450000000
1!
1%
1-
12
#450460000000
0!
0%
b11 *
0-
02
b11 6
#450470000000
1!
1%
1-
12
15
#450480000000
0!
0%
b100 *
0-
02
b100 6
#450490000000
1!
1%
1-
12
#450500000000
0!
0%
b101 *
0-
02
b101 6
#450510000000
1!
1%
1-
12
#450520000000
0!
0%
b110 *
0-
02
b110 6
#450530000000
1!
1%
1-
12
#450540000000
0!
0%
b111 *
0-
02
b111 6
#450550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#450560000000
0!
0%
b0 *
0-
02
b0 6
#450570000000
1!
1%
1-
12
#450580000000
0!
0%
b1 *
0-
02
b1 6
#450590000000
1!
1%
1-
12
#450600000000
0!
0%
b10 *
0-
02
b10 6
#450610000000
1!
1%
1-
12
#450620000000
0!
0%
b11 *
0-
02
b11 6
#450630000000
1!
1%
1-
12
15
#450640000000
0!
0%
b100 *
0-
02
b100 6
#450650000000
1!
1%
1-
12
#450660000000
0!
0%
b101 *
0-
02
b101 6
#450670000000
1!
1%
1-
12
#450680000000
0!
0%
b110 *
0-
02
b110 6
#450690000000
1!
1%
1-
12
#450700000000
0!
0%
b111 *
0-
02
b111 6
#450710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#450720000000
0!
0%
b0 *
0-
02
b0 6
#450730000000
1!
1%
1-
12
#450740000000
0!
0%
b1 *
0-
02
b1 6
#450750000000
1!
1%
1-
12
#450760000000
0!
0%
b10 *
0-
02
b10 6
#450770000000
1!
1%
1-
12
#450780000000
0!
0%
b11 *
0-
02
b11 6
#450790000000
1!
1%
1-
12
15
#450800000000
0!
0%
b100 *
0-
02
b100 6
#450810000000
1!
1%
1-
12
#450820000000
0!
0%
b101 *
0-
02
b101 6
#450830000000
1!
1%
1-
12
#450840000000
0!
0%
b110 *
0-
02
b110 6
#450850000000
1!
1%
1-
12
#450860000000
0!
0%
b111 *
0-
02
b111 6
#450870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#450880000000
0!
0%
b0 *
0-
02
b0 6
#450890000000
1!
1%
1-
12
#450900000000
0!
0%
b1 *
0-
02
b1 6
#450910000000
1!
1%
1-
12
#450920000000
0!
0%
b10 *
0-
02
b10 6
#450930000000
1!
1%
1-
12
#450940000000
0!
0%
b11 *
0-
02
b11 6
#450950000000
1!
1%
1-
12
15
#450960000000
0!
0%
b100 *
0-
02
b100 6
#450970000000
1!
1%
1-
12
#450980000000
0!
0%
b101 *
0-
02
b101 6
#450990000000
1!
1%
1-
12
#451000000000
0!
0%
b110 *
0-
02
b110 6
#451010000000
1!
1%
1-
12
#451020000000
0!
0%
b111 *
0-
02
b111 6
#451030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#451040000000
0!
0%
b0 *
0-
02
b0 6
#451050000000
1!
1%
1-
12
#451060000000
0!
0%
b1 *
0-
02
b1 6
#451070000000
1!
1%
1-
12
#451080000000
0!
0%
b10 *
0-
02
b10 6
#451090000000
1!
1%
1-
12
#451100000000
0!
0%
b11 *
0-
02
b11 6
#451110000000
1!
1%
1-
12
15
#451120000000
0!
0%
b100 *
0-
02
b100 6
#451130000000
1!
1%
1-
12
#451140000000
0!
0%
b101 *
0-
02
b101 6
#451150000000
1!
1%
1-
12
#451160000000
0!
0%
b110 *
0-
02
b110 6
#451170000000
1!
1%
1-
12
#451180000000
0!
0%
b111 *
0-
02
b111 6
#451190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#451200000000
0!
0%
b0 *
0-
02
b0 6
#451210000000
1!
1%
1-
12
#451220000000
0!
0%
b1 *
0-
02
b1 6
#451230000000
1!
1%
1-
12
#451240000000
0!
0%
b10 *
0-
02
b10 6
#451250000000
1!
1%
1-
12
#451260000000
0!
0%
b11 *
0-
02
b11 6
#451270000000
1!
1%
1-
12
15
#451280000000
0!
0%
b100 *
0-
02
b100 6
#451290000000
1!
1%
1-
12
#451300000000
0!
0%
b101 *
0-
02
b101 6
#451310000000
1!
1%
1-
12
#451320000000
0!
0%
b110 *
0-
02
b110 6
#451330000000
1!
1%
1-
12
#451340000000
0!
0%
b111 *
0-
02
b111 6
#451350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#451360000000
0!
0%
b0 *
0-
02
b0 6
#451370000000
1!
1%
1-
12
#451380000000
0!
0%
b1 *
0-
02
b1 6
#451390000000
1!
1%
1-
12
#451400000000
0!
0%
b10 *
0-
02
b10 6
#451410000000
1!
1%
1-
12
#451420000000
0!
0%
b11 *
0-
02
b11 6
#451430000000
1!
1%
1-
12
15
#451440000000
0!
0%
b100 *
0-
02
b100 6
#451450000000
1!
1%
1-
12
#451460000000
0!
0%
b101 *
0-
02
b101 6
#451470000000
1!
1%
1-
12
#451480000000
0!
0%
b110 *
0-
02
b110 6
#451490000000
1!
1%
1-
12
#451500000000
0!
0%
b111 *
0-
02
b111 6
#451510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#451520000000
0!
0%
b0 *
0-
02
b0 6
#451530000000
1!
1%
1-
12
#451540000000
0!
0%
b1 *
0-
02
b1 6
#451550000000
1!
1%
1-
12
#451560000000
0!
0%
b10 *
0-
02
b10 6
#451570000000
1!
1%
1-
12
#451580000000
0!
0%
b11 *
0-
02
b11 6
#451590000000
1!
1%
1-
12
15
#451600000000
0!
0%
b100 *
0-
02
b100 6
#451610000000
1!
1%
1-
12
#451620000000
0!
0%
b101 *
0-
02
b101 6
#451630000000
1!
1%
1-
12
#451640000000
0!
0%
b110 *
0-
02
b110 6
#451650000000
1!
1%
1-
12
#451660000000
0!
0%
b111 *
0-
02
b111 6
#451670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#451680000000
0!
0%
b0 *
0-
02
b0 6
#451690000000
1!
1%
1-
12
#451700000000
0!
0%
b1 *
0-
02
b1 6
#451710000000
1!
1%
1-
12
#451720000000
0!
0%
b10 *
0-
02
b10 6
#451730000000
1!
1%
1-
12
#451740000000
0!
0%
b11 *
0-
02
b11 6
#451750000000
1!
1%
1-
12
15
#451760000000
0!
0%
b100 *
0-
02
b100 6
#451770000000
1!
1%
1-
12
#451780000000
0!
0%
b101 *
0-
02
b101 6
#451790000000
1!
1%
1-
12
#451800000000
0!
0%
b110 *
0-
02
b110 6
#451810000000
1!
1%
1-
12
#451820000000
0!
0%
b111 *
0-
02
b111 6
#451830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#451840000000
0!
0%
b0 *
0-
02
b0 6
#451850000000
1!
1%
1-
12
#451860000000
0!
0%
b1 *
0-
02
b1 6
#451870000000
1!
1%
1-
12
#451880000000
0!
0%
b10 *
0-
02
b10 6
#451890000000
1!
1%
1-
12
#451900000000
0!
0%
b11 *
0-
02
b11 6
#451910000000
1!
1%
1-
12
15
#451920000000
0!
0%
b100 *
0-
02
b100 6
#451930000000
1!
1%
1-
12
#451940000000
0!
0%
b101 *
0-
02
b101 6
#451950000000
1!
1%
1-
12
#451960000000
0!
0%
b110 *
0-
02
b110 6
#451970000000
1!
1%
1-
12
#451980000000
0!
0%
b111 *
0-
02
b111 6
#451990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#452000000000
0!
0%
b0 *
0-
02
b0 6
#452010000000
1!
1%
1-
12
#452020000000
0!
0%
b1 *
0-
02
b1 6
#452030000000
1!
1%
1-
12
#452040000000
0!
0%
b10 *
0-
02
b10 6
#452050000000
1!
1%
1-
12
#452060000000
0!
0%
b11 *
0-
02
b11 6
#452070000000
1!
1%
1-
12
15
#452080000000
0!
0%
b100 *
0-
02
b100 6
#452090000000
1!
1%
1-
12
#452100000000
0!
0%
b101 *
0-
02
b101 6
#452110000000
1!
1%
1-
12
#452120000000
0!
0%
b110 *
0-
02
b110 6
#452130000000
1!
1%
1-
12
#452140000000
0!
0%
b111 *
0-
02
b111 6
#452150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#452160000000
0!
0%
b0 *
0-
02
b0 6
#452170000000
1!
1%
1-
12
#452180000000
0!
0%
b1 *
0-
02
b1 6
#452190000000
1!
1%
1-
12
#452200000000
0!
0%
b10 *
0-
02
b10 6
#452210000000
1!
1%
1-
12
#452220000000
0!
0%
b11 *
0-
02
b11 6
#452230000000
1!
1%
1-
12
15
#452240000000
0!
0%
b100 *
0-
02
b100 6
#452250000000
1!
1%
1-
12
#452260000000
0!
0%
b101 *
0-
02
b101 6
#452270000000
1!
1%
1-
12
#452280000000
0!
0%
b110 *
0-
02
b110 6
#452290000000
1!
1%
1-
12
#452300000000
0!
0%
b111 *
0-
02
b111 6
#452310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#452320000000
0!
0%
b0 *
0-
02
b0 6
#452330000000
1!
1%
1-
12
#452340000000
0!
0%
b1 *
0-
02
b1 6
#452350000000
1!
1%
1-
12
#452360000000
0!
0%
b10 *
0-
02
b10 6
#452370000000
1!
1%
1-
12
#452380000000
0!
0%
b11 *
0-
02
b11 6
#452390000000
1!
1%
1-
12
15
#452400000000
0!
0%
b100 *
0-
02
b100 6
#452410000000
1!
1%
1-
12
#452420000000
0!
0%
b101 *
0-
02
b101 6
#452430000000
1!
1%
1-
12
#452440000000
0!
0%
b110 *
0-
02
b110 6
#452450000000
1!
1%
1-
12
#452460000000
0!
0%
b111 *
0-
02
b111 6
#452470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#452480000000
0!
0%
b0 *
0-
02
b0 6
#452490000000
1!
1%
1-
12
#452500000000
0!
0%
b1 *
0-
02
b1 6
#452510000000
1!
1%
1-
12
#452520000000
0!
0%
b10 *
0-
02
b10 6
#452530000000
1!
1%
1-
12
#452540000000
0!
0%
b11 *
0-
02
b11 6
#452550000000
1!
1%
1-
12
15
#452560000000
0!
0%
b100 *
0-
02
b100 6
#452570000000
1!
1%
1-
12
#452580000000
0!
0%
b101 *
0-
02
b101 6
#452590000000
1!
1%
1-
12
#452600000000
0!
0%
b110 *
0-
02
b110 6
#452610000000
1!
1%
1-
12
#452620000000
0!
0%
b111 *
0-
02
b111 6
#452630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#452640000000
0!
0%
b0 *
0-
02
b0 6
#452650000000
1!
1%
1-
12
#452660000000
0!
0%
b1 *
0-
02
b1 6
#452670000000
1!
1%
1-
12
#452680000000
0!
0%
b10 *
0-
02
b10 6
#452690000000
1!
1%
1-
12
#452700000000
0!
0%
b11 *
0-
02
b11 6
#452710000000
1!
1%
1-
12
15
#452720000000
0!
0%
b100 *
0-
02
b100 6
#452730000000
1!
1%
1-
12
#452740000000
0!
0%
b101 *
0-
02
b101 6
#452750000000
1!
1%
1-
12
#452760000000
0!
0%
b110 *
0-
02
b110 6
#452770000000
1!
1%
1-
12
#452780000000
0!
0%
b111 *
0-
02
b111 6
#452790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#452800000000
0!
0%
b0 *
0-
02
b0 6
#452810000000
1!
1%
1-
12
#452820000000
0!
0%
b1 *
0-
02
b1 6
#452830000000
1!
1%
1-
12
#452840000000
0!
0%
b10 *
0-
02
b10 6
#452850000000
1!
1%
1-
12
#452860000000
0!
0%
b11 *
0-
02
b11 6
#452870000000
1!
1%
1-
12
15
#452880000000
0!
0%
b100 *
0-
02
b100 6
#452890000000
1!
1%
1-
12
#452900000000
0!
0%
b101 *
0-
02
b101 6
#452910000000
1!
1%
1-
12
#452920000000
0!
0%
b110 *
0-
02
b110 6
#452930000000
1!
1%
1-
12
#452940000000
0!
0%
b111 *
0-
02
b111 6
#452950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#452960000000
0!
0%
b0 *
0-
02
b0 6
#452970000000
1!
1%
1-
12
#452980000000
0!
0%
b1 *
0-
02
b1 6
#452990000000
1!
1%
1-
12
#453000000000
0!
0%
b10 *
0-
02
b10 6
#453010000000
1!
1%
1-
12
#453020000000
0!
0%
b11 *
0-
02
b11 6
#453030000000
1!
1%
1-
12
15
#453040000000
0!
0%
b100 *
0-
02
b100 6
#453050000000
1!
1%
1-
12
#453060000000
0!
0%
b101 *
0-
02
b101 6
#453070000000
1!
1%
1-
12
#453080000000
0!
0%
b110 *
0-
02
b110 6
#453090000000
1!
1%
1-
12
#453100000000
0!
0%
b111 *
0-
02
b111 6
#453110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#453120000000
0!
0%
b0 *
0-
02
b0 6
#453130000000
1!
1%
1-
12
#453140000000
0!
0%
b1 *
0-
02
b1 6
#453150000000
1!
1%
1-
12
#453160000000
0!
0%
b10 *
0-
02
b10 6
#453170000000
1!
1%
1-
12
#453180000000
0!
0%
b11 *
0-
02
b11 6
#453190000000
1!
1%
1-
12
15
#453200000000
0!
0%
b100 *
0-
02
b100 6
#453210000000
1!
1%
1-
12
#453220000000
0!
0%
b101 *
0-
02
b101 6
#453230000000
1!
1%
1-
12
#453240000000
0!
0%
b110 *
0-
02
b110 6
#453250000000
1!
1%
1-
12
#453260000000
0!
0%
b111 *
0-
02
b111 6
#453270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#453280000000
0!
0%
b0 *
0-
02
b0 6
#453290000000
1!
1%
1-
12
#453300000000
0!
0%
b1 *
0-
02
b1 6
#453310000000
1!
1%
1-
12
#453320000000
0!
0%
b10 *
0-
02
b10 6
#453330000000
1!
1%
1-
12
#453340000000
0!
0%
b11 *
0-
02
b11 6
#453350000000
1!
1%
1-
12
15
#453360000000
0!
0%
b100 *
0-
02
b100 6
#453370000000
1!
1%
1-
12
#453380000000
0!
0%
b101 *
0-
02
b101 6
#453390000000
1!
1%
1-
12
#453400000000
0!
0%
b110 *
0-
02
b110 6
#453410000000
1!
1%
1-
12
#453420000000
0!
0%
b111 *
0-
02
b111 6
#453430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#453440000000
0!
0%
b0 *
0-
02
b0 6
#453450000000
1!
1%
1-
12
#453460000000
0!
0%
b1 *
0-
02
b1 6
#453470000000
1!
1%
1-
12
#453480000000
0!
0%
b10 *
0-
02
b10 6
#453490000000
1!
1%
1-
12
#453500000000
0!
0%
b11 *
0-
02
b11 6
#453510000000
1!
1%
1-
12
15
#453520000000
0!
0%
b100 *
0-
02
b100 6
#453530000000
1!
1%
1-
12
#453540000000
0!
0%
b101 *
0-
02
b101 6
#453550000000
1!
1%
1-
12
#453560000000
0!
0%
b110 *
0-
02
b110 6
#453570000000
1!
1%
1-
12
#453580000000
0!
0%
b111 *
0-
02
b111 6
#453590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#453600000000
0!
0%
b0 *
0-
02
b0 6
#453610000000
1!
1%
1-
12
#453620000000
0!
0%
b1 *
0-
02
b1 6
#453630000000
1!
1%
1-
12
#453640000000
0!
0%
b10 *
0-
02
b10 6
#453650000000
1!
1%
1-
12
#453660000000
0!
0%
b11 *
0-
02
b11 6
#453670000000
1!
1%
1-
12
15
#453680000000
0!
0%
b100 *
0-
02
b100 6
#453690000000
1!
1%
1-
12
#453700000000
0!
0%
b101 *
0-
02
b101 6
#453710000000
1!
1%
1-
12
#453720000000
0!
0%
b110 *
0-
02
b110 6
#453730000000
1!
1%
1-
12
#453740000000
0!
0%
b111 *
0-
02
b111 6
#453750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#453760000000
0!
0%
b0 *
0-
02
b0 6
#453770000000
1!
1%
1-
12
#453780000000
0!
0%
b1 *
0-
02
b1 6
#453790000000
1!
1%
1-
12
#453800000000
0!
0%
b10 *
0-
02
b10 6
#453810000000
1!
1%
1-
12
#453820000000
0!
0%
b11 *
0-
02
b11 6
#453830000000
1!
1%
1-
12
15
#453840000000
0!
0%
b100 *
0-
02
b100 6
#453850000000
1!
1%
1-
12
#453860000000
0!
0%
b101 *
0-
02
b101 6
#453870000000
1!
1%
1-
12
#453880000000
0!
0%
b110 *
0-
02
b110 6
#453890000000
1!
1%
1-
12
#453900000000
0!
0%
b111 *
0-
02
b111 6
#453910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#453920000000
0!
0%
b0 *
0-
02
b0 6
#453930000000
1!
1%
1-
12
#453940000000
0!
0%
b1 *
0-
02
b1 6
#453950000000
1!
1%
1-
12
#453960000000
0!
0%
b10 *
0-
02
b10 6
#453970000000
1!
1%
1-
12
#453980000000
0!
0%
b11 *
0-
02
b11 6
#453990000000
1!
1%
1-
12
15
#454000000000
0!
0%
b100 *
0-
02
b100 6
#454010000000
1!
1%
1-
12
#454020000000
0!
0%
b101 *
0-
02
b101 6
#454030000000
1!
1%
1-
12
#454040000000
0!
0%
b110 *
0-
02
b110 6
#454050000000
1!
1%
1-
12
#454060000000
0!
0%
b111 *
0-
02
b111 6
#454070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#454080000000
0!
0%
b0 *
0-
02
b0 6
#454090000000
1!
1%
1-
12
#454100000000
0!
0%
b1 *
0-
02
b1 6
#454110000000
1!
1%
1-
12
#454120000000
0!
0%
b10 *
0-
02
b10 6
#454130000000
1!
1%
1-
12
#454140000000
0!
0%
b11 *
0-
02
b11 6
#454150000000
1!
1%
1-
12
15
#454160000000
0!
0%
b100 *
0-
02
b100 6
#454170000000
1!
1%
1-
12
#454180000000
0!
0%
b101 *
0-
02
b101 6
#454190000000
1!
1%
1-
12
#454200000000
0!
0%
b110 *
0-
02
b110 6
#454210000000
1!
1%
1-
12
#454220000000
0!
0%
b111 *
0-
02
b111 6
#454230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#454240000000
0!
0%
b0 *
0-
02
b0 6
#454250000000
1!
1%
1-
12
#454260000000
0!
0%
b1 *
0-
02
b1 6
#454270000000
1!
1%
1-
12
#454280000000
0!
0%
b10 *
0-
02
b10 6
#454290000000
1!
1%
1-
12
#454300000000
0!
0%
b11 *
0-
02
b11 6
#454310000000
1!
1%
1-
12
15
#454320000000
0!
0%
b100 *
0-
02
b100 6
#454330000000
1!
1%
1-
12
#454340000000
0!
0%
b101 *
0-
02
b101 6
#454350000000
1!
1%
1-
12
#454360000000
0!
0%
b110 *
0-
02
b110 6
#454370000000
1!
1%
1-
12
#454380000000
0!
0%
b111 *
0-
02
b111 6
#454390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#454400000000
0!
0%
b0 *
0-
02
b0 6
#454410000000
1!
1%
1-
12
#454420000000
0!
0%
b1 *
0-
02
b1 6
#454430000000
1!
1%
1-
12
#454440000000
0!
0%
b10 *
0-
02
b10 6
#454450000000
1!
1%
1-
12
#454460000000
0!
0%
b11 *
0-
02
b11 6
#454470000000
1!
1%
1-
12
15
#454480000000
0!
0%
b100 *
0-
02
b100 6
#454490000000
1!
1%
1-
12
#454500000000
0!
0%
b101 *
0-
02
b101 6
#454510000000
1!
1%
1-
12
#454520000000
0!
0%
b110 *
0-
02
b110 6
#454530000000
1!
1%
1-
12
#454540000000
0!
0%
b111 *
0-
02
b111 6
#454550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#454560000000
0!
0%
b0 *
0-
02
b0 6
#454570000000
1!
1%
1-
12
#454580000000
0!
0%
b1 *
0-
02
b1 6
#454590000000
1!
1%
1-
12
#454600000000
0!
0%
b10 *
0-
02
b10 6
#454610000000
1!
1%
1-
12
#454620000000
0!
0%
b11 *
0-
02
b11 6
#454630000000
1!
1%
1-
12
15
#454640000000
0!
0%
b100 *
0-
02
b100 6
#454650000000
1!
1%
1-
12
#454660000000
0!
0%
b101 *
0-
02
b101 6
#454670000000
1!
1%
1-
12
#454680000000
0!
0%
b110 *
0-
02
b110 6
#454690000000
1!
1%
1-
12
#454700000000
0!
0%
b111 *
0-
02
b111 6
#454710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#454720000000
0!
0%
b0 *
0-
02
b0 6
#454730000000
1!
1%
1-
12
#454740000000
0!
0%
b1 *
0-
02
b1 6
#454750000000
1!
1%
1-
12
#454760000000
0!
0%
b10 *
0-
02
b10 6
#454770000000
1!
1%
1-
12
#454780000000
0!
0%
b11 *
0-
02
b11 6
#454790000000
1!
1%
1-
12
15
#454800000000
0!
0%
b100 *
0-
02
b100 6
#454810000000
1!
1%
1-
12
#454820000000
0!
0%
b101 *
0-
02
b101 6
#454830000000
1!
1%
1-
12
#454840000000
0!
0%
b110 *
0-
02
b110 6
#454850000000
1!
1%
1-
12
#454860000000
0!
0%
b111 *
0-
02
b111 6
#454870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#454880000000
0!
0%
b0 *
0-
02
b0 6
#454890000000
1!
1%
1-
12
#454900000000
0!
0%
b1 *
0-
02
b1 6
#454910000000
1!
1%
1-
12
#454920000000
0!
0%
b10 *
0-
02
b10 6
#454930000000
1!
1%
1-
12
#454940000000
0!
0%
b11 *
0-
02
b11 6
#454950000000
1!
1%
1-
12
15
#454960000000
0!
0%
b100 *
0-
02
b100 6
#454970000000
1!
1%
1-
12
#454980000000
0!
0%
b101 *
0-
02
b101 6
#454990000000
1!
1%
1-
12
#455000000000
0!
0%
b110 *
0-
02
b110 6
#455010000000
1!
1%
1-
12
#455020000000
0!
0%
b111 *
0-
02
b111 6
#455030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#455040000000
0!
0%
b0 *
0-
02
b0 6
#455050000000
1!
1%
1-
12
#455060000000
0!
0%
b1 *
0-
02
b1 6
#455070000000
1!
1%
1-
12
#455080000000
0!
0%
b10 *
0-
02
b10 6
#455090000000
1!
1%
1-
12
#455100000000
0!
0%
b11 *
0-
02
b11 6
#455110000000
1!
1%
1-
12
15
#455120000000
0!
0%
b100 *
0-
02
b100 6
#455130000000
1!
1%
1-
12
#455140000000
0!
0%
b101 *
0-
02
b101 6
#455150000000
1!
1%
1-
12
#455160000000
0!
0%
b110 *
0-
02
b110 6
#455170000000
1!
1%
1-
12
#455180000000
0!
0%
b111 *
0-
02
b111 6
#455190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#455200000000
0!
0%
b0 *
0-
02
b0 6
#455210000000
1!
1%
1-
12
#455220000000
0!
0%
b1 *
0-
02
b1 6
#455230000000
1!
1%
1-
12
#455240000000
0!
0%
b10 *
0-
02
b10 6
#455250000000
1!
1%
1-
12
#455260000000
0!
0%
b11 *
0-
02
b11 6
#455270000000
1!
1%
1-
12
15
#455280000000
0!
0%
b100 *
0-
02
b100 6
#455290000000
1!
1%
1-
12
#455300000000
0!
0%
b101 *
0-
02
b101 6
#455310000000
1!
1%
1-
12
#455320000000
0!
0%
b110 *
0-
02
b110 6
#455330000000
1!
1%
1-
12
#455340000000
0!
0%
b111 *
0-
02
b111 6
#455350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#455360000000
0!
0%
b0 *
0-
02
b0 6
#455370000000
1!
1%
1-
12
#455380000000
0!
0%
b1 *
0-
02
b1 6
#455390000000
1!
1%
1-
12
#455400000000
0!
0%
b10 *
0-
02
b10 6
#455410000000
1!
1%
1-
12
#455420000000
0!
0%
b11 *
0-
02
b11 6
#455430000000
1!
1%
1-
12
15
#455440000000
0!
0%
b100 *
0-
02
b100 6
#455450000000
1!
1%
1-
12
#455460000000
0!
0%
b101 *
0-
02
b101 6
#455470000000
1!
1%
1-
12
#455480000000
0!
0%
b110 *
0-
02
b110 6
#455490000000
1!
1%
1-
12
#455500000000
0!
0%
b111 *
0-
02
b111 6
#455510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#455520000000
0!
0%
b0 *
0-
02
b0 6
#455530000000
1!
1%
1-
12
#455540000000
0!
0%
b1 *
0-
02
b1 6
#455550000000
1!
1%
1-
12
#455560000000
0!
0%
b10 *
0-
02
b10 6
#455570000000
1!
1%
1-
12
#455580000000
0!
0%
b11 *
0-
02
b11 6
#455590000000
1!
1%
1-
12
15
#455600000000
0!
0%
b100 *
0-
02
b100 6
#455610000000
1!
1%
1-
12
#455620000000
0!
0%
b101 *
0-
02
b101 6
#455630000000
1!
1%
1-
12
#455640000000
0!
0%
b110 *
0-
02
b110 6
#455650000000
1!
1%
1-
12
#455660000000
0!
0%
b111 *
0-
02
b111 6
#455670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#455680000000
0!
0%
b0 *
0-
02
b0 6
#455690000000
1!
1%
1-
12
#455700000000
0!
0%
b1 *
0-
02
b1 6
#455710000000
1!
1%
1-
12
#455720000000
0!
0%
b10 *
0-
02
b10 6
#455730000000
1!
1%
1-
12
#455740000000
0!
0%
b11 *
0-
02
b11 6
#455750000000
1!
1%
1-
12
15
#455760000000
0!
0%
b100 *
0-
02
b100 6
#455770000000
1!
1%
1-
12
#455780000000
0!
0%
b101 *
0-
02
b101 6
#455790000000
1!
1%
1-
12
#455800000000
0!
0%
b110 *
0-
02
b110 6
#455810000000
1!
1%
1-
12
#455820000000
0!
0%
b111 *
0-
02
b111 6
#455830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#455840000000
0!
0%
b0 *
0-
02
b0 6
#455850000000
1!
1%
1-
12
#455860000000
0!
0%
b1 *
0-
02
b1 6
#455870000000
1!
1%
1-
12
#455880000000
0!
0%
b10 *
0-
02
b10 6
#455890000000
1!
1%
1-
12
#455900000000
0!
0%
b11 *
0-
02
b11 6
#455910000000
1!
1%
1-
12
15
#455920000000
0!
0%
b100 *
0-
02
b100 6
#455930000000
1!
1%
1-
12
#455940000000
0!
0%
b101 *
0-
02
b101 6
#455950000000
1!
1%
1-
12
#455960000000
0!
0%
b110 *
0-
02
b110 6
#455970000000
1!
1%
1-
12
#455980000000
0!
0%
b111 *
0-
02
b111 6
#455990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#456000000000
0!
0%
b0 *
0-
02
b0 6
#456010000000
1!
1%
1-
12
#456020000000
0!
0%
b1 *
0-
02
b1 6
#456030000000
1!
1%
1-
12
#456040000000
0!
0%
b10 *
0-
02
b10 6
#456050000000
1!
1%
1-
12
#456060000000
0!
0%
b11 *
0-
02
b11 6
#456070000000
1!
1%
1-
12
15
#456080000000
0!
0%
b100 *
0-
02
b100 6
#456090000000
1!
1%
1-
12
#456100000000
0!
0%
b101 *
0-
02
b101 6
#456110000000
1!
1%
1-
12
#456120000000
0!
0%
b110 *
0-
02
b110 6
#456130000000
1!
1%
1-
12
#456140000000
0!
0%
b111 *
0-
02
b111 6
#456150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#456160000000
0!
0%
b0 *
0-
02
b0 6
#456170000000
1!
1%
1-
12
#456180000000
0!
0%
b1 *
0-
02
b1 6
#456190000000
1!
1%
1-
12
#456200000000
0!
0%
b10 *
0-
02
b10 6
#456210000000
1!
1%
1-
12
#456220000000
0!
0%
b11 *
0-
02
b11 6
#456230000000
1!
1%
1-
12
15
#456240000000
0!
0%
b100 *
0-
02
b100 6
#456250000000
1!
1%
1-
12
#456260000000
0!
0%
b101 *
0-
02
b101 6
#456270000000
1!
1%
1-
12
#456280000000
0!
0%
b110 *
0-
02
b110 6
#456290000000
1!
1%
1-
12
#456300000000
0!
0%
b111 *
0-
02
b111 6
#456310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#456320000000
0!
0%
b0 *
0-
02
b0 6
#456330000000
1!
1%
1-
12
#456340000000
0!
0%
b1 *
0-
02
b1 6
#456350000000
1!
1%
1-
12
#456360000000
0!
0%
b10 *
0-
02
b10 6
#456370000000
1!
1%
1-
12
#456380000000
0!
0%
b11 *
0-
02
b11 6
#456390000000
1!
1%
1-
12
15
#456400000000
0!
0%
b100 *
0-
02
b100 6
#456410000000
1!
1%
1-
12
#456420000000
0!
0%
b101 *
0-
02
b101 6
#456430000000
1!
1%
1-
12
#456440000000
0!
0%
b110 *
0-
02
b110 6
#456450000000
1!
1%
1-
12
#456460000000
0!
0%
b111 *
0-
02
b111 6
#456470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#456480000000
0!
0%
b0 *
0-
02
b0 6
#456490000000
1!
1%
1-
12
#456500000000
0!
0%
b1 *
0-
02
b1 6
#456510000000
1!
1%
1-
12
#456520000000
0!
0%
b10 *
0-
02
b10 6
#456530000000
1!
1%
1-
12
#456540000000
0!
0%
b11 *
0-
02
b11 6
#456550000000
1!
1%
1-
12
15
#456560000000
0!
0%
b100 *
0-
02
b100 6
#456570000000
1!
1%
1-
12
#456580000000
0!
0%
b101 *
0-
02
b101 6
#456590000000
1!
1%
1-
12
#456600000000
0!
0%
b110 *
0-
02
b110 6
#456610000000
1!
1%
1-
12
#456620000000
0!
0%
b111 *
0-
02
b111 6
#456630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#456640000000
0!
0%
b0 *
0-
02
b0 6
#456650000000
1!
1%
1-
12
#456660000000
0!
0%
b1 *
0-
02
b1 6
#456670000000
1!
1%
1-
12
#456680000000
0!
0%
b10 *
0-
02
b10 6
#456690000000
1!
1%
1-
12
#456700000000
0!
0%
b11 *
0-
02
b11 6
#456710000000
1!
1%
1-
12
15
#456720000000
0!
0%
b100 *
0-
02
b100 6
#456730000000
1!
1%
1-
12
#456740000000
0!
0%
b101 *
0-
02
b101 6
#456750000000
1!
1%
1-
12
#456760000000
0!
0%
b110 *
0-
02
b110 6
#456770000000
1!
1%
1-
12
#456780000000
0!
0%
b111 *
0-
02
b111 6
#456790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#456800000000
0!
0%
b0 *
0-
02
b0 6
#456810000000
1!
1%
1-
12
#456820000000
0!
0%
b1 *
0-
02
b1 6
#456830000000
1!
1%
1-
12
#456840000000
0!
0%
b10 *
0-
02
b10 6
#456850000000
1!
1%
1-
12
#456860000000
0!
0%
b11 *
0-
02
b11 6
#456870000000
1!
1%
1-
12
15
#456880000000
0!
0%
b100 *
0-
02
b100 6
#456890000000
1!
1%
1-
12
#456900000000
0!
0%
b101 *
0-
02
b101 6
#456910000000
1!
1%
1-
12
#456920000000
0!
0%
b110 *
0-
02
b110 6
#456930000000
1!
1%
1-
12
#456940000000
0!
0%
b111 *
0-
02
b111 6
#456950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#456960000000
0!
0%
b0 *
0-
02
b0 6
#456970000000
1!
1%
1-
12
#456980000000
0!
0%
b1 *
0-
02
b1 6
#456990000000
1!
1%
1-
12
#457000000000
0!
0%
b10 *
0-
02
b10 6
#457010000000
1!
1%
1-
12
#457020000000
0!
0%
b11 *
0-
02
b11 6
#457030000000
1!
1%
1-
12
15
#457040000000
0!
0%
b100 *
0-
02
b100 6
#457050000000
1!
1%
1-
12
#457060000000
0!
0%
b101 *
0-
02
b101 6
#457070000000
1!
1%
1-
12
#457080000000
0!
0%
b110 *
0-
02
b110 6
#457090000000
1!
1%
1-
12
#457100000000
0!
0%
b111 *
0-
02
b111 6
#457110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#457120000000
0!
0%
b0 *
0-
02
b0 6
#457130000000
1!
1%
1-
12
#457140000000
0!
0%
b1 *
0-
02
b1 6
#457150000000
1!
1%
1-
12
#457160000000
0!
0%
b10 *
0-
02
b10 6
#457170000000
1!
1%
1-
12
#457180000000
0!
0%
b11 *
0-
02
b11 6
#457190000000
1!
1%
1-
12
15
#457200000000
0!
0%
b100 *
0-
02
b100 6
#457210000000
1!
1%
1-
12
#457220000000
0!
0%
b101 *
0-
02
b101 6
#457230000000
1!
1%
1-
12
#457240000000
0!
0%
b110 *
0-
02
b110 6
#457250000000
1!
1%
1-
12
#457260000000
0!
0%
b111 *
0-
02
b111 6
#457270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#457280000000
0!
0%
b0 *
0-
02
b0 6
#457290000000
1!
1%
1-
12
#457300000000
0!
0%
b1 *
0-
02
b1 6
#457310000000
1!
1%
1-
12
#457320000000
0!
0%
b10 *
0-
02
b10 6
#457330000000
1!
1%
1-
12
#457340000000
0!
0%
b11 *
0-
02
b11 6
#457350000000
1!
1%
1-
12
15
#457360000000
0!
0%
b100 *
0-
02
b100 6
#457370000000
1!
1%
1-
12
#457380000000
0!
0%
b101 *
0-
02
b101 6
#457390000000
1!
1%
1-
12
#457400000000
0!
0%
b110 *
0-
02
b110 6
#457410000000
1!
1%
1-
12
#457420000000
0!
0%
b111 *
0-
02
b111 6
#457430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#457440000000
0!
0%
b0 *
0-
02
b0 6
#457450000000
1!
1%
1-
12
#457460000000
0!
0%
b1 *
0-
02
b1 6
#457470000000
1!
1%
1-
12
#457480000000
0!
0%
b10 *
0-
02
b10 6
#457490000000
1!
1%
1-
12
#457500000000
0!
0%
b11 *
0-
02
b11 6
#457510000000
1!
1%
1-
12
15
#457520000000
0!
0%
b100 *
0-
02
b100 6
#457530000000
1!
1%
1-
12
#457540000000
0!
0%
b101 *
0-
02
b101 6
#457550000000
1!
1%
1-
12
#457560000000
0!
0%
b110 *
0-
02
b110 6
#457570000000
1!
1%
1-
12
#457580000000
0!
0%
b111 *
0-
02
b111 6
#457590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#457600000000
0!
0%
b0 *
0-
02
b0 6
#457610000000
1!
1%
1-
12
#457620000000
0!
0%
b1 *
0-
02
b1 6
#457630000000
1!
1%
1-
12
#457640000000
0!
0%
b10 *
0-
02
b10 6
#457650000000
1!
1%
1-
12
#457660000000
0!
0%
b11 *
0-
02
b11 6
#457670000000
1!
1%
1-
12
15
#457680000000
0!
0%
b100 *
0-
02
b100 6
#457690000000
1!
1%
1-
12
#457700000000
0!
0%
b101 *
0-
02
b101 6
#457710000000
1!
1%
1-
12
#457720000000
0!
0%
b110 *
0-
02
b110 6
#457730000000
1!
1%
1-
12
#457740000000
0!
0%
b111 *
0-
02
b111 6
#457750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#457760000000
0!
0%
b0 *
0-
02
b0 6
#457770000000
1!
1%
1-
12
#457780000000
0!
0%
b1 *
0-
02
b1 6
#457790000000
1!
1%
1-
12
#457800000000
0!
0%
b10 *
0-
02
b10 6
#457810000000
1!
1%
1-
12
#457820000000
0!
0%
b11 *
0-
02
b11 6
#457830000000
1!
1%
1-
12
15
#457840000000
0!
0%
b100 *
0-
02
b100 6
#457850000000
1!
1%
1-
12
#457860000000
0!
0%
b101 *
0-
02
b101 6
#457870000000
1!
1%
1-
12
#457880000000
0!
0%
b110 *
0-
02
b110 6
#457890000000
1!
1%
1-
12
#457900000000
0!
0%
b111 *
0-
02
b111 6
#457910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#457920000000
0!
0%
b0 *
0-
02
b0 6
#457930000000
1!
1%
1-
12
#457940000000
0!
0%
b1 *
0-
02
b1 6
#457950000000
1!
1%
1-
12
#457960000000
0!
0%
b10 *
0-
02
b10 6
#457970000000
1!
1%
1-
12
#457980000000
0!
0%
b11 *
0-
02
b11 6
#457990000000
1!
1%
1-
12
15
#458000000000
0!
0%
b100 *
0-
02
b100 6
#458010000000
1!
1%
1-
12
#458020000000
0!
0%
b101 *
0-
02
b101 6
#458030000000
1!
1%
1-
12
#458040000000
0!
0%
b110 *
0-
02
b110 6
#458050000000
1!
1%
1-
12
#458060000000
0!
0%
b111 *
0-
02
b111 6
#458070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#458080000000
0!
0%
b0 *
0-
02
b0 6
#458090000000
1!
1%
1-
12
#458100000000
0!
0%
b1 *
0-
02
b1 6
#458110000000
1!
1%
1-
12
#458120000000
0!
0%
b10 *
0-
02
b10 6
#458130000000
1!
1%
1-
12
#458140000000
0!
0%
b11 *
0-
02
b11 6
#458150000000
1!
1%
1-
12
15
#458160000000
0!
0%
b100 *
0-
02
b100 6
#458170000000
1!
1%
1-
12
#458180000000
0!
0%
b101 *
0-
02
b101 6
#458190000000
1!
1%
1-
12
#458200000000
0!
0%
b110 *
0-
02
b110 6
#458210000000
1!
1%
1-
12
#458220000000
0!
0%
b111 *
0-
02
b111 6
#458230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#458240000000
0!
0%
b0 *
0-
02
b0 6
#458250000000
1!
1%
1-
12
#458260000000
0!
0%
b1 *
0-
02
b1 6
#458270000000
1!
1%
1-
12
#458280000000
0!
0%
b10 *
0-
02
b10 6
#458290000000
1!
1%
1-
12
#458300000000
0!
0%
b11 *
0-
02
b11 6
#458310000000
1!
1%
1-
12
15
#458320000000
0!
0%
b100 *
0-
02
b100 6
#458330000000
1!
1%
1-
12
#458340000000
0!
0%
b101 *
0-
02
b101 6
#458350000000
1!
1%
1-
12
#458360000000
0!
0%
b110 *
0-
02
b110 6
#458370000000
1!
1%
1-
12
#458380000000
0!
0%
b111 *
0-
02
b111 6
#458390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#458400000000
0!
0%
b0 *
0-
02
b0 6
#458410000000
1!
1%
1-
12
#458420000000
0!
0%
b1 *
0-
02
b1 6
#458430000000
1!
1%
1-
12
#458440000000
0!
0%
b10 *
0-
02
b10 6
#458450000000
1!
1%
1-
12
#458460000000
0!
0%
b11 *
0-
02
b11 6
#458470000000
1!
1%
1-
12
15
#458480000000
0!
0%
b100 *
0-
02
b100 6
#458490000000
1!
1%
1-
12
#458500000000
0!
0%
b101 *
0-
02
b101 6
#458510000000
1!
1%
1-
12
#458520000000
0!
0%
b110 *
0-
02
b110 6
#458530000000
1!
1%
1-
12
#458540000000
0!
0%
b111 *
0-
02
b111 6
#458550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#458560000000
0!
0%
b0 *
0-
02
b0 6
#458570000000
1!
1%
1-
12
#458580000000
0!
0%
b1 *
0-
02
b1 6
#458590000000
1!
1%
1-
12
#458600000000
0!
0%
b10 *
0-
02
b10 6
#458610000000
1!
1%
1-
12
#458620000000
0!
0%
b11 *
0-
02
b11 6
#458630000000
1!
1%
1-
12
15
#458640000000
0!
0%
b100 *
0-
02
b100 6
#458650000000
1!
1%
1-
12
#458660000000
0!
0%
b101 *
0-
02
b101 6
#458670000000
1!
1%
1-
12
#458680000000
0!
0%
b110 *
0-
02
b110 6
#458690000000
1!
1%
1-
12
#458700000000
0!
0%
b111 *
0-
02
b111 6
#458710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#458720000000
0!
0%
b0 *
0-
02
b0 6
#458730000000
1!
1%
1-
12
#458740000000
0!
0%
b1 *
0-
02
b1 6
#458750000000
1!
1%
1-
12
#458760000000
0!
0%
b10 *
0-
02
b10 6
#458770000000
1!
1%
1-
12
#458780000000
0!
0%
b11 *
0-
02
b11 6
#458790000000
1!
1%
1-
12
15
#458800000000
0!
0%
b100 *
0-
02
b100 6
#458810000000
1!
1%
1-
12
#458820000000
0!
0%
b101 *
0-
02
b101 6
#458830000000
1!
1%
1-
12
#458840000000
0!
0%
b110 *
0-
02
b110 6
#458850000000
1!
1%
1-
12
#458860000000
0!
0%
b111 *
0-
02
b111 6
#458870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#458880000000
0!
0%
b0 *
0-
02
b0 6
#458890000000
1!
1%
1-
12
#458900000000
0!
0%
b1 *
0-
02
b1 6
#458910000000
1!
1%
1-
12
#458920000000
0!
0%
b10 *
0-
02
b10 6
#458930000000
1!
1%
1-
12
#458940000000
0!
0%
b11 *
0-
02
b11 6
#458950000000
1!
1%
1-
12
15
#458960000000
0!
0%
b100 *
0-
02
b100 6
#458970000000
1!
1%
1-
12
#458980000000
0!
0%
b101 *
0-
02
b101 6
#458990000000
1!
1%
1-
12
#459000000000
0!
0%
b110 *
0-
02
b110 6
#459010000000
1!
1%
1-
12
#459020000000
0!
0%
b111 *
0-
02
b111 6
#459030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#459040000000
0!
0%
b0 *
0-
02
b0 6
#459050000000
1!
1%
1-
12
#459060000000
0!
0%
b1 *
0-
02
b1 6
#459070000000
1!
1%
1-
12
#459080000000
0!
0%
b10 *
0-
02
b10 6
#459090000000
1!
1%
1-
12
#459100000000
0!
0%
b11 *
0-
02
b11 6
#459110000000
1!
1%
1-
12
15
#459120000000
0!
0%
b100 *
0-
02
b100 6
#459130000000
1!
1%
1-
12
#459140000000
0!
0%
b101 *
0-
02
b101 6
#459150000000
1!
1%
1-
12
#459160000000
0!
0%
b110 *
0-
02
b110 6
#459170000000
1!
1%
1-
12
#459180000000
0!
0%
b111 *
0-
02
b111 6
#459190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#459200000000
0!
0%
b0 *
0-
02
b0 6
#459210000000
1!
1%
1-
12
#459220000000
0!
0%
b1 *
0-
02
b1 6
#459230000000
1!
1%
1-
12
#459240000000
0!
0%
b10 *
0-
02
b10 6
#459250000000
1!
1%
1-
12
#459260000000
0!
0%
b11 *
0-
02
b11 6
#459270000000
1!
1%
1-
12
15
#459280000000
0!
0%
b100 *
0-
02
b100 6
#459290000000
1!
1%
1-
12
#459300000000
0!
0%
b101 *
0-
02
b101 6
#459310000000
1!
1%
1-
12
#459320000000
0!
0%
b110 *
0-
02
b110 6
#459330000000
1!
1%
1-
12
#459340000000
0!
0%
b111 *
0-
02
b111 6
#459350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#459360000000
0!
0%
b0 *
0-
02
b0 6
#459370000000
1!
1%
1-
12
#459380000000
0!
0%
b1 *
0-
02
b1 6
#459390000000
1!
1%
1-
12
#459400000000
0!
0%
b10 *
0-
02
b10 6
#459410000000
1!
1%
1-
12
#459420000000
0!
0%
b11 *
0-
02
b11 6
#459430000000
1!
1%
1-
12
15
#459440000000
0!
0%
b100 *
0-
02
b100 6
#459450000000
1!
1%
1-
12
#459460000000
0!
0%
b101 *
0-
02
b101 6
#459470000000
1!
1%
1-
12
#459480000000
0!
0%
b110 *
0-
02
b110 6
#459490000000
1!
1%
1-
12
#459500000000
0!
0%
b111 *
0-
02
b111 6
#459510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#459520000000
0!
0%
b0 *
0-
02
b0 6
#459530000000
1!
1%
1-
12
#459540000000
0!
0%
b1 *
0-
02
b1 6
#459550000000
1!
1%
1-
12
#459560000000
0!
0%
b10 *
0-
02
b10 6
#459570000000
1!
1%
1-
12
#459580000000
0!
0%
b11 *
0-
02
b11 6
#459590000000
1!
1%
1-
12
15
#459600000000
0!
0%
b100 *
0-
02
b100 6
#459610000000
1!
1%
1-
12
#459620000000
0!
0%
b101 *
0-
02
b101 6
#459630000000
1!
1%
1-
12
#459640000000
0!
0%
b110 *
0-
02
b110 6
#459650000000
1!
1%
1-
12
#459660000000
0!
0%
b111 *
0-
02
b111 6
#459670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#459680000000
0!
0%
b0 *
0-
02
b0 6
#459690000000
1!
1%
1-
12
#459700000000
0!
0%
b1 *
0-
02
b1 6
#459710000000
1!
1%
1-
12
#459720000000
0!
0%
b10 *
0-
02
b10 6
#459730000000
1!
1%
1-
12
#459740000000
0!
0%
b11 *
0-
02
b11 6
#459750000000
1!
1%
1-
12
15
#459760000000
0!
0%
b100 *
0-
02
b100 6
#459770000000
1!
1%
1-
12
#459780000000
0!
0%
b101 *
0-
02
b101 6
#459790000000
1!
1%
1-
12
#459800000000
0!
0%
b110 *
0-
02
b110 6
#459810000000
1!
1%
1-
12
#459820000000
0!
0%
b111 *
0-
02
b111 6
#459830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#459840000000
0!
0%
b0 *
0-
02
b0 6
#459850000000
1!
1%
1-
12
#459860000000
0!
0%
b1 *
0-
02
b1 6
#459870000000
1!
1%
1-
12
#459880000000
0!
0%
b10 *
0-
02
b10 6
#459890000000
1!
1%
1-
12
#459900000000
0!
0%
b11 *
0-
02
b11 6
#459910000000
1!
1%
1-
12
15
#459920000000
0!
0%
b100 *
0-
02
b100 6
#459930000000
1!
1%
1-
12
#459940000000
0!
0%
b101 *
0-
02
b101 6
#459950000000
1!
1%
1-
12
#459960000000
0!
0%
b110 *
0-
02
b110 6
#459970000000
1!
1%
1-
12
#459980000000
0!
0%
b111 *
0-
02
b111 6
#459990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#460000000000
0!
0%
b0 *
0-
02
b0 6
#460010000000
1!
1%
1-
12
#460020000000
0!
0%
b1 *
0-
02
b1 6
#460030000000
1!
1%
1-
12
#460040000000
0!
0%
b10 *
0-
02
b10 6
#460050000000
1!
1%
1-
12
#460060000000
0!
0%
b11 *
0-
02
b11 6
#460070000000
1!
1%
1-
12
15
#460080000000
0!
0%
b100 *
0-
02
b100 6
#460090000000
1!
1%
1-
12
#460100000000
0!
0%
b101 *
0-
02
b101 6
#460110000000
1!
1%
1-
12
#460120000000
0!
0%
b110 *
0-
02
b110 6
#460130000000
1!
1%
1-
12
#460140000000
0!
0%
b111 *
0-
02
b111 6
#460150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#460160000000
0!
0%
b0 *
0-
02
b0 6
#460170000000
1!
1%
1-
12
#460180000000
0!
0%
b1 *
0-
02
b1 6
#460190000000
1!
1%
1-
12
#460200000000
0!
0%
b10 *
0-
02
b10 6
#460210000000
1!
1%
1-
12
#460220000000
0!
0%
b11 *
0-
02
b11 6
#460230000000
1!
1%
1-
12
15
#460240000000
0!
0%
b100 *
0-
02
b100 6
#460250000000
1!
1%
1-
12
#460260000000
0!
0%
b101 *
0-
02
b101 6
#460270000000
1!
1%
1-
12
#460280000000
0!
0%
b110 *
0-
02
b110 6
#460290000000
1!
1%
1-
12
#460300000000
0!
0%
b111 *
0-
02
b111 6
#460310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#460320000000
0!
0%
b0 *
0-
02
b0 6
#460330000000
1!
1%
1-
12
#460340000000
0!
0%
b1 *
0-
02
b1 6
#460350000000
1!
1%
1-
12
#460360000000
0!
0%
b10 *
0-
02
b10 6
#460370000000
1!
1%
1-
12
#460380000000
0!
0%
b11 *
0-
02
b11 6
#460390000000
1!
1%
1-
12
15
#460400000000
0!
0%
b100 *
0-
02
b100 6
#460410000000
1!
1%
1-
12
#460420000000
0!
0%
b101 *
0-
02
b101 6
#460430000000
1!
1%
1-
12
#460440000000
0!
0%
b110 *
0-
02
b110 6
#460450000000
1!
1%
1-
12
#460460000000
0!
0%
b111 *
0-
02
b111 6
#460470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#460480000000
0!
0%
b0 *
0-
02
b0 6
#460490000000
1!
1%
1-
12
#460500000000
0!
0%
b1 *
0-
02
b1 6
#460510000000
1!
1%
1-
12
#460520000000
0!
0%
b10 *
0-
02
b10 6
#460530000000
1!
1%
1-
12
#460540000000
0!
0%
b11 *
0-
02
b11 6
#460550000000
1!
1%
1-
12
15
#460560000000
0!
0%
b100 *
0-
02
b100 6
#460570000000
1!
1%
1-
12
#460580000000
0!
0%
b101 *
0-
02
b101 6
#460590000000
1!
1%
1-
12
#460600000000
0!
0%
b110 *
0-
02
b110 6
#460610000000
1!
1%
1-
12
#460620000000
0!
0%
b111 *
0-
02
b111 6
#460630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#460640000000
0!
0%
b0 *
0-
02
b0 6
#460650000000
1!
1%
1-
12
#460660000000
0!
0%
b1 *
0-
02
b1 6
#460670000000
1!
1%
1-
12
#460680000000
0!
0%
b10 *
0-
02
b10 6
#460690000000
1!
1%
1-
12
#460700000000
0!
0%
b11 *
0-
02
b11 6
#460710000000
1!
1%
1-
12
15
#460720000000
0!
0%
b100 *
0-
02
b100 6
#460730000000
1!
1%
1-
12
#460740000000
0!
0%
b101 *
0-
02
b101 6
#460750000000
1!
1%
1-
12
#460760000000
0!
0%
b110 *
0-
02
b110 6
#460770000000
1!
1%
1-
12
#460780000000
0!
0%
b111 *
0-
02
b111 6
#460790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#460800000000
0!
0%
b0 *
0-
02
b0 6
#460810000000
1!
1%
1-
12
#460820000000
0!
0%
b1 *
0-
02
b1 6
#460830000000
1!
1%
1-
12
#460840000000
0!
0%
b10 *
0-
02
b10 6
#460850000000
1!
1%
1-
12
#460860000000
0!
0%
b11 *
0-
02
b11 6
#460870000000
1!
1%
1-
12
15
#460880000000
0!
0%
b100 *
0-
02
b100 6
#460890000000
1!
1%
1-
12
#460900000000
0!
0%
b101 *
0-
02
b101 6
#460910000000
1!
1%
1-
12
#460920000000
0!
0%
b110 *
0-
02
b110 6
#460930000000
1!
1%
1-
12
#460940000000
0!
0%
b111 *
0-
02
b111 6
#460950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#460960000000
0!
0%
b0 *
0-
02
b0 6
#460970000000
1!
1%
1-
12
#460980000000
0!
0%
b1 *
0-
02
b1 6
#460990000000
1!
1%
1-
12
#461000000000
0!
0%
b10 *
0-
02
b10 6
#461010000000
1!
1%
1-
12
#461020000000
0!
0%
b11 *
0-
02
b11 6
#461030000000
1!
1%
1-
12
15
#461040000000
0!
0%
b100 *
0-
02
b100 6
#461050000000
1!
1%
1-
12
#461060000000
0!
0%
b101 *
0-
02
b101 6
#461070000000
1!
1%
1-
12
#461080000000
0!
0%
b110 *
0-
02
b110 6
#461090000000
1!
1%
1-
12
#461100000000
0!
0%
b111 *
0-
02
b111 6
#461110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#461120000000
0!
0%
b0 *
0-
02
b0 6
#461130000000
1!
1%
1-
12
#461140000000
0!
0%
b1 *
0-
02
b1 6
#461150000000
1!
1%
1-
12
#461160000000
0!
0%
b10 *
0-
02
b10 6
#461170000000
1!
1%
1-
12
#461180000000
0!
0%
b11 *
0-
02
b11 6
#461190000000
1!
1%
1-
12
15
#461200000000
0!
0%
b100 *
0-
02
b100 6
#461210000000
1!
1%
1-
12
#461220000000
0!
0%
b101 *
0-
02
b101 6
#461230000000
1!
1%
1-
12
#461240000000
0!
0%
b110 *
0-
02
b110 6
#461250000000
1!
1%
1-
12
#461260000000
0!
0%
b111 *
0-
02
b111 6
#461270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#461280000000
0!
0%
b0 *
0-
02
b0 6
#461290000000
1!
1%
1-
12
#461300000000
0!
0%
b1 *
0-
02
b1 6
#461310000000
1!
1%
1-
12
#461320000000
0!
0%
b10 *
0-
02
b10 6
#461330000000
1!
1%
1-
12
#461340000000
0!
0%
b11 *
0-
02
b11 6
#461350000000
1!
1%
1-
12
15
#461360000000
0!
0%
b100 *
0-
02
b100 6
#461370000000
1!
1%
1-
12
#461380000000
0!
0%
b101 *
0-
02
b101 6
#461390000000
1!
1%
1-
12
#461400000000
0!
0%
b110 *
0-
02
b110 6
#461410000000
1!
1%
1-
12
#461420000000
0!
0%
b111 *
0-
02
b111 6
#461430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#461440000000
0!
0%
b0 *
0-
02
b0 6
#461450000000
1!
1%
1-
12
#461460000000
0!
0%
b1 *
0-
02
b1 6
#461470000000
1!
1%
1-
12
#461480000000
0!
0%
b10 *
0-
02
b10 6
#461490000000
1!
1%
1-
12
#461500000000
0!
0%
b11 *
0-
02
b11 6
#461510000000
1!
1%
1-
12
15
#461520000000
0!
0%
b100 *
0-
02
b100 6
#461530000000
1!
1%
1-
12
#461540000000
0!
0%
b101 *
0-
02
b101 6
#461550000000
1!
1%
1-
12
#461560000000
0!
0%
b110 *
0-
02
b110 6
#461570000000
1!
1%
1-
12
#461580000000
0!
0%
b111 *
0-
02
b111 6
#461590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#461600000000
0!
0%
b0 *
0-
02
b0 6
#461610000000
1!
1%
1-
12
#461620000000
0!
0%
b1 *
0-
02
b1 6
#461630000000
1!
1%
1-
12
#461640000000
0!
0%
b10 *
0-
02
b10 6
#461650000000
1!
1%
1-
12
#461660000000
0!
0%
b11 *
0-
02
b11 6
#461670000000
1!
1%
1-
12
15
#461680000000
0!
0%
b100 *
0-
02
b100 6
#461690000000
1!
1%
1-
12
#461700000000
0!
0%
b101 *
0-
02
b101 6
#461710000000
1!
1%
1-
12
#461720000000
0!
0%
b110 *
0-
02
b110 6
#461730000000
1!
1%
1-
12
#461740000000
0!
0%
b111 *
0-
02
b111 6
#461750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#461760000000
0!
0%
b0 *
0-
02
b0 6
#461770000000
1!
1%
1-
12
#461780000000
0!
0%
b1 *
0-
02
b1 6
#461790000000
1!
1%
1-
12
#461800000000
0!
0%
b10 *
0-
02
b10 6
#461810000000
1!
1%
1-
12
#461820000000
0!
0%
b11 *
0-
02
b11 6
#461830000000
1!
1%
1-
12
15
#461840000000
0!
0%
b100 *
0-
02
b100 6
#461850000000
1!
1%
1-
12
#461860000000
0!
0%
b101 *
0-
02
b101 6
#461870000000
1!
1%
1-
12
#461880000000
0!
0%
b110 *
0-
02
b110 6
#461890000000
1!
1%
1-
12
#461900000000
0!
0%
b111 *
0-
02
b111 6
#461910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#461920000000
0!
0%
b0 *
0-
02
b0 6
#461930000000
1!
1%
1-
12
#461940000000
0!
0%
b1 *
0-
02
b1 6
#461950000000
1!
1%
1-
12
#461960000000
0!
0%
b10 *
0-
02
b10 6
#461970000000
1!
1%
1-
12
#461980000000
0!
0%
b11 *
0-
02
b11 6
#461990000000
1!
1%
1-
12
15
#462000000000
0!
0%
b100 *
0-
02
b100 6
#462010000000
1!
1%
1-
12
#462020000000
0!
0%
b101 *
0-
02
b101 6
#462030000000
1!
1%
1-
12
#462040000000
0!
0%
b110 *
0-
02
b110 6
#462050000000
1!
1%
1-
12
#462060000000
0!
0%
b111 *
0-
02
b111 6
#462070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#462080000000
0!
0%
b0 *
0-
02
b0 6
#462090000000
1!
1%
1-
12
#462100000000
0!
0%
b1 *
0-
02
b1 6
#462110000000
1!
1%
1-
12
#462120000000
0!
0%
b10 *
0-
02
b10 6
#462130000000
1!
1%
1-
12
#462140000000
0!
0%
b11 *
0-
02
b11 6
#462150000000
1!
1%
1-
12
15
#462160000000
0!
0%
b100 *
0-
02
b100 6
#462170000000
1!
1%
1-
12
#462180000000
0!
0%
b101 *
0-
02
b101 6
#462190000000
1!
1%
1-
12
#462200000000
0!
0%
b110 *
0-
02
b110 6
#462210000000
1!
1%
1-
12
#462220000000
0!
0%
b111 *
0-
02
b111 6
#462230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#462240000000
0!
0%
b0 *
0-
02
b0 6
#462250000000
1!
1%
1-
12
#462260000000
0!
0%
b1 *
0-
02
b1 6
#462270000000
1!
1%
1-
12
#462280000000
0!
0%
b10 *
0-
02
b10 6
#462290000000
1!
1%
1-
12
#462300000000
0!
0%
b11 *
0-
02
b11 6
#462310000000
1!
1%
1-
12
15
#462320000000
0!
0%
b100 *
0-
02
b100 6
#462330000000
1!
1%
1-
12
#462340000000
0!
0%
b101 *
0-
02
b101 6
#462350000000
1!
1%
1-
12
#462360000000
0!
0%
b110 *
0-
02
b110 6
#462370000000
1!
1%
1-
12
#462380000000
0!
0%
b111 *
0-
02
b111 6
#462390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#462400000000
0!
0%
b0 *
0-
02
b0 6
#462410000000
1!
1%
1-
12
#462420000000
0!
0%
b1 *
0-
02
b1 6
#462430000000
1!
1%
1-
12
#462440000000
0!
0%
b10 *
0-
02
b10 6
#462450000000
1!
1%
1-
12
#462460000000
0!
0%
b11 *
0-
02
b11 6
#462470000000
1!
1%
1-
12
15
#462480000000
0!
0%
b100 *
0-
02
b100 6
#462490000000
1!
1%
1-
12
#462500000000
0!
0%
b101 *
0-
02
b101 6
#462510000000
1!
1%
1-
12
#462520000000
0!
0%
b110 *
0-
02
b110 6
#462530000000
1!
1%
1-
12
#462540000000
0!
0%
b111 *
0-
02
b111 6
#462550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#462560000000
0!
0%
b0 *
0-
02
b0 6
#462570000000
1!
1%
1-
12
#462580000000
0!
0%
b1 *
0-
02
b1 6
#462590000000
1!
1%
1-
12
#462600000000
0!
0%
b10 *
0-
02
b10 6
#462610000000
1!
1%
1-
12
#462620000000
0!
0%
b11 *
0-
02
b11 6
#462630000000
1!
1%
1-
12
15
#462640000000
0!
0%
b100 *
0-
02
b100 6
#462650000000
1!
1%
1-
12
#462660000000
0!
0%
b101 *
0-
02
b101 6
#462670000000
1!
1%
1-
12
#462680000000
0!
0%
b110 *
0-
02
b110 6
#462690000000
1!
1%
1-
12
#462700000000
0!
0%
b111 *
0-
02
b111 6
#462710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#462720000000
0!
0%
b0 *
0-
02
b0 6
#462730000000
1!
1%
1-
12
#462740000000
0!
0%
b1 *
0-
02
b1 6
#462750000000
1!
1%
1-
12
#462760000000
0!
0%
b10 *
0-
02
b10 6
#462770000000
1!
1%
1-
12
#462780000000
0!
0%
b11 *
0-
02
b11 6
#462790000000
1!
1%
1-
12
15
#462800000000
0!
0%
b100 *
0-
02
b100 6
#462810000000
1!
1%
1-
12
#462820000000
0!
0%
b101 *
0-
02
b101 6
#462830000000
1!
1%
1-
12
#462840000000
0!
0%
b110 *
0-
02
b110 6
#462850000000
1!
1%
1-
12
#462860000000
0!
0%
b111 *
0-
02
b111 6
#462870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#462880000000
0!
0%
b0 *
0-
02
b0 6
#462890000000
1!
1%
1-
12
#462900000000
0!
0%
b1 *
0-
02
b1 6
#462910000000
1!
1%
1-
12
#462920000000
0!
0%
b10 *
0-
02
b10 6
#462930000000
1!
1%
1-
12
#462940000000
0!
0%
b11 *
0-
02
b11 6
#462950000000
1!
1%
1-
12
15
#462960000000
0!
0%
b100 *
0-
02
b100 6
#462970000000
1!
1%
1-
12
#462980000000
0!
0%
b101 *
0-
02
b101 6
#462990000000
1!
1%
1-
12
#463000000000
0!
0%
b110 *
0-
02
b110 6
#463010000000
1!
1%
1-
12
#463020000000
0!
0%
b111 *
0-
02
b111 6
#463030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#463040000000
0!
0%
b0 *
0-
02
b0 6
#463050000000
1!
1%
1-
12
#463060000000
0!
0%
b1 *
0-
02
b1 6
#463070000000
1!
1%
1-
12
#463080000000
0!
0%
b10 *
0-
02
b10 6
#463090000000
1!
1%
1-
12
#463100000000
0!
0%
b11 *
0-
02
b11 6
#463110000000
1!
1%
1-
12
15
#463120000000
0!
0%
b100 *
0-
02
b100 6
#463130000000
1!
1%
1-
12
#463140000000
0!
0%
b101 *
0-
02
b101 6
#463150000000
1!
1%
1-
12
#463160000000
0!
0%
b110 *
0-
02
b110 6
#463170000000
1!
1%
1-
12
#463180000000
0!
0%
b111 *
0-
02
b111 6
#463190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#463200000000
0!
0%
b0 *
0-
02
b0 6
#463210000000
1!
1%
1-
12
#463220000000
0!
0%
b1 *
0-
02
b1 6
#463230000000
1!
1%
1-
12
#463240000000
0!
0%
b10 *
0-
02
b10 6
#463250000000
1!
1%
1-
12
#463260000000
0!
0%
b11 *
0-
02
b11 6
#463270000000
1!
1%
1-
12
15
#463280000000
0!
0%
b100 *
0-
02
b100 6
#463290000000
1!
1%
1-
12
#463300000000
0!
0%
b101 *
0-
02
b101 6
#463310000000
1!
1%
1-
12
#463320000000
0!
0%
b110 *
0-
02
b110 6
#463330000000
1!
1%
1-
12
#463340000000
0!
0%
b111 *
0-
02
b111 6
#463350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#463360000000
0!
0%
b0 *
0-
02
b0 6
#463370000000
1!
1%
1-
12
#463380000000
0!
0%
b1 *
0-
02
b1 6
#463390000000
1!
1%
1-
12
#463400000000
0!
0%
b10 *
0-
02
b10 6
#463410000000
1!
1%
1-
12
#463420000000
0!
0%
b11 *
0-
02
b11 6
#463430000000
1!
1%
1-
12
15
#463440000000
0!
0%
b100 *
0-
02
b100 6
#463450000000
1!
1%
1-
12
#463460000000
0!
0%
b101 *
0-
02
b101 6
#463470000000
1!
1%
1-
12
#463480000000
0!
0%
b110 *
0-
02
b110 6
#463490000000
1!
1%
1-
12
#463500000000
0!
0%
b111 *
0-
02
b111 6
#463510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#463520000000
0!
0%
b0 *
0-
02
b0 6
#463530000000
1!
1%
1-
12
#463540000000
0!
0%
b1 *
0-
02
b1 6
#463550000000
1!
1%
1-
12
#463560000000
0!
0%
b10 *
0-
02
b10 6
#463570000000
1!
1%
1-
12
#463580000000
0!
0%
b11 *
0-
02
b11 6
#463590000000
1!
1%
1-
12
15
#463600000000
0!
0%
b100 *
0-
02
b100 6
#463610000000
1!
1%
1-
12
#463620000000
0!
0%
b101 *
0-
02
b101 6
#463630000000
1!
1%
1-
12
#463640000000
0!
0%
b110 *
0-
02
b110 6
#463650000000
1!
1%
1-
12
#463660000000
0!
0%
b111 *
0-
02
b111 6
#463670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#463680000000
0!
0%
b0 *
0-
02
b0 6
#463690000000
1!
1%
1-
12
#463700000000
0!
0%
b1 *
0-
02
b1 6
#463710000000
1!
1%
1-
12
#463720000000
0!
0%
b10 *
0-
02
b10 6
#463730000000
1!
1%
1-
12
#463740000000
0!
0%
b11 *
0-
02
b11 6
#463750000000
1!
1%
1-
12
15
#463760000000
0!
0%
b100 *
0-
02
b100 6
#463770000000
1!
1%
1-
12
#463780000000
0!
0%
b101 *
0-
02
b101 6
#463790000000
1!
1%
1-
12
#463800000000
0!
0%
b110 *
0-
02
b110 6
#463810000000
1!
1%
1-
12
#463820000000
0!
0%
b111 *
0-
02
b111 6
#463830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#463840000000
0!
0%
b0 *
0-
02
b0 6
#463850000000
1!
1%
1-
12
#463860000000
0!
0%
b1 *
0-
02
b1 6
#463870000000
1!
1%
1-
12
#463880000000
0!
0%
b10 *
0-
02
b10 6
#463890000000
1!
1%
1-
12
#463900000000
0!
0%
b11 *
0-
02
b11 6
#463910000000
1!
1%
1-
12
15
#463920000000
0!
0%
b100 *
0-
02
b100 6
#463930000000
1!
1%
1-
12
#463940000000
0!
0%
b101 *
0-
02
b101 6
#463950000000
1!
1%
1-
12
#463960000000
0!
0%
b110 *
0-
02
b110 6
#463970000000
1!
1%
1-
12
#463980000000
0!
0%
b111 *
0-
02
b111 6
#463990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#464000000000
0!
0%
b0 *
0-
02
b0 6
#464010000000
1!
1%
1-
12
#464020000000
0!
0%
b1 *
0-
02
b1 6
#464030000000
1!
1%
1-
12
#464040000000
0!
0%
b10 *
0-
02
b10 6
#464050000000
1!
1%
1-
12
#464060000000
0!
0%
b11 *
0-
02
b11 6
#464070000000
1!
1%
1-
12
15
#464080000000
0!
0%
b100 *
0-
02
b100 6
#464090000000
1!
1%
1-
12
#464100000000
0!
0%
b101 *
0-
02
b101 6
#464110000000
1!
1%
1-
12
#464120000000
0!
0%
b110 *
0-
02
b110 6
#464130000000
1!
1%
1-
12
#464140000000
0!
0%
b111 *
0-
02
b111 6
#464150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#464160000000
0!
0%
b0 *
0-
02
b0 6
#464170000000
1!
1%
1-
12
#464180000000
0!
0%
b1 *
0-
02
b1 6
#464190000000
1!
1%
1-
12
#464200000000
0!
0%
b10 *
0-
02
b10 6
#464210000000
1!
1%
1-
12
#464220000000
0!
0%
b11 *
0-
02
b11 6
#464230000000
1!
1%
1-
12
15
#464240000000
0!
0%
b100 *
0-
02
b100 6
#464250000000
1!
1%
1-
12
#464260000000
0!
0%
b101 *
0-
02
b101 6
#464270000000
1!
1%
1-
12
#464280000000
0!
0%
b110 *
0-
02
b110 6
#464290000000
1!
1%
1-
12
#464300000000
0!
0%
b111 *
0-
02
b111 6
#464310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#464320000000
0!
0%
b0 *
0-
02
b0 6
#464330000000
1!
1%
1-
12
#464340000000
0!
0%
b1 *
0-
02
b1 6
#464350000000
1!
1%
1-
12
#464360000000
0!
0%
b10 *
0-
02
b10 6
#464370000000
1!
1%
1-
12
#464380000000
0!
0%
b11 *
0-
02
b11 6
#464390000000
1!
1%
1-
12
15
#464400000000
0!
0%
b100 *
0-
02
b100 6
#464410000000
1!
1%
1-
12
#464420000000
0!
0%
b101 *
0-
02
b101 6
#464430000000
1!
1%
1-
12
#464440000000
0!
0%
b110 *
0-
02
b110 6
#464450000000
1!
1%
1-
12
#464460000000
0!
0%
b111 *
0-
02
b111 6
#464470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#464480000000
0!
0%
b0 *
0-
02
b0 6
#464490000000
1!
1%
1-
12
#464500000000
0!
0%
b1 *
0-
02
b1 6
#464510000000
1!
1%
1-
12
#464520000000
0!
0%
b10 *
0-
02
b10 6
#464530000000
1!
1%
1-
12
#464540000000
0!
0%
b11 *
0-
02
b11 6
#464550000000
1!
1%
1-
12
15
#464560000000
0!
0%
b100 *
0-
02
b100 6
#464570000000
1!
1%
1-
12
#464580000000
0!
0%
b101 *
0-
02
b101 6
#464590000000
1!
1%
1-
12
#464600000000
0!
0%
b110 *
0-
02
b110 6
#464610000000
1!
1%
1-
12
#464620000000
0!
0%
b111 *
0-
02
b111 6
#464630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#464640000000
0!
0%
b0 *
0-
02
b0 6
#464650000000
1!
1%
1-
12
#464660000000
0!
0%
b1 *
0-
02
b1 6
#464670000000
1!
1%
1-
12
#464680000000
0!
0%
b10 *
0-
02
b10 6
#464690000000
1!
1%
1-
12
#464700000000
0!
0%
b11 *
0-
02
b11 6
#464710000000
1!
1%
1-
12
15
#464720000000
0!
0%
b100 *
0-
02
b100 6
#464730000000
1!
1%
1-
12
#464740000000
0!
0%
b101 *
0-
02
b101 6
#464750000000
1!
1%
1-
12
#464760000000
0!
0%
b110 *
0-
02
b110 6
#464770000000
1!
1%
1-
12
#464780000000
0!
0%
b111 *
0-
02
b111 6
#464790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#464800000000
0!
0%
b0 *
0-
02
b0 6
#464810000000
1!
1%
1-
12
#464820000000
0!
0%
b1 *
0-
02
b1 6
#464830000000
1!
1%
1-
12
#464840000000
0!
0%
b10 *
0-
02
b10 6
#464850000000
1!
1%
1-
12
#464860000000
0!
0%
b11 *
0-
02
b11 6
#464870000000
1!
1%
1-
12
15
#464880000000
0!
0%
b100 *
0-
02
b100 6
#464890000000
1!
1%
1-
12
#464900000000
0!
0%
b101 *
0-
02
b101 6
#464910000000
1!
1%
1-
12
#464920000000
0!
0%
b110 *
0-
02
b110 6
#464930000000
1!
1%
1-
12
#464940000000
0!
0%
b111 *
0-
02
b111 6
#464950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#464960000000
0!
0%
b0 *
0-
02
b0 6
#464970000000
1!
1%
1-
12
#464980000000
0!
0%
b1 *
0-
02
b1 6
#464990000000
1!
1%
1-
12
#465000000000
0!
0%
b10 *
0-
02
b10 6
#465010000000
1!
1%
1-
12
#465020000000
0!
0%
b11 *
0-
02
b11 6
#465030000000
1!
1%
1-
12
15
#465040000000
0!
0%
b100 *
0-
02
b100 6
#465050000000
1!
1%
1-
12
#465060000000
0!
0%
b101 *
0-
02
b101 6
#465070000000
1!
1%
1-
12
#465080000000
0!
0%
b110 *
0-
02
b110 6
#465090000000
1!
1%
1-
12
#465100000000
0!
0%
b111 *
0-
02
b111 6
#465110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#465120000000
0!
0%
b0 *
0-
02
b0 6
#465130000000
1!
1%
1-
12
#465140000000
0!
0%
b1 *
0-
02
b1 6
#465150000000
1!
1%
1-
12
#465160000000
0!
0%
b10 *
0-
02
b10 6
#465170000000
1!
1%
1-
12
#465180000000
0!
0%
b11 *
0-
02
b11 6
#465190000000
1!
1%
1-
12
15
#465200000000
0!
0%
b100 *
0-
02
b100 6
#465210000000
1!
1%
1-
12
#465220000000
0!
0%
b101 *
0-
02
b101 6
#465230000000
1!
1%
1-
12
#465240000000
0!
0%
b110 *
0-
02
b110 6
#465250000000
1!
1%
1-
12
#465260000000
0!
0%
b111 *
0-
02
b111 6
#465270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#465280000000
0!
0%
b0 *
0-
02
b0 6
#465290000000
1!
1%
1-
12
#465300000000
0!
0%
b1 *
0-
02
b1 6
#465310000000
1!
1%
1-
12
#465320000000
0!
0%
b10 *
0-
02
b10 6
#465330000000
1!
1%
1-
12
#465340000000
0!
0%
b11 *
0-
02
b11 6
#465350000000
1!
1%
1-
12
15
#465360000000
0!
0%
b100 *
0-
02
b100 6
#465370000000
1!
1%
1-
12
#465380000000
0!
0%
b101 *
0-
02
b101 6
#465390000000
1!
1%
1-
12
#465400000000
0!
0%
b110 *
0-
02
b110 6
#465410000000
1!
1%
1-
12
#465420000000
0!
0%
b111 *
0-
02
b111 6
#465430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#465440000000
0!
0%
b0 *
0-
02
b0 6
#465450000000
1!
1%
1-
12
#465460000000
0!
0%
b1 *
0-
02
b1 6
#465470000000
1!
1%
1-
12
#465480000000
0!
0%
b10 *
0-
02
b10 6
#465490000000
1!
1%
1-
12
#465500000000
0!
0%
b11 *
0-
02
b11 6
#465510000000
1!
1%
1-
12
15
#465520000000
0!
0%
b100 *
0-
02
b100 6
#465530000000
1!
1%
1-
12
#465540000000
0!
0%
b101 *
0-
02
b101 6
#465550000000
1!
1%
1-
12
#465560000000
0!
0%
b110 *
0-
02
b110 6
#465570000000
1!
1%
1-
12
#465580000000
0!
0%
b111 *
0-
02
b111 6
#465590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#465600000000
0!
0%
b0 *
0-
02
b0 6
#465610000000
1!
1%
1-
12
#465620000000
0!
0%
b1 *
0-
02
b1 6
#465630000000
1!
1%
1-
12
#465640000000
0!
0%
b10 *
0-
02
b10 6
#465650000000
1!
1%
1-
12
#465660000000
0!
0%
b11 *
0-
02
b11 6
#465670000000
1!
1%
1-
12
15
#465680000000
0!
0%
b100 *
0-
02
b100 6
#465690000000
1!
1%
1-
12
#465700000000
0!
0%
b101 *
0-
02
b101 6
#465710000000
1!
1%
1-
12
#465720000000
0!
0%
b110 *
0-
02
b110 6
#465730000000
1!
1%
1-
12
#465740000000
0!
0%
b111 *
0-
02
b111 6
#465750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#465760000000
0!
0%
b0 *
0-
02
b0 6
#465770000000
1!
1%
1-
12
#465780000000
0!
0%
b1 *
0-
02
b1 6
#465790000000
1!
1%
1-
12
#465800000000
0!
0%
b10 *
0-
02
b10 6
#465810000000
1!
1%
1-
12
#465820000000
0!
0%
b11 *
0-
02
b11 6
#465830000000
1!
1%
1-
12
15
#465840000000
0!
0%
b100 *
0-
02
b100 6
#465850000000
1!
1%
1-
12
#465860000000
0!
0%
b101 *
0-
02
b101 6
#465870000000
1!
1%
1-
12
#465880000000
0!
0%
b110 *
0-
02
b110 6
#465890000000
1!
1%
1-
12
#465900000000
0!
0%
b111 *
0-
02
b111 6
#465910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#465920000000
0!
0%
b0 *
0-
02
b0 6
#465930000000
1!
1%
1-
12
#465940000000
0!
0%
b1 *
0-
02
b1 6
#465950000000
1!
1%
1-
12
#465960000000
0!
0%
b10 *
0-
02
b10 6
#465970000000
1!
1%
1-
12
#465980000000
0!
0%
b11 *
0-
02
b11 6
#465990000000
1!
1%
1-
12
15
#466000000000
0!
0%
b100 *
0-
02
b100 6
#466010000000
1!
1%
1-
12
#466020000000
0!
0%
b101 *
0-
02
b101 6
#466030000000
1!
1%
1-
12
#466040000000
0!
0%
b110 *
0-
02
b110 6
#466050000000
1!
1%
1-
12
#466060000000
0!
0%
b111 *
0-
02
b111 6
#466070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#466080000000
0!
0%
b0 *
0-
02
b0 6
#466090000000
1!
1%
1-
12
#466100000000
0!
0%
b1 *
0-
02
b1 6
#466110000000
1!
1%
1-
12
#466120000000
0!
0%
b10 *
0-
02
b10 6
#466130000000
1!
1%
1-
12
#466140000000
0!
0%
b11 *
0-
02
b11 6
#466150000000
1!
1%
1-
12
15
#466160000000
0!
0%
b100 *
0-
02
b100 6
#466170000000
1!
1%
1-
12
#466180000000
0!
0%
b101 *
0-
02
b101 6
#466190000000
1!
1%
1-
12
#466200000000
0!
0%
b110 *
0-
02
b110 6
#466210000000
1!
1%
1-
12
#466220000000
0!
0%
b111 *
0-
02
b111 6
#466230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#466240000000
0!
0%
b0 *
0-
02
b0 6
#466250000000
1!
1%
1-
12
#466260000000
0!
0%
b1 *
0-
02
b1 6
#466270000000
1!
1%
1-
12
#466280000000
0!
0%
b10 *
0-
02
b10 6
#466290000000
1!
1%
1-
12
#466300000000
0!
0%
b11 *
0-
02
b11 6
#466310000000
1!
1%
1-
12
15
#466320000000
0!
0%
b100 *
0-
02
b100 6
#466330000000
1!
1%
1-
12
#466340000000
0!
0%
b101 *
0-
02
b101 6
#466350000000
1!
1%
1-
12
#466360000000
0!
0%
b110 *
0-
02
b110 6
#466370000000
1!
1%
1-
12
#466380000000
0!
0%
b111 *
0-
02
b111 6
#466390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#466400000000
0!
0%
b0 *
0-
02
b0 6
#466410000000
1!
1%
1-
12
#466420000000
0!
0%
b1 *
0-
02
b1 6
#466430000000
1!
1%
1-
12
#466440000000
0!
0%
b10 *
0-
02
b10 6
#466450000000
1!
1%
1-
12
#466460000000
0!
0%
b11 *
0-
02
b11 6
#466470000000
1!
1%
1-
12
15
#466480000000
0!
0%
b100 *
0-
02
b100 6
#466490000000
1!
1%
1-
12
#466500000000
0!
0%
b101 *
0-
02
b101 6
#466510000000
1!
1%
1-
12
#466520000000
0!
0%
b110 *
0-
02
b110 6
#466530000000
1!
1%
1-
12
#466540000000
0!
0%
b111 *
0-
02
b111 6
#466550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#466560000000
0!
0%
b0 *
0-
02
b0 6
#466570000000
1!
1%
1-
12
#466580000000
0!
0%
b1 *
0-
02
b1 6
#466590000000
1!
1%
1-
12
#466600000000
0!
0%
b10 *
0-
02
b10 6
#466610000000
1!
1%
1-
12
#466620000000
0!
0%
b11 *
0-
02
b11 6
#466630000000
1!
1%
1-
12
15
#466640000000
0!
0%
b100 *
0-
02
b100 6
#466650000000
1!
1%
1-
12
#466660000000
0!
0%
b101 *
0-
02
b101 6
#466670000000
1!
1%
1-
12
#466680000000
0!
0%
b110 *
0-
02
b110 6
#466690000000
1!
1%
1-
12
#466700000000
0!
0%
b111 *
0-
02
b111 6
#466710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#466720000000
0!
0%
b0 *
0-
02
b0 6
#466730000000
1!
1%
1-
12
#466740000000
0!
0%
b1 *
0-
02
b1 6
#466750000000
1!
1%
1-
12
#466760000000
0!
0%
b10 *
0-
02
b10 6
#466770000000
1!
1%
1-
12
#466780000000
0!
0%
b11 *
0-
02
b11 6
#466790000000
1!
1%
1-
12
15
#466800000000
0!
0%
b100 *
0-
02
b100 6
#466810000000
1!
1%
1-
12
#466820000000
0!
0%
b101 *
0-
02
b101 6
#466830000000
1!
1%
1-
12
#466840000000
0!
0%
b110 *
0-
02
b110 6
#466850000000
1!
1%
1-
12
#466860000000
0!
0%
b111 *
0-
02
b111 6
#466870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#466880000000
0!
0%
b0 *
0-
02
b0 6
#466890000000
1!
1%
1-
12
#466900000000
0!
0%
b1 *
0-
02
b1 6
#466910000000
1!
1%
1-
12
#466920000000
0!
0%
b10 *
0-
02
b10 6
#466930000000
1!
1%
1-
12
#466940000000
0!
0%
b11 *
0-
02
b11 6
#466950000000
1!
1%
1-
12
15
#466960000000
0!
0%
b100 *
0-
02
b100 6
#466970000000
1!
1%
1-
12
#466980000000
0!
0%
b101 *
0-
02
b101 6
#466990000000
1!
1%
1-
12
#467000000000
0!
0%
b110 *
0-
02
b110 6
#467010000000
1!
1%
1-
12
#467020000000
0!
0%
b111 *
0-
02
b111 6
#467030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#467040000000
0!
0%
b0 *
0-
02
b0 6
#467050000000
1!
1%
1-
12
#467060000000
0!
0%
b1 *
0-
02
b1 6
#467070000000
1!
1%
1-
12
#467080000000
0!
0%
b10 *
0-
02
b10 6
#467090000000
1!
1%
1-
12
#467100000000
0!
0%
b11 *
0-
02
b11 6
#467110000000
1!
1%
1-
12
15
#467120000000
0!
0%
b100 *
0-
02
b100 6
#467130000000
1!
1%
1-
12
#467140000000
0!
0%
b101 *
0-
02
b101 6
#467150000000
1!
1%
1-
12
#467160000000
0!
0%
b110 *
0-
02
b110 6
#467170000000
1!
1%
1-
12
#467180000000
0!
0%
b111 *
0-
02
b111 6
#467190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#467200000000
0!
0%
b0 *
0-
02
b0 6
#467210000000
1!
1%
1-
12
#467220000000
0!
0%
b1 *
0-
02
b1 6
#467230000000
1!
1%
1-
12
#467240000000
0!
0%
b10 *
0-
02
b10 6
#467250000000
1!
1%
1-
12
#467260000000
0!
0%
b11 *
0-
02
b11 6
#467270000000
1!
1%
1-
12
15
#467280000000
0!
0%
b100 *
0-
02
b100 6
#467290000000
1!
1%
1-
12
#467300000000
0!
0%
b101 *
0-
02
b101 6
#467310000000
1!
1%
1-
12
#467320000000
0!
0%
b110 *
0-
02
b110 6
#467330000000
1!
1%
1-
12
#467340000000
0!
0%
b111 *
0-
02
b111 6
#467350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#467360000000
0!
0%
b0 *
0-
02
b0 6
#467370000000
1!
1%
1-
12
#467380000000
0!
0%
b1 *
0-
02
b1 6
#467390000000
1!
1%
1-
12
#467400000000
0!
0%
b10 *
0-
02
b10 6
#467410000000
1!
1%
1-
12
#467420000000
0!
0%
b11 *
0-
02
b11 6
#467430000000
1!
1%
1-
12
15
#467440000000
0!
0%
b100 *
0-
02
b100 6
#467450000000
1!
1%
1-
12
#467460000000
0!
0%
b101 *
0-
02
b101 6
#467470000000
1!
1%
1-
12
#467480000000
0!
0%
b110 *
0-
02
b110 6
#467490000000
1!
1%
1-
12
#467500000000
0!
0%
b111 *
0-
02
b111 6
#467510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#467520000000
0!
0%
b0 *
0-
02
b0 6
#467530000000
1!
1%
1-
12
#467540000000
0!
0%
b1 *
0-
02
b1 6
#467550000000
1!
1%
1-
12
#467560000000
0!
0%
b10 *
0-
02
b10 6
#467570000000
1!
1%
1-
12
#467580000000
0!
0%
b11 *
0-
02
b11 6
#467590000000
1!
1%
1-
12
15
#467600000000
0!
0%
b100 *
0-
02
b100 6
#467610000000
1!
1%
1-
12
#467620000000
0!
0%
b101 *
0-
02
b101 6
#467630000000
1!
1%
1-
12
#467640000000
0!
0%
b110 *
0-
02
b110 6
#467650000000
1!
1%
1-
12
#467660000000
0!
0%
b111 *
0-
02
b111 6
#467670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#467680000000
0!
0%
b0 *
0-
02
b0 6
#467690000000
1!
1%
1-
12
#467700000000
0!
0%
b1 *
0-
02
b1 6
#467710000000
1!
1%
1-
12
#467720000000
0!
0%
b10 *
0-
02
b10 6
#467730000000
1!
1%
1-
12
#467740000000
0!
0%
b11 *
0-
02
b11 6
#467750000000
1!
1%
1-
12
15
#467760000000
0!
0%
b100 *
0-
02
b100 6
#467770000000
1!
1%
1-
12
#467780000000
0!
0%
b101 *
0-
02
b101 6
#467790000000
1!
1%
1-
12
#467800000000
0!
0%
b110 *
0-
02
b110 6
#467810000000
1!
1%
1-
12
#467820000000
0!
0%
b111 *
0-
02
b111 6
#467830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#467840000000
0!
0%
b0 *
0-
02
b0 6
#467850000000
1!
1%
1-
12
#467860000000
0!
0%
b1 *
0-
02
b1 6
#467870000000
1!
1%
1-
12
#467880000000
0!
0%
b10 *
0-
02
b10 6
#467890000000
1!
1%
1-
12
#467900000000
0!
0%
b11 *
0-
02
b11 6
#467910000000
1!
1%
1-
12
15
#467920000000
0!
0%
b100 *
0-
02
b100 6
#467930000000
1!
1%
1-
12
#467940000000
0!
0%
b101 *
0-
02
b101 6
#467950000000
1!
1%
1-
12
#467960000000
0!
0%
b110 *
0-
02
b110 6
#467970000000
1!
1%
1-
12
#467980000000
0!
0%
b111 *
0-
02
b111 6
#467990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#468000000000
0!
0%
b0 *
0-
02
b0 6
#468010000000
1!
1%
1-
12
#468020000000
0!
0%
b1 *
0-
02
b1 6
#468030000000
1!
1%
1-
12
#468040000000
0!
0%
b10 *
0-
02
b10 6
#468050000000
1!
1%
1-
12
#468060000000
0!
0%
b11 *
0-
02
b11 6
#468070000000
1!
1%
1-
12
15
#468080000000
0!
0%
b100 *
0-
02
b100 6
#468090000000
1!
1%
1-
12
#468100000000
0!
0%
b101 *
0-
02
b101 6
#468110000000
1!
1%
1-
12
#468120000000
0!
0%
b110 *
0-
02
b110 6
#468130000000
1!
1%
1-
12
#468140000000
0!
0%
b111 *
0-
02
b111 6
#468150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#468160000000
0!
0%
b0 *
0-
02
b0 6
#468170000000
1!
1%
1-
12
#468180000000
0!
0%
b1 *
0-
02
b1 6
#468190000000
1!
1%
1-
12
#468200000000
0!
0%
b10 *
0-
02
b10 6
#468210000000
1!
1%
1-
12
#468220000000
0!
0%
b11 *
0-
02
b11 6
#468230000000
1!
1%
1-
12
15
#468240000000
0!
0%
b100 *
0-
02
b100 6
#468250000000
1!
1%
1-
12
#468260000000
0!
0%
b101 *
0-
02
b101 6
#468270000000
1!
1%
1-
12
#468280000000
0!
0%
b110 *
0-
02
b110 6
#468290000000
1!
1%
1-
12
#468300000000
0!
0%
b111 *
0-
02
b111 6
#468310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#468320000000
0!
0%
b0 *
0-
02
b0 6
#468330000000
1!
1%
1-
12
#468340000000
0!
0%
b1 *
0-
02
b1 6
#468350000000
1!
1%
1-
12
#468360000000
0!
0%
b10 *
0-
02
b10 6
#468370000000
1!
1%
1-
12
#468380000000
0!
0%
b11 *
0-
02
b11 6
#468390000000
1!
1%
1-
12
15
#468400000000
0!
0%
b100 *
0-
02
b100 6
#468410000000
1!
1%
1-
12
#468420000000
0!
0%
b101 *
0-
02
b101 6
#468430000000
1!
1%
1-
12
#468440000000
0!
0%
b110 *
0-
02
b110 6
#468450000000
1!
1%
1-
12
#468460000000
0!
0%
b111 *
0-
02
b111 6
#468470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#468480000000
0!
0%
b0 *
0-
02
b0 6
#468490000000
1!
1%
1-
12
#468500000000
0!
0%
b1 *
0-
02
b1 6
#468510000000
1!
1%
1-
12
#468520000000
0!
0%
b10 *
0-
02
b10 6
#468530000000
1!
1%
1-
12
#468540000000
0!
0%
b11 *
0-
02
b11 6
#468550000000
1!
1%
1-
12
15
#468560000000
0!
0%
b100 *
0-
02
b100 6
#468570000000
1!
1%
1-
12
#468580000000
0!
0%
b101 *
0-
02
b101 6
#468590000000
1!
1%
1-
12
#468600000000
0!
0%
b110 *
0-
02
b110 6
#468610000000
1!
1%
1-
12
#468620000000
0!
0%
b111 *
0-
02
b111 6
#468630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#468640000000
0!
0%
b0 *
0-
02
b0 6
#468650000000
1!
1%
1-
12
#468660000000
0!
0%
b1 *
0-
02
b1 6
#468670000000
1!
1%
1-
12
#468680000000
0!
0%
b10 *
0-
02
b10 6
#468690000000
1!
1%
1-
12
#468700000000
0!
0%
b11 *
0-
02
b11 6
#468710000000
1!
1%
1-
12
15
#468720000000
0!
0%
b100 *
0-
02
b100 6
#468730000000
1!
1%
1-
12
#468740000000
0!
0%
b101 *
0-
02
b101 6
#468750000000
1!
1%
1-
12
#468760000000
0!
0%
b110 *
0-
02
b110 6
#468770000000
1!
1%
1-
12
#468780000000
0!
0%
b111 *
0-
02
b111 6
#468790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#468800000000
0!
0%
b0 *
0-
02
b0 6
#468810000000
1!
1%
1-
12
#468820000000
0!
0%
b1 *
0-
02
b1 6
#468830000000
1!
1%
1-
12
#468840000000
0!
0%
b10 *
0-
02
b10 6
#468850000000
1!
1%
1-
12
#468860000000
0!
0%
b11 *
0-
02
b11 6
#468870000000
1!
1%
1-
12
15
#468880000000
0!
0%
b100 *
0-
02
b100 6
#468890000000
1!
1%
1-
12
#468900000000
0!
0%
b101 *
0-
02
b101 6
#468910000000
1!
1%
1-
12
#468920000000
0!
0%
b110 *
0-
02
b110 6
#468930000000
1!
1%
1-
12
#468940000000
0!
0%
b111 *
0-
02
b111 6
#468950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#468960000000
0!
0%
b0 *
0-
02
b0 6
#468970000000
1!
1%
1-
12
#468980000000
0!
0%
b1 *
0-
02
b1 6
#468990000000
1!
1%
1-
12
#469000000000
0!
0%
b10 *
0-
02
b10 6
#469010000000
1!
1%
1-
12
#469020000000
0!
0%
b11 *
0-
02
b11 6
#469030000000
1!
1%
1-
12
15
#469040000000
0!
0%
b100 *
0-
02
b100 6
#469050000000
1!
1%
1-
12
#469060000000
0!
0%
b101 *
0-
02
b101 6
#469070000000
1!
1%
1-
12
#469080000000
0!
0%
b110 *
0-
02
b110 6
#469090000000
1!
1%
1-
12
#469100000000
0!
0%
b111 *
0-
02
b111 6
#469110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#469120000000
0!
0%
b0 *
0-
02
b0 6
#469130000000
1!
1%
1-
12
#469140000000
0!
0%
b1 *
0-
02
b1 6
#469150000000
1!
1%
1-
12
#469160000000
0!
0%
b10 *
0-
02
b10 6
#469170000000
1!
1%
1-
12
#469180000000
0!
0%
b11 *
0-
02
b11 6
#469190000000
1!
1%
1-
12
15
#469200000000
0!
0%
b100 *
0-
02
b100 6
#469210000000
1!
1%
1-
12
#469220000000
0!
0%
b101 *
0-
02
b101 6
#469230000000
1!
1%
1-
12
#469240000000
0!
0%
b110 *
0-
02
b110 6
#469250000000
1!
1%
1-
12
#469260000000
0!
0%
b111 *
0-
02
b111 6
#469270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#469280000000
0!
0%
b0 *
0-
02
b0 6
#469290000000
1!
1%
1-
12
#469300000000
0!
0%
b1 *
0-
02
b1 6
#469310000000
1!
1%
1-
12
#469320000000
0!
0%
b10 *
0-
02
b10 6
#469330000000
1!
1%
1-
12
#469340000000
0!
0%
b11 *
0-
02
b11 6
#469350000000
1!
1%
1-
12
15
#469360000000
0!
0%
b100 *
0-
02
b100 6
#469370000000
1!
1%
1-
12
#469380000000
0!
0%
b101 *
0-
02
b101 6
#469390000000
1!
1%
1-
12
#469400000000
0!
0%
b110 *
0-
02
b110 6
#469410000000
1!
1%
1-
12
#469420000000
0!
0%
b111 *
0-
02
b111 6
#469430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#469440000000
0!
0%
b0 *
0-
02
b0 6
#469450000000
1!
1%
1-
12
#469460000000
0!
0%
b1 *
0-
02
b1 6
#469470000000
1!
1%
1-
12
#469480000000
0!
0%
b10 *
0-
02
b10 6
#469490000000
1!
1%
1-
12
#469500000000
0!
0%
b11 *
0-
02
b11 6
#469510000000
1!
1%
1-
12
15
#469520000000
0!
0%
b100 *
0-
02
b100 6
#469530000000
1!
1%
1-
12
#469540000000
0!
0%
b101 *
0-
02
b101 6
#469550000000
1!
1%
1-
12
#469560000000
0!
0%
b110 *
0-
02
b110 6
#469570000000
1!
1%
1-
12
#469580000000
0!
0%
b111 *
0-
02
b111 6
#469590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#469600000000
0!
0%
b0 *
0-
02
b0 6
#469610000000
1!
1%
1-
12
#469620000000
0!
0%
b1 *
0-
02
b1 6
#469630000000
1!
1%
1-
12
#469640000000
0!
0%
b10 *
0-
02
b10 6
#469650000000
1!
1%
1-
12
#469660000000
0!
0%
b11 *
0-
02
b11 6
#469670000000
1!
1%
1-
12
15
#469680000000
0!
0%
b100 *
0-
02
b100 6
#469690000000
1!
1%
1-
12
#469700000000
0!
0%
b101 *
0-
02
b101 6
#469710000000
1!
1%
1-
12
#469720000000
0!
0%
b110 *
0-
02
b110 6
#469730000000
1!
1%
1-
12
#469740000000
0!
0%
b111 *
0-
02
b111 6
#469750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#469760000000
0!
0%
b0 *
0-
02
b0 6
#469770000000
1!
1%
1-
12
#469780000000
0!
0%
b1 *
0-
02
b1 6
#469790000000
1!
1%
1-
12
#469800000000
0!
0%
b10 *
0-
02
b10 6
#469810000000
1!
1%
1-
12
#469820000000
0!
0%
b11 *
0-
02
b11 6
#469830000000
1!
1%
1-
12
15
#469840000000
0!
0%
b100 *
0-
02
b100 6
#469850000000
1!
1%
1-
12
#469860000000
0!
0%
b101 *
0-
02
b101 6
#469870000000
1!
1%
1-
12
#469880000000
0!
0%
b110 *
0-
02
b110 6
#469890000000
1!
1%
1-
12
#469900000000
0!
0%
b111 *
0-
02
b111 6
#469910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#469920000000
0!
0%
b0 *
0-
02
b0 6
#469930000000
1!
1%
1-
12
#469940000000
0!
0%
b1 *
0-
02
b1 6
#469950000000
1!
1%
1-
12
#469960000000
0!
0%
b10 *
0-
02
b10 6
#469970000000
1!
1%
1-
12
#469980000000
0!
0%
b11 *
0-
02
b11 6
#469990000000
1!
1%
1-
12
15
#470000000000
0!
0%
b100 *
0-
02
b100 6
#470010000000
1!
1%
1-
12
#470020000000
0!
0%
b101 *
0-
02
b101 6
#470030000000
1!
1%
1-
12
#470040000000
0!
0%
b110 *
0-
02
b110 6
#470050000000
1!
1%
1-
12
#470060000000
0!
0%
b111 *
0-
02
b111 6
#470070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#470080000000
0!
0%
b0 *
0-
02
b0 6
#470090000000
1!
1%
1-
12
#470100000000
0!
0%
b1 *
0-
02
b1 6
#470110000000
1!
1%
1-
12
#470120000000
0!
0%
b10 *
0-
02
b10 6
#470130000000
1!
1%
1-
12
#470140000000
0!
0%
b11 *
0-
02
b11 6
#470150000000
1!
1%
1-
12
15
#470160000000
0!
0%
b100 *
0-
02
b100 6
#470170000000
1!
1%
1-
12
#470180000000
0!
0%
b101 *
0-
02
b101 6
#470190000000
1!
1%
1-
12
#470200000000
0!
0%
b110 *
0-
02
b110 6
#470210000000
1!
1%
1-
12
#470220000000
0!
0%
b111 *
0-
02
b111 6
#470230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#470240000000
0!
0%
b0 *
0-
02
b0 6
#470250000000
1!
1%
1-
12
#470260000000
0!
0%
b1 *
0-
02
b1 6
#470270000000
1!
1%
1-
12
#470280000000
0!
0%
b10 *
0-
02
b10 6
#470290000000
1!
1%
1-
12
#470300000000
0!
0%
b11 *
0-
02
b11 6
#470310000000
1!
1%
1-
12
15
#470320000000
0!
0%
b100 *
0-
02
b100 6
#470330000000
1!
1%
1-
12
#470340000000
0!
0%
b101 *
0-
02
b101 6
#470350000000
1!
1%
1-
12
#470360000000
0!
0%
b110 *
0-
02
b110 6
#470370000000
1!
1%
1-
12
#470380000000
0!
0%
b111 *
0-
02
b111 6
#470390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#470400000000
0!
0%
b0 *
0-
02
b0 6
#470410000000
1!
1%
1-
12
#470420000000
0!
0%
b1 *
0-
02
b1 6
#470430000000
1!
1%
1-
12
#470440000000
0!
0%
b10 *
0-
02
b10 6
#470450000000
1!
1%
1-
12
#470460000000
0!
0%
b11 *
0-
02
b11 6
#470470000000
1!
1%
1-
12
15
#470480000000
0!
0%
b100 *
0-
02
b100 6
#470490000000
1!
1%
1-
12
#470500000000
0!
0%
b101 *
0-
02
b101 6
#470510000000
1!
1%
1-
12
#470520000000
0!
0%
b110 *
0-
02
b110 6
#470530000000
1!
1%
1-
12
#470540000000
0!
0%
b111 *
0-
02
b111 6
#470550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#470560000000
0!
0%
b0 *
0-
02
b0 6
#470570000000
1!
1%
1-
12
#470580000000
0!
0%
b1 *
0-
02
b1 6
#470590000000
1!
1%
1-
12
#470600000000
0!
0%
b10 *
0-
02
b10 6
#470610000000
1!
1%
1-
12
#470620000000
0!
0%
b11 *
0-
02
b11 6
#470630000000
1!
1%
1-
12
15
#470640000000
0!
0%
b100 *
0-
02
b100 6
#470650000000
1!
1%
1-
12
#470660000000
0!
0%
b101 *
0-
02
b101 6
#470670000000
1!
1%
1-
12
#470680000000
0!
0%
b110 *
0-
02
b110 6
#470690000000
1!
1%
1-
12
#470700000000
0!
0%
b111 *
0-
02
b111 6
#470710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#470720000000
0!
0%
b0 *
0-
02
b0 6
#470730000000
1!
1%
1-
12
#470740000000
0!
0%
b1 *
0-
02
b1 6
#470750000000
1!
1%
1-
12
#470760000000
0!
0%
b10 *
0-
02
b10 6
#470770000000
1!
1%
1-
12
#470780000000
0!
0%
b11 *
0-
02
b11 6
#470790000000
1!
1%
1-
12
15
#470800000000
0!
0%
b100 *
0-
02
b100 6
#470810000000
1!
1%
1-
12
#470820000000
0!
0%
b101 *
0-
02
b101 6
#470830000000
1!
1%
1-
12
#470840000000
0!
0%
b110 *
0-
02
b110 6
#470850000000
1!
1%
1-
12
#470860000000
0!
0%
b111 *
0-
02
b111 6
#470870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#470880000000
0!
0%
b0 *
0-
02
b0 6
#470890000000
1!
1%
1-
12
#470900000000
0!
0%
b1 *
0-
02
b1 6
#470910000000
1!
1%
1-
12
#470920000000
0!
0%
b10 *
0-
02
b10 6
#470930000000
1!
1%
1-
12
#470940000000
0!
0%
b11 *
0-
02
b11 6
#470950000000
1!
1%
1-
12
15
#470960000000
0!
0%
b100 *
0-
02
b100 6
#470970000000
1!
1%
1-
12
#470980000000
0!
0%
b101 *
0-
02
b101 6
#470990000000
1!
1%
1-
12
#471000000000
0!
0%
b110 *
0-
02
b110 6
#471010000000
1!
1%
1-
12
#471020000000
0!
0%
b111 *
0-
02
b111 6
#471030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#471040000000
0!
0%
b0 *
0-
02
b0 6
#471050000000
1!
1%
1-
12
#471060000000
0!
0%
b1 *
0-
02
b1 6
#471070000000
1!
1%
1-
12
#471080000000
0!
0%
b10 *
0-
02
b10 6
#471090000000
1!
1%
1-
12
#471100000000
0!
0%
b11 *
0-
02
b11 6
#471110000000
1!
1%
1-
12
15
#471120000000
0!
0%
b100 *
0-
02
b100 6
#471130000000
1!
1%
1-
12
#471140000000
0!
0%
b101 *
0-
02
b101 6
#471150000000
1!
1%
1-
12
#471160000000
0!
0%
b110 *
0-
02
b110 6
#471170000000
1!
1%
1-
12
#471180000000
0!
0%
b111 *
0-
02
b111 6
#471190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#471200000000
0!
0%
b0 *
0-
02
b0 6
#471210000000
1!
1%
1-
12
#471220000000
0!
0%
b1 *
0-
02
b1 6
#471230000000
1!
1%
1-
12
#471240000000
0!
0%
b10 *
0-
02
b10 6
#471250000000
1!
1%
1-
12
#471260000000
0!
0%
b11 *
0-
02
b11 6
#471270000000
1!
1%
1-
12
15
#471280000000
0!
0%
b100 *
0-
02
b100 6
#471290000000
1!
1%
1-
12
#471300000000
0!
0%
b101 *
0-
02
b101 6
#471310000000
1!
1%
1-
12
#471320000000
0!
0%
b110 *
0-
02
b110 6
#471330000000
1!
1%
1-
12
#471340000000
0!
0%
b111 *
0-
02
b111 6
#471350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#471360000000
0!
0%
b0 *
0-
02
b0 6
#471370000000
1!
1%
1-
12
#471380000000
0!
0%
b1 *
0-
02
b1 6
#471390000000
1!
1%
1-
12
#471400000000
0!
0%
b10 *
0-
02
b10 6
#471410000000
1!
1%
1-
12
#471420000000
0!
0%
b11 *
0-
02
b11 6
#471430000000
1!
1%
1-
12
15
#471440000000
0!
0%
b100 *
0-
02
b100 6
#471450000000
1!
1%
1-
12
#471460000000
0!
0%
b101 *
0-
02
b101 6
#471470000000
1!
1%
1-
12
#471480000000
0!
0%
b110 *
0-
02
b110 6
#471490000000
1!
1%
1-
12
#471500000000
0!
0%
b111 *
0-
02
b111 6
#471510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#471520000000
0!
0%
b0 *
0-
02
b0 6
#471530000000
1!
1%
1-
12
#471540000000
0!
0%
b1 *
0-
02
b1 6
#471550000000
1!
1%
1-
12
#471560000000
0!
0%
b10 *
0-
02
b10 6
#471570000000
1!
1%
1-
12
#471580000000
0!
0%
b11 *
0-
02
b11 6
#471590000000
1!
1%
1-
12
15
#471600000000
0!
0%
b100 *
0-
02
b100 6
#471610000000
1!
1%
1-
12
#471620000000
0!
0%
b101 *
0-
02
b101 6
#471630000000
1!
1%
1-
12
#471640000000
0!
0%
b110 *
0-
02
b110 6
#471650000000
1!
1%
1-
12
#471660000000
0!
0%
b111 *
0-
02
b111 6
#471670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#471680000000
0!
0%
b0 *
0-
02
b0 6
#471690000000
1!
1%
1-
12
#471700000000
0!
0%
b1 *
0-
02
b1 6
#471710000000
1!
1%
1-
12
#471720000000
0!
0%
b10 *
0-
02
b10 6
#471730000000
1!
1%
1-
12
#471740000000
0!
0%
b11 *
0-
02
b11 6
#471750000000
1!
1%
1-
12
15
#471760000000
0!
0%
b100 *
0-
02
b100 6
#471770000000
1!
1%
1-
12
#471780000000
0!
0%
b101 *
0-
02
b101 6
#471790000000
1!
1%
1-
12
#471800000000
0!
0%
b110 *
0-
02
b110 6
#471810000000
1!
1%
1-
12
#471820000000
0!
0%
b111 *
0-
02
b111 6
#471830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#471840000000
0!
0%
b0 *
0-
02
b0 6
#471850000000
1!
1%
1-
12
#471860000000
0!
0%
b1 *
0-
02
b1 6
#471870000000
1!
1%
1-
12
#471880000000
0!
0%
b10 *
0-
02
b10 6
#471890000000
1!
1%
1-
12
#471900000000
0!
0%
b11 *
0-
02
b11 6
#471910000000
1!
1%
1-
12
15
#471920000000
0!
0%
b100 *
0-
02
b100 6
#471930000000
1!
1%
1-
12
#471940000000
0!
0%
b101 *
0-
02
b101 6
#471950000000
1!
1%
1-
12
#471960000000
0!
0%
b110 *
0-
02
b110 6
#471970000000
1!
1%
1-
12
#471980000000
0!
0%
b111 *
0-
02
b111 6
#471990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#472000000000
0!
0%
b0 *
0-
02
b0 6
#472010000000
1!
1%
1-
12
#472020000000
0!
0%
b1 *
0-
02
b1 6
#472030000000
1!
1%
1-
12
#472040000000
0!
0%
b10 *
0-
02
b10 6
#472050000000
1!
1%
1-
12
#472060000000
0!
0%
b11 *
0-
02
b11 6
#472070000000
1!
1%
1-
12
15
#472080000000
0!
0%
b100 *
0-
02
b100 6
#472090000000
1!
1%
1-
12
#472100000000
0!
0%
b101 *
0-
02
b101 6
#472110000000
1!
1%
1-
12
#472120000000
0!
0%
b110 *
0-
02
b110 6
#472130000000
1!
1%
1-
12
#472140000000
0!
0%
b111 *
0-
02
b111 6
#472150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#472160000000
0!
0%
b0 *
0-
02
b0 6
#472170000000
1!
1%
1-
12
#472180000000
0!
0%
b1 *
0-
02
b1 6
#472190000000
1!
1%
1-
12
#472200000000
0!
0%
b10 *
0-
02
b10 6
#472210000000
1!
1%
1-
12
#472220000000
0!
0%
b11 *
0-
02
b11 6
#472230000000
1!
1%
1-
12
15
#472240000000
0!
0%
b100 *
0-
02
b100 6
#472250000000
1!
1%
1-
12
#472260000000
0!
0%
b101 *
0-
02
b101 6
#472270000000
1!
1%
1-
12
#472280000000
0!
0%
b110 *
0-
02
b110 6
#472290000000
1!
1%
1-
12
#472300000000
0!
0%
b111 *
0-
02
b111 6
#472310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#472320000000
0!
0%
b0 *
0-
02
b0 6
#472330000000
1!
1%
1-
12
#472340000000
0!
0%
b1 *
0-
02
b1 6
#472350000000
1!
1%
1-
12
#472360000000
0!
0%
b10 *
0-
02
b10 6
#472370000000
1!
1%
1-
12
#472380000000
0!
0%
b11 *
0-
02
b11 6
#472390000000
1!
1%
1-
12
15
#472400000000
0!
0%
b100 *
0-
02
b100 6
#472410000000
1!
1%
1-
12
#472420000000
0!
0%
b101 *
0-
02
b101 6
#472430000000
1!
1%
1-
12
#472440000000
0!
0%
b110 *
0-
02
b110 6
#472450000000
1!
1%
1-
12
#472460000000
0!
0%
b111 *
0-
02
b111 6
#472470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#472480000000
0!
0%
b0 *
0-
02
b0 6
#472490000000
1!
1%
1-
12
#472500000000
0!
0%
b1 *
0-
02
b1 6
#472510000000
1!
1%
1-
12
#472520000000
0!
0%
b10 *
0-
02
b10 6
#472530000000
1!
1%
1-
12
#472540000000
0!
0%
b11 *
0-
02
b11 6
#472550000000
1!
1%
1-
12
15
#472560000000
0!
0%
b100 *
0-
02
b100 6
#472570000000
1!
1%
1-
12
#472580000000
0!
0%
b101 *
0-
02
b101 6
#472590000000
1!
1%
1-
12
#472600000000
0!
0%
b110 *
0-
02
b110 6
#472610000000
1!
1%
1-
12
#472620000000
0!
0%
b111 *
0-
02
b111 6
#472630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#472640000000
0!
0%
b0 *
0-
02
b0 6
#472650000000
1!
1%
1-
12
#472660000000
0!
0%
b1 *
0-
02
b1 6
#472670000000
1!
1%
1-
12
#472680000000
0!
0%
b10 *
0-
02
b10 6
#472690000000
1!
1%
1-
12
#472700000000
0!
0%
b11 *
0-
02
b11 6
#472710000000
1!
1%
1-
12
15
#472720000000
0!
0%
b100 *
0-
02
b100 6
#472730000000
1!
1%
1-
12
#472740000000
0!
0%
b101 *
0-
02
b101 6
#472750000000
1!
1%
1-
12
#472760000000
0!
0%
b110 *
0-
02
b110 6
#472770000000
1!
1%
1-
12
#472780000000
0!
0%
b111 *
0-
02
b111 6
#472790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#472800000000
0!
0%
b0 *
0-
02
b0 6
#472810000000
1!
1%
1-
12
#472820000000
0!
0%
b1 *
0-
02
b1 6
#472830000000
1!
1%
1-
12
#472840000000
0!
0%
b10 *
0-
02
b10 6
#472850000000
1!
1%
1-
12
#472860000000
0!
0%
b11 *
0-
02
b11 6
#472870000000
1!
1%
1-
12
15
#472880000000
0!
0%
b100 *
0-
02
b100 6
#472890000000
1!
1%
1-
12
#472900000000
0!
0%
b101 *
0-
02
b101 6
#472910000000
1!
1%
1-
12
#472920000000
0!
0%
b110 *
0-
02
b110 6
#472930000000
1!
1%
1-
12
#472940000000
0!
0%
b111 *
0-
02
b111 6
#472950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#472960000000
0!
0%
b0 *
0-
02
b0 6
#472970000000
1!
1%
1-
12
#472980000000
0!
0%
b1 *
0-
02
b1 6
#472990000000
1!
1%
1-
12
#473000000000
0!
0%
b10 *
0-
02
b10 6
#473010000000
1!
1%
1-
12
#473020000000
0!
0%
b11 *
0-
02
b11 6
#473030000000
1!
1%
1-
12
15
#473040000000
0!
0%
b100 *
0-
02
b100 6
#473050000000
1!
1%
1-
12
#473060000000
0!
0%
b101 *
0-
02
b101 6
#473070000000
1!
1%
1-
12
#473080000000
0!
0%
b110 *
0-
02
b110 6
#473090000000
1!
1%
1-
12
#473100000000
0!
0%
b111 *
0-
02
b111 6
#473110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#473120000000
0!
0%
b0 *
0-
02
b0 6
#473130000000
1!
1%
1-
12
#473140000000
0!
0%
b1 *
0-
02
b1 6
#473150000000
1!
1%
1-
12
#473160000000
0!
0%
b10 *
0-
02
b10 6
#473170000000
1!
1%
1-
12
#473180000000
0!
0%
b11 *
0-
02
b11 6
#473190000000
1!
1%
1-
12
15
#473200000000
0!
0%
b100 *
0-
02
b100 6
#473210000000
1!
1%
1-
12
#473220000000
0!
0%
b101 *
0-
02
b101 6
#473230000000
1!
1%
1-
12
#473240000000
0!
0%
b110 *
0-
02
b110 6
#473250000000
1!
1%
1-
12
#473260000000
0!
0%
b111 *
0-
02
b111 6
#473270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#473280000000
0!
0%
b0 *
0-
02
b0 6
#473290000000
1!
1%
1-
12
#473300000000
0!
0%
b1 *
0-
02
b1 6
#473310000000
1!
1%
1-
12
#473320000000
0!
0%
b10 *
0-
02
b10 6
#473330000000
1!
1%
1-
12
#473340000000
0!
0%
b11 *
0-
02
b11 6
#473350000000
1!
1%
1-
12
15
#473360000000
0!
0%
b100 *
0-
02
b100 6
#473370000000
1!
1%
1-
12
#473380000000
0!
0%
b101 *
0-
02
b101 6
#473390000000
1!
1%
1-
12
#473400000000
0!
0%
b110 *
0-
02
b110 6
#473410000000
1!
1%
1-
12
#473420000000
0!
0%
b111 *
0-
02
b111 6
#473430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#473440000000
0!
0%
b0 *
0-
02
b0 6
#473450000000
1!
1%
1-
12
#473460000000
0!
0%
b1 *
0-
02
b1 6
#473470000000
1!
1%
1-
12
#473480000000
0!
0%
b10 *
0-
02
b10 6
#473490000000
1!
1%
1-
12
#473500000000
0!
0%
b11 *
0-
02
b11 6
#473510000000
1!
1%
1-
12
15
#473520000000
0!
0%
b100 *
0-
02
b100 6
#473530000000
1!
1%
1-
12
#473540000000
0!
0%
b101 *
0-
02
b101 6
#473550000000
1!
1%
1-
12
#473560000000
0!
0%
b110 *
0-
02
b110 6
#473570000000
1!
1%
1-
12
#473580000000
0!
0%
b111 *
0-
02
b111 6
#473590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#473600000000
0!
0%
b0 *
0-
02
b0 6
#473610000000
1!
1%
1-
12
#473620000000
0!
0%
b1 *
0-
02
b1 6
#473630000000
1!
1%
1-
12
#473640000000
0!
0%
b10 *
0-
02
b10 6
#473650000000
1!
1%
1-
12
#473660000000
0!
0%
b11 *
0-
02
b11 6
#473670000000
1!
1%
1-
12
15
#473680000000
0!
0%
b100 *
0-
02
b100 6
#473690000000
1!
1%
1-
12
#473700000000
0!
0%
b101 *
0-
02
b101 6
#473710000000
1!
1%
1-
12
#473720000000
0!
0%
b110 *
0-
02
b110 6
#473730000000
1!
1%
1-
12
#473740000000
0!
0%
b111 *
0-
02
b111 6
#473750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#473760000000
0!
0%
b0 *
0-
02
b0 6
#473770000000
1!
1%
1-
12
#473780000000
0!
0%
b1 *
0-
02
b1 6
#473790000000
1!
1%
1-
12
#473800000000
0!
0%
b10 *
0-
02
b10 6
#473810000000
1!
1%
1-
12
#473820000000
0!
0%
b11 *
0-
02
b11 6
#473830000000
1!
1%
1-
12
15
#473840000000
0!
0%
b100 *
0-
02
b100 6
#473850000000
1!
1%
1-
12
#473860000000
0!
0%
b101 *
0-
02
b101 6
#473870000000
1!
1%
1-
12
#473880000000
0!
0%
b110 *
0-
02
b110 6
#473890000000
1!
1%
1-
12
#473900000000
0!
0%
b111 *
0-
02
b111 6
#473910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#473920000000
0!
0%
b0 *
0-
02
b0 6
#473930000000
1!
1%
1-
12
#473940000000
0!
0%
b1 *
0-
02
b1 6
#473950000000
1!
1%
1-
12
#473960000000
0!
0%
b10 *
0-
02
b10 6
#473970000000
1!
1%
1-
12
#473980000000
0!
0%
b11 *
0-
02
b11 6
#473990000000
1!
1%
1-
12
15
#474000000000
0!
0%
b100 *
0-
02
b100 6
#474010000000
1!
1%
1-
12
#474020000000
0!
0%
b101 *
0-
02
b101 6
#474030000000
1!
1%
1-
12
#474040000000
0!
0%
b110 *
0-
02
b110 6
#474050000000
1!
1%
1-
12
#474060000000
0!
0%
b111 *
0-
02
b111 6
#474070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#474080000000
0!
0%
b0 *
0-
02
b0 6
#474090000000
1!
1%
1-
12
#474100000000
0!
0%
b1 *
0-
02
b1 6
#474110000000
1!
1%
1-
12
#474120000000
0!
0%
b10 *
0-
02
b10 6
#474130000000
1!
1%
1-
12
#474140000000
0!
0%
b11 *
0-
02
b11 6
#474150000000
1!
1%
1-
12
15
#474160000000
0!
0%
b100 *
0-
02
b100 6
#474170000000
1!
1%
1-
12
#474180000000
0!
0%
b101 *
0-
02
b101 6
#474190000000
1!
1%
1-
12
#474200000000
0!
0%
b110 *
0-
02
b110 6
#474210000000
1!
1%
1-
12
#474220000000
0!
0%
b111 *
0-
02
b111 6
#474230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#474240000000
0!
0%
b0 *
0-
02
b0 6
#474250000000
1!
1%
1-
12
#474260000000
0!
0%
b1 *
0-
02
b1 6
#474270000000
1!
1%
1-
12
#474280000000
0!
0%
b10 *
0-
02
b10 6
#474290000000
1!
1%
1-
12
#474300000000
0!
0%
b11 *
0-
02
b11 6
#474310000000
1!
1%
1-
12
15
#474320000000
0!
0%
b100 *
0-
02
b100 6
#474330000000
1!
1%
1-
12
#474340000000
0!
0%
b101 *
0-
02
b101 6
#474350000000
1!
1%
1-
12
#474360000000
0!
0%
b110 *
0-
02
b110 6
#474370000000
1!
1%
1-
12
#474380000000
0!
0%
b111 *
0-
02
b111 6
#474390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#474400000000
0!
0%
b0 *
0-
02
b0 6
#474410000000
1!
1%
1-
12
#474420000000
0!
0%
b1 *
0-
02
b1 6
#474430000000
1!
1%
1-
12
#474440000000
0!
0%
b10 *
0-
02
b10 6
#474450000000
1!
1%
1-
12
#474460000000
0!
0%
b11 *
0-
02
b11 6
#474470000000
1!
1%
1-
12
15
#474480000000
0!
0%
b100 *
0-
02
b100 6
#474490000000
1!
1%
1-
12
#474500000000
0!
0%
b101 *
0-
02
b101 6
#474510000000
1!
1%
1-
12
#474520000000
0!
0%
b110 *
0-
02
b110 6
#474530000000
1!
1%
1-
12
#474540000000
0!
0%
b111 *
0-
02
b111 6
#474550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#474560000000
0!
0%
b0 *
0-
02
b0 6
#474570000000
1!
1%
1-
12
#474580000000
0!
0%
b1 *
0-
02
b1 6
#474590000000
1!
1%
1-
12
#474600000000
0!
0%
b10 *
0-
02
b10 6
#474610000000
1!
1%
1-
12
#474620000000
0!
0%
b11 *
0-
02
b11 6
#474630000000
1!
1%
1-
12
15
#474640000000
0!
0%
b100 *
0-
02
b100 6
#474650000000
1!
1%
1-
12
#474660000000
0!
0%
b101 *
0-
02
b101 6
#474670000000
1!
1%
1-
12
#474680000000
0!
0%
b110 *
0-
02
b110 6
#474690000000
1!
1%
1-
12
#474700000000
0!
0%
b111 *
0-
02
b111 6
#474710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#474720000000
0!
0%
b0 *
0-
02
b0 6
#474730000000
1!
1%
1-
12
#474740000000
0!
0%
b1 *
0-
02
b1 6
#474750000000
1!
1%
1-
12
#474760000000
0!
0%
b10 *
0-
02
b10 6
#474770000000
1!
1%
1-
12
#474780000000
0!
0%
b11 *
0-
02
b11 6
#474790000000
1!
1%
1-
12
15
#474800000000
0!
0%
b100 *
0-
02
b100 6
#474810000000
1!
1%
1-
12
#474820000000
0!
0%
b101 *
0-
02
b101 6
#474830000000
1!
1%
1-
12
#474840000000
0!
0%
b110 *
0-
02
b110 6
#474850000000
1!
1%
1-
12
#474860000000
0!
0%
b111 *
0-
02
b111 6
#474870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#474880000000
0!
0%
b0 *
0-
02
b0 6
#474890000000
1!
1%
1-
12
#474900000000
0!
0%
b1 *
0-
02
b1 6
#474910000000
1!
1%
1-
12
#474920000000
0!
0%
b10 *
0-
02
b10 6
#474930000000
1!
1%
1-
12
#474940000000
0!
0%
b11 *
0-
02
b11 6
#474950000000
1!
1%
1-
12
15
#474960000000
0!
0%
b100 *
0-
02
b100 6
#474970000000
1!
1%
1-
12
#474980000000
0!
0%
b101 *
0-
02
b101 6
#474990000000
1!
1%
1-
12
#475000000000
0!
0%
b110 *
0-
02
b110 6
#475010000000
1!
1%
1-
12
#475020000000
0!
0%
b111 *
0-
02
b111 6
#475030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#475040000000
0!
0%
b0 *
0-
02
b0 6
#475050000000
1!
1%
1-
12
#475060000000
0!
0%
b1 *
0-
02
b1 6
#475070000000
1!
1%
1-
12
#475080000000
0!
0%
b10 *
0-
02
b10 6
#475090000000
1!
1%
1-
12
#475100000000
0!
0%
b11 *
0-
02
b11 6
#475110000000
1!
1%
1-
12
15
#475120000000
0!
0%
b100 *
0-
02
b100 6
#475130000000
1!
1%
1-
12
#475140000000
0!
0%
b101 *
0-
02
b101 6
#475150000000
1!
1%
1-
12
#475160000000
0!
0%
b110 *
0-
02
b110 6
#475170000000
1!
1%
1-
12
#475180000000
0!
0%
b111 *
0-
02
b111 6
#475190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#475200000000
0!
0%
b0 *
0-
02
b0 6
#475210000000
1!
1%
1-
12
#475220000000
0!
0%
b1 *
0-
02
b1 6
#475230000000
1!
1%
1-
12
#475240000000
0!
0%
b10 *
0-
02
b10 6
#475250000000
1!
1%
1-
12
#475260000000
0!
0%
b11 *
0-
02
b11 6
#475270000000
1!
1%
1-
12
15
#475280000000
0!
0%
b100 *
0-
02
b100 6
#475290000000
1!
1%
1-
12
#475300000000
0!
0%
b101 *
0-
02
b101 6
#475310000000
1!
1%
1-
12
#475320000000
0!
0%
b110 *
0-
02
b110 6
#475330000000
1!
1%
1-
12
#475340000000
0!
0%
b111 *
0-
02
b111 6
#475350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#475360000000
0!
0%
b0 *
0-
02
b0 6
#475370000000
1!
1%
1-
12
#475380000000
0!
0%
b1 *
0-
02
b1 6
#475390000000
1!
1%
1-
12
#475400000000
0!
0%
b10 *
0-
02
b10 6
#475410000000
1!
1%
1-
12
#475420000000
0!
0%
b11 *
0-
02
b11 6
#475430000000
1!
1%
1-
12
15
#475440000000
0!
0%
b100 *
0-
02
b100 6
#475450000000
1!
1%
1-
12
#475460000000
0!
0%
b101 *
0-
02
b101 6
#475470000000
1!
1%
1-
12
#475480000000
0!
0%
b110 *
0-
02
b110 6
#475490000000
1!
1%
1-
12
#475500000000
0!
0%
b111 *
0-
02
b111 6
#475510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#475520000000
0!
0%
b0 *
0-
02
b0 6
#475530000000
1!
1%
1-
12
#475540000000
0!
0%
b1 *
0-
02
b1 6
#475550000000
1!
1%
1-
12
#475560000000
0!
0%
b10 *
0-
02
b10 6
#475570000000
1!
1%
1-
12
#475580000000
0!
0%
b11 *
0-
02
b11 6
#475590000000
1!
1%
1-
12
15
#475600000000
0!
0%
b100 *
0-
02
b100 6
#475610000000
1!
1%
1-
12
#475620000000
0!
0%
b101 *
0-
02
b101 6
#475630000000
1!
1%
1-
12
#475640000000
0!
0%
b110 *
0-
02
b110 6
#475650000000
1!
1%
1-
12
#475660000000
0!
0%
b111 *
0-
02
b111 6
#475670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#475680000000
0!
0%
b0 *
0-
02
b0 6
#475690000000
1!
1%
1-
12
#475700000000
0!
0%
b1 *
0-
02
b1 6
#475710000000
1!
1%
1-
12
#475720000000
0!
0%
b10 *
0-
02
b10 6
#475730000000
1!
1%
1-
12
#475740000000
0!
0%
b11 *
0-
02
b11 6
#475750000000
1!
1%
1-
12
15
#475760000000
0!
0%
b100 *
0-
02
b100 6
#475770000000
1!
1%
1-
12
#475780000000
0!
0%
b101 *
0-
02
b101 6
#475790000000
1!
1%
1-
12
#475800000000
0!
0%
b110 *
0-
02
b110 6
#475810000000
1!
1%
1-
12
#475820000000
0!
0%
b111 *
0-
02
b111 6
#475830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#475840000000
0!
0%
b0 *
0-
02
b0 6
#475850000000
1!
1%
1-
12
#475860000000
0!
0%
b1 *
0-
02
b1 6
#475870000000
1!
1%
1-
12
#475880000000
0!
0%
b10 *
0-
02
b10 6
#475890000000
1!
1%
1-
12
#475900000000
0!
0%
b11 *
0-
02
b11 6
#475910000000
1!
1%
1-
12
15
#475920000000
0!
0%
b100 *
0-
02
b100 6
#475930000000
1!
1%
1-
12
#475940000000
0!
0%
b101 *
0-
02
b101 6
#475950000000
1!
1%
1-
12
#475960000000
0!
0%
b110 *
0-
02
b110 6
#475970000000
1!
1%
1-
12
#475980000000
0!
0%
b111 *
0-
02
b111 6
#475990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#476000000000
0!
0%
b0 *
0-
02
b0 6
#476010000000
1!
1%
1-
12
#476020000000
0!
0%
b1 *
0-
02
b1 6
#476030000000
1!
1%
1-
12
#476040000000
0!
0%
b10 *
0-
02
b10 6
#476050000000
1!
1%
1-
12
#476060000000
0!
0%
b11 *
0-
02
b11 6
#476070000000
1!
1%
1-
12
15
#476080000000
0!
0%
b100 *
0-
02
b100 6
#476090000000
1!
1%
1-
12
#476100000000
0!
0%
b101 *
0-
02
b101 6
#476110000000
1!
1%
1-
12
#476120000000
0!
0%
b110 *
0-
02
b110 6
#476130000000
1!
1%
1-
12
#476140000000
0!
0%
b111 *
0-
02
b111 6
#476150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#476160000000
0!
0%
b0 *
0-
02
b0 6
#476170000000
1!
1%
1-
12
#476180000000
0!
0%
b1 *
0-
02
b1 6
#476190000000
1!
1%
1-
12
#476200000000
0!
0%
b10 *
0-
02
b10 6
#476210000000
1!
1%
1-
12
#476220000000
0!
0%
b11 *
0-
02
b11 6
#476230000000
1!
1%
1-
12
15
#476240000000
0!
0%
b100 *
0-
02
b100 6
#476250000000
1!
1%
1-
12
#476260000000
0!
0%
b101 *
0-
02
b101 6
#476270000000
1!
1%
1-
12
#476280000000
0!
0%
b110 *
0-
02
b110 6
#476290000000
1!
1%
1-
12
#476300000000
0!
0%
b111 *
0-
02
b111 6
#476310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#476320000000
0!
0%
b0 *
0-
02
b0 6
#476330000000
1!
1%
1-
12
#476340000000
0!
0%
b1 *
0-
02
b1 6
#476350000000
1!
1%
1-
12
#476360000000
0!
0%
b10 *
0-
02
b10 6
#476370000000
1!
1%
1-
12
#476380000000
0!
0%
b11 *
0-
02
b11 6
#476390000000
1!
1%
1-
12
15
#476400000000
0!
0%
b100 *
0-
02
b100 6
#476410000000
1!
1%
1-
12
#476420000000
0!
0%
b101 *
0-
02
b101 6
#476430000000
1!
1%
1-
12
#476440000000
0!
0%
b110 *
0-
02
b110 6
#476450000000
1!
1%
1-
12
#476460000000
0!
0%
b111 *
0-
02
b111 6
#476470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#476480000000
0!
0%
b0 *
0-
02
b0 6
#476490000000
1!
1%
1-
12
#476500000000
0!
0%
b1 *
0-
02
b1 6
#476510000000
1!
1%
1-
12
#476520000000
0!
0%
b10 *
0-
02
b10 6
#476530000000
1!
1%
1-
12
#476540000000
0!
0%
b11 *
0-
02
b11 6
#476550000000
1!
1%
1-
12
15
#476560000000
0!
0%
b100 *
0-
02
b100 6
#476570000000
1!
1%
1-
12
#476580000000
0!
0%
b101 *
0-
02
b101 6
#476590000000
1!
1%
1-
12
#476600000000
0!
0%
b110 *
0-
02
b110 6
#476610000000
1!
1%
1-
12
#476620000000
0!
0%
b111 *
0-
02
b111 6
#476630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#476640000000
0!
0%
b0 *
0-
02
b0 6
#476650000000
1!
1%
1-
12
#476660000000
0!
0%
b1 *
0-
02
b1 6
#476670000000
1!
1%
1-
12
#476680000000
0!
0%
b10 *
0-
02
b10 6
#476690000000
1!
1%
1-
12
#476700000000
0!
0%
b11 *
0-
02
b11 6
#476710000000
1!
1%
1-
12
15
#476720000000
0!
0%
b100 *
0-
02
b100 6
#476730000000
1!
1%
1-
12
#476740000000
0!
0%
b101 *
0-
02
b101 6
#476750000000
1!
1%
1-
12
#476760000000
0!
0%
b110 *
0-
02
b110 6
#476770000000
1!
1%
1-
12
#476780000000
0!
0%
b111 *
0-
02
b111 6
#476790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#476800000000
0!
0%
b0 *
0-
02
b0 6
#476810000000
1!
1%
1-
12
#476820000000
0!
0%
b1 *
0-
02
b1 6
#476830000000
1!
1%
1-
12
#476840000000
0!
0%
b10 *
0-
02
b10 6
#476850000000
1!
1%
1-
12
#476860000000
0!
0%
b11 *
0-
02
b11 6
#476870000000
1!
1%
1-
12
15
#476880000000
0!
0%
b100 *
0-
02
b100 6
#476890000000
1!
1%
1-
12
#476900000000
0!
0%
b101 *
0-
02
b101 6
#476910000000
1!
1%
1-
12
#476920000000
0!
0%
b110 *
0-
02
b110 6
#476930000000
1!
1%
1-
12
#476940000000
0!
0%
b111 *
0-
02
b111 6
#476950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#476960000000
0!
0%
b0 *
0-
02
b0 6
#476970000000
1!
1%
1-
12
#476980000000
0!
0%
b1 *
0-
02
b1 6
#476990000000
1!
1%
1-
12
#477000000000
0!
0%
b10 *
0-
02
b10 6
#477010000000
1!
1%
1-
12
#477020000000
0!
0%
b11 *
0-
02
b11 6
#477030000000
1!
1%
1-
12
15
#477040000000
0!
0%
b100 *
0-
02
b100 6
#477050000000
1!
1%
1-
12
#477060000000
0!
0%
b101 *
0-
02
b101 6
#477070000000
1!
1%
1-
12
#477080000000
0!
0%
b110 *
0-
02
b110 6
#477090000000
1!
1%
1-
12
#477100000000
0!
0%
b111 *
0-
02
b111 6
#477110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#477120000000
0!
0%
b0 *
0-
02
b0 6
#477130000000
1!
1%
1-
12
#477140000000
0!
0%
b1 *
0-
02
b1 6
#477150000000
1!
1%
1-
12
#477160000000
0!
0%
b10 *
0-
02
b10 6
#477170000000
1!
1%
1-
12
#477180000000
0!
0%
b11 *
0-
02
b11 6
#477190000000
1!
1%
1-
12
15
#477200000000
0!
0%
b100 *
0-
02
b100 6
#477210000000
1!
1%
1-
12
#477220000000
0!
0%
b101 *
0-
02
b101 6
#477230000000
1!
1%
1-
12
#477240000000
0!
0%
b110 *
0-
02
b110 6
#477250000000
1!
1%
1-
12
#477260000000
0!
0%
b111 *
0-
02
b111 6
#477270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#477280000000
0!
0%
b0 *
0-
02
b0 6
#477290000000
1!
1%
1-
12
#477300000000
0!
0%
b1 *
0-
02
b1 6
#477310000000
1!
1%
1-
12
#477320000000
0!
0%
b10 *
0-
02
b10 6
#477330000000
1!
1%
1-
12
#477340000000
0!
0%
b11 *
0-
02
b11 6
#477350000000
1!
1%
1-
12
15
#477360000000
0!
0%
b100 *
0-
02
b100 6
#477370000000
1!
1%
1-
12
#477380000000
0!
0%
b101 *
0-
02
b101 6
#477390000000
1!
1%
1-
12
#477400000000
0!
0%
b110 *
0-
02
b110 6
#477410000000
1!
1%
1-
12
#477420000000
0!
0%
b111 *
0-
02
b111 6
#477430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#477440000000
0!
0%
b0 *
0-
02
b0 6
#477450000000
1!
1%
1-
12
#477460000000
0!
0%
b1 *
0-
02
b1 6
#477470000000
1!
1%
1-
12
#477480000000
0!
0%
b10 *
0-
02
b10 6
#477490000000
1!
1%
1-
12
#477500000000
0!
0%
b11 *
0-
02
b11 6
#477510000000
1!
1%
1-
12
15
#477520000000
0!
0%
b100 *
0-
02
b100 6
#477530000000
1!
1%
1-
12
#477540000000
0!
0%
b101 *
0-
02
b101 6
#477550000000
1!
1%
1-
12
#477560000000
0!
0%
b110 *
0-
02
b110 6
#477570000000
1!
1%
1-
12
#477580000000
0!
0%
b111 *
0-
02
b111 6
#477590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#477600000000
0!
0%
b0 *
0-
02
b0 6
#477610000000
1!
1%
1-
12
#477620000000
0!
0%
b1 *
0-
02
b1 6
#477630000000
1!
1%
1-
12
#477640000000
0!
0%
b10 *
0-
02
b10 6
#477650000000
1!
1%
1-
12
#477660000000
0!
0%
b11 *
0-
02
b11 6
#477670000000
1!
1%
1-
12
15
#477680000000
0!
0%
b100 *
0-
02
b100 6
#477690000000
1!
1%
1-
12
#477700000000
0!
0%
b101 *
0-
02
b101 6
#477710000000
1!
1%
1-
12
#477720000000
0!
0%
b110 *
0-
02
b110 6
#477730000000
1!
1%
1-
12
#477740000000
0!
0%
b111 *
0-
02
b111 6
#477750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#477760000000
0!
0%
b0 *
0-
02
b0 6
#477770000000
1!
1%
1-
12
#477780000000
0!
0%
b1 *
0-
02
b1 6
#477790000000
1!
1%
1-
12
#477800000000
0!
0%
b10 *
0-
02
b10 6
#477810000000
1!
1%
1-
12
#477820000000
0!
0%
b11 *
0-
02
b11 6
#477830000000
1!
1%
1-
12
15
#477840000000
0!
0%
b100 *
0-
02
b100 6
#477850000000
1!
1%
1-
12
#477860000000
0!
0%
b101 *
0-
02
b101 6
#477870000000
1!
1%
1-
12
#477880000000
0!
0%
b110 *
0-
02
b110 6
#477890000000
1!
1%
1-
12
#477900000000
0!
0%
b111 *
0-
02
b111 6
#477910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#477920000000
0!
0%
b0 *
0-
02
b0 6
#477930000000
1!
1%
1-
12
#477940000000
0!
0%
b1 *
0-
02
b1 6
#477950000000
1!
1%
1-
12
#477960000000
0!
0%
b10 *
0-
02
b10 6
#477970000000
1!
1%
1-
12
#477980000000
0!
0%
b11 *
0-
02
b11 6
#477990000000
1!
1%
1-
12
15
#478000000000
0!
0%
b100 *
0-
02
b100 6
#478010000000
1!
1%
1-
12
#478020000000
0!
0%
b101 *
0-
02
b101 6
#478030000000
1!
1%
1-
12
#478040000000
0!
0%
b110 *
0-
02
b110 6
#478050000000
1!
1%
1-
12
#478060000000
0!
0%
b111 *
0-
02
b111 6
#478070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#478080000000
0!
0%
b0 *
0-
02
b0 6
#478090000000
1!
1%
1-
12
#478100000000
0!
0%
b1 *
0-
02
b1 6
#478110000000
1!
1%
1-
12
#478120000000
0!
0%
b10 *
0-
02
b10 6
#478130000000
1!
1%
1-
12
#478140000000
0!
0%
b11 *
0-
02
b11 6
#478150000000
1!
1%
1-
12
15
#478160000000
0!
0%
b100 *
0-
02
b100 6
#478170000000
1!
1%
1-
12
#478180000000
0!
0%
b101 *
0-
02
b101 6
#478190000000
1!
1%
1-
12
#478200000000
0!
0%
b110 *
0-
02
b110 6
#478210000000
1!
1%
1-
12
#478220000000
0!
0%
b111 *
0-
02
b111 6
#478230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#478240000000
0!
0%
b0 *
0-
02
b0 6
#478250000000
1!
1%
1-
12
#478260000000
0!
0%
b1 *
0-
02
b1 6
#478270000000
1!
1%
1-
12
#478280000000
0!
0%
b10 *
0-
02
b10 6
#478290000000
1!
1%
1-
12
#478300000000
0!
0%
b11 *
0-
02
b11 6
#478310000000
1!
1%
1-
12
15
#478320000000
0!
0%
b100 *
0-
02
b100 6
#478330000000
1!
1%
1-
12
#478340000000
0!
0%
b101 *
0-
02
b101 6
#478350000000
1!
1%
1-
12
#478360000000
0!
0%
b110 *
0-
02
b110 6
#478370000000
1!
1%
1-
12
#478380000000
0!
0%
b111 *
0-
02
b111 6
#478390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#478400000000
0!
0%
b0 *
0-
02
b0 6
#478410000000
1!
1%
1-
12
#478420000000
0!
0%
b1 *
0-
02
b1 6
#478430000000
1!
1%
1-
12
#478440000000
0!
0%
b10 *
0-
02
b10 6
#478450000000
1!
1%
1-
12
#478460000000
0!
0%
b11 *
0-
02
b11 6
#478470000000
1!
1%
1-
12
15
#478480000000
0!
0%
b100 *
0-
02
b100 6
#478490000000
1!
1%
1-
12
#478500000000
0!
0%
b101 *
0-
02
b101 6
#478510000000
1!
1%
1-
12
#478520000000
0!
0%
b110 *
0-
02
b110 6
#478530000000
1!
1%
1-
12
#478540000000
0!
0%
b111 *
0-
02
b111 6
#478550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#478560000000
0!
0%
b0 *
0-
02
b0 6
#478570000000
1!
1%
1-
12
#478580000000
0!
0%
b1 *
0-
02
b1 6
#478590000000
1!
1%
1-
12
#478600000000
0!
0%
b10 *
0-
02
b10 6
#478610000000
1!
1%
1-
12
#478620000000
0!
0%
b11 *
0-
02
b11 6
#478630000000
1!
1%
1-
12
15
#478640000000
0!
0%
b100 *
0-
02
b100 6
#478650000000
1!
1%
1-
12
#478660000000
0!
0%
b101 *
0-
02
b101 6
#478670000000
1!
1%
1-
12
#478680000000
0!
0%
b110 *
0-
02
b110 6
#478690000000
1!
1%
1-
12
#478700000000
0!
0%
b111 *
0-
02
b111 6
#478710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#478720000000
0!
0%
b0 *
0-
02
b0 6
#478730000000
1!
1%
1-
12
#478740000000
0!
0%
b1 *
0-
02
b1 6
#478750000000
1!
1%
1-
12
#478760000000
0!
0%
b10 *
0-
02
b10 6
#478770000000
1!
1%
1-
12
#478780000000
0!
0%
b11 *
0-
02
b11 6
#478790000000
1!
1%
1-
12
15
#478800000000
0!
0%
b100 *
0-
02
b100 6
#478810000000
1!
1%
1-
12
#478820000000
0!
0%
b101 *
0-
02
b101 6
#478830000000
1!
1%
1-
12
#478840000000
0!
0%
b110 *
0-
02
b110 6
#478850000000
1!
1%
1-
12
#478860000000
0!
0%
b111 *
0-
02
b111 6
#478870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#478880000000
0!
0%
b0 *
0-
02
b0 6
#478890000000
1!
1%
1-
12
#478900000000
0!
0%
b1 *
0-
02
b1 6
#478910000000
1!
1%
1-
12
#478920000000
0!
0%
b10 *
0-
02
b10 6
#478930000000
1!
1%
1-
12
#478940000000
0!
0%
b11 *
0-
02
b11 6
#478950000000
1!
1%
1-
12
15
#478960000000
0!
0%
b100 *
0-
02
b100 6
#478970000000
1!
1%
1-
12
#478980000000
0!
0%
b101 *
0-
02
b101 6
#478990000000
1!
1%
1-
12
#479000000000
0!
0%
b110 *
0-
02
b110 6
#479010000000
1!
1%
1-
12
#479020000000
0!
0%
b111 *
0-
02
b111 6
#479030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#479040000000
0!
0%
b0 *
0-
02
b0 6
#479050000000
1!
1%
1-
12
#479060000000
0!
0%
b1 *
0-
02
b1 6
#479070000000
1!
1%
1-
12
#479080000000
0!
0%
b10 *
0-
02
b10 6
#479090000000
1!
1%
1-
12
#479100000000
0!
0%
b11 *
0-
02
b11 6
#479110000000
1!
1%
1-
12
15
#479120000000
0!
0%
b100 *
0-
02
b100 6
#479130000000
1!
1%
1-
12
#479140000000
0!
0%
b101 *
0-
02
b101 6
#479150000000
1!
1%
1-
12
#479160000000
0!
0%
b110 *
0-
02
b110 6
#479170000000
1!
1%
1-
12
#479180000000
0!
0%
b111 *
0-
02
b111 6
#479190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#479200000000
0!
0%
b0 *
0-
02
b0 6
#479210000000
1!
1%
1-
12
#479220000000
0!
0%
b1 *
0-
02
b1 6
#479230000000
1!
1%
1-
12
#479240000000
0!
0%
b10 *
0-
02
b10 6
#479250000000
1!
1%
1-
12
#479260000000
0!
0%
b11 *
0-
02
b11 6
#479270000000
1!
1%
1-
12
15
#479280000000
0!
0%
b100 *
0-
02
b100 6
#479290000000
1!
1%
1-
12
#479300000000
0!
0%
b101 *
0-
02
b101 6
#479310000000
1!
1%
1-
12
#479320000000
0!
0%
b110 *
0-
02
b110 6
#479330000000
1!
1%
1-
12
#479340000000
0!
0%
b111 *
0-
02
b111 6
#479350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#479360000000
0!
0%
b0 *
0-
02
b0 6
#479370000000
1!
1%
1-
12
#479380000000
0!
0%
b1 *
0-
02
b1 6
#479390000000
1!
1%
1-
12
#479400000000
0!
0%
b10 *
0-
02
b10 6
#479410000000
1!
1%
1-
12
#479420000000
0!
0%
b11 *
0-
02
b11 6
#479430000000
1!
1%
1-
12
15
#479440000000
0!
0%
b100 *
0-
02
b100 6
#479450000000
1!
1%
1-
12
#479460000000
0!
0%
b101 *
0-
02
b101 6
#479470000000
1!
1%
1-
12
#479480000000
0!
0%
b110 *
0-
02
b110 6
#479490000000
1!
1%
1-
12
#479500000000
0!
0%
b111 *
0-
02
b111 6
#479510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#479520000000
0!
0%
b0 *
0-
02
b0 6
#479530000000
1!
1%
1-
12
#479540000000
0!
0%
b1 *
0-
02
b1 6
#479550000000
1!
1%
1-
12
#479560000000
0!
0%
b10 *
0-
02
b10 6
#479570000000
1!
1%
1-
12
#479580000000
0!
0%
b11 *
0-
02
b11 6
#479590000000
1!
1%
1-
12
15
#479600000000
0!
0%
b100 *
0-
02
b100 6
#479610000000
1!
1%
1-
12
#479620000000
0!
0%
b101 *
0-
02
b101 6
#479630000000
1!
1%
1-
12
#479640000000
0!
0%
b110 *
0-
02
b110 6
#479650000000
1!
1%
1-
12
#479660000000
0!
0%
b111 *
0-
02
b111 6
#479670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#479680000000
0!
0%
b0 *
0-
02
b0 6
#479690000000
1!
1%
1-
12
#479700000000
0!
0%
b1 *
0-
02
b1 6
#479710000000
1!
1%
1-
12
#479720000000
0!
0%
b10 *
0-
02
b10 6
#479730000000
1!
1%
1-
12
#479740000000
0!
0%
b11 *
0-
02
b11 6
#479750000000
1!
1%
1-
12
15
#479760000000
0!
0%
b100 *
0-
02
b100 6
#479770000000
1!
1%
1-
12
#479780000000
0!
0%
b101 *
0-
02
b101 6
#479790000000
1!
1%
1-
12
#479800000000
0!
0%
b110 *
0-
02
b110 6
#479810000000
1!
1%
1-
12
#479820000000
0!
0%
b111 *
0-
02
b111 6
#479830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#479840000000
0!
0%
b0 *
0-
02
b0 6
#479850000000
1!
1%
1-
12
#479860000000
0!
0%
b1 *
0-
02
b1 6
#479870000000
1!
1%
1-
12
#479880000000
0!
0%
b10 *
0-
02
b10 6
#479890000000
1!
1%
1-
12
#479900000000
0!
0%
b11 *
0-
02
b11 6
#479910000000
1!
1%
1-
12
15
#479920000000
0!
0%
b100 *
0-
02
b100 6
#479930000000
1!
1%
1-
12
#479940000000
0!
0%
b101 *
0-
02
b101 6
#479950000000
1!
1%
1-
12
#479960000000
0!
0%
b110 *
0-
02
b110 6
#479970000000
1!
1%
1-
12
#479980000000
0!
0%
b111 *
0-
02
b111 6
#479990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#480000000000
0!
0%
b0 *
0-
02
b0 6
#480010000000
1!
1%
1-
12
#480020000000
0!
0%
b1 *
0-
02
b1 6
#480030000000
1!
1%
1-
12
#480040000000
0!
0%
b10 *
0-
02
b10 6
#480050000000
1!
1%
1-
12
#480060000000
0!
0%
b11 *
0-
02
b11 6
#480070000000
1!
1%
1-
12
15
#480080000000
0!
0%
b100 *
0-
02
b100 6
#480090000000
1!
1%
1-
12
#480100000000
0!
0%
b101 *
0-
02
b101 6
#480110000000
1!
1%
1-
12
#480120000000
0!
0%
b110 *
0-
02
b110 6
#480130000000
1!
1%
1-
12
#480140000000
0!
0%
b111 *
0-
02
b111 6
#480150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#480160000000
0!
0%
b0 *
0-
02
b0 6
#480170000000
1!
1%
1-
12
#480180000000
0!
0%
b1 *
0-
02
b1 6
#480190000000
1!
1%
1-
12
#480200000000
0!
0%
b10 *
0-
02
b10 6
#480210000000
1!
1%
1-
12
#480220000000
0!
0%
b11 *
0-
02
b11 6
#480230000000
1!
1%
1-
12
15
#480240000000
0!
0%
b100 *
0-
02
b100 6
#480250000000
1!
1%
1-
12
#480260000000
0!
0%
b101 *
0-
02
b101 6
#480270000000
1!
1%
1-
12
#480280000000
0!
0%
b110 *
0-
02
b110 6
#480290000000
1!
1%
1-
12
#480300000000
0!
0%
b111 *
0-
02
b111 6
#480310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#480320000000
0!
0%
b0 *
0-
02
b0 6
#480330000000
1!
1%
1-
12
#480340000000
0!
0%
b1 *
0-
02
b1 6
#480350000000
1!
1%
1-
12
#480360000000
0!
0%
b10 *
0-
02
b10 6
#480370000000
1!
1%
1-
12
#480380000000
0!
0%
b11 *
0-
02
b11 6
#480390000000
1!
1%
1-
12
15
#480400000000
0!
0%
b100 *
0-
02
b100 6
#480410000000
1!
1%
1-
12
#480420000000
0!
0%
b101 *
0-
02
b101 6
#480430000000
1!
1%
1-
12
#480440000000
0!
0%
b110 *
0-
02
b110 6
#480450000000
1!
1%
1-
12
#480460000000
0!
0%
b111 *
0-
02
b111 6
#480470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#480480000000
0!
0%
b0 *
0-
02
b0 6
#480490000000
1!
1%
1-
12
#480500000000
0!
0%
b1 *
0-
02
b1 6
#480510000000
1!
1%
1-
12
#480520000000
0!
0%
b10 *
0-
02
b10 6
#480530000000
1!
1%
1-
12
#480540000000
0!
0%
b11 *
0-
02
b11 6
#480550000000
1!
1%
1-
12
15
#480560000000
0!
0%
b100 *
0-
02
b100 6
#480570000000
1!
1%
1-
12
#480580000000
0!
0%
b101 *
0-
02
b101 6
#480590000000
1!
1%
1-
12
#480600000000
0!
0%
b110 *
0-
02
b110 6
#480610000000
1!
1%
1-
12
#480620000000
0!
0%
b111 *
0-
02
b111 6
#480630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#480640000000
0!
0%
b0 *
0-
02
b0 6
#480650000000
1!
1%
1-
12
#480660000000
0!
0%
b1 *
0-
02
b1 6
#480670000000
1!
1%
1-
12
#480680000000
0!
0%
b10 *
0-
02
b10 6
#480690000000
1!
1%
1-
12
#480700000000
0!
0%
b11 *
0-
02
b11 6
#480710000000
1!
1%
1-
12
15
#480720000000
0!
0%
b100 *
0-
02
b100 6
#480730000000
1!
1%
1-
12
#480740000000
0!
0%
b101 *
0-
02
b101 6
#480750000000
1!
1%
1-
12
#480760000000
0!
0%
b110 *
0-
02
b110 6
#480770000000
1!
1%
1-
12
#480780000000
0!
0%
b111 *
0-
02
b111 6
#480790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#480800000000
0!
0%
b0 *
0-
02
b0 6
#480810000000
1!
1%
1-
12
#480820000000
0!
0%
b1 *
0-
02
b1 6
#480830000000
1!
1%
1-
12
#480840000000
0!
0%
b10 *
0-
02
b10 6
#480850000000
1!
1%
1-
12
#480860000000
0!
0%
b11 *
0-
02
b11 6
#480870000000
1!
1%
1-
12
15
#480880000000
0!
0%
b100 *
0-
02
b100 6
#480890000000
1!
1%
1-
12
#480900000000
0!
0%
b101 *
0-
02
b101 6
#480910000000
1!
1%
1-
12
#480920000000
0!
0%
b110 *
0-
02
b110 6
#480930000000
1!
1%
1-
12
#480940000000
0!
0%
b111 *
0-
02
b111 6
#480950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#480960000000
0!
0%
b0 *
0-
02
b0 6
#480970000000
1!
1%
1-
12
#480980000000
0!
0%
b1 *
0-
02
b1 6
#480990000000
1!
1%
1-
12
#481000000000
0!
0%
b10 *
0-
02
b10 6
#481010000000
1!
1%
1-
12
#481020000000
0!
0%
b11 *
0-
02
b11 6
#481030000000
1!
1%
1-
12
15
#481040000000
0!
0%
b100 *
0-
02
b100 6
#481050000000
1!
1%
1-
12
#481060000000
0!
0%
b101 *
0-
02
b101 6
#481070000000
1!
1%
1-
12
#481080000000
0!
0%
b110 *
0-
02
b110 6
#481090000000
1!
1%
1-
12
#481100000000
0!
0%
b111 *
0-
02
b111 6
#481110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#481120000000
0!
0%
b0 *
0-
02
b0 6
#481130000000
1!
1%
1-
12
#481140000000
0!
0%
b1 *
0-
02
b1 6
#481150000000
1!
1%
1-
12
#481160000000
0!
0%
b10 *
0-
02
b10 6
#481170000000
1!
1%
1-
12
#481180000000
0!
0%
b11 *
0-
02
b11 6
#481190000000
1!
1%
1-
12
15
#481200000000
0!
0%
b100 *
0-
02
b100 6
#481210000000
1!
1%
1-
12
#481220000000
0!
0%
b101 *
0-
02
b101 6
#481230000000
1!
1%
1-
12
#481240000000
0!
0%
b110 *
0-
02
b110 6
#481250000000
1!
1%
1-
12
#481260000000
0!
0%
b111 *
0-
02
b111 6
#481270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#481280000000
0!
0%
b0 *
0-
02
b0 6
#481290000000
1!
1%
1-
12
#481300000000
0!
0%
b1 *
0-
02
b1 6
#481310000000
1!
1%
1-
12
#481320000000
0!
0%
b10 *
0-
02
b10 6
#481330000000
1!
1%
1-
12
#481340000000
0!
0%
b11 *
0-
02
b11 6
#481350000000
1!
1%
1-
12
15
#481360000000
0!
0%
b100 *
0-
02
b100 6
#481370000000
1!
1%
1-
12
#481380000000
0!
0%
b101 *
0-
02
b101 6
#481390000000
1!
1%
1-
12
#481400000000
0!
0%
b110 *
0-
02
b110 6
#481410000000
1!
1%
1-
12
#481420000000
0!
0%
b111 *
0-
02
b111 6
#481430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#481440000000
0!
0%
b0 *
0-
02
b0 6
#481450000000
1!
1%
1-
12
#481460000000
0!
0%
b1 *
0-
02
b1 6
#481470000000
1!
1%
1-
12
#481480000000
0!
0%
b10 *
0-
02
b10 6
#481490000000
1!
1%
1-
12
#481500000000
0!
0%
b11 *
0-
02
b11 6
#481510000000
1!
1%
1-
12
15
#481520000000
0!
0%
b100 *
0-
02
b100 6
#481530000000
1!
1%
1-
12
#481540000000
0!
0%
b101 *
0-
02
b101 6
#481550000000
1!
1%
1-
12
#481560000000
0!
0%
b110 *
0-
02
b110 6
#481570000000
1!
1%
1-
12
#481580000000
0!
0%
b111 *
0-
02
b111 6
#481590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#481600000000
0!
0%
b0 *
0-
02
b0 6
#481610000000
1!
1%
1-
12
#481620000000
0!
0%
b1 *
0-
02
b1 6
#481630000000
1!
1%
1-
12
#481640000000
0!
0%
b10 *
0-
02
b10 6
#481650000000
1!
1%
1-
12
#481660000000
0!
0%
b11 *
0-
02
b11 6
#481670000000
1!
1%
1-
12
15
#481680000000
0!
0%
b100 *
0-
02
b100 6
#481690000000
1!
1%
1-
12
#481700000000
0!
0%
b101 *
0-
02
b101 6
#481710000000
1!
1%
1-
12
#481720000000
0!
0%
b110 *
0-
02
b110 6
#481730000000
1!
1%
1-
12
#481740000000
0!
0%
b111 *
0-
02
b111 6
#481750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#481760000000
0!
0%
b0 *
0-
02
b0 6
#481770000000
1!
1%
1-
12
#481780000000
0!
0%
b1 *
0-
02
b1 6
#481790000000
1!
1%
1-
12
#481800000000
0!
0%
b10 *
0-
02
b10 6
#481810000000
1!
1%
1-
12
#481820000000
0!
0%
b11 *
0-
02
b11 6
#481830000000
1!
1%
1-
12
15
#481840000000
0!
0%
b100 *
0-
02
b100 6
#481850000000
1!
1%
1-
12
#481860000000
0!
0%
b101 *
0-
02
b101 6
#481870000000
1!
1%
1-
12
#481880000000
0!
0%
b110 *
0-
02
b110 6
#481890000000
1!
1%
1-
12
#481900000000
0!
0%
b111 *
0-
02
b111 6
#481910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#481920000000
0!
0%
b0 *
0-
02
b0 6
#481930000000
1!
1%
1-
12
#481940000000
0!
0%
b1 *
0-
02
b1 6
#481950000000
1!
1%
1-
12
#481960000000
0!
0%
b10 *
0-
02
b10 6
#481970000000
1!
1%
1-
12
#481980000000
0!
0%
b11 *
0-
02
b11 6
#481990000000
1!
1%
1-
12
15
#482000000000
0!
0%
b100 *
0-
02
b100 6
#482010000000
1!
1%
1-
12
#482020000000
0!
0%
b101 *
0-
02
b101 6
#482030000000
1!
1%
1-
12
#482040000000
0!
0%
b110 *
0-
02
b110 6
#482050000000
1!
1%
1-
12
#482060000000
0!
0%
b111 *
0-
02
b111 6
#482070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#482080000000
0!
0%
b0 *
0-
02
b0 6
#482090000000
1!
1%
1-
12
#482100000000
0!
0%
b1 *
0-
02
b1 6
#482110000000
1!
1%
1-
12
#482120000000
0!
0%
b10 *
0-
02
b10 6
#482130000000
1!
1%
1-
12
#482140000000
0!
0%
b11 *
0-
02
b11 6
#482150000000
1!
1%
1-
12
15
#482160000000
0!
0%
b100 *
0-
02
b100 6
#482170000000
1!
1%
1-
12
#482180000000
0!
0%
b101 *
0-
02
b101 6
#482190000000
1!
1%
1-
12
#482200000000
0!
0%
b110 *
0-
02
b110 6
#482210000000
1!
1%
1-
12
#482220000000
0!
0%
b111 *
0-
02
b111 6
#482230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#482240000000
0!
0%
b0 *
0-
02
b0 6
#482250000000
1!
1%
1-
12
#482260000000
0!
0%
b1 *
0-
02
b1 6
#482270000000
1!
1%
1-
12
#482280000000
0!
0%
b10 *
0-
02
b10 6
#482290000000
1!
1%
1-
12
#482300000000
0!
0%
b11 *
0-
02
b11 6
#482310000000
1!
1%
1-
12
15
#482320000000
0!
0%
b100 *
0-
02
b100 6
#482330000000
1!
1%
1-
12
#482340000000
0!
0%
b101 *
0-
02
b101 6
#482350000000
1!
1%
1-
12
#482360000000
0!
0%
b110 *
0-
02
b110 6
#482370000000
1!
1%
1-
12
#482380000000
0!
0%
b111 *
0-
02
b111 6
#482390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#482400000000
0!
0%
b0 *
0-
02
b0 6
#482410000000
1!
1%
1-
12
#482420000000
0!
0%
b1 *
0-
02
b1 6
#482430000000
1!
1%
1-
12
#482440000000
0!
0%
b10 *
0-
02
b10 6
#482450000000
1!
1%
1-
12
#482460000000
0!
0%
b11 *
0-
02
b11 6
#482470000000
1!
1%
1-
12
15
#482480000000
0!
0%
b100 *
0-
02
b100 6
#482490000000
1!
1%
1-
12
#482500000000
0!
0%
b101 *
0-
02
b101 6
#482510000000
1!
1%
1-
12
#482520000000
0!
0%
b110 *
0-
02
b110 6
#482530000000
1!
1%
1-
12
#482540000000
0!
0%
b111 *
0-
02
b111 6
#482550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#482560000000
0!
0%
b0 *
0-
02
b0 6
#482570000000
1!
1%
1-
12
#482580000000
0!
0%
b1 *
0-
02
b1 6
#482590000000
1!
1%
1-
12
#482600000000
0!
0%
b10 *
0-
02
b10 6
#482610000000
1!
1%
1-
12
#482620000000
0!
0%
b11 *
0-
02
b11 6
#482630000000
1!
1%
1-
12
15
#482640000000
0!
0%
b100 *
0-
02
b100 6
#482650000000
1!
1%
1-
12
#482660000000
0!
0%
b101 *
0-
02
b101 6
#482670000000
1!
1%
1-
12
#482680000000
0!
0%
b110 *
0-
02
b110 6
#482690000000
1!
1%
1-
12
#482700000000
0!
0%
b111 *
0-
02
b111 6
#482710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#482720000000
0!
0%
b0 *
0-
02
b0 6
#482730000000
1!
1%
1-
12
#482740000000
0!
0%
b1 *
0-
02
b1 6
#482750000000
1!
1%
1-
12
#482760000000
0!
0%
b10 *
0-
02
b10 6
#482770000000
1!
1%
1-
12
#482780000000
0!
0%
b11 *
0-
02
b11 6
#482790000000
1!
1%
1-
12
15
#482800000000
0!
0%
b100 *
0-
02
b100 6
#482810000000
1!
1%
1-
12
#482820000000
0!
0%
b101 *
0-
02
b101 6
#482830000000
1!
1%
1-
12
#482840000000
0!
0%
b110 *
0-
02
b110 6
#482850000000
1!
1%
1-
12
#482860000000
0!
0%
b111 *
0-
02
b111 6
#482870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#482880000000
0!
0%
b0 *
0-
02
b0 6
#482890000000
1!
1%
1-
12
#482900000000
0!
0%
b1 *
0-
02
b1 6
#482910000000
1!
1%
1-
12
#482920000000
0!
0%
b10 *
0-
02
b10 6
#482930000000
1!
1%
1-
12
#482940000000
0!
0%
b11 *
0-
02
b11 6
#482950000000
1!
1%
1-
12
15
#482960000000
0!
0%
b100 *
0-
02
b100 6
#482970000000
1!
1%
1-
12
#482980000000
0!
0%
b101 *
0-
02
b101 6
#482990000000
1!
1%
1-
12
#483000000000
0!
0%
b110 *
0-
02
b110 6
#483010000000
1!
1%
1-
12
#483020000000
0!
0%
b111 *
0-
02
b111 6
#483030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#483040000000
0!
0%
b0 *
0-
02
b0 6
#483050000000
1!
1%
1-
12
#483060000000
0!
0%
b1 *
0-
02
b1 6
#483070000000
1!
1%
1-
12
#483080000000
0!
0%
b10 *
0-
02
b10 6
#483090000000
1!
1%
1-
12
#483100000000
0!
0%
b11 *
0-
02
b11 6
#483110000000
1!
1%
1-
12
15
#483120000000
0!
0%
b100 *
0-
02
b100 6
#483130000000
1!
1%
1-
12
#483140000000
0!
0%
b101 *
0-
02
b101 6
#483150000000
1!
1%
1-
12
#483160000000
0!
0%
b110 *
0-
02
b110 6
#483170000000
1!
1%
1-
12
#483180000000
0!
0%
b111 *
0-
02
b111 6
#483190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#483200000000
0!
0%
b0 *
0-
02
b0 6
#483210000000
1!
1%
1-
12
#483220000000
0!
0%
b1 *
0-
02
b1 6
#483230000000
1!
1%
1-
12
#483240000000
0!
0%
b10 *
0-
02
b10 6
#483250000000
1!
1%
1-
12
#483260000000
0!
0%
b11 *
0-
02
b11 6
#483270000000
1!
1%
1-
12
15
#483280000000
0!
0%
b100 *
0-
02
b100 6
#483290000000
1!
1%
1-
12
#483300000000
0!
0%
b101 *
0-
02
b101 6
#483310000000
1!
1%
1-
12
#483320000000
0!
0%
b110 *
0-
02
b110 6
#483330000000
1!
1%
1-
12
#483340000000
0!
0%
b111 *
0-
02
b111 6
#483350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#483360000000
0!
0%
b0 *
0-
02
b0 6
#483370000000
1!
1%
1-
12
#483380000000
0!
0%
b1 *
0-
02
b1 6
#483390000000
1!
1%
1-
12
#483400000000
0!
0%
b10 *
0-
02
b10 6
#483410000000
1!
1%
1-
12
#483420000000
0!
0%
b11 *
0-
02
b11 6
#483430000000
1!
1%
1-
12
15
#483440000000
0!
0%
b100 *
0-
02
b100 6
#483450000000
1!
1%
1-
12
#483460000000
0!
0%
b101 *
0-
02
b101 6
#483470000000
1!
1%
1-
12
#483480000000
0!
0%
b110 *
0-
02
b110 6
#483490000000
1!
1%
1-
12
#483500000000
0!
0%
b111 *
0-
02
b111 6
#483510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#483520000000
0!
0%
b0 *
0-
02
b0 6
#483530000000
1!
1%
1-
12
#483540000000
0!
0%
b1 *
0-
02
b1 6
#483550000000
1!
1%
1-
12
#483560000000
0!
0%
b10 *
0-
02
b10 6
#483570000000
1!
1%
1-
12
#483580000000
0!
0%
b11 *
0-
02
b11 6
#483590000000
1!
1%
1-
12
15
#483600000000
0!
0%
b100 *
0-
02
b100 6
#483610000000
1!
1%
1-
12
#483620000000
0!
0%
b101 *
0-
02
b101 6
#483630000000
1!
1%
1-
12
#483640000000
0!
0%
b110 *
0-
02
b110 6
#483650000000
1!
1%
1-
12
#483660000000
0!
0%
b111 *
0-
02
b111 6
#483670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#483680000000
0!
0%
b0 *
0-
02
b0 6
#483690000000
1!
1%
1-
12
#483700000000
0!
0%
b1 *
0-
02
b1 6
#483710000000
1!
1%
1-
12
#483720000000
0!
0%
b10 *
0-
02
b10 6
#483730000000
1!
1%
1-
12
#483740000000
0!
0%
b11 *
0-
02
b11 6
#483750000000
1!
1%
1-
12
15
#483760000000
0!
0%
b100 *
0-
02
b100 6
#483770000000
1!
1%
1-
12
#483780000000
0!
0%
b101 *
0-
02
b101 6
#483790000000
1!
1%
1-
12
#483800000000
0!
0%
b110 *
0-
02
b110 6
#483810000000
1!
1%
1-
12
#483820000000
0!
0%
b111 *
0-
02
b111 6
#483830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#483840000000
0!
0%
b0 *
0-
02
b0 6
#483850000000
1!
1%
1-
12
#483860000000
0!
0%
b1 *
0-
02
b1 6
#483870000000
1!
1%
1-
12
#483880000000
0!
0%
b10 *
0-
02
b10 6
#483890000000
1!
1%
1-
12
#483900000000
0!
0%
b11 *
0-
02
b11 6
#483910000000
1!
1%
1-
12
15
#483920000000
0!
0%
b100 *
0-
02
b100 6
#483930000000
1!
1%
1-
12
#483940000000
0!
0%
b101 *
0-
02
b101 6
#483950000000
1!
1%
1-
12
#483960000000
0!
0%
b110 *
0-
02
b110 6
#483970000000
1!
1%
1-
12
#483980000000
0!
0%
b111 *
0-
02
b111 6
#483990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#484000000000
0!
0%
b0 *
0-
02
b0 6
#484010000000
1!
1%
1-
12
#484020000000
0!
0%
b1 *
0-
02
b1 6
#484030000000
1!
1%
1-
12
#484040000000
0!
0%
b10 *
0-
02
b10 6
#484050000000
1!
1%
1-
12
#484060000000
0!
0%
b11 *
0-
02
b11 6
#484070000000
1!
1%
1-
12
15
#484080000000
0!
0%
b100 *
0-
02
b100 6
#484090000000
1!
1%
1-
12
#484100000000
0!
0%
b101 *
0-
02
b101 6
#484110000000
1!
1%
1-
12
#484120000000
0!
0%
b110 *
0-
02
b110 6
#484130000000
1!
1%
1-
12
#484140000000
0!
0%
b111 *
0-
02
b111 6
#484150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#484160000000
0!
0%
b0 *
0-
02
b0 6
#484170000000
1!
1%
1-
12
#484180000000
0!
0%
b1 *
0-
02
b1 6
#484190000000
1!
1%
1-
12
#484200000000
0!
0%
b10 *
0-
02
b10 6
#484210000000
1!
1%
1-
12
#484220000000
0!
0%
b11 *
0-
02
b11 6
#484230000000
1!
1%
1-
12
15
#484240000000
0!
0%
b100 *
0-
02
b100 6
#484250000000
1!
1%
1-
12
#484260000000
0!
0%
b101 *
0-
02
b101 6
#484270000000
1!
1%
1-
12
#484280000000
0!
0%
b110 *
0-
02
b110 6
#484290000000
1!
1%
1-
12
#484300000000
0!
0%
b111 *
0-
02
b111 6
#484310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#484320000000
0!
0%
b0 *
0-
02
b0 6
#484330000000
1!
1%
1-
12
#484340000000
0!
0%
b1 *
0-
02
b1 6
#484350000000
1!
1%
1-
12
#484360000000
0!
0%
b10 *
0-
02
b10 6
#484370000000
1!
1%
1-
12
#484380000000
0!
0%
b11 *
0-
02
b11 6
#484390000000
1!
1%
1-
12
15
#484400000000
0!
0%
b100 *
0-
02
b100 6
#484410000000
1!
1%
1-
12
#484420000000
0!
0%
b101 *
0-
02
b101 6
#484430000000
1!
1%
1-
12
#484440000000
0!
0%
b110 *
0-
02
b110 6
#484450000000
1!
1%
1-
12
#484460000000
0!
0%
b111 *
0-
02
b111 6
#484470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#484480000000
0!
0%
b0 *
0-
02
b0 6
#484490000000
1!
1%
1-
12
#484500000000
0!
0%
b1 *
0-
02
b1 6
#484510000000
1!
1%
1-
12
#484520000000
0!
0%
b10 *
0-
02
b10 6
#484530000000
1!
1%
1-
12
#484540000000
0!
0%
b11 *
0-
02
b11 6
#484550000000
1!
1%
1-
12
15
#484560000000
0!
0%
b100 *
0-
02
b100 6
#484570000000
1!
1%
1-
12
#484580000000
0!
0%
b101 *
0-
02
b101 6
#484590000000
1!
1%
1-
12
#484600000000
0!
0%
b110 *
0-
02
b110 6
#484610000000
1!
1%
1-
12
#484620000000
0!
0%
b111 *
0-
02
b111 6
#484630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#484640000000
0!
0%
b0 *
0-
02
b0 6
#484650000000
1!
1%
1-
12
#484660000000
0!
0%
b1 *
0-
02
b1 6
#484670000000
1!
1%
1-
12
#484680000000
0!
0%
b10 *
0-
02
b10 6
#484690000000
1!
1%
1-
12
#484700000000
0!
0%
b11 *
0-
02
b11 6
#484710000000
1!
1%
1-
12
15
#484720000000
0!
0%
b100 *
0-
02
b100 6
#484730000000
1!
1%
1-
12
#484740000000
0!
0%
b101 *
0-
02
b101 6
#484750000000
1!
1%
1-
12
#484760000000
0!
0%
b110 *
0-
02
b110 6
#484770000000
1!
1%
1-
12
#484780000000
0!
0%
b111 *
0-
02
b111 6
#484790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#484800000000
0!
0%
b0 *
0-
02
b0 6
#484810000000
1!
1%
1-
12
#484820000000
0!
0%
b1 *
0-
02
b1 6
#484830000000
1!
1%
1-
12
#484840000000
0!
0%
b10 *
0-
02
b10 6
#484850000000
1!
1%
1-
12
#484860000000
0!
0%
b11 *
0-
02
b11 6
#484870000000
1!
1%
1-
12
15
#484880000000
0!
0%
b100 *
0-
02
b100 6
#484890000000
1!
1%
1-
12
#484900000000
0!
0%
b101 *
0-
02
b101 6
#484910000000
1!
1%
1-
12
#484920000000
0!
0%
b110 *
0-
02
b110 6
#484930000000
1!
1%
1-
12
#484940000000
0!
0%
b111 *
0-
02
b111 6
#484950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#484960000000
0!
0%
b0 *
0-
02
b0 6
#484970000000
1!
1%
1-
12
#484980000000
0!
0%
b1 *
0-
02
b1 6
#484990000000
1!
1%
1-
12
#485000000000
0!
0%
b10 *
0-
02
b10 6
#485010000000
1!
1%
1-
12
#485020000000
0!
0%
b11 *
0-
02
b11 6
#485030000000
1!
1%
1-
12
15
#485040000000
0!
0%
b100 *
0-
02
b100 6
#485050000000
1!
1%
1-
12
#485060000000
0!
0%
b101 *
0-
02
b101 6
#485070000000
1!
1%
1-
12
#485080000000
0!
0%
b110 *
0-
02
b110 6
#485090000000
1!
1%
1-
12
#485100000000
0!
0%
b111 *
0-
02
b111 6
#485110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#485120000000
0!
0%
b0 *
0-
02
b0 6
#485130000000
1!
1%
1-
12
#485140000000
0!
0%
b1 *
0-
02
b1 6
#485150000000
1!
1%
1-
12
#485160000000
0!
0%
b10 *
0-
02
b10 6
#485170000000
1!
1%
1-
12
#485180000000
0!
0%
b11 *
0-
02
b11 6
#485190000000
1!
1%
1-
12
15
#485200000000
0!
0%
b100 *
0-
02
b100 6
#485210000000
1!
1%
1-
12
#485220000000
0!
0%
b101 *
0-
02
b101 6
#485230000000
1!
1%
1-
12
#485240000000
0!
0%
b110 *
0-
02
b110 6
#485250000000
1!
1%
1-
12
#485260000000
0!
0%
b111 *
0-
02
b111 6
#485270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#485280000000
0!
0%
b0 *
0-
02
b0 6
#485290000000
1!
1%
1-
12
#485300000000
0!
0%
b1 *
0-
02
b1 6
#485310000000
1!
1%
1-
12
#485320000000
0!
0%
b10 *
0-
02
b10 6
#485330000000
1!
1%
1-
12
#485340000000
0!
0%
b11 *
0-
02
b11 6
#485350000000
1!
1%
1-
12
15
#485360000000
0!
0%
b100 *
0-
02
b100 6
#485370000000
1!
1%
1-
12
#485380000000
0!
0%
b101 *
0-
02
b101 6
#485390000000
1!
1%
1-
12
#485400000000
0!
0%
b110 *
0-
02
b110 6
#485410000000
1!
1%
1-
12
#485420000000
0!
0%
b111 *
0-
02
b111 6
#485430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#485440000000
0!
0%
b0 *
0-
02
b0 6
#485450000000
1!
1%
1-
12
#485460000000
0!
0%
b1 *
0-
02
b1 6
#485470000000
1!
1%
1-
12
#485480000000
0!
0%
b10 *
0-
02
b10 6
#485490000000
1!
1%
1-
12
#485500000000
0!
0%
b11 *
0-
02
b11 6
#485510000000
1!
1%
1-
12
15
#485520000000
0!
0%
b100 *
0-
02
b100 6
#485530000000
1!
1%
1-
12
#485540000000
0!
0%
b101 *
0-
02
b101 6
#485550000000
1!
1%
1-
12
#485560000000
0!
0%
b110 *
0-
02
b110 6
#485570000000
1!
1%
1-
12
#485580000000
0!
0%
b111 *
0-
02
b111 6
#485590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#485600000000
0!
0%
b0 *
0-
02
b0 6
#485610000000
1!
1%
1-
12
#485620000000
0!
0%
b1 *
0-
02
b1 6
#485630000000
1!
1%
1-
12
#485640000000
0!
0%
b10 *
0-
02
b10 6
#485650000000
1!
1%
1-
12
#485660000000
0!
0%
b11 *
0-
02
b11 6
#485670000000
1!
1%
1-
12
15
#485680000000
0!
0%
b100 *
0-
02
b100 6
#485690000000
1!
1%
1-
12
#485700000000
0!
0%
b101 *
0-
02
b101 6
#485710000000
1!
1%
1-
12
#485720000000
0!
0%
b110 *
0-
02
b110 6
#485730000000
1!
1%
1-
12
#485740000000
0!
0%
b111 *
0-
02
b111 6
#485750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#485760000000
0!
0%
b0 *
0-
02
b0 6
#485770000000
1!
1%
1-
12
#485780000000
0!
0%
b1 *
0-
02
b1 6
#485790000000
1!
1%
1-
12
#485800000000
0!
0%
b10 *
0-
02
b10 6
#485810000000
1!
1%
1-
12
#485820000000
0!
0%
b11 *
0-
02
b11 6
#485830000000
1!
1%
1-
12
15
#485840000000
0!
0%
b100 *
0-
02
b100 6
#485850000000
1!
1%
1-
12
#485860000000
0!
0%
b101 *
0-
02
b101 6
#485870000000
1!
1%
1-
12
#485880000000
0!
0%
b110 *
0-
02
b110 6
#485890000000
1!
1%
1-
12
#485900000000
0!
0%
b111 *
0-
02
b111 6
#485910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#485920000000
0!
0%
b0 *
0-
02
b0 6
#485930000000
1!
1%
1-
12
#485940000000
0!
0%
b1 *
0-
02
b1 6
#485950000000
1!
1%
1-
12
#485960000000
0!
0%
b10 *
0-
02
b10 6
#485970000000
1!
1%
1-
12
#485980000000
0!
0%
b11 *
0-
02
b11 6
#485990000000
1!
1%
1-
12
15
#486000000000
0!
0%
b100 *
0-
02
b100 6
#486010000000
1!
1%
1-
12
#486020000000
0!
0%
b101 *
0-
02
b101 6
#486030000000
1!
1%
1-
12
#486040000000
0!
0%
b110 *
0-
02
b110 6
#486050000000
1!
1%
1-
12
#486060000000
0!
0%
b111 *
0-
02
b111 6
#486070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#486080000000
0!
0%
b0 *
0-
02
b0 6
#486090000000
1!
1%
1-
12
#486100000000
0!
0%
b1 *
0-
02
b1 6
#486110000000
1!
1%
1-
12
#486120000000
0!
0%
b10 *
0-
02
b10 6
#486130000000
1!
1%
1-
12
#486140000000
0!
0%
b11 *
0-
02
b11 6
#486150000000
1!
1%
1-
12
15
#486160000000
0!
0%
b100 *
0-
02
b100 6
#486170000000
1!
1%
1-
12
#486180000000
0!
0%
b101 *
0-
02
b101 6
#486190000000
1!
1%
1-
12
#486200000000
0!
0%
b110 *
0-
02
b110 6
#486210000000
1!
1%
1-
12
#486220000000
0!
0%
b111 *
0-
02
b111 6
#486230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#486240000000
0!
0%
b0 *
0-
02
b0 6
#486250000000
1!
1%
1-
12
#486260000000
0!
0%
b1 *
0-
02
b1 6
#486270000000
1!
1%
1-
12
#486280000000
0!
0%
b10 *
0-
02
b10 6
#486290000000
1!
1%
1-
12
#486300000000
0!
0%
b11 *
0-
02
b11 6
#486310000000
1!
1%
1-
12
15
#486320000000
0!
0%
b100 *
0-
02
b100 6
#486330000000
1!
1%
1-
12
#486340000000
0!
0%
b101 *
0-
02
b101 6
#486350000000
1!
1%
1-
12
#486360000000
0!
0%
b110 *
0-
02
b110 6
#486370000000
1!
1%
1-
12
#486380000000
0!
0%
b111 *
0-
02
b111 6
#486390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#486400000000
0!
0%
b0 *
0-
02
b0 6
#486410000000
1!
1%
1-
12
#486420000000
0!
0%
b1 *
0-
02
b1 6
#486430000000
1!
1%
1-
12
#486440000000
0!
0%
b10 *
0-
02
b10 6
#486450000000
1!
1%
1-
12
#486460000000
0!
0%
b11 *
0-
02
b11 6
#486470000000
1!
1%
1-
12
15
#486480000000
0!
0%
b100 *
0-
02
b100 6
#486490000000
1!
1%
1-
12
#486500000000
0!
0%
b101 *
0-
02
b101 6
#486510000000
1!
1%
1-
12
#486520000000
0!
0%
b110 *
0-
02
b110 6
#486530000000
1!
1%
1-
12
#486540000000
0!
0%
b111 *
0-
02
b111 6
#486550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#486560000000
0!
0%
b0 *
0-
02
b0 6
#486570000000
1!
1%
1-
12
#486580000000
0!
0%
b1 *
0-
02
b1 6
#486590000000
1!
1%
1-
12
#486600000000
0!
0%
b10 *
0-
02
b10 6
#486610000000
1!
1%
1-
12
#486620000000
0!
0%
b11 *
0-
02
b11 6
#486630000000
1!
1%
1-
12
15
#486640000000
0!
0%
b100 *
0-
02
b100 6
#486650000000
1!
1%
1-
12
#486660000000
0!
0%
b101 *
0-
02
b101 6
#486670000000
1!
1%
1-
12
#486680000000
0!
0%
b110 *
0-
02
b110 6
#486690000000
1!
1%
1-
12
#486700000000
0!
0%
b111 *
0-
02
b111 6
#486710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#486720000000
0!
0%
b0 *
0-
02
b0 6
#486730000000
1!
1%
1-
12
#486740000000
0!
0%
b1 *
0-
02
b1 6
#486750000000
1!
1%
1-
12
#486760000000
0!
0%
b10 *
0-
02
b10 6
#486770000000
1!
1%
1-
12
#486780000000
0!
0%
b11 *
0-
02
b11 6
#486790000000
1!
1%
1-
12
15
#486800000000
0!
0%
b100 *
0-
02
b100 6
#486810000000
1!
1%
1-
12
#486820000000
0!
0%
b101 *
0-
02
b101 6
#486830000000
1!
1%
1-
12
#486840000000
0!
0%
b110 *
0-
02
b110 6
#486850000000
1!
1%
1-
12
#486860000000
0!
0%
b111 *
0-
02
b111 6
#486870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#486880000000
0!
0%
b0 *
0-
02
b0 6
#486890000000
1!
1%
1-
12
#486900000000
0!
0%
b1 *
0-
02
b1 6
#486910000000
1!
1%
1-
12
#486920000000
0!
0%
b10 *
0-
02
b10 6
#486930000000
1!
1%
1-
12
#486940000000
0!
0%
b11 *
0-
02
b11 6
#486950000000
1!
1%
1-
12
15
#486960000000
0!
0%
b100 *
0-
02
b100 6
#486970000000
1!
1%
1-
12
#486980000000
0!
0%
b101 *
0-
02
b101 6
#486990000000
1!
1%
1-
12
#487000000000
0!
0%
b110 *
0-
02
b110 6
#487010000000
1!
1%
1-
12
#487020000000
0!
0%
b111 *
0-
02
b111 6
#487030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#487040000000
0!
0%
b0 *
0-
02
b0 6
#487050000000
1!
1%
1-
12
#487060000000
0!
0%
b1 *
0-
02
b1 6
#487070000000
1!
1%
1-
12
#487080000000
0!
0%
b10 *
0-
02
b10 6
#487090000000
1!
1%
1-
12
#487100000000
0!
0%
b11 *
0-
02
b11 6
#487110000000
1!
1%
1-
12
15
#487120000000
0!
0%
b100 *
0-
02
b100 6
#487130000000
1!
1%
1-
12
#487140000000
0!
0%
b101 *
0-
02
b101 6
#487150000000
1!
1%
1-
12
#487160000000
0!
0%
b110 *
0-
02
b110 6
#487170000000
1!
1%
1-
12
#487180000000
0!
0%
b111 *
0-
02
b111 6
#487190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#487200000000
0!
0%
b0 *
0-
02
b0 6
#487210000000
1!
1%
1-
12
#487220000000
0!
0%
b1 *
0-
02
b1 6
#487230000000
1!
1%
1-
12
#487240000000
0!
0%
b10 *
0-
02
b10 6
#487250000000
1!
1%
1-
12
#487260000000
0!
0%
b11 *
0-
02
b11 6
#487270000000
1!
1%
1-
12
15
#487280000000
0!
0%
b100 *
0-
02
b100 6
#487290000000
1!
1%
1-
12
#487300000000
0!
0%
b101 *
0-
02
b101 6
#487310000000
1!
1%
1-
12
#487320000000
0!
0%
b110 *
0-
02
b110 6
#487330000000
1!
1%
1-
12
#487340000000
0!
0%
b111 *
0-
02
b111 6
#487350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#487360000000
0!
0%
b0 *
0-
02
b0 6
#487370000000
1!
1%
1-
12
#487380000000
0!
0%
b1 *
0-
02
b1 6
#487390000000
1!
1%
1-
12
#487400000000
0!
0%
b10 *
0-
02
b10 6
#487410000000
1!
1%
1-
12
#487420000000
0!
0%
b11 *
0-
02
b11 6
#487430000000
1!
1%
1-
12
15
#487440000000
0!
0%
b100 *
0-
02
b100 6
#487450000000
1!
1%
1-
12
#487460000000
0!
0%
b101 *
0-
02
b101 6
#487470000000
1!
1%
1-
12
#487480000000
0!
0%
b110 *
0-
02
b110 6
#487490000000
1!
1%
1-
12
#487500000000
0!
0%
b111 *
0-
02
b111 6
#487510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#487520000000
0!
0%
b0 *
0-
02
b0 6
#487530000000
1!
1%
1-
12
#487540000000
0!
0%
b1 *
0-
02
b1 6
#487550000000
1!
1%
1-
12
#487560000000
0!
0%
b10 *
0-
02
b10 6
#487570000000
1!
1%
1-
12
#487580000000
0!
0%
b11 *
0-
02
b11 6
#487590000000
1!
1%
1-
12
15
#487600000000
0!
0%
b100 *
0-
02
b100 6
#487610000000
1!
1%
1-
12
#487620000000
0!
0%
b101 *
0-
02
b101 6
#487630000000
1!
1%
1-
12
#487640000000
0!
0%
b110 *
0-
02
b110 6
#487650000000
1!
1%
1-
12
#487660000000
0!
0%
b111 *
0-
02
b111 6
#487670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#487680000000
0!
0%
b0 *
0-
02
b0 6
#487690000000
1!
1%
1-
12
#487700000000
0!
0%
b1 *
0-
02
b1 6
#487710000000
1!
1%
1-
12
#487720000000
0!
0%
b10 *
0-
02
b10 6
#487730000000
1!
1%
1-
12
#487740000000
0!
0%
b11 *
0-
02
b11 6
#487750000000
1!
1%
1-
12
15
#487760000000
0!
0%
b100 *
0-
02
b100 6
#487770000000
1!
1%
1-
12
#487780000000
0!
0%
b101 *
0-
02
b101 6
#487790000000
1!
1%
1-
12
#487800000000
0!
0%
b110 *
0-
02
b110 6
#487810000000
1!
1%
1-
12
#487820000000
0!
0%
b111 *
0-
02
b111 6
#487830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#487840000000
0!
0%
b0 *
0-
02
b0 6
#487850000000
1!
1%
1-
12
#487860000000
0!
0%
b1 *
0-
02
b1 6
#487870000000
1!
1%
1-
12
#487880000000
0!
0%
b10 *
0-
02
b10 6
#487890000000
1!
1%
1-
12
#487900000000
0!
0%
b11 *
0-
02
b11 6
#487910000000
1!
1%
1-
12
15
#487920000000
0!
0%
b100 *
0-
02
b100 6
#487930000000
1!
1%
1-
12
#487940000000
0!
0%
b101 *
0-
02
b101 6
#487950000000
1!
1%
1-
12
#487960000000
0!
0%
b110 *
0-
02
b110 6
#487970000000
1!
1%
1-
12
#487980000000
0!
0%
b111 *
0-
02
b111 6
#487990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#488000000000
0!
0%
b0 *
0-
02
b0 6
#488010000000
1!
1%
1-
12
#488020000000
0!
0%
b1 *
0-
02
b1 6
#488030000000
1!
1%
1-
12
#488040000000
0!
0%
b10 *
0-
02
b10 6
#488050000000
1!
1%
1-
12
#488060000000
0!
0%
b11 *
0-
02
b11 6
#488070000000
1!
1%
1-
12
15
#488080000000
0!
0%
b100 *
0-
02
b100 6
#488090000000
1!
1%
1-
12
#488100000000
0!
0%
b101 *
0-
02
b101 6
#488110000000
1!
1%
1-
12
#488120000000
0!
0%
b110 *
0-
02
b110 6
#488130000000
1!
1%
1-
12
#488140000000
0!
0%
b111 *
0-
02
b111 6
#488150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#488160000000
0!
0%
b0 *
0-
02
b0 6
#488170000000
1!
1%
1-
12
#488180000000
0!
0%
b1 *
0-
02
b1 6
#488190000000
1!
1%
1-
12
#488200000000
0!
0%
b10 *
0-
02
b10 6
#488210000000
1!
1%
1-
12
#488220000000
0!
0%
b11 *
0-
02
b11 6
#488230000000
1!
1%
1-
12
15
#488240000000
0!
0%
b100 *
0-
02
b100 6
#488250000000
1!
1%
1-
12
#488260000000
0!
0%
b101 *
0-
02
b101 6
#488270000000
1!
1%
1-
12
#488280000000
0!
0%
b110 *
0-
02
b110 6
#488290000000
1!
1%
1-
12
#488300000000
0!
0%
b111 *
0-
02
b111 6
#488310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#488320000000
0!
0%
b0 *
0-
02
b0 6
#488330000000
1!
1%
1-
12
#488340000000
0!
0%
b1 *
0-
02
b1 6
#488350000000
1!
1%
1-
12
#488360000000
0!
0%
b10 *
0-
02
b10 6
#488370000000
1!
1%
1-
12
#488380000000
0!
0%
b11 *
0-
02
b11 6
#488390000000
1!
1%
1-
12
15
#488400000000
0!
0%
b100 *
0-
02
b100 6
#488410000000
1!
1%
1-
12
#488420000000
0!
0%
b101 *
0-
02
b101 6
#488430000000
1!
1%
1-
12
#488440000000
0!
0%
b110 *
0-
02
b110 6
#488450000000
1!
1%
1-
12
#488460000000
0!
0%
b111 *
0-
02
b111 6
#488470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#488480000000
0!
0%
b0 *
0-
02
b0 6
#488490000000
1!
1%
1-
12
#488500000000
0!
0%
b1 *
0-
02
b1 6
#488510000000
1!
1%
1-
12
#488520000000
0!
0%
b10 *
0-
02
b10 6
#488530000000
1!
1%
1-
12
#488540000000
0!
0%
b11 *
0-
02
b11 6
#488550000000
1!
1%
1-
12
15
#488560000000
0!
0%
b100 *
0-
02
b100 6
#488570000000
1!
1%
1-
12
#488580000000
0!
0%
b101 *
0-
02
b101 6
#488590000000
1!
1%
1-
12
#488600000000
0!
0%
b110 *
0-
02
b110 6
#488610000000
1!
1%
1-
12
#488620000000
0!
0%
b111 *
0-
02
b111 6
#488630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#488640000000
0!
0%
b0 *
0-
02
b0 6
#488650000000
1!
1%
1-
12
#488660000000
0!
0%
b1 *
0-
02
b1 6
#488670000000
1!
1%
1-
12
#488680000000
0!
0%
b10 *
0-
02
b10 6
#488690000000
1!
1%
1-
12
#488700000000
0!
0%
b11 *
0-
02
b11 6
#488710000000
1!
1%
1-
12
15
#488720000000
0!
0%
b100 *
0-
02
b100 6
#488730000000
1!
1%
1-
12
#488740000000
0!
0%
b101 *
0-
02
b101 6
#488750000000
1!
1%
1-
12
#488760000000
0!
0%
b110 *
0-
02
b110 6
#488770000000
1!
1%
1-
12
#488780000000
0!
0%
b111 *
0-
02
b111 6
#488790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#488800000000
0!
0%
b0 *
0-
02
b0 6
#488810000000
1!
1%
1-
12
#488820000000
0!
0%
b1 *
0-
02
b1 6
#488830000000
1!
1%
1-
12
#488840000000
0!
0%
b10 *
0-
02
b10 6
#488850000000
1!
1%
1-
12
#488860000000
0!
0%
b11 *
0-
02
b11 6
#488870000000
1!
1%
1-
12
15
#488880000000
0!
0%
b100 *
0-
02
b100 6
#488890000000
1!
1%
1-
12
#488900000000
0!
0%
b101 *
0-
02
b101 6
#488910000000
1!
1%
1-
12
#488920000000
0!
0%
b110 *
0-
02
b110 6
#488930000000
1!
1%
1-
12
#488940000000
0!
0%
b111 *
0-
02
b111 6
#488950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#488960000000
0!
0%
b0 *
0-
02
b0 6
#488970000000
1!
1%
1-
12
#488980000000
0!
0%
b1 *
0-
02
b1 6
#488990000000
1!
1%
1-
12
#489000000000
0!
0%
b10 *
0-
02
b10 6
#489010000000
1!
1%
1-
12
#489020000000
0!
0%
b11 *
0-
02
b11 6
#489030000000
1!
1%
1-
12
15
#489040000000
0!
0%
b100 *
0-
02
b100 6
#489050000000
1!
1%
1-
12
#489060000000
0!
0%
b101 *
0-
02
b101 6
#489070000000
1!
1%
1-
12
#489080000000
0!
0%
b110 *
0-
02
b110 6
#489090000000
1!
1%
1-
12
#489100000000
0!
0%
b111 *
0-
02
b111 6
#489110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#489120000000
0!
0%
b0 *
0-
02
b0 6
#489130000000
1!
1%
1-
12
#489140000000
0!
0%
b1 *
0-
02
b1 6
#489150000000
1!
1%
1-
12
#489160000000
0!
0%
b10 *
0-
02
b10 6
#489170000000
1!
1%
1-
12
#489180000000
0!
0%
b11 *
0-
02
b11 6
#489190000000
1!
1%
1-
12
15
#489200000000
0!
0%
b100 *
0-
02
b100 6
#489210000000
1!
1%
1-
12
#489220000000
0!
0%
b101 *
0-
02
b101 6
#489230000000
1!
1%
1-
12
#489240000000
0!
0%
b110 *
0-
02
b110 6
#489250000000
1!
1%
1-
12
#489260000000
0!
0%
b111 *
0-
02
b111 6
#489270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#489280000000
0!
0%
b0 *
0-
02
b0 6
#489290000000
1!
1%
1-
12
#489300000000
0!
0%
b1 *
0-
02
b1 6
#489310000000
1!
1%
1-
12
#489320000000
0!
0%
b10 *
0-
02
b10 6
#489330000000
1!
1%
1-
12
#489340000000
0!
0%
b11 *
0-
02
b11 6
#489350000000
1!
1%
1-
12
15
#489360000000
0!
0%
b100 *
0-
02
b100 6
#489370000000
1!
1%
1-
12
#489380000000
0!
0%
b101 *
0-
02
b101 6
#489390000000
1!
1%
1-
12
#489400000000
0!
0%
b110 *
0-
02
b110 6
#489410000000
1!
1%
1-
12
#489420000000
0!
0%
b111 *
0-
02
b111 6
#489430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#489440000000
0!
0%
b0 *
0-
02
b0 6
#489450000000
1!
1%
1-
12
#489460000000
0!
0%
b1 *
0-
02
b1 6
#489470000000
1!
1%
1-
12
#489480000000
0!
0%
b10 *
0-
02
b10 6
#489490000000
1!
1%
1-
12
#489500000000
0!
0%
b11 *
0-
02
b11 6
#489510000000
1!
1%
1-
12
15
#489520000000
0!
0%
b100 *
0-
02
b100 6
#489530000000
1!
1%
1-
12
#489540000000
0!
0%
b101 *
0-
02
b101 6
#489550000000
1!
1%
1-
12
#489560000000
0!
0%
b110 *
0-
02
b110 6
#489570000000
1!
1%
1-
12
#489580000000
0!
0%
b111 *
0-
02
b111 6
#489590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#489600000000
0!
0%
b0 *
0-
02
b0 6
#489610000000
1!
1%
1-
12
#489620000000
0!
0%
b1 *
0-
02
b1 6
#489630000000
1!
1%
1-
12
#489640000000
0!
0%
b10 *
0-
02
b10 6
#489650000000
1!
1%
1-
12
#489660000000
0!
0%
b11 *
0-
02
b11 6
#489670000000
1!
1%
1-
12
15
#489680000000
0!
0%
b100 *
0-
02
b100 6
#489690000000
1!
1%
1-
12
#489700000000
0!
0%
b101 *
0-
02
b101 6
#489710000000
1!
1%
1-
12
#489720000000
0!
0%
b110 *
0-
02
b110 6
#489730000000
1!
1%
1-
12
#489740000000
0!
0%
b111 *
0-
02
b111 6
#489750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#489760000000
0!
0%
b0 *
0-
02
b0 6
#489770000000
1!
1%
1-
12
#489780000000
0!
0%
b1 *
0-
02
b1 6
#489790000000
1!
1%
1-
12
#489800000000
0!
0%
b10 *
0-
02
b10 6
#489810000000
1!
1%
1-
12
#489820000000
0!
0%
b11 *
0-
02
b11 6
#489830000000
1!
1%
1-
12
15
#489840000000
0!
0%
b100 *
0-
02
b100 6
#489850000000
1!
1%
1-
12
#489860000000
0!
0%
b101 *
0-
02
b101 6
#489870000000
1!
1%
1-
12
#489880000000
0!
0%
b110 *
0-
02
b110 6
#489890000000
1!
1%
1-
12
#489900000000
0!
0%
b111 *
0-
02
b111 6
#489910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#489920000000
0!
0%
b0 *
0-
02
b0 6
#489930000000
1!
1%
1-
12
#489940000000
0!
0%
b1 *
0-
02
b1 6
#489950000000
1!
1%
1-
12
#489960000000
0!
0%
b10 *
0-
02
b10 6
#489970000000
1!
1%
1-
12
#489980000000
0!
0%
b11 *
0-
02
b11 6
#489990000000
1!
1%
1-
12
15
#490000000000
0!
0%
b100 *
0-
02
b100 6
#490010000000
1!
1%
1-
12
#490020000000
0!
0%
b101 *
0-
02
b101 6
#490030000000
1!
1%
1-
12
#490040000000
0!
0%
b110 *
0-
02
b110 6
#490050000000
1!
1%
1-
12
#490060000000
0!
0%
b111 *
0-
02
b111 6
#490070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#490080000000
0!
0%
b0 *
0-
02
b0 6
#490090000000
1!
1%
1-
12
#490100000000
0!
0%
b1 *
0-
02
b1 6
#490110000000
1!
1%
1-
12
#490120000000
0!
0%
b10 *
0-
02
b10 6
#490130000000
1!
1%
1-
12
#490140000000
0!
0%
b11 *
0-
02
b11 6
#490150000000
1!
1%
1-
12
15
#490160000000
0!
0%
b100 *
0-
02
b100 6
#490170000000
1!
1%
1-
12
#490180000000
0!
0%
b101 *
0-
02
b101 6
#490190000000
1!
1%
1-
12
#490200000000
0!
0%
b110 *
0-
02
b110 6
#490210000000
1!
1%
1-
12
#490220000000
0!
0%
b111 *
0-
02
b111 6
#490230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#490240000000
0!
0%
b0 *
0-
02
b0 6
#490250000000
1!
1%
1-
12
#490260000000
0!
0%
b1 *
0-
02
b1 6
#490270000000
1!
1%
1-
12
#490280000000
0!
0%
b10 *
0-
02
b10 6
#490290000000
1!
1%
1-
12
#490300000000
0!
0%
b11 *
0-
02
b11 6
#490310000000
1!
1%
1-
12
15
#490320000000
0!
0%
b100 *
0-
02
b100 6
#490330000000
1!
1%
1-
12
#490340000000
0!
0%
b101 *
0-
02
b101 6
#490350000000
1!
1%
1-
12
#490360000000
0!
0%
b110 *
0-
02
b110 6
#490370000000
1!
1%
1-
12
#490380000000
0!
0%
b111 *
0-
02
b111 6
#490390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#490400000000
0!
0%
b0 *
0-
02
b0 6
#490410000000
1!
1%
1-
12
#490420000000
0!
0%
b1 *
0-
02
b1 6
#490430000000
1!
1%
1-
12
#490440000000
0!
0%
b10 *
0-
02
b10 6
#490450000000
1!
1%
1-
12
#490460000000
0!
0%
b11 *
0-
02
b11 6
#490470000000
1!
1%
1-
12
15
#490480000000
0!
0%
b100 *
0-
02
b100 6
#490490000000
1!
1%
1-
12
#490500000000
0!
0%
b101 *
0-
02
b101 6
#490510000000
1!
1%
1-
12
#490520000000
0!
0%
b110 *
0-
02
b110 6
#490530000000
1!
1%
1-
12
#490540000000
0!
0%
b111 *
0-
02
b111 6
#490550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#490560000000
0!
0%
b0 *
0-
02
b0 6
#490570000000
1!
1%
1-
12
#490580000000
0!
0%
b1 *
0-
02
b1 6
#490590000000
1!
1%
1-
12
#490600000000
0!
0%
b10 *
0-
02
b10 6
#490610000000
1!
1%
1-
12
#490620000000
0!
0%
b11 *
0-
02
b11 6
#490630000000
1!
1%
1-
12
15
#490640000000
0!
0%
b100 *
0-
02
b100 6
#490650000000
1!
1%
1-
12
#490660000000
0!
0%
b101 *
0-
02
b101 6
#490670000000
1!
1%
1-
12
#490680000000
0!
0%
b110 *
0-
02
b110 6
#490690000000
1!
1%
1-
12
#490700000000
0!
0%
b111 *
0-
02
b111 6
#490710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#490720000000
0!
0%
b0 *
0-
02
b0 6
#490730000000
1!
1%
1-
12
#490740000000
0!
0%
b1 *
0-
02
b1 6
#490750000000
1!
1%
1-
12
#490760000000
0!
0%
b10 *
0-
02
b10 6
#490770000000
1!
1%
1-
12
#490780000000
0!
0%
b11 *
0-
02
b11 6
#490790000000
1!
1%
1-
12
15
#490800000000
0!
0%
b100 *
0-
02
b100 6
#490810000000
1!
1%
1-
12
#490820000000
0!
0%
b101 *
0-
02
b101 6
#490830000000
1!
1%
1-
12
#490840000000
0!
0%
b110 *
0-
02
b110 6
#490850000000
1!
1%
1-
12
#490860000000
0!
0%
b111 *
0-
02
b111 6
#490870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#490880000000
0!
0%
b0 *
0-
02
b0 6
#490890000000
1!
1%
1-
12
#490900000000
0!
0%
b1 *
0-
02
b1 6
#490910000000
1!
1%
1-
12
#490920000000
0!
0%
b10 *
0-
02
b10 6
#490930000000
1!
1%
1-
12
#490940000000
0!
0%
b11 *
0-
02
b11 6
#490950000000
1!
1%
1-
12
15
#490960000000
0!
0%
b100 *
0-
02
b100 6
#490970000000
1!
1%
1-
12
#490980000000
0!
0%
b101 *
0-
02
b101 6
#490990000000
1!
1%
1-
12
#491000000000
0!
0%
b110 *
0-
02
b110 6
#491010000000
1!
1%
1-
12
#491020000000
0!
0%
b111 *
0-
02
b111 6
#491030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#491040000000
0!
0%
b0 *
0-
02
b0 6
#491050000000
1!
1%
1-
12
#491060000000
0!
0%
b1 *
0-
02
b1 6
#491070000000
1!
1%
1-
12
#491080000000
0!
0%
b10 *
0-
02
b10 6
#491090000000
1!
1%
1-
12
#491100000000
0!
0%
b11 *
0-
02
b11 6
#491110000000
1!
1%
1-
12
15
#491120000000
0!
0%
b100 *
0-
02
b100 6
#491130000000
1!
1%
1-
12
#491140000000
0!
0%
b101 *
0-
02
b101 6
#491150000000
1!
1%
1-
12
#491160000000
0!
0%
b110 *
0-
02
b110 6
#491170000000
1!
1%
1-
12
#491180000000
0!
0%
b111 *
0-
02
b111 6
#491190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#491200000000
0!
0%
b0 *
0-
02
b0 6
#491210000000
1!
1%
1-
12
#491220000000
0!
0%
b1 *
0-
02
b1 6
#491230000000
1!
1%
1-
12
#491240000000
0!
0%
b10 *
0-
02
b10 6
#491250000000
1!
1%
1-
12
#491260000000
0!
0%
b11 *
0-
02
b11 6
#491270000000
1!
1%
1-
12
15
#491280000000
0!
0%
b100 *
0-
02
b100 6
#491290000000
1!
1%
1-
12
#491300000000
0!
0%
b101 *
0-
02
b101 6
#491310000000
1!
1%
1-
12
#491320000000
0!
0%
b110 *
0-
02
b110 6
#491330000000
1!
1%
1-
12
#491340000000
0!
0%
b111 *
0-
02
b111 6
#491350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#491360000000
0!
0%
b0 *
0-
02
b0 6
#491370000000
1!
1%
1-
12
#491380000000
0!
0%
b1 *
0-
02
b1 6
#491390000000
1!
1%
1-
12
#491400000000
0!
0%
b10 *
0-
02
b10 6
#491410000000
1!
1%
1-
12
#491420000000
0!
0%
b11 *
0-
02
b11 6
#491430000000
1!
1%
1-
12
15
#491440000000
0!
0%
b100 *
0-
02
b100 6
#491450000000
1!
1%
1-
12
#491460000000
0!
0%
b101 *
0-
02
b101 6
#491470000000
1!
1%
1-
12
#491480000000
0!
0%
b110 *
0-
02
b110 6
#491490000000
1!
1%
1-
12
#491500000000
0!
0%
b111 *
0-
02
b111 6
#491510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#491520000000
0!
0%
b0 *
0-
02
b0 6
#491530000000
1!
1%
1-
12
#491540000000
0!
0%
b1 *
0-
02
b1 6
#491550000000
1!
1%
1-
12
#491560000000
0!
0%
b10 *
0-
02
b10 6
#491570000000
1!
1%
1-
12
#491580000000
0!
0%
b11 *
0-
02
b11 6
#491590000000
1!
1%
1-
12
15
#491600000000
0!
0%
b100 *
0-
02
b100 6
#491610000000
1!
1%
1-
12
#491620000000
0!
0%
b101 *
0-
02
b101 6
#491630000000
1!
1%
1-
12
#491640000000
0!
0%
b110 *
0-
02
b110 6
#491650000000
1!
1%
1-
12
#491660000000
0!
0%
b111 *
0-
02
b111 6
#491670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#491680000000
0!
0%
b0 *
0-
02
b0 6
#491690000000
1!
1%
1-
12
#491700000000
0!
0%
b1 *
0-
02
b1 6
#491710000000
1!
1%
1-
12
#491720000000
0!
0%
b10 *
0-
02
b10 6
#491730000000
1!
1%
1-
12
#491740000000
0!
0%
b11 *
0-
02
b11 6
#491750000000
1!
1%
1-
12
15
#491760000000
0!
0%
b100 *
0-
02
b100 6
#491770000000
1!
1%
1-
12
#491780000000
0!
0%
b101 *
0-
02
b101 6
#491790000000
1!
1%
1-
12
#491800000000
0!
0%
b110 *
0-
02
b110 6
#491810000000
1!
1%
1-
12
#491820000000
0!
0%
b111 *
0-
02
b111 6
#491830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#491840000000
0!
0%
b0 *
0-
02
b0 6
#491850000000
1!
1%
1-
12
#491860000000
0!
0%
b1 *
0-
02
b1 6
#491870000000
1!
1%
1-
12
#491880000000
0!
0%
b10 *
0-
02
b10 6
#491890000000
1!
1%
1-
12
#491900000000
0!
0%
b11 *
0-
02
b11 6
#491910000000
1!
1%
1-
12
15
#491920000000
0!
0%
b100 *
0-
02
b100 6
#491930000000
1!
1%
1-
12
#491940000000
0!
0%
b101 *
0-
02
b101 6
#491950000000
1!
1%
1-
12
#491960000000
0!
0%
b110 *
0-
02
b110 6
#491970000000
1!
1%
1-
12
#491980000000
0!
0%
b111 *
0-
02
b111 6
#491990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#492000000000
0!
0%
b0 *
0-
02
b0 6
#492010000000
1!
1%
1-
12
#492020000000
0!
0%
b1 *
0-
02
b1 6
#492030000000
1!
1%
1-
12
#492040000000
0!
0%
b10 *
0-
02
b10 6
#492050000000
1!
1%
1-
12
#492060000000
0!
0%
b11 *
0-
02
b11 6
#492070000000
1!
1%
1-
12
15
#492080000000
0!
0%
b100 *
0-
02
b100 6
#492090000000
1!
1%
1-
12
#492100000000
0!
0%
b101 *
0-
02
b101 6
#492110000000
1!
1%
1-
12
#492120000000
0!
0%
b110 *
0-
02
b110 6
#492130000000
1!
1%
1-
12
#492140000000
0!
0%
b111 *
0-
02
b111 6
#492150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#492160000000
0!
0%
b0 *
0-
02
b0 6
#492170000000
1!
1%
1-
12
#492180000000
0!
0%
b1 *
0-
02
b1 6
#492190000000
1!
1%
1-
12
#492200000000
0!
0%
b10 *
0-
02
b10 6
#492210000000
1!
1%
1-
12
#492220000000
0!
0%
b11 *
0-
02
b11 6
#492230000000
1!
1%
1-
12
15
#492240000000
0!
0%
b100 *
0-
02
b100 6
#492250000000
1!
1%
1-
12
#492260000000
0!
0%
b101 *
0-
02
b101 6
#492270000000
1!
1%
1-
12
#492280000000
0!
0%
b110 *
0-
02
b110 6
#492290000000
1!
1%
1-
12
#492300000000
0!
0%
b111 *
0-
02
b111 6
#492310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#492320000000
0!
0%
b0 *
0-
02
b0 6
#492330000000
1!
1%
1-
12
#492340000000
0!
0%
b1 *
0-
02
b1 6
#492350000000
1!
1%
1-
12
#492360000000
0!
0%
b10 *
0-
02
b10 6
#492370000000
1!
1%
1-
12
#492380000000
0!
0%
b11 *
0-
02
b11 6
#492390000000
1!
1%
1-
12
15
#492400000000
0!
0%
b100 *
0-
02
b100 6
#492410000000
1!
1%
1-
12
#492420000000
0!
0%
b101 *
0-
02
b101 6
#492430000000
1!
1%
1-
12
#492440000000
0!
0%
b110 *
0-
02
b110 6
#492450000000
1!
1%
1-
12
#492460000000
0!
0%
b111 *
0-
02
b111 6
#492470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#492480000000
0!
0%
b0 *
0-
02
b0 6
#492490000000
1!
1%
1-
12
#492500000000
0!
0%
b1 *
0-
02
b1 6
#492510000000
1!
1%
1-
12
#492520000000
0!
0%
b10 *
0-
02
b10 6
#492530000000
1!
1%
1-
12
#492540000000
0!
0%
b11 *
0-
02
b11 6
#492550000000
1!
1%
1-
12
15
#492560000000
0!
0%
b100 *
0-
02
b100 6
#492570000000
1!
1%
1-
12
#492580000000
0!
0%
b101 *
0-
02
b101 6
#492590000000
1!
1%
1-
12
#492600000000
0!
0%
b110 *
0-
02
b110 6
#492610000000
1!
1%
1-
12
#492620000000
0!
0%
b111 *
0-
02
b111 6
#492630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#492640000000
0!
0%
b0 *
0-
02
b0 6
#492650000000
1!
1%
1-
12
#492660000000
0!
0%
b1 *
0-
02
b1 6
#492670000000
1!
1%
1-
12
#492680000000
0!
0%
b10 *
0-
02
b10 6
#492690000000
1!
1%
1-
12
#492700000000
0!
0%
b11 *
0-
02
b11 6
#492710000000
1!
1%
1-
12
15
#492720000000
0!
0%
b100 *
0-
02
b100 6
#492730000000
1!
1%
1-
12
#492740000000
0!
0%
b101 *
0-
02
b101 6
#492750000000
1!
1%
1-
12
#492760000000
0!
0%
b110 *
0-
02
b110 6
#492770000000
1!
1%
1-
12
#492780000000
0!
0%
b111 *
0-
02
b111 6
#492790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#492800000000
0!
0%
b0 *
0-
02
b0 6
#492810000000
1!
1%
1-
12
#492820000000
0!
0%
b1 *
0-
02
b1 6
#492830000000
1!
1%
1-
12
#492840000000
0!
0%
b10 *
0-
02
b10 6
#492850000000
1!
1%
1-
12
#492860000000
0!
0%
b11 *
0-
02
b11 6
#492870000000
1!
1%
1-
12
15
#492880000000
0!
0%
b100 *
0-
02
b100 6
#492890000000
1!
1%
1-
12
#492900000000
0!
0%
b101 *
0-
02
b101 6
#492910000000
1!
1%
1-
12
#492920000000
0!
0%
b110 *
0-
02
b110 6
#492930000000
1!
1%
1-
12
#492940000000
0!
0%
b111 *
0-
02
b111 6
#492950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#492960000000
0!
0%
b0 *
0-
02
b0 6
#492970000000
1!
1%
1-
12
#492980000000
0!
0%
b1 *
0-
02
b1 6
#492990000000
1!
1%
1-
12
#493000000000
0!
0%
b10 *
0-
02
b10 6
#493010000000
1!
1%
1-
12
#493020000000
0!
0%
b11 *
0-
02
b11 6
#493030000000
1!
1%
1-
12
15
#493040000000
0!
0%
b100 *
0-
02
b100 6
#493050000000
1!
1%
1-
12
#493060000000
0!
0%
b101 *
0-
02
b101 6
#493070000000
1!
1%
1-
12
#493080000000
0!
0%
b110 *
0-
02
b110 6
#493090000000
1!
1%
1-
12
#493100000000
0!
0%
b111 *
0-
02
b111 6
#493110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#493120000000
0!
0%
b0 *
0-
02
b0 6
#493130000000
1!
1%
1-
12
#493140000000
0!
0%
b1 *
0-
02
b1 6
#493150000000
1!
1%
1-
12
#493160000000
0!
0%
b10 *
0-
02
b10 6
#493170000000
1!
1%
1-
12
#493180000000
0!
0%
b11 *
0-
02
b11 6
#493190000000
1!
1%
1-
12
15
#493200000000
0!
0%
b100 *
0-
02
b100 6
#493210000000
1!
1%
1-
12
#493220000000
0!
0%
b101 *
0-
02
b101 6
#493230000000
1!
1%
1-
12
#493240000000
0!
0%
b110 *
0-
02
b110 6
#493250000000
1!
1%
1-
12
#493260000000
0!
0%
b111 *
0-
02
b111 6
#493270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#493280000000
0!
0%
b0 *
0-
02
b0 6
#493290000000
1!
1%
1-
12
#493300000000
0!
0%
b1 *
0-
02
b1 6
#493310000000
1!
1%
1-
12
#493320000000
0!
0%
b10 *
0-
02
b10 6
#493330000000
1!
1%
1-
12
#493340000000
0!
0%
b11 *
0-
02
b11 6
#493350000000
1!
1%
1-
12
15
#493360000000
0!
0%
b100 *
0-
02
b100 6
#493370000000
1!
1%
1-
12
#493380000000
0!
0%
b101 *
0-
02
b101 6
#493390000000
1!
1%
1-
12
#493400000000
0!
0%
b110 *
0-
02
b110 6
#493410000000
1!
1%
1-
12
#493420000000
0!
0%
b111 *
0-
02
b111 6
#493430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#493440000000
0!
0%
b0 *
0-
02
b0 6
#493450000000
1!
1%
1-
12
#493460000000
0!
0%
b1 *
0-
02
b1 6
#493470000000
1!
1%
1-
12
#493480000000
0!
0%
b10 *
0-
02
b10 6
#493490000000
1!
1%
1-
12
#493500000000
0!
0%
b11 *
0-
02
b11 6
#493510000000
1!
1%
1-
12
15
#493520000000
0!
0%
b100 *
0-
02
b100 6
#493530000000
1!
1%
1-
12
#493540000000
0!
0%
b101 *
0-
02
b101 6
#493550000000
1!
1%
1-
12
#493560000000
0!
0%
b110 *
0-
02
b110 6
#493570000000
1!
1%
1-
12
#493580000000
0!
0%
b111 *
0-
02
b111 6
#493590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#493600000000
0!
0%
b0 *
0-
02
b0 6
#493610000000
1!
1%
1-
12
#493620000000
0!
0%
b1 *
0-
02
b1 6
#493630000000
1!
1%
1-
12
#493640000000
0!
0%
b10 *
0-
02
b10 6
#493650000000
1!
1%
1-
12
#493660000000
0!
0%
b11 *
0-
02
b11 6
#493670000000
1!
1%
1-
12
15
#493680000000
0!
0%
b100 *
0-
02
b100 6
#493690000000
1!
1%
1-
12
#493700000000
0!
0%
b101 *
0-
02
b101 6
#493710000000
1!
1%
1-
12
#493720000000
0!
0%
b110 *
0-
02
b110 6
#493730000000
1!
1%
1-
12
#493740000000
0!
0%
b111 *
0-
02
b111 6
#493750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#493760000000
0!
0%
b0 *
0-
02
b0 6
#493770000000
1!
1%
1-
12
#493780000000
0!
0%
b1 *
0-
02
b1 6
#493790000000
1!
1%
1-
12
#493800000000
0!
0%
b10 *
0-
02
b10 6
#493810000000
1!
1%
1-
12
#493820000000
0!
0%
b11 *
0-
02
b11 6
#493830000000
1!
1%
1-
12
15
#493840000000
0!
0%
b100 *
0-
02
b100 6
#493850000000
1!
1%
1-
12
#493860000000
0!
0%
b101 *
0-
02
b101 6
#493870000000
1!
1%
1-
12
#493880000000
0!
0%
b110 *
0-
02
b110 6
#493890000000
1!
1%
1-
12
#493900000000
0!
0%
b111 *
0-
02
b111 6
#493910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#493920000000
0!
0%
b0 *
0-
02
b0 6
#493930000000
1!
1%
1-
12
#493940000000
0!
0%
b1 *
0-
02
b1 6
#493950000000
1!
1%
1-
12
#493960000000
0!
0%
b10 *
0-
02
b10 6
#493970000000
1!
1%
1-
12
#493980000000
0!
0%
b11 *
0-
02
b11 6
#493990000000
1!
1%
1-
12
15
#494000000000
0!
0%
b100 *
0-
02
b100 6
#494010000000
1!
1%
1-
12
#494020000000
0!
0%
b101 *
0-
02
b101 6
#494030000000
1!
1%
1-
12
#494040000000
0!
0%
b110 *
0-
02
b110 6
#494050000000
1!
1%
1-
12
#494060000000
0!
0%
b111 *
0-
02
b111 6
#494070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#494080000000
0!
0%
b0 *
0-
02
b0 6
#494090000000
1!
1%
1-
12
#494100000000
0!
0%
b1 *
0-
02
b1 6
#494110000000
1!
1%
1-
12
#494120000000
0!
0%
b10 *
0-
02
b10 6
#494130000000
1!
1%
1-
12
#494140000000
0!
0%
b11 *
0-
02
b11 6
#494150000000
1!
1%
1-
12
15
#494160000000
0!
0%
b100 *
0-
02
b100 6
#494170000000
1!
1%
1-
12
#494180000000
0!
0%
b101 *
0-
02
b101 6
#494190000000
1!
1%
1-
12
#494200000000
0!
0%
b110 *
0-
02
b110 6
#494210000000
1!
1%
1-
12
#494220000000
0!
0%
b111 *
0-
02
b111 6
#494230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#494240000000
0!
0%
b0 *
0-
02
b0 6
#494250000000
1!
1%
1-
12
#494260000000
0!
0%
b1 *
0-
02
b1 6
#494270000000
1!
1%
1-
12
#494280000000
0!
0%
b10 *
0-
02
b10 6
#494290000000
1!
1%
1-
12
#494300000000
0!
0%
b11 *
0-
02
b11 6
#494310000000
1!
1%
1-
12
15
#494320000000
0!
0%
b100 *
0-
02
b100 6
#494330000000
1!
1%
1-
12
#494340000000
0!
0%
b101 *
0-
02
b101 6
#494350000000
1!
1%
1-
12
#494360000000
0!
0%
b110 *
0-
02
b110 6
#494370000000
1!
1%
1-
12
#494380000000
0!
0%
b111 *
0-
02
b111 6
#494390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#494400000000
0!
0%
b0 *
0-
02
b0 6
#494410000000
1!
1%
1-
12
#494420000000
0!
0%
b1 *
0-
02
b1 6
#494430000000
1!
1%
1-
12
#494440000000
0!
0%
b10 *
0-
02
b10 6
#494450000000
1!
1%
1-
12
#494460000000
0!
0%
b11 *
0-
02
b11 6
#494470000000
1!
1%
1-
12
15
#494480000000
0!
0%
b100 *
0-
02
b100 6
#494490000000
1!
1%
1-
12
#494500000000
0!
0%
b101 *
0-
02
b101 6
#494510000000
1!
1%
1-
12
#494520000000
0!
0%
b110 *
0-
02
b110 6
#494530000000
1!
1%
1-
12
#494540000000
0!
0%
b111 *
0-
02
b111 6
#494550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#494560000000
0!
0%
b0 *
0-
02
b0 6
#494570000000
1!
1%
1-
12
#494580000000
0!
0%
b1 *
0-
02
b1 6
#494590000000
1!
1%
1-
12
#494600000000
0!
0%
b10 *
0-
02
b10 6
#494610000000
1!
1%
1-
12
#494620000000
0!
0%
b11 *
0-
02
b11 6
#494630000000
1!
1%
1-
12
15
#494640000000
0!
0%
b100 *
0-
02
b100 6
#494650000000
1!
1%
1-
12
#494660000000
0!
0%
b101 *
0-
02
b101 6
#494670000000
1!
1%
1-
12
#494680000000
0!
0%
b110 *
0-
02
b110 6
#494690000000
1!
1%
1-
12
#494700000000
0!
0%
b111 *
0-
02
b111 6
#494710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#494720000000
0!
0%
b0 *
0-
02
b0 6
#494730000000
1!
1%
1-
12
#494740000000
0!
0%
b1 *
0-
02
b1 6
#494750000000
1!
1%
1-
12
#494760000000
0!
0%
b10 *
0-
02
b10 6
#494770000000
1!
1%
1-
12
#494780000000
0!
0%
b11 *
0-
02
b11 6
#494790000000
1!
1%
1-
12
15
#494800000000
0!
0%
b100 *
0-
02
b100 6
#494810000000
1!
1%
1-
12
#494820000000
0!
0%
b101 *
0-
02
b101 6
#494830000000
1!
1%
1-
12
#494840000000
0!
0%
b110 *
0-
02
b110 6
#494850000000
1!
1%
1-
12
#494860000000
0!
0%
b111 *
0-
02
b111 6
#494870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#494880000000
0!
0%
b0 *
0-
02
b0 6
#494890000000
1!
1%
1-
12
#494900000000
0!
0%
b1 *
0-
02
b1 6
#494910000000
1!
1%
1-
12
#494920000000
0!
0%
b10 *
0-
02
b10 6
#494930000000
1!
1%
1-
12
#494940000000
0!
0%
b11 *
0-
02
b11 6
#494950000000
1!
1%
1-
12
15
#494960000000
0!
0%
b100 *
0-
02
b100 6
#494970000000
1!
1%
1-
12
#494980000000
0!
0%
b101 *
0-
02
b101 6
#494990000000
1!
1%
1-
12
#495000000000
0!
0%
b110 *
0-
02
b110 6
#495010000000
1!
1%
1-
12
#495020000000
0!
0%
b111 *
0-
02
b111 6
#495030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#495040000000
0!
0%
b0 *
0-
02
b0 6
#495050000000
1!
1%
1-
12
#495060000000
0!
0%
b1 *
0-
02
b1 6
#495070000000
1!
1%
1-
12
#495080000000
0!
0%
b10 *
0-
02
b10 6
#495090000000
1!
1%
1-
12
#495100000000
0!
0%
b11 *
0-
02
b11 6
#495110000000
1!
1%
1-
12
15
#495120000000
0!
0%
b100 *
0-
02
b100 6
#495130000000
1!
1%
1-
12
#495140000000
0!
0%
b101 *
0-
02
b101 6
#495150000000
1!
1%
1-
12
#495160000000
0!
0%
b110 *
0-
02
b110 6
#495170000000
1!
1%
1-
12
#495180000000
0!
0%
b111 *
0-
02
b111 6
#495190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#495200000000
0!
0%
b0 *
0-
02
b0 6
#495210000000
1!
1%
1-
12
#495220000000
0!
0%
b1 *
0-
02
b1 6
#495230000000
1!
1%
1-
12
#495240000000
0!
0%
b10 *
0-
02
b10 6
#495250000000
1!
1%
1-
12
#495260000000
0!
0%
b11 *
0-
02
b11 6
#495270000000
1!
1%
1-
12
15
#495280000000
0!
0%
b100 *
0-
02
b100 6
#495290000000
1!
1%
1-
12
#495300000000
0!
0%
b101 *
0-
02
b101 6
#495310000000
1!
1%
1-
12
#495320000000
0!
0%
b110 *
0-
02
b110 6
#495330000000
1!
1%
1-
12
#495340000000
0!
0%
b111 *
0-
02
b111 6
#495350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#495360000000
0!
0%
b0 *
0-
02
b0 6
#495370000000
1!
1%
1-
12
#495380000000
0!
0%
b1 *
0-
02
b1 6
#495390000000
1!
1%
1-
12
#495400000000
0!
0%
b10 *
0-
02
b10 6
#495410000000
1!
1%
1-
12
#495420000000
0!
0%
b11 *
0-
02
b11 6
#495430000000
1!
1%
1-
12
15
#495440000000
0!
0%
b100 *
0-
02
b100 6
#495450000000
1!
1%
1-
12
#495460000000
0!
0%
b101 *
0-
02
b101 6
#495470000000
1!
1%
1-
12
#495480000000
0!
0%
b110 *
0-
02
b110 6
#495490000000
1!
1%
1-
12
#495500000000
0!
0%
b111 *
0-
02
b111 6
#495510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#495520000000
0!
0%
b0 *
0-
02
b0 6
#495530000000
1!
1%
1-
12
#495540000000
0!
0%
b1 *
0-
02
b1 6
#495550000000
1!
1%
1-
12
#495560000000
0!
0%
b10 *
0-
02
b10 6
#495570000000
1!
1%
1-
12
#495580000000
0!
0%
b11 *
0-
02
b11 6
#495590000000
1!
1%
1-
12
15
#495600000000
0!
0%
b100 *
0-
02
b100 6
#495610000000
1!
1%
1-
12
#495620000000
0!
0%
b101 *
0-
02
b101 6
#495630000000
1!
1%
1-
12
#495640000000
0!
0%
b110 *
0-
02
b110 6
#495650000000
1!
1%
1-
12
#495660000000
0!
0%
b111 *
0-
02
b111 6
#495670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#495680000000
0!
0%
b0 *
0-
02
b0 6
#495690000000
1!
1%
1-
12
#495700000000
0!
0%
b1 *
0-
02
b1 6
#495710000000
1!
1%
1-
12
#495720000000
0!
0%
b10 *
0-
02
b10 6
#495730000000
1!
1%
1-
12
#495740000000
0!
0%
b11 *
0-
02
b11 6
#495750000000
1!
1%
1-
12
15
#495760000000
0!
0%
b100 *
0-
02
b100 6
#495770000000
1!
1%
1-
12
#495780000000
0!
0%
b101 *
0-
02
b101 6
#495790000000
1!
1%
1-
12
#495800000000
0!
0%
b110 *
0-
02
b110 6
#495810000000
1!
1%
1-
12
#495820000000
0!
0%
b111 *
0-
02
b111 6
#495830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#495840000000
0!
0%
b0 *
0-
02
b0 6
#495850000000
1!
1%
1-
12
#495860000000
0!
0%
b1 *
0-
02
b1 6
#495870000000
1!
1%
1-
12
#495880000000
0!
0%
b10 *
0-
02
b10 6
#495890000000
1!
1%
1-
12
#495900000000
0!
0%
b11 *
0-
02
b11 6
#495910000000
1!
1%
1-
12
15
#495920000000
0!
0%
b100 *
0-
02
b100 6
#495930000000
1!
1%
1-
12
#495940000000
0!
0%
b101 *
0-
02
b101 6
#495950000000
1!
1%
1-
12
#495960000000
0!
0%
b110 *
0-
02
b110 6
#495970000000
1!
1%
1-
12
#495980000000
0!
0%
b111 *
0-
02
b111 6
#495990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#496000000000
0!
0%
b0 *
0-
02
b0 6
#496010000000
1!
1%
1-
12
#496020000000
0!
0%
b1 *
0-
02
b1 6
#496030000000
1!
1%
1-
12
#496040000000
0!
0%
b10 *
0-
02
b10 6
#496050000000
1!
1%
1-
12
#496060000000
0!
0%
b11 *
0-
02
b11 6
#496070000000
1!
1%
1-
12
15
#496080000000
0!
0%
b100 *
0-
02
b100 6
#496090000000
1!
1%
1-
12
#496100000000
0!
0%
b101 *
0-
02
b101 6
#496110000000
1!
1%
1-
12
#496120000000
0!
0%
b110 *
0-
02
b110 6
#496130000000
1!
1%
1-
12
#496140000000
0!
0%
b111 *
0-
02
b111 6
#496150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#496160000000
0!
0%
b0 *
0-
02
b0 6
#496170000000
1!
1%
1-
12
#496180000000
0!
0%
b1 *
0-
02
b1 6
#496190000000
1!
1%
1-
12
#496200000000
0!
0%
b10 *
0-
02
b10 6
#496210000000
1!
1%
1-
12
#496220000000
0!
0%
b11 *
0-
02
b11 6
#496230000000
1!
1%
1-
12
15
#496240000000
0!
0%
b100 *
0-
02
b100 6
#496250000000
1!
1%
1-
12
#496260000000
0!
0%
b101 *
0-
02
b101 6
#496270000000
1!
1%
1-
12
#496280000000
0!
0%
b110 *
0-
02
b110 6
#496290000000
1!
1%
1-
12
#496300000000
0!
0%
b111 *
0-
02
b111 6
#496310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#496320000000
0!
0%
b0 *
0-
02
b0 6
#496330000000
1!
1%
1-
12
#496340000000
0!
0%
b1 *
0-
02
b1 6
#496350000000
1!
1%
1-
12
#496360000000
0!
0%
b10 *
0-
02
b10 6
#496370000000
1!
1%
1-
12
#496380000000
0!
0%
b11 *
0-
02
b11 6
#496390000000
1!
1%
1-
12
15
#496400000000
0!
0%
b100 *
0-
02
b100 6
#496410000000
1!
1%
1-
12
#496420000000
0!
0%
b101 *
0-
02
b101 6
#496430000000
1!
1%
1-
12
#496440000000
0!
0%
b110 *
0-
02
b110 6
#496450000000
1!
1%
1-
12
#496460000000
0!
0%
b111 *
0-
02
b111 6
#496470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#496480000000
0!
0%
b0 *
0-
02
b0 6
#496490000000
1!
1%
1-
12
#496500000000
0!
0%
b1 *
0-
02
b1 6
#496510000000
1!
1%
1-
12
#496520000000
0!
0%
b10 *
0-
02
b10 6
#496530000000
1!
1%
1-
12
#496540000000
0!
0%
b11 *
0-
02
b11 6
#496550000000
1!
1%
1-
12
15
#496560000000
0!
0%
b100 *
0-
02
b100 6
#496570000000
1!
1%
1-
12
#496580000000
0!
0%
b101 *
0-
02
b101 6
#496590000000
1!
1%
1-
12
#496600000000
0!
0%
b110 *
0-
02
b110 6
#496610000000
1!
1%
1-
12
#496620000000
0!
0%
b111 *
0-
02
b111 6
#496630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#496640000000
0!
0%
b0 *
0-
02
b0 6
#496650000000
1!
1%
1-
12
#496660000000
0!
0%
b1 *
0-
02
b1 6
#496670000000
1!
1%
1-
12
#496680000000
0!
0%
b10 *
0-
02
b10 6
#496690000000
1!
1%
1-
12
#496700000000
0!
0%
b11 *
0-
02
b11 6
#496710000000
1!
1%
1-
12
15
#496720000000
0!
0%
b100 *
0-
02
b100 6
#496730000000
1!
1%
1-
12
#496740000000
0!
0%
b101 *
0-
02
b101 6
#496750000000
1!
1%
1-
12
#496760000000
0!
0%
b110 *
0-
02
b110 6
#496770000000
1!
1%
1-
12
#496780000000
0!
0%
b111 *
0-
02
b111 6
#496790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#496800000000
0!
0%
b0 *
0-
02
b0 6
#496810000000
1!
1%
1-
12
#496820000000
0!
0%
b1 *
0-
02
b1 6
#496830000000
1!
1%
1-
12
#496840000000
0!
0%
b10 *
0-
02
b10 6
#496850000000
1!
1%
1-
12
#496860000000
0!
0%
b11 *
0-
02
b11 6
#496870000000
1!
1%
1-
12
15
#496880000000
0!
0%
b100 *
0-
02
b100 6
#496890000000
1!
1%
1-
12
#496900000000
0!
0%
b101 *
0-
02
b101 6
#496910000000
1!
1%
1-
12
#496920000000
0!
0%
b110 *
0-
02
b110 6
#496930000000
1!
1%
1-
12
#496940000000
0!
0%
b111 *
0-
02
b111 6
#496950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#496960000000
0!
0%
b0 *
0-
02
b0 6
#496970000000
1!
1%
1-
12
#496980000000
0!
0%
b1 *
0-
02
b1 6
#496990000000
1!
1%
1-
12
#497000000000
0!
0%
b10 *
0-
02
b10 6
#497010000000
1!
1%
1-
12
#497020000000
0!
0%
b11 *
0-
02
b11 6
#497030000000
1!
1%
1-
12
15
#497040000000
0!
0%
b100 *
0-
02
b100 6
#497050000000
1!
1%
1-
12
#497060000000
0!
0%
b101 *
0-
02
b101 6
#497070000000
1!
1%
1-
12
#497080000000
0!
0%
b110 *
0-
02
b110 6
#497090000000
1!
1%
1-
12
#497100000000
0!
0%
b111 *
0-
02
b111 6
#497110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#497120000000
0!
0%
b0 *
0-
02
b0 6
#497130000000
1!
1%
1-
12
#497140000000
0!
0%
b1 *
0-
02
b1 6
#497150000000
1!
1%
1-
12
#497160000000
0!
0%
b10 *
0-
02
b10 6
#497170000000
1!
1%
1-
12
#497180000000
0!
0%
b11 *
0-
02
b11 6
#497190000000
1!
1%
1-
12
15
#497200000000
0!
0%
b100 *
0-
02
b100 6
#497210000000
1!
1%
1-
12
#497220000000
0!
0%
b101 *
0-
02
b101 6
#497230000000
1!
1%
1-
12
#497240000000
0!
0%
b110 *
0-
02
b110 6
#497250000000
1!
1%
1-
12
#497260000000
0!
0%
b111 *
0-
02
b111 6
#497270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#497280000000
0!
0%
b0 *
0-
02
b0 6
#497290000000
1!
1%
1-
12
#497300000000
0!
0%
b1 *
0-
02
b1 6
#497310000000
1!
1%
1-
12
#497320000000
0!
0%
b10 *
0-
02
b10 6
#497330000000
1!
1%
1-
12
#497340000000
0!
0%
b11 *
0-
02
b11 6
#497350000000
1!
1%
1-
12
15
#497360000000
0!
0%
b100 *
0-
02
b100 6
#497370000000
1!
1%
1-
12
#497380000000
0!
0%
b101 *
0-
02
b101 6
#497390000000
1!
1%
1-
12
#497400000000
0!
0%
b110 *
0-
02
b110 6
#497410000000
1!
1%
1-
12
#497420000000
0!
0%
b111 *
0-
02
b111 6
#497430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#497440000000
0!
0%
b0 *
0-
02
b0 6
#497450000000
1!
1%
1-
12
#497460000000
0!
0%
b1 *
0-
02
b1 6
#497470000000
1!
1%
1-
12
#497480000000
0!
0%
b10 *
0-
02
b10 6
#497490000000
1!
1%
1-
12
#497500000000
0!
0%
b11 *
0-
02
b11 6
#497510000000
1!
1%
1-
12
15
#497520000000
0!
0%
b100 *
0-
02
b100 6
#497530000000
1!
1%
1-
12
#497540000000
0!
0%
b101 *
0-
02
b101 6
#497550000000
1!
1%
1-
12
#497560000000
0!
0%
b110 *
0-
02
b110 6
#497570000000
1!
1%
1-
12
#497580000000
0!
0%
b111 *
0-
02
b111 6
#497590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#497600000000
0!
0%
b0 *
0-
02
b0 6
#497610000000
1!
1%
1-
12
#497620000000
0!
0%
b1 *
0-
02
b1 6
#497630000000
1!
1%
1-
12
#497640000000
0!
0%
b10 *
0-
02
b10 6
#497650000000
1!
1%
1-
12
#497660000000
0!
0%
b11 *
0-
02
b11 6
#497670000000
1!
1%
1-
12
15
#497680000000
0!
0%
b100 *
0-
02
b100 6
#497690000000
1!
1%
1-
12
#497700000000
0!
0%
b101 *
0-
02
b101 6
#497710000000
1!
1%
1-
12
#497720000000
0!
0%
b110 *
0-
02
b110 6
#497730000000
1!
1%
1-
12
#497740000000
0!
0%
b111 *
0-
02
b111 6
#497750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#497760000000
0!
0%
b0 *
0-
02
b0 6
#497770000000
1!
1%
1-
12
#497780000000
0!
0%
b1 *
0-
02
b1 6
#497790000000
1!
1%
1-
12
#497800000000
0!
0%
b10 *
0-
02
b10 6
#497810000000
1!
1%
1-
12
#497820000000
0!
0%
b11 *
0-
02
b11 6
#497830000000
1!
1%
1-
12
15
#497840000000
0!
0%
b100 *
0-
02
b100 6
#497850000000
1!
1%
1-
12
#497860000000
0!
0%
b101 *
0-
02
b101 6
#497870000000
1!
1%
1-
12
#497880000000
0!
0%
b110 *
0-
02
b110 6
#497890000000
1!
1%
1-
12
#497900000000
0!
0%
b111 *
0-
02
b111 6
#497910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#497920000000
0!
0%
b0 *
0-
02
b0 6
#497930000000
1!
1%
1-
12
#497940000000
0!
0%
b1 *
0-
02
b1 6
#497950000000
1!
1%
1-
12
#497960000000
0!
0%
b10 *
0-
02
b10 6
#497970000000
1!
1%
1-
12
#497980000000
0!
0%
b11 *
0-
02
b11 6
#497990000000
1!
1%
1-
12
15
#498000000000
0!
0%
b100 *
0-
02
b100 6
#498010000000
1!
1%
1-
12
#498020000000
0!
0%
b101 *
0-
02
b101 6
#498030000000
1!
1%
1-
12
#498040000000
0!
0%
b110 *
0-
02
b110 6
#498050000000
1!
1%
1-
12
#498060000000
0!
0%
b111 *
0-
02
b111 6
#498070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#498080000000
0!
0%
b0 *
0-
02
b0 6
#498090000000
1!
1%
1-
12
#498100000000
0!
0%
b1 *
0-
02
b1 6
#498110000000
1!
1%
1-
12
#498120000000
0!
0%
b10 *
0-
02
b10 6
#498130000000
1!
1%
1-
12
#498140000000
0!
0%
b11 *
0-
02
b11 6
#498150000000
1!
1%
1-
12
15
#498160000000
0!
0%
b100 *
0-
02
b100 6
#498170000000
1!
1%
1-
12
#498180000000
0!
0%
b101 *
0-
02
b101 6
#498190000000
1!
1%
1-
12
#498200000000
0!
0%
b110 *
0-
02
b110 6
#498210000000
1!
1%
1-
12
#498220000000
0!
0%
b111 *
0-
02
b111 6
#498230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#498240000000
0!
0%
b0 *
0-
02
b0 6
#498250000000
1!
1%
1-
12
#498260000000
0!
0%
b1 *
0-
02
b1 6
#498270000000
1!
1%
1-
12
#498280000000
0!
0%
b10 *
0-
02
b10 6
#498290000000
1!
1%
1-
12
#498300000000
0!
0%
b11 *
0-
02
b11 6
#498310000000
1!
1%
1-
12
15
#498320000000
0!
0%
b100 *
0-
02
b100 6
#498330000000
1!
1%
1-
12
#498340000000
0!
0%
b101 *
0-
02
b101 6
#498350000000
1!
1%
1-
12
#498360000000
0!
0%
b110 *
0-
02
b110 6
#498370000000
1!
1%
1-
12
#498380000000
0!
0%
b111 *
0-
02
b111 6
#498390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#498400000000
0!
0%
b0 *
0-
02
b0 6
#498410000000
1!
1%
1-
12
#498420000000
0!
0%
b1 *
0-
02
b1 6
#498430000000
1!
1%
1-
12
#498440000000
0!
0%
b10 *
0-
02
b10 6
#498450000000
1!
1%
1-
12
#498460000000
0!
0%
b11 *
0-
02
b11 6
#498470000000
1!
1%
1-
12
15
#498480000000
0!
0%
b100 *
0-
02
b100 6
#498490000000
1!
1%
1-
12
#498500000000
0!
0%
b101 *
0-
02
b101 6
#498510000000
1!
1%
1-
12
#498520000000
0!
0%
b110 *
0-
02
b110 6
#498530000000
1!
1%
1-
12
#498540000000
0!
0%
b111 *
0-
02
b111 6
#498550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#498560000000
0!
0%
b0 *
0-
02
b0 6
#498570000000
1!
1%
1-
12
#498580000000
0!
0%
b1 *
0-
02
b1 6
#498590000000
1!
1%
1-
12
#498600000000
0!
0%
b10 *
0-
02
b10 6
#498610000000
1!
1%
1-
12
#498620000000
0!
0%
b11 *
0-
02
b11 6
#498630000000
1!
1%
1-
12
15
#498640000000
0!
0%
b100 *
0-
02
b100 6
#498650000000
1!
1%
1-
12
#498660000000
0!
0%
b101 *
0-
02
b101 6
#498670000000
1!
1%
1-
12
#498680000000
0!
0%
b110 *
0-
02
b110 6
#498690000000
1!
1%
1-
12
#498700000000
0!
0%
b111 *
0-
02
b111 6
#498710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#498720000000
0!
0%
b0 *
0-
02
b0 6
#498730000000
1!
1%
1-
12
#498740000000
0!
0%
b1 *
0-
02
b1 6
#498750000000
1!
1%
1-
12
#498760000000
0!
0%
b10 *
0-
02
b10 6
#498770000000
1!
1%
1-
12
#498780000000
0!
0%
b11 *
0-
02
b11 6
#498790000000
1!
1%
1-
12
15
#498800000000
0!
0%
b100 *
0-
02
b100 6
#498810000000
1!
1%
1-
12
#498820000000
0!
0%
b101 *
0-
02
b101 6
#498830000000
1!
1%
1-
12
#498840000000
0!
0%
b110 *
0-
02
b110 6
#498850000000
1!
1%
1-
12
#498860000000
0!
0%
b111 *
0-
02
b111 6
#498870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#498880000000
0!
0%
b0 *
0-
02
b0 6
#498890000000
1!
1%
1-
12
#498900000000
0!
0%
b1 *
0-
02
b1 6
#498910000000
1!
1%
1-
12
#498920000000
0!
0%
b10 *
0-
02
b10 6
#498930000000
1!
1%
1-
12
#498940000000
0!
0%
b11 *
0-
02
b11 6
#498950000000
1!
1%
1-
12
15
#498960000000
0!
0%
b100 *
0-
02
b100 6
#498970000000
1!
1%
1-
12
#498980000000
0!
0%
b101 *
0-
02
b101 6
#498990000000
1!
1%
1-
12
#499000000000
0!
0%
b110 *
0-
02
b110 6
#499010000000
1!
1%
1-
12
#499020000000
0!
0%
b111 *
0-
02
b111 6
#499030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#499040000000
0!
0%
b0 *
0-
02
b0 6
#499050000000
1!
1%
1-
12
#499060000000
0!
0%
b1 *
0-
02
b1 6
#499070000000
1!
1%
1-
12
#499080000000
0!
0%
b10 *
0-
02
b10 6
#499090000000
1!
1%
1-
12
#499100000000
0!
0%
b11 *
0-
02
b11 6
#499110000000
1!
1%
1-
12
15
#499120000000
0!
0%
b100 *
0-
02
b100 6
#499130000000
1!
1%
1-
12
#499140000000
0!
0%
b101 *
0-
02
b101 6
#499150000000
1!
1%
1-
12
#499160000000
0!
0%
b110 *
0-
02
b110 6
#499170000000
1!
1%
1-
12
#499180000000
0!
0%
b111 *
0-
02
b111 6
#499190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#499200000000
0!
0%
b0 *
0-
02
b0 6
#499210000000
1!
1%
1-
12
#499220000000
0!
0%
b1 *
0-
02
b1 6
#499230000000
1!
1%
1-
12
#499240000000
0!
0%
b10 *
0-
02
b10 6
#499250000000
1!
1%
1-
12
#499260000000
0!
0%
b11 *
0-
02
b11 6
#499270000000
1!
1%
1-
12
15
#499280000000
0!
0%
b100 *
0-
02
b100 6
#499290000000
1!
1%
1-
12
#499300000000
0!
0%
b101 *
0-
02
b101 6
#499310000000
1!
1%
1-
12
#499320000000
0!
0%
b110 *
0-
02
b110 6
#499330000000
1!
1%
1-
12
#499340000000
0!
0%
b111 *
0-
02
b111 6
#499350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#499360000000
0!
0%
b0 *
0-
02
b0 6
#499370000000
1!
1%
1-
12
#499380000000
0!
0%
b1 *
0-
02
b1 6
#499390000000
1!
1%
1-
12
#499400000000
0!
0%
b10 *
0-
02
b10 6
#499410000000
1!
1%
1-
12
#499420000000
0!
0%
b11 *
0-
02
b11 6
#499430000000
1!
1%
1-
12
15
#499440000000
0!
0%
b100 *
0-
02
b100 6
#499450000000
1!
1%
1-
12
#499460000000
0!
0%
b101 *
0-
02
b101 6
#499470000000
1!
1%
1-
12
#499480000000
0!
0%
b110 *
0-
02
b110 6
#499490000000
1!
1%
1-
12
#499500000000
0!
0%
b111 *
0-
02
b111 6
#499510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#499520000000
0!
0%
b0 *
0-
02
b0 6
#499530000000
1!
1%
1-
12
#499540000000
0!
0%
b1 *
0-
02
b1 6
#499550000000
1!
1%
1-
12
#499560000000
0!
0%
b10 *
0-
02
b10 6
#499570000000
1!
1%
1-
12
#499580000000
0!
0%
b11 *
0-
02
b11 6
#499590000000
1!
1%
1-
12
15
#499600000000
0!
0%
b100 *
0-
02
b100 6
#499610000000
1!
1%
1-
12
#499620000000
0!
0%
b101 *
0-
02
b101 6
#499630000000
1!
1%
1-
12
#499640000000
0!
0%
b110 *
0-
02
b110 6
#499650000000
1!
1%
1-
12
#499660000000
0!
0%
b111 *
0-
02
b111 6
#499670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#499680000000
0!
0%
b0 *
0-
02
b0 6
#499690000000
1!
1%
1-
12
#499700000000
0!
0%
b1 *
0-
02
b1 6
#499710000000
1!
1%
1-
12
#499720000000
0!
0%
b10 *
0-
02
b10 6
#499730000000
1!
1%
1-
12
#499740000000
0!
0%
b11 *
0-
02
b11 6
#499750000000
1!
1%
1-
12
15
#499760000000
0!
0%
b100 *
0-
02
b100 6
#499770000000
1!
1%
1-
12
#499780000000
0!
0%
b101 *
0-
02
b101 6
#499790000000
1!
1%
1-
12
#499800000000
0!
0%
b110 *
0-
02
b110 6
#499810000000
1!
1%
1-
12
#499820000000
0!
0%
b111 *
0-
02
b111 6
#499830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#499840000000
0!
0%
b0 *
0-
02
b0 6
#499850000000
1!
1%
1-
12
#499860000000
0!
0%
b1 *
0-
02
b1 6
#499870000000
1!
1%
1-
12
#499880000000
0!
0%
b10 *
0-
02
b10 6
#499890000000
1!
1%
1-
12
#499900000000
0!
0%
b11 *
0-
02
b11 6
#499910000000
1!
1%
1-
12
15
#499920000000
0!
0%
b100 *
0-
02
b100 6
#499930000000
1!
1%
1-
12
#499940000000
0!
0%
b101 *
0-
02
b101 6
#499950000000
1!
1%
1-
12
#499960000000
0!
0%
b110 *
0-
02
b110 6
#499970000000
1!
1%
1-
12
#499980000000
0!
0%
b111 *
0-
02
b111 6
#499990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#500000000000
0!
0%
b0 *
0-
02
b0 6
#500010000000
1!
1%
1-
12
#500020000000
0!
0%
b1 *
0-
02
b1 6
#500030000000
1!
1%
1-
12
#500040000000
0!
0%
b10 *
0-
02
b10 6
#500050000000
1!
1%
1-
12
#500060000000
0!
0%
b11 *
0-
02
b11 6
#500070000000
1!
1%
1-
12
15
#500080000000
0!
0%
b100 *
0-
02
b100 6
#500090000000
1!
1%
1-
12
#500100000000
0!
0%
b101 *
0-
02
b101 6
#500110000000
1!
1%
1-
12
#500120000000
0!
0%
b110 *
0-
02
b110 6
#500130000000
1!
1%
1-
12
#500140000000
0!
0%
b111 *
0-
02
b111 6
#500150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#500160000000
0!
0%
b0 *
0-
02
b0 6
#500170000000
1!
1%
1-
12
#500180000000
0!
0%
b1 *
0-
02
b1 6
#500190000000
1!
1%
1-
12
#500200000000
0!
0%
b10 *
0-
02
b10 6
#500210000000
1!
1%
1-
12
#500220000000
0!
0%
b11 *
0-
02
b11 6
#500230000000
1!
1%
1-
12
15
#500240000000
0!
0%
b100 *
0-
02
b100 6
#500250000000
1!
1%
1-
12
#500260000000
0!
0%
b101 *
0-
02
b101 6
#500270000000
1!
1%
1-
12
#500280000000
0!
0%
b110 *
0-
02
b110 6
#500290000000
1!
1%
1-
12
#500300000000
0!
0%
b111 *
0-
02
b111 6
#500310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#500320000000
0!
0%
b0 *
0-
02
b0 6
#500330000000
1!
1%
1-
12
#500340000000
0!
0%
b1 *
0-
02
b1 6
#500350000000
1!
1%
1-
12
#500360000000
0!
0%
b10 *
0-
02
b10 6
#500370000000
1!
1%
1-
12
#500380000000
0!
0%
b11 *
0-
02
b11 6
#500390000000
1!
1%
1-
12
15
#500400000000
0!
0%
b100 *
0-
02
b100 6
#500410000000
1!
1%
1-
12
#500420000000
0!
0%
b101 *
0-
02
b101 6
#500430000000
1!
1%
1-
12
#500440000000
0!
0%
b110 *
0-
02
b110 6
#500450000000
1!
1%
1-
12
#500460000000
0!
0%
b111 *
0-
02
b111 6
#500470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#500480000000
0!
0%
b0 *
0-
02
b0 6
#500490000000
1!
1%
1-
12
#500500000000
0!
0%
b1 *
0-
02
b1 6
#500510000000
1!
1%
1-
12
#500520000000
0!
0%
b10 *
0-
02
b10 6
#500530000000
1!
1%
1-
12
#500540000000
0!
0%
b11 *
0-
02
b11 6
#500550000000
1!
1%
1-
12
15
#500560000000
0!
0%
b100 *
0-
02
b100 6
#500570000000
1!
1%
1-
12
#500580000000
0!
0%
b101 *
0-
02
b101 6
#500590000000
1!
1%
1-
12
#500600000000
0!
0%
b110 *
0-
02
b110 6
#500610000000
1!
1%
1-
12
#500620000000
0!
0%
b111 *
0-
02
b111 6
#500630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#500640000000
0!
0%
b0 *
0-
02
b0 6
#500650000000
1!
1%
1-
12
#500660000000
0!
0%
b1 *
0-
02
b1 6
#500670000000
1!
1%
1-
12
#500680000000
0!
0%
b10 *
0-
02
b10 6
#500690000000
1!
1%
1-
12
#500700000000
0!
0%
b11 *
0-
02
b11 6
#500710000000
1!
1%
1-
12
15
#500720000000
0!
0%
b100 *
0-
02
b100 6
#500730000000
1!
1%
1-
12
#500740000000
0!
0%
b101 *
0-
02
b101 6
#500750000000
1!
1%
1-
12
#500760000000
0!
0%
b110 *
0-
02
b110 6
#500770000000
1!
1%
1-
12
#500780000000
0!
0%
b111 *
0-
02
b111 6
#500790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#500800000000
0!
0%
b0 *
0-
02
b0 6
#500810000000
1!
1%
1-
12
#500820000000
0!
0%
b1 *
0-
02
b1 6
#500830000000
1!
1%
1-
12
#500840000000
0!
0%
b10 *
0-
02
b10 6
#500850000000
1!
1%
1-
12
#500860000000
0!
0%
b11 *
0-
02
b11 6
#500870000000
1!
1%
1-
12
15
#500880000000
0!
0%
b100 *
0-
02
b100 6
#500890000000
1!
1%
1-
12
#500900000000
0!
0%
b101 *
0-
02
b101 6
#500910000000
1!
1%
1-
12
#500920000000
0!
0%
b110 *
0-
02
b110 6
#500930000000
1!
1%
1-
12
#500940000000
0!
0%
b111 *
0-
02
b111 6
#500950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#500960000000
0!
0%
b0 *
0-
02
b0 6
#500970000000
1!
1%
1-
12
#500980000000
0!
0%
b1 *
0-
02
b1 6
#500990000000
1!
1%
1-
12
#501000000000
0!
0%
b10 *
0-
02
b10 6
#501010000000
1!
1%
1-
12
#501020000000
0!
0%
b11 *
0-
02
b11 6
#501030000000
1!
1%
1-
12
15
#501040000000
0!
0%
b100 *
0-
02
b100 6
#501050000000
1!
1%
1-
12
#501060000000
0!
0%
b101 *
0-
02
b101 6
#501070000000
1!
1%
1-
12
#501080000000
0!
0%
b110 *
0-
02
b110 6
#501090000000
1!
1%
1-
12
#501100000000
0!
0%
b111 *
0-
02
b111 6
#501110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#501120000000
0!
0%
b0 *
0-
02
b0 6
#501130000000
1!
1%
1-
12
#501140000000
0!
0%
b1 *
0-
02
b1 6
#501150000000
1!
1%
1-
12
#501160000000
0!
0%
b10 *
0-
02
b10 6
#501170000000
1!
1%
1-
12
#501180000000
0!
0%
b11 *
0-
02
b11 6
#501190000000
1!
1%
1-
12
15
#501200000000
0!
0%
b100 *
0-
02
b100 6
#501210000000
1!
1%
1-
12
#501220000000
0!
0%
b101 *
0-
02
b101 6
#501230000000
1!
1%
1-
12
#501240000000
0!
0%
b110 *
0-
02
b110 6
#501250000000
1!
1%
1-
12
#501260000000
0!
0%
b111 *
0-
02
b111 6
#501270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#501280000000
0!
0%
b0 *
0-
02
b0 6
#501290000000
1!
1%
1-
12
#501300000000
0!
0%
b1 *
0-
02
b1 6
#501310000000
1!
1%
1-
12
#501320000000
0!
0%
b10 *
0-
02
b10 6
#501330000000
1!
1%
1-
12
#501340000000
0!
0%
b11 *
0-
02
b11 6
#501350000000
1!
1%
1-
12
15
#501360000000
0!
0%
b100 *
0-
02
b100 6
#501370000000
1!
1%
1-
12
#501380000000
0!
0%
b101 *
0-
02
b101 6
#501390000000
1!
1%
1-
12
#501400000000
0!
0%
b110 *
0-
02
b110 6
#501410000000
1!
1%
1-
12
#501420000000
0!
0%
b111 *
0-
02
b111 6
#501430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#501440000000
0!
0%
b0 *
0-
02
b0 6
#501450000000
1!
1%
1-
12
#501460000000
0!
0%
b1 *
0-
02
b1 6
#501470000000
1!
1%
1-
12
#501480000000
0!
0%
b10 *
0-
02
b10 6
#501490000000
1!
1%
1-
12
#501500000000
0!
0%
b11 *
0-
02
b11 6
#501510000000
1!
1%
1-
12
15
#501520000000
0!
0%
b100 *
0-
02
b100 6
#501530000000
1!
1%
1-
12
#501540000000
0!
0%
b101 *
0-
02
b101 6
#501550000000
1!
1%
1-
12
#501560000000
0!
0%
b110 *
0-
02
b110 6
#501570000000
1!
1%
1-
12
#501580000000
0!
0%
b111 *
0-
02
b111 6
#501590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#501600000000
0!
0%
b0 *
0-
02
b0 6
#501610000000
1!
1%
1-
12
#501620000000
0!
0%
b1 *
0-
02
b1 6
#501630000000
1!
1%
1-
12
#501640000000
0!
0%
b10 *
0-
02
b10 6
#501650000000
1!
1%
1-
12
#501660000000
0!
0%
b11 *
0-
02
b11 6
#501670000000
1!
1%
1-
12
15
#501680000000
0!
0%
b100 *
0-
02
b100 6
#501690000000
1!
1%
1-
12
#501700000000
0!
0%
b101 *
0-
02
b101 6
#501710000000
1!
1%
1-
12
#501720000000
0!
0%
b110 *
0-
02
b110 6
#501730000000
1!
1%
1-
12
#501740000000
0!
0%
b111 *
0-
02
b111 6
#501750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#501760000000
0!
0%
b0 *
0-
02
b0 6
#501770000000
1!
1%
1-
12
#501780000000
0!
0%
b1 *
0-
02
b1 6
#501790000000
1!
1%
1-
12
#501800000000
0!
0%
b10 *
0-
02
b10 6
#501810000000
1!
1%
1-
12
#501820000000
0!
0%
b11 *
0-
02
b11 6
#501830000000
1!
1%
1-
12
15
#501840000000
0!
0%
b100 *
0-
02
b100 6
#501850000000
1!
1%
1-
12
#501860000000
0!
0%
b101 *
0-
02
b101 6
#501870000000
1!
1%
1-
12
#501880000000
0!
0%
b110 *
0-
02
b110 6
#501890000000
1!
1%
1-
12
#501900000000
0!
0%
b111 *
0-
02
b111 6
#501910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#501920000000
0!
0%
b0 *
0-
02
b0 6
#501930000000
1!
1%
1-
12
#501940000000
0!
0%
b1 *
0-
02
b1 6
#501950000000
1!
1%
1-
12
#501960000000
0!
0%
b10 *
0-
02
b10 6
#501970000000
1!
1%
1-
12
#501980000000
0!
0%
b11 *
0-
02
b11 6
#501990000000
1!
1%
1-
12
15
#502000000000
0!
0%
b100 *
0-
02
b100 6
#502010000000
1!
1%
1-
12
#502020000000
0!
0%
b101 *
0-
02
b101 6
#502030000000
1!
1%
1-
12
#502040000000
0!
0%
b110 *
0-
02
b110 6
#502050000000
1!
1%
1-
12
#502060000000
0!
0%
b111 *
0-
02
b111 6
#502070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#502080000000
0!
0%
b0 *
0-
02
b0 6
#502090000000
1!
1%
1-
12
#502100000000
0!
0%
b1 *
0-
02
b1 6
#502110000000
1!
1%
1-
12
#502120000000
0!
0%
b10 *
0-
02
b10 6
#502130000000
1!
1%
1-
12
#502140000000
0!
0%
b11 *
0-
02
b11 6
#502150000000
1!
1%
1-
12
15
#502160000000
0!
0%
b100 *
0-
02
b100 6
#502170000000
1!
1%
1-
12
#502180000000
0!
0%
b101 *
0-
02
b101 6
#502190000000
1!
1%
1-
12
#502200000000
0!
0%
b110 *
0-
02
b110 6
#502210000000
1!
1%
1-
12
#502220000000
0!
0%
b111 *
0-
02
b111 6
#502230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#502240000000
0!
0%
b0 *
0-
02
b0 6
#502250000000
1!
1%
1-
12
#502260000000
0!
0%
b1 *
0-
02
b1 6
#502270000000
1!
1%
1-
12
#502280000000
0!
0%
b10 *
0-
02
b10 6
#502290000000
1!
1%
1-
12
#502300000000
0!
0%
b11 *
0-
02
b11 6
#502310000000
1!
1%
1-
12
15
#502320000000
0!
0%
b100 *
0-
02
b100 6
#502330000000
1!
1%
1-
12
#502340000000
0!
0%
b101 *
0-
02
b101 6
#502350000000
1!
1%
1-
12
#502360000000
0!
0%
b110 *
0-
02
b110 6
#502370000000
1!
1%
1-
12
#502380000000
0!
0%
b111 *
0-
02
b111 6
#502390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#502400000000
0!
0%
b0 *
0-
02
b0 6
#502410000000
1!
1%
1-
12
#502420000000
0!
0%
b1 *
0-
02
b1 6
#502430000000
1!
1%
1-
12
#502440000000
0!
0%
b10 *
0-
02
b10 6
#502450000000
1!
1%
1-
12
#502460000000
0!
0%
b11 *
0-
02
b11 6
#502470000000
1!
1%
1-
12
15
#502480000000
0!
0%
b100 *
0-
02
b100 6
#502490000000
1!
1%
1-
12
#502500000000
0!
0%
b101 *
0-
02
b101 6
#502510000000
1!
1%
1-
12
#502520000000
0!
0%
b110 *
0-
02
b110 6
#502530000000
1!
1%
1-
12
#502540000000
0!
0%
b111 *
0-
02
b111 6
#502550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#502560000000
0!
0%
b0 *
0-
02
b0 6
#502570000000
1!
1%
1-
12
#502580000000
0!
0%
b1 *
0-
02
b1 6
#502590000000
1!
1%
1-
12
#502600000000
0!
0%
b10 *
0-
02
b10 6
#502610000000
1!
1%
1-
12
#502620000000
0!
0%
b11 *
0-
02
b11 6
#502630000000
1!
1%
1-
12
15
#502640000000
0!
0%
b100 *
0-
02
b100 6
#502650000000
1!
1%
1-
12
#502660000000
0!
0%
b101 *
0-
02
b101 6
#502670000000
1!
1%
1-
12
#502680000000
0!
0%
b110 *
0-
02
b110 6
#502690000000
1!
1%
1-
12
#502700000000
0!
0%
b111 *
0-
02
b111 6
#502710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#502720000000
0!
0%
b0 *
0-
02
b0 6
#502730000000
1!
1%
1-
12
#502740000000
0!
0%
b1 *
0-
02
b1 6
#502750000000
1!
1%
1-
12
#502760000000
0!
0%
b10 *
0-
02
b10 6
#502770000000
1!
1%
1-
12
#502780000000
0!
0%
b11 *
0-
02
b11 6
#502790000000
1!
1%
1-
12
15
#502800000000
0!
0%
b100 *
0-
02
b100 6
#502810000000
1!
1%
1-
12
#502820000000
0!
0%
b101 *
0-
02
b101 6
#502830000000
1!
1%
1-
12
#502840000000
0!
0%
b110 *
0-
02
b110 6
#502850000000
1!
1%
1-
12
#502860000000
0!
0%
b111 *
0-
02
b111 6
#502870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#502880000000
0!
0%
b0 *
0-
02
b0 6
#502890000000
1!
1%
1-
12
#502900000000
0!
0%
b1 *
0-
02
b1 6
#502910000000
1!
1%
1-
12
#502920000000
0!
0%
b10 *
0-
02
b10 6
#502930000000
1!
1%
1-
12
#502940000000
0!
0%
b11 *
0-
02
b11 6
#502950000000
1!
1%
1-
12
15
#502960000000
0!
0%
b100 *
0-
02
b100 6
#502970000000
1!
1%
1-
12
#502980000000
0!
0%
b101 *
0-
02
b101 6
#502990000000
1!
1%
1-
12
#503000000000
0!
0%
b110 *
0-
02
b110 6
#503010000000
1!
1%
1-
12
#503020000000
0!
0%
b111 *
0-
02
b111 6
#503030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#503040000000
0!
0%
b0 *
0-
02
b0 6
#503050000000
1!
1%
1-
12
#503060000000
0!
0%
b1 *
0-
02
b1 6
#503070000000
1!
1%
1-
12
#503080000000
0!
0%
b10 *
0-
02
b10 6
#503090000000
1!
1%
1-
12
#503100000000
0!
0%
b11 *
0-
02
b11 6
#503110000000
1!
1%
1-
12
15
#503120000000
0!
0%
b100 *
0-
02
b100 6
#503130000000
1!
1%
1-
12
#503140000000
0!
0%
b101 *
0-
02
b101 6
#503150000000
1!
1%
1-
12
#503160000000
0!
0%
b110 *
0-
02
b110 6
#503170000000
1!
1%
1-
12
#503180000000
0!
0%
b111 *
0-
02
b111 6
#503190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#503200000000
0!
0%
b0 *
0-
02
b0 6
#503210000000
1!
1%
1-
12
#503220000000
0!
0%
b1 *
0-
02
b1 6
#503230000000
1!
1%
1-
12
#503240000000
0!
0%
b10 *
0-
02
b10 6
#503250000000
1!
1%
1-
12
#503260000000
0!
0%
b11 *
0-
02
b11 6
#503270000000
1!
1%
1-
12
15
#503280000000
0!
0%
b100 *
0-
02
b100 6
#503290000000
1!
1%
1-
12
#503300000000
0!
0%
b101 *
0-
02
b101 6
#503310000000
1!
1%
1-
12
#503320000000
0!
0%
b110 *
0-
02
b110 6
#503330000000
1!
1%
1-
12
#503340000000
0!
0%
b111 *
0-
02
b111 6
#503350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#503360000000
0!
0%
b0 *
0-
02
b0 6
#503370000000
1!
1%
1-
12
#503380000000
0!
0%
b1 *
0-
02
b1 6
#503390000000
1!
1%
1-
12
#503400000000
0!
0%
b10 *
0-
02
b10 6
#503410000000
1!
1%
1-
12
#503420000000
0!
0%
b11 *
0-
02
b11 6
#503430000000
1!
1%
1-
12
15
#503440000000
0!
0%
b100 *
0-
02
b100 6
#503450000000
1!
1%
1-
12
#503460000000
0!
0%
b101 *
0-
02
b101 6
#503470000000
1!
1%
1-
12
#503480000000
0!
0%
b110 *
0-
02
b110 6
#503490000000
1!
1%
1-
12
#503500000000
0!
0%
b111 *
0-
02
b111 6
#503510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#503520000000
0!
0%
b0 *
0-
02
b0 6
#503530000000
1!
1%
1-
12
#503540000000
0!
0%
b1 *
0-
02
b1 6
#503550000000
1!
1%
1-
12
#503560000000
0!
0%
b10 *
0-
02
b10 6
#503570000000
1!
1%
1-
12
#503580000000
0!
0%
b11 *
0-
02
b11 6
#503590000000
1!
1%
1-
12
15
#503600000000
0!
0%
b100 *
0-
02
b100 6
#503610000000
1!
1%
1-
12
#503620000000
0!
0%
b101 *
0-
02
b101 6
#503630000000
1!
1%
1-
12
#503640000000
0!
0%
b110 *
0-
02
b110 6
#503650000000
1!
1%
1-
12
#503660000000
0!
0%
b111 *
0-
02
b111 6
#503670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#503680000000
0!
0%
b0 *
0-
02
b0 6
#503690000000
1!
1%
1-
12
#503700000000
0!
0%
b1 *
0-
02
b1 6
#503710000000
1!
1%
1-
12
#503720000000
0!
0%
b10 *
0-
02
b10 6
#503730000000
1!
1%
1-
12
#503740000000
0!
0%
b11 *
0-
02
b11 6
#503750000000
1!
1%
1-
12
15
#503760000000
0!
0%
b100 *
0-
02
b100 6
#503770000000
1!
1%
1-
12
#503780000000
0!
0%
b101 *
0-
02
b101 6
#503790000000
1!
1%
1-
12
#503800000000
0!
0%
b110 *
0-
02
b110 6
#503810000000
1!
1%
1-
12
#503820000000
0!
0%
b111 *
0-
02
b111 6
#503830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#503840000000
0!
0%
b0 *
0-
02
b0 6
#503850000000
1!
1%
1-
12
#503860000000
0!
0%
b1 *
0-
02
b1 6
#503870000000
1!
1%
1-
12
#503880000000
0!
0%
b10 *
0-
02
b10 6
#503890000000
1!
1%
1-
12
#503900000000
0!
0%
b11 *
0-
02
b11 6
#503910000000
1!
1%
1-
12
15
#503920000000
0!
0%
b100 *
0-
02
b100 6
#503930000000
1!
1%
1-
12
#503940000000
0!
0%
b101 *
0-
02
b101 6
#503950000000
1!
1%
1-
12
#503960000000
0!
0%
b110 *
0-
02
b110 6
#503970000000
1!
1%
1-
12
#503980000000
0!
0%
b111 *
0-
02
b111 6
#503990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#504000000000
0!
0%
b0 *
0-
02
b0 6
#504010000000
1!
1%
1-
12
#504020000000
0!
0%
b1 *
0-
02
b1 6
#504030000000
1!
1%
1-
12
#504040000000
0!
0%
b10 *
0-
02
b10 6
#504050000000
1!
1%
1-
12
#504060000000
0!
0%
b11 *
0-
02
b11 6
#504070000000
1!
1%
1-
12
15
#504080000000
0!
0%
b100 *
0-
02
b100 6
#504090000000
1!
1%
1-
12
#504100000000
0!
0%
b101 *
0-
02
b101 6
#504110000000
1!
1%
1-
12
#504120000000
0!
0%
b110 *
0-
02
b110 6
#504130000000
1!
1%
1-
12
#504140000000
0!
0%
b111 *
0-
02
b111 6
#504150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#504160000000
0!
0%
b0 *
0-
02
b0 6
#504170000000
1!
1%
1-
12
#504180000000
0!
0%
b1 *
0-
02
b1 6
#504190000000
1!
1%
1-
12
#504200000000
0!
0%
b10 *
0-
02
b10 6
#504210000000
1!
1%
1-
12
#504220000000
0!
0%
b11 *
0-
02
b11 6
#504230000000
1!
1%
1-
12
15
#504240000000
0!
0%
b100 *
0-
02
b100 6
#504250000000
1!
1%
1-
12
#504260000000
0!
0%
b101 *
0-
02
b101 6
#504270000000
1!
1%
1-
12
#504280000000
0!
0%
b110 *
0-
02
b110 6
#504290000000
1!
1%
1-
12
#504300000000
0!
0%
b111 *
0-
02
b111 6
#504310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#504320000000
0!
0%
b0 *
0-
02
b0 6
#504330000000
1!
1%
1-
12
#504340000000
0!
0%
b1 *
0-
02
b1 6
#504350000000
1!
1%
1-
12
#504360000000
0!
0%
b10 *
0-
02
b10 6
#504370000000
1!
1%
1-
12
#504380000000
0!
0%
b11 *
0-
02
b11 6
#504390000000
1!
1%
1-
12
15
#504400000000
0!
0%
b100 *
0-
02
b100 6
#504410000000
1!
1%
1-
12
#504420000000
0!
0%
b101 *
0-
02
b101 6
#504430000000
1!
1%
1-
12
#504440000000
0!
0%
b110 *
0-
02
b110 6
#504450000000
1!
1%
1-
12
#504460000000
0!
0%
b111 *
0-
02
b111 6
#504470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#504480000000
0!
0%
b0 *
0-
02
b0 6
#504490000000
1!
1%
1-
12
#504500000000
0!
0%
b1 *
0-
02
b1 6
#504510000000
1!
1%
1-
12
#504520000000
0!
0%
b10 *
0-
02
b10 6
#504530000000
1!
1%
1-
12
#504540000000
0!
0%
b11 *
0-
02
b11 6
#504550000000
1!
1%
1-
12
15
#504560000000
0!
0%
b100 *
0-
02
b100 6
#504570000000
1!
1%
1-
12
#504580000000
0!
0%
b101 *
0-
02
b101 6
#504590000000
1!
1%
1-
12
#504600000000
0!
0%
b110 *
0-
02
b110 6
#504610000000
1!
1%
1-
12
#504620000000
0!
0%
b111 *
0-
02
b111 6
#504630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#504640000000
0!
0%
b0 *
0-
02
b0 6
#504650000000
1!
1%
1-
12
#504660000000
0!
0%
b1 *
0-
02
b1 6
#504670000000
1!
1%
1-
12
#504680000000
0!
0%
b10 *
0-
02
b10 6
#504690000000
1!
1%
1-
12
#504700000000
0!
0%
b11 *
0-
02
b11 6
#504710000000
1!
1%
1-
12
15
#504720000000
0!
0%
b100 *
0-
02
b100 6
#504730000000
1!
1%
1-
12
#504740000000
0!
0%
b101 *
0-
02
b101 6
#504750000000
1!
1%
1-
12
#504760000000
0!
0%
b110 *
0-
02
b110 6
#504770000000
1!
1%
1-
12
#504780000000
0!
0%
b111 *
0-
02
b111 6
#504790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#504800000000
0!
0%
b0 *
0-
02
b0 6
#504810000000
1!
1%
1-
12
#504820000000
0!
0%
b1 *
0-
02
b1 6
#504830000000
1!
1%
1-
12
#504840000000
0!
0%
b10 *
0-
02
b10 6
#504850000000
1!
1%
1-
12
#504860000000
0!
0%
b11 *
0-
02
b11 6
#504870000000
1!
1%
1-
12
15
#504880000000
0!
0%
b100 *
0-
02
b100 6
#504890000000
1!
1%
1-
12
#504900000000
0!
0%
b101 *
0-
02
b101 6
#504910000000
1!
1%
1-
12
#504920000000
0!
0%
b110 *
0-
02
b110 6
#504930000000
1!
1%
1-
12
#504940000000
0!
0%
b111 *
0-
02
b111 6
#504950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#504960000000
0!
0%
b0 *
0-
02
b0 6
#504970000000
1!
1%
1-
12
#504980000000
0!
0%
b1 *
0-
02
b1 6
#504990000000
1!
1%
1-
12
#505000000000
0!
0%
b10 *
0-
02
b10 6
#505010000000
1!
1%
1-
12
#505020000000
0!
0%
b11 *
0-
02
b11 6
#505030000000
1!
1%
1-
12
15
#505040000000
0!
0%
b100 *
0-
02
b100 6
#505050000000
1!
1%
1-
12
#505060000000
0!
0%
b101 *
0-
02
b101 6
#505070000000
1!
1%
1-
12
#505080000000
0!
0%
b110 *
0-
02
b110 6
#505090000000
1!
1%
1-
12
#505100000000
0!
0%
b111 *
0-
02
b111 6
#505110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#505120000000
0!
0%
b0 *
0-
02
b0 6
#505130000000
1!
1%
1-
12
#505140000000
0!
0%
b1 *
0-
02
b1 6
#505150000000
1!
1%
1-
12
#505160000000
0!
0%
b10 *
0-
02
b10 6
#505170000000
1!
1%
1-
12
#505180000000
0!
0%
b11 *
0-
02
b11 6
#505190000000
1!
1%
1-
12
15
#505200000000
0!
0%
b100 *
0-
02
b100 6
#505210000000
1!
1%
1-
12
#505220000000
0!
0%
b101 *
0-
02
b101 6
#505230000000
1!
1%
1-
12
#505240000000
0!
0%
b110 *
0-
02
b110 6
#505250000000
1!
1%
1-
12
#505260000000
0!
0%
b111 *
0-
02
b111 6
#505270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#505280000000
0!
0%
b0 *
0-
02
b0 6
#505290000000
1!
1%
1-
12
#505300000000
0!
0%
b1 *
0-
02
b1 6
#505310000000
1!
1%
1-
12
#505320000000
0!
0%
b10 *
0-
02
b10 6
#505330000000
1!
1%
1-
12
#505340000000
0!
0%
b11 *
0-
02
b11 6
#505350000000
1!
1%
1-
12
15
#505360000000
0!
0%
b100 *
0-
02
b100 6
#505370000000
1!
1%
1-
12
#505380000000
0!
0%
b101 *
0-
02
b101 6
#505390000000
1!
1%
1-
12
#505400000000
0!
0%
b110 *
0-
02
b110 6
#505410000000
1!
1%
1-
12
#505420000000
0!
0%
b111 *
0-
02
b111 6
#505430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#505440000000
0!
0%
b0 *
0-
02
b0 6
#505450000000
1!
1%
1-
12
#505460000000
0!
0%
b1 *
0-
02
b1 6
#505470000000
1!
1%
1-
12
#505480000000
0!
0%
b10 *
0-
02
b10 6
#505490000000
1!
1%
1-
12
#505500000000
0!
0%
b11 *
0-
02
b11 6
#505510000000
1!
1%
1-
12
15
#505520000000
0!
0%
b100 *
0-
02
b100 6
#505530000000
1!
1%
1-
12
#505540000000
0!
0%
b101 *
0-
02
b101 6
#505550000000
1!
1%
1-
12
#505560000000
0!
0%
b110 *
0-
02
b110 6
#505570000000
1!
1%
1-
12
#505580000000
0!
0%
b111 *
0-
02
b111 6
#505590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#505600000000
0!
0%
b0 *
0-
02
b0 6
#505610000000
1!
1%
1-
12
#505620000000
0!
0%
b1 *
0-
02
b1 6
#505630000000
1!
1%
1-
12
#505640000000
0!
0%
b10 *
0-
02
b10 6
#505650000000
1!
1%
1-
12
#505660000000
0!
0%
b11 *
0-
02
b11 6
#505670000000
1!
1%
1-
12
15
#505680000000
0!
0%
b100 *
0-
02
b100 6
#505690000000
1!
1%
1-
12
#505700000000
0!
0%
b101 *
0-
02
b101 6
#505710000000
1!
1%
1-
12
#505720000000
0!
0%
b110 *
0-
02
b110 6
#505730000000
1!
1%
1-
12
#505740000000
0!
0%
b111 *
0-
02
b111 6
#505750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#505760000000
0!
0%
b0 *
0-
02
b0 6
#505770000000
1!
1%
1-
12
#505780000000
0!
0%
b1 *
0-
02
b1 6
#505790000000
1!
1%
1-
12
#505800000000
0!
0%
b10 *
0-
02
b10 6
#505810000000
1!
1%
1-
12
#505820000000
0!
0%
b11 *
0-
02
b11 6
#505830000000
1!
1%
1-
12
15
#505840000000
0!
0%
b100 *
0-
02
b100 6
#505850000000
1!
1%
1-
12
#505860000000
0!
0%
b101 *
0-
02
b101 6
#505870000000
1!
1%
1-
12
#505880000000
0!
0%
b110 *
0-
02
b110 6
#505890000000
1!
1%
1-
12
#505900000000
0!
0%
b111 *
0-
02
b111 6
#505910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#505920000000
0!
0%
b0 *
0-
02
b0 6
#505930000000
1!
1%
1-
12
#505940000000
0!
0%
b1 *
0-
02
b1 6
#505950000000
1!
1%
1-
12
#505960000000
0!
0%
b10 *
0-
02
b10 6
#505970000000
1!
1%
1-
12
#505980000000
0!
0%
b11 *
0-
02
b11 6
#505990000000
1!
1%
1-
12
15
#506000000000
0!
0%
b100 *
0-
02
b100 6
#506010000000
1!
1%
1-
12
#506020000000
0!
0%
b101 *
0-
02
b101 6
#506030000000
1!
1%
1-
12
#506040000000
0!
0%
b110 *
0-
02
b110 6
#506050000000
1!
1%
1-
12
#506060000000
0!
0%
b111 *
0-
02
b111 6
#506070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#506080000000
0!
0%
b0 *
0-
02
b0 6
#506090000000
1!
1%
1-
12
#506100000000
0!
0%
b1 *
0-
02
b1 6
#506110000000
1!
1%
1-
12
#506120000000
0!
0%
b10 *
0-
02
b10 6
#506130000000
1!
1%
1-
12
#506140000000
0!
0%
b11 *
0-
02
b11 6
#506150000000
1!
1%
1-
12
15
#506160000000
0!
0%
b100 *
0-
02
b100 6
#506170000000
1!
1%
1-
12
#506180000000
0!
0%
b101 *
0-
02
b101 6
#506190000000
1!
1%
1-
12
#506200000000
0!
0%
b110 *
0-
02
b110 6
#506210000000
1!
1%
1-
12
#506220000000
0!
0%
b111 *
0-
02
b111 6
#506230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#506240000000
0!
0%
b0 *
0-
02
b0 6
#506250000000
1!
1%
1-
12
#506260000000
0!
0%
b1 *
0-
02
b1 6
#506270000000
1!
1%
1-
12
#506280000000
0!
0%
b10 *
0-
02
b10 6
#506290000000
1!
1%
1-
12
#506300000000
0!
0%
b11 *
0-
02
b11 6
#506310000000
1!
1%
1-
12
15
#506320000000
0!
0%
b100 *
0-
02
b100 6
#506330000000
1!
1%
1-
12
#506340000000
0!
0%
b101 *
0-
02
b101 6
#506350000000
1!
1%
1-
12
#506360000000
0!
0%
b110 *
0-
02
b110 6
#506370000000
1!
1%
1-
12
#506380000000
0!
0%
b111 *
0-
02
b111 6
#506390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#506400000000
0!
0%
b0 *
0-
02
b0 6
#506410000000
1!
1%
1-
12
#506420000000
0!
0%
b1 *
0-
02
b1 6
#506430000000
1!
1%
1-
12
#506440000000
0!
0%
b10 *
0-
02
b10 6
#506450000000
1!
1%
1-
12
#506460000000
0!
0%
b11 *
0-
02
b11 6
#506470000000
1!
1%
1-
12
15
#506480000000
0!
0%
b100 *
0-
02
b100 6
#506490000000
1!
1%
1-
12
#506500000000
0!
0%
b101 *
0-
02
b101 6
#506510000000
1!
1%
1-
12
#506520000000
0!
0%
b110 *
0-
02
b110 6
#506530000000
1!
1%
1-
12
#506540000000
0!
0%
b111 *
0-
02
b111 6
#506550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#506560000000
0!
0%
b0 *
0-
02
b0 6
#506570000000
1!
1%
1-
12
#506580000000
0!
0%
b1 *
0-
02
b1 6
#506590000000
1!
1%
1-
12
#506600000000
0!
0%
b10 *
0-
02
b10 6
#506610000000
1!
1%
1-
12
#506620000000
0!
0%
b11 *
0-
02
b11 6
#506630000000
1!
1%
1-
12
15
#506640000000
0!
0%
b100 *
0-
02
b100 6
#506650000000
1!
1%
1-
12
#506660000000
0!
0%
b101 *
0-
02
b101 6
#506670000000
1!
1%
1-
12
#506680000000
0!
0%
b110 *
0-
02
b110 6
#506690000000
1!
1%
1-
12
#506700000000
0!
0%
b111 *
0-
02
b111 6
#506710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#506720000000
0!
0%
b0 *
0-
02
b0 6
#506730000000
1!
1%
1-
12
#506740000000
0!
0%
b1 *
0-
02
b1 6
#506750000000
1!
1%
1-
12
#506760000000
0!
0%
b10 *
0-
02
b10 6
#506770000000
1!
1%
1-
12
#506780000000
0!
0%
b11 *
0-
02
b11 6
#506790000000
1!
1%
1-
12
15
#506800000000
0!
0%
b100 *
0-
02
b100 6
#506810000000
1!
1%
1-
12
#506820000000
0!
0%
b101 *
0-
02
b101 6
#506830000000
1!
1%
1-
12
#506840000000
0!
0%
b110 *
0-
02
b110 6
#506850000000
1!
1%
1-
12
#506860000000
0!
0%
b111 *
0-
02
b111 6
#506870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#506880000000
0!
0%
b0 *
0-
02
b0 6
#506890000000
1!
1%
1-
12
#506900000000
0!
0%
b1 *
0-
02
b1 6
#506910000000
1!
1%
1-
12
#506920000000
0!
0%
b10 *
0-
02
b10 6
#506930000000
1!
1%
1-
12
#506940000000
0!
0%
b11 *
0-
02
b11 6
#506950000000
1!
1%
1-
12
15
#506960000000
0!
0%
b100 *
0-
02
b100 6
#506970000000
1!
1%
1-
12
#506980000000
0!
0%
b101 *
0-
02
b101 6
#506990000000
1!
1%
1-
12
#507000000000
0!
0%
b110 *
0-
02
b110 6
#507010000000
1!
1%
1-
12
#507020000000
0!
0%
b111 *
0-
02
b111 6
#507030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#507040000000
0!
0%
b0 *
0-
02
b0 6
#507050000000
1!
1%
1-
12
#507060000000
0!
0%
b1 *
0-
02
b1 6
#507070000000
1!
1%
1-
12
#507080000000
0!
0%
b10 *
0-
02
b10 6
#507090000000
1!
1%
1-
12
#507100000000
0!
0%
b11 *
0-
02
b11 6
#507110000000
1!
1%
1-
12
15
#507120000000
0!
0%
b100 *
0-
02
b100 6
#507130000000
1!
1%
1-
12
#507140000000
0!
0%
b101 *
0-
02
b101 6
#507150000000
1!
1%
1-
12
#507160000000
0!
0%
b110 *
0-
02
b110 6
#507170000000
1!
1%
1-
12
#507180000000
0!
0%
b111 *
0-
02
b111 6
#507190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#507200000000
0!
0%
b0 *
0-
02
b0 6
#507210000000
1!
1%
1-
12
#507220000000
0!
0%
b1 *
0-
02
b1 6
#507230000000
1!
1%
1-
12
#507240000000
0!
0%
b10 *
0-
02
b10 6
#507250000000
1!
1%
1-
12
#507260000000
0!
0%
b11 *
0-
02
b11 6
#507270000000
1!
1%
1-
12
15
#507280000000
0!
0%
b100 *
0-
02
b100 6
#507290000000
1!
1%
1-
12
#507300000000
0!
0%
b101 *
0-
02
b101 6
#507310000000
1!
1%
1-
12
#507320000000
0!
0%
b110 *
0-
02
b110 6
#507330000000
1!
1%
1-
12
#507340000000
0!
0%
b111 *
0-
02
b111 6
#507350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#507360000000
0!
0%
b0 *
0-
02
b0 6
#507370000000
1!
1%
1-
12
#507380000000
0!
0%
b1 *
0-
02
b1 6
#507390000000
1!
1%
1-
12
#507400000000
0!
0%
b10 *
0-
02
b10 6
#507410000000
1!
1%
1-
12
#507420000000
0!
0%
b11 *
0-
02
b11 6
#507430000000
1!
1%
1-
12
15
#507440000000
0!
0%
b100 *
0-
02
b100 6
#507450000000
1!
1%
1-
12
#507460000000
0!
0%
b101 *
0-
02
b101 6
#507470000000
1!
1%
1-
12
#507480000000
0!
0%
b110 *
0-
02
b110 6
#507490000000
1!
1%
1-
12
#507500000000
0!
0%
b111 *
0-
02
b111 6
#507510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#507520000000
0!
0%
b0 *
0-
02
b0 6
#507530000000
1!
1%
1-
12
#507540000000
0!
0%
b1 *
0-
02
b1 6
#507550000000
1!
1%
1-
12
#507560000000
0!
0%
b10 *
0-
02
b10 6
#507570000000
1!
1%
1-
12
#507580000000
0!
0%
b11 *
0-
02
b11 6
#507590000000
1!
1%
1-
12
15
#507600000000
0!
0%
b100 *
0-
02
b100 6
#507610000000
1!
1%
1-
12
#507620000000
0!
0%
b101 *
0-
02
b101 6
#507630000000
1!
1%
1-
12
#507640000000
0!
0%
b110 *
0-
02
b110 6
#507650000000
1!
1%
1-
12
#507660000000
0!
0%
b111 *
0-
02
b111 6
#507670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#507680000000
0!
0%
b0 *
0-
02
b0 6
#507690000000
1!
1%
1-
12
#507700000000
0!
0%
b1 *
0-
02
b1 6
#507710000000
1!
1%
1-
12
#507720000000
0!
0%
b10 *
0-
02
b10 6
#507730000000
1!
1%
1-
12
#507740000000
0!
0%
b11 *
0-
02
b11 6
#507750000000
1!
1%
1-
12
15
#507760000000
0!
0%
b100 *
0-
02
b100 6
#507770000000
1!
1%
1-
12
#507780000000
0!
0%
b101 *
0-
02
b101 6
#507790000000
1!
1%
1-
12
#507800000000
0!
0%
b110 *
0-
02
b110 6
#507810000000
1!
1%
1-
12
#507820000000
0!
0%
b111 *
0-
02
b111 6
#507830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#507840000000
0!
0%
b0 *
0-
02
b0 6
#507850000000
1!
1%
1-
12
#507860000000
0!
0%
b1 *
0-
02
b1 6
#507870000000
1!
1%
1-
12
#507880000000
0!
0%
b10 *
0-
02
b10 6
#507890000000
1!
1%
1-
12
#507900000000
0!
0%
b11 *
0-
02
b11 6
#507910000000
1!
1%
1-
12
15
#507920000000
0!
0%
b100 *
0-
02
b100 6
#507930000000
1!
1%
1-
12
#507940000000
0!
0%
b101 *
0-
02
b101 6
#507950000000
1!
1%
1-
12
#507960000000
0!
0%
b110 *
0-
02
b110 6
#507970000000
1!
1%
1-
12
#507980000000
0!
0%
b111 *
0-
02
b111 6
#507990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#508000000000
0!
0%
b0 *
0-
02
b0 6
#508010000000
1!
1%
1-
12
#508020000000
0!
0%
b1 *
0-
02
b1 6
#508030000000
1!
1%
1-
12
#508040000000
0!
0%
b10 *
0-
02
b10 6
#508050000000
1!
1%
1-
12
#508060000000
0!
0%
b11 *
0-
02
b11 6
#508070000000
1!
1%
1-
12
15
#508080000000
0!
0%
b100 *
0-
02
b100 6
#508090000000
1!
1%
1-
12
#508100000000
0!
0%
b101 *
0-
02
b101 6
#508110000000
1!
1%
1-
12
#508120000000
0!
0%
b110 *
0-
02
b110 6
#508130000000
1!
1%
1-
12
#508140000000
0!
0%
b111 *
0-
02
b111 6
#508150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#508160000000
0!
0%
b0 *
0-
02
b0 6
#508170000000
1!
1%
1-
12
#508180000000
0!
0%
b1 *
0-
02
b1 6
#508190000000
1!
1%
1-
12
#508200000000
0!
0%
b10 *
0-
02
b10 6
#508210000000
1!
1%
1-
12
#508220000000
0!
0%
b11 *
0-
02
b11 6
#508230000000
1!
1%
1-
12
15
#508240000000
0!
0%
b100 *
0-
02
b100 6
#508250000000
1!
1%
1-
12
#508260000000
0!
0%
b101 *
0-
02
b101 6
#508270000000
1!
1%
1-
12
#508280000000
0!
0%
b110 *
0-
02
b110 6
#508290000000
1!
1%
1-
12
#508300000000
0!
0%
b111 *
0-
02
b111 6
#508310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#508320000000
0!
0%
b0 *
0-
02
b0 6
#508330000000
1!
1%
1-
12
#508340000000
0!
0%
b1 *
0-
02
b1 6
#508350000000
1!
1%
1-
12
#508360000000
0!
0%
b10 *
0-
02
b10 6
#508370000000
1!
1%
1-
12
#508380000000
0!
0%
b11 *
0-
02
b11 6
#508390000000
1!
1%
1-
12
15
#508400000000
0!
0%
b100 *
0-
02
b100 6
#508410000000
1!
1%
1-
12
#508420000000
0!
0%
b101 *
0-
02
b101 6
#508430000000
1!
1%
1-
12
#508440000000
0!
0%
b110 *
0-
02
b110 6
#508450000000
1!
1%
1-
12
#508460000000
0!
0%
b111 *
0-
02
b111 6
#508470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#508480000000
0!
0%
b0 *
0-
02
b0 6
#508490000000
1!
1%
1-
12
#508500000000
0!
0%
b1 *
0-
02
b1 6
#508510000000
1!
1%
1-
12
#508520000000
0!
0%
b10 *
0-
02
b10 6
#508530000000
1!
1%
1-
12
#508540000000
0!
0%
b11 *
0-
02
b11 6
#508550000000
1!
1%
1-
12
15
#508560000000
0!
0%
b100 *
0-
02
b100 6
#508570000000
1!
1%
1-
12
#508580000000
0!
0%
b101 *
0-
02
b101 6
#508590000000
1!
1%
1-
12
#508600000000
0!
0%
b110 *
0-
02
b110 6
#508610000000
1!
1%
1-
12
#508620000000
0!
0%
b111 *
0-
02
b111 6
#508630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#508640000000
0!
0%
b0 *
0-
02
b0 6
#508650000000
1!
1%
1-
12
#508660000000
0!
0%
b1 *
0-
02
b1 6
#508670000000
1!
1%
1-
12
#508680000000
0!
0%
b10 *
0-
02
b10 6
#508690000000
1!
1%
1-
12
#508700000000
0!
0%
b11 *
0-
02
b11 6
#508710000000
1!
1%
1-
12
15
#508720000000
0!
0%
b100 *
0-
02
b100 6
#508730000000
1!
1%
1-
12
#508740000000
0!
0%
b101 *
0-
02
b101 6
#508750000000
1!
1%
1-
12
#508760000000
0!
0%
b110 *
0-
02
b110 6
#508770000000
1!
1%
1-
12
#508780000000
0!
0%
b111 *
0-
02
b111 6
#508790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#508800000000
0!
0%
b0 *
0-
02
b0 6
#508810000000
1!
1%
1-
12
#508820000000
0!
0%
b1 *
0-
02
b1 6
#508830000000
1!
1%
1-
12
#508840000000
0!
0%
b10 *
0-
02
b10 6
#508850000000
1!
1%
1-
12
#508860000000
0!
0%
b11 *
0-
02
b11 6
#508870000000
1!
1%
1-
12
15
#508880000000
0!
0%
b100 *
0-
02
b100 6
#508890000000
1!
1%
1-
12
#508900000000
0!
0%
b101 *
0-
02
b101 6
#508910000000
1!
1%
1-
12
#508920000000
0!
0%
b110 *
0-
02
b110 6
#508930000000
1!
1%
1-
12
#508940000000
0!
0%
b111 *
0-
02
b111 6
#508950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#508960000000
0!
0%
b0 *
0-
02
b0 6
#508970000000
1!
1%
1-
12
#508980000000
0!
0%
b1 *
0-
02
b1 6
#508990000000
1!
1%
1-
12
#509000000000
0!
0%
b10 *
0-
02
b10 6
#509010000000
1!
1%
1-
12
#509020000000
0!
0%
b11 *
0-
02
b11 6
#509030000000
1!
1%
1-
12
15
#509040000000
0!
0%
b100 *
0-
02
b100 6
#509050000000
1!
1%
1-
12
#509060000000
0!
0%
b101 *
0-
02
b101 6
#509070000000
1!
1%
1-
12
#509080000000
0!
0%
b110 *
0-
02
b110 6
#509090000000
1!
1%
1-
12
#509100000000
0!
0%
b111 *
0-
02
b111 6
#509110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#509120000000
0!
0%
b0 *
0-
02
b0 6
#509130000000
1!
1%
1-
12
#509140000000
0!
0%
b1 *
0-
02
b1 6
#509150000000
1!
1%
1-
12
#509160000000
0!
0%
b10 *
0-
02
b10 6
#509170000000
1!
1%
1-
12
#509180000000
0!
0%
b11 *
0-
02
b11 6
#509190000000
1!
1%
1-
12
15
#509200000000
0!
0%
b100 *
0-
02
b100 6
#509210000000
1!
1%
1-
12
#509220000000
0!
0%
b101 *
0-
02
b101 6
#509230000000
1!
1%
1-
12
#509240000000
0!
0%
b110 *
0-
02
b110 6
#509250000000
1!
1%
1-
12
#509260000000
0!
0%
b111 *
0-
02
b111 6
#509270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#509280000000
0!
0%
b0 *
0-
02
b0 6
#509290000000
1!
1%
1-
12
#509300000000
0!
0%
b1 *
0-
02
b1 6
#509310000000
1!
1%
1-
12
#509320000000
0!
0%
b10 *
0-
02
b10 6
#509330000000
1!
1%
1-
12
#509340000000
0!
0%
b11 *
0-
02
b11 6
#509350000000
1!
1%
1-
12
15
#509360000000
0!
0%
b100 *
0-
02
b100 6
#509370000000
1!
1%
1-
12
#509380000000
0!
0%
b101 *
0-
02
b101 6
#509390000000
1!
1%
1-
12
#509400000000
0!
0%
b110 *
0-
02
b110 6
#509410000000
1!
1%
1-
12
#509420000000
0!
0%
b111 *
0-
02
b111 6
#509430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#509440000000
0!
0%
b0 *
0-
02
b0 6
#509450000000
1!
1%
1-
12
#509460000000
0!
0%
b1 *
0-
02
b1 6
#509470000000
1!
1%
1-
12
#509480000000
0!
0%
b10 *
0-
02
b10 6
#509490000000
1!
1%
1-
12
#509500000000
0!
0%
b11 *
0-
02
b11 6
#509510000000
1!
1%
1-
12
15
#509520000000
0!
0%
b100 *
0-
02
b100 6
#509530000000
1!
1%
1-
12
#509540000000
0!
0%
b101 *
0-
02
b101 6
#509550000000
1!
1%
1-
12
#509560000000
0!
0%
b110 *
0-
02
b110 6
#509570000000
1!
1%
1-
12
#509580000000
0!
0%
b111 *
0-
02
b111 6
#509590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#509600000000
0!
0%
b0 *
0-
02
b0 6
#509610000000
1!
1%
1-
12
#509620000000
0!
0%
b1 *
0-
02
b1 6
#509630000000
1!
1%
1-
12
#509640000000
0!
0%
b10 *
0-
02
b10 6
#509650000000
1!
1%
1-
12
#509660000000
0!
0%
b11 *
0-
02
b11 6
#509670000000
1!
1%
1-
12
15
#509680000000
0!
0%
b100 *
0-
02
b100 6
#509690000000
1!
1%
1-
12
#509700000000
0!
0%
b101 *
0-
02
b101 6
#509710000000
1!
1%
1-
12
#509720000000
0!
0%
b110 *
0-
02
b110 6
#509730000000
1!
1%
1-
12
#509740000000
0!
0%
b111 *
0-
02
b111 6
#509750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#509760000000
0!
0%
b0 *
0-
02
b0 6
#509770000000
1!
1%
1-
12
#509780000000
0!
0%
b1 *
0-
02
b1 6
#509790000000
1!
1%
1-
12
#509800000000
0!
0%
b10 *
0-
02
b10 6
#509810000000
1!
1%
1-
12
#509820000000
0!
0%
b11 *
0-
02
b11 6
#509830000000
1!
1%
1-
12
15
#509840000000
0!
0%
b100 *
0-
02
b100 6
#509850000000
1!
1%
1-
12
#509860000000
0!
0%
b101 *
0-
02
b101 6
#509870000000
1!
1%
1-
12
#509880000000
0!
0%
b110 *
0-
02
b110 6
#509890000000
1!
1%
1-
12
#509900000000
0!
0%
b111 *
0-
02
b111 6
#509910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#509920000000
0!
0%
b0 *
0-
02
b0 6
#509930000000
1!
1%
1-
12
#509940000000
0!
0%
b1 *
0-
02
b1 6
#509950000000
1!
1%
1-
12
#509960000000
0!
0%
b10 *
0-
02
b10 6
#509970000000
1!
1%
1-
12
#509980000000
0!
0%
b11 *
0-
02
b11 6
#509990000000
1!
1%
1-
12
15
#510000000000
0!
0%
b100 *
0-
02
b100 6
#510010000000
1!
1%
1-
12
#510020000000
0!
0%
b101 *
0-
02
b101 6
#510030000000
1!
1%
1-
12
#510040000000
0!
0%
b110 *
0-
02
b110 6
#510050000000
1!
1%
1-
12
#510060000000
0!
0%
b111 *
0-
02
b111 6
#510070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#510080000000
0!
0%
b0 *
0-
02
b0 6
#510090000000
1!
1%
1-
12
#510100000000
0!
0%
b1 *
0-
02
b1 6
#510110000000
1!
1%
1-
12
#510120000000
0!
0%
b10 *
0-
02
b10 6
#510130000000
1!
1%
1-
12
#510140000000
0!
0%
b11 *
0-
02
b11 6
#510150000000
1!
1%
1-
12
15
#510160000000
0!
0%
b100 *
0-
02
b100 6
#510170000000
1!
1%
1-
12
#510180000000
0!
0%
b101 *
0-
02
b101 6
#510190000000
1!
1%
1-
12
#510200000000
0!
0%
b110 *
0-
02
b110 6
#510210000000
1!
1%
1-
12
#510220000000
0!
0%
b111 *
0-
02
b111 6
#510230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#510240000000
0!
0%
b0 *
0-
02
b0 6
#510250000000
1!
1%
1-
12
#510260000000
0!
0%
b1 *
0-
02
b1 6
#510270000000
1!
1%
1-
12
#510280000000
0!
0%
b10 *
0-
02
b10 6
#510290000000
1!
1%
1-
12
#510300000000
0!
0%
b11 *
0-
02
b11 6
#510310000000
1!
1%
1-
12
15
#510320000000
0!
0%
b100 *
0-
02
b100 6
#510330000000
1!
1%
1-
12
#510340000000
0!
0%
b101 *
0-
02
b101 6
#510350000000
1!
1%
1-
12
#510360000000
0!
0%
b110 *
0-
02
b110 6
#510370000000
1!
1%
1-
12
#510380000000
0!
0%
b111 *
0-
02
b111 6
#510390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#510400000000
0!
0%
b0 *
0-
02
b0 6
#510410000000
1!
1%
1-
12
#510420000000
0!
0%
b1 *
0-
02
b1 6
#510430000000
1!
1%
1-
12
#510440000000
0!
0%
b10 *
0-
02
b10 6
#510450000000
1!
1%
1-
12
#510460000000
0!
0%
b11 *
0-
02
b11 6
#510470000000
1!
1%
1-
12
15
#510480000000
0!
0%
b100 *
0-
02
b100 6
#510490000000
1!
1%
1-
12
#510500000000
0!
0%
b101 *
0-
02
b101 6
#510510000000
1!
1%
1-
12
#510520000000
0!
0%
b110 *
0-
02
b110 6
#510530000000
1!
1%
1-
12
#510540000000
0!
0%
b111 *
0-
02
b111 6
#510550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#510560000000
0!
0%
b0 *
0-
02
b0 6
#510570000000
1!
1%
1-
12
#510580000000
0!
0%
b1 *
0-
02
b1 6
#510590000000
1!
1%
1-
12
#510600000000
0!
0%
b10 *
0-
02
b10 6
#510610000000
1!
1%
1-
12
#510620000000
0!
0%
b11 *
0-
02
b11 6
#510630000000
1!
1%
1-
12
15
#510640000000
0!
0%
b100 *
0-
02
b100 6
#510650000000
1!
1%
1-
12
#510660000000
0!
0%
b101 *
0-
02
b101 6
#510670000000
1!
1%
1-
12
#510680000000
0!
0%
b110 *
0-
02
b110 6
#510690000000
1!
1%
1-
12
#510700000000
0!
0%
b111 *
0-
02
b111 6
#510710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#510720000000
0!
0%
b0 *
0-
02
b0 6
#510730000000
1!
1%
1-
12
#510740000000
0!
0%
b1 *
0-
02
b1 6
#510750000000
1!
1%
1-
12
#510760000000
0!
0%
b10 *
0-
02
b10 6
#510770000000
1!
1%
1-
12
#510780000000
0!
0%
b11 *
0-
02
b11 6
#510790000000
1!
1%
1-
12
15
#510800000000
0!
0%
b100 *
0-
02
b100 6
#510810000000
1!
1%
1-
12
#510820000000
0!
0%
b101 *
0-
02
b101 6
#510830000000
1!
1%
1-
12
#510840000000
0!
0%
b110 *
0-
02
b110 6
#510850000000
1!
1%
1-
12
#510860000000
0!
0%
b111 *
0-
02
b111 6
#510870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#510880000000
0!
0%
b0 *
0-
02
b0 6
#510890000000
1!
1%
1-
12
#510900000000
0!
0%
b1 *
0-
02
b1 6
#510910000000
1!
1%
1-
12
#510920000000
0!
0%
b10 *
0-
02
b10 6
#510930000000
1!
1%
1-
12
#510940000000
0!
0%
b11 *
0-
02
b11 6
#510950000000
1!
1%
1-
12
15
#510960000000
0!
0%
b100 *
0-
02
b100 6
#510970000000
1!
1%
1-
12
#510980000000
0!
0%
b101 *
0-
02
b101 6
#510990000000
1!
1%
1-
12
#511000000000
0!
0%
b110 *
0-
02
b110 6
#511010000000
1!
1%
1-
12
#511020000000
0!
0%
b111 *
0-
02
b111 6
#511030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#511040000000
0!
0%
b0 *
0-
02
b0 6
#511050000000
1!
1%
1-
12
#511060000000
0!
0%
b1 *
0-
02
b1 6
#511070000000
1!
1%
1-
12
#511080000000
0!
0%
b10 *
0-
02
b10 6
#511090000000
1!
1%
1-
12
#511100000000
0!
0%
b11 *
0-
02
b11 6
#511110000000
1!
1%
1-
12
15
#511120000000
0!
0%
b100 *
0-
02
b100 6
#511130000000
1!
1%
1-
12
#511140000000
0!
0%
b101 *
0-
02
b101 6
#511150000000
1!
1%
1-
12
#511160000000
0!
0%
b110 *
0-
02
b110 6
#511170000000
1!
1%
1-
12
#511180000000
0!
0%
b111 *
0-
02
b111 6
#511190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#511200000000
0!
0%
b0 *
0-
02
b0 6
#511210000000
1!
1%
1-
12
#511220000000
0!
0%
b1 *
0-
02
b1 6
#511230000000
1!
1%
1-
12
#511240000000
0!
0%
b10 *
0-
02
b10 6
#511250000000
1!
1%
1-
12
#511260000000
0!
0%
b11 *
0-
02
b11 6
#511270000000
1!
1%
1-
12
15
#511280000000
0!
0%
b100 *
0-
02
b100 6
#511290000000
1!
1%
1-
12
#511300000000
0!
0%
b101 *
0-
02
b101 6
#511310000000
1!
1%
1-
12
#511320000000
0!
0%
b110 *
0-
02
b110 6
#511330000000
1!
1%
1-
12
#511340000000
0!
0%
b111 *
0-
02
b111 6
#511350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#511360000000
0!
0%
b0 *
0-
02
b0 6
#511370000000
1!
1%
1-
12
#511380000000
0!
0%
b1 *
0-
02
b1 6
#511390000000
1!
1%
1-
12
#511400000000
0!
0%
b10 *
0-
02
b10 6
#511410000000
1!
1%
1-
12
#511420000000
0!
0%
b11 *
0-
02
b11 6
#511430000000
1!
1%
1-
12
15
#511440000000
0!
0%
b100 *
0-
02
b100 6
#511450000000
1!
1%
1-
12
#511460000000
0!
0%
b101 *
0-
02
b101 6
#511470000000
1!
1%
1-
12
#511480000000
0!
0%
b110 *
0-
02
b110 6
#511490000000
1!
1%
1-
12
#511500000000
0!
0%
b111 *
0-
02
b111 6
#511510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#511520000000
0!
0%
b0 *
0-
02
b0 6
#511530000000
1!
1%
1-
12
#511540000000
0!
0%
b1 *
0-
02
b1 6
#511550000000
1!
1%
1-
12
#511560000000
0!
0%
b10 *
0-
02
b10 6
#511570000000
1!
1%
1-
12
#511580000000
0!
0%
b11 *
0-
02
b11 6
#511590000000
1!
1%
1-
12
15
#511600000000
0!
0%
b100 *
0-
02
b100 6
#511610000000
1!
1%
1-
12
#511620000000
0!
0%
b101 *
0-
02
b101 6
#511630000000
1!
1%
1-
12
#511640000000
0!
0%
b110 *
0-
02
b110 6
#511650000000
1!
1%
1-
12
#511660000000
0!
0%
b111 *
0-
02
b111 6
#511670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#511680000000
0!
0%
b0 *
0-
02
b0 6
#511690000000
1!
1%
1-
12
#511700000000
0!
0%
b1 *
0-
02
b1 6
#511710000000
1!
1%
1-
12
#511720000000
0!
0%
b10 *
0-
02
b10 6
#511730000000
1!
1%
1-
12
#511740000000
0!
0%
b11 *
0-
02
b11 6
#511750000000
1!
1%
1-
12
15
#511760000000
0!
0%
b100 *
0-
02
b100 6
#511770000000
1!
1%
1-
12
#511780000000
0!
0%
b101 *
0-
02
b101 6
#511790000000
1!
1%
1-
12
#511800000000
0!
0%
b110 *
0-
02
b110 6
#511810000000
1!
1%
1-
12
#511820000000
0!
0%
b111 *
0-
02
b111 6
#511830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#511840000000
0!
0%
b0 *
0-
02
b0 6
#511850000000
1!
1%
1-
12
#511860000000
0!
0%
b1 *
0-
02
b1 6
#511870000000
1!
1%
1-
12
#511880000000
0!
0%
b10 *
0-
02
b10 6
#511890000000
1!
1%
1-
12
#511900000000
0!
0%
b11 *
0-
02
b11 6
#511910000000
1!
1%
1-
12
15
#511920000000
0!
0%
b100 *
0-
02
b100 6
#511930000000
1!
1%
1-
12
#511940000000
0!
0%
b101 *
0-
02
b101 6
#511950000000
1!
1%
1-
12
#511960000000
0!
0%
b110 *
0-
02
b110 6
#511970000000
1!
1%
1-
12
#511980000000
0!
0%
b111 *
0-
02
b111 6
#511990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#512000000000
0!
0%
b0 *
0-
02
b0 6
#512010000000
1!
1%
1-
12
#512020000000
0!
0%
b1 *
0-
02
b1 6
#512030000000
1!
1%
1-
12
#512040000000
0!
0%
b10 *
0-
02
b10 6
#512050000000
1!
1%
1-
12
#512060000000
0!
0%
b11 *
0-
02
b11 6
#512070000000
1!
1%
1-
12
15
#512080000000
0!
0%
b100 *
0-
02
b100 6
#512090000000
1!
1%
1-
12
#512100000000
0!
0%
b101 *
0-
02
b101 6
#512110000000
1!
1%
1-
12
#512120000000
0!
0%
b110 *
0-
02
b110 6
#512130000000
1!
1%
1-
12
#512140000000
0!
0%
b111 *
0-
02
b111 6
#512150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#512160000000
0!
0%
b0 *
0-
02
b0 6
#512170000000
1!
1%
1-
12
#512180000000
0!
0%
b1 *
0-
02
b1 6
#512190000000
1!
1%
1-
12
#512200000000
0!
0%
b10 *
0-
02
b10 6
#512210000000
1!
1%
1-
12
#512220000000
0!
0%
b11 *
0-
02
b11 6
#512230000000
1!
1%
1-
12
15
#512240000000
0!
0%
b100 *
0-
02
b100 6
#512250000000
1!
1%
1-
12
#512260000000
0!
0%
b101 *
0-
02
b101 6
#512270000000
1!
1%
1-
12
#512280000000
0!
0%
b110 *
0-
02
b110 6
#512290000000
1!
1%
1-
12
#512300000000
0!
0%
b111 *
0-
02
b111 6
#512310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#512320000000
0!
0%
b0 *
0-
02
b0 6
#512330000000
1!
1%
1-
12
#512340000000
0!
0%
b1 *
0-
02
b1 6
#512350000000
1!
1%
1-
12
#512360000000
0!
0%
b10 *
0-
02
b10 6
#512370000000
1!
1%
1-
12
#512380000000
0!
0%
b11 *
0-
02
b11 6
#512390000000
1!
1%
1-
12
15
#512400000000
0!
0%
b100 *
0-
02
b100 6
#512410000000
1!
1%
1-
12
#512420000000
0!
0%
b101 *
0-
02
b101 6
#512430000000
1!
1%
1-
12
#512440000000
0!
0%
b110 *
0-
02
b110 6
#512450000000
1!
1%
1-
12
#512460000000
0!
0%
b111 *
0-
02
b111 6
#512470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#512480000000
0!
0%
b0 *
0-
02
b0 6
#512490000000
1!
1%
1-
12
#512500000000
0!
0%
b1 *
0-
02
b1 6
#512510000000
1!
1%
1-
12
#512520000000
0!
0%
b10 *
0-
02
b10 6
#512530000000
1!
1%
1-
12
#512540000000
0!
0%
b11 *
0-
02
b11 6
#512550000000
1!
1%
1-
12
15
#512560000000
0!
0%
b100 *
0-
02
b100 6
#512570000000
1!
1%
1-
12
#512580000000
0!
0%
b101 *
0-
02
b101 6
#512590000000
1!
1%
1-
12
#512600000000
0!
0%
b110 *
0-
02
b110 6
#512610000000
1!
1%
1-
12
#512620000000
0!
0%
b111 *
0-
02
b111 6
#512630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#512640000000
0!
0%
b0 *
0-
02
b0 6
#512650000000
1!
1%
1-
12
#512660000000
0!
0%
b1 *
0-
02
b1 6
#512670000000
1!
1%
1-
12
#512680000000
0!
0%
b10 *
0-
02
b10 6
#512690000000
1!
1%
1-
12
#512700000000
0!
0%
b11 *
0-
02
b11 6
#512710000000
1!
1%
1-
12
15
#512720000000
0!
0%
b100 *
0-
02
b100 6
#512730000000
1!
1%
1-
12
#512740000000
0!
0%
b101 *
0-
02
b101 6
#512750000000
1!
1%
1-
12
#512760000000
0!
0%
b110 *
0-
02
b110 6
#512770000000
1!
1%
1-
12
#512780000000
0!
0%
b111 *
0-
02
b111 6
#512790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#512800000000
0!
0%
b0 *
0-
02
b0 6
#512810000000
1!
1%
1-
12
#512820000000
0!
0%
b1 *
0-
02
b1 6
#512830000000
1!
1%
1-
12
#512840000000
0!
0%
b10 *
0-
02
b10 6
#512850000000
1!
1%
1-
12
#512860000000
0!
0%
b11 *
0-
02
b11 6
#512870000000
1!
1%
1-
12
15
#512880000000
0!
0%
b100 *
0-
02
b100 6
#512890000000
1!
1%
1-
12
#512900000000
0!
0%
b101 *
0-
02
b101 6
#512910000000
1!
1%
1-
12
#512920000000
0!
0%
b110 *
0-
02
b110 6
#512930000000
1!
1%
1-
12
#512940000000
0!
0%
b111 *
0-
02
b111 6
#512950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#512960000000
0!
0%
b0 *
0-
02
b0 6
#512970000000
1!
1%
1-
12
#512980000000
0!
0%
b1 *
0-
02
b1 6
#512990000000
1!
1%
1-
12
#513000000000
0!
0%
b10 *
0-
02
b10 6
#513010000000
1!
1%
1-
12
#513020000000
0!
0%
b11 *
0-
02
b11 6
#513030000000
1!
1%
1-
12
15
#513040000000
0!
0%
b100 *
0-
02
b100 6
#513050000000
1!
1%
1-
12
#513060000000
0!
0%
b101 *
0-
02
b101 6
#513070000000
1!
1%
1-
12
#513080000000
0!
0%
b110 *
0-
02
b110 6
#513090000000
1!
1%
1-
12
#513100000000
0!
0%
b111 *
0-
02
b111 6
#513110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#513120000000
0!
0%
b0 *
0-
02
b0 6
#513130000000
1!
1%
1-
12
#513140000000
0!
0%
b1 *
0-
02
b1 6
#513150000000
1!
1%
1-
12
#513160000000
0!
0%
b10 *
0-
02
b10 6
#513170000000
1!
1%
1-
12
#513180000000
0!
0%
b11 *
0-
02
b11 6
#513190000000
1!
1%
1-
12
15
#513200000000
0!
0%
b100 *
0-
02
b100 6
#513210000000
1!
1%
1-
12
#513220000000
0!
0%
b101 *
0-
02
b101 6
#513230000000
1!
1%
1-
12
#513240000000
0!
0%
b110 *
0-
02
b110 6
#513250000000
1!
1%
1-
12
#513260000000
0!
0%
b111 *
0-
02
b111 6
#513270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#513280000000
0!
0%
b0 *
0-
02
b0 6
#513290000000
1!
1%
1-
12
#513300000000
0!
0%
b1 *
0-
02
b1 6
#513310000000
1!
1%
1-
12
#513320000000
0!
0%
b10 *
0-
02
b10 6
#513330000000
1!
1%
1-
12
#513340000000
0!
0%
b11 *
0-
02
b11 6
#513350000000
1!
1%
1-
12
15
#513360000000
0!
0%
b100 *
0-
02
b100 6
#513370000000
1!
1%
1-
12
#513380000000
0!
0%
b101 *
0-
02
b101 6
#513390000000
1!
1%
1-
12
#513400000000
0!
0%
b110 *
0-
02
b110 6
#513410000000
1!
1%
1-
12
#513420000000
0!
0%
b111 *
0-
02
b111 6
#513430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#513440000000
0!
0%
b0 *
0-
02
b0 6
#513450000000
1!
1%
1-
12
#513460000000
0!
0%
b1 *
0-
02
b1 6
#513470000000
1!
1%
1-
12
#513480000000
0!
0%
b10 *
0-
02
b10 6
#513490000000
1!
1%
1-
12
#513500000000
0!
0%
b11 *
0-
02
b11 6
#513510000000
1!
1%
1-
12
15
#513520000000
0!
0%
b100 *
0-
02
b100 6
#513530000000
1!
1%
1-
12
#513540000000
0!
0%
b101 *
0-
02
b101 6
#513550000000
1!
1%
1-
12
#513560000000
0!
0%
b110 *
0-
02
b110 6
#513570000000
1!
1%
1-
12
#513580000000
0!
0%
b111 *
0-
02
b111 6
#513590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#513600000000
0!
0%
b0 *
0-
02
b0 6
#513610000000
1!
1%
1-
12
#513620000000
0!
0%
b1 *
0-
02
b1 6
#513630000000
1!
1%
1-
12
#513640000000
0!
0%
b10 *
0-
02
b10 6
#513650000000
1!
1%
1-
12
#513660000000
0!
0%
b11 *
0-
02
b11 6
#513670000000
1!
1%
1-
12
15
#513680000000
0!
0%
b100 *
0-
02
b100 6
#513690000000
1!
1%
1-
12
#513700000000
0!
0%
b101 *
0-
02
b101 6
#513710000000
1!
1%
1-
12
#513720000000
0!
0%
b110 *
0-
02
b110 6
#513730000000
1!
1%
1-
12
#513740000000
0!
0%
b111 *
0-
02
b111 6
#513750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#513760000000
0!
0%
b0 *
0-
02
b0 6
#513770000000
1!
1%
1-
12
#513780000000
0!
0%
b1 *
0-
02
b1 6
#513790000000
1!
1%
1-
12
#513800000000
0!
0%
b10 *
0-
02
b10 6
#513810000000
1!
1%
1-
12
#513820000000
0!
0%
b11 *
0-
02
b11 6
#513830000000
1!
1%
1-
12
15
#513840000000
0!
0%
b100 *
0-
02
b100 6
#513850000000
1!
1%
1-
12
#513860000000
0!
0%
b101 *
0-
02
b101 6
#513870000000
1!
1%
1-
12
#513880000000
0!
0%
b110 *
0-
02
b110 6
#513890000000
1!
1%
1-
12
#513900000000
0!
0%
b111 *
0-
02
b111 6
#513910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#513920000000
0!
0%
b0 *
0-
02
b0 6
#513930000000
1!
1%
1-
12
#513940000000
0!
0%
b1 *
0-
02
b1 6
#513950000000
1!
1%
1-
12
#513960000000
0!
0%
b10 *
0-
02
b10 6
#513970000000
1!
1%
1-
12
#513980000000
0!
0%
b11 *
0-
02
b11 6
#513990000000
1!
1%
1-
12
15
#514000000000
0!
0%
b100 *
0-
02
b100 6
#514010000000
1!
1%
1-
12
#514020000000
0!
0%
b101 *
0-
02
b101 6
#514030000000
1!
1%
1-
12
#514040000000
0!
0%
b110 *
0-
02
b110 6
#514050000000
1!
1%
1-
12
#514060000000
0!
0%
b111 *
0-
02
b111 6
#514070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#514080000000
0!
0%
b0 *
0-
02
b0 6
#514090000000
1!
1%
1-
12
#514100000000
0!
0%
b1 *
0-
02
b1 6
#514110000000
1!
1%
1-
12
#514120000000
0!
0%
b10 *
0-
02
b10 6
#514130000000
1!
1%
1-
12
#514140000000
0!
0%
b11 *
0-
02
b11 6
#514150000000
1!
1%
1-
12
15
#514160000000
0!
0%
b100 *
0-
02
b100 6
#514170000000
1!
1%
1-
12
#514180000000
0!
0%
b101 *
0-
02
b101 6
#514190000000
1!
1%
1-
12
#514200000000
0!
0%
b110 *
0-
02
b110 6
#514210000000
1!
1%
1-
12
#514220000000
0!
0%
b111 *
0-
02
b111 6
#514230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#514240000000
0!
0%
b0 *
0-
02
b0 6
#514250000000
1!
1%
1-
12
#514260000000
0!
0%
b1 *
0-
02
b1 6
#514270000000
1!
1%
1-
12
#514280000000
0!
0%
b10 *
0-
02
b10 6
#514290000000
1!
1%
1-
12
#514300000000
0!
0%
b11 *
0-
02
b11 6
#514310000000
1!
1%
1-
12
15
#514320000000
0!
0%
b100 *
0-
02
b100 6
#514330000000
1!
1%
1-
12
#514340000000
0!
0%
b101 *
0-
02
b101 6
#514350000000
1!
1%
1-
12
#514360000000
0!
0%
b110 *
0-
02
b110 6
#514370000000
1!
1%
1-
12
#514380000000
0!
0%
b111 *
0-
02
b111 6
#514390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#514400000000
0!
0%
b0 *
0-
02
b0 6
#514410000000
1!
1%
1-
12
#514420000000
0!
0%
b1 *
0-
02
b1 6
#514430000000
1!
1%
1-
12
#514440000000
0!
0%
b10 *
0-
02
b10 6
#514450000000
1!
1%
1-
12
#514460000000
0!
0%
b11 *
0-
02
b11 6
#514470000000
1!
1%
1-
12
15
#514480000000
0!
0%
b100 *
0-
02
b100 6
#514490000000
1!
1%
1-
12
#514500000000
0!
0%
b101 *
0-
02
b101 6
#514510000000
1!
1%
1-
12
#514520000000
0!
0%
b110 *
0-
02
b110 6
#514530000000
1!
1%
1-
12
#514540000000
0!
0%
b111 *
0-
02
b111 6
#514550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#514560000000
0!
0%
b0 *
0-
02
b0 6
#514570000000
1!
1%
1-
12
#514580000000
0!
0%
b1 *
0-
02
b1 6
#514590000000
1!
1%
1-
12
#514600000000
0!
0%
b10 *
0-
02
b10 6
#514610000000
1!
1%
1-
12
#514620000000
0!
0%
b11 *
0-
02
b11 6
#514630000000
1!
1%
1-
12
15
#514640000000
0!
0%
b100 *
0-
02
b100 6
#514650000000
1!
1%
1-
12
#514660000000
0!
0%
b101 *
0-
02
b101 6
#514670000000
1!
1%
1-
12
#514680000000
0!
0%
b110 *
0-
02
b110 6
#514690000000
1!
1%
1-
12
#514700000000
0!
0%
b111 *
0-
02
b111 6
#514710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#514720000000
0!
0%
b0 *
0-
02
b0 6
#514730000000
1!
1%
1-
12
#514740000000
0!
0%
b1 *
0-
02
b1 6
#514750000000
1!
1%
1-
12
#514760000000
0!
0%
b10 *
0-
02
b10 6
#514770000000
1!
1%
1-
12
#514780000000
0!
0%
b11 *
0-
02
b11 6
#514790000000
1!
1%
1-
12
15
#514800000000
0!
0%
b100 *
0-
02
b100 6
#514810000000
1!
1%
1-
12
#514820000000
0!
0%
b101 *
0-
02
b101 6
#514830000000
1!
1%
1-
12
#514840000000
0!
0%
b110 *
0-
02
b110 6
#514850000000
1!
1%
1-
12
#514860000000
0!
0%
b111 *
0-
02
b111 6
#514870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#514880000000
0!
0%
b0 *
0-
02
b0 6
#514890000000
1!
1%
1-
12
#514900000000
0!
0%
b1 *
0-
02
b1 6
#514910000000
1!
1%
1-
12
#514920000000
0!
0%
b10 *
0-
02
b10 6
#514930000000
1!
1%
1-
12
#514940000000
0!
0%
b11 *
0-
02
b11 6
#514950000000
1!
1%
1-
12
15
#514960000000
0!
0%
b100 *
0-
02
b100 6
#514970000000
1!
1%
1-
12
#514980000000
0!
0%
b101 *
0-
02
b101 6
#514990000000
1!
1%
1-
12
#515000000000
0!
0%
b110 *
0-
02
b110 6
#515010000000
1!
1%
1-
12
#515020000000
0!
0%
b111 *
0-
02
b111 6
#515030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#515040000000
0!
0%
b0 *
0-
02
b0 6
#515050000000
1!
1%
1-
12
#515060000000
0!
0%
b1 *
0-
02
b1 6
#515070000000
1!
1%
1-
12
#515080000000
0!
0%
b10 *
0-
02
b10 6
#515090000000
1!
1%
1-
12
#515100000000
0!
0%
b11 *
0-
02
b11 6
#515110000000
1!
1%
1-
12
15
#515120000000
0!
0%
b100 *
0-
02
b100 6
#515130000000
1!
1%
1-
12
#515140000000
0!
0%
b101 *
0-
02
b101 6
#515150000000
1!
1%
1-
12
#515160000000
0!
0%
b110 *
0-
02
b110 6
#515170000000
1!
1%
1-
12
#515180000000
0!
0%
b111 *
0-
02
b111 6
#515190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#515200000000
0!
0%
b0 *
0-
02
b0 6
#515210000000
1!
1%
1-
12
#515220000000
0!
0%
b1 *
0-
02
b1 6
#515230000000
1!
1%
1-
12
#515240000000
0!
0%
b10 *
0-
02
b10 6
#515250000000
1!
1%
1-
12
#515260000000
0!
0%
b11 *
0-
02
b11 6
#515270000000
1!
1%
1-
12
15
#515280000000
0!
0%
b100 *
0-
02
b100 6
#515290000000
1!
1%
1-
12
#515300000000
0!
0%
b101 *
0-
02
b101 6
#515310000000
1!
1%
1-
12
#515320000000
0!
0%
b110 *
0-
02
b110 6
#515330000000
1!
1%
1-
12
#515340000000
0!
0%
b111 *
0-
02
b111 6
#515350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#515360000000
0!
0%
b0 *
0-
02
b0 6
#515370000000
1!
1%
1-
12
#515380000000
0!
0%
b1 *
0-
02
b1 6
#515390000000
1!
1%
1-
12
#515400000000
0!
0%
b10 *
0-
02
b10 6
#515410000000
1!
1%
1-
12
#515420000000
0!
0%
b11 *
0-
02
b11 6
#515430000000
1!
1%
1-
12
15
#515440000000
0!
0%
b100 *
0-
02
b100 6
#515450000000
1!
1%
1-
12
#515460000000
0!
0%
b101 *
0-
02
b101 6
#515470000000
1!
1%
1-
12
#515480000000
0!
0%
b110 *
0-
02
b110 6
#515490000000
1!
1%
1-
12
#515500000000
0!
0%
b111 *
0-
02
b111 6
#515510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#515520000000
0!
0%
b0 *
0-
02
b0 6
#515530000000
1!
1%
1-
12
#515540000000
0!
0%
b1 *
0-
02
b1 6
#515550000000
1!
1%
1-
12
#515560000000
0!
0%
b10 *
0-
02
b10 6
#515570000000
1!
1%
1-
12
#515580000000
0!
0%
b11 *
0-
02
b11 6
#515590000000
1!
1%
1-
12
15
#515600000000
0!
0%
b100 *
0-
02
b100 6
#515610000000
1!
1%
1-
12
#515620000000
0!
0%
b101 *
0-
02
b101 6
#515630000000
1!
1%
1-
12
#515640000000
0!
0%
b110 *
0-
02
b110 6
#515650000000
1!
1%
1-
12
#515660000000
0!
0%
b111 *
0-
02
b111 6
#515670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#515680000000
0!
0%
b0 *
0-
02
b0 6
#515690000000
1!
1%
1-
12
#515700000000
0!
0%
b1 *
0-
02
b1 6
#515710000000
1!
1%
1-
12
#515720000000
0!
0%
b10 *
0-
02
b10 6
#515730000000
1!
1%
1-
12
#515740000000
0!
0%
b11 *
0-
02
b11 6
#515750000000
1!
1%
1-
12
15
#515760000000
0!
0%
b100 *
0-
02
b100 6
#515770000000
1!
1%
1-
12
#515780000000
0!
0%
b101 *
0-
02
b101 6
#515790000000
1!
1%
1-
12
#515800000000
0!
0%
b110 *
0-
02
b110 6
#515810000000
1!
1%
1-
12
#515820000000
0!
0%
b111 *
0-
02
b111 6
#515830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#515840000000
0!
0%
b0 *
0-
02
b0 6
#515850000000
1!
1%
1-
12
#515860000000
0!
0%
b1 *
0-
02
b1 6
#515870000000
1!
1%
1-
12
#515880000000
0!
0%
b10 *
0-
02
b10 6
#515890000000
1!
1%
1-
12
#515900000000
0!
0%
b11 *
0-
02
b11 6
#515910000000
1!
1%
1-
12
15
#515920000000
0!
0%
b100 *
0-
02
b100 6
#515930000000
1!
1%
1-
12
#515940000000
0!
0%
b101 *
0-
02
b101 6
#515950000000
1!
1%
1-
12
#515960000000
0!
0%
b110 *
0-
02
b110 6
#515970000000
1!
1%
1-
12
#515980000000
0!
0%
b111 *
0-
02
b111 6
#515990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#516000000000
0!
0%
b0 *
0-
02
b0 6
#516010000000
1!
1%
1-
12
#516020000000
0!
0%
b1 *
0-
02
b1 6
#516030000000
1!
1%
1-
12
#516040000000
0!
0%
b10 *
0-
02
b10 6
#516050000000
1!
1%
1-
12
#516060000000
0!
0%
b11 *
0-
02
b11 6
#516070000000
1!
1%
1-
12
15
#516080000000
0!
0%
b100 *
0-
02
b100 6
#516090000000
1!
1%
1-
12
#516100000000
0!
0%
b101 *
0-
02
b101 6
#516110000000
1!
1%
1-
12
#516120000000
0!
0%
b110 *
0-
02
b110 6
#516130000000
1!
1%
1-
12
#516140000000
0!
0%
b111 *
0-
02
b111 6
#516150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#516160000000
0!
0%
b0 *
0-
02
b0 6
#516170000000
1!
1%
1-
12
#516180000000
0!
0%
b1 *
0-
02
b1 6
#516190000000
1!
1%
1-
12
#516200000000
0!
0%
b10 *
0-
02
b10 6
#516210000000
1!
1%
1-
12
#516220000000
0!
0%
b11 *
0-
02
b11 6
#516230000000
1!
1%
1-
12
15
#516240000000
0!
0%
b100 *
0-
02
b100 6
#516250000000
1!
1%
1-
12
#516260000000
0!
0%
b101 *
0-
02
b101 6
#516270000000
1!
1%
1-
12
#516280000000
0!
0%
b110 *
0-
02
b110 6
#516290000000
1!
1%
1-
12
#516300000000
0!
0%
b111 *
0-
02
b111 6
#516310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#516320000000
0!
0%
b0 *
0-
02
b0 6
#516330000000
1!
1%
1-
12
#516340000000
0!
0%
b1 *
0-
02
b1 6
#516350000000
1!
1%
1-
12
#516360000000
0!
0%
b10 *
0-
02
b10 6
#516370000000
1!
1%
1-
12
#516380000000
0!
0%
b11 *
0-
02
b11 6
#516390000000
1!
1%
1-
12
15
#516400000000
0!
0%
b100 *
0-
02
b100 6
#516410000000
1!
1%
1-
12
#516420000000
0!
0%
b101 *
0-
02
b101 6
#516430000000
1!
1%
1-
12
#516440000000
0!
0%
b110 *
0-
02
b110 6
#516450000000
1!
1%
1-
12
#516460000000
0!
0%
b111 *
0-
02
b111 6
#516470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#516480000000
0!
0%
b0 *
0-
02
b0 6
#516490000000
1!
1%
1-
12
#516500000000
0!
0%
b1 *
0-
02
b1 6
#516510000000
1!
1%
1-
12
#516520000000
0!
0%
b10 *
0-
02
b10 6
#516530000000
1!
1%
1-
12
#516540000000
0!
0%
b11 *
0-
02
b11 6
#516550000000
1!
1%
1-
12
15
#516560000000
0!
0%
b100 *
0-
02
b100 6
#516570000000
1!
1%
1-
12
#516580000000
0!
0%
b101 *
0-
02
b101 6
#516590000000
1!
1%
1-
12
#516600000000
0!
0%
b110 *
0-
02
b110 6
#516610000000
1!
1%
1-
12
#516620000000
0!
0%
b111 *
0-
02
b111 6
#516630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#516640000000
0!
0%
b0 *
0-
02
b0 6
#516650000000
1!
1%
1-
12
#516660000000
0!
0%
b1 *
0-
02
b1 6
#516670000000
1!
1%
1-
12
#516680000000
0!
0%
b10 *
0-
02
b10 6
#516690000000
1!
1%
1-
12
#516700000000
0!
0%
b11 *
0-
02
b11 6
#516710000000
1!
1%
1-
12
15
#516720000000
0!
0%
b100 *
0-
02
b100 6
#516730000000
1!
1%
1-
12
#516740000000
0!
0%
b101 *
0-
02
b101 6
#516750000000
1!
1%
1-
12
#516760000000
0!
0%
b110 *
0-
02
b110 6
#516770000000
1!
1%
1-
12
#516780000000
0!
0%
b111 *
0-
02
b111 6
#516790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#516800000000
0!
0%
b0 *
0-
02
b0 6
#516810000000
1!
1%
1-
12
#516820000000
0!
0%
b1 *
0-
02
b1 6
#516830000000
1!
1%
1-
12
#516840000000
0!
0%
b10 *
0-
02
b10 6
#516850000000
1!
1%
1-
12
#516860000000
0!
0%
b11 *
0-
02
b11 6
#516870000000
1!
1%
1-
12
15
#516880000000
0!
0%
b100 *
0-
02
b100 6
#516890000000
1!
1%
1-
12
#516900000000
0!
0%
b101 *
0-
02
b101 6
#516910000000
1!
1%
1-
12
#516920000000
0!
0%
b110 *
0-
02
b110 6
#516930000000
1!
1%
1-
12
#516940000000
0!
0%
b111 *
0-
02
b111 6
#516950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#516960000000
0!
0%
b0 *
0-
02
b0 6
#516970000000
1!
1%
1-
12
#516980000000
0!
0%
b1 *
0-
02
b1 6
#516990000000
1!
1%
1-
12
#517000000000
0!
0%
b10 *
0-
02
b10 6
#517010000000
1!
1%
1-
12
#517020000000
0!
0%
b11 *
0-
02
b11 6
#517030000000
1!
1%
1-
12
15
#517040000000
0!
0%
b100 *
0-
02
b100 6
#517050000000
1!
1%
1-
12
#517060000000
0!
0%
b101 *
0-
02
b101 6
#517070000000
1!
1%
1-
12
#517080000000
0!
0%
b110 *
0-
02
b110 6
#517090000000
1!
1%
1-
12
#517100000000
0!
0%
b111 *
0-
02
b111 6
#517110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#517120000000
0!
0%
b0 *
0-
02
b0 6
#517130000000
1!
1%
1-
12
#517140000000
0!
0%
b1 *
0-
02
b1 6
#517150000000
1!
1%
1-
12
#517160000000
0!
0%
b10 *
0-
02
b10 6
#517170000000
1!
1%
1-
12
#517180000000
0!
0%
b11 *
0-
02
b11 6
#517190000000
1!
1%
1-
12
15
#517200000000
0!
0%
b100 *
0-
02
b100 6
#517210000000
1!
1%
1-
12
#517220000000
0!
0%
b101 *
0-
02
b101 6
#517230000000
1!
1%
1-
12
#517240000000
0!
0%
b110 *
0-
02
b110 6
#517250000000
1!
1%
1-
12
#517260000000
0!
0%
b111 *
0-
02
b111 6
#517270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#517280000000
0!
0%
b0 *
0-
02
b0 6
#517290000000
1!
1%
1-
12
#517300000000
0!
0%
b1 *
0-
02
b1 6
#517310000000
1!
1%
1-
12
#517320000000
0!
0%
b10 *
0-
02
b10 6
#517330000000
1!
1%
1-
12
#517340000000
0!
0%
b11 *
0-
02
b11 6
#517350000000
1!
1%
1-
12
15
#517360000000
0!
0%
b100 *
0-
02
b100 6
#517370000000
1!
1%
1-
12
#517380000000
0!
0%
b101 *
0-
02
b101 6
#517390000000
1!
1%
1-
12
#517400000000
0!
0%
b110 *
0-
02
b110 6
#517410000000
1!
1%
1-
12
#517420000000
0!
0%
b111 *
0-
02
b111 6
#517430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#517440000000
0!
0%
b0 *
0-
02
b0 6
#517450000000
1!
1%
1-
12
#517460000000
0!
0%
b1 *
0-
02
b1 6
#517470000000
1!
1%
1-
12
#517480000000
0!
0%
b10 *
0-
02
b10 6
#517490000000
1!
1%
1-
12
#517500000000
0!
0%
b11 *
0-
02
b11 6
#517510000000
1!
1%
1-
12
15
#517520000000
0!
0%
b100 *
0-
02
b100 6
#517530000000
1!
1%
1-
12
#517540000000
0!
0%
b101 *
0-
02
b101 6
#517550000000
1!
1%
1-
12
#517560000000
0!
0%
b110 *
0-
02
b110 6
#517570000000
1!
1%
1-
12
#517580000000
0!
0%
b111 *
0-
02
b111 6
#517590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#517600000000
0!
0%
b0 *
0-
02
b0 6
#517610000000
1!
1%
1-
12
#517620000000
0!
0%
b1 *
0-
02
b1 6
#517630000000
1!
1%
1-
12
#517640000000
0!
0%
b10 *
0-
02
b10 6
#517650000000
1!
1%
1-
12
#517660000000
0!
0%
b11 *
0-
02
b11 6
#517670000000
1!
1%
1-
12
15
#517680000000
0!
0%
b100 *
0-
02
b100 6
#517690000000
1!
1%
1-
12
#517700000000
0!
0%
b101 *
0-
02
b101 6
#517710000000
1!
1%
1-
12
#517720000000
0!
0%
b110 *
0-
02
b110 6
#517730000000
1!
1%
1-
12
#517740000000
0!
0%
b111 *
0-
02
b111 6
#517750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#517760000000
0!
0%
b0 *
0-
02
b0 6
#517770000000
1!
1%
1-
12
#517780000000
0!
0%
b1 *
0-
02
b1 6
#517790000000
1!
1%
1-
12
#517800000000
0!
0%
b10 *
0-
02
b10 6
#517810000000
1!
1%
1-
12
#517820000000
0!
0%
b11 *
0-
02
b11 6
#517830000000
1!
1%
1-
12
15
#517840000000
0!
0%
b100 *
0-
02
b100 6
#517850000000
1!
1%
1-
12
#517860000000
0!
0%
b101 *
0-
02
b101 6
#517870000000
1!
1%
1-
12
#517880000000
0!
0%
b110 *
0-
02
b110 6
#517890000000
1!
1%
1-
12
#517900000000
0!
0%
b111 *
0-
02
b111 6
#517910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#517920000000
0!
0%
b0 *
0-
02
b0 6
#517930000000
1!
1%
1-
12
#517940000000
0!
0%
b1 *
0-
02
b1 6
#517950000000
1!
1%
1-
12
#517960000000
0!
0%
b10 *
0-
02
b10 6
#517970000000
1!
1%
1-
12
#517980000000
0!
0%
b11 *
0-
02
b11 6
#517990000000
1!
1%
1-
12
15
#518000000000
0!
0%
b100 *
0-
02
b100 6
#518010000000
1!
1%
1-
12
#518020000000
0!
0%
b101 *
0-
02
b101 6
#518030000000
1!
1%
1-
12
#518040000000
0!
0%
b110 *
0-
02
b110 6
#518050000000
1!
1%
1-
12
#518060000000
0!
0%
b111 *
0-
02
b111 6
#518070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#518080000000
0!
0%
b0 *
0-
02
b0 6
#518090000000
1!
1%
1-
12
#518100000000
0!
0%
b1 *
0-
02
b1 6
#518110000000
1!
1%
1-
12
#518120000000
0!
0%
b10 *
0-
02
b10 6
#518130000000
1!
1%
1-
12
#518140000000
0!
0%
b11 *
0-
02
b11 6
#518150000000
1!
1%
1-
12
15
#518160000000
0!
0%
b100 *
0-
02
b100 6
#518170000000
1!
1%
1-
12
#518180000000
0!
0%
b101 *
0-
02
b101 6
#518190000000
1!
1%
1-
12
#518200000000
0!
0%
b110 *
0-
02
b110 6
#518210000000
1!
1%
1-
12
#518220000000
0!
0%
b111 *
0-
02
b111 6
#518230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#518240000000
0!
0%
b0 *
0-
02
b0 6
#518250000000
1!
1%
1-
12
#518260000000
0!
0%
b1 *
0-
02
b1 6
#518270000000
1!
1%
1-
12
#518280000000
0!
0%
b10 *
0-
02
b10 6
#518290000000
1!
1%
1-
12
#518300000000
0!
0%
b11 *
0-
02
b11 6
#518310000000
1!
1%
1-
12
15
#518320000000
0!
0%
b100 *
0-
02
b100 6
#518330000000
1!
1%
1-
12
#518340000000
0!
0%
b101 *
0-
02
b101 6
#518350000000
1!
1%
1-
12
#518360000000
0!
0%
b110 *
0-
02
b110 6
#518370000000
1!
1%
1-
12
#518380000000
0!
0%
b111 *
0-
02
b111 6
#518390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#518400000000
0!
0%
b0 *
0-
02
b0 6
#518410000000
1!
1%
1-
12
#518420000000
0!
0%
b1 *
0-
02
b1 6
#518430000000
1!
1%
1-
12
#518440000000
0!
0%
b10 *
0-
02
b10 6
#518450000000
1!
1%
1-
12
#518460000000
0!
0%
b11 *
0-
02
b11 6
#518470000000
1!
1%
1-
12
15
#518480000000
0!
0%
b100 *
0-
02
b100 6
#518490000000
1!
1%
1-
12
#518500000000
0!
0%
b101 *
0-
02
b101 6
#518510000000
1!
1%
1-
12
#518520000000
0!
0%
b110 *
0-
02
b110 6
#518530000000
1!
1%
1-
12
#518540000000
0!
0%
b111 *
0-
02
b111 6
#518550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#518560000000
0!
0%
b0 *
0-
02
b0 6
#518570000000
1!
1%
1-
12
#518580000000
0!
0%
b1 *
0-
02
b1 6
#518590000000
1!
1%
1-
12
#518600000000
0!
0%
b10 *
0-
02
b10 6
#518610000000
1!
1%
1-
12
#518620000000
0!
0%
b11 *
0-
02
b11 6
#518630000000
1!
1%
1-
12
15
#518640000000
0!
0%
b100 *
0-
02
b100 6
#518650000000
1!
1%
1-
12
#518660000000
0!
0%
b101 *
0-
02
b101 6
#518670000000
1!
1%
1-
12
#518680000000
0!
0%
b110 *
0-
02
b110 6
#518690000000
1!
1%
1-
12
#518700000000
0!
0%
b111 *
0-
02
b111 6
#518710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#518720000000
0!
0%
b0 *
0-
02
b0 6
#518730000000
1!
1%
1-
12
#518740000000
0!
0%
b1 *
0-
02
b1 6
#518750000000
1!
1%
1-
12
#518760000000
0!
0%
b10 *
0-
02
b10 6
#518770000000
1!
1%
1-
12
#518780000000
0!
0%
b11 *
0-
02
b11 6
#518790000000
1!
1%
1-
12
15
#518800000000
0!
0%
b100 *
0-
02
b100 6
#518810000000
1!
1%
1-
12
#518820000000
0!
0%
b101 *
0-
02
b101 6
#518830000000
1!
1%
1-
12
#518840000000
0!
0%
b110 *
0-
02
b110 6
#518850000000
1!
1%
1-
12
#518860000000
0!
0%
b111 *
0-
02
b111 6
#518870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#518880000000
0!
0%
b0 *
0-
02
b0 6
#518890000000
1!
1%
1-
12
#518900000000
0!
0%
b1 *
0-
02
b1 6
#518910000000
1!
1%
1-
12
#518920000000
0!
0%
b10 *
0-
02
b10 6
#518930000000
1!
1%
1-
12
#518940000000
0!
0%
b11 *
0-
02
b11 6
#518950000000
1!
1%
1-
12
15
#518960000000
0!
0%
b100 *
0-
02
b100 6
#518970000000
1!
1%
1-
12
#518980000000
0!
0%
b101 *
0-
02
b101 6
#518990000000
1!
1%
1-
12
#519000000000
0!
0%
b110 *
0-
02
b110 6
#519010000000
1!
1%
1-
12
#519020000000
0!
0%
b111 *
0-
02
b111 6
#519030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#519040000000
0!
0%
b0 *
0-
02
b0 6
#519050000000
1!
1%
1-
12
#519060000000
0!
0%
b1 *
0-
02
b1 6
#519070000000
1!
1%
1-
12
#519080000000
0!
0%
b10 *
0-
02
b10 6
#519090000000
1!
1%
1-
12
#519100000000
0!
0%
b11 *
0-
02
b11 6
#519110000000
1!
1%
1-
12
15
#519120000000
0!
0%
b100 *
0-
02
b100 6
#519130000000
1!
1%
1-
12
#519140000000
0!
0%
b101 *
0-
02
b101 6
#519150000000
1!
1%
1-
12
#519160000000
0!
0%
b110 *
0-
02
b110 6
#519170000000
1!
1%
1-
12
#519180000000
0!
0%
b111 *
0-
02
b111 6
#519190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#519200000000
0!
0%
b0 *
0-
02
b0 6
#519210000000
1!
1%
1-
12
#519220000000
0!
0%
b1 *
0-
02
b1 6
#519230000000
1!
1%
1-
12
#519240000000
0!
0%
b10 *
0-
02
b10 6
#519250000000
1!
1%
1-
12
#519260000000
0!
0%
b11 *
0-
02
b11 6
#519270000000
1!
1%
1-
12
15
#519280000000
0!
0%
b100 *
0-
02
b100 6
#519290000000
1!
1%
1-
12
#519300000000
0!
0%
b101 *
0-
02
b101 6
#519310000000
1!
1%
1-
12
#519320000000
0!
0%
b110 *
0-
02
b110 6
#519330000000
1!
1%
1-
12
#519340000000
0!
0%
b111 *
0-
02
b111 6
#519350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#519360000000
0!
0%
b0 *
0-
02
b0 6
#519370000000
1!
1%
1-
12
#519380000000
0!
0%
b1 *
0-
02
b1 6
#519390000000
1!
1%
1-
12
#519400000000
0!
0%
b10 *
0-
02
b10 6
#519410000000
1!
1%
1-
12
#519420000000
0!
0%
b11 *
0-
02
b11 6
#519430000000
1!
1%
1-
12
15
#519440000000
0!
0%
b100 *
0-
02
b100 6
#519450000000
1!
1%
1-
12
#519460000000
0!
0%
b101 *
0-
02
b101 6
#519470000000
1!
1%
1-
12
#519480000000
0!
0%
b110 *
0-
02
b110 6
#519490000000
1!
1%
1-
12
#519500000000
0!
0%
b111 *
0-
02
b111 6
#519510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#519520000000
0!
0%
b0 *
0-
02
b0 6
#519530000000
1!
1%
1-
12
#519540000000
0!
0%
b1 *
0-
02
b1 6
#519550000000
1!
1%
1-
12
#519560000000
0!
0%
b10 *
0-
02
b10 6
#519570000000
1!
1%
1-
12
#519580000000
0!
0%
b11 *
0-
02
b11 6
#519590000000
1!
1%
1-
12
15
#519600000000
0!
0%
b100 *
0-
02
b100 6
#519610000000
1!
1%
1-
12
#519620000000
0!
0%
b101 *
0-
02
b101 6
#519630000000
1!
1%
1-
12
#519640000000
0!
0%
b110 *
0-
02
b110 6
#519650000000
1!
1%
1-
12
#519660000000
0!
0%
b111 *
0-
02
b111 6
#519670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#519680000000
0!
0%
b0 *
0-
02
b0 6
#519690000000
1!
1%
1-
12
#519700000000
0!
0%
b1 *
0-
02
b1 6
#519710000000
1!
1%
1-
12
#519720000000
0!
0%
b10 *
0-
02
b10 6
#519730000000
1!
1%
1-
12
#519740000000
0!
0%
b11 *
0-
02
b11 6
#519750000000
1!
1%
1-
12
15
#519760000000
0!
0%
b100 *
0-
02
b100 6
#519770000000
1!
1%
1-
12
#519780000000
0!
0%
b101 *
0-
02
b101 6
#519790000000
1!
1%
1-
12
#519800000000
0!
0%
b110 *
0-
02
b110 6
#519810000000
1!
1%
1-
12
#519820000000
0!
0%
b111 *
0-
02
b111 6
#519830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#519840000000
0!
0%
b0 *
0-
02
b0 6
#519850000000
1!
1%
1-
12
#519860000000
0!
0%
b1 *
0-
02
b1 6
#519870000000
1!
1%
1-
12
#519880000000
0!
0%
b10 *
0-
02
b10 6
#519890000000
1!
1%
1-
12
#519900000000
0!
0%
b11 *
0-
02
b11 6
#519910000000
1!
1%
1-
12
15
#519920000000
0!
0%
b100 *
0-
02
b100 6
#519930000000
1!
1%
1-
12
#519940000000
0!
0%
b101 *
0-
02
b101 6
#519950000000
1!
1%
1-
12
#519960000000
0!
0%
b110 *
0-
02
b110 6
#519970000000
1!
1%
1-
12
#519980000000
0!
0%
b111 *
0-
02
b111 6
#519990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#520000000000
0!
0%
b0 *
0-
02
b0 6
#520010000000
1!
1%
1-
12
#520020000000
0!
0%
b1 *
0-
02
b1 6
#520030000000
1!
1%
1-
12
#520040000000
0!
0%
b10 *
0-
02
b10 6
#520050000000
1!
1%
1-
12
#520060000000
0!
0%
b11 *
0-
02
b11 6
#520070000000
1!
1%
1-
12
15
#520080000000
0!
0%
b100 *
0-
02
b100 6
#520090000000
1!
1%
1-
12
#520100000000
0!
0%
b101 *
0-
02
b101 6
#520110000000
1!
1%
1-
12
#520120000000
0!
0%
b110 *
0-
02
b110 6
#520130000000
1!
1%
1-
12
#520140000000
0!
0%
b111 *
0-
02
b111 6
#520150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#520160000000
0!
0%
b0 *
0-
02
b0 6
#520170000000
1!
1%
1-
12
#520180000000
0!
0%
b1 *
0-
02
b1 6
#520190000000
1!
1%
1-
12
#520200000000
0!
0%
b10 *
0-
02
b10 6
#520210000000
1!
1%
1-
12
#520220000000
0!
0%
b11 *
0-
02
b11 6
#520230000000
1!
1%
1-
12
15
#520240000000
0!
0%
b100 *
0-
02
b100 6
#520250000000
1!
1%
1-
12
#520260000000
0!
0%
b101 *
0-
02
b101 6
#520270000000
1!
1%
1-
12
#520280000000
0!
0%
b110 *
0-
02
b110 6
#520290000000
1!
1%
1-
12
#520300000000
0!
0%
b111 *
0-
02
b111 6
#520310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#520320000000
0!
0%
b0 *
0-
02
b0 6
#520330000000
1!
1%
1-
12
#520340000000
0!
0%
b1 *
0-
02
b1 6
#520350000000
1!
1%
1-
12
#520360000000
0!
0%
b10 *
0-
02
b10 6
#520370000000
1!
1%
1-
12
#520380000000
0!
0%
b11 *
0-
02
b11 6
#520390000000
1!
1%
1-
12
15
#520400000000
0!
0%
b100 *
0-
02
b100 6
#520410000000
1!
1%
1-
12
#520420000000
0!
0%
b101 *
0-
02
b101 6
#520430000000
1!
1%
1-
12
#520440000000
0!
0%
b110 *
0-
02
b110 6
#520450000000
1!
1%
1-
12
#520460000000
0!
0%
b111 *
0-
02
b111 6
#520470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#520480000000
0!
0%
b0 *
0-
02
b0 6
#520490000000
1!
1%
1-
12
#520500000000
0!
0%
b1 *
0-
02
b1 6
#520510000000
1!
1%
1-
12
#520520000000
0!
0%
b10 *
0-
02
b10 6
#520530000000
1!
1%
1-
12
#520540000000
0!
0%
b11 *
0-
02
b11 6
#520550000000
1!
1%
1-
12
15
#520560000000
0!
0%
b100 *
0-
02
b100 6
#520570000000
1!
1%
1-
12
#520580000000
0!
0%
b101 *
0-
02
b101 6
#520590000000
1!
1%
1-
12
#520600000000
0!
0%
b110 *
0-
02
b110 6
#520610000000
1!
1%
1-
12
#520620000000
0!
0%
b111 *
0-
02
b111 6
#520630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#520640000000
0!
0%
b0 *
0-
02
b0 6
#520650000000
1!
1%
1-
12
#520660000000
0!
0%
b1 *
0-
02
b1 6
#520670000000
1!
1%
1-
12
#520680000000
0!
0%
b10 *
0-
02
b10 6
#520690000000
1!
1%
1-
12
#520700000000
0!
0%
b11 *
0-
02
b11 6
#520710000000
1!
1%
1-
12
15
#520720000000
0!
0%
b100 *
0-
02
b100 6
#520730000000
1!
1%
1-
12
#520740000000
0!
0%
b101 *
0-
02
b101 6
#520750000000
1!
1%
1-
12
#520760000000
0!
0%
b110 *
0-
02
b110 6
#520770000000
1!
1%
1-
12
#520780000000
0!
0%
b111 *
0-
02
b111 6
#520790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#520800000000
0!
0%
b0 *
0-
02
b0 6
#520810000000
1!
1%
1-
12
#520820000000
0!
0%
b1 *
0-
02
b1 6
#520830000000
1!
1%
1-
12
#520840000000
0!
0%
b10 *
0-
02
b10 6
#520850000000
1!
1%
1-
12
#520860000000
0!
0%
b11 *
0-
02
b11 6
#520870000000
1!
1%
1-
12
15
#520880000000
0!
0%
b100 *
0-
02
b100 6
#520890000000
1!
1%
1-
12
#520900000000
0!
0%
b101 *
0-
02
b101 6
#520910000000
1!
1%
1-
12
#520920000000
0!
0%
b110 *
0-
02
b110 6
#520930000000
1!
1%
1-
12
#520940000000
0!
0%
b111 *
0-
02
b111 6
#520950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#520960000000
0!
0%
b0 *
0-
02
b0 6
#520970000000
1!
1%
1-
12
#520980000000
0!
0%
b1 *
0-
02
b1 6
#520990000000
1!
1%
1-
12
#521000000000
0!
0%
b10 *
0-
02
b10 6
#521010000000
1!
1%
1-
12
#521020000000
0!
0%
b11 *
0-
02
b11 6
#521030000000
1!
1%
1-
12
15
#521040000000
0!
0%
b100 *
0-
02
b100 6
#521050000000
1!
1%
1-
12
#521060000000
0!
0%
b101 *
0-
02
b101 6
#521070000000
1!
1%
1-
12
#521080000000
0!
0%
b110 *
0-
02
b110 6
#521090000000
1!
1%
1-
12
#521100000000
0!
0%
b111 *
0-
02
b111 6
#521110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#521120000000
0!
0%
b0 *
0-
02
b0 6
#521130000000
1!
1%
1-
12
#521140000000
0!
0%
b1 *
0-
02
b1 6
#521150000000
1!
1%
1-
12
#521160000000
0!
0%
b10 *
0-
02
b10 6
#521170000000
1!
1%
1-
12
#521180000000
0!
0%
b11 *
0-
02
b11 6
#521190000000
1!
1%
1-
12
15
#521200000000
0!
0%
b100 *
0-
02
b100 6
#521210000000
1!
1%
1-
12
#521220000000
0!
0%
b101 *
0-
02
b101 6
#521230000000
1!
1%
1-
12
#521240000000
0!
0%
b110 *
0-
02
b110 6
#521250000000
1!
1%
1-
12
#521260000000
0!
0%
b111 *
0-
02
b111 6
#521270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#521280000000
0!
0%
b0 *
0-
02
b0 6
#521290000000
1!
1%
1-
12
#521300000000
0!
0%
b1 *
0-
02
b1 6
#521310000000
1!
1%
1-
12
#521320000000
0!
0%
b10 *
0-
02
b10 6
#521330000000
1!
1%
1-
12
#521340000000
0!
0%
b11 *
0-
02
b11 6
#521350000000
1!
1%
1-
12
15
#521360000000
0!
0%
b100 *
0-
02
b100 6
#521370000000
1!
1%
1-
12
#521380000000
0!
0%
b101 *
0-
02
b101 6
#521390000000
1!
1%
1-
12
#521400000000
0!
0%
b110 *
0-
02
b110 6
#521410000000
1!
1%
1-
12
#521420000000
0!
0%
b111 *
0-
02
b111 6
#521430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#521440000000
0!
0%
b0 *
0-
02
b0 6
#521450000000
1!
1%
1-
12
#521460000000
0!
0%
b1 *
0-
02
b1 6
#521470000000
1!
1%
1-
12
#521480000000
0!
0%
b10 *
0-
02
b10 6
#521490000000
1!
1%
1-
12
#521500000000
0!
0%
b11 *
0-
02
b11 6
#521510000000
1!
1%
1-
12
15
#521520000000
0!
0%
b100 *
0-
02
b100 6
#521530000000
1!
1%
1-
12
#521540000000
0!
0%
b101 *
0-
02
b101 6
#521550000000
1!
1%
1-
12
#521560000000
0!
0%
b110 *
0-
02
b110 6
#521570000000
1!
1%
1-
12
#521580000000
0!
0%
b111 *
0-
02
b111 6
#521590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#521600000000
0!
0%
b0 *
0-
02
b0 6
#521610000000
1!
1%
1-
12
#521620000000
0!
0%
b1 *
0-
02
b1 6
#521630000000
1!
1%
1-
12
#521640000000
0!
0%
b10 *
0-
02
b10 6
#521650000000
1!
1%
1-
12
#521660000000
0!
0%
b11 *
0-
02
b11 6
#521670000000
1!
1%
1-
12
15
#521680000000
0!
0%
b100 *
0-
02
b100 6
#521690000000
1!
1%
1-
12
#521700000000
0!
0%
b101 *
0-
02
b101 6
#521710000000
1!
1%
1-
12
#521720000000
0!
0%
b110 *
0-
02
b110 6
#521730000000
1!
1%
1-
12
#521740000000
0!
0%
b111 *
0-
02
b111 6
#521750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#521760000000
0!
0%
b0 *
0-
02
b0 6
#521770000000
1!
1%
1-
12
#521780000000
0!
0%
b1 *
0-
02
b1 6
#521790000000
1!
1%
1-
12
#521800000000
0!
0%
b10 *
0-
02
b10 6
#521810000000
1!
1%
1-
12
#521820000000
0!
0%
b11 *
0-
02
b11 6
#521830000000
1!
1%
1-
12
15
#521840000000
0!
0%
b100 *
0-
02
b100 6
#521850000000
1!
1%
1-
12
#521860000000
0!
0%
b101 *
0-
02
b101 6
#521870000000
1!
1%
1-
12
#521880000000
0!
0%
b110 *
0-
02
b110 6
#521890000000
1!
1%
1-
12
#521900000000
0!
0%
b111 *
0-
02
b111 6
#521910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#521920000000
0!
0%
b0 *
0-
02
b0 6
#521930000000
1!
1%
1-
12
#521940000000
0!
0%
b1 *
0-
02
b1 6
#521950000000
1!
1%
1-
12
#521960000000
0!
0%
b10 *
0-
02
b10 6
#521970000000
1!
1%
1-
12
#521980000000
0!
0%
b11 *
0-
02
b11 6
#521990000000
1!
1%
1-
12
15
#522000000000
0!
0%
b100 *
0-
02
b100 6
#522010000000
1!
1%
1-
12
#522020000000
0!
0%
b101 *
0-
02
b101 6
#522030000000
1!
1%
1-
12
#522040000000
0!
0%
b110 *
0-
02
b110 6
#522050000000
1!
1%
1-
12
#522060000000
0!
0%
b111 *
0-
02
b111 6
#522070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#522080000000
0!
0%
b0 *
0-
02
b0 6
#522090000000
1!
1%
1-
12
#522100000000
0!
0%
b1 *
0-
02
b1 6
#522110000000
1!
1%
1-
12
#522120000000
0!
0%
b10 *
0-
02
b10 6
#522130000000
1!
1%
1-
12
#522140000000
0!
0%
b11 *
0-
02
b11 6
#522150000000
1!
1%
1-
12
15
#522160000000
0!
0%
b100 *
0-
02
b100 6
#522170000000
1!
1%
1-
12
#522180000000
0!
0%
b101 *
0-
02
b101 6
#522190000000
1!
1%
1-
12
#522200000000
0!
0%
b110 *
0-
02
b110 6
#522210000000
1!
1%
1-
12
#522220000000
0!
0%
b111 *
0-
02
b111 6
#522230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#522240000000
0!
0%
b0 *
0-
02
b0 6
#522250000000
1!
1%
1-
12
#522260000000
0!
0%
b1 *
0-
02
b1 6
#522270000000
1!
1%
1-
12
#522280000000
0!
0%
b10 *
0-
02
b10 6
#522290000000
1!
1%
1-
12
#522300000000
0!
0%
b11 *
0-
02
b11 6
#522310000000
1!
1%
1-
12
15
#522320000000
0!
0%
b100 *
0-
02
b100 6
#522330000000
1!
1%
1-
12
#522340000000
0!
0%
b101 *
0-
02
b101 6
#522350000000
1!
1%
1-
12
#522360000000
0!
0%
b110 *
0-
02
b110 6
#522370000000
1!
1%
1-
12
#522380000000
0!
0%
b111 *
0-
02
b111 6
#522390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#522400000000
0!
0%
b0 *
0-
02
b0 6
#522410000000
1!
1%
1-
12
#522420000000
0!
0%
b1 *
0-
02
b1 6
#522430000000
1!
1%
1-
12
#522440000000
0!
0%
b10 *
0-
02
b10 6
#522450000000
1!
1%
1-
12
#522460000000
0!
0%
b11 *
0-
02
b11 6
#522470000000
1!
1%
1-
12
15
#522480000000
0!
0%
b100 *
0-
02
b100 6
#522490000000
1!
1%
1-
12
#522500000000
0!
0%
b101 *
0-
02
b101 6
#522510000000
1!
1%
1-
12
#522520000000
0!
0%
b110 *
0-
02
b110 6
#522530000000
1!
1%
1-
12
#522540000000
0!
0%
b111 *
0-
02
b111 6
#522550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#522560000000
0!
0%
b0 *
0-
02
b0 6
#522570000000
1!
1%
1-
12
#522580000000
0!
0%
b1 *
0-
02
b1 6
#522590000000
1!
1%
1-
12
#522600000000
0!
0%
b10 *
0-
02
b10 6
#522610000000
1!
1%
1-
12
#522620000000
0!
0%
b11 *
0-
02
b11 6
#522630000000
1!
1%
1-
12
15
#522640000000
0!
0%
b100 *
0-
02
b100 6
#522650000000
1!
1%
1-
12
#522660000000
0!
0%
b101 *
0-
02
b101 6
#522670000000
1!
1%
1-
12
#522680000000
0!
0%
b110 *
0-
02
b110 6
#522690000000
1!
1%
1-
12
#522700000000
0!
0%
b111 *
0-
02
b111 6
#522710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#522720000000
0!
0%
b0 *
0-
02
b0 6
#522730000000
1!
1%
1-
12
#522740000000
0!
0%
b1 *
0-
02
b1 6
#522750000000
1!
1%
1-
12
#522760000000
0!
0%
b10 *
0-
02
b10 6
#522770000000
1!
1%
1-
12
#522780000000
0!
0%
b11 *
0-
02
b11 6
#522790000000
1!
1%
1-
12
15
#522800000000
0!
0%
b100 *
0-
02
b100 6
#522810000000
1!
1%
1-
12
#522820000000
0!
0%
b101 *
0-
02
b101 6
#522830000000
1!
1%
1-
12
#522840000000
0!
0%
b110 *
0-
02
b110 6
#522850000000
1!
1%
1-
12
#522860000000
0!
0%
b111 *
0-
02
b111 6
#522870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#522880000000
0!
0%
b0 *
0-
02
b0 6
#522890000000
1!
1%
1-
12
#522900000000
0!
0%
b1 *
0-
02
b1 6
#522910000000
1!
1%
1-
12
#522920000000
0!
0%
b10 *
0-
02
b10 6
#522930000000
1!
1%
1-
12
#522940000000
0!
0%
b11 *
0-
02
b11 6
#522950000000
1!
1%
1-
12
15
#522960000000
0!
0%
b100 *
0-
02
b100 6
#522970000000
1!
1%
1-
12
#522980000000
0!
0%
b101 *
0-
02
b101 6
#522990000000
1!
1%
1-
12
#523000000000
0!
0%
b110 *
0-
02
b110 6
#523010000000
1!
1%
1-
12
#523020000000
0!
0%
b111 *
0-
02
b111 6
#523030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#523040000000
0!
0%
b0 *
0-
02
b0 6
#523050000000
1!
1%
1-
12
#523060000000
0!
0%
b1 *
0-
02
b1 6
#523070000000
1!
1%
1-
12
#523080000000
0!
0%
b10 *
0-
02
b10 6
#523090000000
1!
1%
1-
12
#523100000000
0!
0%
b11 *
0-
02
b11 6
#523110000000
1!
1%
1-
12
15
#523120000000
0!
0%
b100 *
0-
02
b100 6
#523130000000
1!
1%
1-
12
#523140000000
0!
0%
b101 *
0-
02
b101 6
#523150000000
1!
1%
1-
12
#523160000000
0!
0%
b110 *
0-
02
b110 6
#523170000000
1!
1%
1-
12
#523180000000
0!
0%
b111 *
0-
02
b111 6
#523190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#523200000000
0!
0%
b0 *
0-
02
b0 6
#523210000000
1!
1%
1-
12
#523220000000
0!
0%
b1 *
0-
02
b1 6
#523230000000
1!
1%
1-
12
#523240000000
0!
0%
b10 *
0-
02
b10 6
#523250000000
1!
1%
1-
12
#523260000000
0!
0%
b11 *
0-
02
b11 6
#523270000000
1!
1%
1-
12
15
#523280000000
0!
0%
b100 *
0-
02
b100 6
#523290000000
1!
1%
1-
12
#523300000000
0!
0%
b101 *
0-
02
b101 6
#523310000000
1!
1%
1-
12
#523320000000
0!
0%
b110 *
0-
02
b110 6
#523330000000
1!
1%
1-
12
#523340000000
0!
0%
b111 *
0-
02
b111 6
#523350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#523360000000
0!
0%
b0 *
0-
02
b0 6
#523370000000
1!
1%
1-
12
#523380000000
0!
0%
b1 *
0-
02
b1 6
#523390000000
1!
1%
1-
12
#523400000000
0!
0%
b10 *
0-
02
b10 6
#523410000000
1!
1%
1-
12
#523420000000
0!
0%
b11 *
0-
02
b11 6
#523430000000
1!
1%
1-
12
15
#523440000000
0!
0%
b100 *
0-
02
b100 6
#523450000000
1!
1%
1-
12
#523460000000
0!
0%
b101 *
0-
02
b101 6
#523470000000
1!
1%
1-
12
#523480000000
0!
0%
b110 *
0-
02
b110 6
#523490000000
1!
1%
1-
12
#523500000000
0!
0%
b111 *
0-
02
b111 6
#523510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#523520000000
0!
0%
b0 *
0-
02
b0 6
#523530000000
1!
1%
1-
12
#523540000000
0!
0%
b1 *
0-
02
b1 6
#523550000000
1!
1%
1-
12
#523560000000
0!
0%
b10 *
0-
02
b10 6
#523570000000
1!
1%
1-
12
#523580000000
0!
0%
b11 *
0-
02
b11 6
#523590000000
1!
1%
1-
12
15
#523600000000
0!
0%
b100 *
0-
02
b100 6
#523610000000
1!
1%
1-
12
#523620000000
0!
0%
b101 *
0-
02
b101 6
#523630000000
1!
1%
1-
12
#523640000000
0!
0%
b110 *
0-
02
b110 6
#523650000000
1!
1%
1-
12
#523660000000
0!
0%
b111 *
0-
02
b111 6
#523670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#523680000000
0!
0%
b0 *
0-
02
b0 6
#523690000000
1!
1%
1-
12
#523700000000
0!
0%
b1 *
0-
02
b1 6
#523710000000
1!
1%
1-
12
#523720000000
0!
0%
b10 *
0-
02
b10 6
#523730000000
1!
1%
1-
12
#523740000000
0!
0%
b11 *
0-
02
b11 6
#523750000000
1!
1%
1-
12
15
#523760000000
0!
0%
b100 *
0-
02
b100 6
#523770000000
1!
1%
1-
12
#523780000000
0!
0%
b101 *
0-
02
b101 6
#523790000000
1!
1%
1-
12
#523800000000
0!
0%
b110 *
0-
02
b110 6
#523810000000
1!
1%
1-
12
#523820000000
0!
0%
b111 *
0-
02
b111 6
#523830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#523840000000
0!
0%
b0 *
0-
02
b0 6
#523850000000
1!
1%
1-
12
#523860000000
0!
0%
b1 *
0-
02
b1 6
#523870000000
1!
1%
1-
12
#523880000000
0!
0%
b10 *
0-
02
b10 6
#523890000000
1!
1%
1-
12
#523900000000
0!
0%
b11 *
0-
02
b11 6
#523910000000
1!
1%
1-
12
15
#523920000000
0!
0%
b100 *
0-
02
b100 6
#523930000000
1!
1%
1-
12
#523940000000
0!
0%
b101 *
0-
02
b101 6
#523950000000
1!
1%
1-
12
#523960000000
0!
0%
b110 *
0-
02
b110 6
#523970000000
1!
1%
1-
12
#523980000000
0!
0%
b111 *
0-
02
b111 6
#523990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#524000000000
0!
0%
b0 *
0-
02
b0 6
#524010000000
1!
1%
1-
12
#524020000000
0!
0%
b1 *
0-
02
b1 6
#524030000000
1!
1%
1-
12
#524040000000
0!
0%
b10 *
0-
02
b10 6
#524050000000
1!
1%
1-
12
#524060000000
0!
0%
b11 *
0-
02
b11 6
#524070000000
1!
1%
1-
12
15
#524080000000
0!
0%
b100 *
0-
02
b100 6
#524090000000
1!
1%
1-
12
#524100000000
0!
0%
b101 *
0-
02
b101 6
#524110000000
1!
1%
1-
12
#524120000000
0!
0%
b110 *
0-
02
b110 6
#524130000000
1!
1%
1-
12
#524140000000
0!
0%
b111 *
0-
02
b111 6
#524150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#524160000000
0!
0%
b0 *
0-
02
b0 6
#524170000000
1!
1%
1-
12
#524180000000
0!
0%
b1 *
0-
02
b1 6
#524190000000
1!
1%
1-
12
#524200000000
0!
0%
b10 *
0-
02
b10 6
#524210000000
1!
1%
1-
12
#524220000000
0!
0%
b11 *
0-
02
b11 6
#524230000000
1!
1%
1-
12
15
#524240000000
0!
0%
b100 *
0-
02
b100 6
#524250000000
1!
1%
1-
12
#524260000000
0!
0%
b101 *
0-
02
b101 6
#524270000000
1!
1%
1-
12
#524280000000
0!
0%
b110 *
0-
02
b110 6
#524290000000
1!
1%
1-
12
#524300000000
0!
0%
b111 *
0-
02
b111 6
#524310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#524320000000
0!
0%
b0 *
0-
02
b0 6
#524330000000
1!
1%
1-
12
#524340000000
0!
0%
b1 *
0-
02
b1 6
#524350000000
1!
1%
1-
12
#524360000000
0!
0%
b10 *
0-
02
b10 6
#524370000000
1!
1%
1-
12
#524380000000
0!
0%
b11 *
0-
02
b11 6
#524390000000
1!
1%
1-
12
15
#524400000000
0!
0%
b100 *
0-
02
b100 6
#524410000000
1!
1%
1-
12
#524420000000
0!
0%
b101 *
0-
02
b101 6
#524430000000
1!
1%
1-
12
#524440000000
0!
0%
b110 *
0-
02
b110 6
#524450000000
1!
1%
1-
12
#524460000000
0!
0%
b111 *
0-
02
b111 6
#524470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#524480000000
0!
0%
b0 *
0-
02
b0 6
#524490000000
1!
1%
1-
12
#524500000000
0!
0%
b1 *
0-
02
b1 6
#524510000000
1!
1%
1-
12
#524520000000
0!
0%
b10 *
0-
02
b10 6
#524530000000
1!
1%
1-
12
#524540000000
0!
0%
b11 *
0-
02
b11 6
#524550000000
1!
1%
1-
12
15
#524560000000
0!
0%
b100 *
0-
02
b100 6
#524570000000
1!
1%
1-
12
#524580000000
0!
0%
b101 *
0-
02
b101 6
#524590000000
1!
1%
1-
12
#524600000000
0!
0%
b110 *
0-
02
b110 6
#524610000000
1!
1%
1-
12
#524620000000
0!
0%
b111 *
0-
02
b111 6
#524630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#524640000000
0!
0%
b0 *
0-
02
b0 6
#524650000000
1!
1%
1-
12
#524660000000
0!
0%
b1 *
0-
02
b1 6
#524670000000
1!
1%
1-
12
#524680000000
0!
0%
b10 *
0-
02
b10 6
#524690000000
1!
1%
1-
12
#524700000000
0!
0%
b11 *
0-
02
b11 6
#524710000000
1!
1%
1-
12
15
#524720000000
0!
0%
b100 *
0-
02
b100 6
#524730000000
1!
1%
1-
12
#524740000000
0!
0%
b101 *
0-
02
b101 6
#524750000000
1!
1%
1-
12
#524760000000
0!
0%
b110 *
0-
02
b110 6
#524770000000
1!
1%
1-
12
#524780000000
0!
0%
b111 *
0-
02
b111 6
#524790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#524800000000
0!
0%
b0 *
0-
02
b0 6
#524810000000
1!
1%
1-
12
#524820000000
0!
0%
b1 *
0-
02
b1 6
#524830000000
1!
1%
1-
12
#524840000000
0!
0%
b10 *
0-
02
b10 6
#524850000000
1!
1%
1-
12
#524860000000
0!
0%
b11 *
0-
02
b11 6
#524870000000
1!
1%
1-
12
15
#524880000000
0!
0%
b100 *
0-
02
b100 6
#524890000000
1!
1%
1-
12
#524900000000
0!
0%
b101 *
0-
02
b101 6
#524910000000
1!
1%
1-
12
#524920000000
0!
0%
b110 *
0-
02
b110 6
#524930000000
1!
1%
1-
12
#524940000000
0!
0%
b111 *
0-
02
b111 6
#524950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#524960000000
0!
0%
b0 *
0-
02
b0 6
#524970000000
1!
1%
1-
12
#524980000000
0!
0%
b1 *
0-
02
b1 6
#524990000000
1!
1%
1-
12
#525000000000
0!
0%
b10 *
0-
02
b10 6
#525010000000
1!
1%
1-
12
#525020000000
0!
0%
b11 *
0-
02
b11 6
#525030000000
1!
1%
1-
12
15
#525040000000
0!
0%
b100 *
0-
02
b100 6
#525050000000
1!
1%
1-
12
#525060000000
0!
0%
b101 *
0-
02
b101 6
#525070000000
1!
1%
1-
12
#525080000000
0!
0%
b110 *
0-
02
b110 6
#525090000000
1!
1%
1-
12
#525100000000
0!
0%
b111 *
0-
02
b111 6
#525110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#525120000000
0!
0%
b0 *
0-
02
b0 6
#525130000000
1!
1%
1-
12
#525140000000
0!
0%
b1 *
0-
02
b1 6
#525150000000
1!
1%
1-
12
#525160000000
0!
0%
b10 *
0-
02
b10 6
#525170000000
1!
1%
1-
12
#525180000000
0!
0%
b11 *
0-
02
b11 6
#525190000000
1!
1%
1-
12
15
#525200000000
0!
0%
b100 *
0-
02
b100 6
#525210000000
1!
1%
1-
12
#525220000000
0!
0%
b101 *
0-
02
b101 6
#525230000000
1!
1%
1-
12
#525240000000
0!
0%
b110 *
0-
02
b110 6
#525250000000
1!
1%
1-
12
#525260000000
0!
0%
b111 *
0-
02
b111 6
#525270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#525280000000
0!
0%
b0 *
0-
02
b0 6
#525290000000
1!
1%
1-
12
#525300000000
0!
0%
b1 *
0-
02
b1 6
#525310000000
1!
1%
1-
12
#525320000000
0!
0%
b10 *
0-
02
b10 6
#525330000000
1!
1%
1-
12
#525340000000
0!
0%
b11 *
0-
02
b11 6
#525350000000
1!
1%
1-
12
15
#525360000000
0!
0%
b100 *
0-
02
b100 6
#525370000000
1!
1%
1-
12
#525380000000
0!
0%
b101 *
0-
02
b101 6
#525390000000
1!
1%
1-
12
#525400000000
0!
0%
b110 *
0-
02
b110 6
#525410000000
1!
1%
1-
12
#525420000000
0!
0%
b111 *
0-
02
b111 6
#525430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#525440000000
0!
0%
b0 *
0-
02
b0 6
#525450000000
1!
1%
1-
12
#525460000000
0!
0%
b1 *
0-
02
b1 6
#525470000000
1!
1%
1-
12
#525480000000
0!
0%
b10 *
0-
02
b10 6
#525490000000
1!
1%
1-
12
#525500000000
0!
0%
b11 *
0-
02
b11 6
#525510000000
1!
1%
1-
12
15
#525520000000
0!
0%
b100 *
0-
02
b100 6
#525530000000
1!
1%
1-
12
#525540000000
0!
0%
b101 *
0-
02
b101 6
#525550000000
1!
1%
1-
12
#525560000000
0!
0%
b110 *
0-
02
b110 6
#525570000000
1!
1%
1-
12
#525580000000
0!
0%
b111 *
0-
02
b111 6
#525590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#525600000000
0!
0%
b0 *
0-
02
b0 6
#525610000000
1!
1%
1-
12
#525620000000
0!
0%
b1 *
0-
02
b1 6
#525630000000
1!
1%
1-
12
#525640000000
0!
0%
b10 *
0-
02
b10 6
#525650000000
1!
1%
1-
12
#525660000000
0!
0%
b11 *
0-
02
b11 6
#525670000000
1!
1%
1-
12
15
#525680000000
0!
0%
b100 *
0-
02
b100 6
#525690000000
1!
1%
1-
12
#525700000000
0!
0%
b101 *
0-
02
b101 6
#525710000000
1!
1%
1-
12
#525720000000
0!
0%
b110 *
0-
02
b110 6
#525730000000
1!
1%
1-
12
#525740000000
0!
0%
b111 *
0-
02
b111 6
#525750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#525760000000
0!
0%
b0 *
0-
02
b0 6
#525770000000
1!
1%
1-
12
#525780000000
0!
0%
b1 *
0-
02
b1 6
#525790000000
1!
1%
1-
12
#525800000000
0!
0%
b10 *
0-
02
b10 6
#525810000000
1!
1%
1-
12
#525820000000
0!
0%
b11 *
0-
02
b11 6
#525830000000
1!
1%
1-
12
15
#525840000000
0!
0%
b100 *
0-
02
b100 6
#525850000000
1!
1%
1-
12
#525860000000
0!
0%
b101 *
0-
02
b101 6
#525870000000
1!
1%
1-
12
#525880000000
0!
0%
b110 *
0-
02
b110 6
#525890000000
1!
1%
1-
12
#525900000000
0!
0%
b111 *
0-
02
b111 6
#525910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#525920000000
0!
0%
b0 *
0-
02
b0 6
#525930000000
1!
1%
1-
12
#525940000000
0!
0%
b1 *
0-
02
b1 6
#525950000000
1!
1%
1-
12
#525960000000
0!
0%
b10 *
0-
02
b10 6
#525970000000
1!
1%
1-
12
#525980000000
0!
0%
b11 *
0-
02
b11 6
#525990000000
1!
1%
1-
12
15
#526000000000
0!
0%
b100 *
0-
02
b100 6
#526010000000
1!
1%
1-
12
#526020000000
0!
0%
b101 *
0-
02
b101 6
#526030000000
1!
1%
1-
12
#526040000000
0!
0%
b110 *
0-
02
b110 6
#526050000000
1!
1%
1-
12
#526060000000
0!
0%
b111 *
0-
02
b111 6
#526070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#526080000000
0!
0%
b0 *
0-
02
b0 6
#526090000000
1!
1%
1-
12
#526100000000
0!
0%
b1 *
0-
02
b1 6
#526110000000
1!
1%
1-
12
#526120000000
0!
0%
b10 *
0-
02
b10 6
#526130000000
1!
1%
1-
12
#526140000000
0!
0%
b11 *
0-
02
b11 6
#526150000000
1!
1%
1-
12
15
#526160000000
0!
0%
b100 *
0-
02
b100 6
#526170000000
1!
1%
1-
12
#526180000000
0!
0%
b101 *
0-
02
b101 6
#526190000000
1!
1%
1-
12
#526200000000
0!
0%
b110 *
0-
02
b110 6
#526210000000
1!
1%
1-
12
#526220000000
0!
0%
b111 *
0-
02
b111 6
#526230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#526240000000
0!
0%
b0 *
0-
02
b0 6
#526250000000
1!
1%
1-
12
#526260000000
0!
0%
b1 *
0-
02
b1 6
#526270000000
1!
1%
1-
12
#526280000000
0!
0%
b10 *
0-
02
b10 6
#526290000000
1!
1%
1-
12
#526300000000
0!
0%
b11 *
0-
02
b11 6
#526310000000
1!
1%
1-
12
15
#526320000000
0!
0%
b100 *
0-
02
b100 6
#526330000000
1!
1%
1-
12
#526340000000
0!
0%
b101 *
0-
02
b101 6
#526350000000
1!
1%
1-
12
#526360000000
0!
0%
b110 *
0-
02
b110 6
#526370000000
1!
1%
1-
12
#526380000000
0!
0%
b111 *
0-
02
b111 6
#526390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#526400000000
0!
0%
b0 *
0-
02
b0 6
#526410000000
1!
1%
1-
12
#526420000000
0!
0%
b1 *
0-
02
b1 6
#526430000000
1!
1%
1-
12
#526440000000
0!
0%
b10 *
0-
02
b10 6
#526450000000
1!
1%
1-
12
#526460000000
0!
0%
b11 *
0-
02
b11 6
#526470000000
1!
1%
1-
12
15
#526480000000
0!
0%
b100 *
0-
02
b100 6
#526490000000
1!
1%
1-
12
#526500000000
0!
0%
b101 *
0-
02
b101 6
#526510000000
1!
1%
1-
12
#526520000000
0!
0%
b110 *
0-
02
b110 6
#526530000000
1!
1%
1-
12
#526540000000
0!
0%
b111 *
0-
02
b111 6
#526550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#526560000000
0!
0%
b0 *
0-
02
b0 6
#526570000000
1!
1%
1-
12
#526580000000
0!
0%
b1 *
0-
02
b1 6
#526590000000
1!
1%
1-
12
#526600000000
0!
0%
b10 *
0-
02
b10 6
#526610000000
1!
1%
1-
12
#526620000000
0!
0%
b11 *
0-
02
b11 6
#526630000000
1!
1%
1-
12
15
#526640000000
0!
0%
b100 *
0-
02
b100 6
#526650000000
1!
1%
1-
12
#526660000000
0!
0%
b101 *
0-
02
b101 6
#526670000000
1!
1%
1-
12
#526680000000
0!
0%
b110 *
0-
02
b110 6
#526690000000
1!
1%
1-
12
#526700000000
0!
0%
b111 *
0-
02
b111 6
#526710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#526720000000
0!
0%
b0 *
0-
02
b0 6
#526730000000
1!
1%
1-
12
#526740000000
0!
0%
b1 *
0-
02
b1 6
#526750000000
1!
1%
1-
12
#526760000000
0!
0%
b10 *
0-
02
b10 6
#526770000000
1!
1%
1-
12
#526780000000
0!
0%
b11 *
0-
02
b11 6
#526790000000
1!
1%
1-
12
15
#526800000000
0!
0%
b100 *
0-
02
b100 6
#526810000000
1!
1%
1-
12
#526820000000
0!
0%
b101 *
0-
02
b101 6
#526830000000
1!
1%
1-
12
#526840000000
0!
0%
b110 *
0-
02
b110 6
#526850000000
1!
1%
1-
12
#526860000000
0!
0%
b111 *
0-
02
b111 6
#526870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#526880000000
0!
0%
b0 *
0-
02
b0 6
#526890000000
1!
1%
1-
12
#526900000000
0!
0%
b1 *
0-
02
b1 6
#526910000000
1!
1%
1-
12
#526920000000
0!
0%
b10 *
0-
02
b10 6
#526930000000
1!
1%
1-
12
#526940000000
0!
0%
b11 *
0-
02
b11 6
#526950000000
1!
1%
1-
12
15
#526960000000
0!
0%
b100 *
0-
02
b100 6
#526970000000
1!
1%
1-
12
#526980000000
0!
0%
b101 *
0-
02
b101 6
#526990000000
1!
1%
1-
12
#527000000000
0!
0%
b110 *
0-
02
b110 6
#527010000000
1!
1%
1-
12
#527020000000
0!
0%
b111 *
0-
02
b111 6
#527030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#527040000000
0!
0%
b0 *
0-
02
b0 6
#527050000000
1!
1%
1-
12
#527060000000
0!
0%
b1 *
0-
02
b1 6
#527070000000
1!
1%
1-
12
#527080000000
0!
0%
b10 *
0-
02
b10 6
#527090000000
1!
1%
1-
12
#527100000000
0!
0%
b11 *
0-
02
b11 6
#527110000000
1!
1%
1-
12
15
#527120000000
0!
0%
b100 *
0-
02
b100 6
#527130000000
1!
1%
1-
12
#527140000000
0!
0%
b101 *
0-
02
b101 6
#527150000000
1!
1%
1-
12
#527160000000
0!
0%
b110 *
0-
02
b110 6
#527170000000
1!
1%
1-
12
#527180000000
0!
0%
b111 *
0-
02
b111 6
#527190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#527200000000
0!
0%
b0 *
0-
02
b0 6
#527210000000
1!
1%
1-
12
#527220000000
0!
0%
b1 *
0-
02
b1 6
#527230000000
1!
1%
1-
12
#527240000000
0!
0%
b10 *
0-
02
b10 6
#527250000000
1!
1%
1-
12
#527260000000
0!
0%
b11 *
0-
02
b11 6
#527270000000
1!
1%
1-
12
15
#527280000000
0!
0%
b100 *
0-
02
b100 6
#527290000000
1!
1%
1-
12
#527300000000
0!
0%
b101 *
0-
02
b101 6
#527310000000
1!
1%
1-
12
#527320000000
0!
0%
b110 *
0-
02
b110 6
#527330000000
1!
1%
1-
12
#527340000000
0!
0%
b111 *
0-
02
b111 6
#527350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#527360000000
0!
0%
b0 *
0-
02
b0 6
#527370000000
1!
1%
1-
12
#527380000000
0!
0%
b1 *
0-
02
b1 6
#527390000000
1!
1%
1-
12
#527400000000
0!
0%
b10 *
0-
02
b10 6
#527410000000
1!
1%
1-
12
#527420000000
0!
0%
b11 *
0-
02
b11 6
#527430000000
1!
1%
1-
12
15
#527440000000
0!
0%
b100 *
0-
02
b100 6
#527450000000
1!
1%
1-
12
#527460000000
0!
0%
b101 *
0-
02
b101 6
#527470000000
1!
1%
1-
12
#527480000000
0!
0%
b110 *
0-
02
b110 6
#527490000000
1!
1%
1-
12
#527500000000
0!
0%
b111 *
0-
02
b111 6
#527510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#527520000000
0!
0%
b0 *
0-
02
b0 6
#527530000000
1!
1%
1-
12
#527540000000
0!
0%
b1 *
0-
02
b1 6
#527550000000
1!
1%
1-
12
#527560000000
0!
0%
b10 *
0-
02
b10 6
#527570000000
1!
1%
1-
12
#527580000000
0!
0%
b11 *
0-
02
b11 6
#527590000000
1!
1%
1-
12
15
#527600000000
0!
0%
b100 *
0-
02
b100 6
#527610000000
1!
1%
1-
12
#527620000000
0!
0%
b101 *
0-
02
b101 6
#527630000000
1!
1%
1-
12
#527640000000
0!
0%
b110 *
0-
02
b110 6
#527650000000
1!
1%
1-
12
#527660000000
0!
0%
b111 *
0-
02
b111 6
#527670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#527680000000
0!
0%
b0 *
0-
02
b0 6
#527690000000
1!
1%
1-
12
#527700000000
0!
0%
b1 *
0-
02
b1 6
#527710000000
1!
1%
1-
12
#527720000000
0!
0%
b10 *
0-
02
b10 6
#527730000000
1!
1%
1-
12
#527740000000
0!
0%
b11 *
0-
02
b11 6
#527750000000
1!
1%
1-
12
15
#527760000000
0!
0%
b100 *
0-
02
b100 6
#527770000000
1!
1%
1-
12
#527780000000
0!
0%
b101 *
0-
02
b101 6
#527790000000
1!
1%
1-
12
#527800000000
0!
0%
b110 *
0-
02
b110 6
#527810000000
1!
1%
1-
12
#527820000000
0!
0%
b111 *
0-
02
b111 6
#527830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#527840000000
0!
0%
b0 *
0-
02
b0 6
#527850000000
1!
1%
1-
12
#527860000000
0!
0%
b1 *
0-
02
b1 6
#527870000000
1!
1%
1-
12
#527880000000
0!
0%
b10 *
0-
02
b10 6
#527890000000
1!
1%
1-
12
#527900000000
0!
0%
b11 *
0-
02
b11 6
#527910000000
1!
1%
1-
12
15
#527920000000
0!
0%
b100 *
0-
02
b100 6
#527930000000
1!
1%
1-
12
#527940000000
0!
0%
b101 *
0-
02
b101 6
#527950000000
1!
1%
1-
12
#527960000000
0!
0%
b110 *
0-
02
b110 6
#527970000000
1!
1%
1-
12
#527980000000
0!
0%
b111 *
0-
02
b111 6
#527990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#528000000000
0!
0%
b0 *
0-
02
b0 6
#528010000000
1!
1%
1-
12
#528020000000
0!
0%
b1 *
0-
02
b1 6
#528030000000
1!
1%
1-
12
#528040000000
0!
0%
b10 *
0-
02
b10 6
#528050000000
1!
1%
1-
12
#528060000000
0!
0%
b11 *
0-
02
b11 6
#528070000000
1!
1%
1-
12
15
#528080000000
0!
0%
b100 *
0-
02
b100 6
#528090000000
1!
1%
1-
12
#528100000000
0!
0%
b101 *
0-
02
b101 6
#528110000000
1!
1%
1-
12
#528120000000
0!
0%
b110 *
0-
02
b110 6
#528130000000
1!
1%
1-
12
#528140000000
0!
0%
b111 *
0-
02
b111 6
#528150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#528160000000
0!
0%
b0 *
0-
02
b0 6
#528170000000
1!
1%
1-
12
#528180000000
0!
0%
b1 *
0-
02
b1 6
#528190000000
1!
1%
1-
12
#528200000000
0!
0%
b10 *
0-
02
b10 6
#528210000000
1!
1%
1-
12
#528220000000
0!
0%
b11 *
0-
02
b11 6
#528230000000
1!
1%
1-
12
15
#528240000000
0!
0%
b100 *
0-
02
b100 6
#528250000000
1!
1%
1-
12
#528260000000
0!
0%
b101 *
0-
02
b101 6
#528270000000
1!
1%
1-
12
#528280000000
0!
0%
b110 *
0-
02
b110 6
#528290000000
1!
1%
1-
12
#528300000000
0!
0%
b111 *
0-
02
b111 6
#528310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#528320000000
0!
0%
b0 *
0-
02
b0 6
#528330000000
1!
1%
1-
12
#528340000000
0!
0%
b1 *
0-
02
b1 6
#528350000000
1!
1%
1-
12
#528360000000
0!
0%
b10 *
0-
02
b10 6
#528370000000
1!
1%
1-
12
#528380000000
0!
0%
b11 *
0-
02
b11 6
#528390000000
1!
1%
1-
12
15
#528400000000
0!
0%
b100 *
0-
02
b100 6
#528410000000
1!
1%
1-
12
#528420000000
0!
0%
b101 *
0-
02
b101 6
#528430000000
1!
1%
1-
12
#528440000000
0!
0%
b110 *
0-
02
b110 6
#528450000000
1!
1%
1-
12
#528460000000
0!
0%
b111 *
0-
02
b111 6
#528470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#528480000000
0!
0%
b0 *
0-
02
b0 6
#528490000000
1!
1%
1-
12
#528500000000
0!
0%
b1 *
0-
02
b1 6
#528510000000
1!
1%
1-
12
#528520000000
0!
0%
b10 *
0-
02
b10 6
#528530000000
1!
1%
1-
12
#528540000000
0!
0%
b11 *
0-
02
b11 6
#528550000000
1!
1%
1-
12
15
#528560000000
0!
0%
b100 *
0-
02
b100 6
#528570000000
1!
1%
1-
12
#528580000000
0!
0%
b101 *
0-
02
b101 6
#528590000000
1!
1%
1-
12
#528600000000
0!
0%
b110 *
0-
02
b110 6
#528610000000
1!
1%
1-
12
#528620000000
0!
0%
b111 *
0-
02
b111 6
#528630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#528640000000
0!
0%
b0 *
0-
02
b0 6
#528650000000
1!
1%
1-
12
#528660000000
0!
0%
b1 *
0-
02
b1 6
#528670000000
1!
1%
1-
12
#528680000000
0!
0%
b10 *
0-
02
b10 6
#528690000000
1!
1%
1-
12
#528700000000
0!
0%
b11 *
0-
02
b11 6
#528710000000
1!
1%
1-
12
15
#528720000000
0!
0%
b100 *
0-
02
b100 6
#528730000000
1!
1%
1-
12
#528740000000
0!
0%
b101 *
0-
02
b101 6
#528750000000
1!
1%
1-
12
#528760000000
0!
0%
b110 *
0-
02
b110 6
#528770000000
1!
1%
1-
12
#528780000000
0!
0%
b111 *
0-
02
b111 6
#528790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#528800000000
0!
0%
b0 *
0-
02
b0 6
#528810000000
1!
1%
1-
12
#528820000000
0!
0%
b1 *
0-
02
b1 6
#528830000000
1!
1%
1-
12
#528840000000
0!
0%
b10 *
0-
02
b10 6
#528850000000
1!
1%
1-
12
#528860000000
0!
0%
b11 *
0-
02
b11 6
#528870000000
1!
1%
1-
12
15
#528880000000
0!
0%
b100 *
0-
02
b100 6
#528890000000
1!
1%
1-
12
#528900000000
0!
0%
b101 *
0-
02
b101 6
#528910000000
1!
1%
1-
12
#528920000000
0!
0%
b110 *
0-
02
b110 6
#528930000000
1!
1%
1-
12
#528940000000
0!
0%
b111 *
0-
02
b111 6
#528950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#528960000000
0!
0%
b0 *
0-
02
b0 6
#528970000000
1!
1%
1-
12
#528980000000
0!
0%
b1 *
0-
02
b1 6
#528990000000
1!
1%
1-
12
#529000000000
0!
0%
b10 *
0-
02
b10 6
#529010000000
1!
1%
1-
12
#529020000000
0!
0%
b11 *
0-
02
b11 6
#529030000000
1!
1%
1-
12
15
#529040000000
0!
0%
b100 *
0-
02
b100 6
#529050000000
1!
1%
1-
12
#529060000000
0!
0%
b101 *
0-
02
b101 6
#529070000000
1!
1%
1-
12
#529080000000
0!
0%
b110 *
0-
02
b110 6
#529090000000
1!
1%
1-
12
#529100000000
0!
0%
b111 *
0-
02
b111 6
#529110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#529120000000
0!
0%
b0 *
0-
02
b0 6
#529130000000
1!
1%
1-
12
#529140000000
0!
0%
b1 *
0-
02
b1 6
#529150000000
1!
1%
1-
12
#529160000000
0!
0%
b10 *
0-
02
b10 6
#529170000000
1!
1%
1-
12
#529180000000
0!
0%
b11 *
0-
02
b11 6
#529190000000
1!
1%
1-
12
15
#529200000000
0!
0%
b100 *
0-
02
b100 6
#529210000000
1!
1%
1-
12
#529220000000
0!
0%
b101 *
0-
02
b101 6
#529230000000
1!
1%
1-
12
#529240000000
0!
0%
b110 *
0-
02
b110 6
#529250000000
1!
1%
1-
12
#529260000000
0!
0%
b111 *
0-
02
b111 6
#529270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#529280000000
0!
0%
b0 *
0-
02
b0 6
#529290000000
1!
1%
1-
12
#529300000000
0!
0%
b1 *
0-
02
b1 6
#529310000000
1!
1%
1-
12
#529320000000
0!
0%
b10 *
0-
02
b10 6
#529330000000
1!
1%
1-
12
#529340000000
0!
0%
b11 *
0-
02
b11 6
#529350000000
1!
1%
1-
12
15
#529360000000
0!
0%
b100 *
0-
02
b100 6
#529370000000
1!
1%
1-
12
#529380000000
0!
0%
b101 *
0-
02
b101 6
#529390000000
1!
1%
1-
12
#529400000000
0!
0%
b110 *
0-
02
b110 6
#529410000000
1!
1%
1-
12
#529420000000
0!
0%
b111 *
0-
02
b111 6
#529430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#529440000000
0!
0%
b0 *
0-
02
b0 6
#529450000000
1!
1%
1-
12
#529460000000
0!
0%
b1 *
0-
02
b1 6
#529470000000
1!
1%
1-
12
#529480000000
0!
0%
b10 *
0-
02
b10 6
#529490000000
1!
1%
1-
12
#529500000000
0!
0%
b11 *
0-
02
b11 6
#529510000000
1!
1%
1-
12
15
#529520000000
0!
0%
b100 *
0-
02
b100 6
#529530000000
1!
1%
1-
12
#529540000000
0!
0%
b101 *
0-
02
b101 6
#529550000000
1!
1%
1-
12
#529560000000
0!
0%
b110 *
0-
02
b110 6
#529570000000
1!
1%
1-
12
#529580000000
0!
0%
b111 *
0-
02
b111 6
#529590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#529600000000
0!
0%
b0 *
0-
02
b0 6
#529610000000
1!
1%
1-
12
#529620000000
0!
0%
b1 *
0-
02
b1 6
#529630000000
1!
1%
1-
12
#529640000000
0!
0%
b10 *
0-
02
b10 6
#529650000000
1!
1%
1-
12
#529660000000
0!
0%
b11 *
0-
02
b11 6
#529670000000
1!
1%
1-
12
15
#529680000000
0!
0%
b100 *
0-
02
b100 6
#529690000000
1!
1%
1-
12
#529700000000
0!
0%
b101 *
0-
02
b101 6
#529710000000
1!
1%
1-
12
#529720000000
0!
0%
b110 *
0-
02
b110 6
#529730000000
1!
1%
1-
12
#529740000000
0!
0%
b111 *
0-
02
b111 6
#529750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#529760000000
0!
0%
b0 *
0-
02
b0 6
#529770000000
1!
1%
1-
12
#529780000000
0!
0%
b1 *
0-
02
b1 6
#529790000000
1!
1%
1-
12
#529800000000
0!
0%
b10 *
0-
02
b10 6
#529810000000
1!
1%
1-
12
#529820000000
0!
0%
b11 *
0-
02
b11 6
#529830000000
1!
1%
1-
12
15
#529840000000
0!
0%
b100 *
0-
02
b100 6
#529850000000
1!
1%
1-
12
#529860000000
0!
0%
b101 *
0-
02
b101 6
#529870000000
1!
1%
1-
12
#529880000000
0!
0%
b110 *
0-
02
b110 6
#529890000000
1!
1%
1-
12
#529900000000
0!
0%
b111 *
0-
02
b111 6
#529910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#529920000000
0!
0%
b0 *
0-
02
b0 6
#529930000000
1!
1%
1-
12
#529940000000
0!
0%
b1 *
0-
02
b1 6
#529950000000
1!
1%
1-
12
#529960000000
0!
0%
b10 *
0-
02
b10 6
#529970000000
1!
1%
1-
12
#529980000000
0!
0%
b11 *
0-
02
b11 6
#529990000000
1!
1%
1-
12
15
#530000000000
0!
0%
b100 *
0-
02
b100 6
#530010000000
1!
1%
1-
12
#530020000000
0!
0%
b101 *
0-
02
b101 6
#530030000000
1!
1%
1-
12
#530040000000
0!
0%
b110 *
0-
02
b110 6
#530050000000
1!
1%
1-
12
#530060000000
0!
0%
b111 *
0-
02
b111 6
#530070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#530080000000
0!
0%
b0 *
0-
02
b0 6
#530090000000
1!
1%
1-
12
#530100000000
0!
0%
b1 *
0-
02
b1 6
#530110000000
1!
1%
1-
12
#530120000000
0!
0%
b10 *
0-
02
b10 6
#530130000000
1!
1%
1-
12
#530140000000
0!
0%
b11 *
0-
02
b11 6
#530150000000
1!
1%
1-
12
15
#530160000000
0!
0%
b100 *
0-
02
b100 6
#530170000000
1!
1%
1-
12
#530180000000
0!
0%
b101 *
0-
02
b101 6
#530190000000
1!
1%
1-
12
#530200000000
0!
0%
b110 *
0-
02
b110 6
#530210000000
1!
1%
1-
12
#530220000000
0!
0%
b111 *
0-
02
b111 6
#530230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#530240000000
0!
0%
b0 *
0-
02
b0 6
#530250000000
1!
1%
1-
12
#530260000000
0!
0%
b1 *
0-
02
b1 6
#530270000000
1!
1%
1-
12
#530280000000
0!
0%
b10 *
0-
02
b10 6
#530290000000
1!
1%
1-
12
#530300000000
0!
0%
b11 *
0-
02
b11 6
#530310000000
1!
1%
1-
12
15
#530320000000
0!
0%
b100 *
0-
02
b100 6
#530330000000
1!
1%
1-
12
#530340000000
0!
0%
b101 *
0-
02
b101 6
#530350000000
1!
1%
1-
12
#530360000000
0!
0%
b110 *
0-
02
b110 6
#530370000000
1!
1%
1-
12
#530380000000
0!
0%
b111 *
0-
02
b111 6
#530390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#530400000000
0!
0%
b0 *
0-
02
b0 6
#530410000000
1!
1%
1-
12
#530420000000
0!
0%
b1 *
0-
02
b1 6
#530430000000
1!
1%
1-
12
#530440000000
0!
0%
b10 *
0-
02
b10 6
#530450000000
1!
1%
1-
12
#530460000000
0!
0%
b11 *
0-
02
b11 6
#530470000000
1!
1%
1-
12
15
#530480000000
0!
0%
b100 *
0-
02
b100 6
#530490000000
1!
1%
1-
12
#530500000000
0!
0%
b101 *
0-
02
b101 6
#530510000000
1!
1%
1-
12
#530520000000
0!
0%
b110 *
0-
02
b110 6
#530530000000
1!
1%
1-
12
#530540000000
0!
0%
b111 *
0-
02
b111 6
#530550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#530560000000
0!
0%
b0 *
0-
02
b0 6
#530570000000
1!
1%
1-
12
#530580000000
0!
0%
b1 *
0-
02
b1 6
#530590000000
1!
1%
1-
12
#530600000000
0!
0%
b10 *
0-
02
b10 6
#530610000000
1!
1%
1-
12
#530620000000
0!
0%
b11 *
0-
02
b11 6
#530630000000
1!
1%
1-
12
15
#530640000000
0!
0%
b100 *
0-
02
b100 6
#530650000000
1!
1%
1-
12
#530660000000
0!
0%
b101 *
0-
02
b101 6
#530670000000
1!
1%
1-
12
#530680000000
0!
0%
b110 *
0-
02
b110 6
#530690000000
1!
1%
1-
12
#530700000000
0!
0%
b111 *
0-
02
b111 6
#530710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#530720000000
0!
0%
b0 *
0-
02
b0 6
#530730000000
1!
1%
1-
12
#530740000000
0!
0%
b1 *
0-
02
b1 6
#530750000000
1!
1%
1-
12
#530760000000
0!
0%
b10 *
0-
02
b10 6
#530770000000
1!
1%
1-
12
#530780000000
0!
0%
b11 *
0-
02
b11 6
#530790000000
1!
1%
1-
12
15
#530800000000
0!
0%
b100 *
0-
02
b100 6
#530810000000
1!
1%
1-
12
#530820000000
0!
0%
b101 *
0-
02
b101 6
#530830000000
1!
1%
1-
12
#530840000000
0!
0%
b110 *
0-
02
b110 6
#530850000000
1!
1%
1-
12
#530860000000
0!
0%
b111 *
0-
02
b111 6
#530870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#530880000000
0!
0%
b0 *
0-
02
b0 6
#530890000000
1!
1%
1-
12
#530900000000
0!
0%
b1 *
0-
02
b1 6
#530910000000
1!
1%
1-
12
#530920000000
0!
0%
b10 *
0-
02
b10 6
#530930000000
1!
1%
1-
12
#530940000000
0!
0%
b11 *
0-
02
b11 6
#530950000000
1!
1%
1-
12
15
#530960000000
0!
0%
b100 *
0-
02
b100 6
#530970000000
1!
1%
1-
12
#530980000000
0!
0%
b101 *
0-
02
b101 6
#530990000000
1!
1%
1-
12
#531000000000
0!
0%
b110 *
0-
02
b110 6
#531010000000
1!
1%
1-
12
#531020000000
0!
0%
b111 *
0-
02
b111 6
#531030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#531040000000
0!
0%
b0 *
0-
02
b0 6
#531050000000
1!
1%
1-
12
#531060000000
0!
0%
b1 *
0-
02
b1 6
#531070000000
1!
1%
1-
12
#531080000000
0!
0%
b10 *
0-
02
b10 6
#531090000000
1!
1%
1-
12
#531100000000
0!
0%
b11 *
0-
02
b11 6
#531110000000
1!
1%
1-
12
15
#531120000000
0!
0%
b100 *
0-
02
b100 6
#531130000000
1!
1%
1-
12
#531140000000
0!
0%
b101 *
0-
02
b101 6
#531150000000
1!
1%
1-
12
#531160000000
0!
0%
b110 *
0-
02
b110 6
#531170000000
1!
1%
1-
12
#531180000000
0!
0%
b111 *
0-
02
b111 6
#531190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#531200000000
0!
0%
b0 *
0-
02
b0 6
#531210000000
1!
1%
1-
12
#531220000000
0!
0%
b1 *
0-
02
b1 6
#531230000000
1!
1%
1-
12
#531240000000
0!
0%
b10 *
0-
02
b10 6
#531250000000
1!
1%
1-
12
#531260000000
0!
0%
b11 *
0-
02
b11 6
#531270000000
1!
1%
1-
12
15
#531280000000
0!
0%
b100 *
0-
02
b100 6
#531290000000
1!
1%
1-
12
#531300000000
0!
0%
b101 *
0-
02
b101 6
#531310000000
1!
1%
1-
12
#531320000000
0!
0%
b110 *
0-
02
b110 6
#531330000000
1!
1%
1-
12
#531340000000
0!
0%
b111 *
0-
02
b111 6
#531350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#531360000000
0!
0%
b0 *
0-
02
b0 6
#531370000000
1!
1%
1-
12
#531380000000
0!
0%
b1 *
0-
02
b1 6
#531390000000
1!
1%
1-
12
#531400000000
0!
0%
b10 *
0-
02
b10 6
#531410000000
1!
1%
1-
12
#531420000000
0!
0%
b11 *
0-
02
b11 6
#531430000000
1!
1%
1-
12
15
#531440000000
0!
0%
b100 *
0-
02
b100 6
#531450000000
1!
1%
1-
12
#531460000000
0!
0%
b101 *
0-
02
b101 6
#531470000000
1!
1%
1-
12
#531480000000
0!
0%
b110 *
0-
02
b110 6
#531490000000
1!
1%
1-
12
#531500000000
0!
0%
b111 *
0-
02
b111 6
#531510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#531520000000
0!
0%
b0 *
0-
02
b0 6
#531530000000
1!
1%
1-
12
#531540000000
0!
0%
b1 *
0-
02
b1 6
#531550000000
1!
1%
1-
12
#531560000000
0!
0%
b10 *
0-
02
b10 6
#531570000000
1!
1%
1-
12
#531580000000
0!
0%
b11 *
0-
02
b11 6
#531590000000
1!
1%
1-
12
15
#531600000000
0!
0%
b100 *
0-
02
b100 6
#531610000000
1!
1%
1-
12
#531620000000
0!
0%
b101 *
0-
02
b101 6
#531630000000
1!
1%
1-
12
#531640000000
0!
0%
b110 *
0-
02
b110 6
#531650000000
1!
1%
1-
12
#531660000000
0!
0%
b111 *
0-
02
b111 6
#531670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#531680000000
0!
0%
b0 *
0-
02
b0 6
#531690000000
1!
1%
1-
12
#531700000000
0!
0%
b1 *
0-
02
b1 6
#531710000000
1!
1%
1-
12
#531720000000
0!
0%
b10 *
0-
02
b10 6
#531730000000
1!
1%
1-
12
#531740000000
0!
0%
b11 *
0-
02
b11 6
#531750000000
1!
1%
1-
12
15
#531760000000
0!
0%
b100 *
0-
02
b100 6
#531770000000
1!
1%
1-
12
#531780000000
0!
0%
b101 *
0-
02
b101 6
#531790000000
1!
1%
1-
12
#531800000000
0!
0%
b110 *
0-
02
b110 6
#531810000000
1!
1%
1-
12
#531820000000
0!
0%
b111 *
0-
02
b111 6
#531830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#531840000000
0!
0%
b0 *
0-
02
b0 6
#531850000000
1!
1%
1-
12
#531860000000
0!
0%
b1 *
0-
02
b1 6
#531870000000
1!
1%
1-
12
#531880000000
0!
0%
b10 *
0-
02
b10 6
#531890000000
1!
1%
1-
12
#531900000000
0!
0%
b11 *
0-
02
b11 6
#531910000000
1!
1%
1-
12
15
#531920000000
0!
0%
b100 *
0-
02
b100 6
#531930000000
1!
1%
1-
12
#531940000000
0!
0%
b101 *
0-
02
b101 6
#531950000000
1!
1%
1-
12
#531960000000
0!
0%
b110 *
0-
02
b110 6
#531970000000
1!
1%
1-
12
#531980000000
0!
0%
b111 *
0-
02
b111 6
#531990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#532000000000
0!
0%
b0 *
0-
02
b0 6
#532010000000
1!
1%
1-
12
#532020000000
0!
0%
b1 *
0-
02
b1 6
#532030000000
1!
1%
1-
12
#532040000000
0!
0%
b10 *
0-
02
b10 6
#532050000000
1!
1%
1-
12
#532060000000
0!
0%
b11 *
0-
02
b11 6
#532070000000
1!
1%
1-
12
15
#532080000000
0!
0%
b100 *
0-
02
b100 6
#532090000000
1!
1%
1-
12
#532100000000
0!
0%
b101 *
0-
02
b101 6
#532110000000
1!
1%
1-
12
#532120000000
0!
0%
b110 *
0-
02
b110 6
#532130000000
1!
1%
1-
12
#532140000000
0!
0%
b111 *
0-
02
b111 6
#532150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#532160000000
0!
0%
b0 *
0-
02
b0 6
#532170000000
1!
1%
1-
12
#532180000000
0!
0%
b1 *
0-
02
b1 6
#532190000000
1!
1%
1-
12
#532200000000
0!
0%
b10 *
0-
02
b10 6
#532210000000
1!
1%
1-
12
#532220000000
0!
0%
b11 *
0-
02
b11 6
#532230000000
1!
1%
1-
12
15
#532240000000
0!
0%
b100 *
0-
02
b100 6
#532250000000
1!
1%
1-
12
#532260000000
0!
0%
b101 *
0-
02
b101 6
#532270000000
1!
1%
1-
12
#532280000000
0!
0%
b110 *
0-
02
b110 6
#532290000000
1!
1%
1-
12
#532300000000
0!
0%
b111 *
0-
02
b111 6
#532310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#532320000000
0!
0%
b0 *
0-
02
b0 6
#532330000000
1!
1%
1-
12
#532340000000
0!
0%
b1 *
0-
02
b1 6
#532350000000
1!
1%
1-
12
#532360000000
0!
0%
b10 *
0-
02
b10 6
#532370000000
1!
1%
1-
12
#532380000000
0!
0%
b11 *
0-
02
b11 6
#532390000000
1!
1%
1-
12
15
#532400000000
0!
0%
b100 *
0-
02
b100 6
#532410000000
1!
1%
1-
12
#532420000000
0!
0%
b101 *
0-
02
b101 6
#532430000000
1!
1%
1-
12
#532440000000
0!
0%
b110 *
0-
02
b110 6
#532450000000
1!
1%
1-
12
#532460000000
0!
0%
b111 *
0-
02
b111 6
#532470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#532480000000
0!
0%
b0 *
0-
02
b0 6
#532490000000
1!
1%
1-
12
#532500000000
0!
0%
b1 *
0-
02
b1 6
#532510000000
1!
1%
1-
12
#532520000000
0!
0%
b10 *
0-
02
b10 6
#532530000000
1!
1%
1-
12
#532540000000
0!
0%
b11 *
0-
02
b11 6
#532550000000
1!
1%
1-
12
15
#532560000000
0!
0%
b100 *
0-
02
b100 6
#532570000000
1!
1%
1-
12
#532580000000
0!
0%
b101 *
0-
02
b101 6
#532590000000
1!
1%
1-
12
#532600000000
0!
0%
b110 *
0-
02
b110 6
#532610000000
1!
1%
1-
12
#532620000000
0!
0%
b111 *
0-
02
b111 6
#532630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#532640000000
0!
0%
b0 *
0-
02
b0 6
#532650000000
1!
1%
1-
12
#532660000000
0!
0%
b1 *
0-
02
b1 6
#532670000000
1!
1%
1-
12
#532680000000
0!
0%
b10 *
0-
02
b10 6
#532690000000
1!
1%
1-
12
#532700000000
0!
0%
b11 *
0-
02
b11 6
#532710000000
1!
1%
1-
12
15
#532720000000
0!
0%
b100 *
0-
02
b100 6
#532730000000
1!
1%
1-
12
#532740000000
0!
0%
b101 *
0-
02
b101 6
#532750000000
1!
1%
1-
12
#532760000000
0!
0%
b110 *
0-
02
b110 6
#532770000000
1!
1%
1-
12
#532780000000
0!
0%
b111 *
0-
02
b111 6
#532790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#532800000000
0!
0%
b0 *
0-
02
b0 6
#532810000000
1!
1%
1-
12
#532820000000
0!
0%
b1 *
0-
02
b1 6
#532830000000
1!
1%
1-
12
#532840000000
0!
0%
b10 *
0-
02
b10 6
#532850000000
1!
1%
1-
12
#532860000000
0!
0%
b11 *
0-
02
b11 6
#532870000000
1!
1%
1-
12
15
#532880000000
0!
0%
b100 *
0-
02
b100 6
#532890000000
1!
1%
1-
12
#532900000000
0!
0%
b101 *
0-
02
b101 6
#532910000000
1!
1%
1-
12
#532920000000
0!
0%
b110 *
0-
02
b110 6
#532930000000
1!
1%
1-
12
#532940000000
0!
0%
b111 *
0-
02
b111 6
#532950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#532960000000
0!
0%
b0 *
0-
02
b0 6
#532970000000
1!
1%
1-
12
#532980000000
0!
0%
b1 *
0-
02
b1 6
#532990000000
1!
1%
1-
12
#533000000000
0!
0%
b10 *
0-
02
b10 6
#533010000000
1!
1%
1-
12
#533020000000
0!
0%
b11 *
0-
02
b11 6
#533030000000
1!
1%
1-
12
15
#533040000000
0!
0%
b100 *
0-
02
b100 6
#533050000000
1!
1%
1-
12
#533060000000
0!
0%
b101 *
0-
02
b101 6
#533070000000
1!
1%
1-
12
#533080000000
0!
0%
b110 *
0-
02
b110 6
#533090000000
1!
1%
1-
12
#533100000000
0!
0%
b111 *
0-
02
b111 6
#533110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#533120000000
0!
0%
b0 *
0-
02
b0 6
#533130000000
1!
1%
1-
12
#533140000000
0!
0%
b1 *
0-
02
b1 6
#533150000000
1!
1%
1-
12
#533160000000
0!
0%
b10 *
0-
02
b10 6
#533170000000
1!
1%
1-
12
#533180000000
0!
0%
b11 *
0-
02
b11 6
#533190000000
1!
1%
1-
12
15
#533200000000
0!
0%
b100 *
0-
02
b100 6
#533210000000
1!
1%
1-
12
#533220000000
0!
0%
b101 *
0-
02
b101 6
#533230000000
1!
1%
1-
12
#533240000000
0!
0%
b110 *
0-
02
b110 6
#533250000000
1!
1%
1-
12
#533260000000
0!
0%
b111 *
0-
02
b111 6
#533270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#533280000000
0!
0%
b0 *
0-
02
b0 6
#533290000000
1!
1%
1-
12
#533300000000
0!
0%
b1 *
0-
02
b1 6
#533310000000
1!
1%
1-
12
#533320000000
0!
0%
b10 *
0-
02
b10 6
#533330000000
1!
1%
1-
12
#533340000000
0!
0%
b11 *
0-
02
b11 6
#533350000000
1!
1%
1-
12
15
#533360000000
0!
0%
b100 *
0-
02
b100 6
#533370000000
1!
1%
1-
12
#533380000000
0!
0%
b101 *
0-
02
b101 6
#533390000000
1!
1%
1-
12
#533400000000
0!
0%
b110 *
0-
02
b110 6
#533410000000
1!
1%
1-
12
#533420000000
0!
0%
b111 *
0-
02
b111 6
#533430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#533440000000
0!
0%
b0 *
0-
02
b0 6
#533450000000
1!
1%
1-
12
#533460000000
0!
0%
b1 *
0-
02
b1 6
#533470000000
1!
1%
1-
12
#533480000000
0!
0%
b10 *
0-
02
b10 6
#533490000000
1!
1%
1-
12
#533500000000
0!
0%
b11 *
0-
02
b11 6
#533510000000
1!
1%
1-
12
15
#533520000000
0!
0%
b100 *
0-
02
b100 6
#533530000000
1!
1%
1-
12
#533540000000
0!
0%
b101 *
0-
02
b101 6
#533550000000
1!
1%
1-
12
#533560000000
0!
0%
b110 *
0-
02
b110 6
#533570000000
1!
1%
1-
12
#533580000000
0!
0%
b111 *
0-
02
b111 6
#533590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#533600000000
0!
0%
b0 *
0-
02
b0 6
#533610000000
1!
1%
1-
12
#533620000000
0!
0%
b1 *
0-
02
b1 6
#533630000000
1!
1%
1-
12
#533640000000
0!
0%
b10 *
0-
02
b10 6
#533650000000
1!
1%
1-
12
#533660000000
0!
0%
b11 *
0-
02
b11 6
#533670000000
1!
1%
1-
12
15
#533680000000
0!
0%
b100 *
0-
02
b100 6
#533690000000
1!
1%
1-
12
#533700000000
0!
0%
b101 *
0-
02
b101 6
#533710000000
1!
1%
1-
12
#533720000000
0!
0%
b110 *
0-
02
b110 6
#533730000000
1!
1%
1-
12
#533740000000
0!
0%
b111 *
0-
02
b111 6
#533750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#533760000000
0!
0%
b0 *
0-
02
b0 6
#533770000000
1!
1%
1-
12
#533780000000
0!
0%
b1 *
0-
02
b1 6
#533790000000
1!
1%
1-
12
#533800000000
0!
0%
b10 *
0-
02
b10 6
#533810000000
1!
1%
1-
12
#533820000000
0!
0%
b11 *
0-
02
b11 6
#533830000000
1!
1%
1-
12
15
#533840000000
0!
0%
b100 *
0-
02
b100 6
#533850000000
1!
1%
1-
12
#533860000000
0!
0%
b101 *
0-
02
b101 6
#533870000000
1!
1%
1-
12
#533880000000
0!
0%
b110 *
0-
02
b110 6
#533890000000
1!
1%
1-
12
#533900000000
0!
0%
b111 *
0-
02
b111 6
#533910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#533920000000
0!
0%
b0 *
0-
02
b0 6
#533930000000
1!
1%
1-
12
#533940000000
0!
0%
b1 *
0-
02
b1 6
#533950000000
1!
1%
1-
12
#533960000000
0!
0%
b10 *
0-
02
b10 6
#533970000000
1!
1%
1-
12
#533980000000
0!
0%
b11 *
0-
02
b11 6
#533990000000
1!
1%
1-
12
15
#534000000000
0!
0%
b100 *
0-
02
b100 6
#534010000000
1!
1%
1-
12
#534020000000
0!
0%
b101 *
0-
02
b101 6
#534030000000
1!
1%
1-
12
#534040000000
0!
0%
b110 *
0-
02
b110 6
#534050000000
1!
1%
1-
12
#534060000000
0!
0%
b111 *
0-
02
b111 6
#534070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#534080000000
0!
0%
b0 *
0-
02
b0 6
#534090000000
1!
1%
1-
12
#534100000000
0!
0%
b1 *
0-
02
b1 6
#534110000000
1!
1%
1-
12
#534120000000
0!
0%
b10 *
0-
02
b10 6
#534130000000
1!
1%
1-
12
#534140000000
0!
0%
b11 *
0-
02
b11 6
#534150000000
1!
1%
1-
12
15
#534160000000
0!
0%
b100 *
0-
02
b100 6
#534170000000
1!
1%
1-
12
#534180000000
0!
0%
b101 *
0-
02
b101 6
#534190000000
1!
1%
1-
12
#534200000000
0!
0%
b110 *
0-
02
b110 6
#534210000000
1!
1%
1-
12
#534220000000
0!
0%
b111 *
0-
02
b111 6
#534230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#534240000000
0!
0%
b0 *
0-
02
b0 6
#534250000000
1!
1%
1-
12
#534260000000
0!
0%
b1 *
0-
02
b1 6
#534270000000
1!
1%
1-
12
#534280000000
0!
0%
b10 *
0-
02
b10 6
#534290000000
1!
1%
1-
12
#534300000000
0!
0%
b11 *
0-
02
b11 6
#534310000000
1!
1%
1-
12
15
#534320000000
0!
0%
b100 *
0-
02
b100 6
#534330000000
1!
1%
1-
12
#534340000000
0!
0%
b101 *
0-
02
b101 6
#534350000000
1!
1%
1-
12
#534360000000
0!
0%
b110 *
0-
02
b110 6
#534370000000
1!
1%
1-
12
#534380000000
0!
0%
b111 *
0-
02
b111 6
#534390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#534400000000
0!
0%
b0 *
0-
02
b0 6
#534410000000
1!
1%
1-
12
#534420000000
0!
0%
b1 *
0-
02
b1 6
#534430000000
1!
1%
1-
12
#534440000000
0!
0%
b10 *
0-
02
b10 6
#534450000000
1!
1%
1-
12
#534460000000
0!
0%
b11 *
0-
02
b11 6
#534470000000
1!
1%
1-
12
15
#534480000000
0!
0%
b100 *
0-
02
b100 6
#534490000000
1!
1%
1-
12
#534500000000
0!
0%
b101 *
0-
02
b101 6
#534510000000
1!
1%
1-
12
#534520000000
0!
0%
b110 *
0-
02
b110 6
#534530000000
1!
1%
1-
12
#534540000000
0!
0%
b111 *
0-
02
b111 6
#534550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#534560000000
0!
0%
b0 *
0-
02
b0 6
#534570000000
1!
1%
1-
12
#534580000000
0!
0%
b1 *
0-
02
b1 6
#534590000000
1!
1%
1-
12
#534600000000
0!
0%
b10 *
0-
02
b10 6
#534610000000
1!
1%
1-
12
#534620000000
0!
0%
b11 *
0-
02
b11 6
#534630000000
1!
1%
1-
12
15
#534640000000
0!
0%
b100 *
0-
02
b100 6
#534650000000
1!
1%
1-
12
#534660000000
0!
0%
b101 *
0-
02
b101 6
#534670000000
1!
1%
1-
12
#534680000000
0!
0%
b110 *
0-
02
b110 6
#534690000000
1!
1%
1-
12
#534700000000
0!
0%
b111 *
0-
02
b111 6
#534710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#534720000000
0!
0%
b0 *
0-
02
b0 6
#534730000000
1!
1%
1-
12
#534740000000
0!
0%
b1 *
0-
02
b1 6
#534750000000
1!
1%
1-
12
#534760000000
0!
0%
b10 *
0-
02
b10 6
#534770000000
1!
1%
1-
12
#534780000000
0!
0%
b11 *
0-
02
b11 6
#534790000000
1!
1%
1-
12
15
#534800000000
0!
0%
b100 *
0-
02
b100 6
#534810000000
1!
1%
1-
12
#534820000000
0!
0%
b101 *
0-
02
b101 6
#534830000000
1!
1%
1-
12
#534840000000
0!
0%
b110 *
0-
02
b110 6
#534850000000
1!
1%
1-
12
#534860000000
0!
0%
b111 *
0-
02
b111 6
#534870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#534880000000
0!
0%
b0 *
0-
02
b0 6
#534890000000
1!
1%
1-
12
#534900000000
0!
0%
b1 *
0-
02
b1 6
#534910000000
1!
1%
1-
12
#534920000000
0!
0%
b10 *
0-
02
b10 6
#534930000000
1!
1%
1-
12
#534940000000
0!
0%
b11 *
0-
02
b11 6
#534950000000
1!
1%
1-
12
15
#534960000000
0!
0%
b100 *
0-
02
b100 6
#534970000000
1!
1%
1-
12
#534980000000
0!
0%
b101 *
0-
02
b101 6
#534990000000
1!
1%
1-
12
#535000000000
0!
0%
b110 *
0-
02
b110 6
#535010000000
1!
1%
1-
12
#535020000000
0!
0%
b111 *
0-
02
b111 6
#535030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#535040000000
0!
0%
b0 *
0-
02
b0 6
#535050000000
1!
1%
1-
12
#535060000000
0!
0%
b1 *
0-
02
b1 6
#535070000000
1!
1%
1-
12
#535080000000
0!
0%
b10 *
0-
02
b10 6
#535090000000
1!
1%
1-
12
#535100000000
0!
0%
b11 *
0-
02
b11 6
#535110000000
1!
1%
1-
12
15
#535120000000
0!
0%
b100 *
0-
02
b100 6
#535130000000
1!
1%
1-
12
#535140000000
0!
0%
b101 *
0-
02
b101 6
#535150000000
1!
1%
1-
12
#535160000000
0!
0%
b110 *
0-
02
b110 6
#535170000000
1!
1%
1-
12
#535180000000
0!
0%
b111 *
0-
02
b111 6
#535190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#535200000000
0!
0%
b0 *
0-
02
b0 6
#535210000000
1!
1%
1-
12
#535220000000
0!
0%
b1 *
0-
02
b1 6
#535230000000
1!
1%
1-
12
#535240000000
0!
0%
b10 *
0-
02
b10 6
#535250000000
1!
1%
1-
12
#535260000000
0!
0%
b11 *
0-
02
b11 6
#535270000000
1!
1%
1-
12
15
#535280000000
0!
0%
b100 *
0-
02
b100 6
#535290000000
1!
1%
1-
12
#535300000000
0!
0%
b101 *
0-
02
b101 6
#535310000000
1!
1%
1-
12
#535320000000
0!
0%
b110 *
0-
02
b110 6
#535330000000
1!
1%
1-
12
#535340000000
0!
0%
b111 *
0-
02
b111 6
#535350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#535360000000
0!
0%
b0 *
0-
02
b0 6
#535370000000
1!
1%
1-
12
#535380000000
0!
0%
b1 *
0-
02
b1 6
#535390000000
1!
1%
1-
12
#535400000000
0!
0%
b10 *
0-
02
b10 6
#535410000000
1!
1%
1-
12
#535420000000
0!
0%
b11 *
0-
02
b11 6
#535430000000
1!
1%
1-
12
15
#535440000000
0!
0%
b100 *
0-
02
b100 6
#535450000000
1!
1%
1-
12
#535460000000
0!
0%
b101 *
0-
02
b101 6
#535470000000
1!
1%
1-
12
#535480000000
0!
0%
b110 *
0-
02
b110 6
#535490000000
1!
1%
1-
12
#535500000000
0!
0%
b111 *
0-
02
b111 6
#535510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#535520000000
0!
0%
b0 *
0-
02
b0 6
#535530000000
1!
1%
1-
12
#535540000000
0!
0%
b1 *
0-
02
b1 6
#535550000000
1!
1%
1-
12
#535560000000
0!
0%
b10 *
0-
02
b10 6
#535570000000
1!
1%
1-
12
#535580000000
0!
0%
b11 *
0-
02
b11 6
#535590000000
1!
1%
1-
12
15
#535600000000
0!
0%
b100 *
0-
02
b100 6
#535610000000
1!
1%
1-
12
#535620000000
0!
0%
b101 *
0-
02
b101 6
#535630000000
1!
1%
1-
12
#535640000000
0!
0%
b110 *
0-
02
b110 6
#535650000000
1!
1%
1-
12
#535660000000
0!
0%
b111 *
0-
02
b111 6
#535670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#535680000000
0!
0%
b0 *
0-
02
b0 6
#535690000000
1!
1%
1-
12
#535700000000
0!
0%
b1 *
0-
02
b1 6
#535710000000
1!
1%
1-
12
#535720000000
0!
0%
b10 *
0-
02
b10 6
#535730000000
1!
1%
1-
12
#535740000000
0!
0%
b11 *
0-
02
b11 6
#535750000000
1!
1%
1-
12
15
#535760000000
0!
0%
b100 *
0-
02
b100 6
#535770000000
1!
1%
1-
12
#535780000000
0!
0%
b101 *
0-
02
b101 6
#535790000000
1!
1%
1-
12
#535800000000
0!
0%
b110 *
0-
02
b110 6
#535810000000
1!
1%
1-
12
#535820000000
0!
0%
b111 *
0-
02
b111 6
#535830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#535840000000
0!
0%
b0 *
0-
02
b0 6
#535850000000
1!
1%
1-
12
#535860000000
0!
0%
b1 *
0-
02
b1 6
#535870000000
1!
1%
1-
12
#535880000000
0!
0%
b10 *
0-
02
b10 6
#535890000000
1!
1%
1-
12
#535900000000
0!
0%
b11 *
0-
02
b11 6
#535910000000
1!
1%
1-
12
15
#535920000000
0!
0%
b100 *
0-
02
b100 6
#535930000000
1!
1%
1-
12
#535940000000
0!
0%
b101 *
0-
02
b101 6
#535950000000
1!
1%
1-
12
#535960000000
0!
0%
b110 *
0-
02
b110 6
#535970000000
1!
1%
1-
12
#535980000000
0!
0%
b111 *
0-
02
b111 6
#535990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#536000000000
0!
0%
b0 *
0-
02
b0 6
#536010000000
1!
1%
1-
12
#536020000000
0!
0%
b1 *
0-
02
b1 6
#536030000000
1!
1%
1-
12
#536040000000
0!
0%
b10 *
0-
02
b10 6
#536050000000
1!
1%
1-
12
#536060000000
0!
0%
b11 *
0-
02
b11 6
#536070000000
1!
1%
1-
12
15
#536080000000
0!
0%
b100 *
0-
02
b100 6
#536090000000
1!
1%
1-
12
#536100000000
0!
0%
b101 *
0-
02
b101 6
#536110000000
1!
1%
1-
12
#536120000000
0!
0%
b110 *
0-
02
b110 6
#536130000000
1!
1%
1-
12
#536140000000
0!
0%
b111 *
0-
02
b111 6
#536150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#536160000000
0!
0%
b0 *
0-
02
b0 6
#536170000000
1!
1%
1-
12
#536180000000
0!
0%
b1 *
0-
02
b1 6
#536190000000
1!
1%
1-
12
#536200000000
0!
0%
b10 *
0-
02
b10 6
#536210000000
1!
1%
1-
12
#536220000000
0!
0%
b11 *
0-
02
b11 6
#536230000000
1!
1%
1-
12
15
#536240000000
0!
0%
b100 *
0-
02
b100 6
#536250000000
1!
1%
1-
12
#536260000000
0!
0%
b101 *
0-
02
b101 6
#536270000000
1!
1%
1-
12
#536280000000
0!
0%
b110 *
0-
02
b110 6
#536290000000
1!
1%
1-
12
#536300000000
0!
0%
b111 *
0-
02
b111 6
#536310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#536320000000
0!
0%
b0 *
0-
02
b0 6
#536330000000
1!
1%
1-
12
#536340000000
0!
0%
b1 *
0-
02
b1 6
#536350000000
1!
1%
1-
12
#536360000000
0!
0%
b10 *
0-
02
b10 6
#536370000000
1!
1%
1-
12
#536380000000
0!
0%
b11 *
0-
02
b11 6
#536390000000
1!
1%
1-
12
15
#536400000000
0!
0%
b100 *
0-
02
b100 6
#536410000000
1!
1%
1-
12
#536420000000
0!
0%
b101 *
0-
02
b101 6
#536430000000
1!
1%
1-
12
#536440000000
0!
0%
b110 *
0-
02
b110 6
#536450000000
1!
1%
1-
12
#536460000000
0!
0%
b111 *
0-
02
b111 6
#536470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#536480000000
0!
0%
b0 *
0-
02
b0 6
#536490000000
1!
1%
1-
12
#536500000000
0!
0%
b1 *
0-
02
b1 6
#536510000000
1!
1%
1-
12
#536520000000
0!
0%
b10 *
0-
02
b10 6
#536530000000
1!
1%
1-
12
#536540000000
0!
0%
b11 *
0-
02
b11 6
#536550000000
1!
1%
1-
12
15
#536560000000
0!
0%
b100 *
0-
02
b100 6
#536570000000
1!
1%
1-
12
#536580000000
0!
0%
b101 *
0-
02
b101 6
#536590000000
1!
1%
1-
12
#536600000000
0!
0%
b110 *
0-
02
b110 6
#536610000000
1!
1%
1-
12
#536620000000
0!
0%
b111 *
0-
02
b111 6
#536630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#536640000000
0!
0%
b0 *
0-
02
b0 6
#536650000000
1!
1%
1-
12
#536660000000
0!
0%
b1 *
0-
02
b1 6
#536670000000
1!
1%
1-
12
#536680000000
0!
0%
b10 *
0-
02
b10 6
#536690000000
1!
1%
1-
12
#536700000000
0!
0%
b11 *
0-
02
b11 6
#536710000000
1!
1%
1-
12
15
#536720000000
0!
0%
b100 *
0-
02
b100 6
#536730000000
1!
1%
1-
12
#536740000000
0!
0%
b101 *
0-
02
b101 6
#536750000000
1!
1%
1-
12
#536760000000
0!
0%
b110 *
0-
02
b110 6
#536770000000
1!
1%
1-
12
#536780000000
0!
0%
b111 *
0-
02
b111 6
#536790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#536800000000
0!
0%
b0 *
0-
02
b0 6
#536810000000
1!
1%
1-
12
#536820000000
0!
0%
b1 *
0-
02
b1 6
#536830000000
1!
1%
1-
12
#536840000000
0!
0%
b10 *
0-
02
b10 6
#536850000000
1!
1%
1-
12
#536860000000
0!
0%
b11 *
0-
02
b11 6
#536870000000
1!
1%
1-
12
15
#536880000000
0!
0%
b100 *
0-
02
b100 6
#536890000000
1!
1%
1-
12
#536900000000
0!
0%
b101 *
0-
02
b101 6
#536910000000
1!
1%
1-
12
#536920000000
0!
0%
b110 *
0-
02
b110 6
#536930000000
1!
1%
1-
12
#536940000000
0!
0%
b111 *
0-
02
b111 6
#536950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#536960000000
0!
0%
b0 *
0-
02
b0 6
#536970000000
1!
1%
1-
12
#536980000000
0!
0%
b1 *
0-
02
b1 6
#536990000000
1!
1%
1-
12
#537000000000
0!
0%
b10 *
0-
02
b10 6
#537010000000
1!
1%
1-
12
#537020000000
0!
0%
b11 *
0-
02
b11 6
#537030000000
1!
1%
1-
12
15
#537040000000
0!
0%
b100 *
0-
02
b100 6
#537050000000
1!
1%
1-
12
#537060000000
0!
0%
b101 *
0-
02
b101 6
#537070000000
1!
1%
1-
12
#537080000000
0!
0%
b110 *
0-
02
b110 6
#537090000000
1!
1%
1-
12
#537100000000
0!
0%
b111 *
0-
02
b111 6
#537110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#537120000000
0!
0%
b0 *
0-
02
b0 6
#537130000000
1!
1%
1-
12
#537140000000
0!
0%
b1 *
0-
02
b1 6
#537150000000
1!
1%
1-
12
#537160000000
0!
0%
b10 *
0-
02
b10 6
#537170000000
1!
1%
1-
12
#537180000000
0!
0%
b11 *
0-
02
b11 6
#537190000000
1!
1%
1-
12
15
#537200000000
0!
0%
b100 *
0-
02
b100 6
#537210000000
1!
1%
1-
12
#537220000000
0!
0%
b101 *
0-
02
b101 6
#537230000000
1!
1%
1-
12
#537240000000
0!
0%
b110 *
0-
02
b110 6
#537250000000
1!
1%
1-
12
#537260000000
0!
0%
b111 *
0-
02
b111 6
#537270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#537280000000
0!
0%
b0 *
0-
02
b0 6
#537290000000
1!
1%
1-
12
#537300000000
0!
0%
b1 *
0-
02
b1 6
#537310000000
1!
1%
1-
12
#537320000000
0!
0%
b10 *
0-
02
b10 6
#537330000000
1!
1%
1-
12
#537340000000
0!
0%
b11 *
0-
02
b11 6
#537350000000
1!
1%
1-
12
15
#537360000000
0!
0%
b100 *
0-
02
b100 6
#537370000000
1!
1%
1-
12
#537380000000
0!
0%
b101 *
0-
02
b101 6
#537390000000
1!
1%
1-
12
#537400000000
0!
0%
b110 *
0-
02
b110 6
#537410000000
1!
1%
1-
12
#537420000000
0!
0%
b111 *
0-
02
b111 6
#537430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#537440000000
0!
0%
b0 *
0-
02
b0 6
#537450000000
1!
1%
1-
12
#537460000000
0!
0%
b1 *
0-
02
b1 6
#537470000000
1!
1%
1-
12
#537480000000
0!
0%
b10 *
0-
02
b10 6
#537490000000
1!
1%
1-
12
#537500000000
0!
0%
b11 *
0-
02
b11 6
#537510000000
1!
1%
1-
12
15
#537520000000
0!
0%
b100 *
0-
02
b100 6
#537530000000
1!
1%
1-
12
#537540000000
0!
0%
b101 *
0-
02
b101 6
#537550000000
1!
1%
1-
12
#537560000000
0!
0%
b110 *
0-
02
b110 6
#537570000000
1!
1%
1-
12
#537580000000
0!
0%
b111 *
0-
02
b111 6
#537590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#537600000000
0!
0%
b0 *
0-
02
b0 6
#537610000000
1!
1%
1-
12
#537620000000
0!
0%
b1 *
0-
02
b1 6
#537630000000
1!
1%
1-
12
#537640000000
0!
0%
b10 *
0-
02
b10 6
#537650000000
1!
1%
1-
12
#537660000000
0!
0%
b11 *
0-
02
b11 6
#537670000000
1!
1%
1-
12
15
#537680000000
0!
0%
b100 *
0-
02
b100 6
#537690000000
1!
1%
1-
12
#537700000000
0!
0%
b101 *
0-
02
b101 6
#537710000000
1!
1%
1-
12
#537720000000
0!
0%
b110 *
0-
02
b110 6
#537730000000
1!
1%
1-
12
#537740000000
0!
0%
b111 *
0-
02
b111 6
#537750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#537760000000
0!
0%
b0 *
0-
02
b0 6
#537770000000
1!
1%
1-
12
#537780000000
0!
0%
b1 *
0-
02
b1 6
#537790000000
1!
1%
1-
12
#537800000000
0!
0%
b10 *
0-
02
b10 6
#537810000000
1!
1%
1-
12
#537820000000
0!
0%
b11 *
0-
02
b11 6
#537830000000
1!
1%
1-
12
15
#537840000000
0!
0%
b100 *
0-
02
b100 6
#537850000000
1!
1%
1-
12
#537860000000
0!
0%
b101 *
0-
02
b101 6
#537870000000
1!
1%
1-
12
#537880000000
0!
0%
b110 *
0-
02
b110 6
#537890000000
1!
1%
1-
12
#537900000000
0!
0%
b111 *
0-
02
b111 6
#537910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#537920000000
0!
0%
b0 *
0-
02
b0 6
#537930000000
1!
1%
1-
12
#537940000000
0!
0%
b1 *
0-
02
b1 6
#537950000000
1!
1%
1-
12
#537960000000
0!
0%
b10 *
0-
02
b10 6
#537970000000
1!
1%
1-
12
#537980000000
0!
0%
b11 *
0-
02
b11 6
#537990000000
1!
1%
1-
12
15
#538000000000
0!
0%
b100 *
0-
02
b100 6
#538010000000
1!
1%
1-
12
#538020000000
0!
0%
b101 *
0-
02
b101 6
#538030000000
1!
1%
1-
12
#538040000000
0!
0%
b110 *
0-
02
b110 6
#538050000000
1!
1%
1-
12
#538060000000
0!
0%
b111 *
0-
02
b111 6
#538070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#538080000000
0!
0%
b0 *
0-
02
b0 6
#538090000000
1!
1%
1-
12
#538100000000
0!
0%
b1 *
0-
02
b1 6
#538110000000
1!
1%
1-
12
#538120000000
0!
0%
b10 *
0-
02
b10 6
#538130000000
1!
1%
1-
12
#538140000000
0!
0%
b11 *
0-
02
b11 6
#538150000000
1!
1%
1-
12
15
#538160000000
0!
0%
b100 *
0-
02
b100 6
#538170000000
1!
1%
1-
12
#538180000000
0!
0%
b101 *
0-
02
b101 6
#538190000000
1!
1%
1-
12
#538200000000
0!
0%
b110 *
0-
02
b110 6
#538210000000
1!
1%
1-
12
#538220000000
0!
0%
b111 *
0-
02
b111 6
#538230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#538240000000
0!
0%
b0 *
0-
02
b0 6
#538250000000
1!
1%
1-
12
#538260000000
0!
0%
b1 *
0-
02
b1 6
#538270000000
1!
1%
1-
12
#538280000000
0!
0%
b10 *
0-
02
b10 6
#538290000000
1!
1%
1-
12
#538300000000
0!
0%
b11 *
0-
02
b11 6
#538310000000
1!
1%
1-
12
15
#538320000000
0!
0%
b100 *
0-
02
b100 6
#538330000000
1!
1%
1-
12
#538340000000
0!
0%
b101 *
0-
02
b101 6
#538350000000
1!
1%
1-
12
#538360000000
0!
0%
b110 *
0-
02
b110 6
#538370000000
1!
1%
1-
12
#538380000000
0!
0%
b111 *
0-
02
b111 6
#538390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#538400000000
0!
0%
b0 *
0-
02
b0 6
#538410000000
1!
1%
1-
12
#538420000000
0!
0%
b1 *
0-
02
b1 6
#538430000000
1!
1%
1-
12
#538440000000
0!
0%
b10 *
0-
02
b10 6
#538450000000
1!
1%
1-
12
#538460000000
0!
0%
b11 *
0-
02
b11 6
#538470000000
1!
1%
1-
12
15
#538480000000
0!
0%
b100 *
0-
02
b100 6
#538490000000
1!
1%
1-
12
#538500000000
0!
0%
b101 *
0-
02
b101 6
#538510000000
1!
1%
1-
12
#538520000000
0!
0%
b110 *
0-
02
b110 6
#538530000000
1!
1%
1-
12
#538540000000
0!
0%
b111 *
0-
02
b111 6
#538550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#538560000000
0!
0%
b0 *
0-
02
b0 6
#538570000000
1!
1%
1-
12
#538580000000
0!
0%
b1 *
0-
02
b1 6
#538590000000
1!
1%
1-
12
#538600000000
0!
0%
b10 *
0-
02
b10 6
#538610000000
1!
1%
1-
12
#538620000000
0!
0%
b11 *
0-
02
b11 6
#538630000000
1!
1%
1-
12
15
#538640000000
0!
0%
b100 *
0-
02
b100 6
#538650000000
1!
1%
1-
12
#538660000000
0!
0%
b101 *
0-
02
b101 6
#538670000000
1!
1%
1-
12
#538680000000
0!
0%
b110 *
0-
02
b110 6
#538690000000
1!
1%
1-
12
#538700000000
0!
0%
b111 *
0-
02
b111 6
#538710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#538720000000
0!
0%
b0 *
0-
02
b0 6
#538730000000
1!
1%
1-
12
#538740000000
0!
0%
b1 *
0-
02
b1 6
#538750000000
1!
1%
1-
12
#538760000000
0!
0%
b10 *
0-
02
b10 6
#538770000000
1!
1%
1-
12
#538780000000
0!
0%
b11 *
0-
02
b11 6
#538790000000
1!
1%
1-
12
15
#538800000000
0!
0%
b100 *
0-
02
b100 6
#538810000000
1!
1%
1-
12
#538820000000
0!
0%
b101 *
0-
02
b101 6
#538830000000
1!
1%
1-
12
#538840000000
0!
0%
b110 *
0-
02
b110 6
#538850000000
1!
1%
1-
12
#538860000000
0!
0%
b111 *
0-
02
b111 6
#538870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#538880000000
0!
0%
b0 *
0-
02
b0 6
#538890000000
1!
1%
1-
12
#538900000000
0!
0%
b1 *
0-
02
b1 6
#538910000000
1!
1%
1-
12
#538920000000
0!
0%
b10 *
0-
02
b10 6
#538930000000
1!
1%
1-
12
#538940000000
0!
0%
b11 *
0-
02
b11 6
#538950000000
1!
1%
1-
12
15
#538960000000
0!
0%
b100 *
0-
02
b100 6
#538970000000
1!
1%
1-
12
#538980000000
0!
0%
b101 *
0-
02
b101 6
#538990000000
1!
1%
1-
12
#539000000000
0!
0%
b110 *
0-
02
b110 6
#539010000000
1!
1%
1-
12
#539020000000
0!
0%
b111 *
0-
02
b111 6
#539030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#539040000000
0!
0%
b0 *
0-
02
b0 6
#539050000000
1!
1%
1-
12
#539060000000
0!
0%
b1 *
0-
02
b1 6
#539070000000
1!
1%
1-
12
#539080000000
0!
0%
b10 *
0-
02
b10 6
#539090000000
1!
1%
1-
12
#539100000000
0!
0%
b11 *
0-
02
b11 6
#539110000000
1!
1%
1-
12
15
#539120000000
0!
0%
b100 *
0-
02
b100 6
#539130000000
1!
1%
1-
12
#539140000000
0!
0%
b101 *
0-
02
b101 6
#539150000000
1!
1%
1-
12
#539160000000
0!
0%
b110 *
0-
02
b110 6
#539170000000
1!
1%
1-
12
#539180000000
0!
0%
b111 *
0-
02
b111 6
#539190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#539200000000
0!
0%
b0 *
0-
02
b0 6
#539210000000
1!
1%
1-
12
#539220000000
0!
0%
b1 *
0-
02
b1 6
#539230000000
1!
1%
1-
12
#539240000000
0!
0%
b10 *
0-
02
b10 6
#539250000000
1!
1%
1-
12
#539260000000
0!
0%
b11 *
0-
02
b11 6
#539270000000
1!
1%
1-
12
15
#539280000000
0!
0%
b100 *
0-
02
b100 6
#539290000000
1!
1%
1-
12
#539300000000
0!
0%
b101 *
0-
02
b101 6
#539310000000
1!
1%
1-
12
#539320000000
0!
0%
b110 *
0-
02
b110 6
#539330000000
1!
1%
1-
12
#539340000000
0!
0%
b111 *
0-
02
b111 6
#539350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#539360000000
0!
0%
b0 *
0-
02
b0 6
#539370000000
1!
1%
1-
12
#539380000000
0!
0%
b1 *
0-
02
b1 6
#539390000000
1!
1%
1-
12
#539400000000
0!
0%
b10 *
0-
02
b10 6
#539410000000
1!
1%
1-
12
#539420000000
0!
0%
b11 *
0-
02
b11 6
#539430000000
1!
1%
1-
12
15
#539440000000
0!
0%
b100 *
0-
02
b100 6
#539450000000
1!
1%
1-
12
#539460000000
0!
0%
b101 *
0-
02
b101 6
#539470000000
1!
1%
1-
12
#539480000000
0!
0%
b110 *
0-
02
b110 6
#539490000000
1!
1%
1-
12
#539500000000
0!
0%
b111 *
0-
02
b111 6
#539510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#539520000000
0!
0%
b0 *
0-
02
b0 6
#539530000000
1!
1%
1-
12
#539540000000
0!
0%
b1 *
0-
02
b1 6
#539550000000
1!
1%
1-
12
#539560000000
0!
0%
b10 *
0-
02
b10 6
#539570000000
1!
1%
1-
12
#539580000000
0!
0%
b11 *
0-
02
b11 6
#539590000000
1!
1%
1-
12
15
#539600000000
0!
0%
b100 *
0-
02
b100 6
#539610000000
1!
1%
1-
12
#539620000000
0!
0%
b101 *
0-
02
b101 6
#539630000000
1!
1%
1-
12
#539640000000
0!
0%
b110 *
0-
02
b110 6
#539650000000
1!
1%
1-
12
#539660000000
0!
0%
b111 *
0-
02
b111 6
#539670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#539680000000
0!
0%
b0 *
0-
02
b0 6
#539690000000
1!
1%
1-
12
#539700000000
0!
0%
b1 *
0-
02
b1 6
#539710000000
1!
1%
1-
12
#539720000000
0!
0%
b10 *
0-
02
b10 6
#539730000000
1!
1%
1-
12
#539740000000
0!
0%
b11 *
0-
02
b11 6
#539750000000
1!
1%
1-
12
15
#539760000000
0!
0%
b100 *
0-
02
b100 6
#539770000000
1!
1%
1-
12
#539780000000
0!
0%
b101 *
0-
02
b101 6
#539790000000
1!
1%
1-
12
#539800000000
0!
0%
b110 *
0-
02
b110 6
#539810000000
1!
1%
1-
12
#539820000000
0!
0%
b111 *
0-
02
b111 6
#539830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#539840000000
0!
0%
b0 *
0-
02
b0 6
#539850000000
1!
1%
1-
12
#539860000000
0!
0%
b1 *
0-
02
b1 6
#539870000000
1!
1%
1-
12
#539880000000
0!
0%
b10 *
0-
02
b10 6
#539890000000
1!
1%
1-
12
#539900000000
0!
0%
b11 *
0-
02
b11 6
#539910000000
1!
1%
1-
12
15
#539920000000
0!
0%
b100 *
0-
02
b100 6
#539930000000
1!
1%
1-
12
#539940000000
0!
0%
b101 *
0-
02
b101 6
#539950000000
1!
1%
1-
12
#539960000000
0!
0%
b110 *
0-
02
b110 6
#539970000000
1!
1%
1-
12
#539980000000
0!
0%
b111 *
0-
02
b111 6
#539990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#540000000000
0!
0%
b0 *
0-
02
b0 6
#540010000000
1!
1%
1-
12
#540020000000
0!
0%
b1 *
0-
02
b1 6
#540030000000
1!
1%
1-
12
#540040000000
0!
0%
b10 *
0-
02
b10 6
#540050000000
1!
1%
1-
12
#540060000000
0!
0%
b11 *
0-
02
b11 6
#540070000000
1!
1%
1-
12
15
#540080000000
0!
0%
b100 *
0-
02
b100 6
#540090000000
1!
1%
1-
12
#540100000000
0!
0%
b101 *
0-
02
b101 6
#540110000000
1!
1%
1-
12
#540120000000
0!
0%
b110 *
0-
02
b110 6
#540130000000
1!
1%
1-
12
#540140000000
0!
0%
b111 *
0-
02
b111 6
#540150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#540160000000
0!
0%
b0 *
0-
02
b0 6
#540170000000
1!
1%
1-
12
#540180000000
0!
0%
b1 *
0-
02
b1 6
#540190000000
1!
1%
1-
12
#540200000000
0!
0%
b10 *
0-
02
b10 6
#540210000000
1!
1%
1-
12
#540220000000
0!
0%
b11 *
0-
02
b11 6
#540230000000
1!
1%
1-
12
15
#540240000000
0!
0%
b100 *
0-
02
b100 6
#540250000000
1!
1%
1-
12
#540260000000
0!
0%
b101 *
0-
02
b101 6
#540270000000
1!
1%
1-
12
#540280000000
0!
0%
b110 *
0-
02
b110 6
#540290000000
1!
1%
1-
12
#540300000000
0!
0%
b111 *
0-
02
b111 6
#540310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#540320000000
0!
0%
b0 *
0-
02
b0 6
#540330000000
1!
1%
1-
12
#540340000000
0!
0%
b1 *
0-
02
b1 6
#540350000000
1!
1%
1-
12
#540360000000
0!
0%
b10 *
0-
02
b10 6
#540370000000
1!
1%
1-
12
#540380000000
0!
0%
b11 *
0-
02
b11 6
#540390000000
1!
1%
1-
12
15
#540400000000
0!
0%
b100 *
0-
02
b100 6
#540410000000
1!
1%
1-
12
#540420000000
0!
0%
b101 *
0-
02
b101 6
#540430000000
1!
1%
1-
12
#540440000000
0!
0%
b110 *
0-
02
b110 6
#540450000000
1!
1%
1-
12
#540460000000
0!
0%
b111 *
0-
02
b111 6
#540470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#540480000000
0!
0%
b0 *
0-
02
b0 6
#540490000000
1!
1%
1-
12
#540500000000
0!
0%
b1 *
0-
02
b1 6
#540510000000
1!
1%
1-
12
#540520000000
0!
0%
b10 *
0-
02
b10 6
#540530000000
1!
1%
1-
12
#540540000000
0!
0%
b11 *
0-
02
b11 6
#540550000000
1!
1%
1-
12
15
#540560000000
0!
0%
b100 *
0-
02
b100 6
#540570000000
1!
1%
1-
12
#540580000000
0!
0%
b101 *
0-
02
b101 6
#540590000000
1!
1%
1-
12
#540600000000
0!
0%
b110 *
0-
02
b110 6
#540610000000
1!
1%
1-
12
#540620000000
0!
0%
b111 *
0-
02
b111 6
#540630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#540640000000
0!
0%
b0 *
0-
02
b0 6
#540650000000
1!
1%
1-
12
#540660000000
0!
0%
b1 *
0-
02
b1 6
#540670000000
1!
1%
1-
12
#540680000000
0!
0%
b10 *
0-
02
b10 6
#540690000000
1!
1%
1-
12
#540700000000
0!
0%
b11 *
0-
02
b11 6
#540710000000
1!
1%
1-
12
15
#540720000000
0!
0%
b100 *
0-
02
b100 6
#540730000000
1!
1%
1-
12
#540740000000
0!
0%
b101 *
0-
02
b101 6
#540750000000
1!
1%
1-
12
#540760000000
0!
0%
b110 *
0-
02
b110 6
#540770000000
1!
1%
1-
12
#540780000000
0!
0%
b111 *
0-
02
b111 6
#540790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#540800000000
0!
0%
b0 *
0-
02
b0 6
#540810000000
1!
1%
1-
12
#540820000000
0!
0%
b1 *
0-
02
b1 6
#540830000000
1!
1%
1-
12
#540840000000
0!
0%
b10 *
0-
02
b10 6
#540850000000
1!
1%
1-
12
#540860000000
0!
0%
b11 *
0-
02
b11 6
#540870000000
1!
1%
1-
12
15
#540880000000
0!
0%
b100 *
0-
02
b100 6
#540890000000
1!
1%
1-
12
#540900000000
0!
0%
b101 *
0-
02
b101 6
#540910000000
1!
1%
1-
12
#540920000000
0!
0%
b110 *
0-
02
b110 6
#540930000000
1!
1%
1-
12
#540940000000
0!
0%
b111 *
0-
02
b111 6
#540950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#540960000000
0!
0%
b0 *
0-
02
b0 6
#540970000000
1!
1%
1-
12
#540980000000
0!
0%
b1 *
0-
02
b1 6
#540990000000
1!
1%
1-
12
#541000000000
0!
0%
b10 *
0-
02
b10 6
#541010000000
1!
1%
1-
12
#541020000000
0!
0%
b11 *
0-
02
b11 6
#541030000000
1!
1%
1-
12
15
#541040000000
0!
0%
b100 *
0-
02
b100 6
#541050000000
1!
1%
1-
12
#541060000000
0!
0%
b101 *
0-
02
b101 6
#541070000000
1!
1%
1-
12
#541080000000
0!
0%
b110 *
0-
02
b110 6
#541090000000
1!
1%
1-
12
#541100000000
0!
0%
b111 *
0-
02
b111 6
#541110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#541120000000
0!
0%
b0 *
0-
02
b0 6
#541130000000
1!
1%
1-
12
#541140000000
0!
0%
b1 *
0-
02
b1 6
#541150000000
1!
1%
1-
12
#541160000000
0!
0%
b10 *
0-
02
b10 6
#541170000000
1!
1%
1-
12
#541180000000
0!
0%
b11 *
0-
02
b11 6
#541190000000
1!
1%
1-
12
15
#541200000000
0!
0%
b100 *
0-
02
b100 6
#541210000000
1!
1%
1-
12
#541220000000
0!
0%
b101 *
0-
02
b101 6
#541230000000
1!
1%
1-
12
#541240000000
0!
0%
b110 *
0-
02
b110 6
#541250000000
1!
1%
1-
12
#541260000000
0!
0%
b111 *
0-
02
b111 6
#541270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#541280000000
0!
0%
b0 *
0-
02
b0 6
#541290000000
1!
1%
1-
12
#541300000000
0!
0%
b1 *
0-
02
b1 6
#541310000000
1!
1%
1-
12
#541320000000
0!
0%
b10 *
0-
02
b10 6
#541330000000
1!
1%
1-
12
#541340000000
0!
0%
b11 *
0-
02
b11 6
#541350000000
1!
1%
1-
12
15
#541360000000
0!
0%
b100 *
0-
02
b100 6
#541370000000
1!
1%
1-
12
#541380000000
0!
0%
b101 *
0-
02
b101 6
#541390000000
1!
1%
1-
12
#541400000000
0!
0%
b110 *
0-
02
b110 6
#541410000000
1!
1%
1-
12
#541420000000
0!
0%
b111 *
0-
02
b111 6
#541430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#541440000000
0!
0%
b0 *
0-
02
b0 6
#541450000000
1!
1%
1-
12
#541460000000
0!
0%
b1 *
0-
02
b1 6
#541470000000
1!
1%
1-
12
#541480000000
0!
0%
b10 *
0-
02
b10 6
#541490000000
1!
1%
1-
12
#541500000000
0!
0%
b11 *
0-
02
b11 6
#541510000000
1!
1%
1-
12
15
#541520000000
0!
0%
b100 *
0-
02
b100 6
#541530000000
1!
1%
1-
12
#541540000000
0!
0%
b101 *
0-
02
b101 6
#541550000000
1!
1%
1-
12
#541560000000
0!
0%
b110 *
0-
02
b110 6
#541570000000
1!
1%
1-
12
#541580000000
0!
0%
b111 *
0-
02
b111 6
#541590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#541600000000
0!
0%
b0 *
0-
02
b0 6
#541610000000
1!
1%
1-
12
#541620000000
0!
0%
b1 *
0-
02
b1 6
#541630000000
1!
1%
1-
12
#541640000000
0!
0%
b10 *
0-
02
b10 6
#541650000000
1!
1%
1-
12
#541660000000
0!
0%
b11 *
0-
02
b11 6
#541670000000
1!
1%
1-
12
15
#541680000000
0!
0%
b100 *
0-
02
b100 6
#541690000000
1!
1%
1-
12
#541700000000
0!
0%
b101 *
0-
02
b101 6
#541710000000
1!
1%
1-
12
#541720000000
0!
0%
b110 *
0-
02
b110 6
#541730000000
1!
1%
1-
12
#541740000000
0!
0%
b111 *
0-
02
b111 6
#541750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#541760000000
0!
0%
b0 *
0-
02
b0 6
#541770000000
1!
1%
1-
12
#541780000000
0!
0%
b1 *
0-
02
b1 6
#541790000000
1!
1%
1-
12
#541800000000
0!
0%
b10 *
0-
02
b10 6
#541810000000
1!
1%
1-
12
#541820000000
0!
0%
b11 *
0-
02
b11 6
#541830000000
1!
1%
1-
12
15
#541840000000
0!
0%
b100 *
0-
02
b100 6
#541850000000
1!
1%
1-
12
#541860000000
0!
0%
b101 *
0-
02
b101 6
#541870000000
1!
1%
1-
12
#541880000000
0!
0%
b110 *
0-
02
b110 6
#541890000000
1!
1%
1-
12
#541900000000
0!
0%
b111 *
0-
02
b111 6
#541910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#541920000000
0!
0%
b0 *
0-
02
b0 6
#541930000000
1!
1%
1-
12
#541940000000
0!
0%
b1 *
0-
02
b1 6
#541950000000
1!
1%
1-
12
#541960000000
0!
0%
b10 *
0-
02
b10 6
#541970000000
1!
1%
1-
12
#541980000000
0!
0%
b11 *
0-
02
b11 6
#541990000000
1!
1%
1-
12
15
#542000000000
0!
0%
b100 *
0-
02
b100 6
#542010000000
1!
1%
1-
12
#542020000000
0!
0%
b101 *
0-
02
b101 6
#542030000000
1!
1%
1-
12
#542040000000
0!
0%
b110 *
0-
02
b110 6
#542050000000
1!
1%
1-
12
#542060000000
0!
0%
b111 *
0-
02
b111 6
#542070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#542080000000
0!
0%
b0 *
0-
02
b0 6
#542090000000
1!
1%
1-
12
#542100000000
0!
0%
b1 *
0-
02
b1 6
#542110000000
1!
1%
1-
12
#542120000000
0!
0%
b10 *
0-
02
b10 6
#542130000000
1!
1%
1-
12
#542140000000
0!
0%
b11 *
0-
02
b11 6
#542150000000
1!
1%
1-
12
15
#542160000000
0!
0%
b100 *
0-
02
b100 6
#542170000000
1!
1%
1-
12
#542180000000
0!
0%
b101 *
0-
02
b101 6
#542190000000
1!
1%
1-
12
#542200000000
0!
0%
b110 *
0-
02
b110 6
#542210000000
1!
1%
1-
12
#542220000000
0!
0%
b111 *
0-
02
b111 6
#542230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#542240000000
0!
0%
b0 *
0-
02
b0 6
#542250000000
1!
1%
1-
12
#542260000000
0!
0%
b1 *
0-
02
b1 6
#542270000000
1!
1%
1-
12
#542280000000
0!
0%
b10 *
0-
02
b10 6
#542290000000
1!
1%
1-
12
#542300000000
0!
0%
b11 *
0-
02
b11 6
#542310000000
1!
1%
1-
12
15
#542320000000
0!
0%
b100 *
0-
02
b100 6
#542330000000
1!
1%
1-
12
#542340000000
0!
0%
b101 *
0-
02
b101 6
#542350000000
1!
1%
1-
12
#542360000000
0!
0%
b110 *
0-
02
b110 6
#542370000000
1!
1%
1-
12
#542380000000
0!
0%
b111 *
0-
02
b111 6
#542390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#542400000000
0!
0%
b0 *
0-
02
b0 6
#542410000000
1!
1%
1-
12
#542420000000
0!
0%
b1 *
0-
02
b1 6
#542430000000
1!
1%
1-
12
#542440000000
0!
0%
b10 *
0-
02
b10 6
#542450000000
1!
1%
1-
12
#542460000000
0!
0%
b11 *
0-
02
b11 6
#542470000000
1!
1%
1-
12
15
#542480000000
0!
0%
b100 *
0-
02
b100 6
#542490000000
1!
1%
1-
12
#542500000000
0!
0%
b101 *
0-
02
b101 6
#542510000000
1!
1%
1-
12
#542520000000
0!
0%
b110 *
0-
02
b110 6
#542530000000
1!
1%
1-
12
#542540000000
0!
0%
b111 *
0-
02
b111 6
#542550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#542560000000
0!
0%
b0 *
0-
02
b0 6
#542570000000
1!
1%
1-
12
#542580000000
0!
0%
b1 *
0-
02
b1 6
#542590000000
1!
1%
1-
12
#542600000000
0!
0%
b10 *
0-
02
b10 6
#542610000000
1!
1%
1-
12
#542620000000
0!
0%
b11 *
0-
02
b11 6
#542630000000
1!
1%
1-
12
15
#542640000000
0!
0%
b100 *
0-
02
b100 6
#542650000000
1!
1%
1-
12
#542660000000
0!
0%
b101 *
0-
02
b101 6
#542670000000
1!
1%
1-
12
#542680000000
0!
0%
b110 *
0-
02
b110 6
#542690000000
1!
1%
1-
12
#542700000000
0!
0%
b111 *
0-
02
b111 6
#542710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#542720000000
0!
0%
b0 *
0-
02
b0 6
#542730000000
1!
1%
1-
12
#542740000000
0!
0%
b1 *
0-
02
b1 6
#542750000000
1!
1%
1-
12
#542760000000
0!
0%
b10 *
0-
02
b10 6
#542770000000
1!
1%
1-
12
#542780000000
0!
0%
b11 *
0-
02
b11 6
#542790000000
1!
1%
1-
12
15
#542800000000
0!
0%
b100 *
0-
02
b100 6
#542810000000
1!
1%
1-
12
#542820000000
0!
0%
b101 *
0-
02
b101 6
#542830000000
1!
1%
1-
12
#542840000000
0!
0%
b110 *
0-
02
b110 6
#542850000000
1!
1%
1-
12
#542860000000
0!
0%
b111 *
0-
02
b111 6
#542870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#542880000000
0!
0%
b0 *
0-
02
b0 6
#542890000000
1!
1%
1-
12
#542900000000
0!
0%
b1 *
0-
02
b1 6
#542910000000
1!
1%
1-
12
#542920000000
0!
0%
b10 *
0-
02
b10 6
#542930000000
1!
1%
1-
12
#542940000000
0!
0%
b11 *
0-
02
b11 6
#542950000000
1!
1%
1-
12
15
#542960000000
0!
0%
b100 *
0-
02
b100 6
#542970000000
1!
1%
1-
12
#542980000000
0!
0%
b101 *
0-
02
b101 6
#542990000000
1!
1%
1-
12
#543000000000
0!
0%
b110 *
0-
02
b110 6
#543010000000
1!
1%
1-
12
#543020000000
0!
0%
b111 *
0-
02
b111 6
#543030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#543040000000
0!
0%
b0 *
0-
02
b0 6
#543050000000
1!
1%
1-
12
#543060000000
0!
0%
b1 *
0-
02
b1 6
#543070000000
1!
1%
1-
12
#543080000000
0!
0%
b10 *
0-
02
b10 6
#543090000000
1!
1%
1-
12
#543100000000
0!
0%
b11 *
0-
02
b11 6
#543110000000
1!
1%
1-
12
15
#543120000000
0!
0%
b100 *
0-
02
b100 6
#543130000000
1!
1%
1-
12
#543140000000
0!
0%
b101 *
0-
02
b101 6
#543150000000
1!
1%
1-
12
#543160000000
0!
0%
b110 *
0-
02
b110 6
#543170000000
1!
1%
1-
12
#543180000000
0!
0%
b111 *
0-
02
b111 6
#543190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#543200000000
0!
0%
b0 *
0-
02
b0 6
#543210000000
1!
1%
1-
12
#543220000000
0!
0%
b1 *
0-
02
b1 6
#543230000000
1!
1%
1-
12
#543240000000
0!
0%
b10 *
0-
02
b10 6
#543250000000
1!
1%
1-
12
#543260000000
0!
0%
b11 *
0-
02
b11 6
#543270000000
1!
1%
1-
12
15
#543280000000
0!
0%
b100 *
0-
02
b100 6
#543290000000
1!
1%
1-
12
#543300000000
0!
0%
b101 *
0-
02
b101 6
#543310000000
1!
1%
1-
12
#543320000000
0!
0%
b110 *
0-
02
b110 6
#543330000000
1!
1%
1-
12
#543340000000
0!
0%
b111 *
0-
02
b111 6
#543350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#543360000000
0!
0%
b0 *
0-
02
b0 6
#543370000000
1!
1%
1-
12
#543380000000
0!
0%
b1 *
0-
02
b1 6
#543390000000
1!
1%
1-
12
#543400000000
0!
0%
b10 *
0-
02
b10 6
#543410000000
1!
1%
1-
12
#543420000000
0!
0%
b11 *
0-
02
b11 6
#543430000000
1!
1%
1-
12
15
#543440000000
0!
0%
b100 *
0-
02
b100 6
#543450000000
1!
1%
1-
12
#543460000000
0!
0%
b101 *
0-
02
b101 6
#543470000000
1!
1%
1-
12
#543480000000
0!
0%
b110 *
0-
02
b110 6
#543490000000
1!
1%
1-
12
#543500000000
0!
0%
b111 *
0-
02
b111 6
#543510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#543520000000
0!
0%
b0 *
0-
02
b0 6
#543530000000
1!
1%
1-
12
#543540000000
0!
0%
b1 *
0-
02
b1 6
#543550000000
1!
1%
1-
12
#543560000000
0!
0%
b10 *
0-
02
b10 6
#543570000000
1!
1%
1-
12
#543580000000
0!
0%
b11 *
0-
02
b11 6
#543590000000
1!
1%
1-
12
15
#543600000000
0!
0%
b100 *
0-
02
b100 6
#543610000000
1!
1%
1-
12
#543620000000
0!
0%
b101 *
0-
02
b101 6
#543630000000
1!
1%
1-
12
#543640000000
0!
0%
b110 *
0-
02
b110 6
#543650000000
1!
1%
1-
12
#543660000000
0!
0%
b111 *
0-
02
b111 6
#543670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#543680000000
0!
0%
b0 *
0-
02
b0 6
#543690000000
1!
1%
1-
12
#543700000000
0!
0%
b1 *
0-
02
b1 6
#543710000000
1!
1%
1-
12
#543720000000
0!
0%
b10 *
0-
02
b10 6
#543730000000
1!
1%
1-
12
#543740000000
0!
0%
b11 *
0-
02
b11 6
#543750000000
1!
1%
1-
12
15
#543760000000
0!
0%
b100 *
0-
02
b100 6
#543770000000
1!
1%
1-
12
#543780000000
0!
0%
b101 *
0-
02
b101 6
#543790000000
1!
1%
1-
12
#543800000000
0!
0%
b110 *
0-
02
b110 6
#543810000000
1!
1%
1-
12
#543820000000
0!
0%
b111 *
0-
02
b111 6
#543830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#543840000000
0!
0%
b0 *
0-
02
b0 6
#543850000000
1!
1%
1-
12
#543860000000
0!
0%
b1 *
0-
02
b1 6
#543870000000
1!
1%
1-
12
#543880000000
0!
0%
b10 *
0-
02
b10 6
#543890000000
1!
1%
1-
12
#543900000000
0!
0%
b11 *
0-
02
b11 6
#543910000000
1!
1%
1-
12
15
#543920000000
0!
0%
b100 *
0-
02
b100 6
#543930000000
1!
1%
1-
12
#543940000000
0!
0%
b101 *
0-
02
b101 6
#543950000000
1!
1%
1-
12
#543960000000
0!
0%
b110 *
0-
02
b110 6
#543970000000
1!
1%
1-
12
#543980000000
0!
0%
b111 *
0-
02
b111 6
#543990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#544000000000
0!
0%
b0 *
0-
02
b0 6
#544010000000
1!
1%
1-
12
#544020000000
0!
0%
b1 *
0-
02
b1 6
#544030000000
1!
1%
1-
12
#544040000000
0!
0%
b10 *
0-
02
b10 6
#544050000000
1!
1%
1-
12
#544060000000
0!
0%
b11 *
0-
02
b11 6
#544070000000
1!
1%
1-
12
15
#544080000000
0!
0%
b100 *
0-
02
b100 6
#544090000000
1!
1%
1-
12
#544100000000
0!
0%
b101 *
0-
02
b101 6
#544110000000
1!
1%
1-
12
#544120000000
0!
0%
b110 *
0-
02
b110 6
#544130000000
1!
1%
1-
12
#544140000000
0!
0%
b111 *
0-
02
b111 6
#544150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#544160000000
0!
0%
b0 *
0-
02
b0 6
#544170000000
1!
1%
1-
12
#544180000000
0!
0%
b1 *
0-
02
b1 6
#544190000000
1!
1%
1-
12
#544200000000
0!
0%
b10 *
0-
02
b10 6
#544210000000
1!
1%
1-
12
#544220000000
0!
0%
b11 *
0-
02
b11 6
#544230000000
1!
1%
1-
12
15
#544240000000
0!
0%
b100 *
0-
02
b100 6
#544250000000
1!
1%
1-
12
#544260000000
0!
0%
b101 *
0-
02
b101 6
#544270000000
1!
1%
1-
12
#544280000000
0!
0%
b110 *
0-
02
b110 6
#544290000000
1!
1%
1-
12
#544300000000
0!
0%
b111 *
0-
02
b111 6
#544310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#544320000000
0!
0%
b0 *
0-
02
b0 6
#544330000000
1!
1%
1-
12
#544340000000
0!
0%
b1 *
0-
02
b1 6
#544350000000
1!
1%
1-
12
#544360000000
0!
0%
b10 *
0-
02
b10 6
#544370000000
1!
1%
1-
12
#544380000000
0!
0%
b11 *
0-
02
b11 6
#544390000000
1!
1%
1-
12
15
#544400000000
0!
0%
b100 *
0-
02
b100 6
#544410000000
1!
1%
1-
12
#544420000000
0!
0%
b101 *
0-
02
b101 6
#544430000000
1!
1%
1-
12
#544440000000
0!
0%
b110 *
0-
02
b110 6
#544450000000
1!
1%
1-
12
#544460000000
0!
0%
b111 *
0-
02
b111 6
#544470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#544480000000
0!
0%
b0 *
0-
02
b0 6
#544490000000
1!
1%
1-
12
#544500000000
0!
0%
b1 *
0-
02
b1 6
#544510000000
1!
1%
1-
12
#544520000000
0!
0%
b10 *
0-
02
b10 6
#544530000000
1!
1%
1-
12
#544540000000
0!
0%
b11 *
0-
02
b11 6
#544550000000
1!
1%
1-
12
15
#544560000000
0!
0%
b100 *
0-
02
b100 6
#544570000000
1!
1%
1-
12
#544580000000
0!
0%
b101 *
0-
02
b101 6
#544590000000
1!
1%
1-
12
#544600000000
0!
0%
b110 *
0-
02
b110 6
#544610000000
1!
1%
1-
12
#544620000000
0!
0%
b111 *
0-
02
b111 6
#544630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#544640000000
0!
0%
b0 *
0-
02
b0 6
#544650000000
1!
1%
1-
12
#544660000000
0!
0%
b1 *
0-
02
b1 6
#544670000000
1!
1%
1-
12
#544680000000
0!
0%
b10 *
0-
02
b10 6
#544690000000
1!
1%
1-
12
#544700000000
0!
0%
b11 *
0-
02
b11 6
#544710000000
1!
1%
1-
12
15
#544720000000
0!
0%
b100 *
0-
02
b100 6
#544730000000
1!
1%
1-
12
#544740000000
0!
0%
b101 *
0-
02
b101 6
#544750000000
1!
1%
1-
12
#544760000000
0!
0%
b110 *
0-
02
b110 6
#544770000000
1!
1%
1-
12
#544780000000
0!
0%
b111 *
0-
02
b111 6
#544790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#544800000000
0!
0%
b0 *
0-
02
b0 6
#544810000000
1!
1%
1-
12
#544820000000
0!
0%
b1 *
0-
02
b1 6
#544830000000
1!
1%
1-
12
#544840000000
0!
0%
b10 *
0-
02
b10 6
#544850000000
1!
1%
1-
12
#544860000000
0!
0%
b11 *
0-
02
b11 6
#544870000000
1!
1%
1-
12
15
#544880000000
0!
0%
b100 *
0-
02
b100 6
#544890000000
1!
1%
1-
12
#544900000000
0!
0%
b101 *
0-
02
b101 6
#544910000000
1!
1%
1-
12
#544920000000
0!
0%
b110 *
0-
02
b110 6
#544930000000
1!
1%
1-
12
#544940000000
0!
0%
b111 *
0-
02
b111 6
#544950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#544960000000
0!
0%
b0 *
0-
02
b0 6
#544970000000
1!
1%
1-
12
#544980000000
0!
0%
b1 *
0-
02
b1 6
#544990000000
1!
1%
1-
12
#545000000000
0!
0%
b10 *
0-
02
b10 6
#545010000000
1!
1%
1-
12
#545020000000
0!
0%
b11 *
0-
02
b11 6
#545030000000
1!
1%
1-
12
15
#545040000000
0!
0%
b100 *
0-
02
b100 6
#545050000000
1!
1%
1-
12
#545060000000
0!
0%
b101 *
0-
02
b101 6
#545070000000
1!
1%
1-
12
#545080000000
0!
0%
b110 *
0-
02
b110 6
#545090000000
1!
1%
1-
12
#545100000000
0!
0%
b111 *
0-
02
b111 6
#545110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#545120000000
0!
0%
b0 *
0-
02
b0 6
#545130000000
1!
1%
1-
12
#545140000000
0!
0%
b1 *
0-
02
b1 6
#545150000000
1!
1%
1-
12
#545160000000
0!
0%
b10 *
0-
02
b10 6
#545170000000
1!
1%
1-
12
#545180000000
0!
0%
b11 *
0-
02
b11 6
#545190000000
1!
1%
1-
12
15
#545200000000
0!
0%
b100 *
0-
02
b100 6
#545210000000
1!
1%
1-
12
#545220000000
0!
0%
b101 *
0-
02
b101 6
#545230000000
1!
1%
1-
12
#545240000000
0!
0%
b110 *
0-
02
b110 6
#545250000000
1!
1%
1-
12
#545260000000
0!
0%
b111 *
0-
02
b111 6
#545270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#545280000000
0!
0%
b0 *
0-
02
b0 6
#545290000000
1!
1%
1-
12
#545300000000
0!
0%
b1 *
0-
02
b1 6
#545310000000
1!
1%
1-
12
#545320000000
0!
0%
b10 *
0-
02
b10 6
#545330000000
1!
1%
1-
12
#545340000000
0!
0%
b11 *
0-
02
b11 6
#545350000000
1!
1%
1-
12
15
#545360000000
0!
0%
b100 *
0-
02
b100 6
#545370000000
1!
1%
1-
12
#545380000000
0!
0%
b101 *
0-
02
b101 6
#545390000000
1!
1%
1-
12
#545400000000
0!
0%
b110 *
0-
02
b110 6
#545410000000
1!
1%
1-
12
#545420000000
0!
0%
b111 *
0-
02
b111 6
#545430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#545440000000
0!
0%
b0 *
0-
02
b0 6
#545450000000
1!
1%
1-
12
#545460000000
0!
0%
b1 *
0-
02
b1 6
#545470000000
1!
1%
1-
12
#545480000000
0!
0%
b10 *
0-
02
b10 6
#545490000000
1!
1%
1-
12
#545500000000
0!
0%
b11 *
0-
02
b11 6
#545510000000
1!
1%
1-
12
15
#545520000000
0!
0%
b100 *
0-
02
b100 6
#545530000000
1!
1%
1-
12
#545540000000
0!
0%
b101 *
0-
02
b101 6
#545550000000
1!
1%
1-
12
#545560000000
0!
0%
b110 *
0-
02
b110 6
#545570000000
1!
1%
1-
12
#545580000000
0!
0%
b111 *
0-
02
b111 6
#545590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#545600000000
0!
0%
b0 *
0-
02
b0 6
#545610000000
1!
1%
1-
12
#545620000000
0!
0%
b1 *
0-
02
b1 6
#545630000000
1!
1%
1-
12
#545640000000
0!
0%
b10 *
0-
02
b10 6
#545650000000
1!
1%
1-
12
#545660000000
0!
0%
b11 *
0-
02
b11 6
#545670000000
1!
1%
1-
12
15
#545680000000
0!
0%
b100 *
0-
02
b100 6
#545690000000
1!
1%
1-
12
#545700000000
0!
0%
b101 *
0-
02
b101 6
#545710000000
1!
1%
1-
12
#545720000000
0!
0%
b110 *
0-
02
b110 6
#545730000000
1!
1%
1-
12
#545740000000
0!
0%
b111 *
0-
02
b111 6
#545750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#545760000000
0!
0%
b0 *
0-
02
b0 6
#545770000000
1!
1%
1-
12
#545780000000
0!
0%
b1 *
0-
02
b1 6
#545790000000
1!
1%
1-
12
#545800000000
0!
0%
b10 *
0-
02
b10 6
#545810000000
1!
1%
1-
12
#545820000000
0!
0%
b11 *
0-
02
b11 6
#545830000000
1!
1%
1-
12
15
#545840000000
0!
0%
b100 *
0-
02
b100 6
#545850000000
1!
1%
1-
12
#545860000000
0!
0%
b101 *
0-
02
b101 6
#545870000000
1!
1%
1-
12
#545880000000
0!
0%
b110 *
0-
02
b110 6
#545890000000
1!
1%
1-
12
#545900000000
0!
0%
b111 *
0-
02
b111 6
#545910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#545920000000
0!
0%
b0 *
0-
02
b0 6
#545930000000
1!
1%
1-
12
#545940000000
0!
0%
b1 *
0-
02
b1 6
#545950000000
1!
1%
1-
12
#545960000000
0!
0%
b10 *
0-
02
b10 6
#545970000000
1!
1%
1-
12
#545980000000
0!
0%
b11 *
0-
02
b11 6
#545990000000
1!
1%
1-
12
15
#546000000000
0!
0%
b100 *
0-
02
b100 6
#546010000000
1!
1%
1-
12
#546020000000
0!
0%
b101 *
0-
02
b101 6
#546030000000
1!
1%
1-
12
#546040000000
0!
0%
b110 *
0-
02
b110 6
#546050000000
1!
1%
1-
12
#546060000000
0!
0%
b111 *
0-
02
b111 6
#546070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#546080000000
0!
0%
b0 *
0-
02
b0 6
#546090000000
1!
1%
1-
12
#546100000000
0!
0%
b1 *
0-
02
b1 6
#546110000000
1!
1%
1-
12
#546120000000
0!
0%
b10 *
0-
02
b10 6
#546130000000
1!
1%
1-
12
#546140000000
0!
0%
b11 *
0-
02
b11 6
#546150000000
1!
1%
1-
12
15
#546160000000
0!
0%
b100 *
0-
02
b100 6
#546170000000
1!
1%
1-
12
#546180000000
0!
0%
b101 *
0-
02
b101 6
#546190000000
1!
1%
1-
12
#546200000000
0!
0%
b110 *
0-
02
b110 6
#546210000000
1!
1%
1-
12
#546220000000
0!
0%
b111 *
0-
02
b111 6
#546230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#546240000000
0!
0%
b0 *
0-
02
b0 6
#546250000000
1!
1%
1-
12
#546260000000
0!
0%
b1 *
0-
02
b1 6
#546270000000
1!
1%
1-
12
#546280000000
0!
0%
b10 *
0-
02
b10 6
#546290000000
1!
1%
1-
12
#546300000000
0!
0%
b11 *
0-
02
b11 6
#546310000000
1!
1%
1-
12
15
#546320000000
0!
0%
b100 *
0-
02
b100 6
#546330000000
1!
1%
1-
12
#546340000000
0!
0%
b101 *
0-
02
b101 6
#546350000000
1!
1%
1-
12
#546360000000
0!
0%
b110 *
0-
02
b110 6
#546370000000
1!
1%
1-
12
#546380000000
0!
0%
b111 *
0-
02
b111 6
#546390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#546400000000
0!
0%
b0 *
0-
02
b0 6
#546410000000
1!
1%
1-
12
#546420000000
0!
0%
b1 *
0-
02
b1 6
#546430000000
1!
1%
1-
12
#546440000000
0!
0%
b10 *
0-
02
b10 6
#546450000000
1!
1%
1-
12
#546460000000
0!
0%
b11 *
0-
02
b11 6
#546470000000
1!
1%
1-
12
15
#546480000000
0!
0%
b100 *
0-
02
b100 6
#546490000000
1!
1%
1-
12
#546500000000
0!
0%
b101 *
0-
02
b101 6
#546510000000
1!
1%
1-
12
#546520000000
0!
0%
b110 *
0-
02
b110 6
#546530000000
1!
1%
1-
12
#546540000000
0!
0%
b111 *
0-
02
b111 6
#546550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#546560000000
0!
0%
b0 *
0-
02
b0 6
#546570000000
1!
1%
1-
12
#546580000000
0!
0%
b1 *
0-
02
b1 6
#546590000000
1!
1%
1-
12
#546600000000
0!
0%
b10 *
0-
02
b10 6
#546610000000
1!
1%
1-
12
#546620000000
0!
0%
b11 *
0-
02
b11 6
#546630000000
1!
1%
1-
12
15
#546640000000
0!
0%
b100 *
0-
02
b100 6
#546650000000
1!
1%
1-
12
#546660000000
0!
0%
b101 *
0-
02
b101 6
#546670000000
1!
1%
1-
12
#546680000000
0!
0%
b110 *
0-
02
b110 6
#546690000000
1!
1%
1-
12
#546700000000
0!
0%
b111 *
0-
02
b111 6
#546710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#546720000000
0!
0%
b0 *
0-
02
b0 6
#546730000000
1!
1%
1-
12
#546740000000
0!
0%
b1 *
0-
02
b1 6
#546750000000
1!
1%
1-
12
#546760000000
0!
0%
b10 *
0-
02
b10 6
#546770000000
1!
1%
1-
12
#546780000000
0!
0%
b11 *
0-
02
b11 6
#546790000000
1!
1%
1-
12
15
#546800000000
0!
0%
b100 *
0-
02
b100 6
#546810000000
1!
1%
1-
12
#546820000000
0!
0%
b101 *
0-
02
b101 6
#546830000000
1!
1%
1-
12
#546840000000
0!
0%
b110 *
0-
02
b110 6
#546850000000
1!
1%
1-
12
#546860000000
0!
0%
b111 *
0-
02
b111 6
#546870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#546880000000
0!
0%
b0 *
0-
02
b0 6
#546890000000
1!
1%
1-
12
#546900000000
0!
0%
b1 *
0-
02
b1 6
#546910000000
1!
1%
1-
12
#546920000000
0!
0%
b10 *
0-
02
b10 6
#546930000000
1!
1%
1-
12
#546940000000
0!
0%
b11 *
0-
02
b11 6
#546950000000
1!
1%
1-
12
15
#546960000000
0!
0%
b100 *
0-
02
b100 6
#546970000000
1!
1%
1-
12
#546980000000
0!
0%
b101 *
0-
02
b101 6
#546990000000
1!
1%
1-
12
#547000000000
0!
0%
b110 *
0-
02
b110 6
#547010000000
1!
1%
1-
12
#547020000000
0!
0%
b111 *
0-
02
b111 6
#547030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#547040000000
0!
0%
b0 *
0-
02
b0 6
#547050000000
1!
1%
1-
12
#547060000000
0!
0%
b1 *
0-
02
b1 6
#547070000000
1!
1%
1-
12
#547080000000
0!
0%
b10 *
0-
02
b10 6
#547090000000
1!
1%
1-
12
#547100000000
0!
0%
b11 *
0-
02
b11 6
#547110000000
1!
1%
1-
12
15
#547120000000
0!
0%
b100 *
0-
02
b100 6
#547130000000
1!
1%
1-
12
#547140000000
0!
0%
b101 *
0-
02
b101 6
#547150000000
1!
1%
1-
12
#547160000000
0!
0%
b110 *
0-
02
b110 6
#547170000000
1!
1%
1-
12
#547180000000
0!
0%
b111 *
0-
02
b111 6
#547190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#547200000000
0!
0%
b0 *
0-
02
b0 6
#547210000000
1!
1%
1-
12
#547220000000
0!
0%
b1 *
0-
02
b1 6
#547230000000
1!
1%
1-
12
#547240000000
0!
0%
b10 *
0-
02
b10 6
#547250000000
1!
1%
1-
12
#547260000000
0!
0%
b11 *
0-
02
b11 6
#547270000000
1!
1%
1-
12
15
#547280000000
0!
0%
b100 *
0-
02
b100 6
#547290000000
1!
1%
1-
12
#547300000000
0!
0%
b101 *
0-
02
b101 6
#547310000000
1!
1%
1-
12
#547320000000
0!
0%
b110 *
0-
02
b110 6
#547330000000
1!
1%
1-
12
#547340000000
0!
0%
b111 *
0-
02
b111 6
#547350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#547360000000
0!
0%
b0 *
0-
02
b0 6
#547370000000
1!
1%
1-
12
#547380000000
0!
0%
b1 *
0-
02
b1 6
#547390000000
1!
1%
1-
12
#547400000000
0!
0%
b10 *
0-
02
b10 6
#547410000000
1!
1%
1-
12
#547420000000
0!
0%
b11 *
0-
02
b11 6
#547430000000
1!
1%
1-
12
15
#547440000000
0!
0%
b100 *
0-
02
b100 6
#547450000000
1!
1%
1-
12
#547460000000
0!
0%
b101 *
0-
02
b101 6
#547470000000
1!
1%
1-
12
#547480000000
0!
0%
b110 *
0-
02
b110 6
#547490000000
1!
1%
1-
12
#547500000000
0!
0%
b111 *
0-
02
b111 6
#547510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#547520000000
0!
0%
b0 *
0-
02
b0 6
#547530000000
1!
1%
1-
12
#547540000000
0!
0%
b1 *
0-
02
b1 6
#547550000000
1!
1%
1-
12
#547560000000
0!
0%
b10 *
0-
02
b10 6
#547570000000
1!
1%
1-
12
#547580000000
0!
0%
b11 *
0-
02
b11 6
#547590000000
1!
1%
1-
12
15
#547600000000
0!
0%
b100 *
0-
02
b100 6
#547610000000
1!
1%
1-
12
#547620000000
0!
0%
b101 *
0-
02
b101 6
#547630000000
1!
1%
1-
12
#547640000000
0!
0%
b110 *
0-
02
b110 6
#547650000000
1!
1%
1-
12
#547660000000
0!
0%
b111 *
0-
02
b111 6
#547670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#547680000000
0!
0%
b0 *
0-
02
b0 6
#547690000000
1!
1%
1-
12
#547700000000
0!
0%
b1 *
0-
02
b1 6
#547710000000
1!
1%
1-
12
#547720000000
0!
0%
b10 *
0-
02
b10 6
#547730000000
1!
1%
1-
12
#547740000000
0!
0%
b11 *
0-
02
b11 6
#547750000000
1!
1%
1-
12
15
#547760000000
0!
0%
b100 *
0-
02
b100 6
#547770000000
1!
1%
1-
12
#547780000000
0!
0%
b101 *
0-
02
b101 6
#547790000000
1!
1%
1-
12
#547800000000
0!
0%
b110 *
0-
02
b110 6
#547810000000
1!
1%
1-
12
#547820000000
0!
0%
b111 *
0-
02
b111 6
#547830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#547840000000
0!
0%
b0 *
0-
02
b0 6
#547850000000
1!
1%
1-
12
#547860000000
0!
0%
b1 *
0-
02
b1 6
#547870000000
1!
1%
1-
12
#547880000000
0!
0%
b10 *
0-
02
b10 6
#547890000000
1!
1%
1-
12
#547900000000
0!
0%
b11 *
0-
02
b11 6
#547910000000
1!
1%
1-
12
15
#547920000000
0!
0%
b100 *
0-
02
b100 6
#547930000000
1!
1%
1-
12
#547940000000
0!
0%
b101 *
0-
02
b101 6
#547950000000
1!
1%
1-
12
#547960000000
0!
0%
b110 *
0-
02
b110 6
#547970000000
1!
1%
1-
12
#547980000000
0!
0%
b111 *
0-
02
b111 6
#547990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#548000000000
0!
0%
b0 *
0-
02
b0 6
#548010000000
1!
1%
1-
12
#548020000000
0!
0%
b1 *
0-
02
b1 6
#548030000000
1!
1%
1-
12
#548040000000
0!
0%
b10 *
0-
02
b10 6
#548050000000
1!
1%
1-
12
#548060000000
0!
0%
b11 *
0-
02
b11 6
#548070000000
1!
1%
1-
12
15
#548080000000
0!
0%
b100 *
0-
02
b100 6
#548090000000
1!
1%
1-
12
#548100000000
0!
0%
b101 *
0-
02
b101 6
#548110000000
1!
1%
1-
12
#548120000000
0!
0%
b110 *
0-
02
b110 6
#548130000000
1!
1%
1-
12
#548140000000
0!
0%
b111 *
0-
02
b111 6
#548150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#548160000000
0!
0%
b0 *
0-
02
b0 6
#548170000000
1!
1%
1-
12
#548180000000
0!
0%
b1 *
0-
02
b1 6
#548190000000
1!
1%
1-
12
#548200000000
0!
0%
b10 *
0-
02
b10 6
#548210000000
1!
1%
1-
12
#548220000000
0!
0%
b11 *
0-
02
b11 6
#548230000000
1!
1%
1-
12
15
#548240000000
0!
0%
b100 *
0-
02
b100 6
#548250000000
1!
1%
1-
12
#548260000000
0!
0%
b101 *
0-
02
b101 6
#548270000000
1!
1%
1-
12
#548280000000
0!
0%
b110 *
0-
02
b110 6
#548290000000
1!
1%
1-
12
#548300000000
0!
0%
b111 *
0-
02
b111 6
#548310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#548320000000
0!
0%
b0 *
0-
02
b0 6
#548330000000
1!
1%
1-
12
#548340000000
0!
0%
b1 *
0-
02
b1 6
#548350000000
1!
1%
1-
12
#548360000000
0!
0%
b10 *
0-
02
b10 6
#548370000000
1!
1%
1-
12
#548380000000
0!
0%
b11 *
0-
02
b11 6
#548390000000
1!
1%
1-
12
15
#548400000000
0!
0%
b100 *
0-
02
b100 6
#548410000000
1!
1%
1-
12
#548420000000
0!
0%
b101 *
0-
02
b101 6
#548430000000
1!
1%
1-
12
#548440000000
0!
0%
b110 *
0-
02
b110 6
#548450000000
1!
1%
1-
12
#548460000000
0!
0%
b111 *
0-
02
b111 6
#548470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#548480000000
0!
0%
b0 *
0-
02
b0 6
#548490000000
1!
1%
1-
12
#548500000000
0!
0%
b1 *
0-
02
b1 6
#548510000000
1!
1%
1-
12
#548520000000
0!
0%
b10 *
0-
02
b10 6
#548530000000
1!
1%
1-
12
#548540000000
0!
0%
b11 *
0-
02
b11 6
#548550000000
1!
1%
1-
12
15
#548560000000
0!
0%
b100 *
0-
02
b100 6
#548570000000
1!
1%
1-
12
#548580000000
0!
0%
b101 *
0-
02
b101 6
#548590000000
1!
1%
1-
12
#548600000000
0!
0%
b110 *
0-
02
b110 6
#548610000000
1!
1%
1-
12
#548620000000
0!
0%
b111 *
0-
02
b111 6
#548630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#548640000000
0!
0%
b0 *
0-
02
b0 6
#548650000000
1!
1%
1-
12
#548660000000
0!
0%
b1 *
0-
02
b1 6
#548670000000
1!
1%
1-
12
#548680000000
0!
0%
b10 *
0-
02
b10 6
#548690000000
1!
1%
1-
12
#548700000000
0!
0%
b11 *
0-
02
b11 6
#548710000000
1!
1%
1-
12
15
#548720000000
0!
0%
b100 *
0-
02
b100 6
#548730000000
1!
1%
1-
12
#548740000000
0!
0%
b101 *
0-
02
b101 6
#548750000000
1!
1%
1-
12
#548760000000
0!
0%
b110 *
0-
02
b110 6
#548770000000
1!
1%
1-
12
#548780000000
0!
0%
b111 *
0-
02
b111 6
#548790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#548800000000
0!
0%
b0 *
0-
02
b0 6
#548810000000
1!
1%
1-
12
#548820000000
0!
0%
b1 *
0-
02
b1 6
#548830000000
1!
1%
1-
12
#548840000000
0!
0%
b10 *
0-
02
b10 6
#548850000000
1!
1%
1-
12
#548860000000
0!
0%
b11 *
0-
02
b11 6
#548870000000
1!
1%
1-
12
15
#548880000000
0!
0%
b100 *
0-
02
b100 6
#548890000000
1!
1%
1-
12
#548900000000
0!
0%
b101 *
0-
02
b101 6
#548910000000
1!
1%
1-
12
#548920000000
0!
0%
b110 *
0-
02
b110 6
#548930000000
1!
1%
1-
12
#548940000000
0!
0%
b111 *
0-
02
b111 6
#548950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#548960000000
0!
0%
b0 *
0-
02
b0 6
#548970000000
1!
1%
1-
12
#548980000000
0!
0%
b1 *
0-
02
b1 6
#548990000000
1!
1%
1-
12
#549000000000
0!
0%
b10 *
0-
02
b10 6
#549010000000
1!
1%
1-
12
#549020000000
0!
0%
b11 *
0-
02
b11 6
#549030000000
1!
1%
1-
12
15
#549040000000
0!
0%
b100 *
0-
02
b100 6
#549050000000
1!
1%
1-
12
#549060000000
0!
0%
b101 *
0-
02
b101 6
#549070000000
1!
1%
1-
12
#549080000000
0!
0%
b110 *
0-
02
b110 6
#549090000000
1!
1%
1-
12
#549100000000
0!
0%
b111 *
0-
02
b111 6
#549110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#549120000000
0!
0%
b0 *
0-
02
b0 6
#549130000000
1!
1%
1-
12
#549140000000
0!
0%
b1 *
0-
02
b1 6
#549150000000
1!
1%
1-
12
#549160000000
0!
0%
b10 *
0-
02
b10 6
#549170000000
1!
1%
1-
12
#549180000000
0!
0%
b11 *
0-
02
b11 6
#549190000000
1!
1%
1-
12
15
#549200000000
0!
0%
b100 *
0-
02
b100 6
#549210000000
1!
1%
1-
12
#549220000000
0!
0%
b101 *
0-
02
b101 6
#549230000000
1!
1%
1-
12
#549240000000
0!
0%
b110 *
0-
02
b110 6
#549250000000
1!
1%
1-
12
#549260000000
0!
0%
b111 *
0-
02
b111 6
#549270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#549280000000
0!
0%
b0 *
0-
02
b0 6
#549290000000
1!
1%
1-
12
#549300000000
0!
0%
b1 *
0-
02
b1 6
#549310000000
1!
1%
1-
12
#549320000000
0!
0%
b10 *
0-
02
b10 6
#549330000000
1!
1%
1-
12
#549340000000
0!
0%
b11 *
0-
02
b11 6
#549350000000
1!
1%
1-
12
15
#549360000000
0!
0%
b100 *
0-
02
b100 6
#549370000000
1!
1%
1-
12
#549380000000
0!
0%
b101 *
0-
02
b101 6
#549390000000
1!
1%
1-
12
#549400000000
0!
0%
b110 *
0-
02
b110 6
#549410000000
1!
1%
1-
12
#549420000000
0!
0%
b111 *
0-
02
b111 6
#549430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#549440000000
0!
0%
b0 *
0-
02
b0 6
#549450000000
1!
1%
1-
12
#549460000000
0!
0%
b1 *
0-
02
b1 6
#549470000000
1!
1%
1-
12
#549480000000
0!
0%
b10 *
0-
02
b10 6
#549490000000
1!
1%
1-
12
#549500000000
0!
0%
b11 *
0-
02
b11 6
#549510000000
1!
1%
1-
12
15
#549520000000
0!
0%
b100 *
0-
02
b100 6
#549530000000
1!
1%
1-
12
#549540000000
0!
0%
b101 *
0-
02
b101 6
#549550000000
1!
1%
1-
12
#549560000000
0!
0%
b110 *
0-
02
b110 6
#549570000000
1!
1%
1-
12
#549580000000
0!
0%
b111 *
0-
02
b111 6
#549590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#549600000000
0!
0%
b0 *
0-
02
b0 6
#549610000000
1!
1%
1-
12
#549620000000
0!
0%
b1 *
0-
02
b1 6
#549630000000
1!
1%
1-
12
#549640000000
0!
0%
b10 *
0-
02
b10 6
#549650000000
1!
1%
1-
12
#549660000000
0!
0%
b11 *
0-
02
b11 6
#549670000000
1!
1%
1-
12
15
#549680000000
0!
0%
b100 *
0-
02
b100 6
#549690000000
1!
1%
1-
12
#549700000000
0!
0%
b101 *
0-
02
b101 6
#549710000000
1!
1%
1-
12
#549720000000
0!
0%
b110 *
0-
02
b110 6
#549730000000
1!
1%
1-
12
#549740000000
0!
0%
b111 *
0-
02
b111 6
#549750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#549760000000
0!
0%
b0 *
0-
02
b0 6
#549770000000
1!
1%
1-
12
#549780000000
0!
0%
b1 *
0-
02
b1 6
#549790000000
1!
1%
1-
12
#549800000000
0!
0%
b10 *
0-
02
b10 6
#549810000000
1!
1%
1-
12
#549820000000
0!
0%
b11 *
0-
02
b11 6
#549830000000
1!
1%
1-
12
15
#549840000000
0!
0%
b100 *
0-
02
b100 6
#549850000000
1!
1%
1-
12
#549860000000
0!
0%
b101 *
0-
02
b101 6
#549870000000
1!
1%
1-
12
#549880000000
0!
0%
b110 *
0-
02
b110 6
#549890000000
1!
1%
1-
12
#549900000000
0!
0%
b111 *
0-
02
b111 6
#549910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#549920000000
0!
0%
b0 *
0-
02
b0 6
#549930000000
1!
1%
1-
12
#549940000000
0!
0%
b1 *
0-
02
b1 6
#549950000000
1!
1%
1-
12
#549960000000
0!
0%
b10 *
0-
02
b10 6
#549970000000
1!
1%
1-
12
#549980000000
0!
0%
b11 *
0-
02
b11 6
#549990000000
1!
1%
1-
12
15
#550000000000
0!
0%
b100 *
0-
02
b100 6
#550010000000
1!
1%
1-
12
#550020000000
0!
0%
b101 *
0-
02
b101 6
#550030000000
1!
1%
1-
12
#550040000000
0!
0%
b110 *
0-
02
b110 6
#550050000000
1!
1%
1-
12
#550060000000
0!
0%
b111 *
0-
02
b111 6
#550070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#550080000000
0!
0%
b0 *
0-
02
b0 6
#550090000000
1!
1%
1-
12
#550100000000
0!
0%
b1 *
0-
02
b1 6
#550110000000
1!
1%
1-
12
#550120000000
0!
0%
b10 *
0-
02
b10 6
#550130000000
1!
1%
1-
12
#550140000000
0!
0%
b11 *
0-
02
b11 6
#550150000000
1!
1%
1-
12
15
#550160000000
0!
0%
b100 *
0-
02
b100 6
#550170000000
1!
1%
1-
12
#550180000000
0!
0%
b101 *
0-
02
b101 6
#550190000000
1!
1%
1-
12
#550200000000
0!
0%
b110 *
0-
02
b110 6
#550210000000
1!
1%
1-
12
#550220000000
0!
0%
b111 *
0-
02
b111 6
#550230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#550240000000
0!
0%
b0 *
0-
02
b0 6
#550250000000
1!
1%
1-
12
#550260000000
0!
0%
b1 *
0-
02
b1 6
#550270000000
1!
1%
1-
12
#550280000000
0!
0%
b10 *
0-
02
b10 6
#550290000000
1!
1%
1-
12
#550300000000
0!
0%
b11 *
0-
02
b11 6
#550310000000
1!
1%
1-
12
15
#550320000000
0!
0%
b100 *
0-
02
b100 6
#550330000000
1!
1%
1-
12
#550340000000
0!
0%
b101 *
0-
02
b101 6
#550350000000
1!
1%
1-
12
#550360000000
0!
0%
b110 *
0-
02
b110 6
#550370000000
1!
1%
1-
12
#550380000000
0!
0%
b111 *
0-
02
b111 6
#550390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#550400000000
0!
0%
b0 *
0-
02
b0 6
#550410000000
1!
1%
1-
12
#550420000000
0!
0%
b1 *
0-
02
b1 6
#550430000000
1!
1%
1-
12
#550440000000
0!
0%
b10 *
0-
02
b10 6
#550450000000
1!
1%
1-
12
#550460000000
0!
0%
b11 *
0-
02
b11 6
#550470000000
1!
1%
1-
12
15
#550480000000
0!
0%
b100 *
0-
02
b100 6
#550490000000
1!
1%
1-
12
#550500000000
0!
0%
b101 *
0-
02
b101 6
#550510000000
1!
1%
1-
12
#550520000000
0!
0%
b110 *
0-
02
b110 6
#550530000000
1!
1%
1-
12
#550540000000
0!
0%
b111 *
0-
02
b111 6
#550550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#550560000000
0!
0%
b0 *
0-
02
b0 6
#550570000000
1!
1%
1-
12
#550580000000
0!
0%
b1 *
0-
02
b1 6
#550590000000
1!
1%
1-
12
#550600000000
0!
0%
b10 *
0-
02
b10 6
#550610000000
1!
1%
1-
12
#550620000000
0!
0%
b11 *
0-
02
b11 6
#550630000000
1!
1%
1-
12
15
#550640000000
0!
0%
b100 *
0-
02
b100 6
#550650000000
1!
1%
1-
12
#550660000000
0!
0%
b101 *
0-
02
b101 6
#550670000000
1!
1%
1-
12
#550680000000
0!
0%
b110 *
0-
02
b110 6
#550690000000
1!
1%
1-
12
#550700000000
0!
0%
b111 *
0-
02
b111 6
#550710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#550720000000
0!
0%
b0 *
0-
02
b0 6
#550730000000
1!
1%
1-
12
#550740000000
0!
0%
b1 *
0-
02
b1 6
#550750000000
1!
1%
1-
12
#550760000000
0!
0%
b10 *
0-
02
b10 6
#550770000000
1!
1%
1-
12
#550780000000
0!
0%
b11 *
0-
02
b11 6
#550790000000
1!
1%
1-
12
15
#550800000000
0!
0%
b100 *
0-
02
b100 6
#550810000000
1!
1%
1-
12
#550820000000
0!
0%
b101 *
0-
02
b101 6
#550830000000
1!
1%
1-
12
#550840000000
0!
0%
b110 *
0-
02
b110 6
#550850000000
1!
1%
1-
12
#550860000000
0!
0%
b111 *
0-
02
b111 6
#550870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#550880000000
0!
0%
b0 *
0-
02
b0 6
#550890000000
1!
1%
1-
12
#550900000000
0!
0%
b1 *
0-
02
b1 6
#550910000000
1!
1%
1-
12
#550920000000
0!
0%
b10 *
0-
02
b10 6
#550930000000
1!
1%
1-
12
#550940000000
0!
0%
b11 *
0-
02
b11 6
#550950000000
1!
1%
1-
12
15
#550960000000
0!
0%
b100 *
0-
02
b100 6
#550970000000
1!
1%
1-
12
#550980000000
0!
0%
b101 *
0-
02
b101 6
#550990000000
1!
1%
1-
12
#551000000000
0!
0%
b110 *
0-
02
b110 6
#551010000000
1!
1%
1-
12
#551020000000
0!
0%
b111 *
0-
02
b111 6
#551030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#551040000000
0!
0%
b0 *
0-
02
b0 6
#551050000000
1!
1%
1-
12
#551060000000
0!
0%
b1 *
0-
02
b1 6
#551070000000
1!
1%
1-
12
#551080000000
0!
0%
b10 *
0-
02
b10 6
#551090000000
1!
1%
1-
12
#551100000000
0!
0%
b11 *
0-
02
b11 6
#551110000000
1!
1%
1-
12
15
#551120000000
0!
0%
b100 *
0-
02
b100 6
#551130000000
1!
1%
1-
12
#551140000000
0!
0%
b101 *
0-
02
b101 6
#551150000000
1!
1%
1-
12
#551160000000
0!
0%
b110 *
0-
02
b110 6
#551170000000
1!
1%
1-
12
#551180000000
0!
0%
b111 *
0-
02
b111 6
#551190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#551200000000
0!
0%
b0 *
0-
02
b0 6
#551210000000
1!
1%
1-
12
#551220000000
0!
0%
b1 *
0-
02
b1 6
#551230000000
1!
1%
1-
12
#551240000000
0!
0%
b10 *
0-
02
b10 6
#551250000000
1!
1%
1-
12
#551260000000
0!
0%
b11 *
0-
02
b11 6
#551270000000
1!
1%
1-
12
15
#551280000000
0!
0%
b100 *
0-
02
b100 6
#551290000000
1!
1%
1-
12
#551300000000
0!
0%
b101 *
0-
02
b101 6
#551310000000
1!
1%
1-
12
#551320000000
0!
0%
b110 *
0-
02
b110 6
#551330000000
1!
1%
1-
12
#551340000000
0!
0%
b111 *
0-
02
b111 6
#551350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#551360000000
0!
0%
b0 *
0-
02
b0 6
#551370000000
1!
1%
1-
12
#551380000000
0!
0%
b1 *
0-
02
b1 6
#551390000000
1!
1%
1-
12
#551400000000
0!
0%
b10 *
0-
02
b10 6
#551410000000
1!
1%
1-
12
#551420000000
0!
0%
b11 *
0-
02
b11 6
#551430000000
1!
1%
1-
12
15
#551440000000
0!
0%
b100 *
0-
02
b100 6
#551450000000
1!
1%
1-
12
#551460000000
0!
0%
b101 *
0-
02
b101 6
#551470000000
1!
1%
1-
12
#551480000000
0!
0%
b110 *
0-
02
b110 6
#551490000000
1!
1%
1-
12
#551500000000
0!
0%
b111 *
0-
02
b111 6
#551510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#551520000000
0!
0%
b0 *
0-
02
b0 6
#551530000000
1!
1%
1-
12
#551540000000
0!
0%
b1 *
0-
02
b1 6
#551550000000
1!
1%
1-
12
#551560000000
0!
0%
b10 *
0-
02
b10 6
#551570000000
1!
1%
1-
12
#551580000000
0!
0%
b11 *
0-
02
b11 6
#551590000000
1!
1%
1-
12
15
#551600000000
0!
0%
b100 *
0-
02
b100 6
#551610000000
1!
1%
1-
12
#551620000000
0!
0%
b101 *
0-
02
b101 6
#551630000000
1!
1%
1-
12
#551640000000
0!
0%
b110 *
0-
02
b110 6
#551650000000
1!
1%
1-
12
#551660000000
0!
0%
b111 *
0-
02
b111 6
#551670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#551680000000
0!
0%
b0 *
0-
02
b0 6
#551690000000
1!
1%
1-
12
#551700000000
0!
0%
b1 *
0-
02
b1 6
#551710000000
1!
1%
1-
12
#551720000000
0!
0%
b10 *
0-
02
b10 6
#551730000000
1!
1%
1-
12
#551740000000
0!
0%
b11 *
0-
02
b11 6
#551750000000
1!
1%
1-
12
15
#551760000000
0!
0%
b100 *
0-
02
b100 6
#551770000000
1!
1%
1-
12
#551780000000
0!
0%
b101 *
0-
02
b101 6
#551790000000
1!
1%
1-
12
#551800000000
0!
0%
b110 *
0-
02
b110 6
#551810000000
1!
1%
1-
12
#551820000000
0!
0%
b111 *
0-
02
b111 6
#551830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#551840000000
0!
0%
b0 *
0-
02
b0 6
#551850000000
1!
1%
1-
12
#551860000000
0!
0%
b1 *
0-
02
b1 6
#551870000000
1!
1%
1-
12
#551880000000
0!
0%
b10 *
0-
02
b10 6
#551890000000
1!
1%
1-
12
#551900000000
0!
0%
b11 *
0-
02
b11 6
#551910000000
1!
1%
1-
12
15
#551920000000
0!
0%
b100 *
0-
02
b100 6
#551930000000
1!
1%
1-
12
#551940000000
0!
0%
b101 *
0-
02
b101 6
#551950000000
1!
1%
1-
12
#551960000000
0!
0%
b110 *
0-
02
b110 6
#551970000000
1!
1%
1-
12
#551980000000
0!
0%
b111 *
0-
02
b111 6
#551990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#552000000000
0!
0%
b0 *
0-
02
b0 6
#552010000000
1!
1%
1-
12
#552020000000
0!
0%
b1 *
0-
02
b1 6
#552030000000
1!
1%
1-
12
#552040000000
0!
0%
b10 *
0-
02
b10 6
#552050000000
1!
1%
1-
12
#552060000000
0!
0%
b11 *
0-
02
b11 6
#552070000000
1!
1%
1-
12
15
#552080000000
0!
0%
b100 *
0-
02
b100 6
#552090000000
1!
1%
1-
12
#552100000000
0!
0%
b101 *
0-
02
b101 6
#552110000000
1!
1%
1-
12
#552120000000
0!
0%
b110 *
0-
02
b110 6
#552130000000
1!
1%
1-
12
#552140000000
0!
0%
b111 *
0-
02
b111 6
#552150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#552160000000
0!
0%
b0 *
0-
02
b0 6
#552170000000
1!
1%
1-
12
#552180000000
0!
0%
b1 *
0-
02
b1 6
#552190000000
1!
1%
1-
12
#552200000000
0!
0%
b10 *
0-
02
b10 6
#552210000000
1!
1%
1-
12
#552220000000
0!
0%
b11 *
0-
02
b11 6
#552230000000
1!
1%
1-
12
15
#552240000000
0!
0%
b100 *
0-
02
b100 6
#552250000000
1!
1%
1-
12
#552260000000
0!
0%
b101 *
0-
02
b101 6
#552270000000
1!
1%
1-
12
#552280000000
0!
0%
b110 *
0-
02
b110 6
#552290000000
1!
1%
1-
12
#552300000000
0!
0%
b111 *
0-
02
b111 6
#552310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#552320000000
0!
0%
b0 *
0-
02
b0 6
#552330000000
1!
1%
1-
12
#552340000000
0!
0%
b1 *
0-
02
b1 6
#552350000000
1!
1%
1-
12
#552360000000
0!
0%
b10 *
0-
02
b10 6
#552370000000
1!
1%
1-
12
#552380000000
0!
0%
b11 *
0-
02
b11 6
#552390000000
1!
1%
1-
12
15
#552400000000
0!
0%
b100 *
0-
02
b100 6
#552410000000
1!
1%
1-
12
#552420000000
0!
0%
b101 *
0-
02
b101 6
#552430000000
1!
1%
1-
12
#552440000000
0!
0%
b110 *
0-
02
b110 6
#552450000000
1!
1%
1-
12
#552460000000
0!
0%
b111 *
0-
02
b111 6
#552470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#552480000000
0!
0%
b0 *
0-
02
b0 6
#552490000000
1!
1%
1-
12
#552500000000
0!
0%
b1 *
0-
02
b1 6
#552510000000
1!
1%
1-
12
#552520000000
0!
0%
b10 *
0-
02
b10 6
#552530000000
1!
1%
1-
12
#552540000000
0!
0%
b11 *
0-
02
b11 6
#552550000000
1!
1%
1-
12
15
#552560000000
0!
0%
b100 *
0-
02
b100 6
#552570000000
1!
1%
1-
12
#552580000000
0!
0%
b101 *
0-
02
b101 6
#552590000000
1!
1%
1-
12
#552600000000
0!
0%
b110 *
0-
02
b110 6
#552610000000
1!
1%
1-
12
#552620000000
0!
0%
b111 *
0-
02
b111 6
#552630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#552640000000
0!
0%
b0 *
0-
02
b0 6
#552650000000
1!
1%
1-
12
#552660000000
0!
0%
b1 *
0-
02
b1 6
#552670000000
1!
1%
1-
12
#552680000000
0!
0%
b10 *
0-
02
b10 6
#552690000000
1!
1%
1-
12
#552700000000
0!
0%
b11 *
0-
02
b11 6
#552710000000
1!
1%
1-
12
15
#552720000000
0!
0%
b100 *
0-
02
b100 6
#552730000000
1!
1%
1-
12
#552740000000
0!
0%
b101 *
0-
02
b101 6
#552750000000
1!
1%
1-
12
#552760000000
0!
0%
b110 *
0-
02
b110 6
#552770000000
1!
1%
1-
12
#552780000000
0!
0%
b111 *
0-
02
b111 6
#552790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#552800000000
0!
0%
b0 *
0-
02
b0 6
#552810000000
1!
1%
1-
12
#552820000000
0!
0%
b1 *
0-
02
b1 6
#552830000000
1!
1%
1-
12
#552840000000
0!
0%
b10 *
0-
02
b10 6
#552850000000
1!
1%
1-
12
#552860000000
0!
0%
b11 *
0-
02
b11 6
#552870000000
1!
1%
1-
12
15
#552880000000
0!
0%
b100 *
0-
02
b100 6
#552890000000
1!
1%
1-
12
#552900000000
0!
0%
b101 *
0-
02
b101 6
#552910000000
1!
1%
1-
12
#552920000000
0!
0%
b110 *
0-
02
b110 6
#552930000000
1!
1%
1-
12
#552940000000
0!
0%
b111 *
0-
02
b111 6
#552950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#552960000000
0!
0%
b0 *
0-
02
b0 6
#552970000000
1!
1%
1-
12
#552980000000
0!
0%
b1 *
0-
02
b1 6
#552990000000
1!
1%
1-
12
#553000000000
0!
0%
b10 *
0-
02
b10 6
#553010000000
1!
1%
1-
12
#553020000000
0!
0%
b11 *
0-
02
b11 6
#553030000000
1!
1%
1-
12
15
#553040000000
0!
0%
b100 *
0-
02
b100 6
#553050000000
1!
1%
1-
12
#553060000000
0!
0%
b101 *
0-
02
b101 6
#553070000000
1!
1%
1-
12
#553080000000
0!
0%
b110 *
0-
02
b110 6
#553090000000
1!
1%
1-
12
#553100000000
0!
0%
b111 *
0-
02
b111 6
#553110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#553120000000
0!
0%
b0 *
0-
02
b0 6
#553130000000
1!
1%
1-
12
#553140000000
0!
0%
b1 *
0-
02
b1 6
#553150000000
1!
1%
1-
12
#553160000000
0!
0%
b10 *
0-
02
b10 6
#553170000000
1!
1%
1-
12
#553180000000
0!
0%
b11 *
0-
02
b11 6
#553190000000
1!
1%
1-
12
15
#553200000000
0!
0%
b100 *
0-
02
b100 6
#553210000000
1!
1%
1-
12
#553220000000
0!
0%
b101 *
0-
02
b101 6
#553230000000
1!
1%
1-
12
#553240000000
0!
0%
b110 *
0-
02
b110 6
#553250000000
1!
1%
1-
12
#553260000000
0!
0%
b111 *
0-
02
b111 6
#553270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#553280000000
0!
0%
b0 *
0-
02
b0 6
#553290000000
1!
1%
1-
12
#553300000000
0!
0%
b1 *
0-
02
b1 6
#553310000000
1!
1%
1-
12
#553320000000
0!
0%
b10 *
0-
02
b10 6
#553330000000
1!
1%
1-
12
#553340000000
0!
0%
b11 *
0-
02
b11 6
#553350000000
1!
1%
1-
12
15
#553360000000
0!
0%
b100 *
0-
02
b100 6
#553370000000
1!
1%
1-
12
#553380000000
0!
0%
b101 *
0-
02
b101 6
#553390000000
1!
1%
1-
12
#553400000000
0!
0%
b110 *
0-
02
b110 6
#553410000000
1!
1%
1-
12
#553420000000
0!
0%
b111 *
0-
02
b111 6
#553430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#553440000000
0!
0%
b0 *
0-
02
b0 6
#553450000000
1!
1%
1-
12
#553460000000
0!
0%
b1 *
0-
02
b1 6
#553470000000
1!
1%
1-
12
#553480000000
0!
0%
b10 *
0-
02
b10 6
#553490000000
1!
1%
1-
12
#553500000000
0!
0%
b11 *
0-
02
b11 6
#553510000000
1!
1%
1-
12
15
#553520000000
0!
0%
b100 *
0-
02
b100 6
#553530000000
1!
1%
1-
12
#553540000000
0!
0%
b101 *
0-
02
b101 6
#553550000000
1!
1%
1-
12
#553560000000
0!
0%
b110 *
0-
02
b110 6
#553570000000
1!
1%
1-
12
#553580000000
0!
0%
b111 *
0-
02
b111 6
#553590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#553600000000
0!
0%
b0 *
0-
02
b0 6
#553610000000
1!
1%
1-
12
#553620000000
0!
0%
b1 *
0-
02
b1 6
#553630000000
1!
1%
1-
12
#553640000000
0!
0%
b10 *
0-
02
b10 6
#553650000000
1!
1%
1-
12
#553660000000
0!
0%
b11 *
0-
02
b11 6
#553670000000
1!
1%
1-
12
15
#553680000000
0!
0%
b100 *
0-
02
b100 6
#553690000000
1!
1%
1-
12
#553700000000
0!
0%
b101 *
0-
02
b101 6
#553710000000
1!
1%
1-
12
#553720000000
0!
0%
b110 *
0-
02
b110 6
#553730000000
1!
1%
1-
12
#553740000000
0!
0%
b111 *
0-
02
b111 6
#553750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#553760000000
0!
0%
b0 *
0-
02
b0 6
#553770000000
1!
1%
1-
12
#553780000000
0!
0%
b1 *
0-
02
b1 6
#553790000000
1!
1%
1-
12
#553800000000
0!
0%
b10 *
0-
02
b10 6
#553810000000
1!
1%
1-
12
#553820000000
0!
0%
b11 *
0-
02
b11 6
#553830000000
1!
1%
1-
12
15
#553840000000
0!
0%
b100 *
0-
02
b100 6
#553850000000
1!
1%
1-
12
#553860000000
0!
0%
b101 *
0-
02
b101 6
#553870000000
1!
1%
1-
12
#553880000000
0!
0%
b110 *
0-
02
b110 6
#553890000000
1!
1%
1-
12
#553900000000
0!
0%
b111 *
0-
02
b111 6
#553910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#553920000000
0!
0%
b0 *
0-
02
b0 6
#553930000000
1!
1%
1-
12
#553940000000
0!
0%
b1 *
0-
02
b1 6
#553950000000
1!
1%
1-
12
#553960000000
0!
0%
b10 *
0-
02
b10 6
#553970000000
1!
1%
1-
12
#553980000000
0!
0%
b11 *
0-
02
b11 6
#553990000000
1!
1%
1-
12
15
#554000000000
0!
0%
b100 *
0-
02
b100 6
#554010000000
1!
1%
1-
12
#554020000000
0!
0%
b101 *
0-
02
b101 6
#554030000000
1!
1%
1-
12
#554040000000
0!
0%
b110 *
0-
02
b110 6
#554050000000
1!
1%
1-
12
#554060000000
0!
0%
b111 *
0-
02
b111 6
#554070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#554080000000
0!
0%
b0 *
0-
02
b0 6
#554090000000
1!
1%
1-
12
#554100000000
0!
0%
b1 *
0-
02
b1 6
#554110000000
1!
1%
1-
12
#554120000000
0!
0%
b10 *
0-
02
b10 6
#554130000000
1!
1%
1-
12
#554140000000
0!
0%
b11 *
0-
02
b11 6
#554150000000
1!
1%
1-
12
15
#554160000000
0!
0%
b100 *
0-
02
b100 6
#554170000000
1!
1%
1-
12
#554180000000
0!
0%
b101 *
0-
02
b101 6
#554190000000
1!
1%
1-
12
#554200000000
0!
0%
b110 *
0-
02
b110 6
#554210000000
1!
1%
1-
12
#554220000000
0!
0%
b111 *
0-
02
b111 6
#554230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#554240000000
0!
0%
b0 *
0-
02
b0 6
#554250000000
1!
1%
1-
12
#554260000000
0!
0%
b1 *
0-
02
b1 6
#554270000000
1!
1%
1-
12
#554280000000
0!
0%
b10 *
0-
02
b10 6
#554290000000
1!
1%
1-
12
#554300000000
0!
0%
b11 *
0-
02
b11 6
#554310000000
1!
1%
1-
12
15
#554320000000
0!
0%
b100 *
0-
02
b100 6
#554330000000
1!
1%
1-
12
#554340000000
0!
0%
b101 *
0-
02
b101 6
#554350000000
1!
1%
1-
12
#554360000000
0!
0%
b110 *
0-
02
b110 6
#554370000000
1!
1%
1-
12
#554380000000
0!
0%
b111 *
0-
02
b111 6
#554390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#554400000000
0!
0%
b0 *
0-
02
b0 6
#554410000000
1!
1%
1-
12
#554420000000
0!
0%
b1 *
0-
02
b1 6
#554430000000
1!
1%
1-
12
#554440000000
0!
0%
b10 *
0-
02
b10 6
#554450000000
1!
1%
1-
12
#554460000000
0!
0%
b11 *
0-
02
b11 6
#554470000000
1!
1%
1-
12
15
#554480000000
0!
0%
b100 *
0-
02
b100 6
#554490000000
1!
1%
1-
12
#554500000000
0!
0%
b101 *
0-
02
b101 6
#554510000000
1!
1%
1-
12
#554520000000
0!
0%
b110 *
0-
02
b110 6
#554530000000
1!
1%
1-
12
#554540000000
0!
0%
b111 *
0-
02
b111 6
#554550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#554560000000
0!
0%
b0 *
0-
02
b0 6
#554570000000
1!
1%
1-
12
#554580000000
0!
0%
b1 *
0-
02
b1 6
#554590000000
1!
1%
1-
12
#554600000000
0!
0%
b10 *
0-
02
b10 6
#554610000000
1!
1%
1-
12
#554620000000
0!
0%
b11 *
0-
02
b11 6
#554630000000
1!
1%
1-
12
15
#554640000000
0!
0%
b100 *
0-
02
b100 6
#554650000000
1!
1%
1-
12
#554660000000
0!
0%
b101 *
0-
02
b101 6
#554670000000
1!
1%
1-
12
#554680000000
0!
0%
b110 *
0-
02
b110 6
#554690000000
1!
1%
1-
12
#554700000000
0!
0%
b111 *
0-
02
b111 6
#554710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#554720000000
0!
0%
b0 *
0-
02
b0 6
#554730000000
1!
1%
1-
12
#554740000000
0!
0%
b1 *
0-
02
b1 6
#554750000000
1!
1%
1-
12
#554760000000
0!
0%
b10 *
0-
02
b10 6
#554770000000
1!
1%
1-
12
#554780000000
0!
0%
b11 *
0-
02
b11 6
#554790000000
1!
1%
1-
12
15
#554800000000
0!
0%
b100 *
0-
02
b100 6
#554810000000
1!
1%
1-
12
#554820000000
0!
0%
b101 *
0-
02
b101 6
#554830000000
1!
1%
1-
12
#554840000000
0!
0%
b110 *
0-
02
b110 6
#554850000000
1!
1%
1-
12
#554860000000
0!
0%
b111 *
0-
02
b111 6
#554870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#554880000000
0!
0%
b0 *
0-
02
b0 6
#554890000000
1!
1%
1-
12
#554900000000
0!
0%
b1 *
0-
02
b1 6
#554910000000
1!
1%
1-
12
#554920000000
0!
0%
b10 *
0-
02
b10 6
#554930000000
1!
1%
1-
12
#554940000000
0!
0%
b11 *
0-
02
b11 6
#554950000000
1!
1%
1-
12
15
#554960000000
0!
0%
b100 *
0-
02
b100 6
#554970000000
1!
1%
1-
12
#554980000000
0!
0%
b101 *
0-
02
b101 6
#554990000000
1!
1%
1-
12
#555000000000
0!
0%
b110 *
0-
02
b110 6
#555010000000
1!
1%
1-
12
#555020000000
0!
0%
b111 *
0-
02
b111 6
#555030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#555040000000
0!
0%
b0 *
0-
02
b0 6
#555050000000
1!
1%
1-
12
#555060000000
0!
0%
b1 *
0-
02
b1 6
#555070000000
1!
1%
1-
12
#555080000000
0!
0%
b10 *
0-
02
b10 6
#555090000000
1!
1%
1-
12
#555100000000
0!
0%
b11 *
0-
02
b11 6
#555110000000
1!
1%
1-
12
15
#555120000000
0!
0%
b100 *
0-
02
b100 6
#555130000000
1!
1%
1-
12
#555140000000
0!
0%
b101 *
0-
02
b101 6
#555150000000
1!
1%
1-
12
#555160000000
0!
0%
b110 *
0-
02
b110 6
#555170000000
1!
1%
1-
12
#555180000000
0!
0%
b111 *
0-
02
b111 6
#555190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#555200000000
0!
0%
b0 *
0-
02
b0 6
#555210000000
1!
1%
1-
12
#555220000000
0!
0%
b1 *
0-
02
b1 6
#555230000000
1!
1%
1-
12
#555240000000
0!
0%
b10 *
0-
02
b10 6
#555250000000
1!
1%
1-
12
#555260000000
0!
0%
b11 *
0-
02
b11 6
#555270000000
1!
1%
1-
12
15
#555280000000
0!
0%
b100 *
0-
02
b100 6
#555290000000
1!
1%
1-
12
#555300000000
0!
0%
b101 *
0-
02
b101 6
#555310000000
1!
1%
1-
12
#555320000000
0!
0%
b110 *
0-
02
b110 6
#555330000000
1!
1%
1-
12
#555340000000
0!
0%
b111 *
0-
02
b111 6
#555350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#555360000000
0!
0%
b0 *
0-
02
b0 6
#555370000000
1!
1%
1-
12
#555380000000
0!
0%
b1 *
0-
02
b1 6
#555390000000
1!
1%
1-
12
#555400000000
0!
0%
b10 *
0-
02
b10 6
#555410000000
1!
1%
1-
12
#555420000000
0!
0%
b11 *
0-
02
b11 6
#555430000000
1!
1%
1-
12
15
#555440000000
0!
0%
b100 *
0-
02
b100 6
#555450000000
1!
1%
1-
12
#555460000000
0!
0%
b101 *
0-
02
b101 6
#555470000000
1!
1%
1-
12
#555480000000
0!
0%
b110 *
0-
02
b110 6
#555490000000
1!
1%
1-
12
#555500000000
0!
0%
b111 *
0-
02
b111 6
#555510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#555520000000
0!
0%
b0 *
0-
02
b0 6
#555530000000
1!
1%
1-
12
#555540000000
0!
0%
b1 *
0-
02
b1 6
#555550000000
1!
1%
1-
12
#555560000000
0!
0%
b10 *
0-
02
b10 6
#555570000000
1!
1%
1-
12
#555580000000
0!
0%
b11 *
0-
02
b11 6
#555590000000
1!
1%
1-
12
15
#555600000000
0!
0%
b100 *
0-
02
b100 6
#555610000000
1!
1%
1-
12
#555620000000
0!
0%
b101 *
0-
02
b101 6
#555630000000
1!
1%
1-
12
#555640000000
0!
0%
b110 *
0-
02
b110 6
#555650000000
1!
1%
1-
12
#555660000000
0!
0%
b111 *
0-
02
b111 6
#555670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#555680000000
0!
0%
b0 *
0-
02
b0 6
#555690000000
1!
1%
1-
12
#555700000000
0!
0%
b1 *
0-
02
b1 6
#555710000000
1!
1%
1-
12
#555720000000
0!
0%
b10 *
0-
02
b10 6
#555730000000
1!
1%
1-
12
#555740000000
0!
0%
b11 *
0-
02
b11 6
#555750000000
1!
1%
1-
12
15
#555760000000
0!
0%
b100 *
0-
02
b100 6
#555770000000
1!
1%
1-
12
#555780000000
0!
0%
b101 *
0-
02
b101 6
#555790000000
1!
1%
1-
12
#555800000000
0!
0%
b110 *
0-
02
b110 6
#555810000000
1!
1%
1-
12
#555820000000
0!
0%
b111 *
0-
02
b111 6
#555830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#555840000000
0!
0%
b0 *
0-
02
b0 6
#555850000000
1!
1%
1-
12
#555860000000
0!
0%
b1 *
0-
02
b1 6
#555870000000
1!
1%
1-
12
#555880000000
0!
0%
b10 *
0-
02
b10 6
#555890000000
1!
1%
1-
12
#555900000000
0!
0%
b11 *
0-
02
b11 6
#555910000000
1!
1%
1-
12
15
#555920000000
0!
0%
b100 *
0-
02
b100 6
#555930000000
1!
1%
1-
12
#555940000000
0!
0%
b101 *
0-
02
b101 6
#555950000000
1!
1%
1-
12
#555960000000
0!
0%
b110 *
0-
02
b110 6
#555970000000
1!
1%
1-
12
#555980000000
0!
0%
b111 *
0-
02
b111 6
#555990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#556000000000
0!
0%
b0 *
0-
02
b0 6
#556010000000
1!
1%
1-
12
#556020000000
0!
0%
b1 *
0-
02
b1 6
#556030000000
1!
1%
1-
12
#556040000000
0!
0%
b10 *
0-
02
b10 6
#556050000000
1!
1%
1-
12
#556060000000
0!
0%
b11 *
0-
02
b11 6
#556070000000
1!
1%
1-
12
15
#556080000000
0!
0%
b100 *
0-
02
b100 6
#556090000000
1!
1%
1-
12
#556100000000
0!
0%
b101 *
0-
02
b101 6
#556110000000
1!
1%
1-
12
#556120000000
0!
0%
b110 *
0-
02
b110 6
#556130000000
1!
1%
1-
12
#556140000000
0!
0%
b111 *
0-
02
b111 6
#556150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#556160000000
0!
0%
b0 *
0-
02
b0 6
#556170000000
1!
1%
1-
12
#556180000000
0!
0%
b1 *
0-
02
b1 6
#556190000000
1!
1%
1-
12
#556200000000
0!
0%
b10 *
0-
02
b10 6
#556210000000
1!
1%
1-
12
#556220000000
0!
0%
b11 *
0-
02
b11 6
#556230000000
1!
1%
1-
12
15
#556240000000
0!
0%
b100 *
0-
02
b100 6
#556250000000
1!
1%
1-
12
#556260000000
0!
0%
b101 *
0-
02
b101 6
#556270000000
1!
1%
1-
12
#556280000000
0!
0%
b110 *
0-
02
b110 6
#556290000000
1!
1%
1-
12
#556300000000
0!
0%
b111 *
0-
02
b111 6
#556310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#556320000000
0!
0%
b0 *
0-
02
b0 6
#556330000000
1!
1%
1-
12
#556340000000
0!
0%
b1 *
0-
02
b1 6
#556350000000
1!
1%
1-
12
#556360000000
0!
0%
b10 *
0-
02
b10 6
#556370000000
1!
1%
1-
12
#556380000000
0!
0%
b11 *
0-
02
b11 6
#556390000000
1!
1%
1-
12
15
#556400000000
0!
0%
b100 *
0-
02
b100 6
#556410000000
1!
1%
1-
12
#556420000000
0!
0%
b101 *
0-
02
b101 6
#556430000000
1!
1%
1-
12
#556440000000
0!
0%
b110 *
0-
02
b110 6
#556450000000
1!
1%
1-
12
#556460000000
0!
0%
b111 *
0-
02
b111 6
#556470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#556480000000
0!
0%
b0 *
0-
02
b0 6
#556490000000
1!
1%
1-
12
#556500000000
0!
0%
b1 *
0-
02
b1 6
#556510000000
1!
1%
1-
12
#556520000000
0!
0%
b10 *
0-
02
b10 6
#556530000000
1!
1%
1-
12
#556540000000
0!
0%
b11 *
0-
02
b11 6
#556550000000
1!
1%
1-
12
15
#556560000000
0!
0%
b100 *
0-
02
b100 6
#556570000000
1!
1%
1-
12
#556580000000
0!
0%
b101 *
0-
02
b101 6
#556590000000
1!
1%
1-
12
#556600000000
0!
0%
b110 *
0-
02
b110 6
#556610000000
1!
1%
1-
12
#556620000000
0!
0%
b111 *
0-
02
b111 6
#556630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#556640000000
0!
0%
b0 *
0-
02
b0 6
#556650000000
1!
1%
1-
12
#556660000000
0!
0%
b1 *
0-
02
b1 6
#556670000000
1!
1%
1-
12
#556680000000
0!
0%
b10 *
0-
02
b10 6
#556690000000
1!
1%
1-
12
#556700000000
0!
0%
b11 *
0-
02
b11 6
#556710000000
1!
1%
1-
12
15
#556720000000
0!
0%
b100 *
0-
02
b100 6
#556730000000
1!
1%
1-
12
#556740000000
0!
0%
b101 *
0-
02
b101 6
#556750000000
1!
1%
1-
12
#556760000000
0!
0%
b110 *
0-
02
b110 6
#556770000000
1!
1%
1-
12
#556780000000
0!
0%
b111 *
0-
02
b111 6
#556790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#556800000000
0!
0%
b0 *
0-
02
b0 6
#556810000000
1!
1%
1-
12
#556820000000
0!
0%
b1 *
0-
02
b1 6
#556830000000
1!
1%
1-
12
#556840000000
0!
0%
b10 *
0-
02
b10 6
#556850000000
1!
1%
1-
12
#556860000000
0!
0%
b11 *
0-
02
b11 6
#556870000000
1!
1%
1-
12
15
#556880000000
0!
0%
b100 *
0-
02
b100 6
#556890000000
1!
1%
1-
12
#556900000000
0!
0%
b101 *
0-
02
b101 6
#556910000000
1!
1%
1-
12
#556920000000
0!
0%
b110 *
0-
02
b110 6
#556930000000
1!
1%
1-
12
#556940000000
0!
0%
b111 *
0-
02
b111 6
#556950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#556960000000
0!
0%
b0 *
0-
02
b0 6
#556970000000
1!
1%
1-
12
#556980000000
0!
0%
b1 *
0-
02
b1 6
#556990000000
1!
1%
1-
12
#557000000000
0!
0%
b10 *
0-
02
b10 6
#557010000000
1!
1%
1-
12
#557020000000
0!
0%
b11 *
0-
02
b11 6
#557030000000
1!
1%
1-
12
15
#557040000000
0!
0%
b100 *
0-
02
b100 6
#557050000000
1!
1%
1-
12
#557060000000
0!
0%
b101 *
0-
02
b101 6
#557070000000
1!
1%
1-
12
#557080000000
0!
0%
b110 *
0-
02
b110 6
#557090000000
1!
1%
1-
12
#557100000000
0!
0%
b111 *
0-
02
b111 6
#557110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#557120000000
0!
0%
b0 *
0-
02
b0 6
#557130000000
1!
1%
1-
12
#557140000000
0!
0%
b1 *
0-
02
b1 6
#557150000000
1!
1%
1-
12
#557160000000
0!
0%
b10 *
0-
02
b10 6
#557170000000
1!
1%
1-
12
#557180000000
0!
0%
b11 *
0-
02
b11 6
#557190000000
1!
1%
1-
12
15
#557200000000
0!
0%
b100 *
0-
02
b100 6
#557210000000
1!
1%
1-
12
#557220000000
0!
0%
b101 *
0-
02
b101 6
#557230000000
1!
1%
1-
12
#557240000000
0!
0%
b110 *
0-
02
b110 6
#557250000000
1!
1%
1-
12
#557260000000
0!
0%
b111 *
0-
02
b111 6
#557270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#557280000000
0!
0%
b0 *
0-
02
b0 6
#557290000000
1!
1%
1-
12
#557300000000
0!
0%
b1 *
0-
02
b1 6
#557310000000
1!
1%
1-
12
#557320000000
0!
0%
b10 *
0-
02
b10 6
#557330000000
1!
1%
1-
12
#557340000000
0!
0%
b11 *
0-
02
b11 6
#557350000000
1!
1%
1-
12
15
#557360000000
0!
0%
b100 *
0-
02
b100 6
#557370000000
1!
1%
1-
12
#557380000000
0!
0%
b101 *
0-
02
b101 6
#557390000000
1!
1%
1-
12
#557400000000
0!
0%
b110 *
0-
02
b110 6
#557410000000
1!
1%
1-
12
#557420000000
0!
0%
b111 *
0-
02
b111 6
#557430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#557440000000
0!
0%
b0 *
0-
02
b0 6
#557450000000
1!
1%
1-
12
#557460000000
0!
0%
b1 *
0-
02
b1 6
#557470000000
1!
1%
1-
12
#557480000000
0!
0%
b10 *
0-
02
b10 6
#557490000000
1!
1%
1-
12
#557500000000
0!
0%
b11 *
0-
02
b11 6
#557510000000
1!
1%
1-
12
15
#557520000000
0!
0%
b100 *
0-
02
b100 6
#557530000000
1!
1%
1-
12
#557540000000
0!
0%
b101 *
0-
02
b101 6
#557550000000
1!
1%
1-
12
#557560000000
0!
0%
b110 *
0-
02
b110 6
#557570000000
1!
1%
1-
12
#557580000000
0!
0%
b111 *
0-
02
b111 6
#557590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#557600000000
0!
0%
b0 *
0-
02
b0 6
#557610000000
1!
1%
1-
12
#557620000000
0!
0%
b1 *
0-
02
b1 6
#557630000000
1!
1%
1-
12
#557640000000
0!
0%
b10 *
0-
02
b10 6
#557650000000
1!
1%
1-
12
#557660000000
0!
0%
b11 *
0-
02
b11 6
#557670000000
1!
1%
1-
12
15
#557680000000
0!
0%
b100 *
0-
02
b100 6
#557690000000
1!
1%
1-
12
#557700000000
0!
0%
b101 *
0-
02
b101 6
#557710000000
1!
1%
1-
12
#557720000000
0!
0%
b110 *
0-
02
b110 6
#557730000000
1!
1%
1-
12
#557740000000
0!
0%
b111 *
0-
02
b111 6
#557750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#557760000000
0!
0%
b0 *
0-
02
b0 6
#557770000000
1!
1%
1-
12
#557780000000
0!
0%
b1 *
0-
02
b1 6
#557790000000
1!
1%
1-
12
#557800000000
0!
0%
b10 *
0-
02
b10 6
#557810000000
1!
1%
1-
12
#557820000000
0!
0%
b11 *
0-
02
b11 6
#557830000000
1!
1%
1-
12
15
#557840000000
0!
0%
b100 *
0-
02
b100 6
#557850000000
1!
1%
1-
12
#557860000000
0!
0%
b101 *
0-
02
b101 6
#557870000000
1!
1%
1-
12
#557880000000
0!
0%
b110 *
0-
02
b110 6
#557890000000
1!
1%
1-
12
#557900000000
0!
0%
b111 *
0-
02
b111 6
#557910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#557920000000
0!
0%
b0 *
0-
02
b0 6
#557930000000
1!
1%
1-
12
#557940000000
0!
0%
b1 *
0-
02
b1 6
#557950000000
1!
1%
1-
12
#557960000000
0!
0%
b10 *
0-
02
b10 6
#557970000000
1!
1%
1-
12
#557980000000
0!
0%
b11 *
0-
02
b11 6
#557990000000
1!
1%
1-
12
15
#558000000000
0!
0%
b100 *
0-
02
b100 6
#558010000000
1!
1%
1-
12
#558020000000
0!
0%
b101 *
0-
02
b101 6
#558030000000
1!
1%
1-
12
#558040000000
0!
0%
b110 *
0-
02
b110 6
#558050000000
1!
1%
1-
12
#558060000000
0!
0%
b111 *
0-
02
b111 6
#558070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#558080000000
0!
0%
b0 *
0-
02
b0 6
#558090000000
1!
1%
1-
12
#558100000000
0!
0%
b1 *
0-
02
b1 6
#558110000000
1!
1%
1-
12
#558120000000
0!
0%
b10 *
0-
02
b10 6
#558130000000
1!
1%
1-
12
#558140000000
0!
0%
b11 *
0-
02
b11 6
#558150000000
1!
1%
1-
12
15
#558160000000
0!
0%
b100 *
0-
02
b100 6
#558170000000
1!
1%
1-
12
#558180000000
0!
0%
b101 *
0-
02
b101 6
#558190000000
1!
1%
1-
12
#558200000000
0!
0%
b110 *
0-
02
b110 6
#558210000000
1!
1%
1-
12
#558220000000
0!
0%
b111 *
0-
02
b111 6
#558230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#558240000000
0!
0%
b0 *
0-
02
b0 6
#558250000000
1!
1%
1-
12
#558260000000
0!
0%
b1 *
0-
02
b1 6
#558270000000
1!
1%
1-
12
#558280000000
0!
0%
b10 *
0-
02
b10 6
#558290000000
1!
1%
1-
12
#558300000000
0!
0%
b11 *
0-
02
b11 6
#558310000000
1!
1%
1-
12
15
#558320000000
0!
0%
b100 *
0-
02
b100 6
#558330000000
1!
1%
1-
12
#558340000000
0!
0%
b101 *
0-
02
b101 6
#558350000000
1!
1%
1-
12
#558360000000
0!
0%
b110 *
0-
02
b110 6
#558370000000
1!
1%
1-
12
#558380000000
0!
0%
b111 *
0-
02
b111 6
#558390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#558400000000
0!
0%
b0 *
0-
02
b0 6
#558410000000
1!
1%
1-
12
#558420000000
0!
0%
b1 *
0-
02
b1 6
#558430000000
1!
1%
1-
12
#558440000000
0!
0%
b10 *
0-
02
b10 6
#558450000000
1!
1%
1-
12
#558460000000
0!
0%
b11 *
0-
02
b11 6
#558470000000
1!
1%
1-
12
15
#558480000000
0!
0%
b100 *
0-
02
b100 6
#558490000000
1!
1%
1-
12
#558500000000
0!
0%
b101 *
0-
02
b101 6
#558510000000
1!
1%
1-
12
#558520000000
0!
0%
b110 *
0-
02
b110 6
#558530000000
1!
1%
1-
12
#558540000000
0!
0%
b111 *
0-
02
b111 6
#558550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#558560000000
0!
0%
b0 *
0-
02
b0 6
#558570000000
1!
1%
1-
12
#558580000000
0!
0%
b1 *
0-
02
b1 6
#558590000000
1!
1%
1-
12
#558600000000
0!
0%
b10 *
0-
02
b10 6
#558610000000
1!
1%
1-
12
#558620000000
0!
0%
b11 *
0-
02
b11 6
#558630000000
1!
1%
1-
12
15
#558640000000
0!
0%
b100 *
0-
02
b100 6
#558650000000
1!
1%
1-
12
#558660000000
0!
0%
b101 *
0-
02
b101 6
#558670000000
1!
1%
1-
12
#558680000000
0!
0%
b110 *
0-
02
b110 6
#558690000000
1!
1%
1-
12
#558700000000
0!
0%
b111 *
0-
02
b111 6
#558710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#558720000000
0!
0%
b0 *
0-
02
b0 6
#558730000000
1!
1%
1-
12
#558740000000
0!
0%
b1 *
0-
02
b1 6
#558750000000
1!
1%
1-
12
#558760000000
0!
0%
b10 *
0-
02
b10 6
#558770000000
1!
1%
1-
12
#558780000000
0!
0%
b11 *
0-
02
b11 6
#558790000000
1!
1%
1-
12
15
#558800000000
0!
0%
b100 *
0-
02
b100 6
#558810000000
1!
1%
1-
12
#558820000000
0!
0%
b101 *
0-
02
b101 6
#558830000000
1!
1%
1-
12
#558840000000
0!
0%
b110 *
0-
02
b110 6
#558850000000
1!
1%
1-
12
#558860000000
0!
0%
b111 *
0-
02
b111 6
#558870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#558880000000
0!
0%
b0 *
0-
02
b0 6
#558890000000
1!
1%
1-
12
#558900000000
0!
0%
b1 *
0-
02
b1 6
#558910000000
1!
1%
1-
12
#558920000000
0!
0%
b10 *
0-
02
b10 6
#558930000000
1!
1%
1-
12
#558940000000
0!
0%
b11 *
0-
02
b11 6
#558950000000
1!
1%
1-
12
15
#558960000000
0!
0%
b100 *
0-
02
b100 6
#558970000000
1!
1%
1-
12
#558980000000
0!
0%
b101 *
0-
02
b101 6
#558990000000
1!
1%
1-
12
#559000000000
0!
0%
b110 *
0-
02
b110 6
#559010000000
1!
1%
1-
12
#559020000000
0!
0%
b111 *
0-
02
b111 6
#559030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#559040000000
0!
0%
b0 *
0-
02
b0 6
#559050000000
1!
1%
1-
12
#559060000000
0!
0%
b1 *
0-
02
b1 6
#559070000000
1!
1%
1-
12
#559080000000
0!
0%
b10 *
0-
02
b10 6
#559090000000
1!
1%
1-
12
#559100000000
0!
0%
b11 *
0-
02
b11 6
#559110000000
1!
1%
1-
12
15
#559120000000
0!
0%
b100 *
0-
02
b100 6
#559130000000
1!
1%
1-
12
#559140000000
0!
0%
b101 *
0-
02
b101 6
#559150000000
1!
1%
1-
12
#559160000000
0!
0%
b110 *
0-
02
b110 6
#559170000000
1!
1%
1-
12
#559180000000
0!
0%
b111 *
0-
02
b111 6
#559190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#559200000000
0!
0%
b0 *
0-
02
b0 6
#559210000000
1!
1%
1-
12
#559220000000
0!
0%
b1 *
0-
02
b1 6
#559230000000
1!
1%
1-
12
#559240000000
0!
0%
b10 *
0-
02
b10 6
#559250000000
1!
1%
1-
12
#559260000000
0!
0%
b11 *
0-
02
b11 6
#559270000000
1!
1%
1-
12
15
#559280000000
0!
0%
b100 *
0-
02
b100 6
#559290000000
1!
1%
1-
12
#559300000000
0!
0%
b101 *
0-
02
b101 6
#559310000000
1!
1%
1-
12
#559320000000
0!
0%
b110 *
0-
02
b110 6
#559330000000
1!
1%
1-
12
#559340000000
0!
0%
b111 *
0-
02
b111 6
#559350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#559360000000
0!
0%
b0 *
0-
02
b0 6
#559370000000
1!
1%
1-
12
#559380000000
0!
0%
b1 *
0-
02
b1 6
#559390000000
1!
1%
1-
12
#559400000000
0!
0%
b10 *
0-
02
b10 6
#559410000000
1!
1%
1-
12
#559420000000
0!
0%
b11 *
0-
02
b11 6
#559430000000
1!
1%
1-
12
15
#559440000000
0!
0%
b100 *
0-
02
b100 6
#559450000000
1!
1%
1-
12
#559460000000
0!
0%
b101 *
0-
02
b101 6
#559470000000
1!
1%
1-
12
#559480000000
0!
0%
b110 *
0-
02
b110 6
#559490000000
1!
1%
1-
12
#559500000000
0!
0%
b111 *
0-
02
b111 6
#559510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#559520000000
0!
0%
b0 *
0-
02
b0 6
#559530000000
1!
1%
1-
12
#559540000000
0!
0%
b1 *
0-
02
b1 6
#559550000000
1!
1%
1-
12
#559560000000
0!
0%
b10 *
0-
02
b10 6
#559570000000
1!
1%
1-
12
#559580000000
0!
0%
b11 *
0-
02
b11 6
#559590000000
1!
1%
1-
12
15
#559600000000
0!
0%
b100 *
0-
02
b100 6
#559610000000
1!
1%
1-
12
#559620000000
0!
0%
b101 *
0-
02
b101 6
#559630000000
1!
1%
1-
12
#559640000000
0!
0%
b110 *
0-
02
b110 6
#559650000000
1!
1%
1-
12
#559660000000
0!
0%
b111 *
0-
02
b111 6
#559670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#559680000000
0!
0%
b0 *
0-
02
b0 6
#559690000000
1!
1%
1-
12
#559700000000
0!
0%
b1 *
0-
02
b1 6
#559710000000
1!
1%
1-
12
#559720000000
0!
0%
b10 *
0-
02
b10 6
#559730000000
1!
1%
1-
12
#559740000000
0!
0%
b11 *
0-
02
b11 6
#559750000000
1!
1%
1-
12
15
#559760000000
0!
0%
b100 *
0-
02
b100 6
#559770000000
1!
1%
1-
12
#559780000000
0!
0%
b101 *
0-
02
b101 6
#559790000000
1!
1%
1-
12
#559800000000
0!
0%
b110 *
0-
02
b110 6
#559810000000
1!
1%
1-
12
#559820000000
0!
0%
b111 *
0-
02
b111 6
#559830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#559840000000
0!
0%
b0 *
0-
02
b0 6
#559850000000
1!
1%
1-
12
#559860000000
0!
0%
b1 *
0-
02
b1 6
#559870000000
1!
1%
1-
12
#559880000000
0!
0%
b10 *
0-
02
b10 6
#559890000000
1!
1%
1-
12
#559900000000
0!
0%
b11 *
0-
02
b11 6
#559910000000
1!
1%
1-
12
15
#559920000000
0!
0%
b100 *
0-
02
b100 6
#559930000000
1!
1%
1-
12
#559940000000
0!
0%
b101 *
0-
02
b101 6
#559950000000
1!
1%
1-
12
#559960000000
0!
0%
b110 *
0-
02
b110 6
#559970000000
1!
1%
1-
12
#559980000000
0!
0%
b111 *
0-
02
b111 6
#559990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#560000000000
0!
0%
b0 *
0-
02
b0 6
#560010000000
1!
1%
1-
12
#560020000000
0!
0%
b1 *
0-
02
b1 6
#560030000000
1!
1%
1-
12
#560040000000
0!
0%
b10 *
0-
02
b10 6
#560050000000
1!
1%
1-
12
#560060000000
0!
0%
b11 *
0-
02
b11 6
#560070000000
1!
1%
1-
12
15
#560080000000
0!
0%
b100 *
0-
02
b100 6
#560090000000
1!
1%
1-
12
#560100000000
0!
0%
b101 *
0-
02
b101 6
#560110000000
1!
1%
1-
12
#560120000000
0!
0%
b110 *
0-
02
b110 6
#560130000000
1!
1%
1-
12
#560140000000
0!
0%
b111 *
0-
02
b111 6
#560150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#560160000000
0!
0%
b0 *
0-
02
b0 6
#560170000000
1!
1%
1-
12
#560180000000
0!
0%
b1 *
0-
02
b1 6
#560190000000
1!
1%
1-
12
#560200000000
0!
0%
b10 *
0-
02
b10 6
#560210000000
1!
1%
1-
12
#560220000000
0!
0%
b11 *
0-
02
b11 6
#560230000000
1!
1%
1-
12
15
#560240000000
0!
0%
b100 *
0-
02
b100 6
#560250000000
1!
1%
1-
12
#560260000000
0!
0%
b101 *
0-
02
b101 6
#560270000000
1!
1%
1-
12
#560280000000
0!
0%
b110 *
0-
02
b110 6
#560290000000
1!
1%
1-
12
#560300000000
0!
0%
b111 *
0-
02
b111 6
#560310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#560320000000
0!
0%
b0 *
0-
02
b0 6
#560330000000
1!
1%
1-
12
#560340000000
0!
0%
b1 *
0-
02
b1 6
#560350000000
1!
1%
1-
12
#560360000000
0!
0%
b10 *
0-
02
b10 6
#560370000000
1!
1%
1-
12
#560380000000
0!
0%
b11 *
0-
02
b11 6
#560390000000
1!
1%
1-
12
15
#560400000000
0!
0%
b100 *
0-
02
b100 6
#560410000000
1!
1%
1-
12
#560420000000
0!
0%
b101 *
0-
02
b101 6
#560430000000
1!
1%
1-
12
#560440000000
0!
0%
b110 *
0-
02
b110 6
#560450000000
1!
1%
1-
12
#560460000000
0!
0%
b111 *
0-
02
b111 6
#560470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#560480000000
0!
0%
b0 *
0-
02
b0 6
#560490000000
1!
1%
1-
12
#560500000000
0!
0%
b1 *
0-
02
b1 6
#560510000000
1!
1%
1-
12
#560520000000
0!
0%
b10 *
0-
02
b10 6
#560530000000
1!
1%
1-
12
#560540000000
0!
0%
b11 *
0-
02
b11 6
#560550000000
1!
1%
1-
12
15
#560560000000
0!
0%
b100 *
0-
02
b100 6
#560570000000
1!
1%
1-
12
#560580000000
0!
0%
b101 *
0-
02
b101 6
#560590000000
1!
1%
1-
12
#560600000000
0!
0%
b110 *
0-
02
b110 6
#560610000000
1!
1%
1-
12
#560620000000
0!
0%
b111 *
0-
02
b111 6
#560630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#560640000000
0!
0%
b0 *
0-
02
b0 6
#560650000000
1!
1%
1-
12
#560660000000
0!
0%
b1 *
0-
02
b1 6
#560670000000
1!
1%
1-
12
#560680000000
0!
0%
b10 *
0-
02
b10 6
#560690000000
1!
1%
1-
12
#560700000000
0!
0%
b11 *
0-
02
b11 6
#560710000000
1!
1%
1-
12
15
#560720000000
0!
0%
b100 *
0-
02
b100 6
#560730000000
1!
1%
1-
12
#560740000000
0!
0%
b101 *
0-
02
b101 6
#560750000000
1!
1%
1-
12
#560760000000
0!
0%
b110 *
0-
02
b110 6
#560770000000
1!
1%
1-
12
#560780000000
0!
0%
b111 *
0-
02
b111 6
#560790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#560800000000
0!
0%
b0 *
0-
02
b0 6
#560810000000
1!
1%
1-
12
#560820000000
0!
0%
b1 *
0-
02
b1 6
#560830000000
1!
1%
1-
12
#560840000000
0!
0%
b10 *
0-
02
b10 6
#560850000000
1!
1%
1-
12
#560860000000
0!
0%
b11 *
0-
02
b11 6
#560870000000
1!
1%
1-
12
15
#560880000000
0!
0%
b100 *
0-
02
b100 6
#560890000000
1!
1%
1-
12
#560900000000
0!
0%
b101 *
0-
02
b101 6
#560910000000
1!
1%
1-
12
#560920000000
0!
0%
b110 *
0-
02
b110 6
#560930000000
1!
1%
1-
12
#560940000000
0!
0%
b111 *
0-
02
b111 6
#560950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#560960000000
0!
0%
b0 *
0-
02
b0 6
#560970000000
1!
1%
1-
12
#560980000000
0!
0%
b1 *
0-
02
b1 6
#560990000000
1!
1%
1-
12
#561000000000
0!
0%
b10 *
0-
02
b10 6
#561010000000
1!
1%
1-
12
#561020000000
0!
0%
b11 *
0-
02
b11 6
#561030000000
1!
1%
1-
12
15
#561040000000
0!
0%
b100 *
0-
02
b100 6
#561050000000
1!
1%
1-
12
#561060000000
0!
0%
b101 *
0-
02
b101 6
#561070000000
1!
1%
1-
12
#561080000000
0!
0%
b110 *
0-
02
b110 6
#561090000000
1!
1%
1-
12
#561100000000
0!
0%
b111 *
0-
02
b111 6
#561110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#561120000000
0!
0%
b0 *
0-
02
b0 6
#561130000000
1!
1%
1-
12
#561140000000
0!
0%
b1 *
0-
02
b1 6
#561150000000
1!
1%
1-
12
#561160000000
0!
0%
b10 *
0-
02
b10 6
#561170000000
1!
1%
1-
12
#561180000000
0!
0%
b11 *
0-
02
b11 6
#561190000000
1!
1%
1-
12
15
#561200000000
0!
0%
b100 *
0-
02
b100 6
#561210000000
1!
1%
1-
12
#561220000000
0!
0%
b101 *
0-
02
b101 6
#561230000000
1!
1%
1-
12
#561240000000
0!
0%
b110 *
0-
02
b110 6
#561250000000
1!
1%
1-
12
#561260000000
0!
0%
b111 *
0-
02
b111 6
#561270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#561280000000
0!
0%
b0 *
0-
02
b0 6
#561290000000
1!
1%
1-
12
#561300000000
0!
0%
b1 *
0-
02
b1 6
#561310000000
1!
1%
1-
12
#561320000000
0!
0%
b10 *
0-
02
b10 6
#561330000000
1!
1%
1-
12
#561340000000
0!
0%
b11 *
0-
02
b11 6
#561350000000
1!
1%
1-
12
15
#561360000000
0!
0%
b100 *
0-
02
b100 6
#561370000000
1!
1%
1-
12
#561380000000
0!
0%
b101 *
0-
02
b101 6
#561390000000
1!
1%
1-
12
#561400000000
0!
0%
b110 *
0-
02
b110 6
#561410000000
1!
1%
1-
12
#561420000000
0!
0%
b111 *
0-
02
b111 6
#561430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#561440000000
0!
0%
b0 *
0-
02
b0 6
#561450000000
1!
1%
1-
12
#561460000000
0!
0%
b1 *
0-
02
b1 6
#561470000000
1!
1%
1-
12
#561480000000
0!
0%
b10 *
0-
02
b10 6
#561490000000
1!
1%
1-
12
#561500000000
0!
0%
b11 *
0-
02
b11 6
#561510000000
1!
1%
1-
12
15
#561520000000
0!
0%
b100 *
0-
02
b100 6
#561530000000
1!
1%
1-
12
#561540000000
0!
0%
b101 *
0-
02
b101 6
#561550000000
1!
1%
1-
12
#561560000000
0!
0%
b110 *
0-
02
b110 6
#561570000000
1!
1%
1-
12
#561580000000
0!
0%
b111 *
0-
02
b111 6
#561590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#561600000000
0!
0%
b0 *
0-
02
b0 6
#561610000000
1!
1%
1-
12
#561620000000
0!
0%
b1 *
0-
02
b1 6
#561630000000
1!
1%
1-
12
#561640000000
0!
0%
b10 *
0-
02
b10 6
#561650000000
1!
1%
1-
12
#561660000000
0!
0%
b11 *
0-
02
b11 6
#561670000000
1!
1%
1-
12
15
#561680000000
0!
0%
b100 *
0-
02
b100 6
#561690000000
1!
1%
1-
12
#561700000000
0!
0%
b101 *
0-
02
b101 6
#561710000000
1!
1%
1-
12
#561720000000
0!
0%
b110 *
0-
02
b110 6
#561730000000
1!
1%
1-
12
#561740000000
0!
0%
b111 *
0-
02
b111 6
#561750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#561760000000
0!
0%
b0 *
0-
02
b0 6
#561770000000
1!
1%
1-
12
#561780000000
0!
0%
b1 *
0-
02
b1 6
#561790000000
1!
1%
1-
12
#561800000000
0!
0%
b10 *
0-
02
b10 6
#561810000000
1!
1%
1-
12
#561820000000
0!
0%
b11 *
0-
02
b11 6
#561830000000
1!
1%
1-
12
15
#561840000000
0!
0%
b100 *
0-
02
b100 6
#561850000000
1!
1%
1-
12
#561860000000
0!
0%
b101 *
0-
02
b101 6
#561870000000
1!
1%
1-
12
#561880000000
0!
0%
b110 *
0-
02
b110 6
#561890000000
1!
1%
1-
12
#561900000000
0!
0%
b111 *
0-
02
b111 6
#561910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#561920000000
0!
0%
b0 *
0-
02
b0 6
#561930000000
1!
1%
1-
12
#561940000000
0!
0%
b1 *
0-
02
b1 6
#561950000000
1!
1%
1-
12
#561960000000
0!
0%
b10 *
0-
02
b10 6
#561970000000
1!
1%
1-
12
#561980000000
0!
0%
b11 *
0-
02
b11 6
#561990000000
1!
1%
1-
12
15
#562000000000
0!
0%
b100 *
0-
02
b100 6
#562010000000
1!
1%
1-
12
#562020000000
0!
0%
b101 *
0-
02
b101 6
#562030000000
1!
1%
1-
12
#562040000000
0!
0%
b110 *
0-
02
b110 6
#562050000000
1!
1%
1-
12
#562060000000
0!
0%
b111 *
0-
02
b111 6
#562070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#562080000000
0!
0%
b0 *
0-
02
b0 6
#562090000000
1!
1%
1-
12
#562100000000
0!
0%
b1 *
0-
02
b1 6
#562110000000
1!
1%
1-
12
#562120000000
0!
0%
b10 *
0-
02
b10 6
#562130000000
1!
1%
1-
12
#562140000000
0!
0%
b11 *
0-
02
b11 6
#562150000000
1!
1%
1-
12
15
#562160000000
0!
0%
b100 *
0-
02
b100 6
#562170000000
1!
1%
1-
12
#562180000000
0!
0%
b101 *
0-
02
b101 6
#562190000000
1!
1%
1-
12
#562200000000
0!
0%
b110 *
0-
02
b110 6
#562210000000
1!
1%
1-
12
#562220000000
0!
0%
b111 *
0-
02
b111 6
#562230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#562240000000
0!
0%
b0 *
0-
02
b0 6
#562250000000
1!
1%
1-
12
#562260000000
0!
0%
b1 *
0-
02
b1 6
#562270000000
1!
1%
1-
12
#562280000000
0!
0%
b10 *
0-
02
b10 6
#562290000000
1!
1%
1-
12
#562300000000
0!
0%
b11 *
0-
02
b11 6
#562310000000
1!
1%
1-
12
15
#562320000000
0!
0%
b100 *
0-
02
b100 6
#562330000000
1!
1%
1-
12
#562340000000
0!
0%
b101 *
0-
02
b101 6
#562350000000
1!
1%
1-
12
#562360000000
0!
0%
b110 *
0-
02
b110 6
#562370000000
1!
1%
1-
12
#562380000000
0!
0%
b111 *
0-
02
b111 6
#562390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#562400000000
0!
0%
b0 *
0-
02
b0 6
#562410000000
1!
1%
1-
12
#562420000000
0!
0%
b1 *
0-
02
b1 6
#562430000000
1!
1%
1-
12
#562440000000
0!
0%
b10 *
0-
02
b10 6
#562450000000
1!
1%
1-
12
#562460000000
0!
0%
b11 *
0-
02
b11 6
#562470000000
1!
1%
1-
12
15
#562480000000
0!
0%
b100 *
0-
02
b100 6
#562490000000
1!
1%
1-
12
#562500000000
0!
0%
b101 *
0-
02
b101 6
#562510000000
1!
1%
1-
12
#562520000000
0!
0%
b110 *
0-
02
b110 6
#562530000000
1!
1%
1-
12
#562540000000
0!
0%
b111 *
0-
02
b111 6
#562550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#562560000000
0!
0%
b0 *
0-
02
b0 6
#562570000000
1!
1%
1-
12
#562580000000
0!
0%
b1 *
0-
02
b1 6
#562590000000
1!
1%
1-
12
#562600000000
0!
0%
b10 *
0-
02
b10 6
#562610000000
1!
1%
1-
12
#562620000000
0!
0%
b11 *
0-
02
b11 6
#562630000000
1!
1%
1-
12
15
#562640000000
0!
0%
b100 *
0-
02
b100 6
#562650000000
1!
1%
1-
12
#562660000000
0!
0%
b101 *
0-
02
b101 6
#562670000000
1!
1%
1-
12
#562680000000
0!
0%
b110 *
0-
02
b110 6
#562690000000
1!
1%
1-
12
#562700000000
0!
0%
b111 *
0-
02
b111 6
#562710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#562720000000
0!
0%
b0 *
0-
02
b0 6
#562730000000
1!
1%
1-
12
#562740000000
0!
0%
b1 *
0-
02
b1 6
#562750000000
1!
1%
1-
12
#562760000000
0!
0%
b10 *
0-
02
b10 6
#562770000000
1!
1%
1-
12
#562780000000
0!
0%
b11 *
0-
02
b11 6
#562790000000
1!
1%
1-
12
15
#562800000000
0!
0%
b100 *
0-
02
b100 6
#562810000000
1!
1%
1-
12
#562820000000
0!
0%
b101 *
0-
02
b101 6
#562830000000
1!
1%
1-
12
#562840000000
0!
0%
b110 *
0-
02
b110 6
#562850000000
1!
1%
1-
12
#562860000000
0!
0%
b111 *
0-
02
b111 6
#562870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#562880000000
0!
0%
b0 *
0-
02
b0 6
#562890000000
1!
1%
1-
12
#562900000000
0!
0%
b1 *
0-
02
b1 6
#562910000000
1!
1%
1-
12
#562920000000
0!
0%
b10 *
0-
02
b10 6
#562930000000
1!
1%
1-
12
#562940000000
0!
0%
b11 *
0-
02
b11 6
#562950000000
1!
1%
1-
12
15
#562960000000
0!
0%
b100 *
0-
02
b100 6
#562970000000
1!
1%
1-
12
#562980000000
0!
0%
b101 *
0-
02
b101 6
#562990000000
1!
1%
1-
12
#563000000000
0!
0%
b110 *
0-
02
b110 6
#563010000000
1!
1%
1-
12
#563020000000
0!
0%
b111 *
0-
02
b111 6
#563030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#563040000000
0!
0%
b0 *
0-
02
b0 6
#563050000000
1!
1%
1-
12
#563060000000
0!
0%
b1 *
0-
02
b1 6
#563070000000
1!
1%
1-
12
#563080000000
0!
0%
b10 *
0-
02
b10 6
#563090000000
1!
1%
1-
12
#563100000000
0!
0%
b11 *
0-
02
b11 6
#563110000000
1!
1%
1-
12
15
#563120000000
0!
0%
b100 *
0-
02
b100 6
#563130000000
1!
1%
1-
12
#563140000000
0!
0%
b101 *
0-
02
b101 6
#563150000000
1!
1%
1-
12
#563160000000
0!
0%
b110 *
0-
02
b110 6
#563170000000
1!
1%
1-
12
#563180000000
0!
0%
b111 *
0-
02
b111 6
#563190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#563200000000
0!
0%
b0 *
0-
02
b0 6
#563210000000
1!
1%
1-
12
#563220000000
0!
0%
b1 *
0-
02
b1 6
#563230000000
1!
1%
1-
12
#563240000000
0!
0%
b10 *
0-
02
b10 6
#563250000000
1!
1%
1-
12
#563260000000
0!
0%
b11 *
0-
02
b11 6
#563270000000
1!
1%
1-
12
15
#563280000000
0!
0%
b100 *
0-
02
b100 6
#563290000000
1!
1%
1-
12
#563300000000
0!
0%
b101 *
0-
02
b101 6
#563310000000
1!
1%
1-
12
#563320000000
0!
0%
b110 *
0-
02
b110 6
#563330000000
1!
1%
1-
12
#563340000000
0!
0%
b111 *
0-
02
b111 6
#563350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#563360000000
0!
0%
b0 *
0-
02
b0 6
#563370000000
1!
1%
1-
12
#563380000000
0!
0%
b1 *
0-
02
b1 6
#563390000000
1!
1%
1-
12
#563400000000
0!
0%
b10 *
0-
02
b10 6
#563410000000
1!
1%
1-
12
#563420000000
0!
0%
b11 *
0-
02
b11 6
#563430000000
1!
1%
1-
12
15
#563440000000
0!
0%
b100 *
0-
02
b100 6
#563450000000
1!
1%
1-
12
#563460000000
0!
0%
b101 *
0-
02
b101 6
#563470000000
1!
1%
1-
12
#563480000000
0!
0%
b110 *
0-
02
b110 6
#563490000000
1!
1%
1-
12
#563500000000
0!
0%
b111 *
0-
02
b111 6
#563510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#563520000000
0!
0%
b0 *
0-
02
b0 6
#563530000000
1!
1%
1-
12
#563540000000
0!
0%
b1 *
0-
02
b1 6
#563550000000
1!
1%
1-
12
#563560000000
0!
0%
b10 *
0-
02
b10 6
#563570000000
1!
1%
1-
12
#563580000000
0!
0%
b11 *
0-
02
b11 6
#563590000000
1!
1%
1-
12
15
#563600000000
0!
0%
b100 *
0-
02
b100 6
#563610000000
1!
1%
1-
12
#563620000000
0!
0%
b101 *
0-
02
b101 6
#563630000000
1!
1%
1-
12
#563640000000
0!
0%
b110 *
0-
02
b110 6
#563650000000
1!
1%
1-
12
#563660000000
0!
0%
b111 *
0-
02
b111 6
#563670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#563680000000
0!
0%
b0 *
0-
02
b0 6
#563690000000
1!
1%
1-
12
#563700000000
0!
0%
b1 *
0-
02
b1 6
#563710000000
1!
1%
1-
12
#563720000000
0!
0%
b10 *
0-
02
b10 6
#563730000000
1!
1%
1-
12
#563740000000
0!
0%
b11 *
0-
02
b11 6
#563750000000
1!
1%
1-
12
15
#563760000000
0!
0%
b100 *
0-
02
b100 6
#563770000000
1!
1%
1-
12
#563780000000
0!
0%
b101 *
0-
02
b101 6
#563790000000
1!
1%
1-
12
#563800000000
0!
0%
b110 *
0-
02
b110 6
#563810000000
1!
1%
1-
12
#563820000000
0!
0%
b111 *
0-
02
b111 6
#563830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#563840000000
0!
0%
b0 *
0-
02
b0 6
#563850000000
1!
1%
1-
12
#563860000000
0!
0%
b1 *
0-
02
b1 6
#563870000000
1!
1%
1-
12
#563880000000
0!
0%
b10 *
0-
02
b10 6
#563890000000
1!
1%
1-
12
#563900000000
0!
0%
b11 *
0-
02
b11 6
#563910000000
1!
1%
1-
12
15
#563920000000
0!
0%
b100 *
0-
02
b100 6
#563930000000
1!
1%
1-
12
#563940000000
0!
0%
b101 *
0-
02
b101 6
#563950000000
1!
1%
1-
12
#563960000000
0!
0%
b110 *
0-
02
b110 6
#563970000000
1!
1%
1-
12
#563980000000
0!
0%
b111 *
0-
02
b111 6
#563990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#564000000000
0!
0%
b0 *
0-
02
b0 6
#564010000000
1!
1%
1-
12
#564020000000
0!
0%
b1 *
0-
02
b1 6
#564030000000
1!
1%
1-
12
#564040000000
0!
0%
b10 *
0-
02
b10 6
#564050000000
1!
1%
1-
12
#564060000000
0!
0%
b11 *
0-
02
b11 6
#564070000000
1!
1%
1-
12
15
#564080000000
0!
0%
b100 *
0-
02
b100 6
#564090000000
1!
1%
1-
12
#564100000000
0!
0%
b101 *
0-
02
b101 6
#564110000000
1!
1%
1-
12
#564120000000
0!
0%
b110 *
0-
02
b110 6
#564130000000
1!
1%
1-
12
#564140000000
0!
0%
b111 *
0-
02
b111 6
#564150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#564160000000
0!
0%
b0 *
0-
02
b0 6
#564170000000
1!
1%
1-
12
#564180000000
0!
0%
b1 *
0-
02
b1 6
#564190000000
1!
1%
1-
12
#564200000000
0!
0%
b10 *
0-
02
b10 6
#564210000000
1!
1%
1-
12
#564220000000
0!
0%
b11 *
0-
02
b11 6
#564230000000
1!
1%
1-
12
15
#564240000000
0!
0%
b100 *
0-
02
b100 6
#564250000000
1!
1%
1-
12
#564260000000
0!
0%
b101 *
0-
02
b101 6
#564270000000
1!
1%
1-
12
#564280000000
0!
0%
b110 *
0-
02
b110 6
#564290000000
1!
1%
1-
12
#564300000000
0!
0%
b111 *
0-
02
b111 6
#564310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#564320000000
0!
0%
b0 *
0-
02
b0 6
#564330000000
1!
1%
1-
12
#564340000000
0!
0%
b1 *
0-
02
b1 6
#564350000000
1!
1%
1-
12
#564360000000
0!
0%
b10 *
0-
02
b10 6
#564370000000
1!
1%
1-
12
#564380000000
0!
0%
b11 *
0-
02
b11 6
#564390000000
1!
1%
1-
12
15
#564400000000
0!
0%
b100 *
0-
02
b100 6
#564410000000
1!
1%
1-
12
#564420000000
0!
0%
b101 *
0-
02
b101 6
#564430000000
1!
1%
1-
12
#564440000000
0!
0%
b110 *
0-
02
b110 6
#564450000000
1!
1%
1-
12
#564460000000
0!
0%
b111 *
0-
02
b111 6
#564470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#564480000000
0!
0%
b0 *
0-
02
b0 6
#564490000000
1!
1%
1-
12
#564500000000
0!
0%
b1 *
0-
02
b1 6
#564510000000
1!
1%
1-
12
#564520000000
0!
0%
b10 *
0-
02
b10 6
#564530000000
1!
1%
1-
12
#564540000000
0!
0%
b11 *
0-
02
b11 6
#564550000000
1!
1%
1-
12
15
#564560000000
0!
0%
b100 *
0-
02
b100 6
#564570000000
1!
1%
1-
12
#564580000000
0!
0%
b101 *
0-
02
b101 6
#564590000000
1!
1%
1-
12
#564600000000
0!
0%
b110 *
0-
02
b110 6
#564610000000
1!
1%
1-
12
#564620000000
0!
0%
b111 *
0-
02
b111 6
#564630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#564640000000
0!
0%
b0 *
0-
02
b0 6
#564650000000
1!
1%
1-
12
#564660000000
0!
0%
b1 *
0-
02
b1 6
#564670000000
1!
1%
1-
12
#564680000000
0!
0%
b10 *
0-
02
b10 6
#564690000000
1!
1%
1-
12
#564700000000
0!
0%
b11 *
0-
02
b11 6
#564710000000
1!
1%
1-
12
15
#564720000000
0!
0%
b100 *
0-
02
b100 6
#564730000000
1!
1%
1-
12
#564740000000
0!
0%
b101 *
0-
02
b101 6
#564750000000
1!
1%
1-
12
#564760000000
0!
0%
b110 *
0-
02
b110 6
#564770000000
1!
1%
1-
12
#564780000000
0!
0%
b111 *
0-
02
b111 6
#564790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#564800000000
0!
0%
b0 *
0-
02
b0 6
#564810000000
1!
1%
1-
12
#564820000000
0!
0%
b1 *
0-
02
b1 6
#564830000000
1!
1%
1-
12
#564840000000
0!
0%
b10 *
0-
02
b10 6
#564850000000
1!
1%
1-
12
#564860000000
0!
0%
b11 *
0-
02
b11 6
#564870000000
1!
1%
1-
12
15
#564880000000
0!
0%
b100 *
0-
02
b100 6
#564890000000
1!
1%
1-
12
#564900000000
0!
0%
b101 *
0-
02
b101 6
#564910000000
1!
1%
1-
12
#564920000000
0!
0%
b110 *
0-
02
b110 6
#564930000000
1!
1%
1-
12
#564940000000
0!
0%
b111 *
0-
02
b111 6
#564950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#564960000000
0!
0%
b0 *
0-
02
b0 6
#564970000000
1!
1%
1-
12
#564980000000
0!
0%
b1 *
0-
02
b1 6
#564990000000
1!
1%
1-
12
#565000000000
0!
0%
b10 *
0-
02
b10 6
#565010000000
1!
1%
1-
12
#565020000000
0!
0%
b11 *
0-
02
b11 6
#565030000000
1!
1%
1-
12
15
#565040000000
0!
0%
b100 *
0-
02
b100 6
#565050000000
1!
1%
1-
12
#565060000000
0!
0%
b101 *
0-
02
b101 6
#565070000000
1!
1%
1-
12
#565080000000
0!
0%
b110 *
0-
02
b110 6
#565090000000
1!
1%
1-
12
#565100000000
0!
0%
b111 *
0-
02
b111 6
#565110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#565120000000
0!
0%
b0 *
0-
02
b0 6
#565130000000
1!
1%
1-
12
#565140000000
0!
0%
b1 *
0-
02
b1 6
#565150000000
1!
1%
1-
12
#565160000000
0!
0%
b10 *
0-
02
b10 6
#565170000000
1!
1%
1-
12
#565180000000
0!
0%
b11 *
0-
02
b11 6
#565190000000
1!
1%
1-
12
15
#565200000000
0!
0%
b100 *
0-
02
b100 6
#565210000000
1!
1%
1-
12
#565220000000
0!
0%
b101 *
0-
02
b101 6
#565230000000
1!
1%
1-
12
#565240000000
0!
0%
b110 *
0-
02
b110 6
#565250000000
1!
1%
1-
12
#565260000000
0!
0%
b111 *
0-
02
b111 6
#565270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#565280000000
0!
0%
b0 *
0-
02
b0 6
#565290000000
1!
1%
1-
12
#565300000000
0!
0%
b1 *
0-
02
b1 6
#565310000000
1!
1%
1-
12
#565320000000
0!
0%
b10 *
0-
02
b10 6
#565330000000
1!
1%
1-
12
#565340000000
0!
0%
b11 *
0-
02
b11 6
#565350000000
1!
1%
1-
12
15
#565360000000
0!
0%
b100 *
0-
02
b100 6
#565370000000
1!
1%
1-
12
#565380000000
0!
0%
b101 *
0-
02
b101 6
#565390000000
1!
1%
1-
12
#565400000000
0!
0%
b110 *
0-
02
b110 6
#565410000000
1!
1%
1-
12
#565420000000
0!
0%
b111 *
0-
02
b111 6
#565430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#565440000000
0!
0%
b0 *
0-
02
b0 6
#565450000000
1!
1%
1-
12
#565460000000
0!
0%
b1 *
0-
02
b1 6
#565470000000
1!
1%
1-
12
#565480000000
0!
0%
b10 *
0-
02
b10 6
#565490000000
1!
1%
1-
12
#565500000000
0!
0%
b11 *
0-
02
b11 6
#565510000000
1!
1%
1-
12
15
#565520000000
0!
0%
b100 *
0-
02
b100 6
#565530000000
1!
1%
1-
12
#565540000000
0!
0%
b101 *
0-
02
b101 6
#565550000000
1!
1%
1-
12
#565560000000
0!
0%
b110 *
0-
02
b110 6
#565570000000
1!
1%
1-
12
#565580000000
0!
0%
b111 *
0-
02
b111 6
#565590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#565600000000
0!
0%
b0 *
0-
02
b0 6
#565610000000
1!
1%
1-
12
#565620000000
0!
0%
b1 *
0-
02
b1 6
#565630000000
1!
1%
1-
12
#565640000000
0!
0%
b10 *
0-
02
b10 6
#565650000000
1!
1%
1-
12
#565660000000
0!
0%
b11 *
0-
02
b11 6
#565670000000
1!
1%
1-
12
15
#565680000000
0!
0%
b100 *
0-
02
b100 6
#565690000000
1!
1%
1-
12
#565700000000
0!
0%
b101 *
0-
02
b101 6
#565710000000
1!
1%
1-
12
#565720000000
0!
0%
b110 *
0-
02
b110 6
#565730000000
1!
1%
1-
12
#565740000000
0!
0%
b111 *
0-
02
b111 6
#565750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#565760000000
0!
0%
b0 *
0-
02
b0 6
#565770000000
1!
1%
1-
12
#565780000000
0!
0%
b1 *
0-
02
b1 6
#565790000000
1!
1%
1-
12
#565800000000
0!
0%
b10 *
0-
02
b10 6
#565810000000
1!
1%
1-
12
#565820000000
0!
0%
b11 *
0-
02
b11 6
#565830000000
1!
1%
1-
12
15
#565840000000
0!
0%
b100 *
0-
02
b100 6
#565850000000
1!
1%
1-
12
#565860000000
0!
0%
b101 *
0-
02
b101 6
#565870000000
1!
1%
1-
12
#565880000000
0!
0%
b110 *
0-
02
b110 6
#565890000000
1!
1%
1-
12
#565900000000
0!
0%
b111 *
0-
02
b111 6
#565910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#565920000000
0!
0%
b0 *
0-
02
b0 6
#565930000000
1!
1%
1-
12
#565940000000
0!
0%
b1 *
0-
02
b1 6
#565950000000
1!
1%
1-
12
#565960000000
0!
0%
b10 *
0-
02
b10 6
#565970000000
1!
1%
1-
12
#565980000000
0!
0%
b11 *
0-
02
b11 6
#565990000000
1!
1%
1-
12
15
#566000000000
0!
0%
b100 *
0-
02
b100 6
#566010000000
1!
1%
1-
12
#566020000000
0!
0%
b101 *
0-
02
b101 6
#566030000000
1!
1%
1-
12
#566040000000
0!
0%
b110 *
0-
02
b110 6
#566050000000
1!
1%
1-
12
#566060000000
0!
0%
b111 *
0-
02
b111 6
#566070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#566080000000
0!
0%
b0 *
0-
02
b0 6
#566090000000
1!
1%
1-
12
#566100000000
0!
0%
b1 *
0-
02
b1 6
#566110000000
1!
1%
1-
12
#566120000000
0!
0%
b10 *
0-
02
b10 6
#566130000000
1!
1%
1-
12
#566140000000
0!
0%
b11 *
0-
02
b11 6
#566150000000
1!
1%
1-
12
15
#566160000000
0!
0%
b100 *
0-
02
b100 6
#566170000000
1!
1%
1-
12
#566180000000
0!
0%
b101 *
0-
02
b101 6
#566190000000
1!
1%
1-
12
#566200000000
0!
0%
b110 *
0-
02
b110 6
#566210000000
1!
1%
1-
12
#566220000000
0!
0%
b111 *
0-
02
b111 6
#566230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#566240000000
0!
0%
b0 *
0-
02
b0 6
#566250000000
1!
1%
1-
12
#566260000000
0!
0%
b1 *
0-
02
b1 6
#566270000000
1!
1%
1-
12
#566280000000
0!
0%
b10 *
0-
02
b10 6
#566290000000
1!
1%
1-
12
#566300000000
0!
0%
b11 *
0-
02
b11 6
#566310000000
1!
1%
1-
12
15
#566320000000
0!
0%
b100 *
0-
02
b100 6
#566330000000
1!
1%
1-
12
#566340000000
0!
0%
b101 *
0-
02
b101 6
#566350000000
1!
1%
1-
12
#566360000000
0!
0%
b110 *
0-
02
b110 6
#566370000000
1!
1%
1-
12
#566380000000
0!
0%
b111 *
0-
02
b111 6
#566390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#566400000000
0!
0%
b0 *
0-
02
b0 6
#566410000000
1!
1%
1-
12
#566420000000
0!
0%
b1 *
0-
02
b1 6
#566430000000
1!
1%
1-
12
#566440000000
0!
0%
b10 *
0-
02
b10 6
#566450000000
1!
1%
1-
12
#566460000000
0!
0%
b11 *
0-
02
b11 6
#566470000000
1!
1%
1-
12
15
#566480000000
0!
0%
b100 *
0-
02
b100 6
#566490000000
1!
1%
1-
12
#566500000000
0!
0%
b101 *
0-
02
b101 6
#566510000000
1!
1%
1-
12
#566520000000
0!
0%
b110 *
0-
02
b110 6
#566530000000
1!
1%
1-
12
#566540000000
0!
0%
b111 *
0-
02
b111 6
#566550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#566560000000
0!
0%
b0 *
0-
02
b0 6
#566570000000
1!
1%
1-
12
#566580000000
0!
0%
b1 *
0-
02
b1 6
#566590000000
1!
1%
1-
12
#566600000000
0!
0%
b10 *
0-
02
b10 6
#566610000000
1!
1%
1-
12
#566620000000
0!
0%
b11 *
0-
02
b11 6
#566630000000
1!
1%
1-
12
15
#566640000000
0!
0%
b100 *
0-
02
b100 6
#566650000000
1!
1%
1-
12
#566660000000
0!
0%
b101 *
0-
02
b101 6
#566670000000
1!
1%
1-
12
#566680000000
0!
0%
b110 *
0-
02
b110 6
#566690000000
1!
1%
1-
12
#566700000000
0!
0%
b111 *
0-
02
b111 6
#566710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#566720000000
0!
0%
b0 *
0-
02
b0 6
#566730000000
1!
1%
1-
12
#566740000000
0!
0%
b1 *
0-
02
b1 6
#566750000000
1!
1%
1-
12
#566760000000
0!
0%
b10 *
0-
02
b10 6
#566770000000
1!
1%
1-
12
#566780000000
0!
0%
b11 *
0-
02
b11 6
#566790000000
1!
1%
1-
12
15
#566800000000
0!
0%
b100 *
0-
02
b100 6
#566810000000
1!
1%
1-
12
#566820000000
0!
0%
b101 *
0-
02
b101 6
#566830000000
1!
1%
1-
12
#566840000000
0!
0%
b110 *
0-
02
b110 6
#566850000000
1!
1%
1-
12
#566860000000
0!
0%
b111 *
0-
02
b111 6
#566870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#566880000000
0!
0%
b0 *
0-
02
b0 6
#566890000000
1!
1%
1-
12
#566900000000
0!
0%
b1 *
0-
02
b1 6
#566910000000
1!
1%
1-
12
#566920000000
0!
0%
b10 *
0-
02
b10 6
#566930000000
1!
1%
1-
12
#566940000000
0!
0%
b11 *
0-
02
b11 6
#566950000000
1!
1%
1-
12
15
#566960000000
0!
0%
b100 *
0-
02
b100 6
#566970000000
1!
1%
1-
12
#566980000000
0!
0%
b101 *
0-
02
b101 6
#566990000000
1!
1%
1-
12
#567000000000
0!
0%
b110 *
0-
02
b110 6
#567010000000
1!
1%
1-
12
#567020000000
0!
0%
b111 *
0-
02
b111 6
#567030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#567040000000
0!
0%
b0 *
0-
02
b0 6
#567050000000
1!
1%
1-
12
#567060000000
0!
0%
b1 *
0-
02
b1 6
#567070000000
1!
1%
1-
12
#567080000000
0!
0%
b10 *
0-
02
b10 6
#567090000000
1!
1%
1-
12
#567100000000
0!
0%
b11 *
0-
02
b11 6
#567110000000
1!
1%
1-
12
15
#567120000000
0!
0%
b100 *
0-
02
b100 6
#567130000000
1!
1%
1-
12
#567140000000
0!
0%
b101 *
0-
02
b101 6
#567150000000
1!
1%
1-
12
#567160000000
0!
0%
b110 *
0-
02
b110 6
#567170000000
1!
1%
1-
12
#567180000000
0!
0%
b111 *
0-
02
b111 6
#567190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#567200000000
0!
0%
b0 *
0-
02
b0 6
#567210000000
1!
1%
1-
12
#567220000000
0!
0%
b1 *
0-
02
b1 6
#567230000000
1!
1%
1-
12
#567240000000
0!
0%
b10 *
0-
02
b10 6
#567250000000
1!
1%
1-
12
#567260000000
0!
0%
b11 *
0-
02
b11 6
#567270000000
1!
1%
1-
12
15
#567280000000
0!
0%
b100 *
0-
02
b100 6
#567290000000
1!
1%
1-
12
#567300000000
0!
0%
b101 *
0-
02
b101 6
#567310000000
1!
1%
1-
12
#567320000000
0!
0%
b110 *
0-
02
b110 6
#567330000000
1!
1%
1-
12
#567340000000
0!
0%
b111 *
0-
02
b111 6
#567350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#567360000000
0!
0%
b0 *
0-
02
b0 6
#567370000000
1!
1%
1-
12
#567380000000
0!
0%
b1 *
0-
02
b1 6
#567390000000
1!
1%
1-
12
#567400000000
0!
0%
b10 *
0-
02
b10 6
#567410000000
1!
1%
1-
12
#567420000000
0!
0%
b11 *
0-
02
b11 6
#567430000000
1!
1%
1-
12
15
#567440000000
0!
0%
b100 *
0-
02
b100 6
#567450000000
1!
1%
1-
12
#567460000000
0!
0%
b101 *
0-
02
b101 6
#567470000000
1!
1%
1-
12
#567480000000
0!
0%
b110 *
0-
02
b110 6
#567490000000
1!
1%
1-
12
#567500000000
0!
0%
b111 *
0-
02
b111 6
#567510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#567520000000
0!
0%
b0 *
0-
02
b0 6
#567530000000
1!
1%
1-
12
#567540000000
0!
0%
b1 *
0-
02
b1 6
#567550000000
1!
1%
1-
12
#567560000000
0!
0%
b10 *
0-
02
b10 6
#567570000000
1!
1%
1-
12
#567580000000
0!
0%
b11 *
0-
02
b11 6
#567590000000
1!
1%
1-
12
15
#567600000000
0!
0%
b100 *
0-
02
b100 6
#567610000000
1!
1%
1-
12
#567620000000
0!
0%
b101 *
0-
02
b101 6
#567630000000
1!
1%
1-
12
#567640000000
0!
0%
b110 *
0-
02
b110 6
#567650000000
1!
1%
1-
12
#567660000000
0!
0%
b111 *
0-
02
b111 6
#567670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#567680000000
0!
0%
b0 *
0-
02
b0 6
#567690000000
1!
1%
1-
12
#567700000000
0!
0%
b1 *
0-
02
b1 6
#567710000000
1!
1%
1-
12
#567720000000
0!
0%
b10 *
0-
02
b10 6
#567730000000
1!
1%
1-
12
#567740000000
0!
0%
b11 *
0-
02
b11 6
#567750000000
1!
1%
1-
12
15
#567760000000
0!
0%
b100 *
0-
02
b100 6
#567770000000
1!
1%
1-
12
#567780000000
0!
0%
b101 *
0-
02
b101 6
#567790000000
1!
1%
1-
12
#567800000000
0!
0%
b110 *
0-
02
b110 6
#567810000000
1!
1%
1-
12
#567820000000
0!
0%
b111 *
0-
02
b111 6
#567830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#567840000000
0!
0%
b0 *
0-
02
b0 6
#567850000000
1!
1%
1-
12
#567860000000
0!
0%
b1 *
0-
02
b1 6
#567870000000
1!
1%
1-
12
#567880000000
0!
0%
b10 *
0-
02
b10 6
#567890000000
1!
1%
1-
12
#567900000000
0!
0%
b11 *
0-
02
b11 6
#567910000000
1!
1%
1-
12
15
#567920000000
0!
0%
b100 *
0-
02
b100 6
#567930000000
1!
1%
1-
12
#567940000000
0!
0%
b101 *
0-
02
b101 6
#567950000000
1!
1%
1-
12
#567960000000
0!
0%
b110 *
0-
02
b110 6
#567970000000
1!
1%
1-
12
#567980000000
0!
0%
b111 *
0-
02
b111 6
#567990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#568000000000
0!
0%
b0 *
0-
02
b0 6
#568010000000
1!
1%
1-
12
#568020000000
0!
0%
b1 *
0-
02
b1 6
#568030000000
1!
1%
1-
12
#568040000000
0!
0%
b10 *
0-
02
b10 6
#568050000000
1!
1%
1-
12
#568060000000
0!
0%
b11 *
0-
02
b11 6
#568070000000
1!
1%
1-
12
15
#568080000000
0!
0%
b100 *
0-
02
b100 6
#568090000000
1!
1%
1-
12
#568100000000
0!
0%
b101 *
0-
02
b101 6
#568110000000
1!
1%
1-
12
#568120000000
0!
0%
b110 *
0-
02
b110 6
#568130000000
1!
1%
1-
12
#568140000000
0!
0%
b111 *
0-
02
b111 6
#568150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#568160000000
0!
0%
b0 *
0-
02
b0 6
#568170000000
1!
1%
1-
12
#568180000000
0!
0%
b1 *
0-
02
b1 6
#568190000000
1!
1%
1-
12
#568200000000
0!
0%
b10 *
0-
02
b10 6
#568210000000
1!
1%
1-
12
#568220000000
0!
0%
b11 *
0-
02
b11 6
#568230000000
1!
1%
1-
12
15
#568240000000
0!
0%
b100 *
0-
02
b100 6
#568250000000
1!
1%
1-
12
#568260000000
0!
0%
b101 *
0-
02
b101 6
#568270000000
1!
1%
1-
12
#568280000000
0!
0%
b110 *
0-
02
b110 6
#568290000000
1!
1%
1-
12
#568300000000
0!
0%
b111 *
0-
02
b111 6
#568310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#568320000000
0!
0%
b0 *
0-
02
b0 6
#568330000000
1!
1%
1-
12
#568340000000
0!
0%
b1 *
0-
02
b1 6
#568350000000
1!
1%
1-
12
#568360000000
0!
0%
b10 *
0-
02
b10 6
#568370000000
1!
1%
1-
12
#568380000000
0!
0%
b11 *
0-
02
b11 6
#568390000000
1!
1%
1-
12
15
#568400000000
0!
0%
b100 *
0-
02
b100 6
#568410000000
1!
1%
1-
12
#568420000000
0!
0%
b101 *
0-
02
b101 6
#568430000000
1!
1%
1-
12
#568440000000
0!
0%
b110 *
0-
02
b110 6
#568450000000
1!
1%
1-
12
#568460000000
0!
0%
b111 *
0-
02
b111 6
#568470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#568480000000
0!
0%
b0 *
0-
02
b0 6
#568490000000
1!
1%
1-
12
#568500000000
0!
0%
b1 *
0-
02
b1 6
#568510000000
1!
1%
1-
12
#568520000000
0!
0%
b10 *
0-
02
b10 6
#568530000000
1!
1%
1-
12
#568540000000
0!
0%
b11 *
0-
02
b11 6
#568550000000
1!
1%
1-
12
15
#568560000000
0!
0%
b100 *
0-
02
b100 6
#568570000000
1!
1%
1-
12
#568580000000
0!
0%
b101 *
0-
02
b101 6
#568590000000
1!
1%
1-
12
#568600000000
0!
0%
b110 *
0-
02
b110 6
#568610000000
1!
1%
1-
12
#568620000000
0!
0%
b111 *
0-
02
b111 6
#568630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#568640000000
0!
0%
b0 *
0-
02
b0 6
#568650000000
1!
1%
1-
12
#568660000000
0!
0%
b1 *
0-
02
b1 6
#568670000000
1!
1%
1-
12
#568680000000
0!
0%
b10 *
0-
02
b10 6
#568690000000
1!
1%
1-
12
#568700000000
0!
0%
b11 *
0-
02
b11 6
#568710000000
1!
1%
1-
12
15
#568720000000
0!
0%
b100 *
0-
02
b100 6
#568730000000
1!
1%
1-
12
#568740000000
0!
0%
b101 *
0-
02
b101 6
#568750000000
1!
1%
1-
12
#568760000000
0!
0%
b110 *
0-
02
b110 6
#568770000000
1!
1%
1-
12
#568780000000
0!
0%
b111 *
0-
02
b111 6
#568790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#568800000000
0!
0%
b0 *
0-
02
b0 6
#568810000000
1!
1%
1-
12
#568820000000
0!
0%
b1 *
0-
02
b1 6
#568830000000
1!
1%
1-
12
#568840000000
0!
0%
b10 *
0-
02
b10 6
#568850000000
1!
1%
1-
12
#568860000000
0!
0%
b11 *
0-
02
b11 6
#568870000000
1!
1%
1-
12
15
#568880000000
0!
0%
b100 *
0-
02
b100 6
#568890000000
1!
1%
1-
12
#568900000000
0!
0%
b101 *
0-
02
b101 6
#568910000000
1!
1%
1-
12
#568920000000
0!
0%
b110 *
0-
02
b110 6
#568930000000
1!
1%
1-
12
#568940000000
0!
0%
b111 *
0-
02
b111 6
#568950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#568960000000
0!
0%
b0 *
0-
02
b0 6
#568970000000
1!
1%
1-
12
#568980000000
0!
0%
b1 *
0-
02
b1 6
#568990000000
1!
1%
1-
12
#569000000000
0!
0%
b10 *
0-
02
b10 6
#569010000000
1!
1%
1-
12
#569020000000
0!
0%
b11 *
0-
02
b11 6
#569030000000
1!
1%
1-
12
15
#569040000000
0!
0%
b100 *
0-
02
b100 6
#569050000000
1!
1%
1-
12
#569060000000
0!
0%
b101 *
0-
02
b101 6
#569070000000
1!
1%
1-
12
#569080000000
0!
0%
b110 *
0-
02
b110 6
#569090000000
1!
1%
1-
12
#569100000000
0!
0%
b111 *
0-
02
b111 6
#569110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#569120000000
0!
0%
b0 *
0-
02
b0 6
#569130000000
1!
1%
1-
12
#569140000000
0!
0%
b1 *
0-
02
b1 6
#569150000000
1!
1%
1-
12
#569160000000
0!
0%
b10 *
0-
02
b10 6
#569170000000
1!
1%
1-
12
#569180000000
0!
0%
b11 *
0-
02
b11 6
#569190000000
1!
1%
1-
12
15
#569200000000
0!
0%
b100 *
0-
02
b100 6
#569210000000
1!
1%
1-
12
#569220000000
0!
0%
b101 *
0-
02
b101 6
#569230000000
1!
1%
1-
12
#569240000000
0!
0%
b110 *
0-
02
b110 6
#569250000000
1!
1%
1-
12
#569260000000
0!
0%
b111 *
0-
02
b111 6
#569270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#569280000000
0!
0%
b0 *
0-
02
b0 6
#569290000000
1!
1%
1-
12
#569300000000
0!
0%
b1 *
0-
02
b1 6
#569310000000
1!
1%
1-
12
#569320000000
0!
0%
b10 *
0-
02
b10 6
#569330000000
1!
1%
1-
12
#569340000000
0!
0%
b11 *
0-
02
b11 6
#569350000000
1!
1%
1-
12
15
#569360000000
0!
0%
b100 *
0-
02
b100 6
#569370000000
1!
1%
1-
12
#569380000000
0!
0%
b101 *
0-
02
b101 6
#569390000000
1!
1%
1-
12
#569400000000
0!
0%
b110 *
0-
02
b110 6
#569410000000
1!
1%
1-
12
#569420000000
0!
0%
b111 *
0-
02
b111 6
#569430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#569440000000
0!
0%
b0 *
0-
02
b0 6
#569450000000
1!
1%
1-
12
#569460000000
0!
0%
b1 *
0-
02
b1 6
#569470000000
1!
1%
1-
12
#569480000000
0!
0%
b10 *
0-
02
b10 6
#569490000000
1!
1%
1-
12
#569500000000
0!
0%
b11 *
0-
02
b11 6
#569510000000
1!
1%
1-
12
15
#569520000000
0!
0%
b100 *
0-
02
b100 6
#569530000000
1!
1%
1-
12
#569540000000
0!
0%
b101 *
0-
02
b101 6
#569550000000
1!
1%
1-
12
#569560000000
0!
0%
b110 *
0-
02
b110 6
#569570000000
1!
1%
1-
12
#569580000000
0!
0%
b111 *
0-
02
b111 6
#569590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#569600000000
0!
0%
b0 *
0-
02
b0 6
#569610000000
1!
1%
1-
12
#569620000000
0!
0%
b1 *
0-
02
b1 6
#569630000000
1!
1%
1-
12
#569640000000
0!
0%
b10 *
0-
02
b10 6
#569650000000
1!
1%
1-
12
#569660000000
0!
0%
b11 *
0-
02
b11 6
#569670000000
1!
1%
1-
12
15
#569680000000
0!
0%
b100 *
0-
02
b100 6
#569690000000
1!
1%
1-
12
#569700000000
0!
0%
b101 *
0-
02
b101 6
#569710000000
1!
1%
1-
12
#569720000000
0!
0%
b110 *
0-
02
b110 6
#569730000000
1!
1%
1-
12
#569740000000
0!
0%
b111 *
0-
02
b111 6
#569750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#569760000000
0!
0%
b0 *
0-
02
b0 6
#569770000000
1!
1%
1-
12
#569780000000
0!
0%
b1 *
0-
02
b1 6
#569790000000
1!
1%
1-
12
#569800000000
0!
0%
b10 *
0-
02
b10 6
#569810000000
1!
1%
1-
12
#569820000000
0!
0%
b11 *
0-
02
b11 6
#569830000000
1!
1%
1-
12
15
#569840000000
0!
0%
b100 *
0-
02
b100 6
#569850000000
1!
1%
1-
12
#569860000000
0!
0%
b101 *
0-
02
b101 6
#569870000000
1!
1%
1-
12
#569880000000
0!
0%
b110 *
0-
02
b110 6
#569890000000
1!
1%
1-
12
#569900000000
0!
0%
b111 *
0-
02
b111 6
#569910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#569920000000
0!
0%
b0 *
0-
02
b0 6
#569930000000
1!
1%
1-
12
#569940000000
0!
0%
b1 *
0-
02
b1 6
#569950000000
1!
1%
1-
12
#569960000000
0!
0%
b10 *
0-
02
b10 6
#569970000000
1!
1%
1-
12
#569980000000
0!
0%
b11 *
0-
02
b11 6
#569990000000
1!
1%
1-
12
15
#570000000000
0!
0%
b100 *
0-
02
b100 6
#570010000000
1!
1%
1-
12
#570020000000
0!
0%
b101 *
0-
02
b101 6
#570030000000
1!
1%
1-
12
#570040000000
0!
0%
b110 *
0-
02
b110 6
#570050000000
1!
1%
1-
12
#570060000000
0!
0%
b111 *
0-
02
b111 6
#570070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#570080000000
0!
0%
b0 *
0-
02
b0 6
#570090000000
1!
1%
1-
12
#570100000000
0!
0%
b1 *
0-
02
b1 6
#570110000000
1!
1%
1-
12
#570120000000
0!
0%
b10 *
0-
02
b10 6
#570130000000
1!
1%
1-
12
#570140000000
0!
0%
b11 *
0-
02
b11 6
#570150000000
1!
1%
1-
12
15
#570160000000
0!
0%
b100 *
0-
02
b100 6
#570170000000
1!
1%
1-
12
#570180000000
0!
0%
b101 *
0-
02
b101 6
#570190000000
1!
1%
1-
12
#570200000000
0!
0%
b110 *
0-
02
b110 6
#570210000000
1!
1%
1-
12
#570220000000
0!
0%
b111 *
0-
02
b111 6
#570230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#570240000000
0!
0%
b0 *
0-
02
b0 6
#570250000000
1!
1%
1-
12
#570260000000
0!
0%
b1 *
0-
02
b1 6
#570270000000
1!
1%
1-
12
#570280000000
0!
0%
b10 *
0-
02
b10 6
#570290000000
1!
1%
1-
12
#570300000000
0!
0%
b11 *
0-
02
b11 6
#570310000000
1!
1%
1-
12
15
#570320000000
0!
0%
b100 *
0-
02
b100 6
#570330000000
1!
1%
1-
12
#570340000000
0!
0%
b101 *
0-
02
b101 6
#570350000000
1!
1%
1-
12
#570360000000
0!
0%
b110 *
0-
02
b110 6
#570370000000
1!
1%
1-
12
#570380000000
0!
0%
b111 *
0-
02
b111 6
#570390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#570400000000
0!
0%
b0 *
0-
02
b0 6
#570410000000
1!
1%
1-
12
#570420000000
0!
0%
b1 *
0-
02
b1 6
#570430000000
1!
1%
1-
12
#570440000000
0!
0%
b10 *
0-
02
b10 6
#570450000000
1!
1%
1-
12
#570460000000
0!
0%
b11 *
0-
02
b11 6
#570470000000
1!
1%
1-
12
15
#570480000000
0!
0%
b100 *
0-
02
b100 6
#570490000000
1!
1%
1-
12
#570500000000
0!
0%
b101 *
0-
02
b101 6
#570510000000
1!
1%
1-
12
#570520000000
0!
0%
b110 *
0-
02
b110 6
#570530000000
1!
1%
1-
12
#570540000000
0!
0%
b111 *
0-
02
b111 6
#570550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#570560000000
0!
0%
b0 *
0-
02
b0 6
#570570000000
1!
1%
1-
12
#570580000000
0!
0%
b1 *
0-
02
b1 6
#570590000000
1!
1%
1-
12
#570600000000
0!
0%
b10 *
0-
02
b10 6
#570610000000
1!
1%
1-
12
#570620000000
0!
0%
b11 *
0-
02
b11 6
#570630000000
1!
1%
1-
12
15
#570640000000
0!
0%
b100 *
0-
02
b100 6
#570650000000
1!
1%
1-
12
#570660000000
0!
0%
b101 *
0-
02
b101 6
#570670000000
1!
1%
1-
12
#570680000000
0!
0%
b110 *
0-
02
b110 6
#570690000000
1!
1%
1-
12
#570700000000
0!
0%
b111 *
0-
02
b111 6
#570710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#570720000000
0!
0%
b0 *
0-
02
b0 6
#570730000000
1!
1%
1-
12
#570740000000
0!
0%
b1 *
0-
02
b1 6
#570750000000
1!
1%
1-
12
#570760000000
0!
0%
b10 *
0-
02
b10 6
#570770000000
1!
1%
1-
12
#570780000000
0!
0%
b11 *
0-
02
b11 6
#570790000000
1!
1%
1-
12
15
#570800000000
0!
0%
b100 *
0-
02
b100 6
#570810000000
1!
1%
1-
12
#570820000000
0!
0%
b101 *
0-
02
b101 6
#570830000000
1!
1%
1-
12
#570840000000
0!
0%
b110 *
0-
02
b110 6
#570850000000
1!
1%
1-
12
#570860000000
0!
0%
b111 *
0-
02
b111 6
#570870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#570880000000
0!
0%
b0 *
0-
02
b0 6
#570890000000
1!
1%
1-
12
#570900000000
0!
0%
b1 *
0-
02
b1 6
#570910000000
1!
1%
1-
12
#570920000000
0!
0%
b10 *
0-
02
b10 6
#570930000000
1!
1%
1-
12
#570940000000
0!
0%
b11 *
0-
02
b11 6
#570950000000
1!
1%
1-
12
15
#570960000000
0!
0%
b100 *
0-
02
b100 6
#570970000000
1!
1%
1-
12
#570980000000
0!
0%
b101 *
0-
02
b101 6
#570990000000
1!
1%
1-
12
#571000000000
0!
0%
b110 *
0-
02
b110 6
#571010000000
1!
1%
1-
12
#571020000000
0!
0%
b111 *
0-
02
b111 6
#571030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#571040000000
0!
0%
b0 *
0-
02
b0 6
#571050000000
1!
1%
1-
12
#571060000000
0!
0%
b1 *
0-
02
b1 6
#571070000000
1!
1%
1-
12
#571080000000
0!
0%
b10 *
0-
02
b10 6
#571090000000
1!
1%
1-
12
#571100000000
0!
0%
b11 *
0-
02
b11 6
#571110000000
1!
1%
1-
12
15
#571120000000
0!
0%
b100 *
0-
02
b100 6
#571130000000
1!
1%
1-
12
#571140000000
0!
0%
b101 *
0-
02
b101 6
#571150000000
1!
1%
1-
12
#571160000000
0!
0%
b110 *
0-
02
b110 6
#571170000000
1!
1%
1-
12
#571180000000
0!
0%
b111 *
0-
02
b111 6
#571190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#571200000000
0!
0%
b0 *
0-
02
b0 6
#571210000000
1!
1%
1-
12
#571220000000
0!
0%
b1 *
0-
02
b1 6
#571230000000
1!
1%
1-
12
#571240000000
0!
0%
b10 *
0-
02
b10 6
#571250000000
1!
1%
1-
12
#571260000000
0!
0%
b11 *
0-
02
b11 6
#571270000000
1!
1%
1-
12
15
#571280000000
0!
0%
b100 *
0-
02
b100 6
#571290000000
1!
1%
1-
12
#571300000000
0!
0%
b101 *
0-
02
b101 6
#571310000000
1!
1%
1-
12
#571320000000
0!
0%
b110 *
0-
02
b110 6
#571330000000
1!
1%
1-
12
#571340000000
0!
0%
b111 *
0-
02
b111 6
#571350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#571360000000
0!
0%
b0 *
0-
02
b0 6
#571370000000
1!
1%
1-
12
#571380000000
0!
0%
b1 *
0-
02
b1 6
#571390000000
1!
1%
1-
12
#571400000000
0!
0%
b10 *
0-
02
b10 6
#571410000000
1!
1%
1-
12
#571420000000
0!
0%
b11 *
0-
02
b11 6
#571430000000
1!
1%
1-
12
15
#571440000000
0!
0%
b100 *
0-
02
b100 6
#571450000000
1!
1%
1-
12
#571460000000
0!
0%
b101 *
0-
02
b101 6
#571470000000
1!
1%
1-
12
#571480000000
0!
0%
b110 *
0-
02
b110 6
#571490000000
1!
1%
1-
12
#571500000000
0!
0%
b111 *
0-
02
b111 6
#571510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#571520000000
0!
0%
b0 *
0-
02
b0 6
#571530000000
1!
1%
1-
12
#571540000000
0!
0%
b1 *
0-
02
b1 6
#571550000000
1!
1%
1-
12
#571560000000
0!
0%
b10 *
0-
02
b10 6
#571570000000
1!
1%
1-
12
#571580000000
0!
0%
b11 *
0-
02
b11 6
#571590000000
1!
1%
1-
12
15
#571600000000
0!
0%
b100 *
0-
02
b100 6
#571610000000
1!
1%
1-
12
#571620000000
0!
0%
b101 *
0-
02
b101 6
#571630000000
1!
1%
1-
12
#571640000000
0!
0%
b110 *
0-
02
b110 6
#571650000000
1!
1%
1-
12
#571660000000
0!
0%
b111 *
0-
02
b111 6
#571670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#571680000000
0!
0%
b0 *
0-
02
b0 6
#571690000000
1!
1%
1-
12
#571700000000
0!
0%
b1 *
0-
02
b1 6
#571710000000
1!
1%
1-
12
#571720000000
0!
0%
b10 *
0-
02
b10 6
#571730000000
1!
1%
1-
12
#571740000000
0!
0%
b11 *
0-
02
b11 6
#571750000000
1!
1%
1-
12
15
#571760000000
0!
0%
b100 *
0-
02
b100 6
#571770000000
1!
1%
1-
12
#571780000000
0!
0%
b101 *
0-
02
b101 6
#571790000000
1!
1%
1-
12
#571800000000
0!
0%
b110 *
0-
02
b110 6
#571810000000
1!
1%
1-
12
#571820000000
0!
0%
b111 *
0-
02
b111 6
#571830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#571840000000
0!
0%
b0 *
0-
02
b0 6
#571850000000
1!
1%
1-
12
#571860000000
0!
0%
b1 *
0-
02
b1 6
#571870000000
1!
1%
1-
12
#571880000000
0!
0%
b10 *
0-
02
b10 6
#571890000000
1!
1%
1-
12
#571900000000
0!
0%
b11 *
0-
02
b11 6
#571910000000
1!
1%
1-
12
15
#571920000000
0!
0%
b100 *
0-
02
b100 6
#571930000000
1!
1%
1-
12
#571940000000
0!
0%
b101 *
0-
02
b101 6
#571950000000
1!
1%
1-
12
#571960000000
0!
0%
b110 *
0-
02
b110 6
#571970000000
1!
1%
1-
12
#571980000000
0!
0%
b111 *
0-
02
b111 6
#571990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#572000000000
0!
0%
b0 *
0-
02
b0 6
#572010000000
1!
1%
1-
12
#572020000000
0!
0%
b1 *
0-
02
b1 6
#572030000000
1!
1%
1-
12
#572040000000
0!
0%
b10 *
0-
02
b10 6
#572050000000
1!
1%
1-
12
#572060000000
0!
0%
b11 *
0-
02
b11 6
#572070000000
1!
1%
1-
12
15
#572080000000
0!
0%
b100 *
0-
02
b100 6
#572090000000
1!
1%
1-
12
#572100000000
0!
0%
b101 *
0-
02
b101 6
#572110000000
1!
1%
1-
12
#572120000000
0!
0%
b110 *
0-
02
b110 6
#572130000000
1!
1%
1-
12
#572140000000
0!
0%
b111 *
0-
02
b111 6
#572150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#572160000000
0!
0%
b0 *
0-
02
b0 6
#572170000000
1!
1%
1-
12
#572180000000
0!
0%
b1 *
0-
02
b1 6
#572190000000
1!
1%
1-
12
#572200000000
0!
0%
b10 *
0-
02
b10 6
#572210000000
1!
1%
1-
12
#572220000000
0!
0%
b11 *
0-
02
b11 6
#572230000000
1!
1%
1-
12
15
#572240000000
0!
0%
b100 *
0-
02
b100 6
#572250000000
1!
1%
1-
12
#572260000000
0!
0%
b101 *
0-
02
b101 6
#572270000000
1!
1%
1-
12
#572280000000
0!
0%
b110 *
0-
02
b110 6
#572290000000
1!
1%
1-
12
#572300000000
0!
0%
b111 *
0-
02
b111 6
#572310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#572320000000
0!
0%
b0 *
0-
02
b0 6
#572330000000
1!
1%
1-
12
#572340000000
0!
0%
b1 *
0-
02
b1 6
#572350000000
1!
1%
1-
12
#572360000000
0!
0%
b10 *
0-
02
b10 6
#572370000000
1!
1%
1-
12
#572380000000
0!
0%
b11 *
0-
02
b11 6
#572390000000
1!
1%
1-
12
15
#572400000000
0!
0%
b100 *
0-
02
b100 6
#572410000000
1!
1%
1-
12
#572420000000
0!
0%
b101 *
0-
02
b101 6
#572430000000
1!
1%
1-
12
#572440000000
0!
0%
b110 *
0-
02
b110 6
#572450000000
1!
1%
1-
12
#572460000000
0!
0%
b111 *
0-
02
b111 6
#572470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#572480000000
0!
0%
b0 *
0-
02
b0 6
#572490000000
1!
1%
1-
12
#572500000000
0!
0%
b1 *
0-
02
b1 6
#572510000000
1!
1%
1-
12
#572520000000
0!
0%
b10 *
0-
02
b10 6
#572530000000
1!
1%
1-
12
#572540000000
0!
0%
b11 *
0-
02
b11 6
#572550000000
1!
1%
1-
12
15
#572560000000
0!
0%
b100 *
0-
02
b100 6
#572570000000
1!
1%
1-
12
#572580000000
0!
0%
b101 *
0-
02
b101 6
#572590000000
1!
1%
1-
12
#572600000000
0!
0%
b110 *
0-
02
b110 6
#572610000000
1!
1%
1-
12
#572620000000
0!
0%
b111 *
0-
02
b111 6
#572630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#572640000000
0!
0%
b0 *
0-
02
b0 6
#572650000000
1!
1%
1-
12
#572660000000
0!
0%
b1 *
0-
02
b1 6
#572670000000
1!
1%
1-
12
#572680000000
0!
0%
b10 *
0-
02
b10 6
#572690000000
1!
1%
1-
12
#572700000000
0!
0%
b11 *
0-
02
b11 6
#572710000000
1!
1%
1-
12
15
#572720000000
0!
0%
b100 *
0-
02
b100 6
#572730000000
1!
1%
1-
12
#572740000000
0!
0%
b101 *
0-
02
b101 6
#572750000000
1!
1%
1-
12
#572760000000
0!
0%
b110 *
0-
02
b110 6
#572770000000
1!
1%
1-
12
#572780000000
0!
0%
b111 *
0-
02
b111 6
#572790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#572800000000
0!
0%
b0 *
0-
02
b0 6
#572810000000
1!
1%
1-
12
#572820000000
0!
0%
b1 *
0-
02
b1 6
#572830000000
1!
1%
1-
12
#572840000000
0!
0%
b10 *
0-
02
b10 6
#572850000000
1!
1%
1-
12
#572860000000
0!
0%
b11 *
0-
02
b11 6
#572870000000
1!
1%
1-
12
15
#572880000000
0!
0%
b100 *
0-
02
b100 6
#572890000000
1!
1%
1-
12
#572900000000
0!
0%
b101 *
0-
02
b101 6
#572910000000
1!
1%
1-
12
#572920000000
0!
0%
b110 *
0-
02
b110 6
#572930000000
1!
1%
1-
12
#572940000000
0!
0%
b111 *
0-
02
b111 6
#572950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#572960000000
0!
0%
b0 *
0-
02
b0 6
#572970000000
1!
1%
1-
12
#572980000000
0!
0%
b1 *
0-
02
b1 6
#572990000000
1!
1%
1-
12
#573000000000
0!
0%
b10 *
0-
02
b10 6
#573010000000
1!
1%
1-
12
#573020000000
0!
0%
b11 *
0-
02
b11 6
#573030000000
1!
1%
1-
12
15
#573040000000
0!
0%
b100 *
0-
02
b100 6
#573050000000
1!
1%
1-
12
#573060000000
0!
0%
b101 *
0-
02
b101 6
#573070000000
1!
1%
1-
12
#573080000000
0!
0%
b110 *
0-
02
b110 6
#573090000000
1!
1%
1-
12
#573100000000
0!
0%
b111 *
0-
02
b111 6
#573110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#573120000000
0!
0%
b0 *
0-
02
b0 6
#573130000000
1!
1%
1-
12
#573140000000
0!
0%
b1 *
0-
02
b1 6
#573150000000
1!
1%
1-
12
#573160000000
0!
0%
b10 *
0-
02
b10 6
#573170000000
1!
1%
1-
12
#573180000000
0!
0%
b11 *
0-
02
b11 6
#573190000000
1!
1%
1-
12
15
#573200000000
0!
0%
b100 *
0-
02
b100 6
#573210000000
1!
1%
1-
12
#573220000000
0!
0%
b101 *
0-
02
b101 6
#573230000000
1!
1%
1-
12
#573240000000
0!
0%
b110 *
0-
02
b110 6
#573250000000
1!
1%
1-
12
#573260000000
0!
0%
b111 *
0-
02
b111 6
#573270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#573280000000
0!
0%
b0 *
0-
02
b0 6
#573290000000
1!
1%
1-
12
#573300000000
0!
0%
b1 *
0-
02
b1 6
#573310000000
1!
1%
1-
12
#573320000000
0!
0%
b10 *
0-
02
b10 6
#573330000000
1!
1%
1-
12
#573340000000
0!
0%
b11 *
0-
02
b11 6
#573350000000
1!
1%
1-
12
15
#573360000000
0!
0%
b100 *
0-
02
b100 6
#573370000000
1!
1%
1-
12
#573380000000
0!
0%
b101 *
0-
02
b101 6
#573390000000
1!
1%
1-
12
#573400000000
0!
0%
b110 *
0-
02
b110 6
#573410000000
1!
1%
1-
12
#573420000000
0!
0%
b111 *
0-
02
b111 6
#573430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#573440000000
0!
0%
b0 *
0-
02
b0 6
#573450000000
1!
1%
1-
12
#573460000000
0!
0%
b1 *
0-
02
b1 6
#573470000000
1!
1%
1-
12
#573480000000
0!
0%
b10 *
0-
02
b10 6
#573490000000
1!
1%
1-
12
#573500000000
0!
0%
b11 *
0-
02
b11 6
#573510000000
1!
1%
1-
12
15
#573520000000
0!
0%
b100 *
0-
02
b100 6
#573530000000
1!
1%
1-
12
#573540000000
0!
0%
b101 *
0-
02
b101 6
#573550000000
1!
1%
1-
12
#573560000000
0!
0%
b110 *
0-
02
b110 6
#573570000000
1!
1%
1-
12
#573580000000
0!
0%
b111 *
0-
02
b111 6
#573590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#573600000000
0!
0%
b0 *
0-
02
b0 6
#573610000000
1!
1%
1-
12
#573620000000
0!
0%
b1 *
0-
02
b1 6
#573630000000
1!
1%
1-
12
#573640000000
0!
0%
b10 *
0-
02
b10 6
#573650000000
1!
1%
1-
12
#573660000000
0!
0%
b11 *
0-
02
b11 6
#573670000000
1!
1%
1-
12
15
#573680000000
0!
0%
b100 *
0-
02
b100 6
#573690000000
1!
1%
1-
12
#573700000000
0!
0%
b101 *
0-
02
b101 6
#573710000000
1!
1%
1-
12
#573720000000
0!
0%
b110 *
0-
02
b110 6
#573730000000
1!
1%
1-
12
#573740000000
0!
0%
b111 *
0-
02
b111 6
#573750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#573760000000
0!
0%
b0 *
0-
02
b0 6
#573770000000
1!
1%
1-
12
#573780000000
0!
0%
b1 *
0-
02
b1 6
#573790000000
1!
1%
1-
12
#573800000000
0!
0%
b10 *
0-
02
b10 6
#573810000000
1!
1%
1-
12
#573820000000
0!
0%
b11 *
0-
02
b11 6
#573830000000
1!
1%
1-
12
15
#573840000000
0!
0%
b100 *
0-
02
b100 6
#573850000000
1!
1%
1-
12
#573860000000
0!
0%
b101 *
0-
02
b101 6
#573870000000
1!
1%
1-
12
#573880000000
0!
0%
b110 *
0-
02
b110 6
#573890000000
1!
1%
1-
12
#573900000000
0!
0%
b111 *
0-
02
b111 6
#573910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#573920000000
0!
0%
b0 *
0-
02
b0 6
#573930000000
1!
1%
1-
12
#573940000000
0!
0%
b1 *
0-
02
b1 6
#573950000000
1!
1%
1-
12
#573960000000
0!
0%
b10 *
0-
02
b10 6
#573970000000
1!
1%
1-
12
#573980000000
0!
0%
b11 *
0-
02
b11 6
#573990000000
1!
1%
1-
12
15
#574000000000
0!
0%
b100 *
0-
02
b100 6
#574010000000
1!
1%
1-
12
#574020000000
0!
0%
b101 *
0-
02
b101 6
#574030000000
1!
1%
1-
12
#574040000000
0!
0%
b110 *
0-
02
b110 6
#574050000000
1!
1%
1-
12
#574060000000
0!
0%
b111 *
0-
02
b111 6
#574070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#574080000000
0!
0%
b0 *
0-
02
b0 6
#574090000000
1!
1%
1-
12
#574100000000
0!
0%
b1 *
0-
02
b1 6
#574110000000
1!
1%
1-
12
#574120000000
0!
0%
b10 *
0-
02
b10 6
#574130000000
1!
1%
1-
12
#574140000000
0!
0%
b11 *
0-
02
b11 6
#574150000000
1!
1%
1-
12
15
#574160000000
0!
0%
b100 *
0-
02
b100 6
#574170000000
1!
1%
1-
12
#574180000000
0!
0%
b101 *
0-
02
b101 6
#574190000000
1!
1%
1-
12
#574200000000
0!
0%
b110 *
0-
02
b110 6
#574210000000
1!
1%
1-
12
#574220000000
0!
0%
b111 *
0-
02
b111 6
#574230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#574240000000
0!
0%
b0 *
0-
02
b0 6
#574250000000
1!
1%
1-
12
#574260000000
0!
0%
b1 *
0-
02
b1 6
#574270000000
1!
1%
1-
12
#574280000000
0!
0%
b10 *
0-
02
b10 6
#574290000000
1!
1%
1-
12
#574300000000
0!
0%
b11 *
0-
02
b11 6
#574310000000
1!
1%
1-
12
15
#574320000000
0!
0%
b100 *
0-
02
b100 6
#574330000000
1!
1%
1-
12
#574340000000
0!
0%
b101 *
0-
02
b101 6
#574350000000
1!
1%
1-
12
#574360000000
0!
0%
b110 *
0-
02
b110 6
#574370000000
1!
1%
1-
12
#574380000000
0!
0%
b111 *
0-
02
b111 6
#574390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#574400000000
0!
0%
b0 *
0-
02
b0 6
#574410000000
1!
1%
1-
12
#574420000000
0!
0%
b1 *
0-
02
b1 6
#574430000000
1!
1%
1-
12
#574440000000
0!
0%
b10 *
0-
02
b10 6
#574450000000
1!
1%
1-
12
#574460000000
0!
0%
b11 *
0-
02
b11 6
#574470000000
1!
1%
1-
12
15
#574480000000
0!
0%
b100 *
0-
02
b100 6
#574490000000
1!
1%
1-
12
#574500000000
0!
0%
b101 *
0-
02
b101 6
#574510000000
1!
1%
1-
12
#574520000000
0!
0%
b110 *
0-
02
b110 6
#574530000000
1!
1%
1-
12
#574540000000
0!
0%
b111 *
0-
02
b111 6
#574550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#574560000000
0!
0%
b0 *
0-
02
b0 6
#574570000000
1!
1%
1-
12
#574580000000
0!
0%
b1 *
0-
02
b1 6
#574590000000
1!
1%
1-
12
#574600000000
0!
0%
b10 *
0-
02
b10 6
#574610000000
1!
1%
1-
12
#574620000000
0!
0%
b11 *
0-
02
b11 6
#574630000000
1!
1%
1-
12
15
#574640000000
0!
0%
b100 *
0-
02
b100 6
#574650000000
1!
1%
1-
12
#574660000000
0!
0%
b101 *
0-
02
b101 6
#574670000000
1!
1%
1-
12
#574680000000
0!
0%
b110 *
0-
02
b110 6
#574690000000
1!
1%
1-
12
#574700000000
0!
0%
b111 *
0-
02
b111 6
#574710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#574720000000
0!
0%
b0 *
0-
02
b0 6
#574730000000
1!
1%
1-
12
#574740000000
0!
0%
b1 *
0-
02
b1 6
#574750000000
1!
1%
1-
12
#574760000000
0!
0%
b10 *
0-
02
b10 6
#574770000000
1!
1%
1-
12
#574780000000
0!
0%
b11 *
0-
02
b11 6
#574790000000
1!
1%
1-
12
15
#574800000000
0!
0%
b100 *
0-
02
b100 6
#574810000000
1!
1%
1-
12
#574820000000
0!
0%
b101 *
0-
02
b101 6
#574830000000
1!
1%
1-
12
#574840000000
0!
0%
b110 *
0-
02
b110 6
#574850000000
1!
1%
1-
12
#574860000000
0!
0%
b111 *
0-
02
b111 6
#574870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#574880000000
0!
0%
b0 *
0-
02
b0 6
#574890000000
1!
1%
1-
12
#574900000000
0!
0%
b1 *
0-
02
b1 6
#574910000000
1!
1%
1-
12
#574920000000
0!
0%
b10 *
0-
02
b10 6
#574930000000
1!
1%
1-
12
#574940000000
0!
0%
b11 *
0-
02
b11 6
#574950000000
1!
1%
1-
12
15
#574960000000
0!
0%
b100 *
0-
02
b100 6
#574970000000
1!
1%
1-
12
#574980000000
0!
0%
b101 *
0-
02
b101 6
#574990000000
1!
1%
1-
12
#575000000000
0!
0%
b110 *
0-
02
b110 6
#575010000000
1!
1%
1-
12
#575020000000
0!
0%
b111 *
0-
02
b111 6
#575030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#575040000000
0!
0%
b0 *
0-
02
b0 6
#575050000000
1!
1%
1-
12
#575060000000
0!
0%
b1 *
0-
02
b1 6
#575070000000
1!
1%
1-
12
#575080000000
0!
0%
b10 *
0-
02
b10 6
#575090000000
1!
1%
1-
12
#575100000000
0!
0%
b11 *
0-
02
b11 6
#575110000000
1!
1%
1-
12
15
#575120000000
0!
0%
b100 *
0-
02
b100 6
#575130000000
1!
1%
1-
12
#575140000000
0!
0%
b101 *
0-
02
b101 6
#575150000000
1!
1%
1-
12
#575160000000
0!
0%
b110 *
0-
02
b110 6
#575170000000
1!
1%
1-
12
#575180000000
0!
0%
b111 *
0-
02
b111 6
#575190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#575200000000
0!
0%
b0 *
0-
02
b0 6
#575210000000
1!
1%
1-
12
#575220000000
0!
0%
b1 *
0-
02
b1 6
#575230000000
1!
1%
1-
12
#575240000000
0!
0%
b10 *
0-
02
b10 6
#575250000000
1!
1%
1-
12
#575260000000
0!
0%
b11 *
0-
02
b11 6
#575270000000
1!
1%
1-
12
15
#575280000000
0!
0%
b100 *
0-
02
b100 6
#575290000000
1!
1%
1-
12
#575300000000
0!
0%
b101 *
0-
02
b101 6
#575310000000
1!
1%
1-
12
#575320000000
0!
0%
b110 *
0-
02
b110 6
#575330000000
1!
1%
1-
12
#575340000000
0!
0%
b111 *
0-
02
b111 6
#575350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#575360000000
0!
0%
b0 *
0-
02
b0 6
#575370000000
1!
1%
1-
12
#575380000000
0!
0%
b1 *
0-
02
b1 6
#575390000000
1!
1%
1-
12
#575400000000
0!
0%
b10 *
0-
02
b10 6
#575410000000
1!
1%
1-
12
#575420000000
0!
0%
b11 *
0-
02
b11 6
#575430000000
1!
1%
1-
12
15
#575440000000
0!
0%
b100 *
0-
02
b100 6
#575450000000
1!
1%
1-
12
#575460000000
0!
0%
b101 *
0-
02
b101 6
#575470000000
1!
1%
1-
12
#575480000000
0!
0%
b110 *
0-
02
b110 6
#575490000000
1!
1%
1-
12
#575500000000
0!
0%
b111 *
0-
02
b111 6
#575510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#575520000000
0!
0%
b0 *
0-
02
b0 6
#575530000000
1!
1%
1-
12
#575540000000
0!
0%
b1 *
0-
02
b1 6
#575550000000
1!
1%
1-
12
#575560000000
0!
0%
b10 *
0-
02
b10 6
#575570000000
1!
1%
1-
12
#575580000000
0!
0%
b11 *
0-
02
b11 6
#575590000000
1!
1%
1-
12
15
#575600000000
0!
0%
b100 *
0-
02
b100 6
#575610000000
1!
1%
1-
12
#575620000000
0!
0%
b101 *
0-
02
b101 6
#575630000000
1!
1%
1-
12
#575640000000
0!
0%
b110 *
0-
02
b110 6
#575650000000
1!
1%
1-
12
#575660000000
0!
0%
b111 *
0-
02
b111 6
#575670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#575680000000
0!
0%
b0 *
0-
02
b0 6
#575690000000
1!
1%
1-
12
#575700000000
0!
0%
b1 *
0-
02
b1 6
#575710000000
1!
1%
1-
12
#575720000000
0!
0%
b10 *
0-
02
b10 6
#575730000000
1!
1%
1-
12
#575740000000
0!
0%
b11 *
0-
02
b11 6
#575750000000
1!
1%
1-
12
15
#575760000000
0!
0%
b100 *
0-
02
b100 6
#575770000000
1!
1%
1-
12
#575780000000
0!
0%
b101 *
0-
02
b101 6
#575790000000
1!
1%
1-
12
#575800000000
0!
0%
b110 *
0-
02
b110 6
#575810000000
1!
1%
1-
12
#575820000000
0!
0%
b111 *
0-
02
b111 6
#575830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#575840000000
0!
0%
b0 *
0-
02
b0 6
#575850000000
1!
1%
1-
12
#575860000000
0!
0%
b1 *
0-
02
b1 6
#575870000000
1!
1%
1-
12
#575880000000
0!
0%
b10 *
0-
02
b10 6
#575890000000
1!
1%
1-
12
#575900000000
0!
0%
b11 *
0-
02
b11 6
#575910000000
1!
1%
1-
12
15
#575920000000
0!
0%
b100 *
0-
02
b100 6
#575930000000
1!
1%
1-
12
#575940000000
0!
0%
b101 *
0-
02
b101 6
#575950000000
1!
1%
1-
12
#575960000000
0!
0%
b110 *
0-
02
b110 6
#575970000000
1!
1%
1-
12
#575980000000
0!
0%
b111 *
0-
02
b111 6
#575990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#576000000000
0!
0%
b0 *
0-
02
b0 6
#576010000000
1!
1%
1-
12
#576020000000
0!
0%
b1 *
0-
02
b1 6
#576030000000
1!
1%
1-
12
#576040000000
0!
0%
b10 *
0-
02
b10 6
#576050000000
1!
1%
1-
12
#576060000000
0!
0%
b11 *
0-
02
b11 6
#576070000000
1!
1%
1-
12
15
#576080000000
0!
0%
b100 *
0-
02
b100 6
#576090000000
1!
1%
1-
12
#576100000000
0!
0%
b101 *
0-
02
b101 6
#576110000000
1!
1%
1-
12
#576120000000
0!
0%
b110 *
0-
02
b110 6
#576130000000
1!
1%
1-
12
#576140000000
0!
0%
b111 *
0-
02
b111 6
#576150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#576160000000
0!
0%
b0 *
0-
02
b0 6
#576170000000
1!
1%
1-
12
#576180000000
0!
0%
b1 *
0-
02
b1 6
#576190000000
1!
1%
1-
12
#576200000000
0!
0%
b10 *
0-
02
b10 6
#576210000000
1!
1%
1-
12
#576220000000
0!
0%
b11 *
0-
02
b11 6
#576230000000
1!
1%
1-
12
15
#576240000000
0!
0%
b100 *
0-
02
b100 6
#576250000000
1!
1%
1-
12
#576260000000
0!
0%
b101 *
0-
02
b101 6
#576270000000
1!
1%
1-
12
#576280000000
0!
0%
b110 *
0-
02
b110 6
#576290000000
1!
1%
1-
12
#576300000000
0!
0%
b111 *
0-
02
b111 6
#576310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#576320000000
0!
0%
b0 *
0-
02
b0 6
#576330000000
1!
1%
1-
12
#576340000000
0!
0%
b1 *
0-
02
b1 6
#576350000000
1!
1%
1-
12
#576360000000
0!
0%
b10 *
0-
02
b10 6
#576370000000
1!
1%
1-
12
#576380000000
0!
0%
b11 *
0-
02
b11 6
#576390000000
1!
1%
1-
12
15
#576400000000
0!
0%
b100 *
0-
02
b100 6
#576410000000
1!
1%
1-
12
#576420000000
0!
0%
b101 *
0-
02
b101 6
#576430000000
1!
1%
1-
12
#576440000000
0!
0%
b110 *
0-
02
b110 6
#576450000000
1!
1%
1-
12
#576460000000
0!
0%
b111 *
0-
02
b111 6
#576470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#576480000000
0!
0%
b0 *
0-
02
b0 6
#576490000000
1!
1%
1-
12
#576500000000
0!
0%
b1 *
0-
02
b1 6
#576510000000
1!
1%
1-
12
#576520000000
0!
0%
b10 *
0-
02
b10 6
#576530000000
1!
1%
1-
12
#576540000000
0!
0%
b11 *
0-
02
b11 6
#576550000000
1!
1%
1-
12
15
#576560000000
0!
0%
b100 *
0-
02
b100 6
#576570000000
1!
1%
1-
12
#576580000000
0!
0%
b101 *
0-
02
b101 6
#576590000000
1!
1%
1-
12
#576600000000
0!
0%
b110 *
0-
02
b110 6
#576610000000
1!
1%
1-
12
#576620000000
0!
0%
b111 *
0-
02
b111 6
#576630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#576640000000
0!
0%
b0 *
0-
02
b0 6
#576650000000
1!
1%
1-
12
#576660000000
0!
0%
b1 *
0-
02
b1 6
#576670000000
1!
1%
1-
12
#576680000000
0!
0%
b10 *
0-
02
b10 6
#576690000000
1!
1%
1-
12
#576700000000
0!
0%
b11 *
0-
02
b11 6
#576710000000
1!
1%
1-
12
15
#576720000000
0!
0%
b100 *
0-
02
b100 6
#576730000000
1!
1%
1-
12
#576740000000
0!
0%
b101 *
0-
02
b101 6
#576750000000
1!
1%
1-
12
#576760000000
0!
0%
b110 *
0-
02
b110 6
#576770000000
1!
1%
1-
12
#576780000000
0!
0%
b111 *
0-
02
b111 6
#576790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#576800000000
0!
0%
b0 *
0-
02
b0 6
#576810000000
1!
1%
1-
12
#576820000000
0!
0%
b1 *
0-
02
b1 6
#576830000000
1!
1%
1-
12
#576840000000
0!
0%
b10 *
0-
02
b10 6
#576850000000
1!
1%
1-
12
#576860000000
0!
0%
b11 *
0-
02
b11 6
#576870000000
1!
1%
1-
12
15
#576880000000
0!
0%
b100 *
0-
02
b100 6
#576890000000
1!
1%
1-
12
#576900000000
0!
0%
b101 *
0-
02
b101 6
#576910000000
1!
1%
1-
12
#576920000000
0!
0%
b110 *
0-
02
b110 6
#576930000000
1!
1%
1-
12
#576940000000
0!
0%
b111 *
0-
02
b111 6
#576950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#576960000000
0!
0%
b0 *
0-
02
b0 6
#576970000000
1!
1%
1-
12
#576980000000
0!
0%
b1 *
0-
02
b1 6
#576990000000
1!
1%
1-
12
#577000000000
0!
0%
b10 *
0-
02
b10 6
#577010000000
1!
1%
1-
12
#577020000000
0!
0%
b11 *
0-
02
b11 6
#577030000000
1!
1%
1-
12
15
#577040000000
0!
0%
b100 *
0-
02
b100 6
#577050000000
1!
1%
1-
12
#577060000000
0!
0%
b101 *
0-
02
b101 6
#577070000000
1!
1%
1-
12
#577080000000
0!
0%
b110 *
0-
02
b110 6
#577090000000
1!
1%
1-
12
#577100000000
0!
0%
b111 *
0-
02
b111 6
#577110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#577120000000
0!
0%
b0 *
0-
02
b0 6
#577130000000
1!
1%
1-
12
#577140000000
0!
0%
b1 *
0-
02
b1 6
#577150000000
1!
1%
1-
12
#577160000000
0!
0%
b10 *
0-
02
b10 6
#577170000000
1!
1%
1-
12
#577180000000
0!
0%
b11 *
0-
02
b11 6
#577190000000
1!
1%
1-
12
15
#577200000000
0!
0%
b100 *
0-
02
b100 6
#577210000000
1!
1%
1-
12
#577220000000
0!
0%
b101 *
0-
02
b101 6
#577230000000
1!
1%
1-
12
#577240000000
0!
0%
b110 *
0-
02
b110 6
#577250000000
1!
1%
1-
12
#577260000000
0!
0%
b111 *
0-
02
b111 6
#577270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#577280000000
0!
0%
b0 *
0-
02
b0 6
#577290000000
1!
1%
1-
12
#577300000000
0!
0%
b1 *
0-
02
b1 6
#577310000000
1!
1%
1-
12
#577320000000
0!
0%
b10 *
0-
02
b10 6
#577330000000
1!
1%
1-
12
#577340000000
0!
0%
b11 *
0-
02
b11 6
#577350000000
1!
1%
1-
12
15
#577360000000
0!
0%
b100 *
0-
02
b100 6
#577370000000
1!
1%
1-
12
#577380000000
0!
0%
b101 *
0-
02
b101 6
#577390000000
1!
1%
1-
12
#577400000000
0!
0%
b110 *
0-
02
b110 6
#577410000000
1!
1%
1-
12
#577420000000
0!
0%
b111 *
0-
02
b111 6
#577430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#577440000000
0!
0%
b0 *
0-
02
b0 6
#577450000000
1!
1%
1-
12
#577460000000
0!
0%
b1 *
0-
02
b1 6
#577470000000
1!
1%
1-
12
#577480000000
0!
0%
b10 *
0-
02
b10 6
#577490000000
1!
1%
1-
12
#577500000000
0!
0%
b11 *
0-
02
b11 6
#577510000000
1!
1%
1-
12
15
#577520000000
0!
0%
b100 *
0-
02
b100 6
#577530000000
1!
1%
1-
12
#577540000000
0!
0%
b101 *
0-
02
b101 6
#577550000000
1!
1%
1-
12
#577560000000
0!
0%
b110 *
0-
02
b110 6
#577570000000
1!
1%
1-
12
#577580000000
0!
0%
b111 *
0-
02
b111 6
#577590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#577600000000
0!
0%
b0 *
0-
02
b0 6
#577610000000
1!
1%
1-
12
#577620000000
0!
0%
b1 *
0-
02
b1 6
#577630000000
1!
1%
1-
12
#577640000000
0!
0%
b10 *
0-
02
b10 6
#577650000000
1!
1%
1-
12
#577660000000
0!
0%
b11 *
0-
02
b11 6
#577670000000
1!
1%
1-
12
15
#577680000000
0!
0%
b100 *
0-
02
b100 6
#577690000000
1!
1%
1-
12
#577700000000
0!
0%
b101 *
0-
02
b101 6
#577710000000
1!
1%
1-
12
#577720000000
0!
0%
b110 *
0-
02
b110 6
#577730000000
1!
1%
1-
12
#577740000000
0!
0%
b111 *
0-
02
b111 6
#577750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#577760000000
0!
0%
b0 *
0-
02
b0 6
#577770000000
1!
1%
1-
12
#577780000000
0!
0%
b1 *
0-
02
b1 6
#577790000000
1!
1%
1-
12
#577800000000
0!
0%
b10 *
0-
02
b10 6
#577810000000
1!
1%
1-
12
#577820000000
0!
0%
b11 *
0-
02
b11 6
#577830000000
1!
1%
1-
12
15
#577840000000
0!
0%
b100 *
0-
02
b100 6
#577850000000
1!
1%
1-
12
#577860000000
0!
0%
b101 *
0-
02
b101 6
#577870000000
1!
1%
1-
12
#577880000000
0!
0%
b110 *
0-
02
b110 6
#577890000000
1!
1%
1-
12
#577900000000
0!
0%
b111 *
0-
02
b111 6
#577910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#577920000000
0!
0%
b0 *
0-
02
b0 6
#577930000000
1!
1%
1-
12
#577940000000
0!
0%
b1 *
0-
02
b1 6
#577950000000
1!
1%
1-
12
#577960000000
0!
0%
b10 *
0-
02
b10 6
#577970000000
1!
1%
1-
12
#577980000000
0!
0%
b11 *
0-
02
b11 6
#577990000000
1!
1%
1-
12
15
#578000000000
0!
0%
b100 *
0-
02
b100 6
#578010000000
1!
1%
1-
12
#578020000000
0!
0%
b101 *
0-
02
b101 6
#578030000000
1!
1%
1-
12
#578040000000
0!
0%
b110 *
0-
02
b110 6
#578050000000
1!
1%
1-
12
#578060000000
0!
0%
b111 *
0-
02
b111 6
#578070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#578080000000
0!
0%
b0 *
0-
02
b0 6
#578090000000
1!
1%
1-
12
#578100000000
0!
0%
b1 *
0-
02
b1 6
#578110000000
1!
1%
1-
12
#578120000000
0!
0%
b10 *
0-
02
b10 6
#578130000000
1!
1%
1-
12
#578140000000
0!
0%
b11 *
0-
02
b11 6
#578150000000
1!
1%
1-
12
15
#578160000000
0!
0%
b100 *
0-
02
b100 6
#578170000000
1!
1%
1-
12
#578180000000
0!
0%
b101 *
0-
02
b101 6
#578190000000
1!
1%
1-
12
#578200000000
0!
0%
b110 *
0-
02
b110 6
#578210000000
1!
1%
1-
12
#578220000000
0!
0%
b111 *
0-
02
b111 6
#578230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#578240000000
0!
0%
b0 *
0-
02
b0 6
#578250000000
1!
1%
1-
12
#578260000000
0!
0%
b1 *
0-
02
b1 6
#578270000000
1!
1%
1-
12
#578280000000
0!
0%
b10 *
0-
02
b10 6
#578290000000
1!
1%
1-
12
#578300000000
0!
0%
b11 *
0-
02
b11 6
#578310000000
1!
1%
1-
12
15
#578320000000
0!
0%
b100 *
0-
02
b100 6
#578330000000
1!
1%
1-
12
#578340000000
0!
0%
b101 *
0-
02
b101 6
#578350000000
1!
1%
1-
12
#578360000000
0!
0%
b110 *
0-
02
b110 6
#578370000000
1!
1%
1-
12
#578380000000
0!
0%
b111 *
0-
02
b111 6
#578390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#578400000000
0!
0%
b0 *
0-
02
b0 6
#578410000000
1!
1%
1-
12
#578420000000
0!
0%
b1 *
0-
02
b1 6
#578430000000
1!
1%
1-
12
#578440000000
0!
0%
b10 *
0-
02
b10 6
#578450000000
1!
1%
1-
12
#578460000000
0!
0%
b11 *
0-
02
b11 6
#578470000000
1!
1%
1-
12
15
#578480000000
0!
0%
b100 *
0-
02
b100 6
#578490000000
1!
1%
1-
12
#578500000000
0!
0%
b101 *
0-
02
b101 6
#578510000000
1!
1%
1-
12
#578520000000
0!
0%
b110 *
0-
02
b110 6
#578530000000
1!
1%
1-
12
#578540000000
0!
0%
b111 *
0-
02
b111 6
#578550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#578560000000
0!
0%
b0 *
0-
02
b0 6
#578570000000
1!
1%
1-
12
#578580000000
0!
0%
b1 *
0-
02
b1 6
#578590000000
1!
1%
1-
12
#578600000000
0!
0%
b10 *
0-
02
b10 6
#578610000000
1!
1%
1-
12
#578620000000
0!
0%
b11 *
0-
02
b11 6
#578630000000
1!
1%
1-
12
15
#578640000000
0!
0%
b100 *
0-
02
b100 6
#578650000000
1!
1%
1-
12
#578660000000
0!
0%
b101 *
0-
02
b101 6
#578670000000
1!
1%
1-
12
#578680000000
0!
0%
b110 *
0-
02
b110 6
#578690000000
1!
1%
1-
12
#578700000000
0!
0%
b111 *
0-
02
b111 6
#578710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#578720000000
0!
0%
b0 *
0-
02
b0 6
#578730000000
1!
1%
1-
12
#578740000000
0!
0%
b1 *
0-
02
b1 6
#578750000000
1!
1%
1-
12
#578760000000
0!
0%
b10 *
0-
02
b10 6
#578770000000
1!
1%
1-
12
#578780000000
0!
0%
b11 *
0-
02
b11 6
#578790000000
1!
1%
1-
12
15
#578800000000
0!
0%
b100 *
0-
02
b100 6
#578810000000
1!
1%
1-
12
#578820000000
0!
0%
b101 *
0-
02
b101 6
#578830000000
1!
1%
1-
12
#578840000000
0!
0%
b110 *
0-
02
b110 6
#578850000000
1!
1%
1-
12
#578860000000
0!
0%
b111 *
0-
02
b111 6
#578870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#578880000000
0!
0%
b0 *
0-
02
b0 6
#578890000000
1!
1%
1-
12
#578900000000
0!
0%
b1 *
0-
02
b1 6
#578910000000
1!
1%
1-
12
#578920000000
0!
0%
b10 *
0-
02
b10 6
#578930000000
1!
1%
1-
12
#578940000000
0!
0%
b11 *
0-
02
b11 6
#578950000000
1!
1%
1-
12
15
#578960000000
0!
0%
b100 *
0-
02
b100 6
#578970000000
1!
1%
1-
12
#578980000000
0!
0%
b101 *
0-
02
b101 6
#578990000000
1!
1%
1-
12
#579000000000
0!
0%
b110 *
0-
02
b110 6
#579010000000
1!
1%
1-
12
#579020000000
0!
0%
b111 *
0-
02
b111 6
#579030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#579040000000
0!
0%
b0 *
0-
02
b0 6
#579050000000
1!
1%
1-
12
#579060000000
0!
0%
b1 *
0-
02
b1 6
#579070000000
1!
1%
1-
12
#579080000000
0!
0%
b10 *
0-
02
b10 6
#579090000000
1!
1%
1-
12
#579100000000
0!
0%
b11 *
0-
02
b11 6
#579110000000
1!
1%
1-
12
15
#579120000000
0!
0%
b100 *
0-
02
b100 6
#579130000000
1!
1%
1-
12
#579140000000
0!
0%
b101 *
0-
02
b101 6
#579150000000
1!
1%
1-
12
#579160000000
0!
0%
b110 *
0-
02
b110 6
#579170000000
1!
1%
1-
12
#579180000000
0!
0%
b111 *
0-
02
b111 6
#579190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#579200000000
0!
0%
b0 *
0-
02
b0 6
#579210000000
1!
1%
1-
12
#579220000000
0!
0%
b1 *
0-
02
b1 6
#579230000000
1!
1%
1-
12
#579240000000
0!
0%
b10 *
0-
02
b10 6
#579250000000
1!
1%
1-
12
#579260000000
0!
0%
b11 *
0-
02
b11 6
#579270000000
1!
1%
1-
12
15
#579280000000
0!
0%
b100 *
0-
02
b100 6
#579290000000
1!
1%
1-
12
#579300000000
0!
0%
b101 *
0-
02
b101 6
#579310000000
1!
1%
1-
12
#579320000000
0!
0%
b110 *
0-
02
b110 6
#579330000000
1!
1%
1-
12
#579340000000
0!
0%
b111 *
0-
02
b111 6
#579350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#579360000000
0!
0%
b0 *
0-
02
b0 6
#579370000000
1!
1%
1-
12
#579380000000
0!
0%
b1 *
0-
02
b1 6
#579390000000
1!
1%
1-
12
#579400000000
0!
0%
b10 *
0-
02
b10 6
#579410000000
1!
1%
1-
12
#579420000000
0!
0%
b11 *
0-
02
b11 6
#579430000000
1!
1%
1-
12
15
#579440000000
0!
0%
b100 *
0-
02
b100 6
#579450000000
1!
1%
1-
12
#579460000000
0!
0%
b101 *
0-
02
b101 6
#579470000000
1!
1%
1-
12
#579480000000
0!
0%
b110 *
0-
02
b110 6
#579490000000
1!
1%
1-
12
#579500000000
0!
0%
b111 *
0-
02
b111 6
#579510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#579520000000
0!
0%
b0 *
0-
02
b0 6
#579530000000
1!
1%
1-
12
#579540000000
0!
0%
b1 *
0-
02
b1 6
#579550000000
1!
1%
1-
12
#579560000000
0!
0%
b10 *
0-
02
b10 6
#579570000000
1!
1%
1-
12
#579580000000
0!
0%
b11 *
0-
02
b11 6
#579590000000
1!
1%
1-
12
15
#579600000000
0!
0%
b100 *
0-
02
b100 6
#579610000000
1!
1%
1-
12
#579620000000
0!
0%
b101 *
0-
02
b101 6
#579630000000
1!
1%
1-
12
#579640000000
0!
0%
b110 *
0-
02
b110 6
#579650000000
1!
1%
1-
12
#579660000000
0!
0%
b111 *
0-
02
b111 6
#579670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#579680000000
0!
0%
b0 *
0-
02
b0 6
#579690000000
1!
1%
1-
12
#579700000000
0!
0%
b1 *
0-
02
b1 6
#579710000000
1!
1%
1-
12
#579720000000
0!
0%
b10 *
0-
02
b10 6
#579730000000
1!
1%
1-
12
#579740000000
0!
0%
b11 *
0-
02
b11 6
#579750000000
1!
1%
1-
12
15
#579760000000
0!
0%
b100 *
0-
02
b100 6
#579770000000
1!
1%
1-
12
#579780000000
0!
0%
b101 *
0-
02
b101 6
#579790000000
1!
1%
1-
12
#579800000000
0!
0%
b110 *
0-
02
b110 6
#579810000000
1!
1%
1-
12
#579820000000
0!
0%
b111 *
0-
02
b111 6
#579830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#579840000000
0!
0%
b0 *
0-
02
b0 6
#579850000000
1!
1%
1-
12
#579860000000
0!
0%
b1 *
0-
02
b1 6
#579870000000
1!
1%
1-
12
#579880000000
0!
0%
b10 *
0-
02
b10 6
#579890000000
1!
1%
1-
12
#579900000000
0!
0%
b11 *
0-
02
b11 6
#579910000000
1!
1%
1-
12
15
#579920000000
0!
0%
b100 *
0-
02
b100 6
#579930000000
1!
1%
1-
12
#579940000000
0!
0%
b101 *
0-
02
b101 6
#579950000000
1!
1%
1-
12
#579960000000
0!
0%
b110 *
0-
02
b110 6
#579970000000
1!
1%
1-
12
#579980000000
0!
0%
b111 *
0-
02
b111 6
#579990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#580000000000
0!
0%
b0 *
0-
02
b0 6
#580010000000
1!
1%
1-
12
#580020000000
0!
0%
b1 *
0-
02
b1 6
#580030000000
1!
1%
1-
12
#580040000000
0!
0%
b10 *
0-
02
b10 6
#580050000000
1!
1%
1-
12
#580060000000
0!
0%
b11 *
0-
02
b11 6
#580070000000
1!
1%
1-
12
15
#580080000000
0!
0%
b100 *
0-
02
b100 6
#580090000000
1!
1%
1-
12
#580100000000
0!
0%
b101 *
0-
02
b101 6
#580110000000
1!
1%
1-
12
#580120000000
0!
0%
b110 *
0-
02
b110 6
#580130000000
1!
1%
1-
12
#580140000000
0!
0%
b111 *
0-
02
b111 6
#580150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#580160000000
0!
0%
b0 *
0-
02
b0 6
#580170000000
1!
1%
1-
12
#580180000000
0!
0%
b1 *
0-
02
b1 6
#580190000000
1!
1%
1-
12
#580200000000
0!
0%
b10 *
0-
02
b10 6
#580210000000
1!
1%
1-
12
#580220000000
0!
0%
b11 *
0-
02
b11 6
#580230000000
1!
1%
1-
12
15
#580240000000
0!
0%
b100 *
0-
02
b100 6
#580250000000
1!
1%
1-
12
#580260000000
0!
0%
b101 *
0-
02
b101 6
#580270000000
1!
1%
1-
12
#580280000000
0!
0%
b110 *
0-
02
b110 6
#580290000000
1!
1%
1-
12
#580300000000
0!
0%
b111 *
0-
02
b111 6
#580310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#580320000000
0!
0%
b0 *
0-
02
b0 6
#580330000000
1!
1%
1-
12
#580340000000
0!
0%
b1 *
0-
02
b1 6
#580350000000
1!
1%
1-
12
#580360000000
0!
0%
b10 *
0-
02
b10 6
#580370000000
1!
1%
1-
12
#580380000000
0!
0%
b11 *
0-
02
b11 6
#580390000000
1!
1%
1-
12
15
#580400000000
0!
0%
b100 *
0-
02
b100 6
#580410000000
1!
1%
1-
12
#580420000000
0!
0%
b101 *
0-
02
b101 6
#580430000000
1!
1%
1-
12
#580440000000
0!
0%
b110 *
0-
02
b110 6
#580450000000
1!
1%
1-
12
#580460000000
0!
0%
b111 *
0-
02
b111 6
#580470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#580480000000
0!
0%
b0 *
0-
02
b0 6
#580490000000
1!
1%
1-
12
#580500000000
0!
0%
b1 *
0-
02
b1 6
#580510000000
1!
1%
1-
12
#580520000000
0!
0%
b10 *
0-
02
b10 6
#580530000000
1!
1%
1-
12
#580540000000
0!
0%
b11 *
0-
02
b11 6
#580550000000
1!
1%
1-
12
15
#580560000000
0!
0%
b100 *
0-
02
b100 6
#580570000000
1!
1%
1-
12
#580580000000
0!
0%
b101 *
0-
02
b101 6
#580590000000
1!
1%
1-
12
#580600000000
0!
0%
b110 *
0-
02
b110 6
#580610000000
1!
1%
1-
12
#580620000000
0!
0%
b111 *
0-
02
b111 6
#580630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#580640000000
0!
0%
b0 *
0-
02
b0 6
#580650000000
1!
1%
1-
12
#580660000000
0!
0%
b1 *
0-
02
b1 6
#580670000000
1!
1%
1-
12
#580680000000
0!
0%
b10 *
0-
02
b10 6
#580690000000
1!
1%
1-
12
#580700000000
0!
0%
b11 *
0-
02
b11 6
#580710000000
1!
1%
1-
12
15
#580720000000
0!
0%
b100 *
0-
02
b100 6
#580730000000
1!
1%
1-
12
#580740000000
0!
0%
b101 *
0-
02
b101 6
#580750000000
1!
1%
1-
12
#580760000000
0!
0%
b110 *
0-
02
b110 6
#580770000000
1!
1%
1-
12
#580780000000
0!
0%
b111 *
0-
02
b111 6
#580790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#580800000000
0!
0%
b0 *
0-
02
b0 6
#580810000000
1!
1%
1-
12
#580820000000
0!
0%
b1 *
0-
02
b1 6
#580830000000
1!
1%
1-
12
#580840000000
0!
0%
b10 *
0-
02
b10 6
#580850000000
1!
1%
1-
12
#580860000000
0!
0%
b11 *
0-
02
b11 6
#580870000000
1!
1%
1-
12
15
#580880000000
0!
0%
b100 *
0-
02
b100 6
#580890000000
1!
1%
1-
12
#580900000000
0!
0%
b101 *
0-
02
b101 6
#580910000000
1!
1%
1-
12
#580920000000
0!
0%
b110 *
0-
02
b110 6
#580930000000
1!
1%
1-
12
#580940000000
0!
0%
b111 *
0-
02
b111 6
#580950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#580960000000
0!
0%
b0 *
0-
02
b0 6
#580970000000
1!
1%
1-
12
#580980000000
0!
0%
b1 *
0-
02
b1 6
#580990000000
1!
1%
1-
12
#581000000000
0!
0%
b10 *
0-
02
b10 6
#581010000000
1!
1%
1-
12
#581020000000
0!
0%
b11 *
0-
02
b11 6
#581030000000
1!
1%
1-
12
15
#581040000000
0!
0%
b100 *
0-
02
b100 6
#581050000000
1!
1%
1-
12
#581060000000
0!
0%
b101 *
0-
02
b101 6
#581070000000
1!
1%
1-
12
#581080000000
0!
0%
b110 *
0-
02
b110 6
#581090000000
1!
1%
1-
12
#581100000000
0!
0%
b111 *
0-
02
b111 6
#581110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#581120000000
0!
0%
b0 *
0-
02
b0 6
#581130000000
1!
1%
1-
12
#581140000000
0!
0%
b1 *
0-
02
b1 6
#581150000000
1!
1%
1-
12
#581160000000
0!
0%
b10 *
0-
02
b10 6
#581170000000
1!
1%
1-
12
#581180000000
0!
0%
b11 *
0-
02
b11 6
#581190000000
1!
1%
1-
12
15
#581200000000
0!
0%
b100 *
0-
02
b100 6
#581210000000
1!
1%
1-
12
#581220000000
0!
0%
b101 *
0-
02
b101 6
#581230000000
1!
1%
1-
12
#581240000000
0!
0%
b110 *
0-
02
b110 6
#581250000000
1!
1%
1-
12
#581260000000
0!
0%
b111 *
0-
02
b111 6
#581270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#581280000000
0!
0%
b0 *
0-
02
b0 6
#581290000000
1!
1%
1-
12
#581300000000
0!
0%
b1 *
0-
02
b1 6
#581310000000
1!
1%
1-
12
#581320000000
0!
0%
b10 *
0-
02
b10 6
#581330000000
1!
1%
1-
12
#581340000000
0!
0%
b11 *
0-
02
b11 6
#581350000000
1!
1%
1-
12
15
#581360000000
0!
0%
b100 *
0-
02
b100 6
#581370000000
1!
1%
1-
12
#581380000000
0!
0%
b101 *
0-
02
b101 6
#581390000000
1!
1%
1-
12
#581400000000
0!
0%
b110 *
0-
02
b110 6
#581410000000
1!
1%
1-
12
#581420000000
0!
0%
b111 *
0-
02
b111 6
#581430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#581440000000
0!
0%
b0 *
0-
02
b0 6
#581450000000
1!
1%
1-
12
#581460000000
0!
0%
b1 *
0-
02
b1 6
#581470000000
1!
1%
1-
12
#581480000000
0!
0%
b10 *
0-
02
b10 6
#581490000000
1!
1%
1-
12
#581500000000
0!
0%
b11 *
0-
02
b11 6
#581510000000
1!
1%
1-
12
15
#581520000000
0!
0%
b100 *
0-
02
b100 6
#581530000000
1!
1%
1-
12
#581540000000
0!
0%
b101 *
0-
02
b101 6
#581550000000
1!
1%
1-
12
#581560000000
0!
0%
b110 *
0-
02
b110 6
#581570000000
1!
1%
1-
12
#581580000000
0!
0%
b111 *
0-
02
b111 6
#581590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#581600000000
0!
0%
b0 *
0-
02
b0 6
#581610000000
1!
1%
1-
12
#581620000000
0!
0%
b1 *
0-
02
b1 6
#581630000000
1!
1%
1-
12
#581640000000
0!
0%
b10 *
0-
02
b10 6
#581650000000
1!
1%
1-
12
#581660000000
0!
0%
b11 *
0-
02
b11 6
#581670000000
1!
1%
1-
12
15
#581680000000
0!
0%
b100 *
0-
02
b100 6
#581690000000
1!
1%
1-
12
#581700000000
0!
0%
b101 *
0-
02
b101 6
#581710000000
1!
1%
1-
12
#581720000000
0!
0%
b110 *
0-
02
b110 6
#581730000000
1!
1%
1-
12
#581740000000
0!
0%
b111 *
0-
02
b111 6
#581750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#581760000000
0!
0%
b0 *
0-
02
b0 6
#581770000000
1!
1%
1-
12
#581780000000
0!
0%
b1 *
0-
02
b1 6
#581790000000
1!
1%
1-
12
#581800000000
0!
0%
b10 *
0-
02
b10 6
#581810000000
1!
1%
1-
12
#581820000000
0!
0%
b11 *
0-
02
b11 6
#581830000000
1!
1%
1-
12
15
#581840000000
0!
0%
b100 *
0-
02
b100 6
#581850000000
1!
1%
1-
12
#581860000000
0!
0%
b101 *
0-
02
b101 6
#581870000000
1!
1%
1-
12
#581880000000
0!
0%
b110 *
0-
02
b110 6
#581890000000
1!
1%
1-
12
#581900000000
0!
0%
b111 *
0-
02
b111 6
#581910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#581920000000
0!
0%
b0 *
0-
02
b0 6
#581930000000
1!
1%
1-
12
#581940000000
0!
0%
b1 *
0-
02
b1 6
#581950000000
1!
1%
1-
12
#581960000000
0!
0%
b10 *
0-
02
b10 6
#581970000000
1!
1%
1-
12
#581980000000
0!
0%
b11 *
0-
02
b11 6
#581990000000
1!
1%
1-
12
15
#582000000000
0!
0%
b100 *
0-
02
b100 6
#582010000000
1!
1%
1-
12
#582020000000
0!
0%
b101 *
0-
02
b101 6
#582030000000
1!
1%
1-
12
#582040000000
0!
0%
b110 *
0-
02
b110 6
#582050000000
1!
1%
1-
12
#582060000000
0!
0%
b111 *
0-
02
b111 6
#582070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#582080000000
0!
0%
b0 *
0-
02
b0 6
#582090000000
1!
1%
1-
12
#582100000000
0!
0%
b1 *
0-
02
b1 6
#582110000000
1!
1%
1-
12
#582120000000
0!
0%
b10 *
0-
02
b10 6
#582130000000
1!
1%
1-
12
#582140000000
0!
0%
b11 *
0-
02
b11 6
#582150000000
1!
1%
1-
12
15
#582160000000
0!
0%
b100 *
0-
02
b100 6
#582170000000
1!
1%
1-
12
#582180000000
0!
0%
b101 *
0-
02
b101 6
#582190000000
1!
1%
1-
12
#582200000000
0!
0%
b110 *
0-
02
b110 6
#582210000000
1!
1%
1-
12
#582220000000
0!
0%
b111 *
0-
02
b111 6
#582230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#582240000000
0!
0%
b0 *
0-
02
b0 6
#582250000000
1!
1%
1-
12
#582260000000
0!
0%
b1 *
0-
02
b1 6
#582270000000
1!
1%
1-
12
#582280000000
0!
0%
b10 *
0-
02
b10 6
#582290000000
1!
1%
1-
12
#582300000000
0!
0%
b11 *
0-
02
b11 6
#582310000000
1!
1%
1-
12
15
#582320000000
0!
0%
b100 *
0-
02
b100 6
#582330000000
1!
1%
1-
12
#582340000000
0!
0%
b101 *
0-
02
b101 6
#582350000000
1!
1%
1-
12
#582360000000
0!
0%
b110 *
0-
02
b110 6
#582370000000
1!
1%
1-
12
#582380000000
0!
0%
b111 *
0-
02
b111 6
#582390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#582400000000
0!
0%
b0 *
0-
02
b0 6
#582410000000
1!
1%
1-
12
#582420000000
0!
0%
b1 *
0-
02
b1 6
#582430000000
1!
1%
1-
12
#582440000000
0!
0%
b10 *
0-
02
b10 6
#582450000000
1!
1%
1-
12
#582460000000
0!
0%
b11 *
0-
02
b11 6
#582470000000
1!
1%
1-
12
15
#582480000000
0!
0%
b100 *
0-
02
b100 6
#582490000000
1!
1%
1-
12
#582500000000
0!
0%
b101 *
0-
02
b101 6
#582510000000
1!
1%
1-
12
#582520000000
0!
0%
b110 *
0-
02
b110 6
#582530000000
1!
1%
1-
12
#582540000000
0!
0%
b111 *
0-
02
b111 6
#582550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#582560000000
0!
0%
b0 *
0-
02
b0 6
#582570000000
1!
1%
1-
12
#582580000000
0!
0%
b1 *
0-
02
b1 6
#582590000000
1!
1%
1-
12
#582600000000
0!
0%
b10 *
0-
02
b10 6
#582610000000
1!
1%
1-
12
#582620000000
0!
0%
b11 *
0-
02
b11 6
#582630000000
1!
1%
1-
12
15
#582640000000
0!
0%
b100 *
0-
02
b100 6
#582650000000
1!
1%
1-
12
#582660000000
0!
0%
b101 *
0-
02
b101 6
#582670000000
1!
1%
1-
12
#582680000000
0!
0%
b110 *
0-
02
b110 6
#582690000000
1!
1%
1-
12
#582700000000
0!
0%
b111 *
0-
02
b111 6
#582710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#582720000000
0!
0%
b0 *
0-
02
b0 6
#582730000000
1!
1%
1-
12
#582740000000
0!
0%
b1 *
0-
02
b1 6
#582750000000
1!
1%
1-
12
#582760000000
0!
0%
b10 *
0-
02
b10 6
#582770000000
1!
1%
1-
12
#582780000000
0!
0%
b11 *
0-
02
b11 6
#582790000000
1!
1%
1-
12
15
#582800000000
0!
0%
b100 *
0-
02
b100 6
#582810000000
1!
1%
1-
12
#582820000000
0!
0%
b101 *
0-
02
b101 6
#582830000000
1!
1%
1-
12
#582840000000
0!
0%
b110 *
0-
02
b110 6
#582850000000
1!
1%
1-
12
#582860000000
0!
0%
b111 *
0-
02
b111 6
#582870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#582880000000
0!
0%
b0 *
0-
02
b0 6
#582890000000
1!
1%
1-
12
#582900000000
0!
0%
b1 *
0-
02
b1 6
#582910000000
1!
1%
1-
12
#582920000000
0!
0%
b10 *
0-
02
b10 6
#582930000000
1!
1%
1-
12
#582940000000
0!
0%
b11 *
0-
02
b11 6
#582950000000
1!
1%
1-
12
15
#582960000000
0!
0%
b100 *
0-
02
b100 6
#582970000000
1!
1%
1-
12
#582980000000
0!
0%
b101 *
0-
02
b101 6
#582990000000
1!
1%
1-
12
#583000000000
0!
0%
b110 *
0-
02
b110 6
#583010000000
1!
1%
1-
12
#583020000000
0!
0%
b111 *
0-
02
b111 6
#583030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#583040000000
0!
0%
b0 *
0-
02
b0 6
#583050000000
1!
1%
1-
12
#583060000000
0!
0%
b1 *
0-
02
b1 6
#583070000000
1!
1%
1-
12
#583080000000
0!
0%
b10 *
0-
02
b10 6
#583090000000
1!
1%
1-
12
#583100000000
0!
0%
b11 *
0-
02
b11 6
#583110000000
1!
1%
1-
12
15
#583120000000
0!
0%
b100 *
0-
02
b100 6
#583130000000
1!
1%
1-
12
#583140000000
0!
0%
b101 *
0-
02
b101 6
#583150000000
1!
1%
1-
12
#583160000000
0!
0%
b110 *
0-
02
b110 6
#583170000000
1!
1%
1-
12
#583180000000
0!
0%
b111 *
0-
02
b111 6
#583190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#583200000000
0!
0%
b0 *
0-
02
b0 6
#583210000000
1!
1%
1-
12
#583220000000
0!
0%
b1 *
0-
02
b1 6
#583230000000
1!
1%
1-
12
#583240000000
0!
0%
b10 *
0-
02
b10 6
#583250000000
1!
1%
1-
12
#583260000000
0!
0%
b11 *
0-
02
b11 6
#583270000000
1!
1%
1-
12
15
#583280000000
0!
0%
b100 *
0-
02
b100 6
#583290000000
1!
1%
1-
12
#583300000000
0!
0%
b101 *
0-
02
b101 6
#583310000000
1!
1%
1-
12
#583320000000
0!
0%
b110 *
0-
02
b110 6
#583330000000
1!
1%
1-
12
#583340000000
0!
0%
b111 *
0-
02
b111 6
#583350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#583360000000
0!
0%
b0 *
0-
02
b0 6
#583370000000
1!
1%
1-
12
#583380000000
0!
0%
b1 *
0-
02
b1 6
#583390000000
1!
1%
1-
12
#583400000000
0!
0%
b10 *
0-
02
b10 6
#583410000000
1!
1%
1-
12
#583420000000
0!
0%
b11 *
0-
02
b11 6
#583430000000
1!
1%
1-
12
15
#583440000000
0!
0%
b100 *
0-
02
b100 6
#583450000000
1!
1%
1-
12
#583460000000
0!
0%
b101 *
0-
02
b101 6
#583470000000
1!
1%
1-
12
#583480000000
0!
0%
b110 *
0-
02
b110 6
#583490000000
1!
1%
1-
12
#583500000000
0!
0%
b111 *
0-
02
b111 6
#583510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#583520000000
0!
0%
b0 *
0-
02
b0 6
#583530000000
1!
1%
1-
12
#583540000000
0!
0%
b1 *
0-
02
b1 6
#583550000000
1!
1%
1-
12
#583560000000
0!
0%
b10 *
0-
02
b10 6
#583570000000
1!
1%
1-
12
#583580000000
0!
0%
b11 *
0-
02
b11 6
#583590000000
1!
1%
1-
12
15
#583600000000
0!
0%
b100 *
0-
02
b100 6
#583610000000
1!
1%
1-
12
#583620000000
0!
0%
b101 *
0-
02
b101 6
#583630000000
1!
1%
1-
12
#583640000000
0!
0%
b110 *
0-
02
b110 6
#583650000000
1!
1%
1-
12
#583660000000
0!
0%
b111 *
0-
02
b111 6
#583670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#583680000000
0!
0%
b0 *
0-
02
b0 6
#583690000000
1!
1%
1-
12
#583700000000
0!
0%
b1 *
0-
02
b1 6
#583710000000
1!
1%
1-
12
#583720000000
0!
0%
b10 *
0-
02
b10 6
#583730000000
1!
1%
1-
12
#583740000000
0!
0%
b11 *
0-
02
b11 6
#583750000000
1!
1%
1-
12
15
#583760000000
0!
0%
b100 *
0-
02
b100 6
#583770000000
1!
1%
1-
12
#583780000000
0!
0%
b101 *
0-
02
b101 6
#583790000000
1!
1%
1-
12
#583800000000
0!
0%
b110 *
0-
02
b110 6
#583810000000
1!
1%
1-
12
#583820000000
0!
0%
b111 *
0-
02
b111 6
#583830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#583840000000
0!
0%
b0 *
0-
02
b0 6
#583850000000
1!
1%
1-
12
#583860000000
0!
0%
b1 *
0-
02
b1 6
#583870000000
1!
1%
1-
12
#583880000000
0!
0%
b10 *
0-
02
b10 6
#583890000000
1!
1%
1-
12
#583900000000
0!
0%
b11 *
0-
02
b11 6
#583910000000
1!
1%
1-
12
15
#583920000000
0!
0%
b100 *
0-
02
b100 6
#583930000000
1!
1%
1-
12
#583940000000
0!
0%
b101 *
0-
02
b101 6
#583950000000
1!
1%
1-
12
#583960000000
0!
0%
b110 *
0-
02
b110 6
#583970000000
1!
1%
1-
12
#583980000000
0!
0%
b111 *
0-
02
b111 6
#583990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#584000000000
0!
0%
b0 *
0-
02
b0 6
#584010000000
1!
1%
1-
12
#584020000000
0!
0%
b1 *
0-
02
b1 6
#584030000000
1!
1%
1-
12
#584040000000
0!
0%
b10 *
0-
02
b10 6
#584050000000
1!
1%
1-
12
#584060000000
0!
0%
b11 *
0-
02
b11 6
#584070000000
1!
1%
1-
12
15
#584080000000
0!
0%
b100 *
0-
02
b100 6
#584090000000
1!
1%
1-
12
#584100000000
0!
0%
b101 *
0-
02
b101 6
#584110000000
1!
1%
1-
12
#584120000000
0!
0%
b110 *
0-
02
b110 6
#584130000000
1!
1%
1-
12
#584140000000
0!
0%
b111 *
0-
02
b111 6
#584150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#584160000000
0!
0%
b0 *
0-
02
b0 6
#584170000000
1!
1%
1-
12
#584180000000
0!
0%
b1 *
0-
02
b1 6
#584190000000
1!
1%
1-
12
#584200000000
0!
0%
b10 *
0-
02
b10 6
#584210000000
1!
1%
1-
12
#584220000000
0!
0%
b11 *
0-
02
b11 6
#584230000000
1!
1%
1-
12
15
#584240000000
0!
0%
b100 *
0-
02
b100 6
#584250000000
1!
1%
1-
12
#584260000000
0!
0%
b101 *
0-
02
b101 6
#584270000000
1!
1%
1-
12
#584280000000
0!
0%
b110 *
0-
02
b110 6
#584290000000
1!
1%
1-
12
#584300000000
0!
0%
b111 *
0-
02
b111 6
#584310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#584320000000
0!
0%
b0 *
0-
02
b0 6
#584330000000
1!
1%
1-
12
#584340000000
0!
0%
b1 *
0-
02
b1 6
#584350000000
1!
1%
1-
12
#584360000000
0!
0%
b10 *
0-
02
b10 6
#584370000000
1!
1%
1-
12
#584380000000
0!
0%
b11 *
0-
02
b11 6
#584390000000
1!
1%
1-
12
15
#584400000000
0!
0%
b100 *
0-
02
b100 6
#584410000000
1!
1%
1-
12
#584420000000
0!
0%
b101 *
0-
02
b101 6
#584430000000
1!
1%
1-
12
#584440000000
0!
0%
b110 *
0-
02
b110 6
#584450000000
1!
1%
1-
12
#584460000000
0!
0%
b111 *
0-
02
b111 6
#584470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#584480000000
0!
0%
b0 *
0-
02
b0 6
#584490000000
1!
1%
1-
12
#584500000000
0!
0%
b1 *
0-
02
b1 6
#584510000000
1!
1%
1-
12
#584520000000
0!
0%
b10 *
0-
02
b10 6
#584530000000
1!
1%
1-
12
#584540000000
0!
0%
b11 *
0-
02
b11 6
#584550000000
1!
1%
1-
12
15
#584560000000
0!
0%
b100 *
0-
02
b100 6
#584570000000
1!
1%
1-
12
#584580000000
0!
0%
b101 *
0-
02
b101 6
#584590000000
1!
1%
1-
12
#584600000000
0!
0%
b110 *
0-
02
b110 6
#584610000000
1!
1%
1-
12
#584620000000
0!
0%
b111 *
0-
02
b111 6
#584630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#584640000000
0!
0%
b0 *
0-
02
b0 6
#584650000000
1!
1%
1-
12
#584660000000
0!
0%
b1 *
0-
02
b1 6
#584670000000
1!
1%
1-
12
#584680000000
0!
0%
b10 *
0-
02
b10 6
#584690000000
1!
1%
1-
12
#584700000000
0!
0%
b11 *
0-
02
b11 6
#584710000000
1!
1%
1-
12
15
#584720000000
0!
0%
b100 *
0-
02
b100 6
#584730000000
1!
1%
1-
12
#584740000000
0!
0%
b101 *
0-
02
b101 6
#584750000000
1!
1%
1-
12
#584760000000
0!
0%
b110 *
0-
02
b110 6
#584770000000
1!
1%
1-
12
#584780000000
0!
0%
b111 *
0-
02
b111 6
#584790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#584800000000
0!
0%
b0 *
0-
02
b0 6
#584810000000
1!
1%
1-
12
#584820000000
0!
0%
b1 *
0-
02
b1 6
#584830000000
1!
1%
1-
12
#584840000000
0!
0%
b10 *
0-
02
b10 6
#584850000000
1!
1%
1-
12
#584860000000
0!
0%
b11 *
0-
02
b11 6
#584870000000
1!
1%
1-
12
15
#584880000000
0!
0%
b100 *
0-
02
b100 6
#584890000000
1!
1%
1-
12
#584900000000
0!
0%
b101 *
0-
02
b101 6
#584910000000
1!
1%
1-
12
#584920000000
0!
0%
b110 *
0-
02
b110 6
#584930000000
1!
1%
1-
12
#584940000000
0!
0%
b111 *
0-
02
b111 6
#584950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#584960000000
0!
0%
b0 *
0-
02
b0 6
#584970000000
1!
1%
1-
12
#584980000000
0!
0%
b1 *
0-
02
b1 6
#584990000000
1!
1%
1-
12
#585000000000
0!
0%
b10 *
0-
02
b10 6
#585010000000
1!
1%
1-
12
#585020000000
0!
0%
b11 *
0-
02
b11 6
#585030000000
1!
1%
1-
12
15
#585040000000
0!
0%
b100 *
0-
02
b100 6
#585050000000
1!
1%
1-
12
#585060000000
0!
0%
b101 *
0-
02
b101 6
#585070000000
1!
1%
1-
12
#585080000000
0!
0%
b110 *
0-
02
b110 6
#585090000000
1!
1%
1-
12
#585100000000
0!
0%
b111 *
0-
02
b111 6
#585110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#585120000000
0!
0%
b0 *
0-
02
b0 6
#585130000000
1!
1%
1-
12
#585140000000
0!
0%
b1 *
0-
02
b1 6
#585150000000
1!
1%
1-
12
#585160000000
0!
0%
b10 *
0-
02
b10 6
#585170000000
1!
1%
1-
12
#585180000000
0!
0%
b11 *
0-
02
b11 6
#585190000000
1!
1%
1-
12
15
#585200000000
0!
0%
b100 *
0-
02
b100 6
#585210000000
1!
1%
1-
12
#585220000000
0!
0%
b101 *
0-
02
b101 6
#585230000000
1!
1%
1-
12
#585240000000
0!
0%
b110 *
0-
02
b110 6
#585250000000
1!
1%
1-
12
#585260000000
0!
0%
b111 *
0-
02
b111 6
#585270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#585280000000
0!
0%
b0 *
0-
02
b0 6
#585290000000
1!
1%
1-
12
#585300000000
0!
0%
b1 *
0-
02
b1 6
#585310000000
1!
1%
1-
12
#585320000000
0!
0%
b10 *
0-
02
b10 6
#585330000000
1!
1%
1-
12
#585340000000
0!
0%
b11 *
0-
02
b11 6
#585350000000
1!
1%
1-
12
15
#585360000000
0!
0%
b100 *
0-
02
b100 6
#585370000000
1!
1%
1-
12
#585380000000
0!
0%
b101 *
0-
02
b101 6
#585390000000
1!
1%
1-
12
#585400000000
0!
0%
b110 *
0-
02
b110 6
#585410000000
1!
1%
1-
12
#585420000000
0!
0%
b111 *
0-
02
b111 6
#585430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#585440000000
0!
0%
b0 *
0-
02
b0 6
#585450000000
1!
1%
1-
12
#585460000000
0!
0%
b1 *
0-
02
b1 6
#585470000000
1!
1%
1-
12
#585480000000
0!
0%
b10 *
0-
02
b10 6
#585490000000
1!
1%
1-
12
#585500000000
0!
0%
b11 *
0-
02
b11 6
#585510000000
1!
1%
1-
12
15
#585520000000
0!
0%
b100 *
0-
02
b100 6
#585530000000
1!
1%
1-
12
#585540000000
0!
0%
b101 *
0-
02
b101 6
#585550000000
1!
1%
1-
12
#585560000000
0!
0%
b110 *
0-
02
b110 6
#585570000000
1!
1%
1-
12
#585580000000
0!
0%
b111 *
0-
02
b111 6
#585590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#585600000000
0!
0%
b0 *
0-
02
b0 6
#585610000000
1!
1%
1-
12
#585620000000
0!
0%
b1 *
0-
02
b1 6
#585630000000
1!
1%
1-
12
#585640000000
0!
0%
b10 *
0-
02
b10 6
#585650000000
1!
1%
1-
12
#585660000000
0!
0%
b11 *
0-
02
b11 6
#585670000000
1!
1%
1-
12
15
#585680000000
0!
0%
b100 *
0-
02
b100 6
#585690000000
1!
1%
1-
12
#585700000000
0!
0%
b101 *
0-
02
b101 6
#585710000000
1!
1%
1-
12
#585720000000
0!
0%
b110 *
0-
02
b110 6
#585730000000
1!
1%
1-
12
#585740000000
0!
0%
b111 *
0-
02
b111 6
#585750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#585760000000
0!
0%
b0 *
0-
02
b0 6
#585770000000
1!
1%
1-
12
#585780000000
0!
0%
b1 *
0-
02
b1 6
#585790000000
1!
1%
1-
12
#585800000000
0!
0%
b10 *
0-
02
b10 6
#585810000000
1!
1%
1-
12
#585820000000
0!
0%
b11 *
0-
02
b11 6
#585830000000
1!
1%
1-
12
15
#585840000000
0!
0%
b100 *
0-
02
b100 6
#585850000000
1!
1%
1-
12
#585860000000
0!
0%
b101 *
0-
02
b101 6
#585870000000
1!
1%
1-
12
#585880000000
0!
0%
b110 *
0-
02
b110 6
#585890000000
1!
1%
1-
12
#585900000000
0!
0%
b111 *
0-
02
b111 6
#585910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#585920000000
0!
0%
b0 *
0-
02
b0 6
#585930000000
1!
1%
1-
12
#585940000000
0!
0%
b1 *
0-
02
b1 6
#585950000000
1!
1%
1-
12
#585960000000
0!
0%
b10 *
0-
02
b10 6
#585970000000
1!
1%
1-
12
#585980000000
0!
0%
b11 *
0-
02
b11 6
#585990000000
1!
1%
1-
12
15
#586000000000
0!
0%
b100 *
0-
02
b100 6
#586010000000
1!
1%
1-
12
#586020000000
0!
0%
b101 *
0-
02
b101 6
#586030000000
1!
1%
1-
12
#586040000000
0!
0%
b110 *
0-
02
b110 6
#586050000000
1!
1%
1-
12
#586060000000
0!
0%
b111 *
0-
02
b111 6
#586070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#586080000000
0!
0%
b0 *
0-
02
b0 6
#586090000000
1!
1%
1-
12
#586100000000
0!
0%
b1 *
0-
02
b1 6
#586110000000
1!
1%
1-
12
#586120000000
0!
0%
b10 *
0-
02
b10 6
#586130000000
1!
1%
1-
12
#586140000000
0!
0%
b11 *
0-
02
b11 6
#586150000000
1!
1%
1-
12
15
#586160000000
0!
0%
b100 *
0-
02
b100 6
#586170000000
1!
1%
1-
12
#586180000000
0!
0%
b101 *
0-
02
b101 6
#586190000000
1!
1%
1-
12
#586200000000
0!
0%
b110 *
0-
02
b110 6
#586210000000
1!
1%
1-
12
#586220000000
0!
0%
b111 *
0-
02
b111 6
#586230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#586240000000
0!
0%
b0 *
0-
02
b0 6
#586250000000
1!
1%
1-
12
#586260000000
0!
0%
b1 *
0-
02
b1 6
#586270000000
1!
1%
1-
12
#586280000000
0!
0%
b10 *
0-
02
b10 6
#586290000000
1!
1%
1-
12
#586300000000
0!
0%
b11 *
0-
02
b11 6
#586310000000
1!
1%
1-
12
15
#586320000000
0!
0%
b100 *
0-
02
b100 6
#586330000000
1!
1%
1-
12
#586340000000
0!
0%
b101 *
0-
02
b101 6
#586350000000
1!
1%
1-
12
#586360000000
0!
0%
b110 *
0-
02
b110 6
#586370000000
1!
1%
1-
12
#586380000000
0!
0%
b111 *
0-
02
b111 6
#586390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#586400000000
0!
0%
b0 *
0-
02
b0 6
#586410000000
1!
1%
1-
12
#586420000000
0!
0%
b1 *
0-
02
b1 6
#586430000000
1!
1%
1-
12
#586440000000
0!
0%
b10 *
0-
02
b10 6
#586450000000
1!
1%
1-
12
#586460000000
0!
0%
b11 *
0-
02
b11 6
#586470000000
1!
1%
1-
12
15
#586480000000
0!
0%
b100 *
0-
02
b100 6
#586490000000
1!
1%
1-
12
#586500000000
0!
0%
b101 *
0-
02
b101 6
#586510000000
1!
1%
1-
12
#586520000000
0!
0%
b110 *
0-
02
b110 6
#586530000000
1!
1%
1-
12
#586540000000
0!
0%
b111 *
0-
02
b111 6
#586550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#586560000000
0!
0%
b0 *
0-
02
b0 6
#586570000000
1!
1%
1-
12
#586580000000
0!
0%
b1 *
0-
02
b1 6
#586590000000
1!
1%
1-
12
#586600000000
0!
0%
b10 *
0-
02
b10 6
#586610000000
1!
1%
1-
12
#586620000000
0!
0%
b11 *
0-
02
b11 6
#586630000000
1!
1%
1-
12
15
#586640000000
0!
0%
b100 *
0-
02
b100 6
#586650000000
1!
1%
1-
12
#586660000000
0!
0%
b101 *
0-
02
b101 6
#586670000000
1!
1%
1-
12
#586680000000
0!
0%
b110 *
0-
02
b110 6
#586690000000
1!
1%
1-
12
#586700000000
0!
0%
b111 *
0-
02
b111 6
#586710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#586720000000
0!
0%
b0 *
0-
02
b0 6
#586730000000
1!
1%
1-
12
#586740000000
0!
0%
b1 *
0-
02
b1 6
#586750000000
1!
1%
1-
12
#586760000000
0!
0%
b10 *
0-
02
b10 6
#586770000000
1!
1%
1-
12
#586780000000
0!
0%
b11 *
0-
02
b11 6
#586790000000
1!
1%
1-
12
15
#586800000000
0!
0%
b100 *
0-
02
b100 6
#586810000000
1!
1%
1-
12
#586820000000
0!
0%
b101 *
0-
02
b101 6
#586830000000
1!
1%
1-
12
#586840000000
0!
0%
b110 *
0-
02
b110 6
#586850000000
1!
1%
1-
12
#586860000000
0!
0%
b111 *
0-
02
b111 6
#586870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#586880000000
0!
0%
b0 *
0-
02
b0 6
#586890000000
1!
1%
1-
12
#586900000000
0!
0%
b1 *
0-
02
b1 6
#586910000000
1!
1%
1-
12
#586920000000
0!
0%
b10 *
0-
02
b10 6
#586930000000
1!
1%
1-
12
#586940000000
0!
0%
b11 *
0-
02
b11 6
#586950000000
1!
1%
1-
12
15
#586960000000
0!
0%
b100 *
0-
02
b100 6
#586970000000
1!
1%
1-
12
#586980000000
0!
0%
b101 *
0-
02
b101 6
#586990000000
1!
1%
1-
12
#587000000000
0!
0%
b110 *
0-
02
b110 6
#587010000000
1!
1%
1-
12
#587020000000
0!
0%
b111 *
0-
02
b111 6
#587030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#587040000000
0!
0%
b0 *
0-
02
b0 6
#587050000000
1!
1%
1-
12
#587060000000
0!
0%
b1 *
0-
02
b1 6
#587070000000
1!
1%
1-
12
#587080000000
0!
0%
b10 *
0-
02
b10 6
#587090000000
1!
1%
1-
12
#587100000000
0!
0%
b11 *
0-
02
b11 6
#587110000000
1!
1%
1-
12
15
#587120000000
0!
0%
b100 *
0-
02
b100 6
#587130000000
1!
1%
1-
12
#587140000000
0!
0%
b101 *
0-
02
b101 6
#587150000000
1!
1%
1-
12
#587160000000
0!
0%
b110 *
0-
02
b110 6
#587170000000
1!
1%
1-
12
#587180000000
0!
0%
b111 *
0-
02
b111 6
#587190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#587200000000
0!
0%
b0 *
0-
02
b0 6
#587210000000
1!
1%
1-
12
#587220000000
0!
0%
b1 *
0-
02
b1 6
#587230000000
1!
1%
1-
12
#587240000000
0!
0%
b10 *
0-
02
b10 6
#587250000000
1!
1%
1-
12
#587260000000
0!
0%
b11 *
0-
02
b11 6
#587270000000
1!
1%
1-
12
15
#587280000000
0!
0%
b100 *
0-
02
b100 6
#587290000000
1!
1%
1-
12
#587300000000
0!
0%
b101 *
0-
02
b101 6
#587310000000
1!
1%
1-
12
#587320000000
0!
0%
b110 *
0-
02
b110 6
#587330000000
1!
1%
1-
12
#587340000000
0!
0%
b111 *
0-
02
b111 6
#587350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#587360000000
0!
0%
b0 *
0-
02
b0 6
#587370000000
1!
1%
1-
12
#587380000000
0!
0%
b1 *
0-
02
b1 6
#587390000000
1!
1%
1-
12
#587400000000
0!
0%
b10 *
0-
02
b10 6
#587410000000
1!
1%
1-
12
#587420000000
0!
0%
b11 *
0-
02
b11 6
#587430000000
1!
1%
1-
12
15
#587440000000
0!
0%
b100 *
0-
02
b100 6
#587450000000
1!
1%
1-
12
#587460000000
0!
0%
b101 *
0-
02
b101 6
#587470000000
1!
1%
1-
12
#587480000000
0!
0%
b110 *
0-
02
b110 6
#587490000000
1!
1%
1-
12
#587500000000
0!
0%
b111 *
0-
02
b111 6
#587510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#587520000000
0!
0%
b0 *
0-
02
b0 6
#587530000000
1!
1%
1-
12
#587540000000
0!
0%
b1 *
0-
02
b1 6
#587550000000
1!
1%
1-
12
#587560000000
0!
0%
b10 *
0-
02
b10 6
#587570000000
1!
1%
1-
12
#587580000000
0!
0%
b11 *
0-
02
b11 6
#587590000000
1!
1%
1-
12
15
#587600000000
0!
0%
b100 *
0-
02
b100 6
#587610000000
1!
1%
1-
12
#587620000000
0!
0%
b101 *
0-
02
b101 6
#587630000000
1!
1%
1-
12
#587640000000
0!
0%
b110 *
0-
02
b110 6
#587650000000
1!
1%
1-
12
#587660000000
0!
0%
b111 *
0-
02
b111 6
#587670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#587680000000
0!
0%
b0 *
0-
02
b0 6
#587690000000
1!
1%
1-
12
#587700000000
0!
0%
b1 *
0-
02
b1 6
#587710000000
1!
1%
1-
12
#587720000000
0!
0%
b10 *
0-
02
b10 6
#587730000000
1!
1%
1-
12
#587740000000
0!
0%
b11 *
0-
02
b11 6
#587750000000
1!
1%
1-
12
15
#587760000000
0!
0%
b100 *
0-
02
b100 6
#587770000000
1!
1%
1-
12
#587780000000
0!
0%
b101 *
0-
02
b101 6
#587790000000
1!
1%
1-
12
#587800000000
0!
0%
b110 *
0-
02
b110 6
#587810000000
1!
1%
1-
12
#587820000000
0!
0%
b111 *
0-
02
b111 6
#587830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#587840000000
0!
0%
b0 *
0-
02
b0 6
#587850000000
1!
1%
1-
12
#587860000000
0!
0%
b1 *
0-
02
b1 6
#587870000000
1!
1%
1-
12
#587880000000
0!
0%
b10 *
0-
02
b10 6
#587890000000
1!
1%
1-
12
#587900000000
0!
0%
b11 *
0-
02
b11 6
#587910000000
1!
1%
1-
12
15
#587920000000
0!
0%
b100 *
0-
02
b100 6
#587930000000
1!
1%
1-
12
#587940000000
0!
0%
b101 *
0-
02
b101 6
#587950000000
1!
1%
1-
12
#587960000000
0!
0%
b110 *
0-
02
b110 6
#587970000000
1!
1%
1-
12
#587980000000
0!
0%
b111 *
0-
02
b111 6
#587990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#588000000000
0!
0%
b0 *
0-
02
b0 6
#588010000000
1!
1%
1-
12
#588020000000
0!
0%
b1 *
0-
02
b1 6
#588030000000
1!
1%
1-
12
#588040000000
0!
0%
b10 *
0-
02
b10 6
#588050000000
1!
1%
1-
12
#588060000000
0!
0%
b11 *
0-
02
b11 6
#588070000000
1!
1%
1-
12
15
#588080000000
0!
0%
b100 *
0-
02
b100 6
#588090000000
1!
1%
1-
12
#588100000000
0!
0%
b101 *
0-
02
b101 6
#588110000000
1!
1%
1-
12
#588120000000
0!
0%
b110 *
0-
02
b110 6
#588130000000
1!
1%
1-
12
#588140000000
0!
0%
b111 *
0-
02
b111 6
#588150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#588160000000
0!
0%
b0 *
0-
02
b0 6
#588170000000
1!
1%
1-
12
#588180000000
0!
0%
b1 *
0-
02
b1 6
#588190000000
1!
1%
1-
12
#588200000000
0!
0%
b10 *
0-
02
b10 6
#588210000000
1!
1%
1-
12
#588220000000
0!
0%
b11 *
0-
02
b11 6
#588230000000
1!
1%
1-
12
15
#588240000000
0!
0%
b100 *
0-
02
b100 6
#588250000000
1!
1%
1-
12
#588260000000
0!
0%
b101 *
0-
02
b101 6
#588270000000
1!
1%
1-
12
#588280000000
0!
0%
b110 *
0-
02
b110 6
#588290000000
1!
1%
1-
12
#588300000000
0!
0%
b111 *
0-
02
b111 6
#588310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#588320000000
0!
0%
b0 *
0-
02
b0 6
#588330000000
1!
1%
1-
12
#588340000000
0!
0%
b1 *
0-
02
b1 6
#588350000000
1!
1%
1-
12
#588360000000
0!
0%
b10 *
0-
02
b10 6
#588370000000
1!
1%
1-
12
#588380000000
0!
0%
b11 *
0-
02
b11 6
#588390000000
1!
1%
1-
12
15
#588400000000
0!
0%
b100 *
0-
02
b100 6
#588410000000
1!
1%
1-
12
#588420000000
0!
0%
b101 *
0-
02
b101 6
#588430000000
1!
1%
1-
12
#588440000000
0!
0%
b110 *
0-
02
b110 6
#588450000000
1!
1%
1-
12
#588460000000
0!
0%
b111 *
0-
02
b111 6
#588470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#588480000000
0!
0%
b0 *
0-
02
b0 6
#588490000000
1!
1%
1-
12
#588500000000
0!
0%
b1 *
0-
02
b1 6
#588510000000
1!
1%
1-
12
#588520000000
0!
0%
b10 *
0-
02
b10 6
#588530000000
1!
1%
1-
12
#588540000000
0!
0%
b11 *
0-
02
b11 6
#588550000000
1!
1%
1-
12
15
#588560000000
0!
0%
b100 *
0-
02
b100 6
#588570000000
1!
1%
1-
12
#588580000000
0!
0%
b101 *
0-
02
b101 6
#588590000000
1!
1%
1-
12
#588600000000
0!
0%
b110 *
0-
02
b110 6
#588610000000
1!
1%
1-
12
#588620000000
0!
0%
b111 *
0-
02
b111 6
#588630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#588640000000
0!
0%
b0 *
0-
02
b0 6
#588650000000
1!
1%
1-
12
#588660000000
0!
0%
b1 *
0-
02
b1 6
#588670000000
1!
1%
1-
12
#588680000000
0!
0%
b10 *
0-
02
b10 6
#588690000000
1!
1%
1-
12
#588700000000
0!
0%
b11 *
0-
02
b11 6
#588710000000
1!
1%
1-
12
15
#588720000000
0!
0%
b100 *
0-
02
b100 6
#588730000000
1!
1%
1-
12
#588740000000
0!
0%
b101 *
0-
02
b101 6
#588750000000
1!
1%
1-
12
#588760000000
0!
0%
b110 *
0-
02
b110 6
#588770000000
1!
1%
1-
12
#588780000000
0!
0%
b111 *
0-
02
b111 6
#588790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#588800000000
0!
0%
b0 *
0-
02
b0 6
#588810000000
1!
1%
1-
12
#588820000000
0!
0%
b1 *
0-
02
b1 6
#588830000000
1!
1%
1-
12
#588840000000
0!
0%
b10 *
0-
02
b10 6
#588850000000
1!
1%
1-
12
#588860000000
0!
0%
b11 *
0-
02
b11 6
#588870000000
1!
1%
1-
12
15
#588880000000
0!
0%
b100 *
0-
02
b100 6
#588890000000
1!
1%
1-
12
#588900000000
0!
0%
b101 *
0-
02
b101 6
#588910000000
1!
1%
1-
12
#588920000000
0!
0%
b110 *
0-
02
b110 6
#588930000000
1!
1%
1-
12
#588940000000
0!
0%
b111 *
0-
02
b111 6
#588950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#588960000000
0!
0%
b0 *
0-
02
b0 6
#588970000000
1!
1%
1-
12
#588980000000
0!
0%
b1 *
0-
02
b1 6
#588990000000
1!
1%
1-
12
#589000000000
0!
0%
b10 *
0-
02
b10 6
#589010000000
1!
1%
1-
12
#589020000000
0!
0%
b11 *
0-
02
b11 6
#589030000000
1!
1%
1-
12
15
#589040000000
0!
0%
b100 *
0-
02
b100 6
#589050000000
1!
1%
1-
12
#589060000000
0!
0%
b101 *
0-
02
b101 6
#589070000000
1!
1%
1-
12
#589080000000
0!
0%
b110 *
0-
02
b110 6
#589090000000
1!
1%
1-
12
#589100000000
0!
0%
b111 *
0-
02
b111 6
#589110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#589120000000
0!
0%
b0 *
0-
02
b0 6
#589130000000
1!
1%
1-
12
#589140000000
0!
0%
b1 *
0-
02
b1 6
#589150000000
1!
1%
1-
12
#589160000000
0!
0%
b10 *
0-
02
b10 6
#589170000000
1!
1%
1-
12
#589180000000
0!
0%
b11 *
0-
02
b11 6
#589190000000
1!
1%
1-
12
15
#589200000000
0!
0%
b100 *
0-
02
b100 6
#589210000000
1!
1%
1-
12
#589220000000
0!
0%
b101 *
0-
02
b101 6
#589230000000
1!
1%
1-
12
#589240000000
0!
0%
b110 *
0-
02
b110 6
#589250000000
1!
1%
1-
12
#589260000000
0!
0%
b111 *
0-
02
b111 6
#589270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#589280000000
0!
0%
b0 *
0-
02
b0 6
#589290000000
1!
1%
1-
12
#589300000000
0!
0%
b1 *
0-
02
b1 6
#589310000000
1!
1%
1-
12
#589320000000
0!
0%
b10 *
0-
02
b10 6
#589330000000
1!
1%
1-
12
#589340000000
0!
0%
b11 *
0-
02
b11 6
#589350000000
1!
1%
1-
12
15
#589360000000
0!
0%
b100 *
0-
02
b100 6
#589370000000
1!
1%
1-
12
#589380000000
0!
0%
b101 *
0-
02
b101 6
#589390000000
1!
1%
1-
12
#589400000000
0!
0%
b110 *
0-
02
b110 6
#589410000000
1!
1%
1-
12
#589420000000
0!
0%
b111 *
0-
02
b111 6
#589430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#589440000000
0!
0%
b0 *
0-
02
b0 6
#589450000000
1!
1%
1-
12
#589460000000
0!
0%
b1 *
0-
02
b1 6
#589470000000
1!
1%
1-
12
#589480000000
0!
0%
b10 *
0-
02
b10 6
#589490000000
1!
1%
1-
12
#589500000000
0!
0%
b11 *
0-
02
b11 6
#589510000000
1!
1%
1-
12
15
#589520000000
0!
0%
b100 *
0-
02
b100 6
#589530000000
1!
1%
1-
12
#589540000000
0!
0%
b101 *
0-
02
b101 6
#589550000000
1!
1%
1-
12
#589560000000
0!
0%
b110 *
0-
02
b110 6
#589570000000
1!
1%
1-
12
#589580000000
0!
0%
b111 *
0-
02
b111 6
#589590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#589600000000
0!
0%
b0 *
0-
02
b0 6
#589610000000
1!
1%
1-
12
#589620000000
0!
0%
b1 *
0-
02
b1 6
#589630000000
1!
1%
1-
12
#589640000000
0!
0%
b10 *
0-
02
b10 6
#589650000000
1!
1%
1-
12
#589660000000
0!
0%
b11 *
0-
02
b11 6
#589670000000
1!
1%
1-
12
15
#589680000000
0!
0%
b100 *
0-
02
b100 6
#589690000000
1!
1%
1-
12
#589700000000
0!
0%
b101 *
0-
02
b101 6
#589710000000
1!
1%
1-
12
#589720000000
0!
0%
b110 *
0-
02
b110 6
#589730000000
1!
1%
1-
12
#589740000000
0!
0%
b111 *
0-
02
b111 6
#589750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#589760000000
0!
0%
b0 *
0-
02
b0 6
#589770000000
1!
1%
1-
12
#589780000000
0!
0%
b1 *
0-
02
b1 6
#589790000000
1!
1%
1-
12
#589800000000
0!
0%
b10 *
0-
02
b10 6
#589810000000
1!
1%
1-
12
#589820000000
0!
0%
b11 *
0-
02
b11 6
#589830000000
1!
1%
1-
12
15
#589840000000
0!
0%
b100 *
0-
02
b100 6
#589850000000
1!
1%
1-
12
#589860000000
0!
0%
b101 *
0-
02
b101 6
#589870000000
1!
1%
1-
12
#589880000000
0!
0%
b110 *
0-
02
b110 6
#589890000000
1!
1%
1-
12
#589900000000
0!
0%
b111 *
0-
02
b111 6
#589910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#589920000000
0!
0%
b0 *
0-
02
b0 6
#589930000000
1!
1%
1-
12
#589940000000
0!
0%
b1 *
0-
02
b1 6
#589950000000
1!
1%
1-
12
#589960000000
0!
0%
b10 *
0-
02
b10 6
#589970000000
1!
1%
1-
12
#589980000000
0!
0%
b11 *
0-
02
b11 6
#589990000000
1!
1%
1-
12
15
#590000000000
0!
0%
b100 *
0-
02
b100 6
#590010000000
1!
1%
1-
12
#590020000000
0!
0%
b101 *
0-
02
b101 6
#590030000000
1!
1%
1-
12
#590040000000
0!
0%
b110 *
0-
02
b110 6
#590050000000
1!
1%
1-
12
#590060000000
0!
0%
b111 *
0-
02
b111 6
#590070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#590080000000
0!
0%
b0 *
0-
02
b0 6
#590090000000
1!
1%
1-
12
#590100000000
0!
0%
b1 *
0-
02
b1 6
#590110000000
1!
1%
1-
12
#590120000000
0!
0%
b10 *
0-
02
b10 6
#590130000000
1!
1%
1-
12
#590140000000
0!
0%
b11 *
0-
02
b11 6
#590150000000
1!
1%
1-
12
15
#590160000000
0!
0%
b100 *
0-
02
b100 6
#590170000000
1!
1%
1-
12
#590180000000
0!
0%
b101 *
0-
02
b101 6
#590190000000
1!
1%
1-
12
#590200000000
0!
0%
b110 *
0-
02
b110 6
#590210000000
1!
1%
1-
12
#590220000000
0!
0%
b111 *
0-
02
b111 6
#590230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#590240000000
0!
0%
b0 *
0-
02
b0 6
#590250000000
1!
1%
1-
12
#590260000000
0!
0%
b1 *
0-
02
b1 6
#590270000000
1!
1%
1-
12
#590280000000
0!
0%
b10 *
0-
02
b10 6
#590290000000
1!
1%
1-
12
#590300000000
0!
0%
b11 *
0-
02
b11 6
#590310000000
1!
1%
1-
12
15
#590320000000
0!
0%
b100 *
0-
02
b100 6
#590330000000
1!
1%
1-
12
#590340000000
0!
0%
b101 *
0-
02
b101 6
#590350000000
1!
1%
1-
12
#590360000000
0!
0%
b110 *
0-
02
b110 6
#590370000000
1!
1%
1-
12
#590380000000
0!
0%
b111 *
0-
02
b111 6
#590390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#590400000000
0!
0%
b0 *
0-
02
b0 6
#590410000000
1!
1%
1-
12
#590420000000
0!
0%
b1 *
0-
02
b1 6
#590430000000
1!
1%
1-
12
#590440000000
0!
0%
b10 *
0-
02
b10 6
#590450000000
1!
1%
1-
12
#590460000000
0!
0%
b11 *
0-
02
b11 6
#590470000000
1!
1%
1-
12
15
#590480000000
0!
0%
b100 *
0-
02
b100 6
#590490000000
1!
1%
1-
12
#590500000000
0!
0%
b101 *
0-
02
b101 6
#590510000000
1!
1%
1-
12
#590520000000
0!
0%
b110 *
0-
02
b110 6
#590530000000
1!
1%
1-
12
#590540000000
0!
0%
b111 *
0-
02
b111 6
#590550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#590560000000
0!
0%
b0 *
0-
02
b0 6
#590570000000
1!
1%
1-
12
#590580000000
0!
0%
b1 *
0-
02
b1 6
#590590000000
1!
1%
1-
12
#590600000000
0!
0%
b10 *
0-
02
b10 6
#590610000000
1!
1%
1-
12
#590620000000
0!
0%
b11 *
0-
02
b11 6
#590630000000
1!
1%
1-
12
15
#590640000000
0!
0%
b100 *
0-
02
b100 6
#590650000000
1!
1%
1-
12
#590660000000
0!
0%
b101 *
0-
02
b101 6
#590670000000
1!
1%
1-
12
#590680000000
0!
0%
b110 *
0-
02
b110 6
#590690000000
1!
1%
1-
12
#590700000000
0!
0%
b111 *
0-
02
b111 6
#590710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#590720000000
0!
0%
b0 *
0-
02
b0 6
#590730000000
1!
1%
1-
12
#590740000000
0!
0%
b1 *
0-
02
b1 6
#590750000000
1!
1%
1-
12
#590760000000
0!
0%
b10 *
0-
02
b10 6
#590770000000
1!
1%
1-
12
#590780000000
0!
0%
b11 *
0-
02
b11 6
#590790000000
1!
1%
1-
12
15
#590800000000
0!
0%
b100 *
0-
02
b100 6
#590810000000
1!
1%
1-
12
#590820000000
0!
0%
b101 *
0-
02
b101 6
#590830000000
1!
1%
1-
12
#590840000000
0!
0%
b110 *
0-
02
b110 6
#590850000000
1!
1%
1-
12
#590860000000
0!
0%
b111 *
0-
02
b111 6
#590870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#590880000000
0!
0%
b0 *
0-
02
b0 6
#590890000000
1!
1%
1-
12
#590900000000
0!
0%
b1 *
0-
02
b1 6
#590910000000
1!
1%
1-
12
#590920000000
0!
0%
b10 *
0-
02
b10 6
#590930000000
1!
1%
1-
12
#590940000000
0!
0%
b11 *
0-
02
b11 6
#590950000000
1!
1%
1-
12
15
#590960000000
0!
0%
b100 *
0-
02
b100 6
#590970000000
1!
1%
1-
12
#590980000000
0!
0%
b101 *
0-
02
b101 6
#590990000000
1!
1%
1-
12
#591000000000
0!
0%
b110 *
0-
02
b110 6
#591010000000
1!
1%
1-
12
#591020000000
0!
0%
b111 *
0-
02
b111 6
#591030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#591040000000
0!
0%
b0 *
0-
02
b0 6
#591050000000
1!
1%
1-
12
#591060000000
0!
0%
b1 *
0-
02
b1 6
#591070000000
1!
1%
1-
12
#591080000000
0!
0%
b10 *
0-
02
b10 6
#591090000000
1!
1%
1-
12
#591100000000
0!
0%
b11 *
0-
02
b11 6
#591110000000
1!
1%
1-
12
15
#591120000000
0!
0%
b100 *
0-
02
b100 6
#591130000000
1!
1%
1-
12
#591140000000
0!
0%
b101 *
0-
02
b101 6
#591150000000
1!
1%
1-
12
#591160000000
0!
0%
b110 *
0-
02
b110 6
#591170000000
1!
1%
1-
12
#591180000000
0!
0%
b111 *
0-
02
b111 6
#591190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#591200000000
0!
0%
b0 *
0-
02
b0 6
#591210000000
1!
1%
1-
12
#591220000000
0!
0%
b1 *
0-
02
b1 6
#591230000000
1!
1%
1-
12
#591240000000
0!
0%
b10 *
0-
02
b10 6
#591250000000
1!
1%
1-
12
#591260000000
0!
0%
b11 *
0-
02
b11 6
#591270000000
1!
1%
1-
12
15
#591280000000
0!
0%
b100 *
0-
02
b100 6
#591290000000
1!
1%
1-
12
#591300000000
0!
0%
b101 *
0-
02
b101 6
#591310000000
1!
1%
1-
12
#591320000000
0!
0%
b110 *
0-
02
b110 6
#591330000000
1!
1%
1-
12
#591340000000
0!
0%
b111 *
0-
02
b111 6
#591350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#591360000000
0!
0%
b0 *
0-
02
b0 6
#591370000000
1!
1%
1-
12
#591380000000
0!
0%
b1 *
0-
02
b1 6
#591390000000
1!
1%
1-
12
#591400000000
0!
0%
b10 *
0-
02
b10 6
#591410000000
1!
1%
1-
12
#591420000000
0!
0%
b11 *
0-
02
b11 6
#591430000000
1!
1%
1-
12
15
#591440000000
0!
0%
b100 *
0-
02
b100 6
#591450000000
1!
1%
1-
12
#591460000000
0!
0%
b101 *
0-
02
b101 6
#591470000000
1!
1%
1-
12
#591480000000
0!
0%
b110 *
0-
02
b110 6
#591490000000
1!
1%
1-
12
#591500000000
0!
0%
b111 *
0-
02
b111 6
#591510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#591520000000
0!
0%
b0 *
0-
02
b0 6
#591530000000
1!
1%
1-
12
#591540000000
0!
0%
b1 *
0-
02
b1 6
#591550000000
1!
1%
1-
12
#591560000000
0!
0%
b10 *
0-
02
b10 6
#591570000000
1!
1%
1-
12
#591580000000
0!
0%
b11 *
0-
02
b11 6
#591590000000
1!
1%
1-
12
15
#591600000000
0!
0%
b100 *
0-
02
b100 6
#591610000000
1!
1%
1-
12
#591620000000
0!
0%
b101 *
0-
02
b101 6
#591630000000
1!
1%
1-
12
#591640000000
0!
0%
b110 *
0-
02
b110 6
#591650000000
1!
1%
1-
12
#591660000000
0!
0%
b111 *
0-
02
b111 6
#591670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#591680000000
0!
0%
b0 *
0-
02
b0 6
#591690000000
1!
1%
1-
12
#591700000000
0!
0%
b1 *
0-
02
b1 6
#591710000000
1!
1%
1-
12
#591720000000
0!
0%
b10 *
0-
02
b10 6
#591730000000
1!
1%
1-
12
#591740000000
0!
0%
b11 *
0-
02
b11 6
#591750000000
1!
1%
1-
12
15
#591760000000
0!
0%
b100 *
0-
02
b100 6
#591770000000
1!
1%
1-
12
#591780000000
0!
0%
b101 *
0-
02
b101 6
#591790000000
1!
1%
1-
12
#591800000000
0!
0%
b110 *
0-
02
b110 6
#591810000000
1!
1%
1-
12
#591820000000
0!
0%
b111 *
0-
02
b111 6
#591830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#591840000000
0!
0%
b0 *
0-
02
b0 6
#591850000000
1!
1%
1-
12
#591860000000
0!
0%
b1 *
0-
02
b1 6
#591870000000
1!
1%
1-
12
#591880000000
0!
0%
b10 *
0-
02
b10 6
#591890000000
1!
1%
1-
12
#591900000000
0!
0%
b11 *
0-
02
b11 6
#591910000000
1!
1%
1-
12
15
#591920000000
0!
0%
b100 *
0-
02
b100 6
#591930000000
1!
1%
1-
12
#591940000000
0!
0%
b101 *
0-
02
b101 6
#591950000000
1!
1%
1-
12
#591960000000
0!
0%
b110 *
0-
02
b110 6
#591970000000
1!
1%
1-
12
#591980000000
0!
0%
b111 *
0-
02
b111 6
#591990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#592000000000
0!
0%
b0 *
0-
02
b0 6
#592010000000
1!
1%
1-
12
#592020000000
0!
0%
b1 *
0-
02
b1 6
#592030000000
1!
1%
1-
12
#592040000000
0!
0%
b10 *
0-
02
b10 6
#592050000000
1!
1%
1-
12
#592060000000
0!
0%
b11 *
0-
02
b11 6
#592070000000
1!
1%
1-
12
15
#592080000000
0!
0%
b100 *
0-
02
b100 6
#592090000000
1!
1%
1-
12
#592100000000
0!
0%
b101 *
0-
02
b101 6
#592110000000
1!
1%
1-
12
#592120000000
0!
0%
b110 *
0-
02
b110 6
#592130000000
1!
1%
1-
12
#592140000000
0!
0%
b111 *
0-
02
b111 6
#592150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#592160000000
0!
0%
b0 *
0-
02
b0 6
#592170000000
1!
1%
1-
12
#592180000000
0!
0%
b1 *
0-
02
b1 6
#592190000000
1!
1%
1-
12
#592200000000
0!
0%
b10 *
0-
02
b10 6
#592210000000
1!
1%
1-
12
#592220000000
0!
0%
b11 *
0-
02
b11 6
#592230000000
1!
1%
1-
12
15
#592240000000
0!
0%
b100 *
0-
02
b100 6
#592250000000
1!
1%
1-
12
#592260000000
0!
0%
b101 *
0-
02
b101 6
#592270000000
1!
1%
1-
12
#592280000000
0!
0%
b110 *
0-
02
b110 6
#592290000000
1!
1%
1-
12
#592300000000
0!
0%
b111 *
0-
02
b111 6
#592310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#592320000000
0!
0%
b0 *
0-
02
b0 6
#592330000000
1!
1%
1-
12
#592340000000
0!
0%
b1 *
0-
02
b1 6
#592350000000
1!
1%
1-
12
#592360000000
0!
0%
b10 *
0-
02
b10 6
#592370000000
1!
1%
1-
12
#592380000000
0!
0%
b11 *
0-
02
b11 6
#592390000000
1!
1%
1-
12
15
#592400000000
0!
0%
b100 *
0-
02
b100 6
#592410000000
1!
1%
1-
12
#592420000000
0!
0%
b101 *
0-
02
b101 6
#592430000000
1!
1%
1-
12
#592440000000
0!
0%
b110 *
0-
02
b110 6
#592450000000
1!
1%
1-
12
#592460000000
0!
0%
b111 *
0-
02
b111 6
#592470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#592480000000
0!
0%
b0 *
0-
02
b0 6
#592490000000
1!
1%
1-
12
#592500000000
0!
0%
b1 *
0-
02
b1 6
#592510000000
1!
1%
1-
12
#592520000000
0!
0%
b10 *
0-
02
b10 6
#592530000000
1!
1%
1-
12
#592540000000
0!
0%
b11 *
0-
02
b11 6
#592550000000
1!
1%
1-
12
15
#592560000000
0!
0%
b100 *
0-
02
b100 6
#592570000000
1!
1%
1-
12
#592580000000
0!
0%
b101 *
0-
02
b101 6
#592590000000
1!
1%
1-
12
#592600000000
0!
0%
b110 *
0-
02
b110 6
#592610000000
1!
1%
1-
12
#592620000000
0!
0%
b111 *
0-
02
b111 6
#592630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#592640000000
0!
0%
b0 *
0-
02
b0 6
#592650000000
1!
1%
1-
12
#592660000000
0!
0%
b1 *
0-
02
b1 6
#592670000000
1!
1%
1-
12
#592680000000
0!
0%
b10 *
0-
02
b10 6
#592690000000
1!
1%
1-
12
#592700000000
0!
0%
b11 *
0-
02
b11 6
#592710000000
1!
1%
1-
12
15
#592720000000
0!
0%
b100 *
0-
02
b100 6
#592730000000
1!
1%
1-
12
#592740000000
0!
0%
b101 *
0-
02
b101 6
#592750000000
1!
1%
1-
12
#592760000000
0!
0%
b110 *
0-
02
b110 6
#592770000000
1!
1%
1-
12
#592780000000
0!
0%
b111 *
0-
02
b111 6
#592790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#592800000000
0!
0%
b0 *
0-
02
b0 6
#592810000000
1!
1%
1-
12
#592820000000
0!
0%
b1 *
0-
02
b1 6
#592830000000
1!
1%
1-
12
#592840000000
0!
0%
b10 *
0-
02
b10 6
#592850000000
1!
1%
1-
12
#592860000000
0!
0%
b11 *
0-
02
b11 6
#592870000000
1!
1%
1-
12
15
#592880000000
0!
0%
b100 *
0-
02
b100 6
#592890000000
1!
1%
1-
12
#592900000000
0!
0%
b101 *
0-
02
b101 6
#592910000000
1!
1%
1-
12
#592920000000
0!
0%
b110 *
0-
02
b110 6
#592930000000
1!
1%
1-
12
#592940000000
0!
0%
b111 *
0-
02
b111 6
#592950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#592960000000
0!
0%
b0 *
0-
02
b0 6
#592970000000
1!
1%
1-
12
#592980000000
0!
0%
b1 *
0-
02
b1 6
#592990000000
1!
1%
1-
12
#593000000000
0!
0%
b10 *
0-
02
b10 6
#593010000000
1!
1%
1-
12
#593020000000
0!
0%
b11 *
0-
02
b11 6
#593030000000
1!
1%
1-
12
15
#593040000000
0!
0%
b100 *
0-
02
b100 6
#593050000000
1!
1%
1-
12
#593060000000
0!
0%
b101 *
0-
02
b101 6
#593070000000
1!
1%
1-
12
#593080000000
0!
0%
b110 *
0-
02
b110 6
#593090000000
1!
1%
1-
12
#593100000000
0!
0%
b111 *
0-
02
b111 6
#593110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#593120000000
0!
0%
b0 *
0-
02
b0 6
#593130000000
1!
1%
1-
12
#593140000000
0!
0%
b1 *
0-
02
b1 6
#593150000000
1!
1%
1-
12
#593160000000
0!
0%
b10 *
0-
02
b10 6
#593170000000
1!
1%
1-
12
#593180000000
0!
0%
b11 *
0-
02
b11 6
#593190000000
1!
1%
1-
12
15
#593200000000
0!
0%
b100 *
0-
02
b100 6
#593210000000
1!
1%
1-
12
#593220000000
0!
0%
b101 *
0-
02
b101 6
#593230000000
1!
1%
1-
12
#593240000000
0!
0%
b110 *
0-
02
b110 6
#593250000000
1!
1%
1-
12
#593260000000
0!
0%
b111 *
0-
02
b111 6
#593270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#593280000000
0!
0%
b0 *
0-
02
b0 6
#593290000000
1!
1%
1-
12
#593300000000
0!
0%
b1 *
0-
02
b1 6
#593310000000
1!
1%
1-
12
#593320000000
0!
0%
b10 *
0-
02
b10 6
#593330000000
1!
1%
1-
12
#593340000000
0!
0%
b11 *
0-
02
b11 6
#593350000000
1!
1%
1-
12
15
#593360000000
0!
0%
b100 *
0-
02
b100 6
#593370000000
1!
1%
1-
12
#593380000000
0!
0%
b101 *
0-
02
b101 6
#593390000000
1!
1%
1-
12
#593400000000
0!
0%
b110 *
0-
02
b110 6
#593410000000
1!
1%
1-
12
#593420000000
0!
0%
b111 *
0-
02
b111 6
#593430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#593440000000
0!
0%
b0 *
0-
02
b0 6
#593450000000
1!
1%
1-
12
#593460000000
0!
0%
b1 *
0-
02
b1 6
#593470000000
1!
1%
1-
12
#593480000000
0!
0%
b10 *
0-
02
b10 6
#593490000000
1!
1%
1-
12
#593500000000
0!
0%
b11 *
0-
02
b11 6
#593510000000
1!
1%
1-
12
15
#593520000000
0!
0%
b100 *
0-
02
b100 6
#593530000000
1!
1%
1-
12
#593540000000
0!
0%
b101 *
0-
02
b101 6
#593550000000
1!
1%
1-
12
#593560000000
0!
0%
b110 *
0-
02
b110 6
#593570000000
1!
1%
1-
12
#593580000000
0!
0%
b111 *
0-
02
b111 6
#593590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#593600000000
0!
0%
b0 *
0-
02
b0 6
#593610000000
1!
1%
1-
12
#593620000000
0!
0%
b1 *
0-
02
b1 6
#593630000000
1!
1%
1-
12
#593640000000
0!
0%
b10 *
0-
02
b10 6
#593650000000
1!
1%
1-
12
#593660000000
0!
0%
b11 *
0-
02
b11 6
#593670000000
1!
1%
1-
12
15
#593680000000
0!
0%
b100 *
0-
02
b100 6
#593690000000
1!
1%
1-
12
#593700000000
0!
0%
b101 *
0-
02
b101 6
#593710000000
1!
1%
1-
12
#593720000000
0!
0%
b110 *
0-
02
b110 6
#593730000000
1!
1%
1-
12
#593740000000
0!
0%
b111 *
0-
02
b111 6
#593750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#593760000000
0!
0%
b0 *
0-
02
b0 6
#593770000000
1!
1%
1-
12
#593780000000
0!
0%
b1 *
0-
02
b1 6
#593790000000
1!
1%
1-
12
#593800000000
0!
0%
b10 *
0-
02
b10 6
#593810000000
1!
1%
1-
12
#593820000000
0!
0%
b11 *
0-
02
b11 6
#593830000000
1!
1%
1-
12
15
#593840000000
0!
0%
b100 *
0-
02
b100 6
#593850000000
1!
1%
1-
12
#593860000000
0!
0%
b101 *
0-
02
b101 6
#593870000000
1!
1%
1-
12
#593880000000
0!
0%
b110 *
0-
02
b110 6
#593890000000
1!
1%
1-
12
#593900000000
0!
0%
b111 *
0-
02
b111 6
#593910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#593920000000
0!
0%
b0 *
0-
02
b0 6
#593930000000
1!
1%
1-
12
#593940000000
0!
0%
b1 *
0-
02
b1 6
#593950000000
1!
1%
1-
12
#593960000000
0!
0%
b10 *
0-
02
b10 6
#593970000000
1!
1%
1-
12
#593980000000
0!
0%
b11 *
0-
02
b11 6
#593990000000
1!
1%
1-
12
15
#594000000000
0!
0%
b100 *
0-
02
b100 6
#594010000000
1!
1%
1-
12
#594020000000
0!
0%
b101 *
0-
02
b101 6
#594030000000
1!
1%
1-
12
#594040000000
0!
0%
b110 *
0-
02
b110 6
#594050000000
1!
1%
1-
12
#594060000000
0!
0%
b111 *
0-
02
b111 6
#594070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#594080000000
0!
0%
b0 *
0-
02
b0 6
#594090000000
1!
1%
1-
12
#594100000000
0!
0%
b1 *
0-
02
b1 6
#594110000000
1!
1%
1-
12
#594120000000
0!
0%
b10 *
0-
02
b10 6
#594130000000
1!
1%
1-
12
#594140000000
0!
0%
b11 *
0-
02
b11 6
#594150000000
1!
1%
1-
12
15
#594160000000
0!
0%
b100 *
0-
02
b100 6
#594170000000
1!
1%
1-
12
#594180000000
0!
0%
b101 *
0-
02
b101 6
#594190000000
1!
1%
1-
12
#594200000000
0!
0%
b110 *
0-
02
b110 6
#594210000000
1!
1%
1-
12
#594220000000
0!
0%
b111 *
0-
02
b111 6
#594230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#594240000000
0!
0%
b0 *
0-
02
b0 6
#594250000000
1!
1%
1-
12
#594260000000
0!
0%
b1 *
0-
02
b1 6
#594270000000
1!
1%
1-
12
#594280000000
0!
0%
b10 *
0-
02
b10 6
#594290000000
1!
1%
1-
12
#594300000000
0!
0%
b11 *
0-
02
b11 6
#594310000000
1!
1%
1-
12
15
#594320000000
0!
0%
b100 *
0-
02
b100 6
#594330000000
1!
1%
1-
12
#594340000000
0!
0%
b101 *
0-
02
b101 6
#594350000000
1!
1%
1-
12
#594360000000
0!
0%
b110 *
0-
02
b110 6
#594370000000
1!
1%
1-
12
#594380000000
0!
0%
b111 *
0-
02
b111 6
#594390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#594400000000
0!
0%
b0 *
0-
02
b0 6
#594410000000
1!
1%
1-
12
#594420000000
0!
0%
b1 *
0-
02
b1 6
#594430000000
1!
1%
1-
12
#594440000000
0!
0%
b10 *
0-
02
b10 6
#594450000000
1!
1%
1-
12
#594460000000
0!
0%
b11 *
0-
02
b11 6
#594470000000
1!
1%
1-
12
15
#594480000000
0!
0%
b100 *
0-
02
b100 6
#594490000000
1!
1%
1-
12
#594500000000
0!
0%
b101 *
0-
02
b101 6
#594510000000
1!
1%
1-
12
#594520000000
0!
0%
b110 *
0-
02
b110 6
#594530000000
1!
1%
1-
12
#594540000000
0!
0%
b111 *
0-
02
b111 6
#594550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#594560000000
0!
0%
b0 *
0-
02
b0 6
#594570000000
1!
1%
1-
12
#594580000000
0!
0%
b1 *
0-
02
b1 6
#594590000000
1!
1%
1-
12
#594600000000
0!
0%
b10 *
0-
02
b10 6
#594610000000
1!
1%
1-
12
#594620000000
0!
0%
b11 *
0-
02
b11 6
#594630000000
1!
1%
1-
12
15
#594640000000
0!
0%
b100 *
0-
02
b100 6
#594650000000
1!
1%
1-
12
#594660000000
0!
0%
b101 *
0-
02
b101 6
#594670000000
1!
1%
1-
12
#594680000000
0!
0%
b110 *
0-
02
b110 6
#594690000000
1!
1%
1-
12
#594700000000
0!
0%
b111 *
0-
02
b111 6
#594710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#594720000000
0!
0%
b0 *
0-
02
b0 6
#594730000000
1!
1%
1-
12
#594740000000
0!
0%
b1 *
0-
02
b1 6
#594750000000
1!
1%
1-
12
#594760000000
0!
0%
b10 *
0-
02
b10 6
#594770000000
1!
1%
1-
12
#594780000000
0!
0%
b11 *
0-
02
b11 6
#594790000000
1!
1%
1-
12
15
#594800000000
0!
0%
b100 *
0-
02
b100 6
#594810000000
1!
1%
1-
12
#594820000000
0!
0%
b101 *
0-
02
b101 6
#594830000000
1!
1%
1-
12
#594840000000
0!
0%
b110 *
0-
02
b110 6
#594850000000
1!
1%
1-
12
#594860000000
0!
0%
b111 *
0-
02
b111 6
#594870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#594880000000
0!
0%
b0 *
0-
02
b0 6
#594890000000
1!
1%
1-
12
#594900000000
0!
0%
b1 *
0-
02
b1 6
#594910000000
1!
1%
1-
12
#594920000000
0!
0%
b10 *
0-
02
b10 6
#594930000000
1!
1%
1-
12
#594940000000
0!
0%
b11 *
0-
02
b11 6
#594950000000
1!
1%
1-
12
15
#594960000000
0!
0%
b100 *
0-
02
b100 6
#594970000000
1!
1%
1-
12
#594980000000
0!
0%
b101 *
0-
02
b101 6
#594990000000
1!
1%
1-
12
#595000000000
0!
0%
b110 *
0-
02
b110 6
#595010000000
1!
1%
1-
12
#595020000000
0!
0%
b111 *
0-
02
b111 6
#595030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#595040000000
0!
0%
b0 *
0-
02
b0 6
#595050000000
1!
1%
1-
12
#595060000000
0!
0%
b1 *
0-
02
b1 6
#595070000000
1!
1%
1-
12
#595080000000
0!
0%
b10 *
0-
02
b10 6
#595090000000
1!
1%
1-
12
#595100000000
0!
0%
b11 *
0-
02
b11 6
#595110000000
1!
1%
1-
12
15
#595120000000
0!
0%
b100 *
0-
02
b100 6
#595130000000
1!
1%
1-
12
#595140000000
0!
0%
b101 *
0-
02
b101 6
#595150000000
1!
1%
1-
12
#595160000000
0!
0%
b110 *
0-
02
b110 6
#595170000000
1!
1%
1-
12
#595180000000
0!
0%
b111 *
0-
02
b111 6
#595190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#595200000000
0!
0%
b0 *
0-
02
b0 6
#595210000000
1!
1%
1-
12
#595220000000
0!
0%
b1 *
0-
02
b1 6
#595230000000
1!
1%
1-
12
#595240000000
0!
0%
b10 *
0-
02
b10 6
#595250000000
1!
1%
1-
12
#595260000000
0!
0%
b11 *
0-
02
b11 6
#595270000000
1!
1%
1-
12
15
#595280000000
0!
0%
b100 *
0-
02
b100 6
#595290000000
1!
1%
1-
12
#595300000000
0!
0%
b101 *
0-
02
b101 6
#595310000000
1!
1%
1-
12
#595320000000
0!
0%
b110 *
0-
02
b110 6
#595330000000
1!
1%
1-
12
#595340000000
0!
0%
b111 *
0-
02
b111 6
#595350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#595360000000
0!
0%
b0 *
0-
02
b0 6
#595370000000
1!
1%
1-
12
#595380000000
0!
0%
b1 *
0-
02
b1 6
#595390000000
1!
1%
1-
12
#595400000000
0!
0%
b10 *
0-
02
b10 6
#595410000000
1!
1%
1-
12
#595420000000
0!
0%
b11 *
0-
02
b11 6
#595430000000
1!
1%
1-
12
15
#595440000000
0!
0%
b100 *
0-
02
b100 6
#595450000000
1!
1%
1-
12
#595460000000
0!
0%
b101 *
0-
02
b101 6
#595470000000
1!
1%
1-
12
#595480000000
0!
0%
b110 *
0-
02
b110 6
#595490000000
1!
1%
1-
12
#595500000000
0!
0%
b111 *
0-
02
b111 6
#595510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#595520000000
0!
0%
b0 *
0-
02
b0 6
#595530000000
1!
1%
1-
12
#595540000000
0!
0%
b1 *
0-
02
b1 6
#595550000000
1!
1%
1-
12
#595560000000
0!
0%
b10 *
0-
02
b10 6
#595570000000
1!
1%
1-
12
#595580000000
0!
0%
b11 *
0-
02
b11 6
#595590000000
1!
1%
1-
12
15
#595600000000
0!
0%
b100 *
0-
02
b100 6
#595610000000
1!
1%
1-
12
#595620000000
0!
0%
b101 *
0-
02
b101 6
#595630000000
1!
1%
1-
12
#595640000000
0!
0%
b110 *
0-
02
b110 6
#595650000000
1!
1%
1-
12
#595660000000
0!
0%
b111 *
0-
02
b111 6
#595670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#595680000000
0!
0%
b0 *
0-
02
b0 6
#595690000000
1!
1%
1-
12
#595700000000
0!
0%
b1 *
0-
02
b1 6
#595710000000
1!
1%
1-
12
#595720000000
0!
0%
b10 *
0-
02
b10 6
#595730000000
1!
1%
1-
12
#595740000000
0!
0%
b11 *
0-
02
b11 6
#595750000000
1!
1%
1-
12
15
#595760000000
0!
0%
b100 *
0-
02
b100 6
#595770000000
1!
1%
1-
12
#595780000000
0!
0%
b101 *
0-
02
b101 6
#595790000000
1!
1%
1-
12
#595800000000
0!
0%
b110 *
0-
02
b110 6
#595810000000
1!
1%
1-
12
#595820000000
0!
0%
b111 *
0-
02
b111 6
#595830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#595840000000
0!
0%
b0 *
0-
02
b0 6
#595850000000
1!
1%
1-
12
#595860000000
0!
0%
b1 *
0-
02
b1 6
#595870000000
1!
1%
1-
12
#595880000000
0!
0%
b10 *
0-
02
b10 6
#595890000000
1!
1%
1-
12
#595900000000
0!
0%
b11 *
0-
02
b11 6
#595910000000
1!
1%
1-
12
15
#595920000000
0!
0%
b100 *
0-
02
b100 6
#595930000000
1!
1%
1-
12
#595940000000
0!
0%
b101 *
0-
02
b101 6
#595950000000
1!
1%
1-
12
#595960000000
0!
0%
b110 *
0-
02
b110 6
#595970000000
1!
1%
1-
12
#595980000000
0!
0%
b111 *
0-
02
b111 6
#595990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#596000000000
0!
0%
b0 *
0-
02
b0 6
#596010000000
1!
1%
1-
12
#596020000000
0!
0%
b1 *
0-
02
b1 6
#596030000000
1!
1%
1-
12
#596040000000
0!
0%
b10 *
0-
02
b10 6
#596050000000
1!
1%
1-
12
#596060000000
0!
0%
b11 *
0-
02
b11 6
#596070000000
1!
1%
1-
12
15
#596080000000
0!
0%
b100 *
0-
02
b100 6
#596090000000
1!
1%
1-
12
#596100000000
0!
0%
b101 *
0-
02
b101 6
#596110000000
1!
1%
1-
12
#596120000000
0!
0%
b110 *
0-
02
b110 6
#596130000000
1!
1%
1-
12
#596140000000
0!
0%
b111 *
0-
02
b111 6
#596150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#596160000000
0!
0%
b0 *
0-
02
b0 6
#596170000000
1!
1%
1-
12
#596180000000
0!
0%
b1 *
0-
02
b1 6
#596190000000
1!
1%
1-
12
#596200000000
0!
0%
b10 *
0-
02
b10 6
#596210000000
1!
1%
1-
12
#596220000000
0!
0%
b11 *
0-
02
b11 6
#596230000000
1!
1%
1-
12
15
#596240000000
0!
0%
b100 *
0-
02
b100 6
#596250000000
1!
1%
1-
12
#596260000000
0!
0%
b101 *
0-
02
b101 6
#596270000000
1!
1%
1-
12
#596280000000
0!
0%
b110 *
0-
02
b110 6
#596290000000
1!
1%
1-
12
#596300000000
0!
0%
b111 *
0-
02
b111 6
#596310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#596320000000
0!
0%
b0 *
0-
02
b0 6
#596330000000
1!
1%
1-
12
#596340000000
0!
0%
b1 *
0-
02
b1 6
#596350000000
1!
1%
1-
12
#596360000000
0!
0%
b10 *
0-
02
b10 6
#596370000000
1!
1%
1-
12
#596380000000
0!
0%
b11 *
0-
02
b11 6
#596390000000
1!
1%
1-
12
15
#596400000000
0!
0%
b100 *
0-
02
b100 6
#596410000000
1!
1%
1-
12
#596420000000
0!
0%
b101 *
0-
02
b101 6
#596430000000
1!
1%
1-
12
#596440000000
0!
0%
b110 *
0-
02
b110 6
#596450000000
1!
1%
1-
12
#596460000000
0!
0%
b111 *
0-
02
b111 6
#596470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#596480000000
0!
0%
b0 *
0-
02
b0 6
#596490000000
1!
1%
1-
12
#596500000000
0!
0%
b1 *
0-
02
b1 6
#596510000000
1!
1%
1-
12
#596520000000
0!
0%
b10 *
0-
02
b10 6
#596530000000
1!
1%
1-
12
#596540000000
0!
0%
b11 *
0-
02
b11 6
#596550000000
1!
1%
1-
12
15
#596560000000
0!
0%
b100 *
0-
02
b100 6
#596570000000
1!
1%
1-
12
#596580000000
0!
0%
b101 *
0-
02
b101 6
#596590000000
1!
1%
1-
12
#596600000000
0!
0%
b110 *
0-
02
b110 6
#596610000000
1!
1%
1-
12
#596620000000
0!
0%
b111 *
0-
02
b111 6
#596630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#596640000000
0!
0%
b0 *
0-
02
b0 6
#596650000000
1!
1%
1-
12
#596660000000
0!
0%
b1 *
0-
02
b1 6
#596670000000
1!
1%
1-
12
#596680000000
0!
0%
b10 *
0-
02
b10 6
#596690000000
1!
1%
1-
12
#596700000000
0!
0%
b11 *
0-
02
b11 6
#596710000000
1!
1%
1-
12
15
#596720000000
0!
0%
b100 *
0-
02
b100 6
#596730000000
1!
1%
1-
12
#596740000000
0!
0%
b101 *
0-
02
b101 6
#596750000000
1!
1%
1-
12
#596760000000
0!
0%
b110 *
0-
02
b110 6
#596770000000
1!
1%
1-
12
#596780000000
0!
0%
b111 *
0-
02
b111 6
#596790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#596800000000
0!
0%
b0 *
0-
02
b0 6
#596810000000
1!
1%
1-
12
#596820000000
0!
0%
b1 *
0-
02
b1 6
#596830000000
1!
1%
1-
12
#596840000000
0!
0%
b10 *
0-
02
b10 6
#596850000000
1!
1%
1-
12
#596860000000
0!
0%
b11 *
0-
02
b11 6
#596870000000
1!
1%
1-
12
15
#596880000000
0!
0%
b100 *
0-
02
b100 6
#596890000000
1!
1%
1-
12
#596900000000
0!
0%
b101 *
0-
02
b101 6
#596910000000
1!
1%
1-
12
#596920000000
0!
0%
b110 *
0-
02
b110 6
#596930000000
1!
1%
1-
12
#596940000000
0!
0%
b111 *
0-
02
b111 6
#596950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#596960000000
0!
0%
b0 *
0-
02
b0 6
#596970000000
1!
1%
1-
12
#596980000000
0!
0%
b1 *
0-
02
b1 6
#596990000000
1!
1%
1-
12
#597000000000
0!
0%
b10 *
0-
02
b10 6
#597010000000
1!
1%
1-
12
#597020000000
0!
0%
b11 *
0-
02
b11 6
#597030000000
1!
1%
1-
12
15
#597040000000
0!
0%
b100 *
0-
02
b100 6
#597050000000
1!
1%
1-
12
#597060000000
0!
0%
b101 *
0-
02
b101 6
#597070000000
1!
1%
1-
12
#597080000000
0!
0%
b110 *
0-
02
b110 6
#597090000000
1!
1%
1-
12
#597100000000
0!
0%
b111 *
0-
02
b111 6
#597110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#597120000000
0!
0%
b0 *
0-
02
b0 6
#597130000000
1!
1%
1-
12
#597140000000
0!
0%
b1 *
0-
02
b1 6
#597150000000
1!
1%
1-
12
#597160000000
0!
0%
b10 *
0-
02
b10 6
#597170000000
1!
1%
1-
12
#597180000000
0!
0%
b11 *
0-
02
b11 6
#597190000000
1!
1%
1-
12
15
#597200000000
0!
0%
b100 *
0-
02
b100 6
#597210000000
1!
1%
1-
12
#597220000000
0!
0%
b101 *
0-
02
b101 6
#597230000000
1!
1%
1-
12
#597240000000
0!
0%
b110 *
0-
02
b110 6
#597250000000
1!
1%
1-
12
#597260000000
0!
0%
b111 *
0-
02
b111 6
#597270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#597280000000
0!
0%
b0 *
0-
02
b0 6
#597290000000
1!
1%
1-
12
#597300000000
0!
0%
b1 *
0-
02
b1 6
#597310000000
1!
1%
1-
12
#597320000000
0!
0%
b10 *
0-
02
b10 6
#597330000000
1!
1%
1-
12
#597340000000
0!
0%
b11 *
0-
02
b11 6
#597350000000
1!
1%
1-
12
15
#597360000000
0!
0%
b100 *
0-
02
b100 6
#597370000000
1!
1%
1-
12
#597380000000
0!
0%
b101 *
0-
02
b101 6
#597390000000
1!
1%
1-
12
#597400000000
0!
0%
b110 *
0-
02
b110 6
#597410000000
1!
1%
1-
12
#597420000000
0!
0%
b111 *
0-
02
b111 6
#597430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#597440000000
0!
0%
b0 *
0-
02
b0 6
#597450000000
1!
1%
1-
12
#597460000000
0!
0%
b1 *
0-
02
b1 6
#597470000000
1!
1%
1-
12
#597480000000
0!
0%
b10 *
0-
02
b10 6
#597490000000
1!
1%
1-
12
#597500000000
0!
0%
b11 *
0-
02
b11 6
#597510000000
1!
1%
1-
12
15
#597520000000
0!
0%
b100 *
0-
02
b100 6
#597530000000
1!
1%
1-
12
#597540000000
0!
0%
b101 *
0-
02
b101 6
#597550000000
1!
1%
1-
12
#597560000000
0!
0%
b110 *
0-
02
b110 6
#597570000000
1!
1%
1-
12
#597580000000
0!
0%
b111 *
0-
02
b111 6
#597590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#597600000000
0!
0%
b0 *
0-
02
b0 6
#597610000000
1!
1%
1-
12
#597620000000
0!
0%
b1 *
0-
02
b1 6
#597630000000
1!
1%
1-
12
#597640000000
0!
0%
b10 *
0-
02
b10 6
#597650000000
1!
1%
1-
12
#597660000000
0!
0%
b11 *
0-
02
b11 6
#597670000000
1!
1%
1-
12
15
#597680000000
0!
0%
b100 *
0-
02
b100 6
#597690000000
1!
1%
1-
12
#597700000000
0!
0%
b101 *
0-
02
b101 6
#597710000000
1!
1%
1-
12
#597720000000
0!
0%
b110 *
0-
02
b110 6
#597730000000
1!
1%
1-
12
#597740000000
0!
0%
b111 *
0-
02
b111 6
#597750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#597760000000
0!
0%
b0 *
0-
02
b0 6
#597770000000
1!
1%
1-
12
#597780000000
0!
0%
b1 *
0-
02
b1 6
#597790000000
1!
1%
1-
12
#597800000000
0!
0%
b10 *
0-
02
b10 6
#597810000000
1!
1%
1-
12
#597820000000
0!
0%
b11 *
0-
02
b11 6
#597830000000
1!
1%
1-
12
15
#597840000000
0!
0%
b100 *
0-
02
b100 6
#597850000000
1!
1%
1-
12
#597860000000
0!
0%
b101 *
0-
02
b101 6
#597870000000
1!
1%
1-
12
#597880000000
0!
0%
b110 *
0-
02
b110 6
#597890000000
1!
1%
1-
12
#597900000000
0!
0%
b111 *
0-
02
b111 6
#597910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#597920000000
0!
0%
b0 *
0-
02
b0 6
#597930000000
1!
1%
1-
12
#597940000000
0!
0%
b1 *
0-
02
b1 6
#597950000000
1!
1%
1-
12
#597960000000
0!
0%
b10 *
0-
02
b10 6
#597970000000
1!
1%
1-
12
#597980000000
0!
0%
b11 *
0-
02
b11 6
#597990000000
1!
1%
1-
12
15
#598000000000
0!
0%
b100 *
0-
02
b100 6
#598010000000
1!
1%
1-
12
#598020000000
0!
0%
b101 *
0-
02
b101 6
#598030000000
1!
1%
1-
12
#598040000000
0!
0%
b110 *
0-
02
b110 6
#598050000000
1!
1%
1-
12
#598060000000
0!
0%
b111 *
0-
02
b111 6
#598070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#598080000000
0!
0%
b0 *
0-
02
b0 6
#598090000000
1!
1%
1-
12
#598100000000
0!
0%
b1 *
0-
02
b1 6
#598110000000
1!
1%
1-
12
#598120000000
0!
0%
b10 *
0-
02
b10 6
#598130000000
1!
1%
1-
12
#598140000000
0!
0%
b11 *
0-
02
b11 6
#598150000000
1!
1%
1-
12
15
#598160000000
0!
0%
b100 *
0-
02
b100 6
#598170000000
1!
1%
1-
12
#598180000000
0!
0%
b101 *
0-
02
b101 6
#598190000000
1!
1%
1-
12
#598200000000
0!
0%
b110 *
0-
02
b110 6
#598210000000
1!
1%
1-
12
#598220000000
0!
0%
b111 *
0-
02
b111 6
#598230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#598240000000
0!
0%
b0 *
0-
02
b0 6
#598250000000
1!
1%
1-
12
#598260000000
0!
0%
b1 *
0-
02
b1 6
#598270000000
1!
1%
1-
12
#598280000000
0!
0%
b10 *
0-
02
b10 6
#598290000000
1!
1%
1-
12
#598300000000
0!
0%
b11 *
0-
02
b11 6
#598310000000
1!
1%
1-
12
15
#598320000000
0!
0%
b100 *
0-
02
b100 6
#598330000000
1!
1%
1-
12
#598340000000
0!
0%
b101 *
0-
02
b101 6
#598350000000
1!
1%
1-
12
#598360000000
0!
0%
b110 *
0-
02
b110 6
#598370000000
1!
1%
1-
12
#598380000000
0!
0%
b111 *
0-
02
b111 6
#598390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#598400000000
0!
0%
b0 *
0-
02
b0 6
#598410000000
1!
1%
1-
12
#598420000000
0!
0%
b1 *
0-
02
b1 6
#598430000000
1!
1%
1-
12
#598440000000
0!
0%
b10 *
0-
02
b10 6
#598450000000
1!
1%
1-
12
#598460000000
0!
0%
b11 *
0-
02
b11 6
#598470000000
1!
1%
1-
12
15
#598480000000
0!
0%
b100 *
0-
02
b100 6
#598490000000
1!
1%
1-
12
#598500000000
0!
0%
b101 *
0-
02
b101 6
#598510000000
1!
1%
1-
12
#598520000000
0!
0%
b110 *
0-
02
b110 6
#598530000000
1!
1%
1-
12
#598540000000
0!
0%
b111 *
0-
02
b111 6
#598550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#598560000000
0!
0%
b0 *
0-
02
b0 6
#598570000000
1!
1%
1-
12
#598580000000
0!
0%
b1 *
0-
02
b1 6
#598590000000
1!
1%
1-
12
#598600000000
0!
0%
b10 *
0-
02
b10 6
#598610000000
1!
1%
1-
12
#598620000000
0!
0%
b11 *
0-
02
b11 6
#598630000000
1!
1%
1-
12
15
#598640000000
0!
0%
b100 *
0-
02
b100 6
#598650000000
1!
1%
1-
12
#598660000000
0!
0%
b101 *
0-
02
b101 6
#598670000000
1!
1%
1-
12
#598680000000
0!
0%
b110 *
0-
02
b110 6
#598690000000
1!
1%
1-
12
#598700000000
0!
0%
b111 *
0-
02
b111 6
#598710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#598720000000
0!
0%
b0 *
0-
02
b0 6
#598730000000
1!
1%
1-
12
#598740000000
0!
0%
b1 *
0-
02
b1 6
#598750000000
1!
1%
1-
12
#598760000000
0!
0%
b10 *
0-
02
b10 6
#598770000000
1!
1%
1-
12
#598780000000
0!
0%
b11 *
0-
02
b11 6
#598790000000
1!
1%
1-
12
15
#598800000000
0!
0%
b100 *
0-
02
b100 6
#598810000000
1!
1%
1-
12
#598820000000
0!
0%
b101 *
0-
02
b101 6
#598830000000
1!
1%
1-
12
#598840000000
0!
0%
b110 *
0-
02
b110 6
#598850000000
1!
1%
1-
12
#598860000000
0!
0%
b111 *
0-
02
b111 6
#598870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#598880000000
0!
0%
b0 *
0-
02
b0 6
#598890000000
1!
1%
1-
12
#598900000000
0!
0%
b1 *
0-
02
b1 6
#598910000000
1!
1%
1-
12
#598920000000
0!
0%
b10 *
0-
02
b10 6
#598930000000
1!
1%
1-
12
#598940000000
0!
0%
b11 *
0-
02
b11 6
#598950000000
1!
1%
1-
12
15
#598960000000
0!
0%
b100 *
0-
02
b100 6
#598970000000
1!
1%
1-
12
#598980000000
0!
0%
b101 *
0-
02
b101 6
#598990000000
1!
1%
1-
12
#599000000000
0!
0%
b110 *
0-
02
b110 6
#599010000000
1!
1%
1-
12
#599020000000
0!
0%
b111 *
0-
02
b111 6
#599030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#599040000000
0!
0%
b0 *
0-
02
b0 6
#599050000000
1!
1%
1-
12
#599060000000
0!
0%
b1 *
0-
02
b1 6
#599070000000
1!
1%
1-
12
#599080000000
0!
0%
b10 *
0-
02
b10 6
#599090000000
1!
1%
1-
12
#599100000000
0!
0%
b11 *
0-
02
b11 6
#599110000000
1!
1%
1-
12
15
#599120000000
0!
0%
b100 *
0-
02
b100 6
#599130000000
1!
1%
1-
12
#599140000000
0!
0%
b101 *
0-
02
b101 6
#599150000000
1!
1%
1-
12
#599160000000
0!
0%
b110 *
0-
02
b110 6
#599170000000
1!
1%
1-
12
#599180000000
0!
0%
b111 *
0-
02
b111 6
#599190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#599200000000
0!
0%
b0 *
0-
02
b0 6
#599210000000
1!
1%
1-
12
#599220000000
0!
0%
b1 *
0-
02
b1 6
#599230000000
1!
1%
1-
12
#599240000000
0!
0%
b10 *
0-
02
b10 6
#599250000000
1!
1%
1-
12
#599260000000
0!
0%
b11 *
0-
02
b11 6
#599270000000
1!
1%
1-
12
15
#599280000000
0!
0%
b100 *
0-
02
b100 6
#599290000000
1!
1%
1-
12
#599300000000
0!
0%
b101 *
0-
02
b101 6
#599310000000
1!
1%
1-
12
#599320000000
0!
0%
b110 *
0-
02
b110 6
#599330000000
1!
1%
1-
12
#599340000000
0!
0%
b111 *
0-
02
b111 6
#599350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#599360000000
0!
0%
b0 *
0-
02
b0 6
#599370000000
1!
1%
1-
12
#599380000000
0!
0%
b1 *
0-
02
b1 6
#599390000000
1!
1%
1-
12
#599400000000
0!
0%
b10 *
0-
02
b10 6
#599410000000
1!
1%
1-
12
#599420000000
0!
0%
b11 *
0-
02
b11 6
#599430000000
1!
1%
1-
12
15
#599440000000
0!
0%
b100 *
0-
02
b100 6
#599450000000
1!
1%
1-
12
#599460000000
0!
0%
b101 *
0-
02
b101 6
#599470000000
1!
1%
1-
12
#599480000000
0!
0%
b110 *
0-
02
b110 6
#599490000000
1!
1%
1-
12
#599500000000
0!
0%
b111 *
0-
02
b111 6
#599510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#599520000000
0!
0%
b0 *
0-
02
b0 6
#599530000000
1!
1%
1-
12
#599540000000
0!
0%
b1 *
0-
02
b1 6
#599550000000
1!
1%
1-
12
#599560000000
0!
0%
b10 *
0-
02
b10 6
#599570000000
1!
1%
1-
12
#599580000000
0!
0%
b11 *
0-
02
b11 6
#599590000000
1!
1%
1-
12
15
#599600000000
0!
0%
b100 *
0-
02
b100 6
#599610000000
1!
1%
1-
12
#599620000000
0!
0%
b101 *
0-
02
b101 6
#599630000000
1!
1%
1-
12
#599640000000
0!
0%
b110 *
0-
02
b110 6
#599650000000
1!
1%
1-
12
#599660000000
0!
0%
b111 *
0-
02
b111 6
#599670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#599680000000
0!
0%
b0 *
0-
02
b0 6
#599690000000
1!
1%
1-
12
#599700000000
0!
0%
b1 *
0-
02
b1 6
#599710000000
1!
1%
1-
12
#599720000000
0!
0%
b10 *
0-
02
b10 6
#599730000000
1!
1%
1-
12
#599740000000
0!
0%
b11 *
0-
02
b11 6
#599750000000
1!
1%
1-
12
15
#599760000000
0!
0%
b100 *
0-
02
b100 6
#599770000000
1!
1%
1-
12
#599780000000
0!
0%
b101 *
0-
02
b101 6
#599790000000
1!
1%
1-
12
#599800000000
0!
0%
b110 *
0-
02
b110 6
#599810000000
1!
1%
1-
12
#599820000000
0!
0%
b111 *
0-
02
b111 6
#599830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#599840000000
0!
0%
b0 *
0-
02
b0 6
#599850000000
1!
1%
1-
12
#599860000000
0!
0%
b1 *
0-
02
b1 6
#599870000000
1!
1%
1-
12
#599880000000
0!
0%
b10 *
0-
02
b10 6
#599890000000
1!
1%
1-
12
#599900000000
0!
0%
b11 *
0-
02
b11 6
#599910000000
1!
1%
1-
12
15
#599920000000
0!
0%
b100 *
0-
02
b100 6
#599930000000
1!
1%
1-
12
#599940000000
0!
0%
b101 *
0-
02
b101 6
#599950000000
1!
1%
1-
12
#599960000000
0!
0%
b110 *
0-
02
b110 6
#599970000000
1!
1%
1-
12
#599980000000
0!
0%
b111 *
0-
02
b111 6
#599990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#600000000000
0!
0%
b0 *
0-
02
b0 6
#600010000000
1!
1%
1-
12
#600020000000
0!
0%
b1 *
0-
02
b1 6
#600030000000
1!
1%
1-
12
#600040000000
0!
0%
b10 *
0-
02
b10 6
#600050000000
1!
1%
1-
12
#600060000000
0!
0%
b11 *
0-
02
b11 6
#600070000000
1!
1%
1-
12
15
#600080000000
0!
0%
b100 *
0-
02
b100 6
#600090000000
1!
1%
1-
12
#600100000000
0!
0%
b101 *
0-
02
b101 6
#600110000000
1!
1%
1-
12
#600120000000
0!
0%
b110 *
0-
02
b110 6
#600130000000
1!
1%
1-
12
#600140000000
0!
0%
b111 *
0-
02
b111 6
#600150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#600160000000
0!
0%
b0 *
0-
02
b0 6
#600170000000
1!
1%
1-
12
#600180000000
0!
0%
b1 *
0-
02
b1 6
#600190000000
1!
1%
1-
12
#600200000000
0!
0%
b10 *
0-
02
b10 6
#600210000000
1!
1%
1-
12
#600220000000
0!
0%
b11 *
0-
02
b11 6
#600230000000
1!
1%
1-
12
15
#600240000000
0!
0%
b100 *
0-
02
b100 6
#600250000000
1!
1%
1-
12
#600260000000
0!
0%
b101 *
0-
02
b101 6
#600270000000
1!
1%
1-
12
#600280000000
0!
0%
b110 *
0-
02
b110 6
#600290000000
1!
1%
1-
12
#600300000000
0!
0%
b111 *
0-
02
b111 6
#600310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#600320000000
0!
0%
b0 *
0-
02
b0 6
#600330000000
1!
1%
1-
12
#600340000000
0!
0%
b1 *
0-
02
b1 6
#600350000000
1!
1%
1-
12
#600360000000
0!
0%
b10 *
0-
02
b10 6
#600370000000
1!
1%
1-
12
#600380000000
0!
0%
b11 *
0-
02
b11 6
#600390000000
1!
1%
1-
12
15
#600400000000
0!
0%
b100 *
0-
02
b100 6
#600410000000
1!
1%
1-
12
#600420000000
0!
0%
b101 *
0-
02
b101 6
#600430000000
1!
1%
1-
12
#600440000000
0!
0%
b110 *
0-
02
b110 6
#600450000000
1!
1%
1-
12
#600460000000
0!
0%
b111 *
0-
02
b111 6
#600470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#600480000000
0!
0%
b0 *
0-
02
b0 6
#600490000000
1!
1%
1-
12
#600500000000
0!
0%
b1 *
0-
02
b1 6
#600510000000
1!
1%
1-
12
#600520000000
0!
0%
b10 *
0-
02
b10 6
#600530000000
1!
1%
1-
12
#600540000000
0!
0%
b11 *
0-
02
b11 6
#600550000000
1!
1%
1-
12
15
#600560000000
0!
0%
b100 *
0-
02
b100 6
#600570000000
1!
1%
1-
12
#600580000000
0!
0%
b101 *
0-
02
b101 6
#600590000000
1!
1%
1-
12
#600600000000
0!
0%
b110 *
0-
02
b110 6
#600610000000
1!
1%
1-
12
#600620000000
0!
0%
b111 *
0-
02
b111 6
#600630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#600640000000
0!
0%
b0 *
0-
02
b0 6
#600650000000
1!
1%
1-
12
#600660000000
0!
0%
b1 *
0-
02
b1 6
#600670000000
1!
1%
1-
12
#600680000000
0!
0%
b10 *
0-
02
b10 6
#600690000000
1!
1%
1-
12
#600700000000
0!
0%
b11 *
0-
02
b11 6
#600710000000
1!
1%
1-
12
15
#600720000000
0!
0%
b100 *
0-
02
b100 6
#600730000000
1!
1%
1-
12
#600740000000
0!
0%
b101 *
0-
02
b101 6
#600750000000
1!
1%
1-
12
#600760000000
0!
0%
b110 *
0-
02
b110 6
#600770000000
1!
1%
1-
12
#600780000000
0!
0%
b111 *
0-
02
b111 6
#600790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#600800000000
0!
0%
b0 *
0-
02
b0 6
#600810000000
1!
1%
1-
12
#600820000000
0!
0%
b1 *
0-
02
b1 6
#600830000000
1!
1%
1-
12
#600840000000
0!
0%
b10 *
0-
02
b10 6
#600850000000
1!
1%
1-
12
#600860000000
0!
0%
b11 *
0-
02
b11 6
#600870000000
1!
1%
1-
12
15
#600880000000
0!
0%
b100 *
0-
02
b100 6
#600890000000
1!
1%
1-
12
#600900000000
0!
0%
b101 *
0-
02
b101 6
#600910000000
1!
1%
1-
12
#600920000000
0!
0%
b110 *
0-
02
b110 6
#600930000000
1!
1%
1-
12
#600940000000
0!
0%
b111 *
0-
02
b111 6
#600950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#600960000000
0!
0%
b0 *
0-
02
b0 6
#600970000000
1!
1%
1-
12
#600980000000
0!
0%
b1 *
0-
02
b1 6
#600990000000
1!
1%
1-
12
#601000000000
0!
0%
b10 *
0-
02
b10 6
#601010000000
1!
1%
1-
12
#601020000000
0!
0%
b11 *
0-
02
b11 6
#601030000000
1!
1%
1-
12
15
#601040000000
0!
0%
b100 *
0-
02
b100 6
#601050000000
1!
1%
1-
12
#601060000000
0!
0%
b101 *
0-
02
b101 6
#601070000000
1!
1%
1-
12
#601080000000
0!
0%
b110 *
0-
02
b110 6
#601090000000
1!
1%
1-
12
#601100000000
0!
0%
b111 *
0-
02
b111 6
#601110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#601120000000
0!
0%
b0 *
0-
02
b0 6
#601130000000
1!
1%
1-
12
#601140000000
0!
0%
b1 *
0-
02
b1 6
#601150000000
1!
1%
1-
12
#601160000000
0!
0%
b10 *
0-
02
b10 6
#601170000000
1!
1%
1-
12
#601180000000
0!
0%
b11 *
0-
02
b11 6
#601190000000
1!
1%
1-
12
15
#601200000000
0!
0%
b100 *
0-
02
b100 6
#601210000000
1!
1%
1-
12
#601220000000
0!
0%
b101 *
0-
02
b101 6
#601230000000
1!
1%
1-
12
#601240000000
0!
0%
b110 *
0-
02
b110 6
#601250000000
1!
1%
1-
12
#601260000000
0!
0%
b111 *
0-
02
b111 6
#601270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#601280000000
0!
0%
b0 *
0-
02
b0 6
#601290000000
1!
1%
1-
12
#601300000000
0!
0%
b1 *
0-
02
b1 6
#601310000000
1!
1%
1-
12
#601320000000
0!
0%
b10 *
0-
02
b10 6
#601330000000
1!
1%
1-
12
#601340000000
0!
0%
b11 *
0-
02
b11 6
#601350000000
1!
1%
1-
12
15
#601360000000
0!
0%
b100 *
0-
02
b100 6
#601370000000
1!
1%
1-
12
#601380000000
0!
0%
b101 *
0-
02
b101 6
#601390000000
1!
1%
1-
12
#601400000000
0!
0%
b110 *
0-
02
b110 6
#601410000000
1!
1%
1-
12
#601420000000
0!
0%
b111 *
0-
02
b111 6
#601430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#601440000000
0!
0%
b0 *
0-
02
b0 6
#601450000000
1!
1%
1-
12
#601460000000
0!
0%
b1 *
0-
02
b1 6
#601470000000
1!
1%
1-
12
#601480000000
0!
0%
b10 *
0-
02
b10 6
#601490000000
1!
1%
1-
12
#601500000000
0!
0%
b11 *
0-
02
b11 6
#601510000000
1!
1%
1-
12
15
#601520000000
0!
0%
b100 *
0-
02
b100 6
#601530000000
1!
1%
1-
12
#601540000000
0!
0%
b101 *
0-
02
b101 6
#601550000000
1!
1%
1-
12
#601560000000
0!
0%
b110 *
0-
02
b110 6
#601570000000
1!
1%
1-
12
#601580000000
0!
0%
b111 *
0-
02
b111 6
#601590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#601600000000
0!
0%
b0 *
0-
02
b0 6
#601610000000
1!
1%
1-
12
#601620000000
0!
0%
b1 *
0-
02
b1 6
#601630000000
1!
1%
1-
12
#601640000000
0!
0%
b10 *
0-
02
b10 6
#601650000000
1!
1%
1-
12
#601660000000
0!
0%
b11 *
0-
02
b11 6
#601670000000
1!
1%
1-
12
15
#601680000000
0!
0%
b100 *
0-
02
b100 6
#601690000000
1!
1%
1-
12
#601700000000
0!
0%
b101 *
0-
02
b101 6
#601710000000
1!
1%
1-
12
#601720000000
0!
0%
b110 *
0-
02
b110 6
#601730000000
1!
1%
1-
12
#601740000000
0!
0%
b111 *
0-
02
b111 6
#601750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#601760000000
0!
0%
b0 *
0-
02
b0 6
#601770000000
1!
1%
1-
12
#601780000000
0!
0%
b1 *
0-
02
b1 6
#601790000000
1!
1%
1-
12
#601800000000
0!
0%
b10 *
0-
02
b10 6
#601810000000
1!
1%
1-
12
#601820000000
0!
0%
b11 *
0-
02
b11 6
#601830000000
1!
1%
1-
12
15
#601840000000
0!
0%
b100 *
0-
02
b100 6
#601850000000
1!
1%
1-
12
#601860000000
0!
0%
b101 *
0-
02
b101 6
#601870000000
1!
1%
1-
12
#601880000000
0!
0%
b110 *
0-
02
b110 6
#601890000000
1!
1%
1-
12
#601900000000
0!
0%
b111 *
0-
02
b111 6
#601910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#601920000000
0!
0%
b0 *
0-
02
b0 6
#601930000000
1!
1%
1-
12
#601940000000
0!
0%
b1 *
0-
02
b1 6
#601950000000
1!
1%
1-
12
#601960000000
0!
0%
b10 *
0-
02
b10 6
#601970000000
1!
1%
1-
12
#601980000000
0!
0%
b11 *
0-
02
b11 6
#601990000000
1!
1%
1-
12
15
#602000000000
0!
0%
b100 *
0-
02
b100 6
#602010000000
1!
1%
1-
12
#602020000000
0!
0%
b101 *
0-
02
b101 6
#602030000000
1!
1%
1-
12
#602040000000
0!
0%
b110 *
0-
02
b110 6
#602050000000
1!
1%
1-
12
#602060000000
0!
0%
b111 *
0-
02
b111 6
#602070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#602080000000
0!
0%
b0 *
0-
02
b0 6
#602090000000
1!
1%
1-
12
#602100000000
0!
0%
b1 *
0-
02
b1 6
#602110000000
1!
1%
1-
12
#602120000000
0!
0%
b10 *
0-
02
b10 6
#602130000000
1!
1%
1-
12
#602140000000
0!
0%
b11 *
0-
02
b11 6
#602150000000
1!
1%
1-
12
15
#602160000000
0!
0%
b100 *
0-
02
b100 6
#602170000000
1!
1%
1-
12
#602180000000
0!
0%
b101 *
0-
02
b101 6
#602190000000
1!
1%
1-
12
#602200000000
0!
0%
b110 *
0-
02
b110 6
#602210000000
1!
1%
1-
12
#602220000000
0!
0%
b111 *
0-
02
b111 6
#602230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#602240000000
0!
0%
b0 *
0-
02
b0 6
#602250000000
1!
1%
1-
12
#602260000000
0!
0%
b1 *
0-
02
b1 6
#602270000000
1!
1%
1-
12
#602280000000
0!
0%
b10 *
0-
02
b10 6
#602290000000
1!
1%
1-
12
#602300000000
0!
0%
b11 *
0-
02
b11 6
#602310000000
1!
1%
1-
12
15
#602320000000
0!
0%
b100 *
0-
02
b100 6
#602330000000
1!
1%
1-
12
#602340000000
0!
0%
b101 *
0-
02
b101 6
#602350000000
1!
1%
1-
12
#602360000000
0!
0%
b110 *
0-
02
b110 6
#602370000000
1!
1%
1-
12
#602380000000
0!
0%
b111 *
0-
02
b111 6
#602390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#602400000000
0!
0%
b0 *
0-
02
b0 6
#602410000000
1!
1%
1-
12
#602420000000
0!
0%
b1 *
0-
02
b1 6
#602430000000
1!
1%
1-
12
#602440000000
0!
0%
b10 *
0-
02
b10 6
#602450000000
1!
1%
1-
12
#602460000000
0!
0%
b11 *
0-
02
b11 6
#602470000000
1!
1%
1-
12
15
#602480000000
0!
0%
b100 *
0-
02
b100 6
#602490000000
1!
1%
1-
12
#602500000000
0!
0%
b101 *
0-
02
b101 6
#602510000000
1!
1%
1-
12
#602520000000
0!
0%
b110 *
0-
02
b110 6
#602530000000
1!
1%
1-
12
#602540000000
0!
0%
b111 *
0-
02
b111 6
#602550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#602560000000
0!
0%
b0 *
0-
02
b0 6
#602570000000
1!
1%
1-
12
#602580000000
0!
0%
b1 *
0-
02
b1 6
#602590000000
1!
1%
1-
12
#602600000000
0!
0%
b10 *
0-
02
b10 6
#602610000000
1!
1%
1-
12
#602620000000
0!
0%
b11 *
0-
02
b11 6
#602630000000
1!
1%
1-
12
15
#602640000000
0!
0%
b100 *
0-
02
b100 6
#602650000000
1!
1%
1-
12
#602660000000
0!
0%
b101 *
0-
02
b101 6
#602670000000
1!
1%
1-
12
#602680000000
0!
0%
b110 *
0-
02
b110 6
#602690000000
1!
1%
1-
12
#602700000000
0!
0%
b111 *
0-
02
b111 6
#602710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#602720000000
0!
0%
b0 *
0-
02
b0 6
#602730000000
1!
1%
1-
12
#602740000000
0!
0%
b1 *
0-
02
b1 6
#602750000000
1!
1%
1-
12
#602760000000
0!
0%
b10 *
0-
02
b10 6
#602770000000
1!
1%
1-
12
#602780000000
0!
0%
b11 *
0-
02
b11 6
#602790000000
1!
1%
1-
12
15
#602800000000
0!
0%
b100 *
0-
02
b100 6
#602810000000
1!
1%
1-
12
#602820000000
0!
0%
b101 *
0-
02
b101 6
#602830000000
1!
1%
1-
12
#602840000000
0!
0%
b110 *
0-
02
b110 6
#602850000000
1!
1%
1-
12
#602860000000
0!
0%
b111 *
0-
02
b111 6
#602870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#602880000000
0!
0%
b0 *
0-
02
b0 6
#602890000000
1!
1%
1-
12
#602900000000
0!
0%
b1 *
0-
02
b1 6
#602910000000
1!
1%
1-
12
#602920000000
0!
0%
b10 *
0-
02
b10 6
#602930000000
1!
1%
1-
12
#602940000000
0!
0%
b11 *
0-
02
b11 6
#602950000000
1!
1%
1-
12
15
#602960000000
0!
0%
b100 *
0-
02
b100 6
#602970000000
1!
1%
1-
12
#602980000000
0!
0%
b101 *
0-
02
b101 6
#602990000000
1!
1%
1-
12
#603000000000
0!
0%
b110 *
0-
02
b110 6
#603010000000
1!
1%
1-
12
#603020000000
0!
0%
b111 *
0-
02
b111 6
#603030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#603040000000
0!
0%
b0 *
0-
02
b0 6
#603050000000
1!
1%
1-
12
#603060000000
0!
0%
b1 *
0-
02
b1 6
#603070000000
1!
1%
1-
12
#603080000000
0!
0%
b10 *
0-
02
b10 6
#603090000000
1!
1%
1-
12
#603100000000
0!
0%
b11 *
0-
02
b11 6
#603110000000
1!
1%
1-
12
15
#603120000000
0!
0%
b100 *
0-
02
b100 6
#603130000000
1!
1%
1-
12
#603140000000
0!
0%
b101 *
0-
02
b101 6
#603150000000
1!
1%
1-
12
#603160000000
0!
0%
b110 *
0-
02
b110 6
#603170000000
1!
1%
1-
12
#603180000000
0!
0%
b111 *
0-
02
b111 6
#603190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#603200000000
0!
0%
b0 *
0-
02
b0 6
#603210000000
1!
1%
1-
12
#603220000000
0!
0%
b1 *
0-
02
b1 6
#603230000000
1!
1%
1-
12
#603240000000
0!
0%
b10 *
0-
02
b10 6
#603250000000
1!
1%
1-
12
#603260000000
0!
0%
b11 *
0-
02
b11 6
#603270000000
1!
1%
1-
12
15
#603280000000
0!
0%
b100 *
0-
02
b100 6
#603290000000
1!
1%
1-
12
#603300000000
0!
0%
b101 *
0-
02
b101 6
#603310000000
1!
1%
1-
12
#603320000000
0!
0%
b110 *
0-
02
b110 6
#603330000000
1!
1%
1-
12
#603340000000
0!
0%
b111 *
0-
02
b111 6
#603350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#603360000000
0!
0%
b0 *
0-
02
b0 6
#603370000000
1!
1%
1-
12
#603380000000
0!
0%
b1 *
0-
02
b1 6
#603390000000
1!
1%
1-
12
#603400000000
0!
0%
b10 *
0-
02
b10 6
#603410000000
1!
1%
1-
12
#603420000000
0!
0%
b11 *
0-
02
b11 6
#603430000000
1!
1%
1-
12
15
#603440000000
0!
0%
b100 *
0-
02
b100 6
#603450000000
1!
1%
1-
12
#603460000000
0!
0%
b101 *
0-
02
b101 6
#603470000000
1!
1%
1-
12
#603480000000
0!
0%
b110 *
0-
02
b110 6
#603490000000
1!
1%
1-
12
#603500000000
0!
0%
b111 *
0-
02
b111 6
#603510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#603520000000
0!
0%
b0 *
0-
02
b0 6
#603530000000
1!
1%
1-
12
#603540000000
0!
0%
b1 *
0-
02
b1 6
#603550000000
1!
1%
1-
12
#603560000000
0!
0%
b10 *
0-
02
b10 6
#603570000000
1!
1%
1-
12
#603580000000
0!
0%
b11 *
0-
02
b11 6
#603590000000
1!
1%
1-
12
15
#603600000000
0!
0%
b100 *
0-
02
b100 6
#603610000000
1!
1%
1-
12
#603620000000
0!
0%
b101 *
0-
02
b101 6
#603630000000
1!
1%
1-
12
#603640000000
0!
0%
b110 *
0-
02
b110 6
#603650000000
1!
1%
1-
12
#603660000000
0!
0%
b111 *
0-
02
b111 6
#603670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#603680000000
0!
0%
b0 *
0-
02
b0 6
#603690000000
1!
1%
1-
12
#603700000000
0!
0%
b1 *
0-
02
b1 6
#603710000000
1!
1%
1-
12
#603720000000
0!
0%
b10 *
0-
02
b10 6
#603730000000
1!
1%
1-
12
#603740000000
0!
0%
b11 *
0-
02
b11 6
#603750000000
1!
1%
1-
12
15
#603760000000
0!
0%
b100 *
0-
02
b100 6
#603770000000
1!
1%
1-
12
#603780000000
0!
0%
b101 *
0-
02
b101 6
#603790000000
1!
1%
1-
12
#603800000000
0!
0%
b110 *
0-
02
b110 6
#603810000000
1!
1%
1-
12
#603820000000
0!
0%
b111 *
0-
02
b111 6
#603830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#603840000000
0!
0%
b0 *
0-
02
b0 6
#603850000000
1!
1%
1-
12
#603860000000
0!
0%
b1 *
0-
02
b1 6
#603870000000
1!
1%
1-
12
#603880000000
0!
0%
b10 *
0-
02
b10 6
#603890000000
1!
1%
1-
12
#603900000000
0!
0%
b11 *
0-
02
b11 6
#603910000000
1!
1%
1-
12
15
#603920000000
0!
0%
b100 *
0-
02
b100 6
#603930000000
1!
1%
1-
12
#603940000000
0!
0%
b101 *
0-
02
b101 6
#603950000000
1!
1%
1-
12
#603960000000
0!
0%
b110 *
0-
02
b110 6
#603970000000
1!
1%
1-
12
#603980000000
0!
0%
b111 *
0-
02
b111 6
#603990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#604000000000
0!
0%
b0 *
0-
02
b0 6
#604010000000
1!
1%
1-
12
#604020000000
0!
0%
b1 *
0-
02
b1 6
#604030000000
1!
1%
1-
12
#604040000000
0!
0%
b10 *
0-
02
b10 6
#604050000000
1!
1%
1-
12
#604060000000
0!
0%
b11 *
0-
02
b11 6
#604070000000
1!
1%
1-
12
15
#604080000000
0!
0%
b100 *
0-
02
b100 6
#604090000000
1!
1%
1-
12
#604100000000
0!
0%
b101 *
0-
02
b101 6
#604110000000
1!
1%
1-
12
#604120000000
0!
0%
b110 *
0-
02
b110 6
#604130000000
1!
1%
1-
12
#604140000000
0!
0%
b111 *
0-
02
b111 6
#604150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#604160000000
0!
0%
b0 *
0-
02
b0 6
#604170000000
1!
1%
1-
12
#604180000000
0!
0%
b1 *
0-
02
b1 6
#604190000000
1!
1%
1-
12
#604200000000
0!
0%
b10 *
0-
02
b10 6
#604210000000
1!
1%
1-
12
#604220000000
0!
0%
b11 *
0-
02
b11 6
#604230000000
1!
1%
1-
12
15
#604240000000
0!
0%
b100 *
0-
02
b100 6
#604250000000
1!
1%
1-
12
#604260000000
0!
0%
b101 *
0-
02
b101 6
#604270000000
1!
1%
1-
12
#604280000000
0!
0%
b110 *
0-
02
b110 6
#604290000000
1!
1%
1-
12
#604300000000
0!
0%
b111 *
0-
02
b111 6
#604310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#604320000000
0!
0%
b0 *
0-
02
b0 6
#604330000000
1!
1%
1-
12
#604340000000
0!
0%
b1 *
0-
02
b1 6
#604350000000
1!
1%
1-
12
#604360000000
0!
0%
b10 *
0-
02
b10 6
#604370000000
1!
1%
1-
12
#604380000000
0!
0%
b11 *
0-
02
b11 6
#604390000000
1!
1%
1-
12
15
#604400000000
0!
0%
b100 *
0-
02
b100 6
#604410000000
1!
1%
1-
12
#604420000000
0!
0%
b101 *
0-
02
b101 6
#604430000000
1!
1%
1-
12
#604440000000
0!
0%
b110 *
0-
02
b110 6
#604450000000
1!
1%
1-
12
#604460000000
0!
0%
b111 *
0-
02
b111 6
#604470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#604480000000
0!
0%
b0 *
0-
02
b0 6
#604490000000
1!
1%
1-
12
#604500000000
0!
0%
b1 *
0-
02
b1 6
#604510000000
1!
1%
1-
12
#604520000000
0!
0%
b10 *
0-
02
b10 6
#604530000000
1!
1%
1-
12
#604540000000
0!
0%
b11 *
0-
02
b11 6
#604550000000
1!
1%
1-
12
15
#604560000000
0!
0%
b100 *
0-
02
b100 6
#604570000000
1!
1%
1-
12
#604580000000
0!
0%
b101 *
0-
02
b101 6
#604590000000
1!
1%
1-
12
#604600000000
0!
0%
b110 *
0-
02
b110 6
#604610000000
1!
1%
1-
12
#604620000000
0!
0%
b111 *
0-
02
b111 6
#604630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#604640000000
0!
0%
b0 *
0-
02
b0 6
#604650000000
1!
1%
1-
12
#604660000000
0!
0%
b1 *
0-
02
b1 6
#604670000000
1!
1%
1-
12
#604680000000
0!
0%
b10 *
0-
02
b10 6
#604690000000
1!
1%
1-
12
#604700000000
0!
0%
b11 *
0-
02
b11 6
#604710000000
1!
1%
1-
12
15
#604720000000
0!
0%
b100 *
0-
02
b100 6
#604730000000
1!
1%
1-
12
#604740000000
0!
0%
b101 *
0-
02
b101 6
#604750000000
1!
1%
1-
12
#604760000000
0!
0%
b110 *
0-
02
b110 6
#604770000000
1!
1%
1-
12
#604780000000
0!
0%
b111 *
0-
02
b111 6
#604790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#604800000000
0!
0%
b0 *
0-
02
b0 6
#604810000000
1!
1%
1-
12
#604820000000
0!
0%
b1 *
0-
02
b1 6
#604830000000
1!
1%
1-
12
#604840000000
0!
0%
b10 *
0-
02
b10 6
#604850000000
1!
1%
1-
12
#604860000000
0!
0%
b11 *
0-
02
b11 6
#604870000000
1!
1%
1-
12
15
#604880000000
0!
0%
b100 *
0-
02
b100 6
#604890000000
1!
1%
1-
12
#604900000000
0!
0%
b101 *
0-
02
b101 6
#604910000000
1!
1%
1-
12
#604920000000
0!
0%
b110 *
0-
02
b110 6
#604930000000
1!
1%
1-
12
#604940000000
0!
0%
b111 *
0-
02
b111 6
#604950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#604960000000
0!
0%
b0 *
0-
02
b0 6
#604970000000
1!
1%
1-
12
#604980000000
0!
0%
b1 *
0-
02
b1 6
#604990000000
1!
1%
1-
12
#605000000000
0!
0%
b10 *
0-
02
b10 6
#605010000000
1!
1%
1-
12
#605020000000
0!
0%
b11 *
0-
02
b11 6
#605030000000
1!
1%
1-
12
15
#605040000000
0!
0%
b100 *
0-
02
b100 6
#605050000000
1!
1%
1-
12
#605060000000
0!
0%
b101 *
0-
02
b101 6
#605070000000
1!
1%
1-
12
#605080000000
0!
0%
b110 *
0-
02
b110 6
#605090000000
1!
1%
1-
12
#605100000000
0!
0%
b111 *
0-
02
b111 6
#605110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#605120000000
0!
0%
b0 *
0-
02
b0 6
#605130000000
1!
1%
1-
12
#605140000000
0!
0%
b1 *
0-
02
b1 6
#605150000000
1!
1%
1-
12
#605160000000
0!
0%
b10 *
0-
02
b10 6
#605170000000
1!
1%
1-
12
#605180000000
0!
0%
b11 *
0-
02
b11 6
#605190000000
1!
1%
1-
12
15
#605200000000
0!
0%
b100 *
0-
02
b100 6
#605210000000
1!
1%
1-
12
#605220000000
0!
0%
b101 *
0-
02
b101 6
#605230000000
1!
1%
1-
12
#605240000000
0!
0%
b110 *
0-
02
b110 6
#605250000000
1!
1%
1-
12
#605260000000
0!
0%
b111 *
0-
02
b111 6
#605270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#605280000000
0!
0%
b0 *
0-
02
b0 6
#605290000000
1!
1%
1-
12
#605300000000
0!
0%
b1 *
0-
02
b1 6
#605310000000
1!
1%
1-
12
#605320000000
0!
0%
b10 *
0-
02
b10 6
#605330000000
1!
1%
1-
12
#605340000000
0!
0%
b11 *
0-
02
b11 6
#605350000000
1!
1%
1-
12
15
#605360000000
0!
0%
b100 *
0-
02
b100 6
#605370000000
1!
1%
1-
12
#605380000000
0!
0%
b101 *
0-
02
b101 6
#605390000000
1!
1%
1-
12
#605400000000
0!
0%
b110 *
0-
02
b110 6
#605410000000
1!
1%
1-
12
#605420000000
0!
0%
b111 *
0-
02
b111 6
#605430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#605440000000
0!
0%
b0 *
0-
02
b0 6
#605450000000
1!
1%
1-
12
#605460000000
0!
0%
b1 *
0-
02
b1 6
#605470000000
1!
1%
1-
12
#605480000000
0!
0%
b10 *
0-
02
b10 6
#605490000000
1!
1%
1-
12
#605500000000
0!
0%
b11 *
0-
02
b11 6
#605510000000
1!
1%
1-
12
15
#605520000000
0!
0%
b100 *
0-
02
b100 6
#605530000000
1!
1%
1-
12
#605540000000
0!
0%
b101 *
0-
02
b101 6
#605550000000
1!
1%
1-
12
#605560000000
0!
0%
b110 *
0-
02
b110 6
#605570000000
1!
1%
1-
12
#605580000000
0!
0%
b111 *
0-
02
b111 6
#605590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#605600000000
0!
0%
b0 *
0-
02
b0 6
#605610000000
1!
1%
1-
12
#605620000000
0!
0%
b1 *
0-
02
b1 6
#605630000000
1!
1%
1-
12
#605640000000
0!
0%
b10 *
0-
02
b10 6
#605650000000
1!
1%
1-
12
#605660000000
0!
0%
b11 *
0-
02
b11 6
#605670000000
1!
1%
1-
12
15
#605680000000
0!
0%
b100 *
0-
02
b100 6
#605690000000
1!
1%
1-
12
#605700000000
0!
0%
b101 *
0-
02
b101 6
#605710000000
1!
1%
1-
12
#605720000000
0!
0%
b110 *
0-
02
b110 6
#605730000000
1!
1%
1-
12
#605740000000
0!
0%
b111 *
0-
02
b111 6
#605750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#605760000000
0!
0%
b0 *
0-
02
b0 6
#605770000000
1!
1%
1-
12
#605780000000
0!
0%
b1 *
0-
02
b1 6
#605790000000
1!
1%
1-
12
#605800000000
0!
0%
b10 *
0-
02
b10 6
#605810000000
1!
1%
1-
12
#605820000000
0!
0%
b11 *
0-
02
b11 6
#605830000000
1!
1%
1-
12
15
#605840000000
0!
0%
b100 *
0-
02
b100 6
#605850000000
1!
1%
1-
12
#605860000000
0!
0%
b101 *
0-
02
b101 6
#605870000000
1!
1%
1-
12
#605880000000
0!
0%
b110 *
0-
02
b110 6
#605890000000
1!
1%
1-
12
#605900000000
0!
0%
b111 *
0-
02
b111 6
#605910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#605920000000
0!
0%
b0 *
0-
02
b0 6
#605930000000
1!
1%
1-
12
#605940000000
0!
0%
b1 *
0-
02
b1 6
#605950000000
1!
1%
1-
12
#605960000000
0!
0%
b10 *
0-
02
b10 6
#605970000000
1!
1%
1-
12
#605980000000
0!
0%
b11 *
0-
02
b11 6
#605990000000
1!
1%
1-
12
15
#606000000000
0!
0%
b100 *
0-
02
b100 6
#606010000000
1!
1%
1-
12
#606020000000
0!
0%
b101 *
0-
02
b101 6
#606030000000
1!
1%
1-
12
#606040000000
0!
0%
b110 *
0-
02
b110 6
#606050000000
1!
1%
1-
12
#606060000000
0!
0%
b111 *
0-
02
b111 6
#606070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#606080000000
0!
0%
b0 *
0-
02
b0 6
#606090000000
1!
1%
1-
12
#606100000000
0!
0%
b1 *
0-
02
b1 6
#606110000000
1!
1%
1-
12
#606120000000
0!
0%
b10 *
0-
02
b10 6
#606130000000
1!
1%
1-
12
#606140000000
0!
0%
b11 *
0-
02
b11 6
#606150000000
1!
1%
1-
12
15
#606160000000
0!
0%
b100 *
0-
02
b100 6
#606170000000
1!
1%
1-
12
#606180000000
0!
0%
b101 *
0-
02
b101 6
#606190000000
1!
1%
1-
12
#606200000000
0!
0%
b110 *
0-
02
b110 6
#606210000000
1!
1%
1-
12
#606220000000
0!
0%
b111 *
0-
02
b111 6
#606230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#606240000000
0!
0%
b0 *
0-
02
b0 6
#606250000000
1!
1%
1-
12
#606260000000
0!
0%
b1 *
0-
02
b1 6
#606270000000
1!
1%
1-
12
#606280000000
0!
0%
b10 *
0-
02
b10 6
#606290000000
1!
1%
1-
12
#606300000000
0!
0%
b11 *
0-
02
b11 6
#606310000000
1!
1%
1-
12
15
#606320000000
0!
0%
b100 *
0-
02
b100 6
#606330000000
1!
1%
1-
12
#606340000000
0!
0%
b101 *
0-
02
b101 6
#606350000000
1!
1%
1-
12
#606360000000
0!
0%
b110 *
0-
02
b110 6
#606370000000
1!
1%
1-
12
#606380000000
0!
0%
b111 *
0-
02
b111 6
#606390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#606400000000
0!
0%
b0 *
0-
02
b0 6
#606410000000
1!
1%
1-
12
#606420000000
0!
0%
b1 *
0-
02
b1 6
#606430000000
1!
1%
1-
12
#606440000000
0!
0%
b10 *
0-
02
b10 6
#606450000000
1!
1%
1-
12
#606460000000
0!
0%
b11 *
0-
02
b11 6
#606470000000
1!
1%
1-
12
15
#606480000000
0!
0%
b100 *
0-
02
b100 6
#606490000000
1!
1%
1-
12
#606500000000
0!
0%
b101 *
0-
02
b101 6
#606510000000
1!
1%
1-
12
#606520000000
0!
0%
b110 *
0-
02
b110 6
#606530000000
1!
1%
1-
12
#606540000000
0!
0%
b111 *
0-
02
b111 6
#606550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#606560000000
0!
0%
b0 *
0-
02
b0 6
#606570000000
1!
1%
1-
12
#606580000000
0!
0%
b1 *
0-
02
b1 6
#606590000000
1!
1%
1-
12
#606600000000
0!
0%
b10 *
0-
02
b10 6
#606610000000
1!
1%
1-
12
#606620000000
0!
0%
b11 *
0-
02
b11 6
#606630000000
1!
1%
1-
12
15
#606640000000
0!
0%
b100 *
0-
02
b100 6
#606650000000
1!
1%
1-
12
#606660000000
0!
0%
b101 *
0-
02
b101 6
#606670000000
1!
1%
1-
12
#606680000000
0!
0%
b110 *
0-
02
b110 6
#606690000000
1!
1%
1-
12
#606700000000
0!
0%
b111 *
0-
02
b111 6
#606710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#606720000000
0!
0%
b0 *
0-
02
b0 6
#606730000000
1!
1%
1-
12
#606740000000
0!
0%
b1 *
0-
02
b1 6
#606750000000
1!
1%
1-
12
#606760000000
0!
0%
b10 *
0-
02
b10 6
#606770000000
1!
1%
1-
12
#606780000000
0!
0%
b11 *
0-
02
b11 6
#606790000000
1!
1%
1-
12
15
#606800000000
0!
0%
b100 *
0-
02
b100 6
#606810000000
1!
1%
1-
12
#606820000000
0!
0%
b101 *
0-
02
b101 6
#606830000000
1!
1%
1-
12
#606840000000
0!
0%
b110 *
0-
02
b110 6
#606850000000
1!
1%
1-
12
#606860000000
0!
0%
b111 *
0-
02
b111 6
#606870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#606880000000
0!
0%
b0 *
0-
02
b0 6
#606890000000
1!
1%
1-
12
#606900000000
0!
0%
b1 *
0-
02
b1 6
#606910000000
1!
1%
1-
12
#606920000000
0!
0%
b10 *
0-
02
b10 6
#606930000000
1!
1%
1-
12
#606940000000
0!
0%
b11 *
0-
02
b11 6
#606950000000
1!
1%
1-
12
15
#606960000000
0!
0%
b100 *
0-
02
b100 6
#606970000000
1!
1%
1-
12
#606980000000
0!
0%
b101 *
0-
02
b101 6
#606990000000
1!
1%
1-
12
#607000000000
0!
0%
b110 *
0-
02
b110 6
#607010000000
1!
1%
1-
12
#607020000000
0!
0%
b111 *
0-
02
b111 6
#607030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#607040000000
0!
0%
b0 *
0-
02
b0 6
#607050000000
1!
1%
1-
12
#607060000000
0!
0%
b1 *
0-
02
b1 6
#607070000000
1!
1%
1-
12
#607080000000
0!
0%
b10 *
0-
02
b10 6
#607090000000
1!
1%
1-
12
#607100000000
0!
0%
b11 *
0-
02
b11 6
#607110000000
1!
1%
1-
12
15
#607120000000
0!
0%
b100 *
0-
02
b100 6
#607130000000
1!
1%
1-
12
#607140000000
0!
0%
b101 *
0-
02
b101 6
#607150000000
1!
1%
1-
12
#607160000000
0!
0%
b110 *
0-
02
b110 6
#607170000000
1!
1%
1-
12
#607180000000
0!
0%
b111 *
0-
02
b111 6
#607190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#607200000000
0!
0%
b0 *
0-
02
b0 6
#607210000000
1!
1%
1-
12
#607220000000
0!
0%
b1 *
0-
02
b1 6
#607230000000
1!
1%
1-
12
#607240000000
0!
0%
b10 *
0-
02
b10 6
#607250000000
1!
1%
1-
12
#607260000000
0!
0%
b11 *
0-
02
b11 6
#607270000000
1!
1%
1-
12
15
#607280000000
0!
0%
b100 *
0-
02
b100 6
#607290000000
1!
1%
1-
12
#607300000000
0!
0%
b101 *
0-
02
b101 6
#607310000000
1!
1%
1-
12
#607320000000
0!
0%
b110 *
0-
02
b110 6
#607330000000
1!
1%
1-
12
#607340000000
0!
0%
b111 *
0-
02
b111 6
#607350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#607360000000
0!
0%
b0 *
0-
02
b0 6
#607370000000
1!
1%
1-
12
#607380000000
0!
0%
b1 *
0-
02
b1 6
#607390000000
1!
1%
1-
12
#607400000000
0!
0%
b10 *
0-
02
b10 6
#607410000000
1!
1%
1-
12
#607420000000
0!
0%
b11 *
0-
02
b11 6
#607430000000
1!
1%
1-
12
15
#607440000000
0!
0%
b100 *
0-
02
b100 6
#607450000000
1!
1%
1-
12
#607460000000
0!
0%
b101 *
0-
02
b101 6
#607470000000
1!
1%
1-
12
#607480000000
0!
0%
b110 *
0-
02
b110 6
#607490000000
1!
1%
1-
12
#607500000000
0!
0%
b111 *
0-
02
b111 6
#607510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#607520000000
0!
0%
b0 *
0-
02
b0 6
#607530000000
1!
1%
1-
12
#607540000000
0!
0%
b1 *
0-
02
b1 6
#607550000000
1!
1%
1-
12
#607560000000
0!
0%
b10 *
0-
02
b10 6
#607570000000
1!
1%
1-
12
#607580000000
0!
0%
b11 *
0-
02
b11 6
#607590000000
1!
1%
1-
12
15
#607600000000
0!
0%
b100 *
0-
02
b100 6
#607610000000
1!
1%
1-
12
#607620000000
0!
0%
b101 *
0-
02
b101 6
#607630000000
1!
1%
1-
12
#607640000000
0!
0%
b110 *
0-
02
b110 6
#607650000000
1!
1%
1-
12
#607660000000
0!
0%
b111 *
0-
02
b111 6
#607670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#607680000000
0!
0%
b0 *
0-
02
b0 6
#607690000000
1!
1%
1-
12
#607700000000
0!
0%
b1 *
0-
02
b1 6
#607710000000
1!
1%
1-
12
#607720000000
0!
0%
b10 *
0-
02
b10 6
#607730000000
1!
1%
1-
12
#607740000000
0!
0%
b11 *
0-
02
b11 6
#607750000000
1!
1%
1-
12
15
#607760000000
0!
0%
b100 *
0-
02
b100 6
#607770000000
1!
1%
1-
12
#607780000000
0!
0%
b101 *
0-
02
b101 6
#607790000000
1!
1%
1-
12
#607800000000
0!
0%
b110 *
0-
02
b110 6
#607810000000
1!
1%
1-
12
#607820000000
0!
0%
b111 *
0-
02
b111 6
#607830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#607840000000
0!
0%
b0 *
0-
02
b0 6
#607850000000
1!
1%
1-
12
#607860000000
0!
0%
b1 *
0-
02
b1 6
#607870000000
1!
1%
1-
12
#607880000000
0!
0%
b10 *
0-
02
b10 6
#607890000000
1!
1%
1-
12
#607900000000
0!
0%
b11 *
0-
02
b11 6
#607910000000
1!
1%
1-
12
15
#607920000000
0!
0%
b100 *
0-
02
b100 6
#607930000000
1!
1%
1-
12
#607940000000
0!
0%
b101 *
0-
02
b101 6
#607950000000
1!
1%
1-
12
#607960000000
0!
0%
b110 *
0-
02
b110 6
#607970000000
1!
1%
1-
12
#607980000000
0!
0%
b111 *
0-
02
b111 6
#607990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#608000000000
0!
0%
b0 *
0-
02
b0 6
#608010000000
1!
1%
1-
12
#608020000000
0!
0%
b1 *
0-
02
b1 6
#608030000000
1!
1%
1-
12
#608040000000
0!
0%
b10 *
0-
02
b10 6
#608050000000
1!
1%
1-
12
#608060000000
0!
0%
b11 *
0-
02
b11 6
#608070000000
1!
1%
1-
12
15
#608080000000
0!
0%
b100 *
0-
02
b100 6
#608090000000
1!
1%
1-
12
#608100000000
0!
0%
b101 *
0-
02
b101 6
#608110000000
1!
1%
1-
12
#608120000000
0!
0%
b110 *
0-
02
b110 6
#608130000000
1!
1%
1-
12
#608140000000
0!
0%
b111 *
0-
02
b111 6
#608150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#608160000000
0!
0%
b0 *
0-
02
b0 6
#608170000000
1!
1%
1-
12
#608180000000
0!
0%
b1 *
0-
02
b1 6
#608190000000
1!
1%
1-
12
#608200000000
0!
0%
b10 *
0-
02
b10 6
#608210000000
1!
1%
1-
12
#608220000000
0!
0%
b11 *
0-
02
b11 6
#608230000000
1!
1%
1-
12
15
#608240000000
0!
0%
b100 *
0-
02
b100 6
#608250000000
1!
1%
1-
12
#608260000000
0!
0%
b101 *
0-
02
b101 6
#608270000000
1!
1%
1-
12
#608280000000
0!
0%
b110 *
0-
02
b110 6
#608290000000
1!
1%
1-
12
#608300000000
0!
0%
b111 *
0-
02
b111 6
#608310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#608320000000
0!
0%
b0 *
0-
02
b0 6
#608330000000
1!
1%
1-
12
#608340000000
0!
0%
b1 *
0-
02
b1 6
#608350000000
1!
1%
1-
12
#608360000000
0!
0%
b10 *
0-
02
b10 6
#608370000000
1!
1%
1-
12
#608380000000
0!
0%
b11 *
0-
02
b11 6
#608390000000
1!
1%
1-
12
15
#608400000000
0!
0%
b100 *
0-
02
b100 6
#608410000000
1!
1%
1-
12
#608420000000
0!
0%
b101 *
0-
02
b101 6
#608430000000
1!
1%
1-
12
#608440000000
0!
0%
b110 *
0-
02
b110 6
#608450000000
1!
1%
1-
12
#608460000000
0!
0%
b111 *
0-
02
b111 6
#608470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#608480000000
0!
0%
b0 *
0-
02
b0 6
#608490000000
1!
1%
1-
12
#608500000000
0!
0%
b1 *
0-
02
b1 6
#608510000000
1!
1%
1-
12
#608520000000
0!
0%
b10 *
0-
02
b10 6
#608530000000
1!
1%
1-
12
#608540000000
0!
0%
b11 *
0-
02
b11 6
#608550000000
1!
1%
1-
12
15
#608560000000
0!
0%
b100 *
0-
02
b100 6
#608570000000
1!
1%
1-
12
#608580000000
0!
0%
b101 *
0-
02
b101 6
#608590000000
1!
1%
1-
12
#608600000000
0!
0%
b110 *
0-
02
b110 6
#608610000000
1!
1%
1-
12
#608620000000
0!
0%
b111 *
0-
02
b111 6
#608630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#608640000000
0!
0%
b0 *
0-
02
b0 6
#608650000000
1!
1%
1-
12
#608660000000
0!
0%
b1 *
0-
02
b1 6
#608670000000
1!
1%
1-
12
#608680000000
0!
0%
b10 *
0-
02
b10 6
#608690000000
1!
1%
1-
12
#608700000000
0!
0%
b11 *
0-
02
b11 6
#608710000000
1!
1%
1-
12
15
#608720000000
0!
0%
b100 *
0-
02
b100 6
#608730000000
1!
1%
1-
12
#608740000000
0!
0%
b101 *
0-
02
b101 6
#608750000000
1!
1%
1-
12
#608760000000
0!
0%
b110 *
0-
02
b110 6
#608770000000
1!
1%
1-
12
#608780000000
0!
0%
b111 *
0-
02
b111 6
#608790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#608800000000
0!
0%
b0 *
0-
02
b0 6
#608810000000
1!
1%
1-
12
#608820000000
0!
0%
b1 *
0-
02
b1 6
#608830000000
1!
1%
1-
12
#608840000000
0!
0%
b10 *
0-
02
b10 6
#608850000000
1!
1%
1-
12
#608860000000
0!
0%
b11 *
0-
02
b11 6
#608870000000
1!
1%
1-
12
15
#608880000000
0!
0%
b100 *
0-
02
b100 6
#608890000000
1!
1%
1-
12
#608900000000
0!
0%
b101 *
0-
02
b101 6
#608910000000
1!
1%
1-
12
#608920000000
0!
0%
b110 *
0-
02
b110 6
#608930000000
1!
1%
1-
12
#608940000000
0!
0%
b111 *
0-
02
b111 6
#608950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#608960000000
0!
0%
b0 *
0-
02
b0 6
#608970000000
1!
1%
1-
12
#608980000000
0!
0%
b1 *
0-
02
b1 6
#608990000000
1!
1%
1-
12
#609000000000
0!
0%
b10 *
0-
02
b10 6
#609010000000
1!
1%
1-
12
#609020000000
0!
0%
b11 *
0-
02
b11 6
#609030000000
1!
1%
1-
12
15
#609040000000
0!
0%
b100 *
0-
02
b100 6
#609050000000
1!
1%
1-
12
#609060000000
0!
0%
b101 *
0-
02
b101 6
#609070000000
1!
1%
1-
12
#609080000000
0!
0%
b110 *
0-
02
b110 6
#609090000000
1!
1%
1-
12
#609100000000
0!
0%
b111 *
0-
02
b111 6
#609110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#609120000000
0!
0%
b0 *
0-
02
b0 6
#609130000000
1!
1%
1-
12
#609140000000
0!
0%
b1 *
0-
02
b1 6
#609150000000
1!
1%
1-
12
#609160000000
0!
0%
b10 *
0-
02
b10 6
#609170000000
1!
1%
1-
12
#609180000000
0!
0%
b11 *
0-
02
b11 6
#609190000000
1!
1%
1-
12
15
#609200000000
0!
0%
b100 *
0-
02
b100 6
#609210000000
1!
1%
1-
12
#609220000000
0!
0%
b101 *
0-
02
b101 6
#609230000000
1!
1%
1-
12
#609240000000
0!
0%
b110 *
0-
02
b110 6
#609250000000
1!
1%
1-
12
#609260000000
0!
0%
b111 *
0-
02
b111 6
#609270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#609280000000
0!
0%
b0 *
0-
02
b0 6
#609290000000
1!
1%
1-
12
#609300000000
0!
0%
b1 *
0-
02
b1 6
#609310000000
1!
1%
1-
12
#609320000000
0!
0%
b10 *
0-
02
b10 6
#609330000000
1!
1%
1-
12
#609340000000
0!
0%
b11 *
0-
02
b11 6
#609350000000
1!
1%
1-
12
15
#609360000000
0!
0%
b100 *
0-
02
b100 6
#609370000000
1!
1%
1-
12
#609380000000
0!
0%
b101 *
0-
02
b101 6
#609390000000
1!
1%
1-
12
#609400000000
0!
0%
b110 *
0-
02
b110 6
#609410000000
1!
1%
1-
12
#609420000000
0!
0%
b111 *
0-
02
b111 6
#609430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#609440000000
0!
0%
b0 *
0-
02
b0 6
#609450000000
1!
1%
1-
12
#609460000000
0!
0%
b1 *
0-
02
b1 6
#609470000000
1!
1%
1-
12
#609480000000
0!
0%
b10 *
0-
02
b10 6
#609490000000
1!
1%
1-
12
#609500000000
0!
0%
b11 *
0-
02
b11 6
#609510000000
1!
1%
1-
12
15
#609520000000
0!
0%
b100 *
0-
02
b100 6
#609530000000
1!
1%
1-
12
#609540000000
0!
0%
b101 *
0-
02
b101 6
#609550000000
1!
1%
1-
12
#609560000000
0!
0%
b110 *
0-
02
b110 6
#609570000000
1!
1%
1-
12
#609580000000
0!
0%
b111 *
0-
02
b111 6
#609590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#609600000000
0!
0%
b0 *
0-
02
b0 6
#609610000000
1!
1%
1-
12
#609620000000
0!
0%
b1 *
0-
02
b1 6
#609630000000
1!
1%
1-
12
#609640000000
0!
0%
b10 *
0-
02
b10 6
#609650000000
1!
1%
1-
12
#609660000000
0!
0%
b11 *
0-
02
b11 6
#609670000000
1!
1%
1-
12
15
#609680000000
0!
0%
b100 *
0-
02
b100 6
#609690000000
1!
1%
1-
12
#609700000000
0!
0%
b101 *
0-
02
b101 6
#609710000000
1!
1%
1-
12
#609720000000
0!
0%
b110 *
0-
02
b110 6
#609730000000
1!
1%
1-
12
#609740000000
0!
0%
b111 *
0-
02
b111 6
#609750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#609760000000
0!
0%
b0 *
0-
02
b0 6
#609770000000
1!
1%
1-
12
#609780000000
0!
0%
b1 *
0-
02
b1 6
#609790000000
1!
1%
1-
12
#609800000000
0!
0%
b10 *
0-
02
b10 6
#609810000000
1!
1%
1-
12
#609820000000
0!
0%
b11 *
0-
02
b11 6
#609830000000
1!
1%
1-
12
15
#609840000000
0!
0%
b100 *
0-
02
b100 6
#609850000000
1!
1%
1-
12
#609860000000
0!
0%
b101 *
0-
02
b101 6
#609870000000
1!
1%
1-
12
#609880000000
0!
0%
b110 *
0-
02
b110 6
#609890000000
1!
1%
1-
12
#609900000000
0!
0%
b111 *
0-
02
b111 6
#609910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#609920000000
0!
0%
b0 *
0-
02
b0 6
#609930000000
1!
1%
1-
12
#609940000000
0!
0%
b1 *
0-
02
b1 6
#609950000000
1!
1%
1-
12
#609960000000
0!
0%
b10 *
0-
02
b10 6
#609970000000
1!
1%
1-
12
#609980000000
0!
0%
b11 *
0-
02
b11 6
#609990000000
1!
1%
1-
12
15
#610000000000
0!
0%
b100 *
0-
02
b100 6
#610010000000
1!
1%
1-
12
#610020000000
0!
0%
b101 *
0-
02
b101 6
#610030000000
1!
1%
1-
12
#610040000000
0!
0%
b110 *
0-
02
b110 6
#610050000000
1!
1%
1-
12
#610060000000
0!
0%
b111 *
0-
02
b111 6
#610070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#610080000000
0!
0%
b0 *
0-
02
b0 6
#610090000000
1!
1%
1-
12
#610100000000
0!
0%
b1 *
0-
02
b1 6
#610110000000
1!
1%
1-
12
#610120000000
0!
0%
b10 *
0-
02
b10 6
#610130000000
1!
1%
1-
12
#610140000000
0!
0%
b11 *
0-
02
b11 6
#610150000000
1!
1%
1-
12
15
#610160000000
0!
0%
b100 *
0-
02
b100 6
#610170000000
1!
1%
1-
12
#610180000000
0!
0%
b101 *
0-
02
b101 6
#610190000000
1!
1%
1-
12
#610200000000
0!
0%
b110 *
0-
02
b110 6
#610210000000
1!
1%
1-
12
#610220000000
0!
0%
b111 *
0-
02
b111 6
#610230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#610240000000
0!
0%
b0 *
0-
02
b0 6
#610250000000
1!
1%
1-
12
#610260000000
0!
0%
b1 *
0-
02
b1 6
#610270000000
1!
1%
1-
12
#610280000000
0!
0%
b10 *
0-
02
b10 6
#610290000000
1!
1%
1-
12
#610300000000
0!
0%
b11 *
0-
02
b11 6
#610310000000
1!
1%
1-
12
15
#610320000000
0!
0%
b100 *
0-
02
b100 6
#610330000000
1!
1%
1-
12
#610340000000
0!
0%
b101 *
0-
02
b101 6
#610350000000
1!
1%
1-
12
#610360000000
0!
0%
b110 *
0-
02
b110 6
#610370000000
1!
1%
1-
12
#610380000000
0!
0%
b111 *
0-
02
b111 6
#610390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#610400000000
0!
0%
b0 *
0-
02
b0 6
#610410000000
1!
1%
1-
12
#610420000000
0!
0%
b1 *
0-
02
b1 6
#610430000000
1!
1%
1-
12
#610440000000
0!
0%
b10 *
0-
02
b10 6
#610450000000
1!
1%
1-
12
#610460000000
0!
0%
b11 *
0-
02
b11 6
#610470000000
1!
1%
1-
12
15
#610480000000
0!
0%
b100 *
0-
02
b100 6
#610490000000
1!
1%
1-
12
#610500000000
0!
0%
b101 *
0-
02
b101 6
#610510000000
1!
1%
1-
12
#610520000000
0!
0%
b110 *
0-
02
b110 6
#610530000000
1!
1%
1-
12
#610540000000
0!
0%
b111 *
0-
02
b111 6
#610550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#610560000000
0!
0%
b0 *
0-
02
b0 6
#610570000000
1!
1%
1-
12
#610580000000
0!
0%
b1 *
0-
02
b1 6
#610590000000
1!
1%
1-
12
#610600000000
0!
0%
b10 *
0-
02
b10 6
#610610000000
1!
1%
1-
12
#610620000000
0!
0%
b11 *
0-
02
b11 6
#610630000000
1!
1%
1-
12
15
#610640000000
0!
0%
b100 *
0-
02
b100 6
#610650000000
1!
1%
1-
12
#610660000000
0!
0%
b101 *
0-
02
b101 6
#610670000000
1!
1%
1-
12
#610680000000
0!
0%
b110 *
0-
02
b110 6
#610690000000
1!
1%
1-
12
#610700000000
0!
0%
b111 *
0-
02
b111 6
#610710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#610720000000
0!
0%
b0 *
0-
02
b0 6
#610730000000
1!
1%
1-
12
#610740000000
0!
0%
b1 *
0-
02
b1 6
#610750000000
1!
1%
1-
12
#610760000000
0!
0%
b10 *
0-
02
b10 6
#610770000000
1!
1%
1-
12
#610780000000
0!
0%
b11 *
0-
02
b11 6
#610790000000
1!
1%
1-
12
15
#610800000000
0!
0%
b100 *
0-
02
b100 6
#610810000000
1!
1%
1-
12
#610820000000
0!
0%
b101 *
0-
02
b101 6
#610830000000
1!
1%
1-
12
#610840000000
0!
0%
b110 *
0-
02
b110 6
#610850000000
1!
1%
1-
12
#610860000000
0!
0%
b111 *
0-
02
b111 6
#610870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#610880000000
0!
0%
b0 *
0-
02
b0 6
#610890000000
1!
1%
1-
12
#610900000000
0!
0%
b1 *
0-
02
b1 6
#610910000000
1!
1%
1-
12
#610920000000
0!
0%
b10 *
0-
02
b10 6
#610930000000
1!
1%
1-
12
#610940000000
0!
0%
b11 *
0-
02
b11 6
#610950000000
1!
1%
1-
12
15
#610960000000
0!
0%
b100 *
0-
02
b100 6
#610970000000
1!
1%
1-
12
#610980000000
0!
0%
b101 *
0-
02
b101 6
#610990000000
1!
1%
1-
12
#611000000000
0!
0%
b110 *
0-
02
b110 6
#611010000000
1!
1%
1-
12
#611020000000
0!
0%
b111 *
0-
02
b111 6
#611030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#611040000000
0!
0%
b0 *
0-
02
b0 6
#611050000000
1!
1%
1-
12
#611060000000
0!
0%
b1 *
0-
02
b1 6
#611070000000
1!
1%
1-
12
#611080000000
0!
0%
b10 *
0-
02
b10 6
#611090000000
1!
1%
1-
12
#611100000000
0!
0%
b11 *
0-
02
b11 6
#611110000000
1!
1%
1-
12
15
#611120000000
0!
0%
b100 *
0-
02
b100 6
#611130000000
1!
1%
1-
12
#611140000000
0!
0%
b101 *
0-
02
b101 6
#611150000000
1!
1%
1-
12
#611160000000
0!
0%
b110 *
0-
02
b110 6
#611170000000
1!
1%
1-
12
#611180000000
0!
0%
b111 *
0-
02
b111 6
#611190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#611200000000
0!
0%
b0 *
0-
02
b0 6
#611210000000
1!
1%
1-
12
#611220000000
0!
0%
b1 *
0-
02
b1 6
#611230000000
1!
1%
1-
12
#611240000000
0!
0%
b10 *
0-
02
b10 6
#611250000000
1!
1%
1-
12
#611260000000
0!
0%
b11 *
0-
02
b11 6
#611270000000
1!
1%
1-
12
15
#611280000000
0!
0%
b100 *
0-
02
b100 6
#611290000000
1!
1%
1-
12
#611300000000
0!
0%
b101 *
0-
02
b101 6
#611310000000
1!
1%
1-
12
#611320000000
0!
0%
b110 *
0-
02
b110 6
#611330000000
1!
1%
1-
12
#611340000000
0!
0%
b111 *
0-
02
b111 6
#611350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#611360000000
0!
0%
b0 *
0-
02
b0 6
#611370000000
1!
1%
1-
12
#611380000000
0!
0%
b1 *
0-
02
b1 6
#611390000000
1!
1%
1-
12
#611400000000
0!
0%
b10 *
0-
02
b10 6
#611410000000
1!
1%
1-
12
#611420000000
0!
0%
b11 *
0-
02
b11 6
#611430000000
1!
1%
1-
12
15
#611440000000
0!
0%
b100 *
0-
02
b100 6
#611450000000
1!
1%
1-
12
#611460000000
0!
0%
b101 *
0-
02
b101 6
#611470000000
1!
1%
1-
12
#611480000000
0!
0%
b110 *
0-
02
b110 6
#611490000000
1!
1%
1-
12
#611500000000
0!
0%
b111 *
0-
02
b111 6
#611510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#611520000000
0!
0%
b0 *
0-
02
b0 6
#611530000000
1!
1%
1-
12
#611540000000
0!
0%
b1 *
0-
02
b1 6
#611550000000
1!
1%
1-
12
#611560000000
0!
0%
b10 *
0-
02
b10 6
#611570000000
1!
1%
1-
12
#611580000000
0!
0%
b11 *
0-
02
b11 6
#611590000000
1!
1%
1-
12
15
#611600000000
0!
0%
b100 *
0-
02
b100 6
#611610000000
1!
1%
1-
12
#611620000000
0!
0%
b101 *
0-
02
b101 6
#611630000000
1!
1%
1-
12
#611640000000
0!
0%
b110 *
0-
02
b110 6
#611650000000
1!
1%
1-
12
#611660000000
0!
0%
b111 *
0-
02
b111 6
#611670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#611680000000
0!
0%
b0 *
0-
02
b0 6
#611690000000
1!
1%
1-
12
#611700000000
0!
0%
b1 *
0-
02
b1 6
#611710000000
1!
1%
1-
12
#611720000000
0!
0%
b10 *
0-
02
b10 6
#611730000000
1!
1%
1-
12
#611740000000
0!
0%
b11 *
0-
02
b11 6
#611750000000
1!
1%
1-
12
15
#611760000000
0!
0%
b100 *
0-
02
b100 6
#611770000000
1!
1%
1-
12
#611780000000
0!
0%
b101 *
0-
02
b101 6
#611790000000
1!
1%
1-
12
#611800000000
0!
0%
b110 *
0-
02
b110 6
#611810000000
1!
1%
1-
12
#611820000000
0!
0%
b111 *
0-
02
b111 6
#611830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#611840000000
0!
0%
b0 *
0-
02
b0 6
#611850000000
1!
1%
1-
12
#611860000000
0!
0%
b1 *
0-
02
b1 6
#611870000000
1!
1%
1-
12
#611880000000
0!
0%
b10 *
0-
02
b10 6
#611890000000
1!
1%
1-
12
#611900000000
0!
0%
b11 *
0-
02
b11 6
#611910000000
1!
1%
1-
12
15
#611920000000
0!
0%
b100 *
0-
02
b100 6
#611930000000
1!
1%
1-
12
#611940000000
0!
0%
b101 *
0-
02
b101 6
#611950000000
1!
1%
1-
12
#611960000000
0!
0%
b110 *
0-
02
b110 6
#611970000000
1!
1%
1-
12
#611980000000
0!
0%
b111 *
0-
02
b111 6
#611990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#612000000000
0!
0%
b0 *
0-
02
b0 6
#612010000000
1!
1%
1-
12
#612020000000
0!
0%
b1 *
0-
02
b1 6
#612030000000
1!
1%
1-
12
#612040000000
0!
0%
b10 *
0-
02
b10 6
#612050000000
1!
1%
1-
12
#612060000000
0!
0%
b11 *
0-
02
b11 6
#612070000000
1!
1%
1-
12
15
#612080000000
0!
0%
b100 *
0-
02
b100 6
#612090000000
1!
1%
1-
12
#612100000000
0!
0%
b101 *
0-
02
b101 6
#612110000000
1!
1%
1-
12
#612120000000
0!
0%
b110 *
0-
02
b110 6
#612130000000
1!
1%
1-
12
#612140000000
0!
0%
b111 *
0-
02
b111 6
#612150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#612160000000
0!
0%
b0 *
0-
02
b0 6
#612170000000
1!
1%
1-
12
#612180000000
0!
0%
b1 *
0-
02
b1 6
#612190000000
1!
1%
1-
12
#612200000000
0!
0%
b10 *
0-
02
b10 6
#612210000000
1!
1%
1-
12
#612220000000
0!
0%
b11 *
0-
02
b11 6
#612230000000
1!
1%
1-
12
15
#612240000000
0!
0%
b100 *
0-
02
b100 6
#612250000000
1!
1%
1-
12
#612260000000
0!
0%
b101 *
0-
02
b101 6
#612270000000
1!
1%
1-
12
#612280000000
0!
0%
b110 *
0-
02
b110 6
#612290000000
1!
1%
1-
12
#612300000000
0!
0%
b111 *
0-
02
b111 6
#612310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#612320000000
0!
0%
b0 *
0-
02
b0 6
#612330000000
1!
1%
1-
12
#612340000000
0!
0%
b1 *
0-
02
b1 6
#612350000000
1!
1%
1-
12
#612360000000
0!
0%
b10 *
0-
02
b10 6
#612370000000
1!
1%
1-
12
#612380000000
0!
0%
b11 *
0-
02
b11 6
#612390000000
1!
1%
1-
12
15
#612400000000
0!
0%
b100 *
0-
02
b100 6
#612410000000
1!
1%
1-
12
#612420000000
0!
0%
b101 *
0-
02
b101 6
#612430000000
1!
1%
1-
12
#612440000000
0!
0%
b110 *
0-
02
b110 6
#612450000000
1!
1%
1-
12
#612460000000
0!
0%
b111 *
0-
02
b111 6
#612470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#612480000000
0!
0%
b0 *
0-
02
b0 6
#612490000000
1!
1%
1-
12
#612500000000
0!
0%
b1 *
0-
02
b1 6
#612510000000
1!
1%
1-
12
#612520000000
0!
0%
b10 *
0-
02
b10 6
#612530000000
1!
1%
1-
12
#612540000000
0!
0%
b11 *
0-
02
b11 6
#612550000000
1!
1%
1-
12
15
#612560000000
0!
0%
b100 *
0-
02
b100 6
#612570000000
1!
1%
1-
12
#612580000000
0!
0%
b101 *
0-
02
b101 6
#612590000000
1!
1%
1-
12
#612600000000
0!
0%
b110 *
0-
02
b110 6
#612610000000
1!
1%
1-
12
#612620000000
0!
0%
b111 *
0-
02
b111 6
#612630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#612640000000
0!
0%
b0 *
0-
02
b0 6
#612650000000
1!
1%
1-
12
#612660000000
0!
0%
b1 *
0-
02
b1 6
#612670000000
1!
1%
1-
12
#612680000000
0!
0%
b10 *
0-
02
b10 6
#612690000000
1!
1%
1-
12
#612700000000
0!
0%
b11 *
0-
02
b11 6
#612710000000
1!
1%
1-
12
15
#612720000000
0!
0%
b100 *
0-
02
b100 6
#612730000000
1!
1%
1-
12
#612740000000
0!
0%
b101 *
0-
02
b101 6
#612750000000
1!
1%
1-
12
#612760000000
0!
0%
b110 *
0-
02
b110 6
#612770000000
1!
1%
1-
12
#612780000000
0!
0%
b111 *
0-
02
b111 6
#612790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#612800000000
0!
0%
b0 *
0-
02
b0 6
#612810000000
1!
1%
1-
12
#612820000000
0!
0%
b1 *
0-
02
b1 6
#612830000000
1!
1%
1-
12
#612840000000
0!
0%
b10 *
0-
02
b10 6
#612850000000
1!
1%
1-
12
#612860000000
0!
0%
b11 *
0-
02
b11 6
#612870000000
1!
1%
1-
12
15
#612880000000
0!
0%
b100 *
0-
02
b100 6
#612890000000
1!
1%
1-
12
#612900000000
0!
0%
b101 *
0-
02
b101 6
#612910000000
1!
1%
1-
12
#612920000000
0!
0%
b110 *
0-
02
b110 6
#612930000000
1!
1%
1-
12
#612940000000
0!
0%
b111 *
0-
02
b111 6
#612950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#612960000000
0!
0%
b0 *
0-
02
b0 6
#612970000000
1!
1%
1-
12
#612980000000
0!
0%
b1 *
0-
02
b1 6
#612990000000
1!
1%
1-
12
#613000000000
0!
0%
b10 *
0-
02
b10 6
#613010000000
1!
1%
1-
12
#613020000000
0!
0%
b11 *
0-
02
b11 6
#613030000000
1!
1%
1-
12
15
#613040000000
0!
0%
b100 *
0-
02
b100 6
#613050000000
1!
1%
1-
12
#613060000000
0!
0%
b101 *
0-
02
b101 6
#613070000000
1!
1%
1-
12
#613080000000
0!
0%
b110 *
0-
02
b110 6
#613090000000
1!
1%
1-
12
#613100000000
0!
0%
b111 *
0-
02
b111 6
#613110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#613120000000
0!
0%
b0 *
0-
02
b0 6
#613130000000
1!
1%
1-
12
#613140000000
0!
0%
b1 *
0-
02
b1 6
#613150000000
1!
1%
1-
12
#613160000000
0!
0%
b10 *
0-
02
b10 6
#613170000000
1!
1%
1-
12
#613180000000
0!
0%
b11 *
0-
02
b11 6
#613190000000
1!
1%
1-
12
15
#613200000000
0!
0%
b100 *
0-
02
b100 6
#613210000000
1!
1%
1-
12
#613220000000
0!
0%
b101 *
0-
02
b101 6
#613230000000
1!
1%
1-
12
#613240000000
0!
0%
b110 *
0-
02
b110 6
#613250000000
1!
1%
1-
12
#613260000000
0!
0%
b111 *
0-
02
b111 6
#613270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#613280000000
0!
0%
b0 *
0-
02
b0 6
#613290000000
1!
1%
1-
12
#613300000000
0!
0%
b1 *
0-
02
b1 6
#613310000000
1!
1%
1-
12
#613320000000
0!
0%
b10 *
0-
02
b10 6
#613330000000
1!
1%
1-
12
#613340000000
0!
0%
b11 *
0-
02
b11 6
#613350000000
1!
1%
1-
12
15
#613360000000
0!
0%
b100 *
0-
02
b100 6
#613370000000
1!
1%
1-
12
#613380000000
0!
0%
b101 *
0-
02
b101 6
#613390000000
1!
1%
1-
12
#613400000000
0!
0%
b110 *
0-
02
b110 6
#613410000000
1!
1%
1-
12
#613420000000
0!
0%
b111 *
0-
02
b111 6
#613430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#613440000000
0!
0%
b0 *
0-
02
b0 6
#613450000000
1!
1%
1-
12
#613460000000
0!
0%
b1 *
0-
02
b1 6
#613470000000
1!
1%
1-
12
#613480000000
0!
0%
b10 *
0-
02
b10 6
#613490000000
1!
1%
1-
12
#613500000000
0!
0%
b11 *
0-
02
b11 6
#613510000000
1!
1%
1-
12
15
#613520000000
0!
0%
b100 *
0-
02
b100 6
#613530000000
1!
1%
1-
12
#613540000000
0!
0%
b101 *
0-
02
b101 6
#613550000000
1!
1%
1-
12
#613560000000
0!
0%
b110 *
0-
02
b110 6
#613570000000
1!
1%
1-
12
#613580000000
0!
0%
b111 *
0-
02
b111 6
#613590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#613600000000
0!
0%
b0 *
0-
02
b0 6
#613610000000
1!
1%
1-
12
#613620000000
0!
0%
b1 *
0-
02
b1 6
#613630000000
1!
1%
1-
12
#613640000000
0!
0%
b10 *
0-
02
b10 6
#613650000000
1!
1%
1-
12
#613660000000
0!
0%
b11 *
0-
02
b11 6
#613670000000
1!
1%
1-
12
15
#613680000000
0!
0%
b100 *
0-
02
b100 6
#613690000000
1!
1%
1-
12
#613700000000
0!
0%
b101 *
0-
02
b101 6
#613710000000
1!
1%
1-
12
#613720000000
0!
0%
b110 *
0-
02
b110 6
#613730000000
1!
1%
1-
12
#613740000000
0!
0%
b111 *
0-
02
b111 6
#613750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#613760000000
0!
0%
b0 *
0-
02
b0 6
#613770000000
1!
1%
1-
12
#613780000000
0!
0%
b1 *
0-
02
b1 6
#613790000000
1!
1%
1-
12
#613800000000
0!
0%
b10 *
0-
02
b10 6
#613810000000
1!
1%
1-
12
#613820000000
0!
0%
b11 *
0-
02
b11 6
#613830000000
1!
1%
1-
12
15
#613840000000
0!
0%
b100 *
0-
02
b100 6
#613850000000
1!
1%
1-
12
#613860000000
0!
0%
b101 *
0-
02
b101 6
#613870000000
1!
1%
1-
12
#613880000000
0!
0%
b110 *
0-
02
b110 6
#613890000000
1!
1%
1-
12
#613900000000
0!
0%
b111 *
0-
02
b111 6
#613910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#613920000000
0!
0%
b0 *
0-
02
b0 6
#613930000000
1!
1%
1-
12
#613940000000
0!
0%
b1 *
0-
02
b1 6
#613950000000
1!
1%
1-
12
#613960000000
0!
0%
b10 *
0-
02
b10 6
#613970000000
1!
1%
1-
12
#613980000000
0!
0%
b11 *
0-
02
b11 6
#613990000000
1!
1%
1-
12
15
#614000000000
0!
0%
b100 *
0-
02
b100 6
#614010000000
1!
1%
1-
12
#614020000000
0!
0%
b101 *
0-
02
b101 6
#614030000000
1!
1%
1-
12
#614040000000
0!
0%
b110 *
0-
02
b110 6
#614050000000
1!
1%
1-
12
#614060000000
0!
0%
b111 *
0-
02
b111 6
#614070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#614080000000
0!
0%
b0 *
0-
02
b0 6
#614090000000
1!
1%
1-
12
#614100000000
0!
0%
b1 *
0-
02
b1 6
#614110000000
1!
1%
1-
12
#614120000000
0!
0%
b10 *
0-
02
b10 6
#614130000000
1!
1%
1-
12
#614140000000
0!
0%
b11 *
0-
02
b11 6
#614150000000
1!
1%
1-
12
15
#614160000000
0!
0%
b100 *
0-
02
b100 6
#614170000000
1!
1%
1-
12
#614180000000
0!
0%
b101 *
0-
02
b101 6
#614190000000
1!
1%
1-
12
#614200000000
0!
0%
b110 *
0-
02
b110 6
#614210000000
1!
1%
1-
12
#614220000000
0!
0%
b111 *
0-
02
b111 6
#614230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#614240000000
0!
0%
b0 *
0-
02
b0 6
#614250000000
1!
1%
1-
12
#614260000000
0!
0%
b1 *
0-
02
b1 6
#614270000000
1!
1%
1-
12
#614280000000
0!
0%
b10 *
0-
02
b10 6
#614290000000
1!
1%
1-
12
#614300000000
0!
0%
b11 *
0-
02
b11 6
#614310000000
1!
1%
1-
12
15
#614320000000
0!
0%
b100 *
0-
02
b100 6
#614330000000
1!
1%
1-
12
#614340000000
0!
0%
b101 *
0-
02
b101 6
#614350000000
1!
1%
1-
12
#614360000000
0!
0%
b110 *
0-
02
b110 6
#614370000000
1!
1%
1-
12
#614380000000
0!
0%
b111 *
0-
02
b111 6
#614390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#614400000000
0!
0%
b0 *
0-
02
b0 6
#614410000000
1!
1%
1-
12
#614420000000
0!
0%
b1 *
0-
02
b1 6
#614430000000
1!
1%
1-
12
#614440000000
0!
0%
b10 *
0-
02
b10 6
#614450000000
1!
1%
1-
12
#614460000000
0!
0%
b11 *
0-
02
b11 6
#614470000000
1!
1%
1-
12
15
#614480000000
0!
0%
b100 *
0-
02
b100 6
#614490000000
1!
1%
1-
12
#614500000000
0!
0%
b101 *
0-
02
b101 6
#614510000000
1!
1%
1-
12
#614520000000
0!
0%
b110 *
0-
02
b110 6
#614530000000
1!
1%
1-
12
#614540000000
0!
0%
b111 *
0-
02
b111 6
#614550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#614560000000
0!
0%
b0 *
0-
02
b0 6
#614570000000
1!
1%
1-
12
#614580000000
0!
0%
b1 *
0-
02
b1 6
#614590000000
1!
1%
1-
12
#614600000000
0!
0%
b10 *
0-
02
b10 6
#614610000000
1!
1%
1-
12
#614620000000
0!
0%
b11 *
0-
02
b11 6
#614630000000
1!
1%
1-
12
15
#614640000000
0!
0%
b100 *
0-
02
b100 6
#614650000000
1!
1%
1-
12
#614660000000
0!
0%
b101 *
0-
02
b101 6
#614670000000
1!
1%
1-
12
#614680000000
0!
0%
b110 *
0-
02
b110 6
#614690000000
1!
1%
1-
12
#614700000000
0!
0%
b111 *
0-
02
b111 6
#614710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#614720000000
0!
0%
b0 *
0-
02
b0 6
#614730000000
1!
1%
1-
12
#614740000000
0!
0%
b1 *
0-
02
b1 6
#614750000000
1!
1%
1-
12
#614760000000
0!
0%
b10 *
0-
02
b10 6
#614770000000
1!
1%
1-
12
#614780000000
0!
0%
b11 *
0-
02
b11 6
#614790000000
1!
1%
1-
12
15
#614800000000
0!
0%
b100 *
0-
02
b100 6
#614810000000
1!
1%
1-
12
#614820000000
0!
0%
b101 *
0-
02
b101 6
#614830000000
1!
1%
1-
12
#614840000000
0!
0%
b110 *
0-
02
b110 6
#614850000000
1!
1%
1-
12
#614860000000
0!
0%
b111 *
0-
02
b111 6
#614870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#614880000000
0!
0%
b0 *
0-
02
b0 6
#614890000000
1!
1%
1-
12
#614900000000
0!
0%
b1 *
0-
02
b1 6
#614910000000
1!
1%
1-
12
#614920000000
0!
0%
b10 *
0-
02
b10 6
#614930000000
1!
1%
1-
12
#614940000000
0!
0%
b11 *
0-
02
b11 6
#614950000000
1!
1%
1-
12
15
#614960000000
0!
0%
b100 *
0-
02
b100 6
#614970000000
1!
1%
1-
12
#614980000000
0!
0%
b101 *
0-
02
b101 6
#614990000000
1!
1%
1-
12
#615000000000
0!
0%
b110 *
0-
02
b110 6
#615010000000
1!
1%
1-
12
#615020000000
0!
0%
b111 *
0-
02
b111 6
#615030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#615040000000
0!
0%
b0 *
0-
02
b0 6
#615050000000
1!
1%
1-
12
#615060000000
0!
0%
b1 *
0-
02
b1 6
#615070000000
1!
1%
1-
12
#615080000000
0!
0%
b10 *
0-
02
b10 6
#615090000000
1!
1%
1-
12
#615100000000
0!
0%
b11 *
0-
02
b11 6
#615110000000
1!
1%
1-
12
15
#615120000000
0!
0%
b100 *
0-
02
b100 6
#615130000000
1!
1%
1-
12
#615140000000
0!
0%
b101 *
0-
02
b101 6
#615150000000
1!
1%
1-
12
#615160000000
0!
0%
b110 *
0-
02
b110 6
#615170000000
1!
1%
1-
12
#615180000000
0!
0%
b111 *
0-
02
b111 6
#615190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#615200000000
0!
0%
b0 *
0-
02
b0 6
#615210000000
1!
1%
1-
12
#615220000000
0!
0%
b1 *
0-
02
b1 6
#615230000000
1!
1%
1-
12
#615240000000
0!
0%
b10 *
0-
02
b10 6
#615250000000
1!
1%
1-
12
#615260000000
0!
0%
b11 *
0-
02
b11 6
#615270000000
1!
1%
1-
12
15
#615280000000
0!
0%
b100 *
0-
02
b100 6
#615290000000
1!
1%
1-
12
#615300000000
0!
0%
b101 *
0-
02
b101 6
#615310000000
1!
1%
1-
12
#615320000000
0!
0%
b110 *
0-
02
b110 6
#615330000000
1!
1%
1-
12
#615340000000
0!
0%
b111 *
0-
02
b111 6
#615350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#615360000000
0!
0%
b0 *
0-
02
b0 6
#615370000000
1!
1%
1-
12
#615380000000
0!
0%
b1 *
0-
02
b1 6
#615390000000
1!
1%
1-
12
#615400000000
0!
0%
b10 *
0-
02
b10 6
#615410000000
1!
1%
1-
12
#615420000000
0!
0%
b11 *
0-
02
b11 6
#615430000000
1!
1%
1-
12
15
#615440000000
0!
0%
b100 *
0-
02
b100 6
#615450000000
1!
1%
1-
12
#615460000000
0!
0%
b101 *
0-
02
b101 6
#615470000000
1!
1%
1-
12
#615480000000
0!
0%
b110 *
0-
02
b110 6
#615490000000
1!
1%
1-
12
#615500000000
0!
0%
b111 *
0-
02
b111 6
#615510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#615520000000
0!
0%
b0 *
0-
02
b0 6
#615530000000
1!
1%
1-
12
#615540000000
0!
0%
b1 *
0-
02
b1 6
#615550000000
1!
1%
1-
12
#615560000000
0!
0%
b10 *
0-
02
b10 6
#615570000000
1!
1%
1-
12
#615580000000
0!
0%
b11 *
0-
02
b11 6
#615590000000
1!
1%
1-
12
15
#615600000000
0!
0%
b100 *
0-
02
b100 6
#615610000000
1!
1%
1-
12
#615620000000
0!
0%
b101 *
0-
02
b101 6
#615630000000
1!
1%
1-
12
#615640000000
0!
0%
b110 *
0-
02
b110 6
#615650000000
1!
1%
1-
12
#615660000000
0!
0%
b111 *
0-
02
b111 6
#615670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#615680000000
0!
0%
b0 *
0-
02
b0 6
#615690000000
1!
1%
1-
12
#615700000000
0!
0%
b1 *
0-
02
b1 6
#615710000000
1!
1%
1-
12
#615720000000
0!
0%
b10 *
0-
02
b10 6
#615730000000
1!
1%
1-
12
#615740000000
0!
0%
b11 *
0-
02
b11 6
#615750000000
1!
1%
1-
12
15
#615760000000
0!
0%
b100 *
0-
02
b100 6
#615770000000
1!
1%
1-
12
#615780000000
0!
0%
b101 *
0-
02
b101 6
#615790000000
1!
1%
1-
12
#615800000000
0!
0%
b110 *
0-
02
b110 6
#615810000000
1!
1%
1-
12
#615820000000
0!
0%
b111 *
0-
02
b111 6
#615830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#615840000000
0!
0%
b0 *
0-
02
b0 6
#615850000000
1!
1%
1-
12
#615860000000
0!
0%
b1 *
0-
02
b1 6
#615870000000
1!
1%
1-
12
#615880000000
0!
0%
b10 *
0-
02
b10 6
#615890000000
1!
1%
1-
12
#615900000000
0!
0%
b11 *
0-
02
b11 6
#615910000000
1!
1%
1-
12
15
#615920000000
0!
0%
b100 *
0-
02
b100 6
#615930000000
1!
1%
1-
12
#615940000000
0!
0%
b101 *
0-
02
b101 6
#615950000000
1!
1%
1-
12
#615960000000
0!
0%
b110 *
0-
02
b110 6
#615970000000
1!
1%
1-
12
#615980000000
0!
0%
b111 *
0-
02
b111 6
#615990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#616000000000
0!
0%
b0 *
0-
02
b0 6
#616010000000
1!
1%
1-
12
#616020000000
0!
0%
b1 *
0-
02
b1 6
#616030000000
1!
1%
1-
12
#616040000000
0!
0%
b10 *
0-
02
b10 6
#616050000000
1!
1%
1-
12
#616060000000
0!
0%
b11 *
0-
02
b11 6
#616070000000
1!
1%
1-
12
15
#616080000000
0!
0%
b100 *
0-
02
b100 6
#616090000000
1!
1%
1-
12
#616100000000
0!
0%
b101 *
0-
02
b101 6
#616110000000
1!
1%
1-
12
#616120000000
0!
0%
b110 *
0-
02
b110 6
#616130000000
1!
1%
1-
12
#616140000000
0!
0%
b111 *
0-
02
b111 6
#616150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#616160000000
0!
0%
b0 *
0-
02
b0 6
#616170000000
1!
1%
1-
12
#616180000000
0!
0%
b1 *
0-
02
b1 6
#616190000000
1!
1%
1-
12
#616200000000
0!
0%
b10 *
0-
02
b10 6
#616210000000
1!
1%
1-
12
#616220000000
0!
0%
b11 *
0-
02
b11 6
#616230000000
1!
1%
1-
12
15
#616240000000
0!
0%
b100 *
0-
02
b100 6
#616250000000
1!
1%
1-
12
#616260000000
0!
0%
b101 *
0-
02
b101 6
#616270000000
1!
1%
1-
12
#616280000000
0!
0%
b110 *
0-
02
b110 6
#616290000000
1!
1%
1-
12
#616300000000
0!
0%
b111 *
0-
02
b111 6
#616310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#616320000000
0!
0%
b0 *
0-
02
b0 6
#616330000000
1!
1%
1-
12
#616340000000
0!
0%
b1 *
0-
02
b1 6
#616350000000
1!
1%
1-
12
#616360000000
0!
0%
b10 *
0-
02
b10 6
#616370000000
1!
1%
1-
12
#616380000000
0!
0%
b11 *
0-
02
b11 6
#616390000000
1!
1%
1-
12
15
#616400000000
0!
0%
b100 *
0-
02
b100 6
#616410000000
1!
1%
1-
12
#616420000000
0!
0%
b101 *
0-
02
b101 6
#616430000000
1!
1%
1-
12
#616440000000
0!
0%
b110 *
0-
02
b110 6
#616450000000
1!
1%
1-
12
#616460000000
0!
0%
b111 *
0-
02
b111 6
#616470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#616480000000
0!
0%
b0 *
0-
02
b0 6
#616490000000
1!
1%
1-
12
#616500000000
0!
0%
b1 *
0-
02
b1 6
#616510000000
1!
1%
1-
12
#616520000000
0!
0%
b10 *
0-
02
b10 6
#616530000000
1!
1%
1-
12
#616540000000
0!
0%
b11 *
0-
02
b11 6
#616550000000
1!
1%
1-
12
15
#616560000000
0!
0%
b100 *
0-
02
b100 6
#616570000000
1!
1%
1-
12
#616580000000
0!
0%
b101 *
0-
02
b101 6
#616590000000
1!
1%
1-
12
#616600000000
0!
0%
b110 *
0-
02
b110 6
#616610000000
1!
1%
1-
12
#616620000000
0!
0%
b111 *
0-
02
b111 6
#616630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#616640000000
0!
0%
b0 *
0-
02
b0 6
#616650000000
1!
1%
1-
12
#616660000000
0!
0%
b1 *
0-
02
b1 6
#616670000000
1!
1%
1-
12
#616680000000
0!
0%
b10 *
0-
02
b10 6
#616690000000
1!
1%
1-
12
#616700000000
0!
0%
b11 *
0-
02
b11 6
#616710000000
1!
1%
1-
12
15
#616720000000
0!
0%
b100 *
0-
02
b100 6
#616730000000
1!
1%
1-
12
#616740000000
0!
0%
b101 *
0-
02
b101 6
#616750000000
1!
1%
1-
12
#616760000000
0!
0%
b110 *
0-
02
b110 6
#616770000000
1!
1%
1-
12
#616780000000
0!
0%
b111 *
0-
02
b111 6
#616790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#616800000000
0!
0%
b0 *
0-
02
b0 6
#616810000000
1!
1%
1-
12
#616820000000
0!
0%
b1 *
0-
02
b1 6
#616830000000
1!
1%
1-
12
#616840000000
0!
0%
b10 *
0-
02
b10 6
#616850000000
1!
1%
1-
12
#616860000000
0!
0%
b11 *
0-
02
b11 6
#616870000000
1!
1%
1-
12
15
#616880000000
0!
0%
b100 *
0-
02
b100 6
#616890000000
1!
1%
1-
12
#616900000000
0!
0%
b101 *
0-
02
b101 6
#616910000000
1!
1%
1-
12
#616920000000
0!
0%
b110 *
0-
02
b110 6
#616930000000
1!
1%
1-
12
#616940000000
0!
0%
b111 *
0-
02
b111 6
#616950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#616960000000
0!
0%
b0 *
0-
02
b0 6
#616970000000
1!
1%
1-
12
#616980000000
0!
0%
b1 *
0-
02
b1 6
#616990000000
1!
1%
1-
12
#617000000000
0!
0%
b10 *
0-
02
b10 6
#617010000000
1!
1%
1-
12
#617020000000
0!
0%
b11 *
0-
02
b11 6
#617030000000
1!
1%
1-
12
15
#617040000000
0!
0%
b100 *
0-
02
b100 6
#617050000000
1!
1%
1-
12
#617060000000
0!
0%
b101 *
0-
02
b101 6
#617070000000
1!
1%
1-
12
#617080000000
0!
0%
b110 *
0-
02
b110 6
#617090000000
1!
1%
1-
12
#617100000000
0!
0%
b111 *
0-
02
b111 6
#617110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#617120000000
0!
0%
b0 *
0-
02
b0 6
#617130000000
1!
1%
1-
12
#617140000000
0!
0%
b1 *
0-
02
b1 6
#617150000000
1!
1%
1-
12
#617160000000
0!
0%
b10 *
0-
02
b10 6
#617170000000
1!
1%
1-
12
#617180000000
0!
0%
b11 *
0-
02
b11 6
#617190000000
1!
1%
1-
12
15
#617200000000
0!
0%
b100 *
0-
02
b100 6
#617210000000
1!
1%
1-
12
#617220000000
0!
0%
b101 *
0-
02
b101 6
#617230000000
1!
1%
1-
12
#617240000000
0!
0%
b110 *
0-
02
b110 6
#617250000000
1!
1%
1-
12
#617260000000
0!
0%
b111 *
0-
02
b111 6
#617270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#617280000000
0!
0%
b0 *
0-
02
b0 6
#617290000000
1!
1%
1-
12
#617300000000
0!
0%
b1 *
0-
02
b1 6
#617310000000
1!
1%
1-
12
#617320000000
0!
0%
b10 *
0-
02
b10 6
#617330000000
1!
1%
1-
12
#617340000000
0!
0%
b11 *
0-
02
b11 6
#617350000000
1!
1%
1-
12
15
#617360000000
0!
0%
b100 *
0-
02
b100 6
#617370000000
1!
1%
1-
12
#617380000000
0!
0%
b101 *
0-
02
b101 6
#617390000000
1!
1%
1-
12
#617400000000
0!
0%
b110 *
0-
02
b110 6
#617410000000
1!
1%
1-
12
#617420000000
0!
0%
b111 *
0-
02
b111 6
#617430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#617440000000
0!
0%
b0 *
0-
02
b0 6
#617450000000
1!
1%
1-
12
#617460000000
0!
0%
b1 *
0-
02
b1 6
#617470000000
1!
1%
1-
12
#617480000000
0!
0%
b10 *
0-
02
b10 6
#617490000000
1!
1%
1-
12
#617500000000
0!
0%
b11 *
0-
02
b11 6
#617510000000
1!
1%
1-
12
15
#617520000000
0!
0%
b100 *
0-
02
b100 6
#617530000000
1!
1%
1-
12
#617540000000
0!
0%
b101 *
0-
02
b101 6
#617550000000
1!
1%
1-
12
#617560000000
0!
0%
b110 *
0-
02
b110 6
#617570000000
1!
1%
1-
12
#617580000000
0!
0%
b111 *
0-
02
b111 6
#617590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#617600000000
0!
0%
b0 *
0-
02
b0 6
#617610000000
1!
1%
1-
12
#617620000000
0!
0%
b1 *
0-
02
b1 6
#617630000000
1!
1%
1-
12
#617640000000
0!
0%
b10 *
0-
02
b10 6
#617650000000
1!
1%
1-
12
#617660000000
0!
0%
b11 *
0-
02
b11 6
#617670000000
1!
1%
1-
12
15
#617680000000
0!
0%
b100 *
0-
02
b100 6
#617690000000
1!
1%
1-
12
#617700000000
0!
0%
b101 *
0-
02
b101 6
#617710000000
1!
1%
1-
12
#617720000000
0!
0%
b110 *
0-
02
b110 6
#617730000000
1!
1%
1-
12
#617740000000
0!
0%
b111 *
0-
02
b111 6
#617750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#617760000000
0!
0%
b0 *
0-
02
b0 6
#617770000000
1!
1%
1-
12
#617780000000
0!
0%
b1 *
0-
02
b1 6
#617790000000
1!
1%
1-
12
#617800000000
0!
0%
b10 *
0-
02
b10 6
#617810000000
1!
1%
1-
12
#617820000000
0!
0%
b11 *
0-
02
b11 6
#617830000000
1!
1%
1-
12
15
#617840000000
0!
0%
b100 *
0-
02
b100 6
#617850000000
1!
1%
1-
12
#617860000000
0!
0%
b101 *
0-
02
b101 6
#617870000000
1!
1%
1-
12
#617880000000
0!
0%
b110 *
0-
02
b110 6
#617890000000
1!
1%
1-
12
#617900000000
0!
0%
b111 *
0-
02
b111 6
#617910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#617920000000
0!
0%
b0 *
0-
02
b0 6
#617930000000
1!
1%
1-
12
#617940000000
0!
0%
b1 *
0-
02
b1 6
#617950000000
1!
1%
1-
12
#617960000000
0!
0%
b10 *
0-
02
b10 6
#617970000000
1!
1%
1-
12
#617980000000
0!
0%
b11 *
0-
02
b11 6
#617990000000
1!
1%
1-
12
15
#618000000000
0!
0%
b100 *
0-
02
b100 6
#618010000000
1!
1%
1-
12
#618020000000
0!
0%
b101 *
0-
02
b101 6
#618030000000
1!
1%
1-
12
#618040000000
0!
0%
b110 *
0-
02
b110 6
#618050000000
1!
1%
1-
12
#618060000000
0!
0%
b111 *
0-
02
b111 6
#618070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#618080000000
0!
0%
b0 *
0-
02
b0 6
#618090000000
1!
1%
1-
12
#618100000000
0!
0%
b1 *
0-
02
b1 6
#618110000000
1!
1%
1-
12
#618120000000
0!
0%
b10 *
0-
02
b10 6
#618130000000
1!
1%
1-
12
#618140000000
0!
0%
b11 *
0-
02
b11 6
#618150000000
1!
1%
1-
12
15
#618160000000
0!
0%
b100 *
0-
02
b100 6
#618170000000
1!
1%
1-
12
#618180000000
0!
0%
b101 *
0-
02
b101 6
#618190000000
1!
1%
1-
12
#618200000000
0!
0%
b110 *
0-
02
b110 6
#618210000000
1!
1%
1-
12
#618220000000
0!
0%
b111 *
0-
02
b111 6
#618230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#618240000000
0!
0%
b0 *
0-
02
b0 6
#618250000000
1!
1%
1-
12
#618260000000
0!
0%
b1 *
0-
02
b1 6
#618270000000
1!
1%
1-
12
#618280000000
0!
0%
b10 *
0-
02
b10 6
#618290000000
1!
1%
1-
12
#618300000000
0!
0%
b11 *
0-
02
b11 6
#618310000000
1!
1%
1-
12
15
#618320000000
0!
0%
b100 *
0-
02
b100 6
#618330000000
1!
1%
1-
12
#618340000000
0!
0%
b101 *
0-
02
b101 6
#618350000000
1!
1%
1-
12
#618360000000
0!
0%
b110 *
0-
02
b110 6
#618370000000
1!
1%
1-
12
#618380000000
0!
0%
b111 *
0-
02
b111 6
#618390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#618400000000
0!
0%
b0 *
0-
02
b0 6
#618410000000
1!
1%
1-
12
#618420000000
0!
0%
b1 *
0-
02
b1 6
#618430000000
1!
1%
1-
12
#618440000000
0!
0%
b10 *
0-
02
b10 6
#618450000000
1!
1%
1-
12
#618460000000
0!
0%
b11 *
0-
02
b11 6
#618470000000
1!
1%
1-
12
15
#618480000000
0!
0%
b100 *
0-
02
b100 6
#618490000000
1!
1%
1-
12
#618500000000
0!
0%
b101 *
0-
02
b101 6
#618510000000
1!
1%
1-
12
#618520000000
0!
0%
b110 *
0-
02
b110 6
#618530000000
1!
1%
1-
12
#618540000000
0!
0%
b111 *
0-
02
b111 6
#618550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#618560000000
0!
0%
b0 *
0-
02
b0 6
#618570000000
1!
1%
1-
12
#618580000000
0!
0%
b1 *
0-
02
b1 6
#618590000000
1!
1%
1-
12
#618600000000
0!
0%
b10 *
0-
02
b10 6
#618610000000
1!
1%
1-
12
#618620000000
0!
0%
b11 *
0-
02
b11 6
#618630000000
1!
1%
1-
12
15
#618640000000
0!
0%
b100 *
0-
02
b100 6
#618650000000
1!
1%
1-
12
#618660000000
0!
0%
b101 *
0-
02
b101 6
#618670000000
1!
1%
1-
12
#618680000000
0!
0%
b110 *
0-
02
b110 6
#618690000000
1!
1%
1-
12
#618700000000
0!
0%
b111 *
0-
02
b111 6
#618710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#618720000000
0!
0%
b0 *
0-
02
b0 6
#618730000000
1!
1%
1-
12
#618740000000
0!
0%
b1 *
0-
02
b1 6
#618750000000
1!
1%
1-
12
#618760000000
0!
0%
b10 *
0-
02
b10 6
#618770000000
1!
1%
1-
12
#618780000000
0!
0%
b11 *
0-
02
b11 6
#618790000000
1!
1%
1-
12
15
#618800000000
0!
0%
b100 *
0-
02
b100 6
#618810000000
1!
1%
1-
12
#618820000000
0!
0%
b101 *
0-
02
b101 6
#618830000000
1!
1%
1-
12
#618840000000
0!
0%
b110 *
0-
02
b110 6
#618850000000
1!
1%
1-
12
#618860000000
0!
0%
b111 *
0-
02
b111 6
#618870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#618880000000
0!
0%
b0 *
0-
02
b0 6
#618890000000
1!
1%
1-
12
#618900000000
0!
0%
b1 *
0-
02
b1 6
#618910000000
1!
1%
1-
12
#618920000000
0!
0%
b10 *
0-
02
b10 6
#618930000000
1!
1%
1-
12
#618940000000
0!
0%
b11 *
0-
02
b11 6
#618950000000
1!
1%
1-
12
15
#618960000000
0!
0%
b100 *
0-
02
b100 6
#618970000000
1!
1%
1-
12
#618980000000
0!
0%
b101 *
0-
02
b101 6
#618990000000
1!
1%
1-
12
#619000000000
0!
0%
b110 *
0-
02
b110 6
#619010000000
1!
1%
1-
12
#619020000000
0!
0%
b111 *
0-
02
b111 6
#619030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#619040000000
0!
0%
b0 *
0-
02
b0 6
#619050000000
1!
1%
1-
12
#619060000000
0!
0%
b1 *
0-
02
b1 6
#619070000000
1!
1%
1-
12
#619080000000
0!
0%
b10 *
0-
02
b10 6
#619090000000
1!
1%
1-
12
#619100000000
0!
0%
b11 *
0-
02
b11 6
#619110000000
1!
1%
1-
12
15
#619120000000
0!
0%
b100 *
0-
02
b100 6
#619130000000
1!
1%
1-
12
#619140000000
0!
0%
b101 *
0-
02
b101 6
#619150000000
1!
1%
1-
12
#619160000000
0!
0%
b110 *
0-
02
b110 6
#619170000000
1!
1%
1-
12
#619180000000
0!
0%
b111 *
0-
02
b111 6
#619190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#619200000000
0!
0%
b0 *
0-
02
b0 6
#619210000000
1!
1%
1-
12
#619220000000
0!
0%
b1 *
0-
02
b1 6
#619230000000
1!
1%
1-
12
#619240000000
0!
0%
b10 *
0-
02
b10 6
#619250000000
1!
1%
1-
12
#619260000000
0!
0%
b11 *
0-
02
b11 6
#619270000000
1!
1%
1-
12
15
#619280000000
0!
0%
b100 *
0-
02
b100 6
#619290000000
1!
1%
1-
12
#619300000000
0!
0%
b101 *
0-
02
b101 6
#619310000000
1!
1%
1-
12
#619320000000
0!
0%
b110 *
0-
02
b110 6
#619330000000
1!
1%
1-
12
#619340000000
0!
0%
b111 *
0-
02
b111 6
#619350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#619360000000
0!
0%
b0 *
0-
02
b0 6
#619370000000
1!
1%
1-
12
#619380000000
0!
0%
b1 *
0-
02
b1 6
#619390000000
1!
1%
1-
12
#619400000000
0!
0%
b10 *
0-
02
b10 6
#619410000000
1!
1%
1-
12
#619420000000
0!
0%
b11 *
0-
02
b11 6
#619430000000
1!
1%
1-
12
15
#619440000000
0!
0%
b100 *
0-
02
b100 6
#619450000000
1!
1%
1-
12
#619460000000
0!
0%
b101 *
0-
02
b101 6
#619470000000
1!
1%
1-
12
#619480000000
0!
0%
b110 *
0-
02
b110 6
#619490000000
1!
1%
1-
12
#619500000000
0!
0%
b111 *
0-
02
b111 6
#619510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#619520000000
0!
0%
b0 *
0-
02
b0 6
#619530000000
1!
1%
1-
12
#619540000000
0!
0%
b1 *
0-
02
b1 6
#619550000000
1!
1%
1-
12
#619560000000
0!
0%
b10 *
0-
02
b10 6
#619570000000
1!
1%
1-
12
#619580000000
0!
0%
b11 *
0-
02
b11 6
#619590000000
1!
1%
1-
12
15
#619600000000
0!
0%
b100 *
0-
02
b100 6
#619610000000
1!
1%
1-
12
#619620000000
0!
0%
b101 *
0-
02
b101 6
#619630000000
1!
1%
1-
12
#619640000000
0!
0%
b110 *
0-
02
b110 6
#619650000000
1!
1%
1-
12
#619660000000
0!
0%
b111 *
0-
02
b111 6
#619670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#619680000000
0!
0%
b0 *
0-
02
b0 6
#619690000000
1!
1%
1-
12
#619700000000
0!
0%
b1 *
0-
02
b1 6
#619710000000
1!
1%
1-
12
#619720000000
0!
0%
b10 *
0-
02
b10 6
#619730000000
1!
1%
1-
12
#619740000000
0!
0%
b11 *
0-
02
b11 6
#619750000000
1!
1%
1-
12
15
#619760000000
0!
0%
b100 *
0-
02
b100 6
#619770000000
1!
1%
1-
12
#619780000000
0!
0%
b101 *
0-
02
b101 6
#619790000000
1!
1%
1-
12
#619800000000
0!
0%
b110 *
0-
02
b110 6
#619810000000
1!
1%
1-
12
#619820000000
0!
0%
b111 *
0-
02
b111 6
#619830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#619840000000
0!
0%
b0 *
0-
02
b0 6
#619850000000
1!
1%
1-
12
#619860000000
0!
0%
b1 *
0-
02
b1 6
#619870000000
1!
1%
1-
12
#619880000000
0!
0%
b10 *
0-
02
b10 6
#619890000000
1!
1%
1-
12
#619900000000
0!
0%
b11 *
0-
02
b11 6
#619910000000
1!
1%
1-
12
15
#619920000000
0!
0%
b100 *
0-
02
b100 6
#619930000000
1!
1%
1-
12
#619940000000
0!
0%
b101 *
0-
02
b101 6
#619950000000
1!
1%
1-
12
#619960000000
0!
0%
b110 *
0-
02
b110 6
#619970000000
1!
1%
1-
12
#619980000000
0!
0%
b111 *
0-
02
b111 6
#619990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#620000000000
0!
0%
b0 *
0-
02
b0 6
#620010000000
1!
1%
1-
12
#620020000000
0!
0%
b1 *
0-
02
b1 6
#620030000000
1!
1%
1-
12
#620040000000
0!
0%
b10 *
0-
02
b10 6
#620050000000
1!
1%
1-
12
#620060000000
0!
0%
b11 *
0-
02
b11 6
#620070000000
1!
1%
1-
12
15
#620080000000
0!
0%
b100 *
0-
02
b100 6
#620090000000
1!
1%
1-
12
#620100000000
0!
0%
b101 *
0-
02
b101 6
#620110000000
1!
1%
1-
12
#620120000000
0!
0%
b110 *
0-
02
b110 6
#620130000000
1!
1%
1-
12
#620140000000
0!
0%
b111 *
0-
02
b111 6
#620150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#620160000000
0!
0%
b0 *
0-
02
b0 6
#620170000000
1!
1%
1-
12
#620180000000
0!
0%
b1 *
0-
02
b1 6
#620190000000
1!
1%
1-
12
#620200000000
0!
0%
b10 *
0-
02
b10 6
#620210000000
1!
1%
1-
12
#620220000000
0!
0%
b11 *
0-
02
b11 6
#620230000000
1!
1%
1-
12
15
#620240000000
0!
0%
b100 *
0-
02
b100 6
#620250000000
1!
1%
1-
12
#620260000000
0!
0%
b101 *
0-
02
b101 6
#620270000000
1!
1%
1-
12
#620280000000
0!
0%
b110 *
0-
02
b110 6
#620290000000
1!
1%
1-
12
#620300000000
0!
0%
b111 *
0-
02
b111 6
#620310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#620320000000
0!
0%
b0 *
0-
02
b0 6
#620330000000
1!
1%
1-
12
#620340000000
0!
0%
b1 *
0-
02
b1 6
#620350000000
1!
1%
1-
12
#620360000000
0!
0%
b10 *
0-
02
b10 6
#620370000000
1!
1%
1-
12
#620380000000
0!
0%
b11 *
0-
02
b11 6
#620390000000
1!
1%
1-
12
15
#620400000000
0!
0%
b100 *
0-
02
b100 6
#620410000000
1!
1%
1-
12
#620420000000
0!
0%
b101 *
0-
02
b101 6
#620430000000
1!
1%
1-
12
#620440000000
0!
0%
b110 *
0-
02
b110 6
#620450000000
1!
1%
1-
12
#620460000000
0!
0%
b111 *
0-
02
b111 6
#620470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#620480000000
0!
0%
b0 *
0-
02
b0 6
#620490000000
1!
1%
1-
12
#620500000000
0!
0%
b1 *
0-
02
b1 6
#620510000000
1!
1%
1-
12
#620520000000
0!
0%
b10 *
0-
02
b10 6
#620530000000
1!
1%
1-
12
#620540000000
0!
0%
b11 *
0-
02
b11 6
#620550000000
1!
1%
1-
12
15
#620560000000
0!
0%
b100 *
0-
02
b100 6
#620570000000
1!
1%
1-
12
#620580000000
0!
0%
b101 *
0-
02
b101 6
#620590000000
1!
1%
1-
12
#620600000000
0!
0%
b110 *
0-
02
b110 6
#620610000000
1!
1%
1-
12
#620620000000
0!
0%
b111 *
0-
02
b111 6
#620630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#620640000000
0!
0%
b0 *
0-
02
b0 6
#620650000000
1!
1%
1-
12
#620660000000
0!
0%
b1 *
0-
02
b1 6
#620670000000
1!
1%
1-
12
#620680000000
0!
0%
b10 *
0-
02
b10 6
#620690000000
1!
1%
1-
12
#620700000000
0!
0%
b11 *
0-
02
b11 6
#620710000000
1!
1%
1-
12
15
#620720000000
0!
0%
b100 *
0-
02
b100 6
#620730000000
1!
1%
1-
12
#620740000000
0!
0%
b101 *
0-
02
b101 6
#620750000000
1!
1%
1-
12
#620760000000
0!
0%
b110 *
0-
02
b110 6
#620770000000
1!
1%
1-
12
#620780000000
0!
0%
b111 *
0-
02
b111 6
#620790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#620800000000
0!
0%
b0 *
0-
02
b0 6
#620810000000
1!
1%
1-
12
#620820000000
0!
0%
b1 *
0-
02
b1 6
#620830000000
1!
1%
1-
12
#620840000000
0!
0%
b10 *
0-
02
b10 6
#620850000000
1!
1%
1-
12
#620860000000
0!
0%
b11 *
0-
02
b11 6
#620870000000
1!
1%
1-
12
15
#620880000000
0!
0%
b100 *
0-
02
b100 6
#620890000000
1!
1%
1-
12
#620900000000
0!
0%
b101 *
0-
02
b101 6
#620910000000
1!
1%
1-
12
#620920000000
0!
0%
b110 *
0-
02
b110 6
#620930000000
1!
1%
1-
12
#620940000000
0!
0%
b111 *
0-
02
b111 6
#620950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#620960000000
0!
0%
b0 *
0-
02
b0 6
#620970000000
1!
1%
1-
12
#620980000000
0!
0%
b1 *
0-
02
b1 6
#620990000000
1!
1%
1-
12
#621000000000
0!
0%
b10 *
0-
02
b10 6
#621010000000
1!
1%
1-
12
#621020000000
0!
0%
b11 *
0-
02
b11 6
#621030000000
1!
1%
1-
12
15
#621040000000
0!
0%
b100 *
0-
02
b100 6
#621050000000
1!
1%
1-
12
#621060000000
0!
0%
b101 *
0-
02
b101 6
#621070000000
1!
1%
1-
12
#621080000000
0!
0%
b110 *
0-
02
b110 6
#621090000000
1!
1%
1-
12
#621100000000
0!
0%
b111 *
0-
02
b111 6
#621110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#621120000000
0!
0%
b0 *
0-
02
b0 6
#621130000000
1!
1%
1-
12
#621140000000
0!
0%
b1 *
0-
02
b1 6
#621150000000
1!
1%
1-
12
#621160000000
0!
0%
b10 *
0-
02
b10 6
#621170000000
1!
1%
1-
12
#621180000000
0!
0%
b11 *
0-
02
b11 6
#621190000000
1!
1%
1-
12
15
#621200000000
0!
0%
b100 *
0-
02
b100 6
#621210000000
1!
1%
1-
12
#621220000000
0!
0%
b101 *
0-
02
b101 6
#621230000000
1!
1%
1-
12
#621240000000
0!
0%
b110 *
0-
02
b110 6
#621250000000
1!
1%
1-
12
#621260000000
0!
0%
b111 *
0-
02
b111 6
#621270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#621280000000
0!
0%
b0 *
0-
02
b0 6
#621290000000
1!
1%
1-
12
#621300000000
0!
0%
b1 *
0-
02
b1 6
#621310000000
1!
1%
1-
12
#621320000000
0!
0%
b10 *
0-
02
b10 6
#621330000000
1!
1%
1-
12
#621340000000
0!
0%
b11 *
0-
02
b11 6
#621350000000
1!
1%
1-
12
15
#621360000000
0!
0%
b100 *
0-
02
b100 6
#621370000000
1!
1%
1-
12
#621380000000
0!
0%
b101 *
0-
02
b101 6
#621390000000
1!
1%
1-
12
#621400000000
0!
0%
b110 *
0-
02
b110 6
#621410000000
1!
1%
1-
12
#621420000000
0!
0%
b111 *
0-
02
b111 6
#621430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#621440000000
0!
0%
b0 *
0-
02
b0 6
#621450000000
1!
1%
1-
12
#621460000000
0!
0%
b1 *
0-
02
b1 6
#621470000000
1!
1%
1-
12
#621480000000
0!
0%
b10 *
0-
02
b10 6
#621490000000
1!
1%
1-
12
#621500000000
0!
0%
b11 *
0-
02
b11 6
#621510000000
1!
1%
1-
12
15
#621520000000
0!
0%
b100 *
0-
02
b100 6
#621530000000
1!
1%
1-
12
#621540000000
0!
0%
b101 *
0-
02
b101 6
#621550000000
1!
1%
1-
12
#621560000000
0!
0%
b110 *
0-
02
b110 6
#621570000000
1!
1%
1-
12
#621580000000
0!
0%
b111 *
0-
02
b111 6
#621590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#621600000000
0!
0%
b0 *
0-
02
b0 6
#621610000000
1!
1%
1-
12
#621620000000
0!
0%
b1 *
0-
02
b1 6
#621630000000
1!
1%
1-
12
#621640000000
0!
0%
b10 *
0-
02
b10 6
#621650000000
1!
1%
1-
12
#621660000000
0!
0%
b11 *
0-
02
b11 6
#621670000000
1!
1%
1-
12
15
#621680000000
0!
0%
b100 *
0-
02
b100 6
#621690000000
1!
1%
1-
12
#621700000000
0!
0%
b101 *
0-
02
b101 6
#621710000000
1!
1%
1-
12
#621720000000
0!
0%
b110 *
0-
02
b110 6
#621730000000
1!
1%
1-
12
#621740000000
0!
0%
b111 *
0-
02
b111 6
#621750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#621760000000
0!
0%
b0 *
0-
02
b0 6
#621770000000
1!
1%
1-
12
#621780000000
0!
0%
b1 *
0-
02
b1 6
#621790000000
1!
1%
1-
12
#621800000000
0!
0%
b10 *
0-
02
b10 6
#621810000000
1!
1%
1-
12
#621820000000
0!
0%
b11 *
0-
02
b11 6
#621830000000
1!
1%
1-
12
15
#621840000000
0!
0%
b100 *
0-
02
b100 6
#621850000000
1!
1%
1-
12
#621860000000
0!
0%
b101 *
0-
02
b101 6
#621870000000
1!
1%
1-
12
#621880000000
0!
0%
b110 *
0-
02
b110 6
#621890000000
1!
1%
1-
12
#621900000000
0!
0%
b111 *
0-
02
b111 6
#621910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#621920000000
0!
0%
b0 *
0-
02
b0 6
#621930000000
1!
1%
1-
12
#621940000000
0!
0%
b1 *
0-
02
b1 6
#621950000000
1!
1%
1-
12
#621960000000
0!
0%
b10 *
0-
02
b10 6
#621970000000
1!
1%
1-
12
#621980000000
0!
0%
b11 *
0-
02
b11 6
#621990000000
1!
1%
1-
12
15
#622000000000
0!
0%
b100 *
0-
02
b100 6
#622010000000
1!
1%
1-
12
#622020000000
0!
0%
b101 *
0-
02
b101 6
#622030000000
1!
1%
1-
12
#622040000000
0!
0%
b110 *
0-
02
b110 6
#622050000000
1!
1%
1-
12
#622060000000
0!
0%
b111 *
0-
02
b111 6
#622070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#622080000000
0!
0%
b0 *
0-
02
b0 6
#622090000000
1!
1%
1-
12
#622100000000
0!
0%
b1 *
0-
02
b1 6
#622110000000
1!
1%
1-
12
#622120000000
0!
0%
b10 *
0-
02
b10 6
#622130000000
1!
1%
1-
12
#622140000000
0!
0%
b11 *
0-
02
b11 6
#622150000000
1!
1%
1-
12
15
#622160000000
0!
0%
b100 *
0-
02
b100 6
#622170000000
1!
1%
1-
12
#622180000000
0!
0%
b101 *
0-
02
b101 6
#622190000000
1!
1%
1-
12
#622200000000
0!
0%
b110 *
0-
02
b110 6
#622210000000
1!
1%
1-
12
#622220000000
0!
0%
b111 *
0-
02
b111 6
#622230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#622240000000
0!
0%
b0 *
0-
02
b0 6
#622250000000
1!
1%
1-
12
#622260000000
0!
0%
b1 *
0-
02
b1 6
#622270000000
1!
1%
1-
12
#622280000000
0!
0%
b10 *
0-
02
b10 6
#622290000000
1!
1%
1-
12
#622300000000
0!
0%
b11 *
0-
02
b11 6
#622310000000
1!
1%
1-
12
15
#622320000000
0!
0%
b100 *
0-
02
b100 6
#622330000000
1!
1%
1-
12
#622340000000
0!
0%
b101 *
0-
02
b101 6
#622350000000
1!
1%
1-
12
#622360000000
0!
0%
b110 *
0-
02
b110 6
#622370000000
1!
1%
1-
12
#622380000000
0!
0%
b111 *
0-
02
b111 6
#622390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#622400000000
0!
0%
b0 *
0-
02
b0 6
#622410000000
1!
1%
1-
12
#622420000000
0!
0%
b1 *
0-
02
b1 6
#622430000000
1!
1%
1-
12
#622440000000
0!
0%
b10 *
0-
02
b10 6
#622450000000
1!
1%
1-
12
#622460000000
0!
0%
b11 *
0-
02
b11 6
#622470000000
1!
1%
1-
12
15
#622480000000
0!
0%
b100 *
0-
02
b100 6
#622490000000
1!
1%
1-
12
#622500000000
0!
0%
b101 *
0-
02
b101 6
#622510000000
1!
1%
1-
12
#622520000000
0!
0%
b110 *
0-
02
b110 6
#622530000000
1!
1%
1-
12
#622540000000
0!
0%
b111 *
0-
02
b111 6
#622550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#622560000000
0!
0%
b0 *
0-
02
b0 6
#622570000000
1!
1%
1-
12
#622580000000
0!
0%
b1 *
0-
02
b1 6
#622590000000
1!
1%
1-
12
#622600000000
0!
0%
b10 *
0-
02
b10 6
#622610000000
1!
1%
1-
12
#622620000000
0!
0%
b11 *
0-
02
b11 6
#622630000000
1!
1%
1-
12
15
#622640000000
0!
0%
b100 *
0-
02
b100 6
#622650000000
1!
1%
1-
12
#622660000000
0!
0%
b101 *
0-
02
b101 6
#622670000000
1!
1%
1-
12
#622680000000
0!
0%
b110 *
0-
02
b110 6
#622690000000
1!
1%
1-
12
#622700000000
0!
0%
b111 *
0-
02
b111 6
#622710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#622720000000
0!
0%
b0 *
0-
02
b0 6
#622730000000
1!
1%
1-
12
#622740000000
0!
0%
b1 *
0-
02
b1 6
#622750000000
1!
1%
1-
12
#622760000000
0!
0%
b10 *
0-
02
b10 6
#622770000000
1!
1%
1-
12
#622780000000
0!
0%
b11 *
0-
02
b11 6
#622790000000
1!
1%
1-
12
15
#622800000000
0!
0%
b100 *
0-
02
b100 6
#622810000000
1!
1%
1-
12
#622820000000
0!
0%
b101 *
0-
02
b101 6
#622830000000
1!
1%
1-
12
#622840000000
0!
0%
b110 *
0-
02
b110 6
#622850000000
1!
1%
1-
12
#622860000000
0!
0%
b111 *
0-
02
b111 6
#622870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#622880000000
0!
0%
b0 *
0-
02
b0 6
#622890000000
1!
1%
1-
12
#622900000000
0!
0%
b1 *
0-
02
b1 6
#622910000000
1!
1%
1-
12
#622920000000
0!
0%
b10 *
0-
02
b10 6
#622930000000
1!
1%
1-
12
#622940000000
0!
0%
b11 *
0-
02
b11 6
#622950000000
1!
1%
1-
12
15
#622960000000
0!
0%
b100 *
0-
02
b100 6
#622970000000
1!
1%
1-
12
#622980000000
0!
0%
b101 *
0-
02
b101 6
#622990000000
1!
1%
1-
12
#623000000000
0!
0%
b110 *
0-
02
b110 6
#623010000000
1!
1%
1-
12
#623020000000
0!
0%
b111 *
0-
02
b111 6
#623030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#623040000000
0!
0%
b0 *
0-
02
b0 6
#623050000000
1!
1%
1-
12
#623060000000
0!
0%
b1 *
0-
02
b1 6
#623070000000
1!
1%
1-
12
#623080000000
0!
0%
b10 *
0-
02
b10 6
#623090000000
1!
1%
1-
12
#623100000000
0!
0%
b11 *
0-
02
b11 6
#623110000000
1!
1%
1-
12
15
#623120000000
0!
0%
b100 *
0-
02
b100 6
#623130000000
1!
1%
1-
12
#623140000000
0!
0%
b101 *
0-
02
b101 6
#623150000000
1!
1%
1-
12
#623160000000
0!
0%
b110 *
0-
02
b110 6
#623170000000
1!
1%
1-
12
#623180000000
0!
0%
b111 *
0-
02
b111 6
#623190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#623200000000
0!
0%
b0 *
0-
02
b0 6
#623210000000
1!
1%
1-
12
#623220000000
0!
0%
b1 *
0-
02
b1 6
#623230000000
1!
1%
1-
12
#623240000000
0!
0%
b10 *
0-
02
b10 6
#623250000000
1!
1%
1-
12
#623260000000
0!
0%
b11 *
0-
02
b11 6
#623270000000
1!
1%
1-
12
15
#623280000000
0!
0%
b100 *
0-
02
b100 6
#623290000000
1!
1%
1-
12
#623300000000
0!
0%
b101 *
0-
02
b101 6
#623310000000
1!
1%
1-
12
#623320000000
0!
0%
b110 *
0-
02
b110 6
#623330000000
1!
1%
1-
12
#623340000000
0!
0%
b111 *
0-
02
b111 6
#623350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#623360000000
0!
0%
b0 *
0-
02
b0 6
#623370000000
1!
1%
1-
12
#623380000000
0!
0%
b1 *
0-
02
b1 6
#623390000000
1!
1%
1-
12
#623400000000
0!
0%
b10 *
0-
02
b10 6
#623410000000
1!
1%
1-
12
#623420000000
0!
0%
b11 *
0-
02
b11 6
#623430000000
1!
1%
1-
12
15
#623440000000
0!
0%
b100 *
0-
02
b100 6
#623450000000
1!
1%
1-
12
#623460000000
0!
0%
b101 *
0-
02
b101 6
#623470000000
1!
1%
1-
12
#623480000000
0!
0%
b110 *
0-
02
b110 6
#623490000000
1!
1%
1-
12
#623500000000
0!
0%
b111 *
0-
02
b111 6
#623510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#623520000000
0!
0%
b0 *
0-
02
b0 6
#623530000000
1!
1%
1-
12
#623540000000
0!
0%
b1 *
0-
02
b1 6
#623550000000
1!
1%
1-
12
#623560000000
0!
0%
b10 *
0-
02
b10 6
#623570000000
1!
1%
1-
12
#623580000000
0!
0%
b11 *
0-
02
b11 6
#623590000000
1!
1%
1-
12
15
#623600000000
0!
0%
b100 *
0-
02
b100 6
#623610000000
1!
1%
1-
12
#623620000000
0!
0%
b101 *
0-
02
b101 6
#623630000000
1!
1%
1-
12
#623640000000
0!
0%
b110 *
0-
02
b110 6
#623650000000
1!
1%
1-
12
#623660000000
0!
0%
b111 *
0-
02
b111 6
#623670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#623680000000
0!
0%
b0 *
0-
02
b0 6
#623690000000
1!
1%
1-
12
#623700000000
0!
0%
b1 *
0-
02
b1 6
#623710000000
1!
1%
1-
12
#623720000000
0!
0%
b10 *
0-
02
b10 6
#623730000000
1!
1%
1-
12
#623740000000
0!
0%
b11 *
0-
02
b11 6
#623750000000
1!
1%
1-
12
15
#623760000000
0!
0%
b100 *
0-
02
b100 6
#623770000000
1!
1%
1-
12
#623780000000
0!
0%
b101 *
0-
02
b101 6
#623790000000
1!
1%
1-
12
#623800000000
0!
0%
b110 *
0-
02
b110 6
#623810000000
1!
1%
1-
12
#623820000000
0!
0%
b111 *
0-
02
b111 6
#623830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#623840000000
0!
0%
b0 *
0-
02
b0 6
#623850000000
1!
1%
1-
12
#623860000000
0!
0%
b1 *
0-
02
b1 6
#623870000000
1!
1%
1-
12
#623880000000
0!
0%
b10 *
0-
02
b10 6
#623890000000
1!
1%
1-
12
#623900000000
0!
0%
b11 *
0-
02
b11 6
#623910000000
1!
1%
1-
12
15
#623920000000
0!
0%
b100 *
0-
02
b100 6
#623930000000
1!
1%
1-
12
#623940000000
0!
0%
b101 *
0-
02
b101 6
#623950000000
1!
1%
1-
12
#623960000000
0!
0%
b110 *
0-
02
b110 6
#623970000000
1!
1%
1-
12
#623980000000
0!
0%
b111 *
0-
02
b111 6
#623990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#624000000000
0!
0%
b0 *
0-
02
b0 6
#624010000000
1!
1%
1-
12
#624020000000
0!
0%
b1 *
0-
02
b1 6
#624030000000
1!
1%
1-
12
#624040000000
0!
0%
b10 *
0-
02
b10 6
#624050000000
1!
1%
1-
12
#624060000000
0!
0%
b11 *
0-
02
b11 6
#624070000000
1!
1%
1-
12
15
#624080000000
0!
0%
b100 *
0-
02
b100 6
#624090000000
1!
1%
1-
12
#624100000000
0!
0%
b101 *
0-
02
b101 6
#624110000000
1!
1%
1-
12
#624120000000
0!
0%
b110 *
0-
02
b110 6
#624130000000
1!
1%
1-
12
#624140000000
0!
0%
b111 *
0-
02
b111 6
#624150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#624160000000
0!
0%
b0 *
0-
02
b0 6
#624170000000
1!
1%
1-
12
#624180000000
0!
0%
b1 *
0-
02
b1 6
#624190000000
1!
1%
1-
12
#624200000000
0!
0%
b10 *
0-
02
b10 6
#624210000000
1!
1%
1-
12
#624220000000
0!
0%
b11 *
0-
02
b11 6
#624230000000
1!
1%
1-
12
15
#624240000000
0!
0%
b100 *
0-
02
b100 6
#624250000000
1!
1%
1-
12
#624260000000
0!
0%
b101 *
0-
02
b101 6
#624270000000
1!
1%
1-
12
#624280000000
0!
0%
b110 *
0-
02
b110 6
#624290000000
1!
1%
1-
12
#624300000000
0!
0%
b111 *
0-
02
b111 6
#624310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#624320000000
0!
0%
b0 *
0-
02
b0 6
#624330000000
1!
1%
1-
12
#624340000000
0!
0%
b1 *
0-
02
b1 6
#624350000000
1!
1%
1-
12
#624360000000
0!
0%
b10 *
0-
02
b10 6
#624370000000
1!
1%
1-
12
#624380000000
0!
0%
b11 *
0-
02
b11 6
#624390000000
1!
1%
1-
12
15
#624400000000
0!
0%
b100 *
0-
02
b100 6
#624410000000
1!
1%
1-
12
#624420000000
0!
0%
b101 *
0-
02
b101 6
#624430000000
1!
1%
1-
12
#624440000000
0!
0%
b110 *
0-
02
b110 6
#624450000000
1!
1%
1-
12
#624460000000
0!
0%
b111 *
0-
02
b111 6
#624470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#624480000000
0!
0%
b0 *
0-
02
b0 6
#624490000000
1!
1%
1-
12
#624500000000
0!
0%
b1 *
0-
02
b1 6
#624510000000
1!
1%
1-
12
#624520000000
0!
0%
b10 *
0-
02
b10 6
#624530000000
1!
1%
1-
12
#624540000000
0!
0%
b11 *
0-
02
b11 6
#624550000000
1!
1%
1-
12
15
#624560000000
0!
0%
b100 *
0-
02
b100 6
#624570000000
1!
1%
1-
12
#624580000000
0!
0%
b101 *
0-
02
b101 6
#624590000000
1!
1%
1-
12
#624600000000
0!
0%
b110 *
0-
02
b110 6
#624610000000
1!
1%
1-
12
#624620000000
0!
0%
b111 *
0-
02
b111 6
#624630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#624640000000
0!
0%
b0 *
0-
02
b0 6
#624650000000
1!
1%
1-
12
#624660000000
0!
0%
b1 *
0-
02
b1 6
#624670000000
1!
1%
1-
12
#624680000000
0!
0%
b10 *
0-
02
b10 6
#624690000000
1!
1%
1-
12
#624700000000
0!
0%
b11 *
0-
02
b11 6
#624710000000
1!
1%
1-
12
15
#624720000000
0!
0%
b100 *
0-
02
b100 6
#624730000000
1!
1%
1-
12
#624740000000
0!
0%
b101 *
0-
02
b101 6
#624750000000
1!
1%
1-
12
#624760000000
0!
0%
b110 *
0-
02
b110 6
#624770000000
1!
1%
1-
12
#624780000000
0!
0%
b111 *
0-
02
b111 6
#624790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#624800000000
0!
0%
b0 *
0-
02
b0 6
#624810000000
1!
1%
1-
12
#624820000000
0!
0%
b1 *
0-
02
b1 6
#624830000000
1!
1%
1-
12
#624840000000
0!
0%
b10 *
0-
02
b10 6
#624850000000
1!
1%
1-
12
#624860000000
0!
0%
b11 *
0-
02
b11 6
#624870000000
1!
1%
1-
12
15
#624880000000
0!
0%
b100 *
0-
02
b100 6
#624890000000
1!
1%
1-
12
#624900000000
0!
0%
b101 *
0-
02
b101 6
#624910000000
1!
1%
1-
12
#624920000000
0!
0%
b110 *
0-
02
b110 6
#624930000000
1!
1%
1-
12
#624940000000
0!
0%
b111 *
0-
02
b111 6
#624950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#624960000000
0!
0%
b0 *
0-
02
b0 6
#624970000000
1!
1%
1-
12
#624980000000
0!
0%
b1 *
0-
02
b1 6
#624990000000
1!
1%
1-
12
#625000000000
0!
0%
b10 *
0-
02
b10 6
#625010000000
1!
1%
1-
12
#625020000000
0!
0%
b11 *
0-
02
b11 6
#625030000000
1!
1%
1-
12
15
#625040000000
0!
0%
b100 *
0-
02
b100 6
#625050000000
1!
1%
1-
12
#625060000000
0!
0%
b101 *
0-
02
b101 6
#625070000000
1!
1%
1-
12
#625080000000
0!
0%
b110 *
0-
02
b110 6
#625090000000
1!
1%
1-
12
#625100000000
0!
0%
b111 *
0-
02
b111 6
#625110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#625120000000
0!
0%
b0 *
0-
02
b0 6
#625130000000
1!
1%
1-
12
#625140000000
0!
0%
b1 *
0-
02
b1 6
#625150000000
1!
1%
1-
12
#625160000000
0!
0%
b10 *
0-
02
b10 6
#625170000000
1!
1%
1-
12
#625180000000
0!
0%
b11 *
0-
02
b11 6
#625190000000
1!
1%
1-
12
15
#625200000000
0!
0%
b100 *
0-
02
b100 6
#625210000000
1!
1%
1-
12
#625220000000
0!
0%
b101 *
0-
02
b101 6
#625230000000
1!
1%
1-
12
#625240000000
0!
0%
b110 *
0-
02
b110 6
#625250000000
1!
1%
1-
12
#625260000000
0!
0%
b111 *
0-
02
b111 6
#625270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#625280000000
0!
0%
b0 *
0-
02
b0 6
#625290000000
1!
1%
1-
12
#625300000000
0!
0%
b1 *
0-
02
b1 6
#625310000000
1!
1%
1-
12
#625320000000
0!
0%
b10 *
0-
02
b10 6
#625330000000
1!
1%
1-
12
#625340000000
0!
0%
b11 *
0-
02
b11 6
#625350000000
1!
1%
1-
12
15
#625360000000
0!
0%
b100 *
0-
02
b100 6
#625370000000
1!
1%
1-
12
#625380000000
0!
0%
b101 *
0-
02
b101 6
#625390000000
1!
1%
1-
12
#625400000000
0!
0%
b110 *
0-
02
b110 6
#625410000000
1!
1%
1-
12
#625420000000
0!
0%
b111 *
0-
02
b111 6
#625430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#625440000000
0!
0%
b0 *
0-
02
b0 6
#625450000000
1!
1%
1-
12
#625460000000
0!
0%
b1 *
0-
02
b1 6
#625470000000
1!
1%
1-
12
#625480000000
0!
0%
b10 *
0-
02
b10 6
#625490000000
1!
1%
1-
12
#625500000000
0!
0%
b11 *
0-
02
b11 6
#625510000000
1!
1%
1-
12
15
#625520000000
0!
0%
b100 *
0-
02
b100 6
#625530000000
1!
1%
1-
12
#625540000000
0!
0%
b101 *
0-
02
b101 6
#625550000000
1!
1%
1-
12
#625560000000
0!
0%
b110 *
0-
02
b110 6
#625570000000
1!
1%
1-
12
#625580000000
0!
0%
b111 *
0-
02
b111 6
#625590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#625600000000
0!
0%
b0 *
0-
02
b0 6
#625610000000
1!
1%
1-
12
#625620000000
0!
0%
b1 *
0-
02
b1 6
#625630000000
1!
1%
1-
12
#625640000000
0!
0%
b10 *
0-
02
b10 6
#625650000000
1!
1%
1-
12
#625660000000
0!
0%
b11 *
0-
02
b11 6
#625670000000
1!
1%
1-
12
15
#625680000000
0!
0%
b100 *
0-
02
b100 6
#625690000000
1!
1%
1-
12
#625700000000
0!
0%
b101 *
0-
02
b101 6
#625710000000
1!
1%
1-
12
#625720000000
0!
0%
b110 *
0-
02
b110 6
#625730000000
1!
1%
1-
12
#625740000000
0!
0%
b111 *
0-
02
b111 6
#625750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#625760000000
0!
0%
b0 *
0-
02
b0 6
#625770000000
1!
1%
1-
12
#625780000000
0!
0%
b1 *
0-
02
b1 6
#625790000000
1!
1%
1-
12
#625800000000
0!
0%
b10 *
0-
02
b10 6
#625810000000
1!
1%
1-
12
#625820000000
0!
0%
b11 *
0-
02
b11 6
#625830000000
1!
1%
1-
12
15
#625840000000
0!
0%
b100 *
0-
02
b100 6
#625850000000
1!
1%
1-
12
#625860000000
0!
0%
b101 *
0-
02
b101 6
#625870000000
1!
1%
1-
12
#625880000000
0!
0%
b110 *
0-
02
b110 6
#625890000000
1!
1%
1-
12
#625900000000
0!
0%
b111 *
0-
02
b111 6
#625910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#625920000000
0!
0%
b0 *
0-
02
b0 6
#625930000000
1!
1%
1-
12
#625940000000
0!
0%
b1 *
0-
02
b1 6
#625950000000
1!
1%
1-
12
#625960000000
0!
0%
b10 *
0-
02
b10 6
#625970000000
1!
1%
1-
12
#625980000000
0!
0%
b11 *
0-
02
b11 6
#625990000000
1!
1%
1-
12
15
#626000000000
0!
0%
b100 *
0-
02
b100 6
#626010000000
1!
1%
1-
12
#626020000000
0!
0%
b101 *
0-
02
b101 6
#626030000000
1!
1%
1-
12
#626040000000
0!
0%
b110 *
0-
02
b110 6
#626050000000
1!
1%
1-
12
#626060000000
0!
0%
b111 *
0-
02
b111 6
#626070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#626080000000
0!
0%
b0 *
0-
02
b0 6
#626090000000
1!
1%
1-
12
#626100000000
0!
0%
b1 *
0-
02
b1 6
#626110000000
1!
1%
1-
12
#626120000000
0!
0%
b10 *
0-
02
b10 6
#626130000000
1!
1%
1-
12
#626140000000
0!
0%
b11 *
0-
02
b11 6
#626150000000
1!
1%
1-
12
15
#626160000000
0!
0%
b100 *
0-
02
b100 6
#626170000000
1!
1%
1-
12
#626180000000
0!
0%
b101 *
0-
02
b101 6
#626190000000
1!
1%
1-
12
#626200000000
0!
0%
b110 *
0-
02
b110 6
#626210000000
1!
1%
1-
12
#626220000000
0!
0%
b111 *
0-
02
b111 6
#626230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#626240000000
0!
0%
b0 *
0-
02
b0 6
#626250000000
1!
1%
1-
12
#626260000000
0!
0%
b1 *
0-
02
b1 6
#626270000000
1!
1%
1-
12
#626280000000
0!
0%
b10 *
0-
02
b10 6
#626290000000
1!
1%
1-
12
#626300000000
0!
0%
b11 *
0-
02
b11 6
#626310000000
1!
1%
1-
12
15
#626320000000
0!
0%
b100 *
0-
02
b100 6
#626330000000
1!
1%
1-
12
#626340000000
0!
0%
b101 *
0-
02
b101 6
#626350000000
1!
1%
1-
12
#626360000000
0!
0%
b110 *
0-
02
b110 6
#626370000000
1!
1%
1-
12
#626380000000
0!
0%
b111 *
0-
02
b111 6
#626390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#626400000000
0!
0%
b0 *
0-
02
b0 6
#626410000000
1!
1%
1-
12
#626420000000
0!
0%
b1 *
0-
02
b1 6
#626430000000
1!
1%
1-
12
#626440000000
0!
0%
b10 *
0-
02
b10 6
#626450000000
1!
1%
1-
12
#626460000000
0!
0%
b11 *
0-
02
b11 6
#626470000000
1!
1%
1-
12
15
#626480000000
0!
0%
b100 *
0-
02
b100 6
#626490000000
1!
1%
1-
12
#626500000000
0!
0%
b101 *
0-
02
b101 6
#626510000000
1!
1%
1-
12
#626520000000
0!
0%
b110 *
0-
02
b110 6
#626530000000
1!
1%
1-
12
#626540000000
0!
0%
b111 *
0-
02
b111 6
#626550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#626560000000
0!
0%
b0 *
0-
02
b0 6
#626570000000
1!
1%
1-
12
#626580000000
0!
0%
b1 *
0-
02
b1 6
#626590000000
1!
1%
1-
12
#626600000000
0!
0%
b10 *
0-
02
b10 6
#626610000000
1!
1%
1-
12
#626620000000
0!
0%
b11 *
0-
02
b11 6
#626630000000
1!
1%
1-
12
15
#626640000000
0!
0%
b100 *
0-
02
b100 6
#626650000000
1!
1%
1-
12
#626660000000
0!
0%
b101 *
0-
02
b101 6
#626670000000
1!
1%
1-
12
#626680000000
0!
0%
b110 *
0-
02
b110 6
#626690000000
1!
1%
1-
12
#626700000000
0!
0%
b111 *
0-
02
b111 6
#626710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#626720000000
0!
0%
b0 *
0-
02
b0 6
#626730000000
1!
1%
1-
12
#626740000000
0!
0%
b1 *
0-
02
b1 6
#626750000000
1!
1%
1-
12
#626760000000
0!
0%
b10 *
0-
02
b10 6
#626770000000
1!
1%
1-
12
#626780000000
0!
0%
b11 *
0-
02
b11 6
#626790000000
1!
1%
1-
12
15
#626800000000
0!
0%
b100 *
0-
02
b100 6
#626810000000
1!
1%
1-
12
#626820000000
0!
0%
b101 *
0-
02
b101 6
#626830000000
1!
1%
1-
12
#626840000000
0!
0%
b110 *
0-
02
b110 6
#626850000000
1!
1%
1-
12
#626860000000
0!
0%
b111 *
0-
02
b111 6
#626870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#626880000000
0!
0%
b0 *
0-
02
b0 6
#626890000000
1!
1%
1-
12
#626900000000
0!
0%
b1 *
0-
02
b1 6
#626910000000
1!
1%
1-
12
#626920000000
0!
0%
b10 *
0-
02
b10 6
#626930000000
1!
1%
1-
12
#626940000000
0!
0%
b11 *
0-
02
b11 6
#626950000000
1!
1%
1-
12
15
#626960000000
0!
0%
b100 *
0-
02
b100 6
#626970000000
1!
1%
1-
12
#626980000000
0!
0%
b101 *
0-
02
b101 6
#626990000000
1!
1%
1-
12
#627000000000
0!
0%
b110 *
0-
02
b110 6
#627010000000
1!
1%
1-
12
#627020000000
0!
0%
b111 *
0-
02
b111 6
#627030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#627040000000
0!
0%
b0 *
0-
02
b0 6
#627050000000
1!
1%
1-
12
#627060000000
0!
0%
b1 *
0-
02
b1 6
#627070000000
1!
1%
1-
12
#627080000000
0!
0%
b10 *
0-
02
b10 6
#627090000000
1!
1%
1-
12
#627100000000
0!
0%
b11 *
0-
02
b11 6
#627110000000
1!
1%
1-
12
15
#627120000000
0!
0%
b100 *
0-
02
b100 6
#627130000000
1!
1%
1-
12
#627140000000
0!
0%
b101 *
0-
02
b101 6
#627150000000
1!
1%
1-
12
#627160000000
0!
0%
b110 *
0-
02
b110 6
#627170000000
1!
1%
1-
12
#627180000000
0!
0%
b111 *
0-
02
b111 6
#627190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#627200000000
0!
0%
b0 *
0-
02
b0 6
#627210000000
1!
1%
1-
12
#627220000000
0!
0%
b1 *
0-
02
b1 6
#627230000000
1!
1%
1-
12
#627240000000
0!
0%
b10 *
0-
02
b10 6
#627250000000
1!
1%
1-
12
#627260000000
0!
0%
b11 *
0-
02
b11 6
#627270000000
1!
1%
1-
12
15
#627280000000
0!
0%
b100 *
0-
02
b100 6
#627290000000
1!
1%
1-
12
#627300000000
0!
0%
b101 *
0-
02
b101 6
#627310000000
1!
1%
1-
12
#627320000000
0!
0%
b110 *
0-
02
b110 6
#627330000000
1!
1%
1-
12
#627340000000
0!
0%
b111 *
0-
02
b111 6
#627350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#627360000000
0!
0%
b0 *
0-
02
b0 6
#627370000000
1!
1%
1-
12
#627380000000
0!
0%
b1 *
0-
02
b1 6
#627390000000
1!
1%
1-
12
#627400000000
0!
0%
b10 *
0-
02
b10 6
#627410000000
1!
1%
1-
12
#627420000000
0!
0%
b11 *
0-
02
b11 6
#627430000000
1!
1%
1-
12
15
#627440000000
0!
0%
b100 *
0-
02
b100 6
#627450000000
1!
1%
1-
12
#627460000000
0!
0%
b101 *
0-
02
b101 6
#627470000000
1!
1%
1-
12
#627480000000
0!
0%
b110 *
0-
02
b110 6
#627490000000
1!
1%
1-
12
#627500000000
0!
0%
b111 *
0-
02
b111 6
#627510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#627520000000
0!
0%
b0 *
0-
02
b0 6
#627530000000
1!
1%
1-
12
#627540000000
0!
0%
b1 *
0-
02
b1 6
#627550000000
1!
1%
1-
12
#627560000000
0!
0%
b10 *
0-
02
b10 6
#627570000000
1!
1%
1-
12
#627580000000
0!
0%
b11 *
0-
02
b11 6
#627590000000
1!
1%
1-
12
15
#627600000000
0!
0%
b100 *
0-
02
b100 6
#627610000000
1!
1%
1-
12
#627620000000
0!
0%
b101 *
0-
02
b101 6
#627630000000
1!
1%
1-
12
#627640000000
0!
0%
b110 *
0-
02
b110 6
#627650000000
1!
1%
1-
12
#627660000000
0!
0%
b111 *
0-
02
b111 6
#627670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#627680000000
0!
0%
b0 *
0-
02
b0 6
#627690000000
1!
1%
1-
12
#627700000000
0!
0%
b1 *
0-
02
b1 6
#627710000000
1!
1%
1-
12
#627720000000
0!
0%
b10 *
0-
02
b10 6
#627730000000
1!
1%
1-
12
#627740000000
0!
0%
b11 *
0-
02
b11 6
#627750000000
1!
1%
1-
12
15
#627760000000
0!
0%
b100 *
0-
02
b100 6
#627770000000
1!
1%
1-
12
#627780000000
0!
0%
b101 *
0-
02
b101 6
#627790000000
1!
1%
1-
12
#627800000000
0!
0%
b110 *
0-
02
b110 6
#627810000000
1!
1%
1-
12
#627820000000
0!
0%
b111 *
0-
02
b111 6
#627830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#627840000000
0!
0%
b0 *
0-
02
b0 6
#627850000000
1!
1%
1-
12
#627860000000
0!
0%
b1 *
0-
02
b1 6
#627870000000
1!
1%
1-
12
#627880000000
0!
0%
b10 *
0-
02
b10 6
#627890000000
1!
1%
1-
12
#627900000000
0!
0%
b11 *
0-
02
b11 6
#627910000000
1!
1%
1-
12
15
#627920000000
0!
0%
b100 *
0-
02
b100 6
#627930000000
1!
1%
1-
12
#627940000000
0!
0%
b101 *
0-
02
b101 6
#627950000000
1!
1%
1-
12
#627960000000
0!
0%
b110 *
0-
02
b110 6
#627970000000
1!
1%
1-
12
#627980000000
0!
0%
b111 *
0-
02
b111 6
#627990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#628000000000
0!
0%
b0 *
0-
02
b0 6
#628010000000
1!
1%
1-
12
#628020000000
0!
0%
b1 *
0-
02
b1 6
#628030000000
1!
1%
1-
12
#628040000000
0!
0%
b10 *
0-
02
b10 6
#628050000000
1!
1%
1-
12
#628060000000
0!
0%
b11 *
0-
02
b11 6
#628070000000
1!
1%
1-
12
15
#628080000000
0!
0%
b100 *
0-
02
b100 6
#628090000000
1!
1%
1-
12
#628100000000
0!
0%
b101 *
0-
02
b101 6
#628110000000
1!
1%
1-
12
#628120000000
0!
0%
b110 *
0-
02
b110 6
#628130000000
1!
1%
1-
12
#628140000000
0!
0%
b111 *
0-
02
b111 6
#628150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#628160000000
0!
0%
b0 *
0-
02
b0 6
#628170000000
1!
1%
1-
12
#628180000000
0!
0%
b1 *
0-
02
b1 6
#628190000000
1!
1%
1-
12
#628200000000
0!
0%
b10 *
0-
02
b10 6
#628210000000
1!
1%
1-
12
#628220000000
0!
0%
b11 *
0-
02
b11 6
#628230000000
1!
1%
1-
12
15
#628240000000
0!
0%
b100 *
0-
02
b100 6
#628250000000
1!
1%
1-
12
#628260000000
0!
0%
b101 *
0-
02
b101 6
#628270000000
1!
1%
1-
12
#628280000000
0!
0%
b110 *
0-
02
b110 6
#628290000000
1!
1%
1-
12
#628300000000
0!
0%
b111 *
0-
02
b111 6
#628310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#628320000000
0!
0%
b0 *
0-
02
b0 6
#628330000000
1!
1%
1-
12
#628340000000
0!
0%
b1 *
0-
02
b1 6
#628350000000
1!
1%
1-
12
#628360000000
0!
0%
b10 *
0-
02
b10 6
#628370000000
1!
1%
1-
12
#628380000000
0!
0%
b11 *
0-
02
b11 6
#628390000000
1!
1%
1-
12
15
#628400000000
0!
0%
b100 *
0-
02
b100 6
#628410000000
1!
1%
1-
12
#628420000000
0!
0%
b101 *
0-
02
b101 6
#628430000000
1!
1%
1-
12
#628440000000
0!
0%
b110 *
0-
02
b110 6
#628450000000
1!
1%
1-
12
#628460000000
0!
0%
b111 *
0-
02
b111 6
#628470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#628480000000
0!
0%
b0 *
0-
02
b0 6
#628490000000
1!
1%
1-
12
#628500000000
0!
0%
b1 *
0-
02
b1 6
#628510000000
1!
1%
1-
12
#628520000000
0!
0%
b10 *
0-
02
b10 6
#628530000000
1!
1%
1-
12
#628540000000
0!
0%
b11 *
0-
02
b11 6
#628550000000
1!
1%
1-
12
15
#628560000000
0!
0%
b100 *
0-
02
b100 6
#628570000000
1!
1%
1-
12
#628580000000
0!
0%
b101 *
0-
02
b101 6
#628590000000
1!
1%
1-
12
#628600000000
0!
0%
b110 *
0-
02
b110 6
#628610000000
1!
1%
1-
12
#628620000000
0!
0%
b111 *
0-
02
b111 6
#628630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#628640000000
0!
0%
b0 *
0-
02
b0 6
#628650000000
1!
1%
1-
12
#628660000000
0!
0%
b1 *
0-
02
b1 6
#628670000000
1!
1%
1-
12
#628680000000
0!
0%
b10 *
0-
02
b10 6
#628690000000
1!
1%
1-
12
#628700000000
0!
0%
b11 *
0-
02
b11 6
#628710000000
1!
1%
1-
12
15
#628720000000
0!
0%
b100 *
0-
02
b100 6
#628730000000
1!
1%
1-
12
#628740000000
0!
0%
b101 *
0-
02
b101 6
#628750000000
1!
1%
1-
12
#628760000000
0!
0%
b110 *
0-
02
b110 6
#628770000000
1!
1%
1-
12
#628780000000
0!
0%
b111 *
0-
02
b111 6
#628790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#628800000000
0!
0%
b0 *
0-
02
b0 6
#628810000000
1!
1%
1-
12
#628820000000
0!
0%
b1 *
0-
02
b1 6
#628830000000
1!
1%
1-
12
#628840000000
0!
0%
b10 *
0-
02
b10 6
#628850000000
1!
1%
1-
12
#628860000000
0!
0%
b11 *
0-
02
b11 6
#628870000000
1!
1%
1-
12
15
#628880000000
0!
0%
b100 *
0-
02
b100 6
#628890000000
1!
1%
1-
12
#628900000000
0!
0%
b101 *
0-
02
b101 6
#628910000000
1!
1%
1-
12
#628920000000
0!
0%
b110 *
0-
02
b110 6
#628930000000
1!
1%
1-
12
#628940000000
0!
0%
b111 *
0-
02
b111 6
#628950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#628960000000
0!
0%
b0 *
0-
02
b0 6
#628970000000
1!
1%
1-
12
#628980000000
0!
0%
b1 *
0-
02
b1 6
#628990000000
1!
1%
1-
12
#629000000000
0!
0%
b10 *
0-
02
b10 6
#629010000000
1!
1%
1-
12
#629020000000
0!
0%
b11 *
0-
02
b11 6
#629030000000
1!
1%
1-
12
15
#629040000000
0!
0%
b100 *
0-
02
b100 6
#629050000000
1!
1%
1-
12
#629060000000
0!
0%
b101 *
0-
02
b101 6
#629070000000
1!
1%
1-
12
#629080000000
0!
0%
b110 *
0-
02
b110 6
#629090000000
1!
1%
1-
12
#629100000000
0!
0%
b111 *
0-
02
b111 6
#629110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#629120000000
0!
0%
b0 *
0-
02
b0 6
#629130000000
1!
1%
1-
12
#629140000000
0!
0%
b1 *
0-
02
b1 6
#629150000000
1!
1%
1-
12
#629160000000
0!
0%
b10 *
0-
02
b10 6
#629170000000
1!
1%
1-
12
#629180000000
0!
0%
b11 *
0-
02
b11 6
#629190000000
1!
1%
1-
12
15
#629200000000
0!
0%
b100 *
0-
02
b100 6
#629210000000
1!
1%
1-
12
#629220000000
0!
0%
b101 *
0-
02
b101 6
#629230000000
1!
1%
1-
12
#629240000000
0!
0%
b110 *
0-
02
b110 6
#629250000000
1!
1%
1-
12
#629260000000
0!
0%
b111 *
0-
02
b111 6
#629270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#629280000000
0!
0%
b0 *
0-
02
b0 6
#629290000000
1!
1%
1-
12
#629300000000
0!
0%
b1 *
0-
02
b1 6
#629310000000
1!
1%
1-
12
#629320000000
0!
0%
b10 *
0-
02
b10 6
#629330000000
1!
1%
1-
12
#629340000000
0!
0%
b11 *
0-
02
b11 6
#629350000000
1!
1%
1-
12
15
#629360000000
0!
0%
b100 *
0-
02
b100 6
#629370000000
1!
1%
1-
12
#629380000000
0!
0%
b101 *
0-
02
b101 6
#629390000000
1!
1%
1-
12
#629400000000
0!
0%
b110 *
0-
02
b110 6
#629410000000
1!
1%
1-
12
#629420000000
0!
0%
b111 *
0-
02
b111 6
#629430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#629440000000
0!
0%
b0 *
0-
02
b0 6
#629450000000
1!
1%
1-
12
#629460000000
0!
0%
b1 *
0-
02
b1 6
#629470000000
1!
1%
1-
12
#629480000000
0!
0%
b10 *
0-
02
b10 6
#629490000000
1!
1%
1-
12
#629500000000
0!
0%
b11 *
0-
02
b11 6
#629510000000
1!
1%
1-
12
15
#629520000000
0!
0%
b100 *
0-
02
b100 6
#629530000000
1!
1%
1-
12
#629540000000
0!
0%
b101 *
0-
02
b101 6
#629550000000
1!
1%
1-
12
#629560000000
0!
0%
b110 *
0-
02
b110 6
#629570000000
1!
1%
1-
12
#629580000000
0!
0%
b111 *
0-
02
b111 6
#629590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#629600000000
0!
0%
b0 *
0-
02
b0 6
#629610000000
1!
1%
1-
12
#629620000000
0!
0%
b1 *
0-
02
b1 6
#629630000000
1!
1%
1-
12
#629640000000
0!
0%
b10 *
0-
02
b10 6
#629650000000
1!
1%
1-
12
#629660000000
0!
0%
b11 *
0-
02
b11 6
#629670000000
1!
1%
1-
12
15
#629680000000
0!
0%
b100 *
0-
02
b100 6
#629690000000
1!
1%
1-
12
#629700000000
0!
0%
b101 *
0-
02
b101 6
#629710000000
1!
1%
1-
12
#629720000000
0!
0%
b110 *
0-
02
b110 6
#629730000000
1!
1%
1-
12
#629740000000
0!
0%
b111 *
0-
02
b111 6
#629750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#629760000000
0!
0%
b0 *
0-
02
b0 6
#629770000000
1!
1%
1-
12
#629780000000
0!
0%
b1 *
0-
02
b1 6
#629790000000
1!
1%
1-
12
#629800000000
0!
0%
b10 *
0-
02
b10 6
#629810000000
1!
1%
1-
12
#629820000000
0!
0%
b11 *
0-
02
b11 6
#629830000000
1!
1%
1-
12
15
#629840000000
0!
0%
b100 *
0-
02
b100 6
#629850000000
1!
1%
1-
12
#629860000000
0!
0%
b101 *
0-
02
b101 6
#629870000000
1!
1%
1-
12
#629880000000
0!
0%
b110 *
0-
02
b110 6
#629890000000
1!
1%
1-
12
#629900000000
0!
0%
b111 *
0-
02
b111 6
#629910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#629920000000
0!
0%
b0 *
0-
02
b0 6
#629930000000
1!
1%
1-
12
#629940000000
0!
0%
b1 *
0-
02
b1 6
#629950000000
1!
1%
1-
12
#629960000000
0!
0%
b10 *
0-
02
b10 6
#629970000000
1!
1%
1-
12
#629980000000
0!
0%
b11 *
0-
02
b11 6
#629990000000
1!
1%
1-
12
15
#630000000000
0!
0%
b100 *
0-
02
b100 6
#630010000000
1!
1%
1-
12
#630020000000
0!
0%
b101 *
0-
02
b101 6
#630030000000
1!
1%
1-
12
#630040000000
0!
0%
b110 *
0-
02
b110 6
#630050000000
1!
1%
1-
12
#630060000000
0!
0%
b111 *
0-
02
b111 6
#630070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#630080000000
0!
0%
b0 *
0-
02
b0 6
#630090000000
1!
1%
1-
12
#630100000000
0!
0%
b1 *
0-
02
b1 6
#630110000000
1!
1%
1-
12
#630120000000
0!
0%
b10 *
0-
02
b10 6
#630130000000
1!
1%
1-
12
#630140000000
0!
0%
b11 *
0-
02
b11 6
#630150000000
1!
1%
1-
12
15
#630160000000
0!
0%
b100 *
0-
02
b100 6
#630170000000
1!
1%
1-
12
#630180000000
0!
0%
b101 *
0-
02
b101 6
#630190000000
1!
1%
1-
12
#630200000000
0!
0%
b110 *
0-
02
b110 6
#630210000000
1!
1%
1-
12
#630220000000
0!
0%
b111 *
0-
02
b111 6
#630230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#630240000000
0!
0%
b0 *
0-
02
b0 6
#630250000000
1!
1%
1-
12
#630260000000
0!
0%
b1 *
0-
02
b1 6
#630270000000
1!
1%
1-
12
#630280000000
0!
0%
b10 *
0-
02
b10 6
#630290000000
1!
1%
1-
12
#630300000000
0!
0%
b11 *
0-
02
b11 6
#630310000000
1!
1%
1-
12
15
#630320000000
0!
0%
b100 *
0-
02
b100 6
#630330000000
1!
1%
1-
12
#630340000000
0!
0%
b101 *
0-
02
b101 6
#630350000000
1!
1%
1-
12
#630360000000
0!
0%
b110 *
0-
02
b110 6
#630370000000
1!
1%
1-
12
#630380000000
0!
0%
b111 *
0-
02
b111 6
#630390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#630400000000
0!
0%
b0 *
0-
02
b0 6
#630410000000
1!
1%
1-
12
#630420000000
0!
0%
b1 *
0-
02
b1 6
#630430000000
1!
1%
1-
12
#630440000000
0!
0%
b10 *
0-
02
b10 6
#630450000000
1!
1%
1-
12
#630460000000
0!
0%
b11 *
0-
02
b11 6
#630470000000
1!
1%
1-
12
15
#630480000000
0!
0%
b100 *
0-
02
b100 6
#630490000000
1!
1%
1-
12
#630500000000
0!
0%
b101 *
0-
02
b101 6
#630510000000
1!
1%
1-
12
#630520000000
0!
0%
b110 *
0-
02
b110 6
#630530000000
1!
1%
1-
12
#630540000000
0!
0%
b111 *
0-
02
b111 6
#630550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#630560000000
0!
0%
b0 *
0-
02
b0 6
#630570000000
1!
1%
1-
12
#630580000000
0!
0%
b1 *
0-
02
b1 6
#630590000000
1!
1%
1-
12
#630600000000
0!
0%
b10 *
0-
02
b10 6
#630610000000
1!
1%
1-
12
#630620000000
0!
0%
b11 *
0-
02
b11 6
#630630000000
1!
1%
1-
12
15
#630640000000
0!
0%
b100 *
0-
02
b100 6
#630650000000
1!
1%
1-
12
#630660000000
0!
0%
b101 *
0-
02
b101 6
#630670000000
1!
1%
1-
12
#630680000000
0!
0%
b110 *
0-
02
b110 6
#630690000000
1!
1%
1-
12
#630700000000
0!
0%
b111 *
0-
02
b111 6
#630710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#630720000000
0!
0%
b0 *
0-
02
b0 6
#630730000000
1!
1%
1-
12
#630740000000
0!
0%
b1 *
0-
02
b1 6
#630750000000
1!
1%
1-
12
#630760000000
0!
0%
b10 *
0-
02
b10 6
#630770000000
1!
1%
1-
12
#630780000000
0!
0%
b11 *
0-
02
b11 6
#630790000000
1!
1%
1-
12
15
#630800000000
0!
0%
b100 *
0-
02
b100 6
#630810000000
1!
1%
1-
12
#630820000000
0!
0%
b101 *
0-
02
b101 6
#630830000000
1!
1%
1-
12
#630840000000
0!
0%
b110 *
0-
02
b110 6
#630850000000
1!
1%
1-
12
#630860000000
0!
0%
b111 *
0-
02
b111 6
#630870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#630880000000
0!
0%
b0 *
0-
02
b0 6
#630890000000
1!
1%
1-
12
#630900000000
0!
0%
b1 *
0-
02
b1 6
#630910000000
1!
1%
1-
12
#630920000000
0!
0%
b10 *
0-
02
b10 6
#630930000000
1!
1%
1-
12
#630940000000
0!
0%
b11 *
0-
02
b11 6
#630950000000
1!
1%
1-
12
15
#630960000000
0!
0%
b100 *
0-
02
b100 6
#630970000000
1!
1%
1-
12
#630980000000
0!
0%
b101 *
0-
02
b101 6
#630990000000
1!
1%
1-
12
#631000000000
0!
0%
b110 *
0-
02
b110 6
#631010000000
1!
1%
1-
12
#631020000000
0!
0%
b111 *
0-
02
b111 6
#631030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#631040000000
0!
0%
b0 *
0-
02
b0 6
#631050000000
1!
1%
1-
12
#631060000000
0!
0%
b1 *
0-
02
b1 6
#631070000000
1!
1%
1-
12
#631080000000
0!
0%
b10 *
0-
02
b10 6
#631090000000
1!
1%
1-
12
#631100000000
0!
0%
b11 *
0-
02
b11 6
#631110000000
1!
1%
1-
12
15
#631120000000
0!
0%
b100 *
0-
02
b100 6
#631130000000
1!
1%
1-
12
#631140000000
0!
0%
b101 *
0-
02
b101 6
#631150000000
1!
1%
1-
12
#631160000000
0!
0%
b110 *
0-
02
b110 6
#631170000000
1!
1%
1-
12
#631180000000
0!
0%
b111 *
0-
02
b111 6
#631190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#631200000000
0!
0%
b0 *
0-
02
b0 6
#631210000000
1!
1%
1-
12
#631220000000
0!
0%
b1 *
0-
02
b1 6
#631230000000
1!
1%
1-
12
#631240000000
0!
0%
b10 *
0-
02
b10 6
#631250000000
1!
1%
1-
12
#631260000000
0!
0%
b11 *
0-
02
b11 6
#631270000000
1!
1%
1-
12
15
#631280000000
0!
0%
b100 *
0-
02
b100 6
#631290000000
1!
1%
1-
12
#631300000000
0!
0%
b101 *
0-
02
b101 6
#631310000000
1!
1%
1-
12
#631320000000
0!
0%
b110 *
0-
02
b110 6
#631330000000
1!
1%
1-
12
#631340000000
0!
0%
b111 *
0-
02
b111 6
#631350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#631360000000
0!
0%
b0 *
0-
02
b0 6
#631370000000
1!
1%
1-
12
#631380000000
0!
0%
b1 *
0-
02
b1 6
#631390000000
1!
1%
1-
12
#631400000000
0!
0%
b10 *
0-
02
b10 6
#631410000000
1!
1%
1-
12
#631420000000
0!
0%
b11 *
0-
02
b11 6
#631430000000
1!
1%
1-
12
15
#631440000000
0!
0%
b100 *
0-
02
b100 6
#631450000000
1!
1%
1-
12
#631460000000
0!
0%
b101 *
0-
02
b101 6
#631470000000
1!
1%
1-
12
#631480000000
0!
0%
b110 *
0-
02
b110 6
#631490000000
1!
1%
1-
12
#631500000000
0!
0%
b111 *
0-
02
b111 6
#631510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#631520000000
0!
0%
b0 *
0-
02
b0 6
#631530000000
1!
1%
1-
12
#631540000000
0!
0%
b1 *
0-
02
b1 6
#631550000000
1!
1%
1-
12
#631560000000
0!
0%
b10 *
0-
02
b10 6
#631570000000
1!
1%
1-
12
#631580000000
0!
0%
b11 *
0-
02
b11 6
#631590000000
1!
1%
1-
12
15
#631600000000
0!
0%
b100 *
0-
02
b100 6
#631610000000
1!
1%
1-
12
#631620000000
0!
0%
b101 *
0-
02
b101 6
#631630000000
1!
1%
1-
12
#631640000000
0!
0%
b110 *
0-
02
b110 6
#631650000000
1!
1%
1-
12
#631660000000
0!
0%
b111 *
0-
02
b111 6
#631670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#631680000000
0!
0%
b0 *
0-
02
b0 6
#631690000000
1!
1%
1-
12
#631700000000
0!
0%
b1 *
0-
02
b1 6
#631710000000
1!
1%
1-
12
#631720000000
0!
0%
b10 *
0-
02
b10 6
#631730000000
1!
1%
1-
12
#631740000000
0!
0%
b11 *
0-
02
b11 6
#631750000000
1!
1%
1-
12
15
#631760000000
0!
0%
b100 *
0-
02
b100 6
#631770000000
1!
1%
1-
12
#631780000000
0!
0%
b101 *
0-
02
b101 6
#631790000000
1!
1%
1-
12
#631800000000
0!
0%
b110 *
0-
02
b110 6
#631810000000
1!
1%
1-
12
#631820000000
0!
0%
b111 *
0-
02
b111 6
#631830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#631840000000
0!
0%
b0 *
0-
02
b0 6
#631850000000
1!
1%
1-
12
#631860000000
0!
0%
b1 *
0-
02
b1 6
#631870000000
1!
1%
1-
12
#631880000000
0!
0%
b10 *
0-
02
b10 6
#631890000000
1!
1%
1-
12
#631900000000
0!
0%
b11 *
0-
02
b11 6
#631910000000
1!
1%
1-
12
15
#631920000000
0!
0%
b100 *
0-
02
b100 6
#631930000000
1!
1%
1-
12
#631940000000
0!
0%
b101 *
0-
02
b101 6
#631950000000
1!
1%
1-
12
#631960000000
0!
0%
b110 *
0-
02
b110 6
#631970000000
1!
1%
1-
12
#631980000000
0!
0%
b111 *
0-
02
b111 6
#631990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#632000000000
0!
0%
b0 *
0-
02
b0 6
#632010000000
1!
1%
1-
12
#632020000000
0!
0%
b1 *
0-
02
b1 6
#632030000000
1!
1%
1-
12
#632040000000
0!
0%
b10 *
0-
02
b10 6
#632050000000
1!
1%
1-
12
#632060000000
0!
0%
b11 *
0-
02
b11 6
#632070000000
1!
1%
1-
12
15
#632080000000
0!
0%
b100 *
0-
02
b100 6
#632090000000
1!
1%
1-
12
#632100000000
0!
0%
b101 *
0-
02
b101 6
#632110000000
1!
1%
1-
12
#632120000000
0!
0%
b110 *
0-
02
b110 6
#632130000000
1!
1%
1-
12
#632140000000
0!
0%
b111 *
0-
02
b111 6
#632150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#632160000000
0!
0%
b0 *
0-
02
b0 6
#632170000000
1!
1%
1-
12
#632180000000
0!
0%
b1 *
0-
02
b1 6
#632190000000
1!
1%
1-
12
#632200000000
0!
0%
b10 *
0-
02
b10 6
#632210000000
1!
1%
1-
12
#632220000000
0!
0%
b11 *
0-
02
b11 6
#632230000000
1!
1%
1-
12
15
#632240000000
0!
0%
b100 *
0-
02
b100 6
#632250000000
1!
1%
1-
12
#632260000000
0!
0%
b101 *
0-
02
b101 6
#632270000000
1!
1%
1-
12
#632280000000
0!
0%
b110 *
0-
02
b110 6
#632290000000
1!
1%
1-
12
#632300000000
0!
0%
b111 *
0-
02
b111 6
#632310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#632320000000
0!
0%
b0 *
0-
02
b0 6
#632330000000
1!
1%
1-
12
#632340000000
0!
0%
b1 *
0-
02
b1 6
#632350000000
1!
1%
1-
12
#632360000000
0!
0%
b10 *
0-
02
b10 6
#632370000000
1!
1%
1-
12
#632380000000
0!
0%
b11 *
0-
02
b11 6
#632390000000
1!
1%
1-
12
15
#632400000000
0!
0%
b100 *
0-
02
b100 6
#632410000000
1!
1%
1-
12
#632420000000
0!
0%
b101 *
0-
02
b101 6
#632430000000
1!
1%
1-
12
#632440000000
0!
0%
b110 *
0-
02
b110 6
#632450000000
1!
1%
1-
12
#632460000000
0!
0%
b111 *
0-
02
b111 6
#632470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#632480000000
0!
0%
b0 *
0-
02
b0 6
#632490000000
1!
1%
1-
12
#632500000000
0!
0%
b1 *
0-
02
b1 6
#632510000000
1!
1%
1-
12
#632520000000
0!
0%
b10 *
0-
02
b10 6
#632530000000
1!
1%
1-
12
#632540000000
0!
0%
b11 *
0-
02
b11 6
#632550000000
1!
1%
1-
12
15
#632560000000
0!
0%
b100 *
0-
02
b100 6
#632570000000
1!
1%
1-
12
#632580000000
0!
0%
b101 *
0-
02
b101 6
#632590000000
1!
1%
1-
12
#632600000000
0!
0%
b110 *
0-
02
b110 6
#632610000000
1!
1%
1-
12
#632620000000
0!
0%
b111 *
0-
02
b111 6
#632630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#632640000000
0!
0%
b0 *
0-
02
b0 6
#632650000000
1!
1%
1-
12
#632660000000
0!
0%
b1 *
0-
02
b1 6
#632670000000
1!
1%
1-
12
#632680000000
0!
0%
b10 *
0-
02
b10 6
#632690000000
1!
1%
1-
12
#632700000000
0!
0%
b11 *
0-
02
b11 6
#632710000000
1!
1%
1-
12
15
#632720000000
0!
0%
b100 *
0-
02
b100 6
#632730000000
1!
1%
1-
12
#632740000000
0!
0%
b101 *
0-
02
b101 6
#632750000000
1!
1%
1-
12
#632760000000
0!
0%
b110 *
0-
02
b110 6
#632770000000
1!
1%
1-
12
#632780000000
0!
0%
b111 *
0-
02
b111 6
#632790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#632800000000
0!
0%
b0 *
0-
02
b0 6
#632810000000
1!
1%
1-
12
#632820000000
0!
0%
b1 *
0-
02
b1 6
#632830000000
1!
1%
1-
12
#632840000000
0!
0%
b10 *
0-
02
b10 6
#632850000000
1!
1%
1-
12
#632860000000
0!
0%
b11 *
0-
02
b11 6
#632870000000
1!
1%
1-
12
15
#632880000000
0!
0%
b100 *
0-
02
b100 6
#632890000000
1!
1%
1-
12
#632900000000
0!
0%
b101 *
0-
02
b101 6
#632910000000
1!
1%
1-
12
#632920000000
0!
0%
b110 *
0-
02
b110 6
#632930000000
1!
1%
1-
12
#632940000000
0!
0%
b111 *
0-
02
b111 6
#632950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#632960000000
0!
0%
b0 *
0-
02
b0 6
#632970000000
1!
1%
1-
12
#632980000000
0!
0%
b1 *
0-
02
b1 6
#632990000000
1!
1%
1-
12
#633000000000
0!
0%
b10 *
0-
02
b10 6
#633010000000
1!
1%
1-
12
#633020000000
0!
0%
b11 *
0-
02
b11 6
#633030000000
1!
1%
1-
12
15
#633040000000
0!
0%
b100 *
0-
02
b100 6
#633050000000
1!
1%
1-
12
#633060000000
0!
0%
b101 *
0-
02
b101 6
#633070000000
1!
1%
1-
12
#633080000000
0!
0%
b110 *
0-
02
b110 6
#633090000000
1!
1%
1-
12
#633100000000
0!
0%
b111 *
0-
02
b111 6
#633110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#633120000000
0!
0%
b0 *
0-
02
b0 6
#633130000000
1!
1%
1-
12
#633140000000
0!
0%
b1 *
0-
02
b1 6
#633150000000
1!
1%
1-
12
#633160000000
0!
0%
b10 *
0-
02
b10 6
#633170000000
1!
1%
1-
12
#633180000000
0!
0%
b11 *
0-
02
b11 6
#633190000000
1!
1%
1-
12
15
#633200000000
0!
0%
b100 *
0-
02
b100 6
#633210000000
1!
1%
1-
12
#633220000000
0!
0%
b101 *
0-
02
b101 6
#633230000000
1!
1%
1-
12
#633240000000
0!
0%
b110 *
0-
02
b110 6
#633250000000
1!
1%
1-
12
#633260000000
0!
0%
b111 *
0-
02
b111 6
#633270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#633280000000
0!
0%
b0 *
0-
02
b0 6
#633290000000
1!
1%
1-
12
#633300000000
0!
0%
b1 *
0-
02
b1 6
#633310000000
1!
1%
1-
12
#633320000000
0!
0%
b10 *
0-
02
b10 6
#633330000000
1!
1%
1-
12
#633340000000
0!
0%
b11 *
0-
02
b11 6
#633350000000
1!
1%
1-
12
15
#633360000000
0!
0%
b100 *
0-
02
b100 6
#633370000000
1!
1%
1-
12
#633380000000
0!
0%
b101 *
0-
02
b101 6
#633390000000
1!
1%
1-
12
#633400000000
0!
0%
b110 *
0-
02
b110 6
#633410000000
1!
1%
1-
12
#633420000000
0!
0%
b111 *
0-
02
b111 6
#633430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#633440000000
0!
0%
b0 *
0-
02
b0 6
#633450000000
1!
1%
1-
12
#633460000000
0!
0%
b1 *
0-
02
b1 6
#633470000000
1!
1%
1-
12
#633480000000
0!
0%
b10 *
0-
02
b10 6
#633490000000
1!
1%
1-
12
#633500000000
0!
0%
b11 *
0-
02
b11 6
#633510000000
1!
1%
1-
12
15
#633520000000
0!
0%
b100 *
0-
02
b100 6
#633530000000
1!
1%
1-
12
#633540000000
0!
0%
b101 *
0-
02
b101 6
#633550000000
1!
1%
1-
12
#633560000000
0!
0%
b110 *
0-
02
b110 6
#633570000000
1!
1%
1-
12
#633580000000
0!
0%
b111 *
0-
02
b111 6
#633590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#633600000000
0!
0%
b0 *
0-
02
b0 6
#633610000000
1!
1%
1-
12
#633620000000
0!
0%
b1 *
0-
02
b1 6
#633630000000
1!
1%
1-
12
#633640000000
0!
0%
b10 *
0-
02
b10 6
#633650000000
1!
1%
1-
12
#633660000000
0!
0%
b11 *
0-
02
b11 6
#633670000000
1!
1%
1-
12
15
#633680000000
0!
0%
b100 *
0-
02
b100 6
#633690000000
1!
1%
1-
12
#633700000000
0!
0%
b101 *
0-
02
b101 6
#633710000000
1!
1%
1-
12
#633720000000
0!
0%
b110 *
0-
02
b110 6
#633730000000
1!
1%
1-
12
#633740000000
0!
0%
b111 *
0-
02
b111 6
#633750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#633760000000
0!
0%
b0 *
0-
02
b0 6
#633770000000
1!
1%
1-
12
#633780000000
0!
0%
b1 *
0-
02
b1 6
#633790000000
1!
1%
1-
12
#633800000000
0!
0%
b10 *
0-
02
b10 6
#633810000000
1!
1%
1-
12
#633820000000
0!
0%
b11 *
0-
02
b11 6
#633830000000
1!
1%
1-
12
15
#633840000000
0!
0%
b100 *
0-
02
b100 6
#633850000000
1!
1%
1-
12
#633860000000
0!
0%
b101 *
0-
02
b101 6
#633870000000
1!
1%
1-
12
#633880000000
0!
0%
b110 *
0-
02
b110 6
#633890000000
1!
1%
1-
12
#633900000000
0!
0%
b111 *
0-
02
b111 6
#633910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#633920000000
0!
0%
b0 *
0-
02
b0 6
#633930000000
1!
1%
1-
12
#633940000000
0!
0%
b1 *
0-
02
b1 6
#633950000000
1!
1%
1-
12
#633960000000
0!
0%
b10 *
0-
02
b10 6
#633970000000
1!
1%
1-
12
#633980000000
0!
0%
b11 *
0-
02
b11 6
#633990000000
1!
1%
1-
12
15
#634000000000
0!
0%
b100 *
0-
02
b100 6
#634010000000
1!
1%
1-
12
#634020000000
0!
0%
b101 *
0-
02
b101 6
#634030000000
1!
1%
1-
12
#634040000000
0!
0%
b110 *
0-
02
b110 6
#634050000000
1!
1%
1-
12
#634060000000
0!
0%
b111 *
0-
02
b111 6
#634070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#634080000000
0!
0%
b0 *
0-
02
b0 6
#634090000000
1!
1%
1-
12
#634100000000
0!
0%
b1 *
0-
02
b1 6
#634110000000
1!
1%
1-
12
#634120000000
0!
0%
b10 *
0-
02
b10 6
#634130000000
1!
1%
1-
12
#634140000000
0!
0%
b11 *
0-
02
b11 6
#634150000000
1!
1%
1-
12
15
#634160000000
0!
0%
b100 *
0-
02
b100 6
#634170000000
1!
1%
1-
12
#634180000000
0!
0%
b101 *
0-
02
b101 6
#634190000000
1!
1%
1-
12
#634200000000
0!
0%
b110 *
0-
02
b110 6
#634210000000
1!
1%
1-
12
#634220000000
0!
0%
b111 *
0-
02
b111 6
#634230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#634240000000
0!
0%
b0 *
0-
02
b0 6
#634250000000
1!
1%
1-
12
#634260000000
0!
0%
b1 *
0-
02
b1 6
#634270000000
1!
1%
1-
12
#634280000000
0!
0%
b10 *
0-
02
b10 6
#634290000000
1!
1%
1-
12
#634300000000
0!
0%
b11 *
0-
02
b11 6
#634310000000
1!
1%
1-
12
15
#634320000000
0!
0%
b100 *
0-
02
b100 6
#634330000000
1!
1%
1-
12
#634340000000
0!
0%
b101 *
0-
02
b101 6
#634350000000
1!
1%
1-
12
#634360000000
0!
0%
b110 *
0-
02
b110 6
#634370000000
1!
1%
1-
12
#634380000000
0!
0%
b111 *
0-
02
b111 6
#634390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#634400000000
0!
0%
b0 *
0-
02
b0 6
#634410000000
1!
1%
1-
12
#634420000000
0!
0%
b1 *
0-
02
b1 6
#634430000000
1!
1%
1-
12
#634440000000
0!
0%
b10 *
0-
02
b10 6
#634450000000
1!
1%
1-
12
#634460000000
0!
0%
b11 *
0-
02
b11 6
#634470000000
1!
1%
1-
12
15
#634480000000
0!
0%
b100 *
0-
02
b100 6
#634490000000
1!
1%
1-
12
#634500000000
0!
0%
b101 *
0-
02
b101 6
#634510000000
1!
1%
1-
12
#634520000000
0!
0%
b110 *
0-
02
b110 6
#634530000000
1!
1%
1-
12
#634540000000
0!
0%
b111 *
0-
02
b111 6
#634550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#634560000000
0!
0%
b0 *
0-
02
b0 6
#634570000000
1!
1%
1-
12
#634580000000
0!
0%
b1 *
0-
02
b1 6
#634590000000
1!
1%
1-
12
#634600000000
0!
0%
b10 *
0-
02
b10 6
#634610000000
1!
1%
1-
12
#634620000000
0!
0%
b11 *
0-
02
b11 6
#634630000000
1!
1%
1-
12
15
#634640000000
0!
0%
b100 *
0-
02
b100 6
#634650000000
1!
1%
1-
12
#634660000000
0!
0%
b101 *
0-
02
b101 6
#634670000000
1!
1%
1-
12
#634680000000
0!
0%
b110 *
0-
02
b110 6
#634690000000
1!
1%
1-
12
#634700000000
0!
0%
b111 *
0-
02
b111 6
#634710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#634720000000
0!
0%
b0 *
0-
02
b0 6
#634730000000
1!
1%
1-
12
#634740000000
0!
0%
b1 *
0-
02
b1 6
#634750000000
1!
1%
1-
12
#634760000000
0!
0%
b10 *
0-
02
b10 6
#634770000000
1!
1%
1-
12
#634780000000
0!
0%
b11 *
0-
02
b11 6
#634790000000
1!
1%
1-
12
15
#634800000000
0!
0%
b100 *
0-
02
b100 6
#634810000000
1!
1%
1-
12
#634820000000
0!
0%
b101 *
0-
02
b101 6
#634830000000
1!
1%
1-
12
#634840000000
0!
0%
b110 *
0-
02
b110 6
#634850000000
1!
1%
1-
12
#634860000000
0!
0%
b111 *
0-
02
b111 6
#634870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#634880000000
0!
0%
b0 *
0-
02
b0 6
#634890000000
1!
1%
1-
12
#634900000000
0!
0%
b1 *
0-
02
b1 6
#634910000000
1!
1%
1-
12
#634920000000
0!
0%
b10 *
0-
02
b10 6
#634930000000
1!
1%
1-
12
#634940000000
0!
0%
b11 *
0-
02
b11 6
#634950000000
1!
1%
1-
12
15
#634960000000
0!
0%
b100 *
0-
02
b100 6
#634970000000
1!
1%
1-
12
#634980000000
0!
0%
b101 *
0-
02
b101 6
#634990000000
1!
1%
1-
12
#635000000000
0!
0%
b110 *
0-
02
b110 6
#635010000000
1!
1%
1-
12
#635020000000
0!
0%
b111 *
0-
02
b111 6
#635030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#635040000000
0!
0%
b0 *
0-
02
b0 6
#635050000000
1!
1%
1-
12
#635060000000
0!
0%
b1 *
0-
02
b1 6
#635070000000
1!
1%
1-
12
#635080000000
0!
0%
b10 *
0-
02
b10 6
#635090000000
1!
1%
1-
12
#635100000000
0!
0%
b11 *
0-
02
b11 6
#635110000000
1!
1%
1-
12
15
#635120000000
0!
0%
b100 *
0-
02
b100 6
#635130000000
1!
1%
1-
12
#635140000000
0!
0%
b101 *
0-
02
b101 6
#635150000000
1!
1%
1-
12
#635160000000
0!
0%
b110 *
0-
02
b110 6
#635170000000
1!
1%
1-
12
#635180000000
0!
0%
b111 *
0-
02
b111 6
#635190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#635200000000
0!
0%
b0 *
0-
02
b0 6
#635210000000
1!
1%
1-
12
#635220000000
0!
0%
b1 *
0-
02
b1 6
#635230000000
1!
1%
1-
12
#635240000000
0!
0%
b10 *
0-
02
b10 6
#635250000000
1!
1%
1-
12
#635260000000
0!
0%
b11 *
0-
02
b11 6
#635270000000
1!
1%
1-
12
15
#635280000000
0!
0%
b100 *
0-
02
b100 6
#635290000000
1!
1%
1-
12
#635300000000
0!
0%
b101 *
0-
02
b101 6
#635310000000
1!
1%
1-
12
#635320000000
0!
0%
b110 *
0-
02
b110 6
#635330000000
1!
1%
1-
12
#635340000000
0!
0%
b111 *
0-
02
b111 6
#635350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#635360000000
0!
0%
b0 *
0-
02
b0 6
#635370000000
1!
1%
1-
12
#635380000000
0!
0%
b1 *
0-
02
b1 6
#635390000000
1!
1%
1-
12
#635400000000
0!
0%
b10 *
0-
02
b10 6
#635410000000
1!
1%
1-
12
#635420000000
0!
0%
b11 *
0-
02
b11 6
#635430000000
1!
1%
1-
12
15
#635440000000
0!
0%
b100 *
0-
02
b100 6
#635450000000
1!
1%
1-
12
#635460000000
0!
0%
b101 *
0-
02
b101 6
#635470000000
1!
1%
1-
12
#635480000000
0!
0%
b110 *
0-
02
b110 6
#635490000000
1!
1%
1-
12
#635500000000
0!
0%
b111 *
0-
02
b111 6
#635510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#635520000000
0!
0%
b0 *
0-
02
b0 6
#635530000000
1!
1%
1-
12
#635540000000
0!
0%
b1 *
0-
02
b1 6
#635550000000
1!
1%
1-
12
#635560000000
0!
0%
b10 *
0-
02
b10 6
#635570000000
1!
1%
1-
12
#635580000000
0!
0%
b11 *
0-
02
b11 6
#635590000000
1!
1%
1-
12
15
#635600000000
0!
0%
b100 *
0-
02
b100 6
#635610000000
1!
1%
1-
12
#635620000000
0!
0%
b101 *
0-
02
b101 6
#635630000000
1!
1%
1-
12
#635640000000
0!
0%
b110 *
0-
02
b110 6
#635650000000
1!
1%
1-
12
#635660000000
0!
0%
b111 *
0-
02
b111 6
#635670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#635680000000
0!
0%
b0 *
0-
02
b0 6
#635690000000
1!
1%
1-
12
#635700000000
0!
0%
b1 *
0-
02
b1 6
#635710000000
1!
1%
1-
12
#635720000000
0!
0%
b10 *
0-
02
b10 6
#635730000000
1!
1%
1-
12
#635740000000
0!
0%
b11 *
0-
02
b11 6
#635750000000
1!
1%
1-
12
15
#635760000000
0!
0%
b100 *
0-
02
b100 6
#635770000000
1!
1%
1-
12
#635780000000
0!
0%
b101 *
0-
02
b101 6
#635790000000
1!
1%
1-
12
#635800000000
0!
0%
b110 *
0-
02
b110 6
#635810000000
1!
1%
1-
12
#635820000000
0!
0%
b111 *
0-
02
b111 6
#635830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#635840000000
0!
0%
b0 *
0-
02
b0 6
#635850000000
1!
1%
1-
12
#635860000000
0!
0%
b1 *
0-
02
b1 6
#635870000000
1!
1%
1-
12
#635880000000
0!
0%
b10 *
0-
02
b10 6
#635890000000
1!
1%
1-
12
#635900000000
0!
0%
b11 *
0-
02
b11 6
#635910000000
1!
1%
1-
12
15
#635920000000
0!
0%
b100 *
0-
02
b100 6
#635930000000
1!
1%
1-
12
#635940000000
0!
0%
b101 *
0-
02
b101 6
#635950000000
1!
1%
1-
12
#635960000000
0!
0%
b110 *
0-
02
b110 6
#635970000000
1!
1%
1-
12
#635980000000
0!
0%
b111 *
0-
02
b111 6
#635990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#636000000000
0!
0%
b0 *
0-
02
b0 6
#636010000000
1!
1%
1-
12
#636020000000
0!
0%
b1 *
0-
02
b1 6
#636030000000
1!
1%
1-
12
#636040000000
0!
0%
b10 *
0-
02
b10 6
#636050000000
1!
1%
1-
12
#636060000000
0!
0%
b11 *
0-
02
b11 6
#636070000000
1!
1%
1-
12
15
#636080000000
0!
0%
b100 *
0-
02
b100 6
#636090000000
1!
1%
1-
12
#636100000000
0!
0%
b101 *
0-
02
b101 6
#636110000000
1!
1%
1-
12
#636120000000
0!
0%
b110 *
0-
02
b110 6
#636130000000
1!
1%
1-
12
#636140000000
0!
0%
b111 *
0-
02
b111 6
#636150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#636160000000
0!
0%
b0 *
0-
02
b0 6
#636170000000
1!
1%
1-
12
#636180000000
0!
0%
b1 *
0-
02
b1 6
#636190000000
1!
1%
1-
12
#636200000000
0!
0%
b10 *
0-
02
b10 6
#636210000000
1!
1%
1-
12
#636220000000
0!
0%
b11 *
0-
02
b11 6
#636230000000
1!
1%
1-
12
15
#636240000000
0!
0%
b100 *
0-
02
b100 6
#636250000000
1!
1%
1-
12
#636260000000
0!
0%
b101 *
0-
02
b101 6
#636270000000
1!
1%
1-
12
#636280000000
0!
0%
b110 *
0-
02
b110 6
#636290000000
1!
1%
1-
12
#636300000000
0!
0%
b111 *
0-
02
b111 6
#636310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#636320000000
0!
0%
b0 *
0-
02
b0 6
#636330000000
1!
1%
1-
12
#636340000000
0!
0%
b1 *
0-
02
b1 6
#636350000000
1!
1%
1-
12
#636360000000
0!
0%
b10 *
0-
02
b10 6
#636370000000
1!
1%
1-
12
#636380000000
0!
0%
b11 *
0-
02
b11 6
#636390000000
1!
1%
1-
12
15
#636400000000
0!
0%
b100 *
0-
02
b100 6
#636410000000
1!
1%
1-
12
#636420000000
0!
0%
b101 *
0-
02
b101 6
#636430000000
1!
1%
1-
12
#636440000000
0!
0%
b110 *
0-
02
b110 6
#636450000000
1!
1%
1-
12
#636460000000
0!
0%
b111 *
0-
02
b111 6
#636470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#636480000000
0!
0%
b0 *
0-
02
b0 6
#636490000000
1!
1%
1-
12
#636500000000
0!
0%
b1 *
0-
02
b1 6
#636510000000
1!
1%
1-
12
#636520000000
0!
0%
b10 *
0-
02
b10 6
#636530000000
1!
1%
1-
12
#636540000000
0!
0%
b11 *
0-
02
b11 6
#636550000000
1!
1%
1-
12
15
#636560000000
0!
0%
b100 *
0-
02
b100 6
#636570000000
1!
1%
1-
12
#636580000000
0!
0%
b101 *
0-
02
b101 6
#636590000000
1!
1%
1-
12
#636600000000
0!
0%
b110 *
0-
02
b110 6
#636610000000
1!
1%
1-
12
#636620000000
0!
0%
b111 *
0-
02
b111 6
#636630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#636640000000
0!
0%
b0 *
0-
02
b0 6
#636650000000
1!
1%
1-
12
#636660000000
0!
0%
b1 *
0-
02
b1 6
#636670000000
1!
1%
1-
12
#636680000000
0!
0%
b10 *
0-
02
b10 6
#636690000000
1!
1%
1-
12
#636700000000
0!
0%
b11 *
0-
02
b11 6
#636710000000
1!
1%
1-
12
15
#636720000000
0!
0%
b100 *
0-
02
b100 6
#636730000000
1!
1%
1-
12
#636740000000
0!
0%
b101 *
0-
02
b101 6
#636750000000
1!
1%
1-
12
#636760000000
0!
0%
b110 *
0-
02
b110 6
#636770000000
1!
1%
1-
12
#636780000000
0!
0%
b111 *
0-
02
b111 6
#636790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#636800000000
0!
0%
b0 *
0-
02
b0 6
#636810000000
1!
1%
1-
12
#636820000000
0!
0%
b1 *
0-
02
b1 6
#636830000000
1!
1%
1-
12
#636840000000
0!
0%
b10 *
0-
02
b10 6
#636850000000
1!
1%
1-
12
#636860000000
0!
0%
b11 *
0-
02
b11 6
#636870000000
1!
1%
1-
12
15
#636880000000
0!
0%
b100 *
0-
02
b100 6
#636890000000
1!
1%
1-
12
#636900000000
0!
0%
b101 *
0-
02
b101 6
#636910000000
1!
1%
1-
12
#636920000000
0!
0%
b110 *
0-
02
b110 6
#636930000000
1!
1%
1-
12
#636940000000
0!
0%
b111 *
0-
02
b111 6
#636950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#636960000000
0!
0%
b0 *
0-
02
b0 6
#636970000000
1!
1%
1-
12
#636980000000
0!
0%
b1 *
0-
02
b1 6
#636990000000
1!
1%
1-
12
#637000000000
0!
0%
b10 *
0-
02
b10 6
#637010000000
1!
1%
1-
12
#637020000000
0!
0%
b11 *
0-
02
b11 6
#637030000000
1!
1%
1-
12
15
#637040000000
0!
0%
b100 *
0-
02
b100 6
#637050000000
1!
1%
1-
12
#637060000000
0!
0%
b101 *
0-
02
b101 6
#637070000000
1!
1%
1-
12
#637080000000
0!
0%
b110 *
0-
02
b110 6
#637090000000
1!
1%
1-
12
#637100000000
0!
0%
b111 *
0-
02
b111 6
#637110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#637120000000
0!
0%
b0 *
0-
02
b0 6
#637130000000
1!
1%
1-
12
#637140000000
0!
0%
b1 *
0-
02
b1 6
#637150000000
1!
1%
1-
12
#637160000000
0!
0%
b10 *
0-
02
b10 6
#637170000000
1!
1%
1-
12
#637180000000
0!
0%
b11 *
0-
02
b11 6
#637190000000
1!
1%
1-
12
15
#637200000000
0!
0%
b100 *
0-
02
b100 6
#637210000000
1!
1%
1-
12
#637220000000
0!
0%
b101 *
0-
02
b101 6
#637230000000
1!
1%
1-
12
#637240000000
0!
0%
b110 *
0-
02
b110 6
#637250000000
1!
1%
1-
12
#637260000000
0!
0%
b111 *
0-
02
b111 6
#637270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#637280000000
0!
0%
b0 *
0-
02
b0 6
#637290000000
1!
1%
1-
12
#637300000000
0!
0%
b1 *
0-
02
b1 6
#637310000000
1!
1%
1-
12
#637320000000
0!
0%
b10 *
0-
02
b10 6
#637330000000
1!
1%
1-
12
#637340000000
0!
0%
b11 *
0-
02
b11 6
#637350000000
1!
1%
1-
12
15
#637360000000
0!
0%
b100 *
0-
02
b100 6
#637370000000
1!
1%
1-
12
#637380000000
0!
0%
b101 *
0-
02
b101 6
#637390000000
1!
1%
1-
12
#637400000000
0!
0%
b110 *
0-
02
b110 6
#637410000000
1!
1%
1-
12
#637420000000
0!
0%
b111 *
0-
02
b111 6
#637430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#637440000000
0!
0%
b0 *
0-
02
b0 6
#637450000000
1!
1%
1-
12
#637460000000
0!
0%
b1 *
0-
02
b1 6
#637470000000
1!
1%
1-
12
#637480000000
0!
0%
b10 *
0-
02
b10 6
#637490000000
1!
1%
1-
12
#637500000000
0!
0%
b11 *
0-
02
b11 6
#637510000000
1!
1%
1-
12
15
#637520000000
0!
0%
b100 *
0-
02
b100 6
#637530000000
1!
1%
1-
12
#637540000000
0!
0%
b101 *
0-
02
b101 6
#637550000000
1!
1%
1-
12
#637560000000
0!
0%
b110 *
0-
02
b110 6
#637570000000
1!
1%
1-
12
#637580000000
0!
0%
b111 *
0-
02
b111 6
#637590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#637600000000
0!
0%
b0 *
0-
02
b0 6
#637610000000
1!
1%
1-
12
#637620000000
0!
0%
b1 *
0-
02
b1 6
#637630000000
1!
1%
1-
12
#637640000000
0!
0%
b10 *
0-
02
b10 6
#637650000000
1!
1%
1-
12
#637660000000
0!
0%
b11 *
0-
02
b11 6
#637670000000
1!
1%
1-
12
15
#637680000000
0!
0%
b100 *
0-
02
b100 6
#637690000000
1!
1%
1-
12
#637700000000
0!
0%
b101 *
0-
02
b101 6
#637710000000
1!
1%
1-
12
#637720000000
0!
0%
b110 *
0-
02
b110 6
#637730000000
1!
1%
1-
12
#637740000000
0!
0%
b111 *
0-
02
b111 6
#637750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#637760000000
0!
0%
b0 *
0-
02
b0 6
#637770000000
1!
1%
1-
12
#637780000000
0!
0%
b1 *
0-
02
b1 6
#637790000000
1!
1%
1-
12
#637800000000
0!
0%
b10 *
0-
02
b10 6
#637810000000
1!
1%
1-
12
#637820000000
0!
0%
b11 *
0-
02
b11 6
#637830000000
1!
1%
1-
12
15
#637840000000
0!
0%
b100 *
0-
02
b100 6
#637850000000
1!
1%
1-
12
#637860000000
0!
0%
b101 *
0-
02
b101 6
#637870000000
1!
1%
1-
12
#637880000000
0!
0%
b110 *
0-
02
b110 6
#637890000000
1!
1%
1-
12
#637900000000
0!
0%
b111 *
0-
02
b111 6
#637910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#637920000000
0!
0%
b0 *
0-
02
b0 6
#637930000000
1!
1%
1-
12
#637940000000
0!
0%
b1 *
0-
02
b1 6
#637950000000
1!
1%
1-
12
#637960000000
0!
0%
b10 *
0-
02
b10 6
#637970000000
1!
1%
1-
12
#637980000000
0!
0%
b11 *
0-
02
b11 6
#637990000000
1!
1%
1-
12
15
#638000000000
0!
0%
b100 *
0-
02
b100 6
#638010000000
1!
1%
1-
12
#638020000000
0!
0%
b101 *
0-
02
b101 6
#638030000000
1!
1%
1-
12
#638040000000
0!
0%
b110 *
0-
02
b110 6
#638050000000
1!
1%
1-
12
#638060000000
0!
0%
b111 *
0-
02
b111 6
#638070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#638080000000
0!
0%
b0 *
0-
02
b0 6
#638090000000
1!
1%
1-
12
#638100000000
0!
0%
b1 *
0-
02
b1 6
#638110000000
1!
1%
1-
12
#638120000000
0!
0%
b10 *
0-
02
b10 6
#638130000000
1!
1%
1-
12
#638140000000
0!
0%
b11 *
0-
02
b11 6
#638150000000
1!
1%
1-
12
15
#638160000000
0!
0%
b100 *
0-
02
b100 6
#638170000000
1!
1%
1-
12
#638180000000
0!
0%
b101 *
0-
02
b101 6
#638190000000
1!
1%
1-
12
#638200000000
0!
0%
b110 *
0-
02
b110 6
#638210000000
1!
1%
1-
12
#638220000000
0!
0%
b111 *
0-
02
b111 6
#638230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#638240000000
0!
0%
b0 *
0-
02
b0 6
#638250000000
1!
1%
1-
12
#638260000000
0!
0%
b1 *
0-
02
b1 6
#638270000000
1!
1%
1-
12
#638280000000
0!
0%
b10 *
0-
02
b10 6
#638290000000
1!
1%
1-
12
#638300000000
0!
0%
b11 *
0-
02
b11 6
#638310000000
1!
1%
1-
12
15
#638320000000
0!
0%
b100 *
0-
02
b100 6
#638330000000
1!
1%
1-
12
#638340000000
0!
0%
b101 *
0-
02
b101 6
#638350000000
1!
1%
1-
12
#638360000000
0!
0%
b110 *
0-
02
b110 6
#638370000000
1!
1%
1-
12
#638380000000
0!
0%
b111 *
0-
02
b111 6
#638390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#638400000000
0!
0%
b0 *
0-
02
b0 6
#638410000000
1!
1%
1-
12
#638420000000
0!
0%
b1 *
0-
02
b1 6
#638430000000
1!
1%
1-
12
#638440000000
0!
0%
b10 *
0-
02
b10 6
#638450000000
1!
1%
1-
12
#638460000000
0!
0%
b11 *
0-
02
b11 6
#638470000000
1!
1%
1-
12
15
#638480000000
0!
0%
b100 *
0-
02
b100 6
#638490000000
1!
1%
1-
12
#638500000000
0!
0%
b101 *
0-
02
b101 6
#638510000000
1!
1%
1-
12
#638520000000
0!
0%
b110 *
0-
02
b110 6
#638530000000
1!
1%
1-
12
#638540000000
0!
0%
b111 *
0-
02
b111 6
#638550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#638560000000
0!
0%
b0 *
0-
02
b0 6
#638570000000
1!
1%
1-
12
#638580000000
0!
0%
b1 *
0-
02
b1 6
#638590000000
1!
1%
1-
12
#638600000000
0!
0%
b10 *
0-
02
b10 6
#638610000000
1!
1%
1-
12
#638620000000
0!
0%
b11 *
0-
02
b11 6
#638630000000
1!
1%
1-
12
15
#638640000000
0!
0%
b100 *
0-
02
b100 6
#638650000000
1!
1%
1-
12
#638660000000
0!
0%
b101 *
0-
02
b101 6
#638670000000
1!
1%
1-
12
#638680000000
0!
0%
b110 *
0-
02
b110 6
#638690000000
1!
1%
1-
12
#638700000000
0!
0%
b111 *
0-
02
b111 6
#638710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#638720000000
0!
0%
b0 *
0-
02
b0 6
#638730000000
1!
1%
1-
12
#638740000000
0!
0%
b1 *
0-
02
b1 6
#638750000000
1!
1%
1-
12
#638760000000
0!
0%
b10 *
0-
02
b10 6
#638770000000
1!
1%
1-
12
#638780000000
0!
0%
b11 *
0-
02
b11 6
#638790000000
1!
1%
1-
12
15
#638800000000
0!
0%
b100 *
0-
02
b100 6
#638810000000
1!
1%
1-
12
#638820000000
0!
0%
b101 *
0-
02
b101 6
#638830000000
1!
1%
1-
12
#638840000000
0!
0%
b110 *
0-
02
b110 6
#638850000000
1!
1%
1-
12
#638860000000
0!
0%
b111 *
0-
02
b111 6
#638870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#638880000000
0!
0%
b0 *
0-
02
b0 6
#638890000000
1!
1%
1-
12
#638900000000
0!
0%
b1 *
0-
02
b1 6
#638910000000
1!
1%
1-
12
#638920000000
0!
0%
b10 *
0-
02
b10 6
#638930000000
1!
1%
1-
12
#638940000000
0!
0%
b11 *
0-
02
b11 6
#638950000000
1!
1%
1-
12
15
#638960000000
0!
0%
b100 *
0-
02
b100 6
#638970000000
1!
1%
1-
12
#638980000000
0!
0%
b101 *
0-
02
b101 6
#638990000000
1!
1%
1-
12
#639000000000
0!
0%
b110 *
0-
02
b110 6
#639010000000
1!
1%
1-
12
#639020000000
0!
0%
b111 *
0-
02
b111 6
#639030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#639040000000
0!
0%
b0 *
0-
02
b0 6
#639050000000
1!
1%
1-
12
#639060000000
0!
0%
b1 *
0-
02
b1 6
#639070000000
1!
1%
1-
12
#639080000000
0!
0%
b10 *
0-
02
b10 6
#639090000000
1!
1%
1-
12
#639100000000
0!
0%
b11 *
0-
02
b11 6
#639110000000
1!
1%
1-
12
15
#639120000000
0!
0%
b100 *
0-
02
b100 6
#639130000000
1!
1%
1-
12
#639140000000
0!
0%
b101 *
0-
02
b101 6
#639150000000
1!
1%
1-
12
#639160000000
0!
0%
b110 *
0-
02
b110 6
#639170000000
1!
1%
1-
12
#639180000000
0!
0%
b111 *
0-
02
b111 6
#639190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#639200000000
0!
0%
b0 *
0-
02
b0 6
#639210000000
1!
1%
1-
12
#639220000000
0!
0%
b1 *
0-
02
b1 6
#639230000000
1!
1%
1-
12
#639240000000
0!
0%
b10 *
0-
02
b10 6
#639250000000
1!
1%
1-
12
#639260000000
0!
0%
b11 *
0-
02
b11 6
#639270000000
1!
1%
1-
12
15
#639280000000
0!
0%
b100 *
0-
02
b100 6
#639290000000
1!
1%
1-
12
#639300000000
0!
0%
b101 *
0-
02
b101 6
#639310000000
1!
1%
1-
12
#639320000000
0!
0%
b110 *
0-
02
b110 6
#639330000000
1!
1%
1-
12
#639340000000
0!
0%
b111 *
0-
02
b111 6
#639350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#639360000000
0!
0%
b0 *
0-
02
b0 6
#639370000000
1!
1%
1-
12
#639380000000
0!
0%
b1 *
0-
02
b1 6
#639390000000
1!
1%
1-
12
#639400000000
0!
0%
b10 *
0-
02
b10 6
#639410000000
1!
1%
1-
12
#639420000000
0!
0%
b11 *
0-
02
b11 6
#639430000000
1!
1%
1-
12
15
#639440000000
0!
0%
b100 *
0-
02
b100 6
#639450000000
1!
1%
1-
12
#639460000000
0!
0%
b101 *
0-
02
b101 6
#639470000000
1!
1%
1-
12
#639480000000
0!
0%
b110 *
0-
02
b110 6
#639490000000
1!
1%
1-
12
#639500000000
0!
0%
b111 *
0-
02
b111 6
#639510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#639520000000
0!
0%
b0 *
0-
02
b0 6
#639530000000
1!
1%
1-
12
#639540000000
0!
0%
b1 *
0-
02
b1 6
#639550000000
1!
1%
1-
12
#639560000000
0!
0%
b10 *
0-
02
b10 6
#639570000000
1!
1%
1-
12
#639580000000
0!
0%
b11 *
0-
02
b11 6
#639590000000
1!
1%
1-
12
15
#639600000000
0!
0%
b100 *
0-
02
b100 6
#639610000000
1!
1%
1-
12
#639620000000
0!
0%
b101 *
0-
02
b101 6
#639630000000
1!
1%
1-
12
#639640000000
0!
0%
b110 *
0-
02
b110 6
#639650000000
1!
1%
1-
12
#639660000000
0!
0%
b111 *
0-
02
b111 6
#639670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#639680000000
0!
0%
b0 *
0-
02
b0 6
#639690000000
1!
1%
1-
12
#639700000000
0!
0%
b1 *
0-
02
b1 6
#639710000000
1!
1%
1-
12
#639720000000
0!
0%
b10 *
0-
02
b10 6
#639730000000
1!
1%
1-
12
#639740000000
0!
0%
b11 *
0-
02
b11 6
#639750000000
1!
1%
1-
12
15
#639760000000
0!
0%
b100 *
0-
02
b100 6
#639770000000
1!
1%
1-
12
#639780000000
0!
0%
b101 *
0-
02
b101 6
#639790000000
1!
1%
1-
12
#639800000000
0!
0%
b110 *
0-
02
b110 6
#639810000000
1!
1%
1-
12
#639820000000
0!
0%
b111 *
0-
02
b111 6
#639830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#639840000000
0!
0%
b0 *
0-
02
b0 6
#639850000000
1!
1%
1-
12
#639860000000
0!
0%
b1 *
0-
02
b1 6
#639870000000
1!
1%
1-
12
#639880000000
0!
0%
b10 *
0-
02
b10 6
#639890000000
1!
1%
1-
12
#639900000000
0!
0%
b11 *
0-
02
b11 6
#639910000000
1!
1%
1-
12
15
#639920000000
0!
0%
b100 *
0-
02
b100 6
#639930000000
1!
1%
1-
12
#639940000000
0!
0%
b101 *
0-
02
b101 6
#639950000000
1!
1%
1-
12
#639960000000
0!
0%
b110 *
0-
02
b110 6
#639970000000
1!
1%
1-
12
#639980000000
0!
0%
b111 *
0-
02
b111 6
#639990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#640000000000
0!
0%
b0 *
0-
02
b0 6
#640010000000
1!
1%
1-
12
#640020000000
0!
0%
b1 *
0-
02
b1 6
#640030000000
1!
1%
1-
12
#640040000000
0!
0%
b10 *
0-
02
b10 6
#640050000000
1!
1%
1-
12
#640060000000
0!
0%
b11 *
0-
02
b11 6
#640070000000
1!
1%
1-
12
15
#640080000000
0!
0%
b100 *
0-
02
b100 6
#640090000000
1!
1%
1-
12
#640100000000
0!
0%
b101 *
0-
02
b101 6
#640110000000
1!
1%
1-
12
#640120000000
0!
0%
b110 *
0-
02
b110 6
#640130000000
1!
1%
1-
12
#640140000000
0!
0%
b111 *
0-
02
b111 6
#640150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#640160000000
0!
0%
b0 *
0-
02
b0 6
#640170000000
1!
1%
1-
12
#640180000000
0!
0%
b1 *
0-
02
b1 6
#640190000000
1!
1%
1-
12
#640200000000
0!
0%
b10 *
0-
02
b10 6
#640210000000
1!
1%
1-
12
#640220000000
0!
0%
b11 *
0-
02
b11 6
#640230000000
1!
1%
1-
12
15
#640240000000
0!
0%
b100 *
0-
02
b100 6
#640250000000
1!
1%
1-
12
#640260000000
0!
0%
b101 *
0-
02
b101 6
#640270000000
1!
1%
1-
12
#640280000000
0!
0%
b110 *
0-
02
b110 6
#640290000000
1!
1%
1-
12
#640300000000
0!
0%
b111 *
0-
02
b111 6
#640310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#640320000000
0!
0%
b0 *
0-
02
b0 6
#640330000000
1!
1%
1-
12
#640340000000
0!
0%
b1 *
0-
02
b1 6
#640350000000
1!
1%
1-
12
#640360000000
0!
0%
b10 *
0-
02
b10 6
#640370000000
1!
1%
1-
12
#640380000000
0!
0%
b11 *
0-
02
b11 6
#640390000000
1!
1%
1-
12
15
#640400000000
0!
0%
b100 *
0-
02
b100 6
#640410000000
1!
1%
1-
12
#640420000000
0!
0%
b101 *
0-
02
b101 6
#640430000000
1!
1%
1-
12
#640440000000
0!
0%
b110 *
0-
02
b110 6
#640450000000
1!
1%
1-
12
#640460000000
0!
0%
b111 *
0-
02
b111 6
#640470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#640480000000
0!
0%
b0 *
0-
02
b0 6
#640490000000
1!
1%
1-
12
#640500000000
0!
0%
b1 *
0-
02
b1 6
#640510000000
1!
1%
1-
12
#640520000000
0!
0%
b10 *
0-
02
b10 6
#640530000000
1!
1%
1-
12
#640540000000
0!
0%
b11 *
0-
02
b11 6
#640550000000
1!
1%
1-
12
15
#640560000000
0!
0%
b100 *
0-
02
b100 6
#640570000000
1!
1%
1-
12
#640580000000
0!
0%
b101 *
0-
02
b101 6
#640590000000
1!
1%
1-
12
#640600000000
0!
0%
b110 *
0-
02
b110 6
#640610000000
1!
1%
1-
12
#640620000000
0!
0%
b111 *
0-
02
b111 6
#640630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#640640000000
0!
0%
b0 *
0-
02
b0 6
#640650000000
1!
1%
1-
12
#640660000000
0!
0%
b1 *
0-
02
b1 6
#640670000000
1!
1%
1-
12
#640680000000
0!
0%
b10 *
0-
02
b10 6
#640690000000
1!
1%
1-
12
#640700000000
0!
0%
b11 *
0-
02
b11 6
#640710000000
1!
1%
1-
12
15
#640720000000
0!
0%
b100 *
0-
02
b100 6
#640730000000
1!
1%
1-
12
#640740000000
0!
0%
b101 *
0-
02
b101 6
#640750000000
1!
1%
1-
12
#640760000000
0!
0%
b110 *
0-
02
b110 6
#640770000000
1!
1%
1-
12
#640780000000
0!
0%
b111 *
0-
02
b111 6
#640790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#640800000000
0!
0%
b0 *
0-
02
b0 6
#640810000000
1!
1%
1-
12
#640820000000
0!
0%
b1 *
0-
02
b1 6
#640830000000
1!
1%
1-
12
#640840000000
0!
0%
b10 *
0-
02
b10 6
#640850000000
1!
1%
1-
12
#640860000000
0!
0%
b11 *
0-
02
b11 6
#640870000000
1!
1%
1-
12
15
#640880000000
0!
0%
b100 *
0-
02
b100 6
#640890000000
1!
1%
1-
12
#640900000000
0!
0%
b101 *
0-
02
b101 6
#640910000000
1!
1%
1-
12
#640920000000
0!
0%
b110 *
0-
02
b110 6
#640930000000
1!
1%
1-
12
#640940000000
0!
0%
b111 *
0-
02
b111 6
#640950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#640960000000
0!
0%
b0 *
0-
02
b0 6
#640970000000
1!
1%
1-
12
#640980000000
0!
0%
b1 *
0-
02
b1 6
#640990000000
1!
1%
1-
12
#641000000000
0!
0%
b10 *
0-
02
b10 6
#641010000000
1!
1%
1-
12
#641020000000
0!
0%
b11 *
0-
02
b11 6
#641030000000
1!
1%
1-
12
15
#641040000000
0!
0%
b100 *
0-
02
b100 6
#641050000000
1!
1%
1-
12
#641060000000
0!
0%
b101 *
0-
02
b101 6
#641070000000
1!
1%
1-
12
#641080000000
0!
0%
b110 *
0-
02
b110 6
#641090000000
1!
1%
1-
12
#641100000000
0!
0%
b111 *
0-
02
b111 6
#641110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#641120000000
0!
0%
b0 *
0-
02
b0 6
#641130000000
1!
1%
1-
12
#641140000000
0!
0%
b1 *
0-
02
b1 6
#641150000000
1!
1%
1-
12
#641160000000
0!
0%
b10 *
0-
02
b10 6
#641170000000
1!
1%
1-
12
#641180000000
0!
0%
b11 *
0-
02
b11 6
#641190000000
1!
1%
1-
12
15
#641200000000
0!
0%
b100 *
0-
02
b100 6
#641210000000
1!
1%
1-
12
#641220000000
0!
0%
b101 *
0-
02
b101 6
#641230000000
1!
1%
1-
12
#641240000000
0!
0%
b110 *
0-
02
b110 6
#641250000000
1!
1%
1-
12
#641260000000
0!
0%
b111 *
0-
02
b111 6
#641270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#641280000000
0!
0%
b0 *
0-
02
b0 6
#641290000000
1!
1%
1-
12
#641300000000
0!
0%
b1 *
0-
02
b1 6
#641310000000
1!
1%
1-
12
#641320000000
0!
0%
b10 *
0-
02
b10 6
#641330000000
1!
1%
1-
12
#641340000000
0!
0%
b11 *
0-
02
b11 6
#641350000000
1!
1%
1-
12
15
#641360000000
0!
0%
b100 *
0-
02
b100 6
#641370000000
1!
1%
1-
12
#641380000000
0!
0%
b101 *
0-
02
b101 6
#641390000000
1!
1%
1-
12
#641400000000
0!
0%
b110 *
0-
02
b110 6
#641410000000
1!
1%
1-
12
#641420000000
0!
0%
b111 *
0-
02
b111 6
#641430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#641440000000
0!
0%
b0 *
0-
02
b0 6
#641450000000
1!
1%
1-
12
#641460000000
0!
0%
b1 *
0-
02
b1 6
#641470000000
1!
1%
1-
12
#641480000000
0!
0%
b10 *
0-
02
b10 6
#641490000000
1!
1%
1-
12
#641500000000
0!
0%
b11 *
0-
02
b11 6
#641510000000
1!
1%
1-
12
15
#641520000000
0!
0%
b100 *
0-
02
b100 6
#641530000000
1!
1%
1-
12
#641540000000
0!
0%
b101 *
0-
02
b101 6
#641550000000
1!
1%
1-
12
#641560000000
0!
0%
b110 *
0-
02
b110 6
#641570000000
1!
1%
1-
12
#641580000000
0!
0%
b111 *
0-
02
b111 6
#641590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#641600000000
0!
0%
b0 *
0-
02
b0 6
#641610000000
1!
1%
1-
12
#641620000000
0!
0%
b1 *
0-
02
b1 6
#641630000000
1!
1%
1-
12
#641640000000
0!
0%
b10 *
0-
02
b10 6
#641650000000
1!
1%
1-
12
#641660000000
0!
0%
b11 *
0-
02
b11 6
#641670000000
1!
1%
1-
12
15
#641680000000
0!
0%
b100 *
0-
02
b100 6
#641690000000
1!
1%
1-
12
#641700000000
0!
0%
b101 *
0-
02
b101 6
#641710000000
1!
1%
1-
12
#641720000000
0!
0%
b110 *
0-
02
b110 6
#641730000000
1!
1%
1-
12
#641740000000
0!
0%
b111 *
0-
02
b111 6
#641750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#641760000000
0!
0%
b0 *
0-
02
b0 6
#641770000000
1!
1%
1-
12
#641780000000
0!
0%
b1 *
0-
02
b1 6
#641790000000
1!
1%
1-
12
#641800000000
0!
0%
b10 *
0-
02
b10 6
#641810000000
1!
1%
1-
12
#641820000000
0!
0%
b11 *
0-
02
b11 6
#641830000000
1!
1%
1-
12
15
#641840000000
0!
0%
b100 *
0-
02
b100 6
#641850000000
1!
1%
1-
12
#641860000000
0!
0%
b101 *
0-
02
b101 6
#641870000000
1!
1%
1-
12
#641880000000
0!
0%
b110 *
0-
02
b110 6
#641890000000
1!
1%
1-
12
#641900000000
0!
0%
b111 *
0-
02
b111 6
#641910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#641920000000
0!
0%
b0 *
0-
02
b0 6
#641930000000
1!
1%
1-
12
#641940000000
0!
0%
b1 *
0-
02
b1 6
#641950000000
1!
1%
1-
12
#641960000000
0!
0%
b10 *
0-
02
b10 6
#641970000000
1!
1%
1-
12
#641980000000
0!
0%
b11 *
0-
02
b11 6
#641990000000
1!
1%
1-
12
15
#642000000000
0!
0%
b100 *
0-
02
b100 6
#642010000000
1!
1%
1-
12
#642020000000
0!
0%
b101 *
0-
02
b101 6
#642030000000
1!
1%
1-
12
#642040000000
0!
0%
b110 *
0-
02
b110 6
#642050000000
1!
1%
1-
12
#642060000000
0!
0%
b111 *
0-
02
b111 6
#642070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#642080000000
0!
0%
b0 *
0-
02
b0 6
#642090000000
1!
1%
1-
12
#642100000000
0!
0%
b1 *
0-
02
b1 6
#642110000000
1!
1%
1-
12
#642120000000
0!
0%
b10 *
0-
02
b10 6
#642130000000
1!
1%
1-
12
#642140000000
0!
0%
b11 *
0-
02
b11 6
#642150000000
1!
1%
1-
12
15
#642160000000
0!
0%
b100 *
0-
02
b100 6
#642170000000
1!
1%
1-
12
#642180000000
0!
0%
b101 *
0-
02
b101 6
#642190000000
1!
1%
1-
12
#642200000000
0!
0%
b110 *
0-
02
b110 6
#642210000000
1!
1%
1-
12
#642220000000
0!
0%
b111 *
0-
02
b111 6
#642230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#642240000000
0!
0%
b0 *
0-
02
b0 6
#642250000000
1!
1%
1-
12
#642260000000
0!
0%
b1 *
0-
02
b1 6
#642270000000
1!
1%
1-
12
#642280000000
0!
0%
b10 *
0-
02
b10 6
#642290000000
1!
1%
1-
12
#642300000000
0!
0%
b11 *
0-
02
b11 6
#642310000000
1!
1%
1-
12
15
#642320000000
0!
0%
b100 *
0-
02
b100 6
#642330000000
1!
1%
1-
12
#642340000000
0!
0%
b101 *
0-
02
b101 6
#642350000000
1!
1%
1-
12
#642360000000
0!
0%
b110 *
0-
02
b110 6
#642370000000
1!
1%
1-
12
#642380000000
0!
0%
b111 *
0-
02
b111 6
#642390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#642400000000
0!
0%
b0 *
0-
02
b0 6
#642410000000
1!
1%
1-
12
#642420000000
0!
0%
b1 *
0-
02
b1 6
#642430000000
1!
1%
1-
12
#642440000000
0!
0%
b10 *
0-
02
b10 6
#642450000000
1!
1%
1-
12
#642460000000
0!
0%
b11 *
0-
02
b11 6
#642470000000
1!
1%
1-
12
15
#642480000000
0!
0%
b100 *
0-
02
b100 6
#642490000000
1!
1%
1-
12
#642500000000
0!
0%
b101 *
0-
02
b101 6
#642510000000
1!
1%
1-
12
#642520000000
0!
0%
b110 *
0-
02
b110 6
#642530000000
1!
1%
1-
12
#642540000000
0!
0%
b111 *
0-
02
b111 6
#642550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#642560000000
0!
0%
b0 *
0-
02
b0 6
#642570000000
1!
1%
1-
12
#642580000000
0!
0%
b1 *
0-
02
b1 6
#642590000000
1!
1%
1-
12
#642600000000
0!
0%
b10 *
0-
02
b10 6
#642610000000
1!
1%
1-
12
#642620000000
0!
0%
b11 *
0-
02
b11 6
#642630000000
1!
1%
1-
12
15
#642640000000
0!
0%
b100 *
0-
02
b100 6
#642650000000
1!
1%
1-
12
#642660000000
0!
0%
b101 *
0-
02
b101 6
#642670000000
1!
1%
1-
12
#642680000000
0!
0%
b110 *
0-
02
b110 6
#642690000000
1!
1%
1-
12
#642700000000
0!
0%
b111 *
0-
02
b111 6
#642710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#642720000000
0!
0%
b0 *
0-
02
b0 6
#642730000000
1!
1%
1-
12
#642740000000
0!
0%
b1 *
0-
02
b1 6
#642750000000
1!
1%
1-
12
#642760000000
0!
0%
b10 *
0-
02
b10 6
#642770000000
1!
1%
1-
12
#642780000000
0!
0%
b11 *
0-
02
b11 6
#642790000000
1!
1%
1-
12
15
#642800000000
0!
0%
b100 *
0-
02
b100 6
#642810000000
1!
1%
1-
12
#642820000000
0!
0%
b101 *
0-
02
b101 6
#642830000000
1!
1%
1-
12
#642840000000
0!
0%
b110 *
0-
02
b110 6
#642850000000
1!
1%
1-
12
#642860000000
0!
0%
b111 *
0-
02
b111 6
#642870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#642880000000
0!
0%
b0 *
0-
02
b0 6
#642890000000
1!
1%
1-
12
#642900000000
0!
0%
b1 *
0-
02
b1 6
#642910000000
1!
1%
1-
12
#642920000000
0!
0%
b10 *
0-
02
b10 6
#642930000000
1!
1%
1-
12
#642940000000
0!
0%
b11 *
0-
02
b11 6
#642950000000
1!
1%
1-
12
15
#642960000000
0!
0%
b100 *
0-
02
b100 6
#642970000000
1!
1%
1-
12
#642980000000
0!
0%
b101 *
0-
02
b101 6
#642990000000
1!
1%
1-
12
#643000000000
0!
0%
b110 *
0-
02
b110 6
#643010000000
1!
1%
1-
12
#643020000000
0!
0%
b111 *
0-
02
b111 6
#643030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#643040000000
0!
0%
b0 *
0-
02
b0 6
#643050000000
1!
1%
1-
12
#643060000000
0!
0%
b1 *
0-
02
b1 6
#643070000000
1!
1%
1-
12
#643080000000
0!
0%
b10 *
0-
02
b10 6
#643090000000
1!
1%
1-
12
#643100000000
0!
0%
b11 *
0-
02
b11 6
#643110000000
1!
1%
1-
12
15
#643120000000
0!
0%
b100 *
0-
02
b100 6
#643130000000
1!
1%
1-
12
#643140000000
0!
0%
b101 *
0-
02
b101 6
#643150000000
1!
1%
1-
12
#643160000000
0!
0%
b110 *
0-
02
b110 6
#643170000000
1!
1%
1-
12
#643180000000
0!
0%
b111 *
0-
02
b111 6
#643190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#643200000000
0!
0%
b0 *
0-
02
b0 6
#643210000000
1!
1%
1-
12
#643220000000
0!
0%
b1 *
0-
02
b1 6
#643230000000
1!
1%
1-
12
#643240000000
0!
0%
b10 *
0-
02
b10 6
#643250000000
1!
1%
1-
12
#643260000000
0!
0%
b11 *
0-
02
b11 6
#643270000000
1!
1%
1-
12
15
#643280000000
0!
0%
b100 *
0-
02
b100 6
#643290000000
1!
1%
1-
12
#643300000000
0!
0%
b101 *
0-
02
b101 6
#643310000000
1!
1%
1-
12
#643320000000
0!
0%
b110 *
0-
02
b110 6
#643330000000
1!
1%
1-
12
#643340000000
0!
0%
b111 *
0-
02
b111 6
#643350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#643360000000
0!
0%
b0 *
0-
02
b0 6
#643370000000
1!
1%
1-
12
#643380000000
0!
0%
b1 *
0-
02
b1 6
#643390000000
1!
1%
1-
12
#643400000000
0!
0%
b10 *
0-
02
b10 6
#643410000000
1!
1%
1-
12
#643420000000
0!
0%
b11 *
0-
02
b11 6
#643430000000
1!
1%
1-
12
15
#643440000000
0!
0%
b100 *
0-
02
b100 6
#643450000000
1!
1%
1-
12
#643460000000
0!
0%
b101 *
0-
02
b101 6
#643470000000
1!
1%
1-
12
#643480000000
0!
0%
b110 *
0-
02
b110 6
#643490000000
1!
1%
1-
12
#643500000000
0!
0%
b111 *
0-
02
b111 6
#643510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#643520000000
0!
0%
b0 *
0-
02
b0 6
#643530000000
1!
1%
1-
12
#643540000000
0!
0%
b1 *
0-
02
b1 6
#643550000000
1!
1%
1-
12
#643560000000
0!
0%
b10 *
0-
02
b10 6
#643570000000
1!
1%
1-
12
#643580000000
0!
0%
b11 *
0-
02
b11 6
#643590000000
1!
1%
1-
12
15
#643600000000
0!
0%
b100 *
0-
02
b100 6
#643610000000
1!
1%
1-
12
#643620000000
0!
0%
b101 *
0-
02
b101 6
#643630000000
1!
1%
1-
12
#643640000000
0!
0%
b110 *
0-
02
b110 6
#643650000000
1!
1%
1-
12
#643660000000
0!
0%
b111 *
0-
02
b111 6
#643670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#643680000000
0!
0%
b0 *
0-
02
b0 6
#643690000000
1!
1%
1-
12
#643700000000
0!
0%
b1 *
0-
02
b1 6
#643710000000
1!
1%
1-
12
#643720000000
0!
0%
b10 *
0-
02
b10 6
#643730000000
1!
1%
1-
12
#643740000000
0!
0%
b11 *
0-
02
b11 6
#643750000000
1!
1%
1-
12
15
#643760000000
0!
0%
b100 *
0-
02
b100 6
#643770000000
1!
1%
1-
12
#643780000000
0!
0%
b101 *
0-
02
b101 6
#643790000000
1!
1%
1-
12
#643800000000
0!
0%
b110 *
0-
02
b110 6
#643810000000
1!
1%
1-
12
#643820000000
0!
0%
b111 *
0-
02
b111 6
#643830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#643840000000
0!
0%
b0 *
0-
02
b0 6
#643850000000
1!
1%
1-
12
#643860000000
0!
0%
b1 *
0-
02
b1 6
#643870000000
1!
1%
1-
12
#643880000000
0!
0%
b10 *
0-
02
b10 6
#643890000000
1!
1%
1-
12
#643900000000
0!
0%
b11 *
0-
02
b11 6
#643910000000
1!
1%
1-
12
15
#643920000000
0!
0%
b100 *
0-
02
b100 6
#643930000000
1!
1%
1-
12
#643940000000
0!
0%
b101 *
0-
02
b101 6
#643950000000
1!
1%
1-
12
#643960000000
0!
0%
b110 *
0-
02
b110 6
#643970000000
1!
1%
1-
12
#643980000000
0!
0%
b111 *
0-
02
b111 6
#643990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#644000000000
0!
0%
b0 *
0-
02
b0 6
#644010000000
1!
1%
1-
12
#644020000000
0!
0%
b1 *
0-
02
b1 6
#644030000000
1!
1%
1-
12
#644040000000
0!
0%
b10 *
0-
02
b10 6
#644050000000
1!
1%
1-
12
#644060000000
0!
0%
b11 *
0-
02
b11 6
#644070000000
1!
1%
1-
12
15
#644080000000
0!
0%
b100 *
0-
02
b100 6
#644090000000
1!
1%
1-
12
#644100000000
0!
0%
b101 *
0-
02
b101 6
#644110000000
1!
1%
1-
12
#644120000000
0!
0%
b110 *
0-
02
b110 6
#644130000000
1!
1%
1-
12
#644140000000
0!
0%
b111 *
0-
02
b111 6
#644150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#644160000000
0!
0%
b0 *
0-
02
b0 6
#644170000000
1!
1%
1-
12
#644180000000
0!
0%
b1 *
0-
02
b1 6
#644190000000
1!
1%
1-
12
#644200000000
0!
0%
b10 *
0-
02
b10 6
#644210000000
1!
1%
1-
12
#644220000000
0!
0%
b11 *
0-
02
b11 6
#644230000000
1!
1%
1-
12
15
#644240000000
0!
0%
b100 *
0-
02
b100 6
#644250000000
1!
1%
1-
12
#644260000000
0!
0%
b101 *
0-
02
b101 6
#644270000000
1!
1%
1-
12
#644280000000
0!
0%
b110 *
0-
02
b110 6
#644290000000
1!
1%
1-
12
#644300000000
0!
0%
b111 *
0-
02
b111 6
#644310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#644320000000
0!
0%
b0 *
0-
02
b0 6
#644330000000
1!
1%
1-
12
#644340000000
0!
0%
b1 *
0-
02
b1 6
#644350000000
1!
1%
1-
12
#644360000000
0!
0%
b10 *
0-
02
b10 6
#644370000000
1!
1%
1-
12
#644380000000
0!
0%
b11 *
0-
02
b11 6
#644390000000
1!
1%
1-
12
15
#644400000000
0!
0%
b100 *
0-
02
b100 6
#644410000000
1!
1%
1-
12
#644420000000
0!
0%
b101 *
0-
02
b101 6
#644430000000
1!
1%
1-
12
#644440000000
0!
0%
b110 *
0-
02
b110 6
#644450000000
1!
1%
1-
12
#644460000000
0!
0%
b111 *
0-
02
b111 6
#644470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#644480000000
0!
0%
b0 *
0-
02
b0 6
#644490000000
1!
1%
1-
12
#644500000000
0!
0%
b1 *
0-
02
b1 6
#644510000000
1!
1%
1-
12
#644520000000
0!
0%
b10 *
0-
02
b10 6
#644530000000
1!
1%
1-
12
#644540000000
0!
0%
b11 *
0-
02
b11 6
#644550000000
1!
1%
1-
12
15
#644560000000
0!
0%
b100 *
0-
02
b100 6
#644570000000
1!
1%
1-
12
#644580000000
0!
0%
b101 *
0-
02
b101 6
#644590000000
1!
1%
1-
12
#644600000000
0!
0%
b110 *
0-
02
b110 6
#644610000000
1!
1%
1-
12
#644620000000
0!
0%
b111 *
0-
02
b111 6
#644630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#644640000000
0!
0%
b0 *
0-
02
b0 6
#644650000000
1!
1%
1-
12
#644660000000
0!
0%
b1 *
0-
02
b1 6
#644670000000
1!
1%
1-
12
#644680000000
0!
0%
b10 *
0-
02
b10 6
#644690000000
1!
1%
1-
12
#644700000000
0!
0%
b11 *
0-
02
b11 6
#644710000000
1!
1%
1-
12
15
#644720000000
0!
0%
b100 *
0-
02
b100 6
#644730000000
1!
1%
1-
12
#644740000000
0!
0%
b101 *
0-
02
b101 6
#644750000000
1!
1%
1-
12
#644760000000
0!
0%
b110 *
0-
02
b110 6
#644770000000
1!
1%
1-
12
#644780000000
0!
0%
b111 *
0-
02
b111 6
#644790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#644800000000
0!
0%
b0 *
0-
02
b0 6
#644810000000
1!
1%
1-
12
#644820000000
0!
0%
b1 *
0-
02
b1 6
#644830000000
1!
1%
1-
12
#644840000000
0!
0%
b10 *
0-
02
b10 6
#644850000000
1!
1%
1-
12
#644860000000
0!
0%
b11 *
0-
02
b11 6
#644870000000
1!
1%
1-
12
15
#644880000000
0!
0%
b100 *
0-
02
b100 6
#644890000000
1!
1%
1-
12
#644900000000
0!
0%
b101 *
0-
02
b101 6
#644910000000
1!
1%
1-
12
#644920000000
0!
0%
b110 *
0-
02
b110 6
#644930000000
1!
1%
1-
12
#644940000000
0!
0%
b111 *
0-
02
b111 6
#644950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#644960000000
0!
0%
b0 *
0-
02
b0 6
#644970000000
1!
1%
1-
12
#644980000000
0!
0%
b1 *
0-
02
b1 6
#644990000000
1!
1%
1-
12
#645000000000
0!
0%
b10 *
0-
02
b10 6
#645010000000
1!
1%
1-
12
#645020000000
0!
0%
b11 *
0-
02
b11 6
#645030000000
1!
1%
1-
12
15
#645040000000
0!
0%
b100 *
0-
02
b100 6
#645050000000
1!
1%
1-
12
#645060000000
0!
0%
b101 *
0-
02
b101 6
#645070000000
1!
1%
1-
12
#645080000000
0!
0%
b110 *
0-
02
b110 6
#645090000000
1!
1%
1-
12
#645100000000
0!
0%
b111 *
0-
02
b111 6
#645110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#645120000000
0!
0%
b0 *
0-
02
b0 6
#645130000000
1!
1%
1-
12
#645140000000
0!
0%
b1 *
0-
02
b1 6
#645150000000
1!
1%
1-
12
#645160000000
0!
0%
b10 *
0-
02
b10 6
#645170000000
1!
1%
1-
12
#645180000000
0!
0%
b11 *
0-
02
b11 6
#645190000000
1!
1%
1-
12
15
#645200000000
0!
0%
b100 *
0-
02
b100 6
#645210000000
1!
1%
1-
12
#645220000000
0!
0%
b101 *
0-
02
b101 6
#645230000000
1!
1%
1-
12
#645240000000
0!
0%
b110 *
0-
02
b110 6
#645250000000
1!
1%
1-
12
#645260000000
0!
0%
b111 *
0-
02
b111 6
#645270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#645280000000
0!
0%
b0 *
0-
02
b0 6
#645290000000
1!
1%
1-
12
#645300000000
0!
0%
b1 *
0-
02
b1 6
#645310000000
1!
1%
1-
12
#645320000000
0!
0%
b10 *
0-
02
b10 6
#645330000000
1!
1%
1-
12
#645340000000
0!
0%
b11 *
0-
02
b11 6
#645350000000
1!
1%
1-
12
15
#645360000000
0!
0%
b100 *
0-
02
b100 6
#645370000000
1!
1%
1-
12
#645380000000
0!
0%
b101 *
0-
02
b101 6
#645390000000
1!
1%
1-
12
#645400000000
0!
0%
b110 *
0-
02
b110 6
#645410000000
1!
1%
1-
12
#645420000000
0!
0%
b111 *
0-
02
b111 6
#645430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#645440000000
0!
0%
b0 *
0-
02
b0 6
#645450000000
1!
1%
1-
12
#645460000000
0!
0%
b1 *
0-
02
b1 6
#645470000000
1!
1%
1-
12
#645480000000
0!
0%
b10 *
0-
02
b10 6
#645490000000
1!
1%
1-
12
#645500000000
0!
0%
b11 *
0-
02
b11 6
#645510000000
1!
1%
1-
12
15
#645520000000
0!
0%
b100 *
0-
02
b100 6
#645530000000
1!
1%
1-
12
#645540000000
0!
0%
b101 *
0-
02
b101 6
#645550000000
1!
1%
1-
12
#645560000000
0!
0%
b110 *
0-
02
b110 6
#645570000000
1!
1%
1-
12
#645580000000
0!
0%
b111 *
0-
02
b111 6
#645590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#645600000000
0!
0%
b0 *
0-
02
b0 6
#645610000000
1!
1%
1-
12
#645620000000
0!
0%
b1 *
0-
02
b1 6
#645630000000
1!
1%
1-
12
#645640000000
0!
0%
b10 *
0-
02
b10 6
#645650000000
1!
1%
1-
12
#645660000000
0!
0%
b11 *
0-
02
b11 6
#645670000000
1!
1%
1-
12
15
#645680000000
0!
0%
b100 *
0-
02
b100 6
#645690000000
1!
1%
1-
12
#645700000000
0!
0%
b101 *
0-
02
b101 6
#645710000000
1!
1%
1-
12
#645720000000
0!
0%
b110 *
0-
02
b110 6
#645730000000
1!
1%
1-
12
#645740000000
0!
0%
b111 *
0-
02
b111 6
#645750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#645760000000
0!
0%
b0 *
0-
02
b0 6
#645770000000
1!
1%
1-
12
#645780000000
0!
0%
b1 *
0-
02
b1 6
#645790000000
1!
1%
1-
12
#645800000000
0!
0%
b10 *
0-
02
b10 6
#645810000000
1!
1%
1-
12
#645820000000
0!
0%
b11 *
0-
02
b11 6
#645830000000
1!
1%
1-
12
15
#645840000000
0!
0%
b100 *
0-
02
b100 6
#645850000000
1!
1%
1-
12
#645860000000
0!
0%
b101 *
0-
02
b101 6
#645870000000
1!
1%
1-
12
#645880000000
0!
0%
b110 *
0-
02
b110 6
#645890000000
1!
1%
1-
12
#645900000000
0!
0%
b111 *
0-
02
b111 6
#645910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#645920000000
0!
0%
b0 *
0-
02
b0 6
#645930000000
1!
1%
1-
12
#645940000000
0!
0%
b1 *
0-
02
b1 6
#645950000000
1!
1%
1-
12
#645960000000
0!
0%
b10 *
0-
02
b10 6
#645970000000
1!
1%
1-
12
#645980000000
0!
0%
b11 *
0-
02
b11 6
#645990000000
1!
1%
1-
12
15
#646000000000
0!
0%
b100 *
0-
02
b100 6
#646010000000
1!
1%
1-
12
#646020000000
0!
0%
b101 *
0-
02
b101 6
#646030000000
1!
1%
1-
12
#646040000000
0!
0%
b110 *
0-
02
b110 6
#646050000000
1!
1%
1-
12
#646060000000
0!
0%
b111 *
0-
02
b111 6
#646070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#646080000000
0!
0%
b0 *
0-
02
b0 6
#646090000000
1!
1%
1-
12
#646100000000
0!
0%
b1 *
0-
02
b1 6
#646110000000
1!
1%
1-
12
#646120000000
0!
0%
b10 *
0-
02
b10 6
#646130000000
1!
1%
1-
12
#646140000000
0!
0%
b11 *
0-
02
b11 6
#646150000000
1!
1%
1-
12
15
#646160000000
0!
0%
b100 *
0-
02
b100 6
#646170000000
1!
1%
1-
12
#646180000000
0!
0%
b101 *
0-
02
b101 6
#646190000000
1!
1%
1-
12
#646200000000
0!
0%
b110 *
0-
02
b110 6
#646210000000
1!
1%
1-
12
#646220000000
0!
0%
b111 *
0-
02
b111 6
#646230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#646240000000
0!
0%
b0 *
0-
02
b0 6
#646250000000
1!
1%
1-
12
#646260000000
0!
0%
b1 *
0-
02
b1 6
#646270000000
1!
1%
1-
12
#646280000000
0!
0%
b10 *
0-
02
b10 6
#646290000000
1!
1%
1-
12
#646300000000
0!
0%
b11 *
0-
02
b11 6
#646310000000
1!
1%
1-
12
15
#646320000000
0!
0%
b100 *
0-
02
b100 6
#646330000000
1!
1%
1-
12
#646340000000
0!
0%
b101 *
0-
02
b101 6
#646350000000
1!
1%
1-
12
#646360000000
0!
0%
b110 *
0-
02
b110 6
#646370000000
1!
1%
1-
12
#646380000000
0!
0%
b111 *
0-
02
b111 6
#646390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#646400000000
0!
0%
b0 *
0-
02
b0 6
#646410000000
1!
1%
1-
12
#646420000000
0!
0%
b1 *
0-
02
b1 6
#646430000000
1!
1%
1-
12
#646440000000
0!
0%
b10 *
0-
02
b10 6
#646450000000
1!
1%
1-
12
#646460000000
0!
0%
b11 *
0-
02
b11 6
#646470000000
1!
1%
1-
12
15
#646480000000
0!
0%
b100 *
0-
02
b100 6
#646490000000
1!
1%
1-
12
#646500000000
0!
0%
b101 *
0-
02
b101 6
#646510000000
1!
1%
1-
12
#646520000000
0!
0%
b110 *
0-
02
b110 6
#646530000000
1!
1%
1-
12
#646540000000
0!
0%
b111 *
0-
02
b111 6
#646550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#646560000000
0!
0%
b0 *
0-
02
b0 6
#646570000000
1!
1%
1-
12
#646580000000
0!
0%
b1 *
0-
02
b1 6
#646590000000
1!
1%
1-
12
#646600000000
0!
0%
b10 *
0-
02
b10 6
#646610000000
1!
1%
1-
12
#646620000000
0!
0%
b11 *
0-
02
b11 6
#646630000000
1!
1%
1-
12
15
#646640000000
0!
0%
b100 *
0-
02
b100 6
#646650000000
1!
1%
1-
12
#646660000000
0!
0%
b101 *
0-
02
b101 6
#646670000000
1!
1%
1-
12
#646680000000
0!
0%
b110 *
0-
02
b110 6
#646690000000
1!
1%
1-
12
#646700000000
0!
0%
b111 *
0-
02
b111 6
#646710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#646720000000
0!
0%
b0 *
0-
02
b0 6
#646730000000
1!
1%
1-
12
#646740000000
0!
0%
b1 *
0-
02
b1 6
#646750000000
1!
1%
1-
12
#646760000000
0!
0%
b10 *
0-
02
b10 6
#646770000000
1!
1%
1-
12
#646780000000
0!
0%
b11 *
0-
02
b11 6
#646790000000
1!
1%
1-
12
15
#646800000000
0!
0%
b100 *
0-
02
b100 6
#646810000000
1!
1%
1-
12
#646820000000
0!
0%
b101 *
0-
02
b101 6
#646830000000
1!
1%
1-
12
#646840000000
0!
0%
b110 *
0-
02
b110 6
#646850000000
1!
1%
1-
12
#646860000000
0!
0%
b111 *
0-
02
b111 6
#646870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#646880000000
0!
0%
b0 *
0-
02
b0 6
#646890000000
1!
1%
1-
12
#646900000000
0!
0%
b1 *
0-
02
b1 6
#646910000000
1!
1%
1-
12
#646920000000
0!
0%
b10 *
0-
02
b10 6
#646930000000
1!
1%
1-
12
#646940000000
0!
0%
b11 *
0-
02
b11 6
#646950000000
1!
1%
1-
12
15
#646960000000
0!
0%
b100 *
0-
02
b100 6
#646970000000
1!
1%
1-
12
#646980000000
0!
0%
b101 *
0-
02
b101 6
#646990000000
1!
1%
1-
12
#647000000000
0!
0%
b110 *
0-
02
b110 6
#647010000000
1!
1%
1-
12
#647020000000
0!
0%
b111 *
0-
02
b111 6
#647030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#647040000000
0!
0%
b0 *
0-
02
b0 6
#647050000000
1!
1%
1-
12
#647060000000
0!
0%
b1 *
0-
02
b1 6
#647070000000
1!
1%
1-
12
#647080000000
0!
0%
b10 *
0-
02
b10 6
#647090000000
1!
1%
1-
12
#647100000000
0!
0%
b11 *
0-
02
b11 6
#647110000000
1!
1%
1-
12
15
#647120000000
0!
0%
b100 *
0-
02
b100 6
#647130000000
1!
1%
1-
12
#647140000000
0!
0%
b101 *
0-
02
b101 6
#647150000000
1!
1%
1-
12
#647160000000
0!
0%
b110 *
0-
02
b110 6
#647170000000
1!
1%
1-
12
#647180000000
0!
0%
b111 *
0-
02
b111 6
#647190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#647200000000
0!
0%
b0 *
0-
02
b0 6
#647210000000
1!
1%
1-
12
#647220000000
0!
0%
b1 *
0-
02
b1 6
#647230000000
1!
1%
1-
12
#647240000000
0!
0%
b10 *
0-
02
b10 6
#647250000000
1!
1%
1-
12
#647260000000
0!
0%
b11 *
0-
02
b11 6
#647270000000
1!
1%
1-
12
15
#647280000000
0!
0%
b100 *
0-
02
b100 6
#647290000000
1!
1%
1-
12
#647300000000
0!
0%
b101 *
0-
02
b101 6
#647310000000
1!
1%
1-
12
#647320000000
0!
0%
b110 *
0-
02
b110 6
#647330000000
1!
1%
1-
12
#647340000000
0!
0%
b111 *
0-
02
b111 6
#647350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#647360000000
0!
0%
b0 *
0-
02
b0 6
#647370000000
1!
1%
1-
12
#647380000000
0!
0%
b1 *
0-
02
b1 6
#647390000000
1!
1%
1-
12
#647400000000
0!
0%
b10 *
0-
02
b10 6
#647410000000
1!
1%
1-
12
#647420000000
0!
0%
b11 *
0-
02
b11 6
#647430000000
1!
1%
1-
12
15
#647440000000
0!
0%
b100 *
0-
02
b100 6
#647450000000
1!
1%
1-
12
#647460000000
0!
0%
b101 *
0-
02
b101 6
#647470000000
1!
1%
1-
12
#647480000000
0!
0%
b110 *
0-
02
b110 6
#647490000000
1!
1%
1-
12
#647500000000
0!
0%
b111 *
0-
02
b111 6
#647510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#647520000000
0!
0%
b0 *
0-
02
b0 6
#647530000000
1!
1%
1-
12
#647540000000
0!
0%
b1 *
0-
02
b1 6
#647550000000
1!
1%
1-
12
#647560000000
0!
0%
b10 *
0-
02
b10 6
#647570000000
1!
1%
1-
12
#647580000000
0!
0%
b11 *
0-
02
b11 6
#647590000000
1!
1%
1-
12
15
#647600000000
0!
0%
b100 *
0-
02
b100 6
#647610000000
1!
1%
1-
12
#647620000000
0!
0%
b101 *
0-
02
b101 6
#647630000000
1!
1%
1-
12
#647640000000
0!
0%
b110 *
0-
02
b110 6
#647650000000
1!
1%
1-
12
#647660000000
0!
0%
b111 *
0-
02
b111 6
#647670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#647680000000
0!
0%
b0 *
0-
02
b0 6
#647690000000
1!
1%
1-
12
#647700000000
0!
0%
b1 *
0-
02
b1 6
#647710000000
1!
1%
1-
12
#647720000000
0!
0%
b10 *
0-
02
b10 6
#647730000000
1!
1%
1-
12
#647740000000
0!
0%
b11 *
0-
02
b11 6
#647750000000
1!
1%
1-
12
15
#647760000000
0!
0%
b100 *
0-
02
b100 6
#647770000000
1!
1%
1-
12
#647780000000
0!
0%
b101 *
0-
02
b101 6
#647790000000
1!
1%
1-
12
#647800000000
0!
0%
b110 *
0-
02
b110 6
#647810000000
1!
1%
1-
12
#647820000000
0!
0%
b111 *
0-
02
b111 6
#647830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#647840000000
0!
0%
b0 *
0-
02
b0 6
#647850000000
1!
1%
1-
12
#647860000000
0!
0%
b1 *
0-
02
b1 6
#647870000000
1!
1%
1-
12
#647880000000
0!
0%
b10 *
0-
02
b10 6
#647890000000
1!
1%
1-
12
#647900000000
0!
0%
b11 *
0-
02
b11 6
#647910000000
1!
1%
1-
12
15
#647920000000
0!
0%
b100 *
0-
02
b100 6
#647930000000
1!
1%
1-
12
#647940000000
0!
0%
b101 *
0-
02
b101 6
#647950000000
1!
1%
1-
12
#647960000000
0!
0%
b110 *
0-
02
b110 6
#647970000000
1!
1%
1-
12
#647980000000
0!
0%
b111 *
0-
02
b111 6
#647990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#648000000000
0!
0%
b0 *
0-
02
b0 6
#648010000000
1!
1%
1-
12
#648020000000
0!
0%
b1 *
0-
02
b1 6
#648030000000
1!
1%
1-
12
#648040000000
0!
0%
b10 *
0-
02
b10 6
#648050000000
1!
1%
1-
12
#648060000000
0!
0%
b11 *
0-
02
b11 6
#648070000000
1!
1%
1-
12
15
#648080000000
0!
0%
b100 *
0-
02
b100 6
#648090000000
1!
1%
1-
12
#648100000000
0!
0%
b101 *
0-
02
b101 6
#648110000000
1!
1%
1-
12
#648120000000
0!
0%
b110 *
0-
02
b110 6
#648130000000
1!
1%
1-
12
#648140000000
0!
0%
b111 *
0-
02
b111 6
#648150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#648160000000
0!
0%
b0 *
0-
02
b0 6
#648170000000
1!
1%
1-
12
#648180000000
0!
0%
b1 *
0-
02
b1 6
#648190000000
1!
1%
1-
12
#648200000000
0!
0%
b10 *
0-
02
b10 6
#648210000000
1!
1%
1-
12
#648220000000
0!
0%
b11 *
0-
02
b11 6
#648230000000
1!
1%
1-
12
15
#648240000000
0!
0%
b100 *
0-
02
b100 6
#648250000000
1!
1%
1-
12
#648260000000
0!
0%
b101 *
0-
02
b101 6
#648270000000
1!
1%
1-
12
#648280000000
0!
0%
b110 *
0-
02
b110 6
#648290000000
1!
1%
1-
12
#648300000000
0!
0%
b111 *
0-
02
b111 6
#648310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#648320000000
0!
0%
b0 *
0-
02
b0 6
#648330000000
1!
1%
1-
12
#648340000000
0!
0%
b1 *
0-
02
b1 6
#648350000000
1!
1%
1-
12
#648360000000
0!
0%
b10 *
0-
02
b10 6
#648370000000
1!
1%
1-
12
#648380000000
0!
0%
b11 *
0-
02
b11 6
#648390000000
1!
1%
1-
12
15
#648400000000
0!
0%
b100 *
0-
02
b100 6
#648410000000
1!
1%
1-
12
#648420000000
0!
0%
b101 *
0-
02
b101 6
#648430000000
1!
1%
1-
12
#648440000000
0!
0%
b110 *
0-
02
b110 6
#648450000000
1!
1%
1-
12
#648460000000
0!
0%
b111 *
0-
02
b111 6
#648470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#648480000000
0!
0%
b0 *
0-
02
b0 6
#648490000000
1!
1%
1-
12
#648500000000
0!
0%
b1 *
0-
02
b1 6
#648510000000
1!
1%
1-
12
#648520000000
0!
0%
b10 *
0-
02
b10 6
#648530000000
1!
1%
1-
12
#648540000000
0!
0%
b11 *
0-
02
b11 6
#648550000000
1!
1%
1-
12
15
#648560000000
0!
0%
b100 *
0-
02
b100 6
#648570000000
1!
1%
1-
12
#648580000000
0!
0%
b101 *
0-
02
b101 6
#648590000000
1!
1%
1-
12
#648600000000
0!
0%
b110 *
0-
02
b110 6
#648610000000
1!
1%
1-
12
#648620000000
0!
0%
b111 *
0-
02
b111 6
#648630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#648640000000
0!
0%
b0 *
0-
02
b0 6
#648650000000
1!
1%
1-
12
#648660000000
0!
0%
b1 *
0-
02
b1 6
#648670000000
1!
1%
1-
12
#648680000000
0!
0%
b10 *
0-
02
b10 6
#648690000000
1!
1%
1-
12
#648700000000
0!
0%
b11 *
0-
02
b11 6
#648710000000
1!
1%
1-
12
15
#648720000000
0!
0%
b100 *
0-
02
b100 6
#648730000000
1!
1%
1-
12
#648740000000
0!
0%
b101 *
0-
02
b101 6
#648750000000
1!
1%
1-
12
#648760000000
0!
0%
b110 *
0-
02
b110 6
#648770000000
1!
1%
1-
12
#648780000000
0!
0%
b111 *
0-
02
b111 6
#648790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#648800000000
0!
0%
b0 *
0-
02
b0 6
#648810000000
1!
1%
1-
12
#648820000000
0!
0%
b1 *
0-
02
b1 6
#648830000000
1!
1%
1-
12
#648840000000
0!
0%
b10 *
0-
02
b10 6
#648850000000
1!
1%
1-
12
#648860000000
0!
0%
b11 *
0-
02
b11 6
#648870000000
1!
1%
1-
12
15
#648880000000
0!
0%
b100 *
0-
02
b100 6
#648890000000
1!
1%
1-
12
#648900000000
0!
0%
b101 *
0-
02
b101 6
#648910000000
1!
1%
1-
12
#648920000000
0!
0%
b110 *
0-
02
b110 6
#648930000000
1!
1%
1-
12
#648940000000
0!
0%
b111 *
0-
02
b111 6
#648950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#648960000000
0!
0%
b0 *
0-
02
b0 6
#648970000000
1!
1%
1-
12
#648980000000
0!
0%
b1 *
0-
02
b1 6
#648990000000
1!
1%
1-
12
#649000000000
0!
0%
b10 *
0-
02
b10 6
#649010000000
1!
1%
1-
12
#649020000000
0!
0%
b11 *
0-
02
b11 6
#649030000000
1!
1%
1-
12
15
#649040000000
0!
0%
b100 *
0-
02
b100 6
#649050000000
1!
1%
1-
12
#649060000000
0!
0%
b101 *
0-
02
b101 6
#649070000000
1!
1%
1-
12
#649080000000
0!
0%
b110 *
0-
02
b110 6
#649090000000
1!
1%
1-
12
#649100000000
0!
0%
b111 *
0-
02
b111 6
#649110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#649120000000
0!
0%
b0 *
0-
02
b0 6
#649130000000
1!
1%
1-
12
#649140000000
0!
0%
b1 *
0-
02
b1 6
#649150000000
1!
1%
1-
12
#649160000000
0!
0%
b10 *
0-
02
b10 6
#649170000000
1!
1%
1-
12
#649180000000
0!
0%
b11 *
0-
02
b11 6
#649190000000
1!
1%
1-
12
15
#649200000000
0!
0%
b100 *
0-
02
b100 6
#649210000000
1!
1%
1-
12
#649220000000
0!
0%
b101 *
0-
02
b101 6
#649230000000
1!
1%
1-
12
#649240000000
0!
0%
b110 *
0-
02
b110 6
#649250000000
1!
1%
1-
12
#649260000000
0!
0%
b111 *
0-
02
b111 6
#649270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#649280000000
0!
0%
b0 *
0-
02
b0 6
#649290000000
1!
1%
1-
12
#649300000000
0!
0%
b1 *
0-
02
b1 6
#649310000000
1!
1%
1-
12
#649320000000
0!
0%
b10 *
0-
02
b10 6
#649330000000
1!
1%
1-
12
#649340000000
0!
0%
b11 *
0-
02
b11 6
#649350000000
1!
1%
1-
12
15
#649360000000
0!
0%
b100 *
0-
02
b100 6
#649370000000
1!
1%
1-
12
#649380000000
0!
0%
b101 *
0-
02
b101 6
#649390000000
1!
1%
1-
12
#649400000000
0!
0%
b110 *
0-
02
b110 6
#649410000000
1!
1%
1-
12
#649420000000
0!
0%
b111 *
0-
02
b111 6
#649430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#649440000000
0!
0%
b0 *
0-
02
b0 6
#649450000000
1!
1%
1-
12
#649460000000
0!
0%
b1 *
0-
02
b1 6
#649470000000
1!
1%
1-
12
#649480000000
0!
0%
b10 *
0-
02
b10 6
#649490000000
1!
1%
1-
12
#649500000000
0!
0%
b11 *
0-
02
b11 6
#649510000000
1!
1%
1-
12
15
#649520000000
0!
0%
b100 *
0-
02
b100 6
#649530000000
1!
1%
1-
12
#649540000000
0!
0%
b101 *
0-
02
b101 6
#649550000000
1!
1%
1-
12
#649560000000
0!
0%
b110 *
0-
02
b110 6
#649570000000
1!
1%
1-
12
#649580000000
0!
0%
b111 *
0-
02
b111 6
#649590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#649600000000
0!
0%
b0 *
0-
02
b0 6
#649610000000
1!
1%
1-
12
#649620000000
0!
0%
b1 *
0-
02
b1 6
#649630000000
1!
1%
1-
12
#649640000000
0!
0%
b10 *
0-
02
b10 6
#649650000000
1!
1%
1-
12
#649660000000
0!
0%
b11 *
0-
02
b11 6
#649670000000
1!
1%
1-
12
15
#649680000000
0!
0%
b100 *
0-
02
b100 6
#649690000000
1!
1%
1-
12
#649700000000
0!
0%
b101 *
0-
02
b101 6
#649710000000
1!
1%
1-
12
#649720000000
0!
0%
b110 *
0-
02
b110 6
#649730000000
1!
1%
1-
12
#649740000000
0!
0%
b111 *
0-
02
b111 6
#649750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#649760000000
0!
0%
b0 *
0-
02
b0 6
#649770000000
1!
1%
1-
12
#649780000000
0!
0%
b1 *
0-
02
b1 6
#649790000000
1!
1%
1-
12
#649800000000
0!
0%
b10 *
0-
02
b10 6
#649810000000
1!
1%
1-
12
#649820000000
0!
0%
b11 *
0-
02
b11 6
#649830000000
1!
1%
1-
12
15
#649840000000
0!
0%
b100 *
0-
02
b100 6
#649850000000
1!
1%
1-
12
#649860000000
0!
0%
b101 *
0-
02
b101 6
#649870000000
1!
1%
1-
12
#649880000000
0!
0%
b110 *
0-
02
b110 6
#649890000000
1!
1%
1-
12
#649900000000
0!
0%
b111 *
0-
02
b111 6
#649910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#649920000000
0!
0%
b0 *
0-
02
b0 6
#649930000000
1!
1%
1-
12
#649940000000
0!
0%
b1 *
0-
02
b1 6
#649950000000
1!
1%
1-
12
#649960000000
0!
0%
b10 *
0-
02
b10 6
#649970000000
1!
1%
1-
12
#649980000000
0!
0%
b11 *
0-
02
b11 6
#649990000000
1!
1%
1-
12
15
#650000000000
0!
0%
b100 *
0-
02
b100 6
#650010000000
1!
1%
1-
12
#650020000000
0!
0%
b101 *
0-
02
b101 6
#650030000000
1!
1%
1-
12
#650040000000
0!
0%
b110 *
0-
02
b110 6
#650050000000
1!
1%
1-
12
#650060000000
0!
0%
b111 *
0-
02
b111 6
#650070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#650080000000
0!
0%
b0 *
0-
02
b0 6
#650090000000
1!
1%
1-
12
#650100000000
0!
0%
b1 *
0-
02
b1 6
#650110000000
1!
1%
1-
12
#650120000000
0!
0%
b10 *
0-
02
b10 6
#650130000000
1!
1%
1-
12
#650140000000
0!
0%
b11 *
0-
02
b11 6
#650150000000
1!
1%
1-
12
15
#650160000000
0!
0%
b100 *
0-
02
b100 6
#650170000000
1!
1%
1-
12
#650180000000
0!
0%
b101 *
0-
02
b101 6
#650190000000
1!
1%
1-
12
#650200000000
0!
0%
b110 *
0-
02
b110 6
#650210000000
1!
1%
1-
12
#650220000000
0!
0%
b111 *
0-
02
b111 6
#650230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#650240000000
0!
0%
b0 *
0-
02
b0 6
#650250000000
1!
1%
1-
12
#650260000000
0!
0%
b1 *
0-
02
b1 6
#650270000000
1!
1%
1-
12
#650280000000
0!
0%
b10 *
0-
02
b10 6
#650290000000
1!
1%
1-
12
#650300000000
0!
0%
b11 *
0-
02
b11 6
#650310000000
1!
1%
1-
12
15
#650320000000
0!
0%
b100 *
0-
02
b100 6
#650330000000
1!
1%
1-
12
#650340000000
0!
0%
b101 *
0-
02
b101 6
#650350000000
1!
1%
1-
12
#650360000000
0!
0%
b110 *
0-
02
b110 6
#650370000000
1!
1%
1-
12
#650380000000
0!
0%
b111 *
0-
02
b111 6
#650390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#650400000000
0!
0%
b0 *
0-
02
b0 6
#650410000000
1!
1%
1-
12
#650420000000
0!
0%
b1 *
0-
02
b1 6
#650430000000
1!
1%
1-
12
#650440000000
0!
0%
b10 *
0-
02
b10 6
#650450000000
1!
1%
1-
12
#650460000000
0!
0%
b11 *
0-
02
b11 6
#650470000000
1!
1%
1-
12
15
#650480000000
0!
0%
b100 *
0-
02
b100 6
#650490000000
1!
1%
1-
12
#650500000000
0!
0%
b101 *
0-
02
b101 6
#650510000000
1!
1%
1-
12
#650520000000
0!
0%
b110 *
0-
02
b110 6
#650530000000
1!
1%
1-
12
#650540000000
0!
0%
b111 *
0-
02
b111 6
#650550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#650560000000
0!
0%
b0 *
0-
02
b0 6
#650570000000
1!
1%
1-
12
#650580000000
0!
0%
b1 *
0-
02
b1 6
#650590000000
1!
1%
1-
12
#650600000000
0!
0%
b10 *
0-
02
b10 6
#650610000000
1!
1%
1-
12
#650620000000
0!
0%
b11 *
0-
02
b11 6
#650630000000
1!
1%
1-
12
15
#650640000000
0!
0%
b100 *
0-
02
b100 6
#650650000000
1!
1%
1-
12
#650660000000
0!
0%
b101 *
0-
02
b101 6
#650670000000
1!
1%
1-
12
#650680000000
0!
0%
b110 *
0-
02
b110 6
#650690000000
1!
1%
1-
12
#650700000000
0!
0%
b111 *
0-
02
b111 6
#650710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#650720000000
0!
0%
b0 *
0-
02
b0 6
#650730000000
1!
1%
1-
12
#650740000000
0!
0%
b1 *
0-
02
b1 6
#650750000000
1!
1%
1-
12
#650760000000
0!
0%
b10 *
0-
02
b10 6
#650770000000
1!
1%
1-
12
#650780000000
0!
0%
b11 *
0-
02
b11 6
#650790000000
1!
1%
1-
12
15
#650800000000
0!
0%
b100 *
0-
02
b100 6
#650810000000
1!
1%
1-
12
#650820000000
0!
0%
b101 *
0-
02
b101 6
#650830000000
1!
1%
1-
12
#650840000000
0!
0%
b110 *
0-
02
b110 6
#650850000000
1!
1%
1-
12
#650860000000
0!
0%
b111 *
0-
02
b111 6
#650870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#650880000000
0!
0%
b0 *
0-
02
b0 6
#650890000000
1!
1%
1-
12
#650900000000
0!
0%
b1 *
0-
02
b1 6
#650910000000
1!
1%
1-
12
#650920000000
0!
0%
b10 *
0-
02
b10 6
#650930000000
1!
1%
1-
12
#650940000000
0!
0%
b11 *
0-
02
b11 6
#650950000000
1!
1%
1-
12
15
#650960000000
0!
0%
b100 *
0-
02
b100 6
#650970000000
1!
1%
1-
12
#650980000000
0!
0%
b101 *
0-
02
b101 6
#650990000000
1!
1%
1-
12
#651000000000
0!
0%
b110 *
0-
02
b110 6
#651010000000
1!
1%
1-
12
#651020000000
0!
0%
b111 *
0-
02
b111 6
#651030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#651040000000
0!
0%
b0 *
0-
02
b0 6
#651050000000
1!
1%
1-
12
#651060000000
0!
0%
b1 *
0-
02
b1 6
#651070000000
1!
1%
1-
12
#651080000000
0!
0%
b10 *
0-
02
b10 6
#651090000000
1!
1%
1-
12
#651100000000
0!
0%
b11 *
0-
02
b11 6
#651110000000
1!
1%
1-
12
15
#651120000000
0!
0%
b100 *
0-
02
b100 6
#651130000000
1!
1%
1-
12
#651140000000
0!
0%
b101 *
0-
02
b101 6
#651150000000
1!
1%
1-
12
#651160000000
0!
0%
b110 *
0-
02
b110 6
#651170000000
1!
1%
1-
12
#651180000000
0!
0%
b111 *
0-
02
b111 6
#651190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#651200000000
0!
0%
b0 *
0-
02
b0 6
#651210000000
1!
1%
1-
12
#651220000000
0!
0%
b1 *
0-
02
b1 6
#651230000000
1!
1%
1-
12
#651240000000
0!
0%
b10 *
0-
02
b10 6
#651250000000
1!
1%
1-
12
#651260000000
0!
0%
b11 *
0-
02
b11 6
#651270000000
1!
1%
1-
12
15
#651280000000
0!
0%
b100 *
0-
02
b100 6
#651290000000
1!
1%
1-
12
#651300000000
0!
0%
b101 *
0-
02
b101 6
#651310000000
1!
1%
1-
12
#651320000000
0!
0%
b110 *
0-
02
b110 6
#651330000000
1!
1%
1-
12
#651340000000
0!
0%
b111 *
0-
02
b111 6
#651350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#651360000000
0!
0%
b0 *
0-
02
b0 6
#651370000000
1!
1%
1-
12
#651380000000
0!
0%
b1 *
0-
02
b1 6
#651390000000
1!
1%
1-
12
#651400000000
0!
0%
b10 *
0-
02
b10 6
#651410000000
1!
1%
1-
12
#651420000000
0!
0%
b11 *
0-
02
b11 6
#651430000000
1!
1%
1-
12
15
#651440000000
0!
0%
b100 *
0-
02
b100 6
#651450000000
1!
1%
1-
12
#651460000000
0!
0%
b101 *
0-
02
b101 6
#651470000000
1!
1%
1-
12
#651480000000
0!
0%
b110 *
0-
02
b110 6
#651490000000
1!
1%
1-
12
#651500000000
0!
0%
b111 *
0-
02
b111 6
#651510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#651520000000
0!
0%
b0 *
0-
02
b0 6
#651530000000
1!
1%
1-
12
#651540000000
0!
0%
b1 *
0-
02
b1 6
#651550000000
1!
1%
1-
12
#651560000000
0!
0%
b10 *
0-
02
b10 6
#651570000000
1!
1%
1-
12
#651580000000
0!
0%
b11 *
0-
02
b11 6
#651590000000
1!
1%
1-
12
15
#651600000000
0!
0%
b100 *
0-
02
b100 6
#651610000000
1!
1%
1-
12
#651620000000
0!
0%
b101 *
0-
02
b101 6
#651630000000
1!
1%
1-
12
#651640000000
0!
0%
b110 *
0-
02
b110 6
#651650000000
1!
1%
1-
12
#651660000000
0!
0%
b111 *
0-
02
b111 6
#651670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#651680000000
0!
0%
b0 *
0-
02
b0 6
#651690000000
1!
1%
1-
12
#651700000000
0!
0%
b1 *
0-
02
b1 6
#651710000000
1!
1%
1-
12
#651720000000
0!
0%
b10 *
0-
02
b10 6
#651730000000
1!
1%
1-
12
#651740000000
0!
0%
b11 *
0-
02
b11 6
#651750000000
1!
1%
1-
12
15
#651760000000
0!
0%
b100 *
0-
02
b100 6
#651770000000
1!
1%
1-
12
#651780000000
0!
0%
b101 *
0-
02
b101 6
#651790000000
1!
1%
1-
12
#651800000000
0!
0%
b110 *
0-
02
b110 6
#651810000000
1!
1%
1-
12
#651820000000
0!
0%
b111 *
0-
02
b111 6
#651830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#651840000000
0!
0%
b0 *
0-
02
b0 6
#651850000000
1!
1%
1-
12
#651860000000
0!
0%
b1 *
0-
02
b1 6
#651870000000
1!
1%
1-
12
#651880000000
0!
0%
b10 *
0-
02
b10 6
#651890000000
1!
1%
1-
12
#651900000000
0!
0%
b11 *
0-
02
b11 6
#651910000000
1!
1%
1-
12
15
#651920000000
0!
0%
b100 *
0-
02
b100 6
#651930000000
1!
1%
1-
12
#651940000000
0!
0%
b101 *
0-
02
b101 6
#651950000000
1!
1%
1-
12
#651960000000
0!
0%
b110 *
0-
02
b110 6
#651970000000
1!
1%
1-
12
#651980000000
0!
0%
b111 *
0-
02
b111 6
#651990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#652000000000
0!
0%
b0 *
0-
02
b0 6
#652010000000
1!
1%
1-
12
#652020000000
0!
0%
b1 *
0-
02
b1 6
#652030000000
1!
1%
1-
12
#652040000000
0!
0%
b10 *
0-
02
b10 6
#652050000000
1!
1%
1-
12
#652060000000
0!
0%
b11 *
0-
02
b11 6
#652070000000
1!
1%
1-
12
15
#652080000000
0!
0%
b100 *
0-
02
b100 6
#652090000000
1!
1%
1-
12
#652100000000
0!
0%
b101 *
0-
02
b101 6
#652110000000
1!
1%
1-
12
#652120000000
0!
0%
b110 *
0-
02
b110 6
#652130000000
1!
1%
1-
12
#652140000000
0!
0%
b111 *
0-
02
b111 6
#652150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#652160000000
0!
0%
b0 *
0-
02
b0 6
#652170000000
1!
1%
1-
12
#652180000000
0!
0%
b1 *
0-
02
b1 6
#652190000000
1!
1%
1-
12
#652200000000
0!
0%
b10 *
0-
02
b10 6
#652210000000
1!
1%
1-
12
#652220000000
0!
0%
b11 *
0-
02
b11 6
#652230000000
1!
1%
1-
12
15
#652240000000
0!
0%
b100 *
0-
02
b100 6
#652250000000
1!
1%
1-
12
#652260000000
0!
0%
b101 *
0-
02
b101 6
#652270000000
1!
1%
1-
12
#652280000000
0!
0%
b110 *
0-
02
b110 6
#652290000000
1!
1%
1-
12
#652300000000
0!
0%
b111 *
0-
02
b111 6
#652310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#652320000000
0!
0%
b0 *
0-
02
b0 6
#652330000000
1!
1%
1-
12
#652340000000
0!
0%
b1 *
0-
02
b1 6
#652350000000
1!
1%
1-
12
#652360000000
0!
0%
b10 *
0-
02
b10 6
#652370000000
1!
1%
1-
12
#652380000000
0!
0%
b11 *
0-
02
b11 6
#652390000000
1!
1%
1-
12
15
#652400000000
0!
0%
b100 *
0-
02
b100 6
#652410000000
1!
1%
1-
12
#652420000000
0!
0%
b101 *
0-
02
b101 6
#652430000000
1!
1%
1-
12
#652440000000
0!
0%
b110 *
0-
02
b110 6
#652450000000
1!
1%
1-
12
#652460000000
0!
0%
b111 *
0-
02
b111 6
#652470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#652480000000
0!
0%
b0 *
0-
02
b0 6
#652490000000
1!
1%
1-
12
#652500000000
0!
0%
b1 *
0-
02
b1 6
#652510000000
1!
1%
1-
12
#652520000000
0!
0%
b10 *
0-
02
b10 6
#652530000000
1!
1%
1-
12
#652540000000
0!
0%
b11 *
0-
02
b11 6
#652550000000
1!
1%
1-
12
15
#652560000000
0!
0%
b100 *
0-
02
b100 6
#652570000000
1!
1%
1-
12
#652580000000
0!
0%
b101 *
0-
02
b101 6
#652590000000
1!
1%
1-
12
#652600000000
0!
0%
b110 *
0-
02
b110 6
#652610000000
1!
1%
1-
12
#652620000000
0!
0%
b111 *
0-
02
b111 6
#652630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#652640000000
0!
0%
b0 *
0-
02
b0 6
#652650000000
1!
1%
1-
12
#652660000000
0!
0%
b1 *
0-
02
b1 6
#652670000000
1!
1%
1-
12
#652680000000
0!
0%
b10 *
0-
02
b10 6
#652690000000
1!
1%
1-
12
#652700000000
0!
0%
b11 *
0-
02
b11 6
#652710000000
1!
1%
1-
12
15
#652720000000
0!
0%
b100 *
0-
02
b100 6
#652730000000
1!
1%
1-
12
#652740000000
0!
0%
b101 *
0-
02
b101 6
#652750000000
1!
1%
1-
12
#652760000000
0!
0%
b110 *
0-
02
b110 6
#652770000000
1!
1%
1-
12
#652780000000
0!
0%
b111 *
0-
02
b111 6
#652790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#652800000000
0!
0%
b0 *
0-
02
b0 6
#652810000000
1!
1%
1-
12
#652820000000
0!
0%
b1 *
0-
02
b1 6
#652830000000
1!
1%
1-
12
#652840000000
0!
0%
b10 *
0-
02
b10 6
#652850000000
1!
1%
1-
12
#652860000000
0!
0%
b11 *
0-
02
b11 6
#652870000000
1!
1%
1-
12
15
#652880000000
0!
0%
b100 *
0-
02
b100 6
#652890000000
1!
1%
1-
12
#652900000000
0!
0%
b101 *
0-
02
b101 6
#652910000000
1!
1%
1-
12
#652920000000
0!
0%
b110 *
0-
02
b110 6
#652930000000
1!
1%
1-
12
#652940000000
0!
0%
b111 *
0-
02
b111 6
#652950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#652960000000
0!
0%
b0 *
0-
02
b0 6
#652970000000
1!
1%
1-
12
#652980000000
0!
0%
b1 *
0-
02
b1 6
#652990000000
1!
1%
1-
12
#653000000000
0!
0%
b10 *
0-
02
b10 6
#653010000000
1!
1%
1-
12
#653020000000
0!
0%
b11 *
0-
02
b11 6
#653030000000
1!
1%
1-
12
15
#653040000000
0!
0%
b100 *
0-
02
b100 6
#653050000000
1!
1%
1-
12
#653060000000
0!
0%
b101 *
0-
02
b101 6
#653070000000
1!
1%
1-
12
#653080000000
0!
0%
b110 *
0-
02
b110 6
#653090000000
1!
1%
1-
12
#653100000000
0!
0%
b111 *
0-
02
b111 6
#653110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#653120000000
0!
0%
b0 *
0-
02
b0 6
#653130000000
1!
1%
1-
12
#653140000000
0!
0%
b1 *
0-
02
b1 6
#653150000000
1!
1%
1-
12
#653160000000
0!
0%
b10 *
0-
02
b10 6
#653170000000
1!
1%
1-
12
#653180000000
0!
0%
b11 *
0-
02
b11 6
#653190000000
1!
1%
1-
12
15
#653200000000
0!
0%
b100 *
0-
02
b100 6
#653210000000
1!
1%
1-
12
#653220000000
0!
0%
b101 *
0-
02
b101 6
#653230000000
1!
1%
1-
12
#653240000000
0!
0%
b110 *
0-
02
b110 6
#653250000000
1!
1%
1-
12
#653260000000
0!
0%
b111 *
0-
02
b111 6
#653270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#653280000000
0!
0%
b0 *
0-
02
b0 6
#653290000000
1!
1%
1-
12
#653300000000
0!
0%
b1 *
0-
02
b1 6
#653310000000
1!
1%
1-
12
#653320000000
0!
0%
b10 *
0-
02
b10 6
#653330000000
1!
1%
1-
12
#653340000000
0!
0%
b11 *
0-
02
b11 6
#653350000000
1!
1%
1-
12
15
#653360000000
0!
0%
b100 *
0-
02
b100 6
#653370000000
1!
1%
1-
12
#653380000000
0!
0%
b101 *
0-
02
b101 6
#653390000000
1!
1%
1-
12
#653400000000
0!
0%
b110 *
0-
02
b110 6
#653410000000
1!
1%
1-
12
#653420000000
0!
0%
b111 *
0-
02
b111 6
#653430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#653440000000
0!
0%
b0 *
0-
02
b0 6
#653450000000
1!
1%
1-
12
#653460000000
0!
0%
b1 *
0-
02
b1 6
#653470000000
1!
1%
1-
12
#653480000000
0!
0%
b10 *
0-
02
b10 6
#653490000000
1!
1%
1-
12
#653500000000
0!
0%
b11 *
0-
02
b11 6
#653510000000
1!
1%
1-
12
15
#653520000000
0!
0%
b100 *
0-
02
b100 6
#653530000000
1!
1%
1-
12
#653540000000
0!
0%
b101 *
0-
02
b101 6
#653550000000
1!
1%
1-
12
#653560000000
0!
0%
b110 *
0-
02
b110 6
#653570000000
1!
1%
1-
12
#653580000000
0!
0%
b111 *
0-
02
b111 6
#653590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#653600000000
0!
0%
b0 *
0-
02
b0 6
#653610000000
1!
1%
1-
12
#653620000000
0!
0%
b1 *
0-
02
b1 6
#653630000000
1!
1%
1-
12
#653640000000
0!
0%
b10 *
0-
02
b10 6
#653650000000
1!
1%
1-
12
#653660000000
0!
0%
b11 *
0-
02
b11 6
#653670000000
1!
1%
1-
12
15
#653680000000
0!
0%
b100 *
0-
02
b100 6
#653690000000
1!
1%
1-
12
#653700000000
0!
0%
b101 *
0-
02
b101 6
#653710000000
1!
1%
1-
12
#653720000000
0!
0%
b110 *
0-
02
b110 6
#653730000000
1!
1%
1-
12
#653740000000
0!
0%
b111 *
0-
02
b111 6
#653750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#653760000000
0!
0%
b0 *
0-
02
b0 6
#653770000000
1!
1%
1-
12
#653780000000
0!
0%
b1 *
0-
02
b1 6
#653790000000
1!
1%
1-
12
#653800000000
0!
0%
b10 *
0-
02
b10 6
#653810000000
1!
1%
1-
12
#653820000000
0!
0%
b11 *
0-
02
b11 6
#653830000000
1!
1%
1-
12
15
#653840000000
0!
0%
b100 *
0-
02
b100 6
#653850000000
1!
1%
1-
12
#653860000000
0!
0%
b101 *
0-
02
b101 6
#653870000000
1!
1%
1-
12
#653880000000
0!
0%
b110 *
0-
02
b110 6
#653890000000
1!
1%
1-
12
#653900000000
0!
0%
b111 *
0-
02
b111 6
#653910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#653920000000
0!
0%
b0 *
0-
02
b0 6
#653930000000
1!
1%
1-
12
#653940000000
0!
0%
b1 *
0-
02
b1 6
#653950000000
1!
1%
1-
12
#653960000000
0!
0%
b10 *
0-
02
b10 6
#653970000000
1!
1%
1-
12
#653980000000
0!
0%
b11 *
0-
02
b11 6
#653990000000
1!
1%
1-
12
15
#654000000000
0!
0%
b100 *
0-
02
b100 6
#654010000000
1!
1%
1-
12
#654020000000
0!
0%
b101 *
0-
02
b101 6
#654030000000
1!
1%
1-
12
#654040000000
0!
0%
b110 *
0-
02
b110 6
#654050000000
1!
1%
1-
12
#654060000000
0!
0%
b111 *
0-
02
b111 6
#654070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#654080000000
0!
0%
b0 *
0-
02
b0 6
#654090000000
1!
1%
1-
12
#654100000000
0!
0%
b1 *
0-
02
b1 6
#654110000000
1!
1%
1-
12
#654120000000
0!
0%
b10 *
0-
02
b10 6
#654130000000
1!
1%
1-
12
#654140000000
0!
0%
b11 *
0-
02
b11 6
#654150000000
1!
1%
1-
12
15
#654160000000
0!
0%
b100 *
0-
02
b100 6
#654170000000
1!
1%
1-
12
#654180000000
0!
0%
b101 *
0-
02
b101 6
#654190000000
1!
1%
1-
12
#654200000000
0!
0%
b110 *
0-
02
b110 6
#654210000000
1!
1%
1-
12
#654220000000
0!
0%
b111 *
0-
02
b111 6
#654230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#654240000000
0!
0%
b0 *
0-
02
b0 6
#654250000000
1!
1%
1-
12
#654260000000
0!
0%
b1 *
0-
02
b1 6
#654270000000
1!
1%
1-
12
#654280000000
0!
0%
b10 *
0-
02
b10 6
#654290000000
1!
1%
1-
12
#654300000000
0!
0%
b11 *
0-
02
b11 6
#654310000000
1!
1%
1-
12
15
#654320000000
0!
0%
b100 *
0-
02
b100 6
#654330000000
1!
1%
1-
12
#654340000000
0!
0%
b101 *
0-
02
b101 6
#654350000000
1!
1%
1-
12
#654360000000
0!
0%
b110 *
0-
02
b110 6
#654370000000
1!
1%
1-
12
#654380000000
0!
0%
b111 *
0-
02
b111 6
#654390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#654400000000
0!
0%
b0 *
0-
02
b0 6
#654410000000
1!
1%
1-
12
#654420000000
0!
0%
b1 *
0-
02
b1 6
#654430000000
1!
1%
1-
12
#654440000000
0!
0%
b10 *
0-
02
b10 6
#654450000000
1!
1%
1-
12
#654460000000
0!
0%
b11 *
0-
02
b11 6
#654470000000
1!
1%
1-
12
15
#654480000000
0!
0%
b100 *
0-
02
b100 6
#654490000000
1!
1%
1-
12
#654500000000
0!
0%
b101 *
0-
02
b101 6
#654510000000
1!
1%
1-
12
#654520000000
0!
0%
b110 *
0-
02
b110 6
#654530000000
1!
1%
1-
12
#654540000000
0!
0%
b111 *
0-
02
b111 6
#654550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#654560000000
0!
0%
b0 *
0-
02
b0 6
#654570000000
1!
1%
1-
12
#654580000000
0!
0%
b1 *
0-
02
b1 6
#654590000000
1!
1%
1-
12
#654600000000
0!
0%
b10 *
0-
02
b10 6
#654610000000
1!
1%
1-
12
#654620000000
0!
0%
b11 *
0-
02
b11 6
#654630000000
1!
1%
1-
12
15
#654640000000
0!
0%
b100 *
0-
02
b100 6
#654650000000
1!
1%
1-
12
#654660000000
0!
0%
b101 *
0-
02
b101 6
#654670000000
1!
1%
1-
12
#654680000000
0!
0%
b110 *
0-
02
b110 6
#654690000000
1!
1%
1-
12
#654700000000
0!
0%
b111 *
0-
02
b111 6
#654710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#654720000000
0!
0%
b0 *
0-
02
b0 6
#654730000000
1!
1%
1-
12
#654740000000
0!
0%
b1 *
0-
02
b1 6
#654750000000
1!
1%
1-
12
#654760000000
0!
0%
b10 *
0-
02
b10 6
#654770000000
1!
1%
1-
12
#654780000000
0!
0%
b11 *
0-
02
b11 6
#654790000000
1!
1%
1-
12
15
#654800000000
0!
0%
b100 *
0-
02
b100 6
#654810000000
1!
1%
1-
12
#654820000000
0!
0%
b101 *
0-
02
b101 6
#654830000000
1!
1%
1-
12
#654840000000
0!
0%
b110 *
0-
02
b110 6
#654850000000
1!
1%
1-
12
#654860000000
0!
0%
b111 *
0-
02
b111 6
#654870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#654880000000
0!
0%
b0 *
0-
02
b0 6
#654890000000
1!
1%
1-
12
#654900000000
0!
0%
b1 *
0-
02
b1 6
#654910000000
1!
1%
1-
12
#654920000000
0!
0%
b10 *
0-
02
b10 6
#654930000000
1!
1%
1-
12
#654940000000
0!
0%
b11 *
0-
02
b11 6
#654950000000
1!
1%
1-
12
15
#654960000000
0!
0%
b100 *
0-
02
b100 6
#654970000000
1!
1%
1-
12
#654980000000
0!
0%
b101 *
0-
02
b101 6
#654990000000
1!
1%
1-
12
#655000000000
0!
0%
b110 *
0-
02
b110 6
#655010000000
1!
1%
1-
12
#655020000000
0!
0%
b111 *
0-
02
b111 6
#655030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#655040000000
0!
0%
b0 *
0-
02
b0 6
#655050000000
1!
1%
1-
12
#655060000000
0!
0%
b1 *
0-
02
b1 6
#655070000000
1!
1%
1-
12
#655080000000
0!
0%
b10 *
0-
02
b10 6
#655090000000
1!
1%
1-
12
#655100000000
0!
0%
b11 *
0-
02
b11 6
#655110000000
1!
1%
1-
12
15
#655120000000
0!
0%
b100 *
0-
02
b100 6
#655130000000
1!
1%
1-
12
#655140000000
0!
0%
b101 *
0-
02
b101 6
#655150000000
1!
1%
1-
12
#655160000000
0!
0%
b110 *
0-
02
b110 6
#655170000000
1!
1%
1-
12
#655180000000
0!
0%
b111 *
0-
02
b111 6
#655190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#655200000000
0!
0%
b0 *
0-
02
b0 6
#655210000000
1!
1%
1-
12
#655220000000
0!
0%
b1 *
0-
02
b1 6
#655230000000
1!
1%
1-
12
#655240000000
0!
0%
b10 *
0-
02
b10 6
#655250000000
1!
1%
1-
12
#655260000000
0!
0%
b11 *
0-
02
b11 6
#655270000000
1!
1%
1-
12
15
#655280000000
0!
0%
b100 *
0-
02
b100 6
#655290000000
1!
1%
1-
12
#655300000000
0!
0%
b101 *
0-
02
b101 6
#655310000000
1!
1%
1-
12
#655320000000
0!
0%
b110 *
0-
02
b110 6
#655330000000
1!
1%
1-
12
#655340000000
0!
0%
b111 *
0-
02
b111 6
#655350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#655360000000
0!
0%
b0 *
0-
02
b0 6
#655370000000
1!
1%
1-
12
#655380000000
0!
0%
b1 *
0-
02
b1 6
#655390000000
1!
1%
1-
12
#655400000000
0!
0%
b10 *
0-
02
b10 6
#655410000000
1!
1%
1-
12
#655420000000
0!
0%
b11 *
0-
02
b11 6
#655430000000
1!
1%
1-
12
15
#655440000000
0!
0%
b100 *
0-
02
b100 6
#655450000000
1!
1%
1-
12
#655460000000
0!
0%
b101 *
0-
02
b101 6
#655470000000
1!
1%
1-
12
#655480000000
0!
0%
b110 *
0-
02
b110 6
#655490000000
1!
1%
1-
12
#655500000000
0!
0%
b111 *
0-
02
b111 6
#655510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#655520000000
0!
0%
b0 *
0-
02
b0 6
#655530000000
1!
1%
1-
12
#655540000000
0!
0%
b1 *
0-
02
b1 6
#655550000000
1!
1%
1-
12
#655560000000
0!
0%
b10 *
0-
02
b10 6
#655570000000
1!
1%
1-
12
#655580000000
0!
0%
b11 *
0-
02
b11 6
#655590000000
1!
1%
1-
12
15
#655600000000
0!
0%
b100 *
0-
02
b100 6
#655610000000
1!
1%
1-
12
#655620000000
0!
0%
b101 *
0-
02
b101 6
#655630000000
1!
1%
1-
12
#655640000000
0!
0%
b110 *
0-
02
b110 6
#655650000000
1!
1%
1-
12
#655660000000
0!
0%
b111 *
0-
02
b111 6
#655670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#655680000000
0!
0%
b0 *
0-
02
b0 6
#655690000000
1!
1%
1-
12
#655700000000
0!
0%
b1 *
0-
02
b1 6
#655710000000
1!
1%
1-
12
#655720000000
0!
0%
b10 *
0-
02
b10 6
#655730000000
1!
1%
1-
12
#655740000000
0!
0%
b11 *
0-
02
b11 6
#655750000000
1!
1%
1-
12
15
#655760000000
0!
0%
b100 *
0-
02
b100 6
#655770000000
1!
1%
1-
12
#655780000000
0!
0%
b101 *
0-
02
b101 6
#655790000000
1!
1%
1-
12
#655800000000
0!
0%
b110 *
0-
02
b110 6
#655810000000
1!
1%
1-
12
#655820000000
0!
0%
b111 *
0-
02
b111 6
#655830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#655840000000
0!
0%
b0 *
0-
02
b0 6
#655850000000
1!
1%
1-
12
#655860000000
0!
0%
b1 *
0-
02
b1 6
#655870000000
1!
1%
1-
12
#655880000000
0!
0%
b10 *
0-
02
b10 6
#655890000000
1!
1%
1-
12
#655900000000
0!
0%
b11 *
0-
02
b11 6
#655910000000
1!
1%
1-
12
15
#655920000000
0!
0%
b100 *
0-
02
b100 6
#655930000000
1!
1%
1-
12
#655940000000
0!
0%
b101 *
0-
02
b101 6
#655950000000
1!
1%
1-
12
#655960000000
0!
0%
b110 *
0-
02
b110 6
#655970000000
1!
1%
1-
12
#655980000000
0!
0%
b111 *
0-
02
b111 6
#655990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#656000000000
0!
0%
b0 *
0-
02
b0 6
#656010000000
1!
1%
1-
12
#656020000000
0!
0%
b1 *
0-
02
b1 6
#656030000000
1!
1%
1-
12
#656040000000
0!
0%
b10 *
0-
02
b10 6
#656050000000
1!
1%
1-
12
#656060000000
0!
0%
b11 *
0-
02
b11 6
#656070000000
1!
1%
1-
12
15
#656080000000
0!
0%
b100 *
0-
02
b100 6
#656090000000
1!
1%
1-
12
#656100000000
0!
0%
b101 *
0-
02
b101 6
#656110000000
1!
1%
1-
12
#656120000000
0!
0%
b110 *
0-
02
b110 6
#656130000000
1!
1%
1-
12
#656140000000
0!
0%
b111 *
0-
02
b111 6
#656150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#656160000000
0!
0%
b0 *
0-
02
b0 6
#656170000000
1!
1%
1-
12
#656180000000
0!
0%
b1 *
0-
02
b1 6
#656190000000
1!
1%
1-
12
#656200000000
0!
0%
b10 *
0-
02
b10 6
#656210000000
1!
1%
1-
12
#656220000000
0!
0%
b11 *
0-
02
b11 6
#656230000000
1!
1%
1-
12
15
#656240000000
0!
0%
b100 *
0-
02
b100 6
#656250000000
1!
1%
1-
12
#656260000000
0!
0%
b101 *
0-
02
b101 6
#656270000000
1!
1%
1-
12
#656280000000
0!
0%
b110 *
0-
02
b110 6
#656290000000
1!
1%
1-
12
#656300000000
0!
0%
b111 *
0-
02
b111 6
#656310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#656320000000
0!
0%
b0 *
0-
02
b0 6
#656330000000
1!
1%
1-
12
#656340000000
0!
0%
b1 *
0-
02
b1 6
#656350000000
1!
1%
1-
12
#656360000000
0!
0%
b10 *
0-
02
b10 6
#656370000000
1!
1%
1-
12
#656380000000
0!
0%
b11 *
0-
02
b11 6
#656390000000
1!
1%
1-
12
15
#656400000000
0!
0%
b100 *
0-
02
b100 6
#656410000000
1!
1%
1-
12
#656420000000
0!
0%
b101 *
0-
02
b101 6
#656430000000
1!
1%
1-
12
#656440000000
0!
0%
b110 *
0-
02
b110 6
#656450000000
1!
1%
1-
12
#656460000000
0!
0%
b111 *
0-
02
b111 6
#656470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#656480000000
0!
0%
b0 *
0-
02
b0 6
#656490000000
1!
1%
1-
12
#656500000000
0!
0%
b1 *
0-
02
b1 6
#656510000000
1!
1%
1-
12
#656520000000
0!
0%
b10 *
0-
02
b10 6
#656530000000
1!
1%
1-
12
#656540000000
0!
0%
b11 *
0-
02
b11 6
#656550000000
1!
1%
1-
12
15
#656560000000
0!
0%
b100 *
0-
02
b100 6
#656570000000
1!
1%
1-
12
#656580000000
0!
0%
b101 *
0-
02
b101 6
#656590000000
1!
1%
1-
12
#656600000000
0!
0%
b110 *
0-
02
b110 6
#656610000000
1!
1%
1-
12
#656620000000
0!
0%
b111 *
0-
02
b111 6
#656630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#656640000000
0!
0%
b0 *
0-
02
b0 6
#656650000000
1!
1%
1-
12
#656660000000
0!
0%
b1 *
0-
02
b1 6
#656670000000
1!
1%
1-
12
#656680000000
0!
0%
b10 *
0-
02
b10 6
#656690000000
1!
1%
1-
12
#656700000000
0!
0%
b11 *
0-
02
b11 6
#656710000000
1!
1%
1-
12
15
#656720000000
0!
0%
b100 *
0-
02
b100 6
#656730000000
1!
1%
1-
12
#656740000000
0!
0%
b101 *
0-
02
b101 6
#656750000000
1!
1%
1-
12
#656760000000
0!
0%
b110 *
0-
02
b110 6
#656770000000
1!
1%
1-
12
#656780000000
0!
0%
b111 *
0-
02
b111 6
#656790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#656800000000
0!
0%
b0 *
0-
02
b0 6
#656810000000
1!
1%
1-
12
#656820000000
0!
0%
b1 *
0-
02
b1 6
#656830000000
1!
1%
1-
12
#656840000000
0!
0%
b10 *
0-
02
b10 6
#656850000000
1!
1%
1-
12
#656860000000
0!
0%
b11 *
0-
02
b11 6
#656870000000
1!
1%
1-
12
15
#656880000000
0!
0%
b100 *
0-
02
b100 6
#656890000000
1!
1%
1-
12
#656900000000
0!
0%
b101 *
0-
02
b101 6
#656910000000
1!
1%
1-
12
#656920000000
0!
0%
b110 *
0-
02
b110 6
#656930000000
1!
1%
1-
12
#656940000000
0!
0%
b111 *
0-
02
b111 6
#656950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#656960000000
0!
0%
b0 *
0-
02
b0 6
#656970000000
1!
1%
1-
12
#656980000000
0!
0%
b1 *
0-
02
b1 6
#656990000000
1!
1%
1-
12
#657000000000
0!
0%
b10 *
0-
02
b10 6
#657010000000
1!
1%
1-
12
#657020000000
0!
0%
b11 *
0-
02
b11 6
#657030000000
1!
1%
1-
12
15
#657040000000
0!
0%
b100 *
0-
02
b100 6
#657050000000
1!
1%
1-
12
#657060000000
0!
0%
b101 *
0-
02
b101 6
#657070000000
1!
1%
1-
12
#657080000000
0!
0%
b110 *
0-
02
b110 6
#657090000000
1!
1%
1-
12
#657100000000
0!
0%
b111 *
0-
02
b111 6
#657110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#657120000000
0!
0%
b0 *
0-
02
b0 6
#657130000000
1!
1%
1-
12
#657140000000
0!
0%
b1 *
0-
02
b1 6
#657150000000
1!
1%
1-
12
#657160000000
0!
0%
b10 *
0-
02
b10 6
#657170000000
1!
1%
1-
12
#657180000000
0!
0%
b11 *
0-
02
b11 6
#657190000000
1!
1%
1-
12
15
#657200000000
0!
0%
b100 *
0-
02
b100 6
#657210000000
1!
1%
1-
12
#657220000000
0!
0%
b101 *
0-
02
b101 6
#657230000000
1!
1%
1-
12
#657240000000
0!
0%
b110 *
0-
02
b110 6
#657250000000
1!
1%
1-
12
#657260000000
0!
0%
b111 *
0-
02
b111 6
#657270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#657280000000
0!
0%
b0 *
0-
02
b0 6
#657290000000
1!
1%
1-
12
#657300000000
0!
0%
b1 *
0-
02
b1 6
#657310000000
1!
1%
1-
12
#657320000000
0!
0%
b10 *
0-
02
b10 6
#657330000000
1!
1%
1-
12
#657340000000
0!
0%
b11 *
0-
02
b11 6
#657350000000
1!
1%
1-
12
15
#657360000000
0!
0%
b100 *
0-
02
b100 6
#657370000000
1!
1%
1-
12
#657380000000
0!
0%
b101 *
0-
02
b101 6
#657390000000
1!
1%
1-
12
#657400000000
0!
0%
b110 *
0-
02
b110 6
#657410000000
1!
1%
1-
12
#657420000000
0!
0%
b111 *
0-
02
b111 6
#657430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#657440000000
0!
0%
b0 *
0-
02
b0 6
#657450000000
1!
1%
1-
12
#657460000000
0!
0%
b1 *
0-
02
b1 6
#657470000000
1!
1%
1-
12
#657480000000
0!
0%
b10 *
0-
02
b10 6
#657490000000
1!
1%
1-
12
#657500000000
0!
0%
b11 *
0-
02
b11 6
#657510000000
1!
1%
1-
12
15
#657520000000
0!
0%
b100 *
0-
02
b100 6
#657530000000
1!
1%
1-
12
#657540000000
0!
0%
b101 *
0-
02
b101 6
#657550000000
1!
1%
1-
12
#657560000000
0!
0%
b110 *
0-
02
b110 6
#657570000000
1!
1%
1-
12
#657580000000
0!
0%
b111 *
0-
02
b111 6
#657590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#657600000000
0!
0%
b0 *
0-
02
b0 6
#657610000000
1!
1%
1-
12
#657620000000
0!
0%
b1 *
0-
02
b1 6
#657630000000
1!
1%
1-
12
#657640000000
0!
0%
b10 *
0-
02
b10 6
#657650000000
1!
1%
1-
12
#657660000000
0!
0%
b11 *
0-
02
b11 6
#657670000000
1!
1%
1-
12
15
#657680000000
0!
0%
b100 *
0-
02
b100 6
#657690000000
1!
1%
1-
12
#657700000000
0!
0%
b101 *
0-
02
b101 6
#657710000000
1!
1%
1-
12
#657720000000
0!
0%
b110 *
0-
02
b110 6
#657730000000
1!
1%
1-
12
#657740000000
0!
0%
b111 *
0-
02
b111 6
#657750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#657760000000
0!
0%
b0 *
0-
02
b0 6
#657770000000
1!
1%
1-
12
#657780000000
0!
0%
b1 *
0-
02
b1 6
#657790000000
1!
1%
1-
12
#657800000000
0!
0%
b10 *
0-
02
b10 6
#657810000000
1!
1%
1-
12
#657820000000
0!
0%
b11 *
0-
02
b11 6
#657830000000
1!
1%
1-
12
15
#657840000000
0!
0%
b100 *
0-
02
b100 6
#657850000000
1!
1%
1-
12
#657860000000
0!
0%
b101 *
0-
02
b101 6
#657870000000
1!
1%
1-
12
#657880000000
0!
0%
b110 *
0-
02
b110 6
#657890000000
1!
1%
1-
12
#657900000000
0!
0%
b111 *
0-
02
b111 6
#657910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#657920000000
0!
0%
b0 *
0-
02
b0 6
#657930000000
1!
1%
1-
12
#657940000000
0!
0%
b1 *
0-
02
b1 6
#657950000000
1!
1%
1-
12
#657960000000
0!
0%
b10 *
0-
02
b10 6
#657970000000
1!
1%
1-
12
#657980000000
0!
0%
b11 *
0-
02
b11 6
#657990000000
1!
1%
1-
12
15
#658000000000
0!
0%
b100 *
0-
02
b100 6
#658010000000
1!
1%
1-
12
#658020000000
0!
0%
b101 *
0-
02
b101 6
#658030000000
1!
1%
1-
12
#658040000000
0!
0%
b110 *
0-
02
b110 6
#658050000000
1!
1%
1-
12
#658060000000
0!
0%
b111 *
0-
02
b111 6
#658070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#658080000000
0!
0%
b0 *
0-
02
b0 6
#658090000000
1!
1%
1-
12
#658100000000
0!
0%
b1 *
0-
02
b1 6
#658110000000
1!
1%
1-
12
#658120000000
0!
0%
b10 *
0-
02
b10 6
#658130000000
1!
1%
1-
12
#658140000000
0!
0%
b11 *
0-
02
b11 6
#658150000000
1!
1%
1-
12
15
#658160000000
0!
0%
b100 *
0-
02
b100 6
#658170000000
1!
1%
1-
12
#658180000000
0!
0%
b101 *
0-
02
b101 6
#658190000000
1!
1%
1-
12
#658200000000
0!
0%
b110 *
0-
02
b110 6
#658210000000
1!
1%
1-
12
#658220000000
0!
0%
b111 *
0-
02
b111 6
#658230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#658240000000
0!
0%
b0 *
0-
02
b0 6
#658250000000
1!
1%
1-
12
#658260000000
0!
0%
b1 *
0-
02
b1 6
#658270000000
1!
1%
1-
12
#658280000000
0!
0%
b10 *
0-
02
b10 6
#658290000000
1!
1%
1-
12
#658300000000
0!
0%
b11 *
0-
02
b11 6
#658310000000
1!
1%
1-
12
15
#658320000000
0!
0%
b100 *
0-
02
b100 6
#658330000000
1!
1%
1-
12
#658340000000
0!
0%
b101 *
0-
02
b101 6
#658350000000
1!
1%
1-
12
#658360000000
0!
0%
b110 *
0-
02
b110 6
#658370000000
1!
1%
1-
12
#658380000000
0!
0%
b111 *
0-
02
b111 6
#658390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#658400000000
0!
0%
b0 *
0-
02
b0 6
#658410000000
1!
1%
1-
12
#658420000000
0!
0%
b1 *
0-
02
b1 6
#658430000000
1!
1%
1-
12
#658440000000
0!
0%
b10 *
0-
02
b10 6
#658450000000
1!
1%
1-
12
#658460000000
0!
0%
b11 *
0-
02
b11 6
#658470000000
1!
1%
1-
12
15
#658480000000
0!
0%
b100 *
0-
02
b100 6
#658490000000
1!
1%
1-
12
#658500000000
0!
0%
b101 *
0-
02
b101 6
#658510000000
1!
1%
1-
12
#658520000000
0!
0%
b110 *
0-
02
b110 6
#658530000000
1!
1%
1-
12
#658540000000
0!
0%
b111 *
0-
02
b111 6
#658550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#658560000000
0!
0%
b0 *
0-
02
b0 6
#658570000000
1!
1%
1-
12
#658580000000
0!
0%
b1 *
0-
02
b1 6
#658590000000
1!
1%
1-
12
#658600000000
0!
0%
b10 *
0-
02
b10 6
#658610000000
1!
1%
1-
12
#658620000000
0!
0%
b11 *
0-
02
b11 6
#658630000000
1!
1%
1-
12
15
#658640000000
0!
0%
b100 *
0-
02
b100 6
#658650000000
1!
1%
1-
12
#658660000000
0!
0%
b101 *
0-
02
b101 6
#658670000000
1!
1%
1-
12
#658680000000
0!
0%
b110 *
0-
02
b110 6
#658690000000
1!
1%
1-
12
#658700000000
0!
0%
b111 *
0-
02
b111 6
#658710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#658720000000
0!
0%
b0 *
0-
02
b0 6
#658730000000
1!
1%
1-
12
#658740000000
0!
0%
b1 *
0-
02
b1 6
#658750000000
1!
1%
1-
12
#658760000000
0!
0%
b10 *
0-
02
b10 6
#658770000000
1!
1%
1-
12
#658780000000
0!
0%
b11 *
0-
02
b11 6
#658790000000
1!
1%
1-
12
15
#658800000000
0!
0%
b100 *
0-
02
b100 6
#658810000000
1!
1%
1-
12
#658820000000
0!
0%
b101 *
0-
02
b101 6
#658830000000
1!
1%
1-
12
#658840000000
0!
0%
b110 *
0-
02
b110 6
#658850000000
1!
1%
1-
12
#658860000000
0!
0%
b111 *
0-
02
b111 6
#658870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#658880000000
0!
0%
b0 *
0-
02
b0 6
#658890000000
1!
1%
1-
12
#658900000000
0!
0%
b1 *
0-
02
b1 6
#658910000000
1!
1%
1-
12
#658920000000
0!
0%
b10 *
0-
02
b10 6
#658930000000
1!
1%
1-
12
#658940000000
0!
0%
b11 *
0-
02
b11 6
#658950000000
1!
1%
1-
12
15
#658960000000
0!
0%
b100 *
0-
02
b100 6
#658970000000
1!
1%
1-
12
#658980000000
0!
0%
b101 *
0-
02
b101 6
#658990000000
1!
1%
1-
12
#659000000000
0!
0%
b110 *
0-
02
b110 6
#659010000000
1!
1%
1-
12
#659020000000
0!
0%
b111 *
0-
02
b111 6
#659030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#659040000000
0!
0%
b0 *
0-
02
b0 6
#659050000000
1!
1%
1-
12
#659060000000
0!
0%
b1 *
0-
02
b1 6
#659070000000
1!
1%
1-
12
#659080000000
0!
0%
b10 *
0-
02
b10 6
#659090000000
1!
1%
1-
12
#659100000000
0!
0%
b11 *
0-
02
b11 6
#659110000000
1!
1%
1-
12
15
#659120000000
0!
0%
b100 *
0-
02
b100 6
#659130000000
1!
1%
1-
12
#659140000000
0!
0%
b101 *
0-
02
b101 6
#659150000000
1!
1%
1-
12
#659160000000
0!
0%
b110 *
0-
02
b110 6
#659170000000
1!
1%
1-
12
#659180000000
0!
0%
b111 *
0-
02
b111 6
#659190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#659200000000
0!
0%
b0 *
0-
02
b0 6
#659210000000
1!
1%
1-
12
#659220000000
0!
0%
b1 *
0-
02
b1 6
#659230000000
1!
1%
1-
12
#659240000000
0!
0%
b10 *
0-
02
b10 6
#659250000000
1!
1%
1-
12
#659260000000
0!
0%
b11 *
0-
02
b11 6
#659270000000
1!
1%
1-
12
15
#659280000000
0!
0%
b100 *
0-
02
b100 6
#659290000000
1!
1%
1-
12
#659300000000
0!
0%
b101 *
0-
02
b101 6
#659310000000
1!
1%
1-
12
#659320000000
0!
0%
b110 *
0-
02
b110 6
#659330000000
1!
1%
1-
12
#659340000000
0!
0%
b111 *
0-
02
b111 6
#659350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#659360000000
0!
0%
b0 *
0-
02
b0 6
#659370000000
1!
1%
1-
12
#659380000000
0!
0%
b1 *
0-
02
b1 6
#659390000000
1!
1%
1-
12
#659400000000
0!
0%
b10 *
0-
02
b10 6
#659410000000
1!
1%
1-
12
#659420000000
0!
0%
b11 *
0-
02
b11 6
#659430000000
1!
1%
1-
12
15
#659440000000
0!
0%
b100 *
0-
02
b100 6
#659450000000
1!
1%
1-
12
#659460000000
0!
0%
b101 *
0-
02
b101 6
#659470000000
1!
1%
1-
12
#659480000000
0!
0%
b110 *
0-
02
b110 6
#659490000000
1!
1%
1-
12
#659500000000
0!
0%
b111 *
0-
02
b111 6
#659510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#659520000000
0!
0%
b0 *
0-
02
b0 6
#659530000000
1!
1%
1-
12
#659540000000
0!
0%
b1 *
0-
02
b1 6
#659550000000
1!
1%
1-
12
#659560000000
0!
0%
b10 *
0-
02
b10 6
#659570000000
1!
1%
1-
12
#659580000000
0!
0%
b11 *
0-
02
b11 6
#659590000000
1!
1%
1-
12
15
#659600000000
0!
0%
b100 *
0-
02
b100 6
#659610000000
1!
1%
1-
12
#659620000000
0!
0%
b101 *
0-
02
b101 6
#659630000000
1!
1%
1-
12
#659640000000
0!
0%
b110 *
0-
02
b110 6
#659650000000
1!
1%
1-
12
#659660000000
0!
0%
b111 *
0-
02
b111 6
#659670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#659680000000
0!
0%
b0 *
0-
02
b0 6
#659690000000
1!
1%
1-
12
#659700000000
0!
0%
b1 *
0-
02
b1 6
#659710000000
1!
1%
1-
12
#659720000000
0!
0%
b10 *
0-
02
b10 6
#659730000000
1!
1%
1-
12
#659740000000
0!
0%
b11 *
0-
02
b11 6
#659750000000
1!
1%
1-
12
15
#659760000000
0!
0%
b100 *
0-
02
b100 6
#659770000000
1!
1%
1-
12
#659780000000
0!
0%
b101 *
0-
02
b101 6
#659790000000
1!
1%
1-
12
#659800000000
0!
0%
b110 *
0-
02
b110 6
#659810000000
1!
1%
1-
12
#659820000000
0!
0%
b111 *
0-
02
b111 6
#659830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#659840000000
0!
0%
b0 *
0-
02
b0 6
#659850000000
1!
1%
1-
12
#659860000000
0!
0%
b1 *
0-
02
b1 6
#659870000000
1!
1%
1-
12
#659880000000
0!
0%
b10 *
0-
02
b10 6
#659890000000
1!
1%
1-
12
#659900000000
0!
0%
b11 *
0-
02
b11 6
#659910000000
1!
1%
1-
12
15
#659920000000
0!
0%
b100 *
0-
02
b100 6
#659930000000
1!
1%
1-
12
#659940000000
0!
0%
b101 *
0-
02
b101 6
#659950000000
1!
1%
1-
12
#659960000000
0!
0%
b110 *
0-
02
b110 6
#659970000000
1!
1%
1-
12
#659980000000
0!
0%
b111 *
0-
02
b111 6
#659990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#660000000000
0!
0%
b0 *
0-
02
b0 6
#660010000000
1!
1%
1-
12
#660020000000
0!
0%
b1 *
0-
02
b1 6
#660030000000
1!
1%
1-
12
#660040000000
0!
0%
b10 *
0-
02
b10 6
#660050000000
1!
1%
1-
12
#660060000000
0!
0%
b11 *
0-
02
b11 6
#660070000000
1!
1%
1-
12
15
#660080000000
0!
0%
b100 *
0-
02
b100 6
#660090000000
1!
1%
1-
12
#660100000000
0!
0%
b101 *
0-
02
b101 6
#660110000000
1!
1%
1-
12
#660120000000
0!
0%
b110 *
0-
02
b110 6
#660130000000
1!
1%
1-
12
#660140000000
0!
0%
b111 *
0-
02
b111 6
#660150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#660160000000
0!
0%
b0 *
0-
02
b0 6
#660170000000
1!
1%
1-
12
#660180000000
0!
0%
b1 *
0-
02
b1 6
#660190000000
1!
1%
1-
12
#660200000000
0!
0%
b10 *
0-
02
b10 6
#660210000000
1!
1%
1-
12
#660220000000
0!
0%
b11 *
0-
02
b11 6
#660230000000
1!
1%
1-
12
15
#660240000000
0!
0%
b100 *
0-
02
b100 6
#660250000000
1!
1%
1-
12
#660260000000
0!
0%
b101 *
0-
02
b101 6
#660270000000
1!
1%
1-
12
#660280000000
0!
0%
b110 *
0-
02
b110 6
#660290000000
1!
1%
1-
12
#660300000000
0!
0%
b111 *
0-
02
b111 6
#660310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#660320000000
0!
0%
b0 *
0-
02
b0 6
#660330000000
1!
1%
1-
12
#660340000000
0!
0%
b1 *
0-
02
b1 6
#660350000000
1!
1%
1-
12
#660360000000
0!
0%
b10 *
0-
02
b10 6
#660370000000
1!
1%
1-
12
#660380000000
0!
0%
b11 *
0-
02
b11 6
#660390000000
1!
1%
1-
12
15
#660400000000
0!
0%
b100 *
0-
02
b100 6
#660410000000
1!
1%
1-
12
#660420000000
0!
0%
b101 *
0-
02
b101 6
#660430000000
1!
1%
1-
12
#660440000000
0!
0%
b110 *
0-
02
b110 6
#660450000000
1!
1%
1-
12
#660460000000
0!
0%
b111 *
0-
02
b111 6
#660470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#660480000000
0!
0%
b0 *
0-
02
b0 6
#660490000000
1!
1%
1-
12
#660500000000
0!
0%
b1 *
0-
02
b1 6
#660510000000
1!
1%
1-
12
#660520000000
0!
0%
b10 *
0-
02
b10 6
#660530000000
1!
1%
1-
12
#660540000000
0!
0%
b11 *
0-
02
b11 6
#660550000000
1!
1%
1-
12
15
#660560000000
0!
0%
b100 *
0-
02
b100 6
#660570000000
1!
1%
1-
12
#660580000000
0!
0%
b101 *
0-
02
b101 6
#660590000000
1!
1%
1-
12
#660600000000
0!
0%
b110 *
0-
02
b110 6
#660610000000
1!
1%
1-
12
#660620000000
0!
0%
b111 *
0-
02
b111 6
#660630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#660640000000
0!
0%
b0 *
0-
02
b0 6
#660650000000
1!
1%
1-
12
#660660000000
0!
0%
b1 *
0-
02
b1 6
#660670000000
1!
1%
1-
12
#660680000000
0!
0%
b10 *
0-
02
b10 6
#660690000000
1!
1%
1-
12
#660700000000
0!
0%
b11 *
0-
02
b11 6
#660710000000
1!
1%
1-
12
15
#660720000000
0!
0%
b100 *
0-
02
b100 6
#660730000000
1!
1%
1-
12
#660740000000
0!
0%
b101 *
0-
02
b101 6
#660750000000
1!
1%
1-
12
#660760000000
0!
0%
b110 *
0-
02
b110 6
#660770000000
1!
1%
1-
12
#660780000000
0!
0%
b111 *
0-
02
b111 6
#660790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#660800000000
0!
0%
b0 *
0-
02
b0 6
#660810000000
1!
1%
1-
12
#660820000000
0!
0%
b1 *
0-
02
b1 6
#660830000000
1!
1%
1-
12
#660840000000
0!
0%
b10 *
0-
02
b10 6
#660850000000
1!
1%
1-
12
#660860000000
0!
0%
b11 *
0-
02
b11 6
#660870000000
1!
1%
1-
12
15
#660880000000
0!
0%
b100 *
0-
02
b100 6
#660890000000
1!
1%
1-
12
#660900000000
0!
0%
b101 *
0-
02
b101 6
#660910000000
1!
1%
1-
12
#660920000000
0!
0%
b110 *
0-
02
b110 6
#660930000000
1!
1%
1-
12
#660940000000
0!
0%
b111 *
0-
02
b111 6
#660950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#660960000000
0!
0%
b0 *
0-
02
b0 6
#660970000000
1!
1%
1-
12
#660980000000
0!
0%
b1 *
0-
02
b1 6
#660990000000
1!
1%
1-
12
#661000000000
0!
0%
b10 *
0-
02
b10 6
#661010000000
1!
1%
1-
12
#661020000000
0!
0%
b11 *
0-
02
b11 6
#661030000000
1!
1%
1-
12
15
#661040000000
0!
0%
b100 *
0-
02
b100 6
#661050000000
1!
1%
1-
12
#661060000000
0!
0%
b101 *
0-
02
b101 6
#661070000000
1!
1%
1-
12
#661080000000
0!
0%
b110 *
0-
02
b110 6
#661090000000
1!
1%
1-
12
#661100000000
0!
0%
b111 *
0-
02
b111 6
#661110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#661120000000
0!
0%
b0 *
0-
02
b0 6
#661130000000
1!
1%
1-
12
#661140000000
0!
0%
b1 *
0-
02
b1 6
#661150000000
1!
1%
1-
12
#661160000000
0!
0%
b10 *
0-
02
b10 6
#661170000000
1!
1%
1-
12
#661180000000
0!
0%
b11 *
0-
02
b11 6
#661190000000
1!
1%
1-
12
15
#661200000000
0!
0%
b100 *
0-
02
b100 6
#661210000000
1!
1%
1-
12
#661220000000
0!
0%
b101 *
0-
02
b101 6
#661230000000
1!
1%
1-
12
#661240000000
0!
0%
b110 *
0-
02
b110 6
#661250000000
1!
1%
1-
12
#661260000000
0!
0%
b111 *
0-
02
b111 6
#661270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#661280000000
0!
0%
b0 *
0-
02
b0 6
#661290000000
1!
1%
1-
12
#661300000000
0!
0%
b1 *
0-
02
b1 6
#661310000000
1!
1%
1-
12
#661320000000
0!
0%
b10 *
0-
02
b10 6
#661330000000
1!
1%
1-
12
#661340000000
0!
0%
b11 *
0-
02
b11 6
#661350000000
1!
1%
1-
12
15
#661360000000
0!
0%
b100 *
0-
02
b100 6
#661370000000
1!
1%
1-
12
#661380000000
0!
0%
b101 *
0-
02
b101 6
#661390000000
1!
1%
1-
12
#661400000000
0!
0%
b110 *
0-
02
b110 6
#661410000000
1!
1%
1-
12
#661420000000
0!
0%
b111 *
0-
02
b111 6
#661430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#661440000000
0!
0%
b0 *
0-
02
b0 6
#661450000000
1!
1%
1-
12
#661460000000
0!
0%
b1 *
0-
02
b1 6
#661470000000
1!
1%
1-
12
#661480000000
0!
0%
b10 *
0-
02
b10 6
#661490000000
1!
1%
1-
12
#661500000000
0!
0%
b11 *
0-
02
b11 6
#661510000000
1!
1%
1-
12
15
#661520000000
0!
0%
b100 *
0-
02
b100 6
#661530000000
1!
1%
1-
12
#661540000000
0!
0%
b101 *
0-
02
b101 6
#661550000000
1!
1%
1-
12
#661560000000
0!
0%
b110 *
0-
02
b110 6
#661570000000
1!
1%
1-
12
#661580000000
0!
0%
b111 *
0-
02
b111 6
#661590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#661600000000
0!
0%
b0 *
0-
02
b0 6
#661610000000
1!
1%
1-
12
#661620000000
0!
0%
b1 *
0-
02
b1 6
#661630000000
1!
1%
1-
12
#661640000000
0!
0%
b10 *
0-
02
b10 6
#661650000000
1!
1%
1-
12
#661660000000
0!
0%
b11 *
0-
02
b11 6
#661670000000
1!
1%
1-
12
15
#661680000000
0!
0%
b100 *
0-
02
b100 6
#661690000000
1!
1%
1-
12
#661700000000
0!
0%
b101 *
0-
02
b101 6
#661710000000
1!
1%
1-
12
#661720000000
0!
0%
b110 *
0-
02
b110 6
#661730000000
1!
1%
1-
12
#661740000000
0!
0%
b111 *
0-
02
b111 6
#661750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#661760000000
0!
0%
b0 *
0-
02
b0 6
#661770000000
1!
1%
1-
12
#661780000000
0!
0%
b1 *
0-
02
b1 6
#661790000000
1!
1%
1-
12
#661800000000
0!
0%
b10 *
0-
02
b10 6
#661810000000
1!
1%
1-
12
#661820000000
0!
0%
b11 *
0-
02
b11 6
#661830000000
1!
1%
1-
12
15
#661840000000
0!
0%
b100 *
0-
02
b100 6
#661850000000
1!
1%
1-
12
#661860000000
0!
0%
b101 *
0-
02
b101 6
#661870000000
1!
1%
1-
12
#661880000000
0!
0%
b110 *
0-
02
b110 6
#661890000000
1!
1%
1-
12
#661900000000
0!
0%
b111 *
0-
02
b111 6
#661910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#661920000000
0!
0%
b0 *
0-
02
b0 6
#661930000000
1!
1%
1-
12
#661940000000
0!
0%
b1 *
0-
02
b1 6
#661950000000
1!
1%
1-
12
#661960000000
0!
0%
b10 *
0-
02
b10 6
#661970000000
1!
1%
1-
12
#661980000000
0!
0%
b11 *
0-
02
b11 6
#661990000000
1!
1%
1-
12
15
#662000000000
0!
0%
b100 *
0-
02
b100 6
#662010000000
1!
1%
1-
12
#662020000000
0!
0%
b101 *
0-
02
b101 6
#662030000000
1!
1%
1-
12
#662040000000
0!
0%
b110 *
0-
02
b110 6
#662050000000
1!
1%
1-
12
#662060000000
0!
0%
b111 *
0-
02
b111 6
#662070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#662080000000
0!
0%
b0 *
0-
02
b0 6
#662090000000
1!
1%
1-
12
#662100000000
0!
0%
b1 *
0-
02
b1 6
#662110000000
1!
1%
1-
12
#662120000000
0!
0%
b10 *
0-
02
b10 6
#662130000000
1!
1%
1-
12
#662140000000
0!
0%
b11 *
0-
02
b11 6
#662150000000
1!
1%
1-
12
15
#662160000000
0!
0%
b100 *
0-
02
b100 6
#662170000000
1!
1%
1-
12
#662180000000
0!
0%
b101 *
0-
02
b101 6
#662190000000
1!
1%
1-
12
#662200000000
0!
0%
b110 *
0-
02
b110 6
#662210000000
1!
1%
1-
12
#662220000000
0!
0%
b111 *
0-
02
b111 6
#662230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#662240000000
0!
0%
b0 *
0-
02
b0 6
#662250000000
1!
1%
1-
12
#662260000000
0!
0%
b1 *
0-
02
b1 6
#662270000000
1!
1%
1-
12
#662280000000
0!
0%
b10 *
0-
02
b10 6
#662290000000
1!
1%
1-
12
#662300000000
0!
0%
b11 *
0-
02
b11 6
#662310000000
1!
1%
1-
12
15
#662320000000
0!
0%
b100 *
0-
02
b100 6
#662330000000
1!
1%
1-
12
#662340000000
0!
0%
b101 *
0-
02
b101 6
#662350000000
1!
1%
1-
12
#662360000000
0!
0%
b110 *
0-
02
b110 6
#662370000000
1!
1%
1-
12
#662380000000
0!
0%
b111 *
0-
02
b111 6
#662390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#662400000000
0!
0%
b0 *
0-
02
b0 6
#662410000000
1!
1%
1-
12
#662420000000
0!
0%
b1 *
0-
02
b1 6
#662430000000
1!
1%
1-
12
#662440000000
0!
0%
b10 *
0-
02
b10 6
#662450000000
1!
1%
1-
12
#662460000000
0!
0%
b11 *
0-
02
b11 6
#662470000000
1!
1%
1-
12
15
#662480000000
0!
0%
b100 *
0-
02
b100 6
#662490000000
1!
1%
1-
12
#662500000000
0!
0%
b101 *
0-
02
b101 6
#662510000000
1!
1%
1-
12
#662520000000
0!
0%
b110 *
0-
02
b110 6
#662530000000
1!
1%
1-
12
#662540000000
0!
0%
b111 *
0-
02
b111 6
#662550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#662560000000
0!
0%
b0 *
0-
02
b0 6
#662570000000
1!
1%
1-
12
#662580000000
0!
0%
b1 *
0-
02
b1 6
#662590000000
1!
1%
1-
12
#662600000000
0!
0%
b10 *
0-
02
b10 6
#662610000000
1!
1%
1-
12
#662620000000
0!
0%
b11 *
0-
02
b11 6
#662630000000
1!
1%
1-
12
15
#662640000000
0!
0%
b100 *
0-
02
b100 6
#662650000000
1!
1%
1-
12
#662660000000
0!
0%
b101 *
0-
02
b101 6
#662670000000
1!
1%
1-
12
#662680000000
0!
0%
b110 *
0-
02
b110 6
#662690000000
1!
1%
1-
12
#662700000000
0!
0%
b111 *
0-
02
b111 6
#662710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#662720000000
0!
0%
b0 *
0-
02
b0 6
#662730000000
1!
1%
1-
12
#662740000000
0!
0%
b1 *
0-
02
b1 6
#662750000000
1!
1%
1-
12
#662760000000
0!
0%
b10 *
0-
02
b10 6
#662770000000
1!
1%
1-
12
#662780000000
0!
0%
b11 *
0-
02
b11 6
#662790000000
1!
1%
1-
12
15
#662800000000
0!
0%
b100 *
0-
02
b100 6
#662810000000
1!
1%
1-
12
#662820000000
0!
0%
b101 *
0-
02
b101 6
#662830000000
1!
1%
1-
12
#662840000000
0!
0%
b110 *
0-
02
b110 6
#662850000000
1!
1%
1-
12
#662860000000
0!
0%
b111 *
0-
02
b111 6
#662870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#662880000000
0!
0%
b0 *
0-
02
b0 6
#662890000000
1!
1%
1-
12
#662900000000
0!
0%
b1 *
0-
02
b1 6
#662910000000
1!
1%
1-
12
#662920000000
0!
0%
b10 *
0-
02
b10 6
#662930000000
1!
1%
1-
12
#662940000000
0!
0%
b11 *
0-
02
b11 6
#662950000000
1!
1%
1-
12
15
#662960000000
0!
0%
b100 *
0-
02
b100 6
#662970000000
1!
1%
1-
12
#662980000000
0!
0%
b101 *
0-
02
b101 6
#662990000000
1!
1%
1-
12
#663000000000
0!
0%
b110 *
0-
02
b110 6
#663010000000
1!
1%
1-
12
#663020000000
0!
0%
b111 *
0-
02
b111 6
#663030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#663040000000
0!
0%
b0 *
0-
02
b0 6
#663050000000
1!
1%
1-
12
#663060000000
0!
0%
b1 *
0-
02
b1 6
#663070000000
1!
1%
1-
12
#663080000000
0!
0%
b10 *
0-
02
b10 6
#663090000000
1!
1%
1-
12
#663100000000
0!
0%
b11 *
0-
02
b11 6
#663110000000
1!
1%
1-
12
15
#663120000000
0!
0%
b100 *
0-
02
b100 6
#663130000000
1!
1%
1-
12
#663140000000
0!
0%
b101 *
0-
02
b101 6
#663150000000
1!
1%
1-
12
#663160000000
0!
0%
b110 *
0-
02
b110 6
#663170000000
1!
1%
1-
12
#663180000000
0!
0%
b111 *
0-
02
b111 6
#663190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#663200000000
0!
0%
b0 *
0-
02
b0 6
#663210000000
1!
1%
1-
12
#663220000000
0!
0%
b1 *
0-
02
b1 6
#663230000000
1!
1%
1-
12
#663240000000
0!
0%
b10 *
0-
02
b10 6
#663250000000
1!
1%
1-
12
#663260000000
0!
0%
b11 *
0-
02
b11 6
#663270000000
1!
1%
1-
12
15
#663280000000
0!
0%
b100 *
0-
02
b100 6
#663290000000
1!
1%
1-
12
#663300000000
0!
0%
b101 *
0-
02
b101 6
#663310000000
1!
1%
1-
12
#663320000000
0!
0%
b110 *
0-
02
b110 6
#663330000000
1!
1%
1-
12
#663340000000
0!
0%
b111 *
0-
02
b111 6
#663350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#663360000000
0!
0%
b0 *
0-
02
b0 6
#663370000000
1!
1%
1-
12
#663380000000
0!
0%
b1 *
0-
02
b1 6
#663390000000
1!
1%
1-
12
#663400000000
0!
0%
b10 *
0-
02
b10 6
#663410000000
1!
1%
1-
12
#663420000000
0!
0%
b11 *
0-
02
b11 6
#663430000000
1!
1%
1-
12
15
#663440000000
0!
0%
b100 *
0-
02
b100 6
#663450000000
1!
1%
1-
12
#663460000000
0!
0%
b101 *
0-
02
b101 6
#663470000000
1!
1%
1-
12
#663480000000
0!
0%
b110 *
0-
02
b110 6
#663490000000
1!
1%
1-
12
#663500000000
0!
0%
b111 *
0-
02
b111 6
#663510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#663520000000
0!
0%
b0 *
0-
02
b0 6
#663530000000
1!
1%
1-
12
#663540000000
0!
0%
b1 *
0-
02
b1 6
#663550000000
1!
1%
1-
12
#663560000000
0!
0%
b10 *
0-
02
b10 6
#663570000000
1!
1%
1-
12
#663580000000
0!
0%
b11 *
0-
02
b11 6
#663590000000
1!
1%
1-
12
15
#663600000000
0!
0%
b100 *
0-
02
b100 6
#663610000000
1!
1%
1-
12
#663620000000
0!
0%
b101 *
0-
02
b101 6
#663630000000
1!
1%
1-
12
#663640000000
0!
0%
b110 *
0-
02
b110 6
#663650000000
1!
1%
1-
12
#663660000000
0!
0%
b111 *
0-
02
b111 6
#663670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#663680000000
0!
0%
b0 *
0-
02
b0 6
#663690000000
1!
1%
1-
12
#663700000000
0!
0%
b1 *
0-
02
b1 6
#663710000000
1!
1%
1-
12
#663720000000
0!
0%
b10 *
0-
02
b10 6
#663730000000
1!
1%
1-
12
#663740000000
0!
0%
b11 *
0-
02
b11 6
#663750000000
1!
1%
1-
12
15
#663760000000
0!
0%
b100 *
0-
02
b100 6
#663770000000
1!
1%
1-
12
#663780000000
0!
0%
b101 *
0-
02
b101 6
#663790000000
1!
1%
1-
12
#663800000000
0!
0%
b110 *
0-
02
b110 6
#663810000000
1!
1%
1-
12
#663820000000
0!
0%
b111 *
0-
02
b111 6
#663830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#663840000000
0!
0%
b0 *
0-
02
b0 6
#663850000000
1!
1%
1-
12
#663860000000
0!
0%
b1 *
0-
02
b1 6
#663870000000
1!
1%
1-
12
#663880000000
0!
0%
b10 *
0-
02
b10 6
#663890000000
1!
1%
1-
12
#663900000000
0!
0%
b11 *
0-
02
b11 6
#663910000000
1!
1%
1-
12
15
#663920000000
0!
0%
b100 *
0-
02
b100 6
#663930000000
1!
1%
1-
12
#663940000000
0!
0%
b101 *
0-
02
b101 6
#663950000000
1!
1%
1-
12
#663960000000
0!
0%
b110 *
0-
02
b110 6
#663970000000
1!
1%
1-
12
#663980000000
0!
0%
b111 *
0-
02
b111 6
#663990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#664000000000
0!
0%
b0 *
0-
02
b0 6
#664010000000
1!
1%
1-
12
#664020000000
0!
0%
b1 *
0-
02
b1 6
#664030000000
1!
1%
1-
12
#664040000000
0!
0%
b10 *
0-
02
b10 6
#664050000000
1!
1%
1-
12
#664060000000
0!
0%
b11 *
0-
02
b11 6
#664070000000
1!
1%
1-
12
15
#664080000000
0!
0%
b100 *
0-
02
b100 6
#664090000000
1!
1%
1-
12
#664100000000
0!
0%
b101 *
0-
02
b101 6
#664110000000
1!
1%
1-
12
#664120000000
0!
0%
b110 *
0-
02
b110 6
#664130000000
1!
1%
1-
12
#664140000000
0!
0%
b111 *
0-
02
b111 6
#664150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#664160000000
0!
0%
b0 *
0-
02
b0 6
#664170000000
1!
1%
1-
12
#664180000000
0!
0%
b1 *
0-
02
b1 6
#664190000000
1!
1%
1-
12
#664200000000
0!
0%
b10 *
0-
02
b10 6
#664210000000
1!
1%
1-
12
#664220000000
0!
0%
b11 *
0-
02
b11 6
#664230000000
1!
1%
1-
12
15
#664240000000
0!
0%
b100 *
0-
02
b100 6
#664250000000
1!
1%
1-
12
#664260000000
0!
0%
b101 *
0-
02
b101 6
#664270000000
1!
1%
1-
12
#664280000000
0!
0%
b110 *
0-
02
b110 6
#664290000000
1!
1%
1-
12
#664300000000
0!
0%
b111 *
0-
02
b111 6
#664310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#664320000000
0!
0%
b0 *
0-
02
b0 6
#664330000000
1!
1%
1-
12
#664340000000
0!
0%
b1 *
0-
02
b1 6
#664350000000
1!
1%
1-
12
#664360000000
0!
0%
b10 *
0-
02
b10 6
#664370000000
1!
1%
1-
12
#664380000000
0!
0%
b11 *
0-
02
b11 6
#664390000000
1!
1%
1-
12
15
#664400000000
0!
0%
b100 *
0-
02
b100 6
#664410000000
1!
1%
1-
12
#664420000000
0!
0%
b101 *
0-
02
b101 6
#664430000000
1!
1%
1-
12
#664440000000
0!
0%
b110 *
0-
02
b110 6
#664450000000
1!
1%
1-
12
#664460000000
0!
0%
b111 *
0-
02
b111 6
#664470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#664480000000
0!
0%
b0 *
0-
02
b0 6
#664490000000
1!
1%
1-
12
#664500000000
0!
0%
b1 *
0-
02
b1 6
#664510000000
1!
1%
1-
12
#664520000000
0!
0%
b10 *
0-
02
b10 6
#664530000000
1!
1%
1-
12
#664540000000
0!
0%
b11 *
0-
02
b11 6
#664550000000
1!
1%
1-
12
15
#664560000000
0!
0%
b100 *
0-
02
b100 6
#664570000000
1!
1%
1-
12
#664580000000
0!
0%
b101 *
0-
02
b101 6
#664590000000
1!
1%
1-
12
#664600000000
0!
0%
b110 *
0-
02
b110 6
#664610000000
1!
1%
1-
12
#664620000000
0!
0%
b111 *
0-
02
b111 6
#664630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#664640000000
0!
0%
b0 *
0-
02
b0 6
#664650000000
1!
1%
1-
12
#664660000000
0!
0%
b1 *
0-
02
b1 6
#664670000000
1!
1%
1-
12
#664680000000
0!
0%
b10 *
0-
02
b10 6
#664690000000
1!
1%
1-
12
#664700000000
0!
0%
b11 *
0-
02
b11 6
#664710000000
1!
1%
1-
12
15
#664720000000
0!
0%
b100 *
0-
02
b100 6
#664730000000
1!
1%
1-
12
#664740000000
0!
0%
b101 *
0-
02
b101 6
#664750000000
1!
1%
1-
12
#664760000000
0!
0%
b110 *
0-
02
b110 6
#664770000000
1!
1%
1-
12
#664780000000
0!
0%
b111 *
0-
02
b111 6
#664790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#664800000000
0!
0%
b0 *
0-
02
b0 6
#664810000000
1!
1%
1-
12
#664820000000
0!
0%
b1 *
0-
02
b1 6
#664830000000
1!
1%
1-
12
#664840000000
0!
0%
b10 *
0-
02
b10 6
#664850000000
1!
1%
1-
12
#664860000000
0!
0%
b11 *
0-
02
b11 6
#664870000000
1!
1%
1-
12
15
#664880000000
0!
0%
b100 *
0-
02
b100 6
#664890000000
1!
1%
1-
12
#664900000000
0!
0%
b101 *
0-
02
b101 6
#664910000000
1!
1%
1-
12
#664920000000
0!
0%
b110 *
0-
02
b110 6
#664930000000
1!
1%
1-
12
#664940000000
0!
0%
b111 *
0-
02
b111 6
#664950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#664960000000
0!
0%
b0 *
0-
02
b0 6
#664970000000
1!
1%
1-
12
#664980000000
0!
0%
b1 *
0-
02
b1 6
#664990000000
1!
1%
1-
12
#665000000000
0!
0%
b10 *
0-
02
b10 6
#665010000000
1!
1%
1-
12
#665020000000
0!
0%
b11 *
0-
02
b11 6
#665030000000
1!
1%
1-
12
15
#665040000000
0!
0%
b100 *
0-
02
b100 6
#665050000000
1!
1%
1-
12
#665060000000
0!
0%
b101 *
0-
02
b101 6
#665070000000
1!
1%
1-
12
#665080000000
0!
0%
b110 *
0-
02
b110 6
#665090000000
1!
1%
1-
12
#665100000000
0!
0%
b111 *
0-
02
b111 6
#665110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#665120000000
0!
0%
b0 *
0-
02
b0 6
#665130000000
1!
1%
1-
12
#665140000000
0!
0%
b1 *
0-
02
b1 6
#665150000000
1!
1%
1-
12
#665160000000
0!
0%
b10 *
0-
02
b10 6
#665170000000
1!
1%
1-
12
#665180000000
0!
0%
b11 *
0-
02
b11 6
#665190000000
1!
1%
1-
12
15
#665200000000
0!
0%
b100 *
0-
02
b100 6
#665210000000
1!
1%
1-
12
#665220000000
0!
0%
b101 *
0-
02
b101 6
#665230000000
1!
1%
1-
12
#665240000000
0!
0%
b110 *
0-
02
b110 6
#665250000000
1!
1%
1-
12
#665260000000
0!
0%
b111 *
0-
02
b111 6
#665270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#665280000000
0!
0%
b0 *
0-
02
b0 6
#665290000000
1!
1%
1-
12
#665300000000
0!
0%
b1 *
0-
02
b1 6
#665310000000
1!
1%
1-
12
#665320000000
0!
0%
b10 *
0-
02
b10 6
#665330000000
1!
1%
1-
12
#665340000000
0!
0%
b11 *
0-
02
b11 6
#665350000000
1!
1%
1-
12
15
#665360000000
0!
0%
b100 *
0-
02
b100 6
#665370000000
1!
1%
1-
12
#665380000000
0!
0%
b101 *
0-
02
b101 6
#665390000000
1!
1%
1-
12
#665400000000
0!
0%
b110 *
0-
02
b110 6
#665410000000
1!
1%
1-
12
#665420000000
0!
0%
b111 *
0-
02
b111 6
#665430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#665440000000
0!
0%
b0 *
0-
02
b0 6
#665450000000
1!
1%
1-
12
#665460000000
0!
0%
b1 *
0-
02
b1 6
#665470000000
1!
1%
1-
12
#665480000000
0!
0%
b10 *
0-
02
b10 6
#665490000000
1!
1%
1-
12
#665500000000
0!
0%
b11 *
0-
02
b11 6
#665510000000
1!
1%
1-
12
15
#665520000000
0!
0%
b100 *
0-
02
b100 6
#665530000000
1!
1%
1-
12
#665540000000
0!
0%
b101 *
0-
02
b101 6
#665550000000
1!
1%
1-
12
#665560000000
0!
0%
b110 *
0-
02
b110 6
#665570000000
1!
1%
1-
12
#665580000000
0!
0%
b111 *
0-
02
b111 6
#665590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#665600000000
0!
0%
b0 *
0-
02
b0 6
#665610000000
1!
1%
1-
12
#665620000000
0!
0%
b1 *
0-
02
b1 6
#665630000000
1!
1%
1-
12
#665640000000
0!
0%
b10 *
0-
02
b10 6
#665650000000
1!
1%
1-
12
#665660000000
0!
0%
b11 *
0-
02
b11 6
#665670000000
1!
1%
1-
12
15
#665680000000
0!
0%
b100 *
0-
02
b100 6
#665690000000
1!
1%
1-
12
#665700000000
0!
0%
b101 *
0-
02
b101 6
#665710000000
1!
1%
1-
12
#665720000000
0!
0%
b110 *
0-
02
b110 6
#665730000000
1!
1%
1-
12
#665740000000
0!
0%
b111 *
0-
02
b111 6
#665750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#665760000000
0!
0%
b0 *
0-
02
b0 6
#665770000000
1!
1%
1-
12
#665780000000
0!
0%
b1 *
0-
02
b1 6
#665790000000
1!
1%
1-
12
#665800000000
0!
0%
b10 *
0-
02
b10 6
#665810000000
1!
1%
1-
12
#665820000000
0!
0%
b11 *
0-
02
b11 6
#665830000000
1!
1%
1-
12
15
#665840000000
0!
0%
b100 *
0-
02
b100 6
#665850000000
1!
1%
1-
12
#665860000000
0!
0%
b101 *
0-
02
b101 6
#665870000000
1!
1%
1-
12
#665880000000
0!
0%
b110 *
0-
02
b110 6
#665890000000
1!
1%
1-
12
#665900000000
0!
0%
b111 *
0-
02
b111 6
#665910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#665920000000
0!
0%
b0 *
0-
02
b0 6
#665930000000
1!
1%
1-
12
#665940000000
0!
0%
b1 *
0-
02
b1 6
#665950000000
1!
1%
1-
12
#665960000000
0!
0%
b10 *
0-
02
b10 6
#665970000000
1!
1%
1-
12
#665980000000
0!
0%
b11 *
0-
02
b11 6
#665990000000
1!
1%
1-
12
15
#666000000000
0!
0%
b100 *
0-
02
b100 6
#666010000000
1!
1%
1-
12
#666020000000
0!
0%
b101 *
0-
02
b101 6
#666030000000
1!
1%
1-
12
#666040000000
0!
0%
b110 *
0-
02
b110 6
#666050000000
1!
1%
1-
12
#666060000000
0!
0%
b111 *
0-
02
b111 6
#666070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#666080000000
0!
0%
b0 *
0-
02
b0 6
#666090000000
1!
1%
1-
12
#666100000000
0!
0%
b1 *
0-
02
b1 6
#666110000000
1!
1%
1-
12
#666120000000
0!
0%
b10 *
0-
02
b10 6
#666130000000
1!
1%
1-
12
#666140000000
0!
0%
b11 *
0-
02
b11 6
#666150000000
1!
1%
1-
12
15
#666160000000
0!
0%
b100 *
0-
02
b100 6
#666170000000
1!
1%
1-
12
#666180000000
0!
0%
b101 *
0-
02
b101 6
#666190000000
1!
1%
1-
12
#666200000000
0!
0%
b110 *
0-
02
b110 6
#666210000000
1!
1%
1-
12
#666220000000
0!
0%
b111 *
0-
02
b111 6
#666230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#666240000000
0!
0%
b0 *
0-
02
b0 6
#666250000000
1!
1%
1-
12
#666260000000
0!
0%
b1 *
0-
02
b1 6
#666270000000
1!
1%
1-
12
#666280000000
0!
0%
b10 *
0-
02
b10 6
#666290000000
1!
1%
1-
12
#666300000000
0!
0%
b11 *
0-
02
b11 6
#666310000000
1!
1%
1-
12
15
#666320000000
0!
0%
b100 *
0-
02
b100 6
#666330000000
1!
1%
1-
12
#666340000000
0!
0%
b101 *
0-
02
b101 6
#666350000000
1!
1%
1-
12
#666360000000
0!
0%
b110 *
0-
02
b110 6
#666370000000
1!
1%
1-
12
#666380000000
0!
0%
b111 *
0-
02
b111 6
#666390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#666400000000
0!
0%
b0 *
0-
02
b0 6
#666410000000
1!
1%
1-
12
#666420000000
0!
0%
b1 *
0-
02
b1 6
#666430000000
1!
1%
1-
12
#666440000000
0!
0%
b10 *
0-
02
b10 6
#666450000000
1!
1%
1-
12
#666460000000
0!
0%
b11 *
0-
02
b11 6
#666470000000
1!
1%
1-
12
15
#666480000000
0!
0%
b100 *
0-
02
b100 6
#666490000000
1!
1%
1-
12
#666500000000
0!
0%
b101 *
0-
02
b101 6
#666510000000
1!
1%
1-
12
#666520000000
0!
0%
b110 *
0-
02
b110 6
#666530000000
1!
1%
1-
12
#666540000000
0!
0%
b111 *
0-
02
b111 6
#666550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#666560000000
0!
0%
b0 *
0-
02
b0 6
#666570000000
1!
1%
1-
12
#666580000000
0!
0%
b1 *
0-
02
b1 6
#666590000000
1!
1%
1-
12
#666600000000
0!
0%
b10 *
0-
02
b10 6
#666610000000
1!
1%
1-
12
#666620000000
0!
0%
b11 *
0-
02
b11 6
#666630000000
1!
1%
1-
12
15
#666640000000
0!
0%
b100 *
0-
02
b100 6
#666650000000
1!
1%
1-
12
#666660000000
0!
0%
b101 *
0-
02
b101 6
#666670000000
1!
1%
1-
12
#666680000000
0!
0%
b110 *
0-
02
b110 6
#666690000000
1!
1%
1-
12
#666700000000
0!
0%
b111 *
0-
02
b111 6
#666710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#666720000000
0!
0%
b0 *
0-
02
b0 6
#666730000000
1!
1%
1-
12
#666740000000
0!
0%
b1 *
0-
02
b1 6
#666750000000
1!
1%
1-
12
#666760000000
0!
0%
b10 *
0-
02
b10 6
#666770000000
1!
1%
1-
12
#666780000000
0!
0%
b11 *
0-
02
b11 6
#666790000000
1!
1%
1-
12
15
#666800000000
0!
0%
b100 *
0-
02
b100 6
#666810000000
1!
1%
1-
12
#666820000000
0!
0%
b101 *
0-
02
b101 6
#666830000000
1!
1%
1-
12
#666840000000
0!
0%
b110 *
0-
02
b110 6
#666850000000
1!
1%
1-
12
#666860000000
0!
0%
b111 *
0-
02
b111 6
#666870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#666880000000
0!
0%
b0 *
0-
02
b0 6
#666890000000
1!
1%
1-
12
#666900000000
0!
0%
b1 *
0-
02
b1 6
#666910000000
1!
1%
1-
12
#666920000000
0!
0%
b10 *
0-
02
b10 6
#666930000000
1!
1%
1-
12
#666940000000
0!
0%
b11 *
0-
02
b11 6
#666950000000
1!
1%
1-
12
15
#666960000000
0!
0%
b100 *
0-
02
b100 6
#666970000000
1!
1%
1-
12
#666980000000
0!
0%
b101 *
0-
02
b101 6
#666990000000
1!
1%
1-
12
#667000000000
0!
0%
b110 *
0-
02
b110 6
#667010000000
1!
1%
1-
12
#667020000000
0!
0%
b111 *
0-
02
b111 6
#667030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#667040000000
0!
0%
b0 *
0-
02
b0 6
#667050000000
1!
1%
1-
12
#667060000000
0!
0%
b1 *
0-
02
b1 6
#667070000000
1!
1%
1-
12
#667080000000
0!
0%
b10 *
0-
02
b10 6
#667090000000
1!
1%
1-
12
#667100000000
0!
0%
b11 *
0-
02
b11 6
#667110000000
1!
1%
1-
12
15
#667120000000
0!
0%
b100 *
0-
02
b100 6
#667130000000
1!
1%
1-
12
#667140000000
0!
0%
b101 *
0-
02
b101 6
#667150000000
1!
1%
1-
12
#667160000000
0!
0%
b110 *
0-
02
b110 6
#667170000000
1!
1%
1-
12
#667180000000
0!
0%
b111 *
0-
02
b111 6
#667190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#667200000000
0!
0%
b0 *
0-
02
b0 6
#667210000000
1!
1%
1-
12
#667220000000
0!
0%
b1 *
0-
02
b1 6
#667230000000
1!
1%
1-
12
#667240000000
0!
0%
b10 *
0-
02
b10 6
#667250000000
1!
1%
1-
12
#667260000000
0!
0%
b11 *
0-
02
b11 6
#667270000000
1!
1%
1-
12
15
#667280000000
0!
0%
b100 *
0-
02
b100 6
#667290000000
1!
1%
1-
12
#667300000000
0!
0%
b101 *
0-
02
b101 6
#667310000000
1!
1%
1-
12
#667320000000
0!
0%
b110 *
0-
02
b110 6
#667330000000
1!
1%
1-
12
#667340000000
0!
0%
b111 *
0-
02
b111 6
#667350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#667360000000
0!
0%
b0 *
0-
02
b0 6
#667370000000
1!
1%
1-
12
#667380000000
0!
0%
b1 *
0-
02
b1 6
#667390000000
1!
1%
1-
12
#667400000000
0!
0%
b10 *
0-
02
b10 6
#667410000000
1!
1%
1-
12
#667420000000
0!
0%
b11 *
0-
02
b11 6
#667430000000
1!
1%
1-
12
15
#667440000000
0!
0%
b100 *
0-
02
b100 6
#667450000000
1!
1%
1-
12
#667460000000
0!
0%
b101 *
0-
02
b101 6
#667470000000
1!
1%
1-
12
#667480000000
0!
0%
b110 *
0-
02
b110 6
#667490000000
1!
1%
1-
12
#667500000000
0!
0%
b111 *
0-
02
b111 6
#667510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#667520000000
0!
0%
b0 *
0-
02
b0 6
#667530000000
1!
1%
1-
12
#667540000000
0!
0%
b1 *
0-
02
b1 6
#667550000000
1!
1%
1-
12
#667560000000
0!
0%
b10 *
0-
02
b10 6
#667570000000
1!
1%
1-
12
#667580000000
0!
0%
b11 *
0-
02
b11 6
#667590000000
1!
1%
1-
12
15
#667600000000
0!
0%
b100 *
0-
02
b100 6
#667610000000
1!
1%
1-
12
#667620000000
0!
0%
b101 *
0-
02
b101 6
#667630000000
1!
1%
1-
12
#667640000000
0!
0%
b110 *
0-
02
b110 6
#667650000000
1!
1%
1-
12
#667660000000
0!
0%
b111 *
0-
02
b111 6
#667670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#667680000000
0!
0%
b0 *
0-
02
b0 6
#667690000000
1!
1%
1-
12
#667700000000
0!
0%
b1 *
0-
02
b1 6
#667710000000
1!
1%
1-
12
#667720000000
0!
0%
b10 *
0-
02
b10 6
#667730000000
1!
1%
1-
12
#667740000000
0!
0%
b11 *
0-
02
b11 6
#667750000000
1!
1%
1-
12
15
#667760000000
0!
0%
b100 *
0-
02
b100 6
#667770000000
1!
1%
1-
12
#667780000000
0!
0%
b101 *
0-
02
b101 6
#667790000000
1!
1%
1-
12
#667800000000
0!
0%
b110 *
0-
02
b110 6
#667810000000
1!
1%
1-
12
#667820000000
0!
0%
b111 *
0-
02
b111 6
#667830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#667840000000
0!
0%
b0 *
0-
02
b0 6
#667850000000
1!
1%
1-
12
#667860000000
0!
0%
b1 *
0-
02
b1 6
#667870000000
1!
1%
1-
12
#667880000000
0!
0%
b10 *
0-
02
b10 6
#667890000000
1!
1%
1-
12
#667900000000
0!
0%
b11 *
0-
02
b11 6
#667910000000
1!
1%
1-
12
15
#667920000000
0!
0%
b100 *
0-
02
b100 6
#667930000000
1!
1%
1-
12
#667940000000
0!
0%
b101 *
0-
02
b101 6
#667950000000
1!
1%
1-
12
#667960000000
0!
0%
b110 *
0-
02
b110 6
#667970000000
1!
1%
1-
12
#667980000000
0!
0%
b111 *
0-
02
b111 6
#667990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#668000000000
0!
0%
b0 *
0-
02
b0 6
#668010000000
1!
1%
1-
12
#668020000000
0!
0%
b1 *
0-
02
b1 6
#668030000000
1!
1%
1-
12
#668040000000
0!
0%
b10 *
0-
02
b10 6
#668050000000
1!
1%
1-
12
#668060000000
0!
0%
b11 *
0-
02
b11 6
#668070000000
1!
1%
1-
12
15
#668080000000
0!
0%
b100 *
0-
02
b100 6
#668090000000
1!
1%
1-
12
#668100000000
0!
0%
b101 *
0-
02
b101 6
#668110000000
1!
1%
1-
12
#668120000000
0!
0%
b110 *
0-
02
b110 6
#668130000000
1!
1%
1-
12
#668140000000
0!
0%
b111 *
0-
02
b111 6
#668150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#668160000000
0!
0%
b0 *
0-
02
b0 6
#668170000000
1!
1%
1-
12
#668180000000
0!
0%
b1 *
0-
02
b1 6
#668190000000
1!
1%
1-
12
#668200000000
0!
0%
b10 *
0-
02
b10 6
#668210000000
1!
1%
1-
12
#668220000000
0!
0%
b11 *
0-
02
b11 6
#668230000000
1!
1%
1-
12
15
#668240000000
0!
0%
b100 *
0-
02
b100 6
#668250000000
1!
1%
1-
12
#668260000000
0!
0%
b101 *
0-
02
b101 6
#668270000000
1!
1%
1-
12
#668280000000
0!
0%
b110 *
0-
02
b110 6
#668290000000
1!
1%
1-
12
#668300000000
0!
0%
b111 *
0-
02
b111 6
#668310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#668320000000
0!
0%
b0 *
0-
02
b0 6
#668330000000
1!
1%
1-
12
#668340000000
0!
0%
b1 *
0-
02
b1 6
#668350000000
1!
1%
1-
12
#668360000000
0!
0%
b10 *
0-
02
b10 6
#668370000000
1!
1%
1-
12
#668380000000
0!
0%
b11 *
0-
02
b11 6
#668390000000
1!
1%
1-
12
15
#668400000000
0!
0%
b100 *
0-
02
b100 6
#668410000000
1!
1%
1-
12
#668420000000
0!
0%
b101 *
0-
02
b101 6
#668430000000
1!
1%
1-
12
#668440000000
0!
0%
b110 *
0-
02
b110 6
#668450000000
1!
1%
1-
12
#668460000000
0!
0%
b111 *
0-
02
b111 6
#668470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#668480000000
0!
0%
b0 *
0-
02
b0 6
#668490000000
1!
1%
1-
12
#668500000000
0!
0%
b1 *
0-
02
b1 6
#668510000000
1!
1%
1-
12
#668520000000
0!
0%
b10 *
0-
02
b10 6
#668530000000
1!
1%
1-
12
#668540000000
0!
0%
b11 *
0-
02
b11 6
#668550000000
1!
1%
1-
12
15
#668560000000
0!
0%
b100 *
0-
02
b100 6
#668570000000
1!
1%
1-
12
#668580000000
0!
0%
b101 *
0-
02
b101 6
#668590000000
1!
1%
1-
12
#668600000000
0!
0%
b110 *
0-
02
b110 6
#668610000000
1!
1%
1-
12
#668620000000
0!
0%
b111 *
0-
02
b111 6
#668630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#668640000000
0!
0%
b0 *
0-
02
b0 6
#668650000000
1!
1%
1-
12
#668660000000
0!
0%
b1 *
0-
02
b1 6
#668670000000
1!
1%
1-
12
#668680000000
0!
0%
b10 *
0-
02
b10 6
#668690000000
1!
1%
1-
12
#668700000000
0!
0%
b11 *
0-
02
b11 6
#668710000000
1!
1%
1-
12
15
#668720000000
0!
0%
b100 *
0-
02
b100 6
#668730000000
1!
1%
1-
12
#668740000000
0!
0%
b101 *
0-
02
b101 6
#668750000000
1!
1%
1-
12
#668760000000
0!
0%
b110 *
0-
02
b110 6
#668770000000
1!
1%
1-
12
#668780000000
0!
0%
b111 *
0-
02
b111 6
#668790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#668800000000
0!
0%
b0 *
0-
02
b0 6
#668810000000
1!
1%
1-
12
#668820000000
0!
0%
b1 *
0-
02
b1 6
#668830000000
1!
1%
1-
12
#668840000000
0!
0%
b10 *
0-
02
b10 6
#668850000000
1!
1%
1-
12
#668860000000
0!
0%
b11 *
0-
02
b11 6
#668870000000
1!
1%
1-
12
15
#668880000000
0!
0%
b100 *
0-
02
b100 6
#668890000000
1!
1%
1-
12
#668900000000
0!
0%
b101 *
0-
02
b101 6
#668910000000
1!
1%
1-
12
#668920000000
0!
0%
b110 *
0-
02
b110 6
#668930000000
1!
1%
1-
12
#668940000000
0!
0%
b111 *
0-
02
b111 6
#668950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#668960000000
0!
0%
b0 *
0-
02
b0 6
#668970000000
1!
1%
1-
12
#668980000000
0!
0%
b1 *
0-
02
b1 6
#668990000000
1!
1%
1-
12
#669000000000
0!
0%
b10 *
0-
02
b10 6
#669010000000
1!
1%
1-
12
#669020000000
0!
0%
b11 *
0-
02
b11 6
#669030000000
1!
1%
1-
12
15
#669040000000
0!
0%
b100 *
0-
02
b100 6
#669050000000
1!
1%
1-
12
#669060000000
0!
0%
b101 *
0-
02
b101 6
#669070000000
1!
1%
1-
12
#669080000000
0!
0%
b110 *
0-
02
b110 6
#669090000000
1!
1%
1-
12
#669100000000
0!
0%
b111 *
0-
02
b111 6
#669110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#669120000000
0!
0%
b0 *
0-
02
b0 6
#669130000000
1!
1%
1-
12
#669140000000
0!
0%
b1 *
0-
02
b1 6
#669150000000
1!
1%
1-
12
#669160000000
0!
0%
b10 *
0-
02
b10 6
#669170000000
1!
1%
1-
12
#669180000000
0!
0%
b11 *
0-
02
b11 6
#669190000000
1!
1%
1-
12
15
#669200000000
0!
0%
b100 *
0-
02
b100 6
#669210000000
1!
1%
1-
12
#669220000000
0!
0%
b101 *
0-
02
b101 6
#669230000000
1!
1%
1-
12
#669240000000
0!
0%
b110 *
0-
02
b110 6
#669250000000
1!
1%
1-
12
#669260000000
0!
0%
b111 *
0-
02
b111 6
#669270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#669280000000
0!
0%
b0 *
0-
02
b0 6
#669290000000
1!
1%
1-
12
#669300000000
0!
0%
b1 *
0-
02
b1 6
#669310000000
1!
1%
1-
12
#669320000000
0!
0%
b10 *
0-
02
b10 6
#669330000000
1!
1%
1-
12
#669340000000
0!
0%
b11 *
0-
02
b11 6
#669350000000
1!
1%
1-
12
15
#669360000000
0!
0%
b100 *
0-
02
b100 6
#669370000000
1!
1%
1-
12
#669380000000
0!
0%
b101 *
0-
02
b101 6
#669390000000
1!
1%
1-
12
#669400000000
0!
0%
b110 *
0-
02
b110 6
#669410000000
1!
1%
1-
12
#669420000000
0!
0%
b111 *
0-
02
b111 6
#669430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#669440000000
0!
0%
b0 *
0-
02
b0 6
#669450000000
1!
1%
1-
12
#669460000000
0!
0%
b1 *
0-
02
b1 6
#669470000000
1!
1%
1-
12
#669480000000
0!
0%
b10 *
0-
02
b10 6
#669490000000
1!
1%
1-
12
#669500000000
0!
0%
b11 *
0-
02
b11 6
#669510000000
1!
1%
1-
12
15
#669520000000
0!
0%
b100 *
0-
02
b100 6
#669530000000
1!
1%
1-
12
#669540000000
0!
0%
b101 *
0-
02
b101 6
#669550000000
1!
1%
1-
12
#669560000000
0!
0%
b110 *
0-
02
b110 6
#669570000000
1!
1%
1-
12
#669580000000
0!
0%
b111 *
0-
02
b111 6
#669590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#669600000000
0!
0%
b0 *
0-
02
b0 6
#669610000000
1!
1%
1-
12
#669620000000
0!
0%
b1 *
0-
02
b1 6
#669630000000
1!
1%
1-
12
#669640000000
0!
0%
b10 *
0-
02
b10 6
#669650000000
1!
1%
1-
12
#669660000000
0!
0%
b11 *
0-
02
b11 6
#669670000000
1!
1%
1-
12
15
#669680000000
0!
0%
b100 *
0-
02
b100 6
#669690000000
1!
1%
1-
12
#669700000000
0!
0%
b101 *
0-
02
b101 6
#669710000000
1!
1%
1-
12
#669720000000
0!
0%
b110 *
0-
02
b110 6
#669730000000
1!
1%
1-
12
#669740000000
0!
0%
b111 *
0-
02
b111 6
#669750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#669760000000
0!
0%
b0 *
0-
02
b0 6
#669770000000
1!
1%
1-
12
#669780000000
0!
0%
b1 *
0-
02
b1 6
#669790000000
1!
1%
1-
12
#669800000000
0!
0%
b10 *
0-
02
b10 6
#669810000000
1!
1%
1-
12
#669820000000
0!
0%
b11 *
0-
02
b11 6
#669830000000
1!
1%
1-
12
15
#669840000000
0!
0%
b100 *
0-
02
b100 6
#669850000000
1!
1%
1-
12
#669860000000
0!
0%
b101 *
0-
02
b101 6
#669870000000
1!
1%
1-
12
#669880000000
0!
0%
b110 *
0-
02
b110 6
#669890000000
1!
1%
1-
12
#669900000000
0!
0%
b111 *
0-
02
b111 6
#669910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#669920000000
0!
0%
b0 *
0-
02
b0 6
#669930000000
1!
1%
1-
12
#669940000000
0!
0%
b1 *
0-
02
b1 6
#669950000000
1!
1%
1-
12
#669960000000
0!
0%
b10 *
0-
02
b10 6
#669970000000
1!
1%
1-
12
#669980000000
0!
0%
b11 *
0-
02
b11 6
#669990000000
1!
1%
1-
12
15
#670000000000
0!
0%
b100 *
0-
02
b100 6
#670010000000
1!
1%
1-
12
#670020000000
0!
0%
b101 *
0-
02
b101 6
#670030000000
1!
1%
1-
12
#670040000000
0!
0%
b110 *
0-
02
b110 6
#670050000000
1!
1%
1-
12
#670060000000
0!
0%
b111 *
0-
02
b111 6
#670070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#670080000000
0!
0%
b0 *
0-
02
b0 6
#670090000000
1!
1%
1-
12
#670100000000
0!
0%
b1 *
0-
02
b1 6
#670110000000
1!
1%
1-
12
#670120000000
0!
0%
b10 *
0-
02
b10 6
#670130000000
1!
1%
1-
12
#670140000000
0!
0%
b11 *
0-
02
b11 6
#670150000000
1!
1%
1-
12
15
#670160000000
0!
0%
b100 *
0-
02
b100 6
#670170000000
1!
1%
1-
12
#670180000000
0!
0%
b101 *
0-
02
b101 6
#670190000000
1!
1%
1-
12
#670200000000
0!
0%
b110 *
0-
02
b110 6
#670210000000
1!
1%
1-
12
#670220000000
0!
0%
b111 *
0-
02
b111 6
#670230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#670240000000
0!
0%
b0 *
0-
02
b0 6
#670250000000
1!
1%
1-
12
#670260000000
0!
0%
b1 *
0-
02
b1 6
#670270000000
1!
1%
1-
12
#670280000000
0!
0%
b10 *
0-
02
b10 6
#670290000000
1!
1%
1-
12
#670300000000
0!
0%
b11 *
0-
02
b11 6
#670310000000
1!
1%
1-
12
15
#670320000000
0!
0%
b100 *
0-
02
b100 6
#670330000000
1!
1%
1-
12
#670340000000
0!
0%
b101 *
0-
02
b101 6
#670350000000
1!
1%
1-
12
#670360000000
0!
0%
b110 *
0-
02
b110 6
#670370000000
1!
1%
1-
12
#670380000000
0!
0%
b111 *
0-
02
b111 6
#670390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#670400000000
0!
0%
b0 *
0-
02
b0 6
#670410000000
1!
1%
1-
12
#670420000000
0!
0%
b1 *
0-
02
b1 6
#670430000000
1!
1%
1-
12
#670440000000
0!
0%
b10 *
0-
02
b10 6
#670450000000
1!
1%
1-
12
#670460000000
0!
0%
b11 *
0-
02
b11 6
#670470000000
1!
1%
1-
12
15
#670480000000
0!
0%
b100 *
0-
02
b100 6
#670490000000
1!
1%
1-
12
#670500000000
0!
0%
b101 *
0-
02
b101 6
#670510000000
1!
1%
1-
12
#670520000000
0!
0%
b110 *
0-
02
b110 6
#670530000000
1!
1%
1-
12
#670540000000
0!
0%
b111 *
0-
02
b111 6
#670550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#670560000000
0!
0%
b0 *
0-
02
b0 6
#670570000000
1!
1%
1-
12
#670580000000
0!
0%
b1 *
0-
02
b1 6
#670590000000
1!
1%
1-
12
#670600000000
0!
0%
b10 *
0-
02
b10 6
#670610000000
1!
1%
1-
12
#670620000000
0!
0%
b11 *
0-
02
b11 6
#670630000000
1!
1%
1-
12
15
#670640000000
0!
0%
b100 *
0-
02
b100 6
#670650000000
1!
1%
1-
12
#670660000000
0!
0%
b101 *
0-
02
b101 6
#670670000000
1!
1%
1-
12
#670680000000
0!
0%
b110 *
0-
02
b110 6
#670690000000
1!
1%
1-
12
#670700000000
0!
0%
b111 *
0-
02
b111 6
#670710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#670720000000
0!
0%
b0 *
0-
02
b0 6
#670730000000
1!
1%
1-
12
#670740000000
0!
0%
b1 *
0-
02
b1 6
#670750000000
1!
1%
1-
12
#670760000000
0!
0%
b10 *
0-
02
b10 6
#670770000000
1!
1%
1-
12
#670780000000
0!
0%
b11 *
0-
02
b11 6
#670790000000
1!
1%
1-
12
15
#670800000000
0!
0%
b100 *
0-
02
b100 6
#670810000000
1!
1%
1-
12
#670820000000
0!
0%
b101 *
0-
02
b101 6
#670830000000
1!
1%
1-
12
#670840000000
0!
0%
b110 *
0-
02
b110 6
#670850000000
1!
1%
1-
12
#670860000000
0!
0%
b111 *
0-
02
b111 6
#670870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#670880000000
0!
0%
b0 *
0-
02
b0 6
#670890000000
1!
1%
1-
12
#670900000000
0!
0%
b1 *
0-
02
b1 6
#670910000000
1!
1%
1-
12
#670920000000
0!
0%
b10 *
0-
02
b10 6
#670930000000
1!
1%
1-
12
#670940000000
0!
0%
b11 *
0-
02
b11 6
#670950000000
1!
1%
1-
12
15
#670960000000
0!
0%
b100 *
0-
02
b100 6
#670970000000
1!
1%
1-
12
#670980000000
0!
0%
b101 *
0-
02
b101 6
#670990000000
1!
1%
1-
12
#671000000000
0!
0%
b110 *
0-
02
b110 6
#671010000000
1!
1%
1-
12
#671020000000
0!
0%
b111 *
0-
02
b111 6
#671030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#671040000000
0!
0%
b0 *
0-
02
b0 6
#671050000000
1!
1%
1-
12
#671060000000
0!
0%
b1 *
0-
02
b1 6
#671070000000
1!
1%
1-
12
#671080000000
0!
0%
b10 *
0-
02
b10 6
#671090000000
1!
1%
1-
12
#671100000000
0!
0%
b11 *
0-
02
b11 6
#671110000000
1!
1%
1-
12
15
#671120000000
0!
0%
b100 *
0-
02
b100 6
#671130000000
1!
1%
1-
12
#671140000000
0!
0%
b101 *
0-
02
b101 6
#671150000000
1!
1%
1-
12
#671160000000
0!
0%
b110 *
0-
02
b110 6
#671170000000
1!
1%
1-
12
#671180000000
0!
0%
b111 *
0-
02
b111 6
#671190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#671200000000
0!
0%
b0 *
0-
02
b0 6
#671210000000
1!
1%
1-
12
#671220000000
0!
0%
b1 *
0-
02
b1 6
#671230000000
1!
1%
1-
12
#671240000000
0!
0%
b10 *
0-
02
b10 6
#671250000000
1!
1%
1-
12
#671260000000
0!
0%
b11 *
0-
02
b11 6
#671270000000
1!
1%
1-
12
15
#671280000000
0!
0%
b100 *
0-
02
b100 6
#671290000000
1!
1%
1-
12
#671300000000
0!
0%
b101 *
0-
02
b101 6
#671310000000
1!
1%
1-
12
#671320000000
0!
0%
b110 *
0-
02
b110 6
#671330000000
1!
1%
1-
12
#671340000000
0!
0%
b111 *
0-
02
b111 6
#671350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#671360000000
0!
0%
b0 *
0-
02
b0 6
#671370000000
1!
1%
1-
12
#671380000000
0!
0%
b1 *
0-
02
b1 6
#671390000000
1!
1%
1-
12
#671400000000
0!
0%
b10 *
0-
02
b10 6
#671410000000
1!
1%
1-
12
#671420000000
0!
0%
b11 *
0-
02
b11 6
#671430000000
1!
1%
1-
12
15
#671440000000
0!
0%
b100 *
0-
02
b100 6
#671450000000
1!
1%
1-
12
#671460000000
0!
0%
b101 *
0-
02
b101 6
#671470000000
1!
1%
1-
12
#671480000000
0!
0%
b110 *
0-
02
b110 6
#671490000000
1!
1%
1-
12
#671500000000
0!
0%
b111 *
0-
02
b111 6
#671510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#671520000000
0!
0%
b0 *
0-
02
b0 6
#671530000000
1!
1%
1-
12
#671540000000
0!
0%
b1 *
0-
02
b1 6
#671550000000
1!
1%
1-
12
#671560000000
0!
0%
b10 *
0-
02
b10 6
#671570000000
1!
1%
1-
12
#671580000000
0!
0%
b11 *
0-
02
b11 6
#671590000000
1!
1%
1-
12
15
#671600000000
0!
0%
b100 *
0-
02
b100 6
#671610000000
1!
1%
1-
12
#671620000000
0!
0%
b101 *
0-
02
b101 6
#671630000000
1!
1%
1-
12
#671640000000
0!
0%
b110 *
0-
02
b110 6
#671650000000
1!
1%
1-
12
#671660000000
0!
0%
b111 *
0-
02
b111 6
#671670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#671680000000
0!
0%
b0 *
0-
02
b0 6
#671690000000
1!
1%
1-
12
#671700000000
0!
0%
b1 *
0-
02
b1 6
#671710000000
1!
1%
1-
12
#671720000000
0!
0%
b10 *
0-
02
b10 6
#671730000000
1!
1%
1-
12
#671740000000
0!
0%
b11 *
0-
02
b11 6
#671750000000
1!
1%
1-
12
15
#671760000000
0!
0%
b100 *
0-
02
b100 6
#671770000000
1!
1%
1-
12
#671780000000
0!
0%
b101 *
0-
02
b101 6
#671790000000
1!
1%
1-
12
#671800000000
0!
0%
b110 *
0-
02
b110 6
#671810000000
1!
1%
1-
12
#671820000000
0!
0%
b111 *
0-
02
b111 6
#671830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#671840000000
0!
0%
b0 *
0-
02
b0 6
#671850000000
1!
1%
1-
12
#671860000000
0!
0%
b1 *
0-
02
b1 6
#671870000000
1!
1%
1-
12
#671880000000
0!
0%
b10 *
0-
02
b10 6
#671890000000
1!
1%
1-
12
#671900000000
0!
0%
b11 *
0-
02
b11 6
#671910000000
1!
1%
1-
12
15
#671920000000
0!
0%
b100 *
0-
02
b100 6
#671930000000
1!
1%
1-
12
#671940000000
0!
0%
b101 *
0-
02
b101 6
#671950000000
1!
1%
1-
12
#671960000000
0!
0%
b110 *
0-
02
b110 6
#671970000000
1!
1%
1-
12
#671980000000
0!
0%
b111 *
0-
02
b111 6
#671990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#672000000000
0!
0%
b0 *
0-
02
b0 6
#672010000000
1!
1%
1-
12
#672020000000
0!
0%
b1 *
0-
02
b1 6
#672030000000
1!
1%
1-
12
#672040000000
0!
0%
b10 *
0-
02
b10 6
#672050000000
1!
1%
1-
12
#672060000000
0!
0%
b11 *
0-
02
b11 6
#672070000000
1!
1%
1-
12
15
#672080000000
0!
0%
b100 *
0-
02
b100 6
#672090000000
1!
1%
1-
12
#672100000000
0!
0%
b101 *
0-
02
b101 6
#672110000000
1!
1%
1-
12
#672120000000
0!
0%
b110 *
0-
02
b110 6
#672130000000
1!
1%
1-
12
#672140000000
0!
0%
b111 *
0-
02
b111 6
#672150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#672160000000
0!
0%
b0 *
0-
02
b0 6
#672170000000
1!
1%
1-
12
#672180000000
0!
0%
b1 *
0-
02
b1 6
#672190000000
1!
1%
1-
12
#672200000000
0!
0%
b10 *
0-
02
b10 6
#672210000000
1!
1%
1-
12
#672220000000
0!
0%
b11 *
0-
02
b11 6
#672230000000
1!
1%
1-
12
15
#672240000000
0!
0%
b100 *
0-
02
b100 6
#672250000000
1!
1%
1-
12
#672260000000
0!
0%
b101 *
0-
02
b101 6
#672270000000
1!
1%
1-
12
#672280000000
0!
0%
b110 *
0-
02
b110 6
#672290000000
1!
1%
1-
12
#672300000000
0!
0%
b111 *
0-
02
b111 6
#672310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#672320000000
0!
0%
b0 *
0-
02
b0 6
#672330000000
1!
1%
1-
12
#672340000000
0!
0%
b1 *
0-
02
b1 6
#672350000000
1!
1%
1-
12
#672360000000
0!
0%
b10 *
0-
02
b10 6
#672370000000
1!
1%
1-
12
#672380000000
0!
0%
b11 *
0-
02
b11 6
#672390000000
1!
1%
1-
12
15
#672400000000
0!
0%
b100 *
0-
02
b100 6
#672410000000
1!
1%
1-
12
#672420000000
0!
0%
b101 *
0-
02
b101 6
#672430000000
1!
1%
1-
12
#672440000000
0!
0%
b110 *
0-
02
b110 6
#672450000000
1!
1%
1-
12
#672460000000
0!
0%
b111 *
0-
02
b111 6
#672470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#672480000000
0!
0%
b0 *
0-
02
b0 6
#672490000000
1!
1%
1-
12
#672500000000
0!
0%
b1 *
0-
02
b1 6
#672510000000
1!
1%
1-
12
#672520000000
0!
0%
b10 *
0-
02
b10 6
#672530000000
1!
1%
1-
12
#672540000000
0!
0%
b11 *
0-
02
b11 6
#672550000000
1!
1%
1-
12
15
#672560000000
0!
0%
b100 *
0-
02
b100 6
#672570000000
1!
1%
1-
12
#672580000000
0!
0%
b101 *
0-
02
b101 6
#672590000000
1!
1%
1-
12
#672600000000
0!
0%
b110 *
0-
02
b110 6
#672610000000
1!
1%
1-
12
#672620000000
0!
0%
b111 *
0-
02
b111 6
#672630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#672640000000
0!
0%
b0 *
0-
02
b0 6
#672650000000
1!
1%
1-
12
#672660000000
0!
0%
b1 *
0-
02
b1 6
#672670000000
1!
1%
1-
12
#672680000000
0!
0%
b10 *
0-
02
b10 6
#672690000000
1!
1%
1-
12
#672700000000
0!
0%
b11 *
0-
02
b11 6
#672710000000
1!
1%
1-
12
15
#672720000000
0!
0%
b100 *
0-
02
b100 6
#672730000000
1!
1%
1-
12
#672740000000
0!
0%
b101 *
0-
02
b101 6
#672750000000
1!
1%
1-
12
#672760000000
0!
0%
b110 *
0-
02
b110 6
#672770000000
1!
1%
1-
12
#672780000000
0!
0%
b111 *
0-
02
b111 6
#672790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#672800000000
0!
0%
b0 *
0-
02
b0 6
#672810000000
1!
1%
1-
12
#672820000000
0!
0%
b1 *
0-
02
b1 6
#672830000000
1!
1%
1-
12
#672840000000
0!
0%
b10 *
0-
02
b10 6
#672850000000
1!
1%
1-
12
#672860000000
0!
0%
b11 *
0-
02
b11 6
#672870000000
1!
1%
1-
12
15
#672880000000
0!
0%
b100 *
0-
02
b100 6
#672890000000
1!
1%
1-
12
#672900000000
0!
0%
b101 *
0-
02
b101 6
#672910000000
1!
1%
1-
12
#672920000000
0!
0%
b110 *
0-
02
b110 6
#672930000000
1!
1%
1-
12
#672940000000
0!
0%
b111 *
0-
02
b111 6
#672950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#672960000000
0!
0%
b0 *
0-
02
b0 6
#672970000000
1!
1%
1-
12
#672980000000
0!
0%
b1 *
0-
02
b1 6
#672990000000
1!
1%
1-
12
#673000000000
0!
0%
b10 *
0-
02
b10 6
#673010000000
1!
1%
1-
12
#673020000000
0!
0%
b11 *
0-
02
b11 6
#673030000000
1!
1%
1-
12
15
#673040000000
0!
0%
b100 *
0-
02
b100 6
#673050000000
1!
1%
1-
12
#673060000000
0!
0%
b101 *
0-
02
b101 6
#673070000000
1!
1%
1-
12
#673080000000
0!
0%
b110 *
0-
02
b110 6
#673090000000
1!
1%
1-
12
#673100000000
0!
0%
b111 *
0-
02
b111 6
#673110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#673120000000
0!
0%
b0 *
0-
02
b0 6
#673130000000
1!
1%
1-
12
#673140000000
0!
0%
b1 *
0-
02
b1 6
#673150000000
1!
1%
1-
12
#673160000000
0!
0%
b10 *
0-
02
b10 6
#673170000000
1!
1%
1-
12
#673180000000
0!
0%
b11 *
0-
02
b11 6
#673190000000
1!
1%
1-
12
15
#673200000000
0!
0%
b100 *
0-
02
b100 6
#673210000000
1!
1%
1-
12
#673220000000
0!
0%
b101 *
0-
02
b101 6
#673230000000
1!
1%
1-
12
#673240000000
0!
0%
b110 *
0-
02
b110 6
#673250000000
1!
1%
1-
12
#673260000000
0!
0%
b111 *
0-
02
b111 6
#673270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#673280000000
0!
0%
b0 *
0-
02
b0 6
#673290000000
1!
1%
1-
12
#673300000000
0!
0%
b1 *
0-
02
b1 6
#673310000000
1!
1%
1-
12
#673320000000
0!
0%
b10 *
0-
02
b10 6
#673330000000
1!
1%
1-
12
#673340000000
0!
0%
b11 *
0-
02
b11 6
#673350000000
1!
1%
1-
12
15
#673360000000
0!
0%
b100 *
0-
02
b100 6
#673370000000
1!
1%
1-
12
#673380000000
0!
0%
b101 *
0-
02
b101 6
#673390000000
1!
1%
1-
12
#673400000000
0!
0%
b110 *
0-
02
b110 6
#673410000000
1!
1%
1-
12
#673420000000
0!
0%
b111 *
0-
02
b111 6
#673430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#673440000000
0!
0%
b0 *
0-
02
b0 6
#673450000000
1!
1%
1-
12
#673460000000
0!
0%
b1 *
0-
02
b1 6
#673470000000
1!
1%
1-
12
#673480000000
0!
0%
b10 *
0-
02
b10 6
#673490000000
1!
1%
1-
12
#673500000000
0!
0%
b11 *
0-
02
b11 6
#673510000000
1!
1%
1-
12
15
#673520000000
0!
0%
b100 *
0-
02
b100 6
#673530000000
1!
1%
1-
12
#673540000000
0!
0%
b101 *
0-
02
b101 6
#673550000000
1!
1%
1-
12
#673560000000
0!
0%
b110 *
0-
02
b110 6
#673570000000
1!
1%
1-
12
#673580000000
0!
0%
b111 *
0-
02
b111 6
#673590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#673600000000
0!
0%
b0 *
0-
02
b0 6
#673610000000
1!
1%
1-
12
#673620000000
0!
0%
b1 *
0-
02
b1 6
#673630000000
1!
1%
1-
12
#673640000000
0!
0%
b10 *
0-
02
b10 6
#673650000000
1!
1%
1-
12
#673660000000
0!
0%
b11 *
0-
02
b11 6
#673670000000
1!
1%
1-
12
15
#673680000000
0!
0%
b100 *
0-
02
b100 6
#673690000000
1!
1%
1-
12
#673700000000
0!
0%
b101 *
0-
02
b101 6
#673710000000
1!
1%
1-
12
#673720000000
0!
0%
b110 *
0-
02
b110 6
#673730000000
1!
1%
1-
12
#673740000000
0!
0%
b111 *
0-
02
b111 6
#673750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#673760000000
0!
0%
b0 *
0-
02
b0 6
#673770000000
1!
1%
1-
12
#673780000000
0!
0%
b1 *
0-
02
b1 6
#673790000000
1!
1%
1-
12
#673800000000
0!
0%
b10 *
0-
02
b10 6
#673810000000
1!
1%
1-
12
#673820000000
0!
0%
b11 *
0-
02
b11 6
#673830000000
1!
1%
1-
12
15
#673840000000
0!
0%
b100 *
0-
02
b100 6
#673850000000
1!
1%
1-
12
#673860000000
0!
0%
b101 *
0-
02
b101 6
#673870000000
1!
1%
1-
12
#673880000000
0!
0%
b110 *
0-
02
b110 6
#673890000000
1!
1%
1-
12
#673900000000
0!
0%
b111 *
0-
02
b111 6
#673910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#673920000000
0!
0%
b0 *
0-
02
b0 6
#673930000000
1!
1%
1-
12
#673940000000
0!
0%
b1 *
0-
02
b1 6
#673950000000
1!
1%
1-
12
#673960000000
0!
0%
b10 *
0-
02
b10 6
#673970000000
1!
1%
1-
12
#673980000000
0!
0%
b11 *
0-
02
b11 6
#673990000000
1!
1%
1-
12
15
#674000000000
0!
0%
b100 *
0-
02
b100 6
#674010000000
1!
1%
1-
12
#674020000000
0!
0%
b101 *
0-
02
b101 6
#674030000000
1!
1%
1-
12
#674040000000
0!
0%
b110 *
0-
02
b110 6
#674050000000
1!
1%
1-
12
#674060000000
0!
0%
b111 *
0-
02
b111 6
#674070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#674080000000
0!
0%
b0 *
0-
02
b0 6
#674090000000
1!
1%
1-
12
#674100000000
0!
0%
b1 *
0-
02
b1 6
#674110000000
1!
1%
1-
12
#674120000000
0!
0%
b10 *
0-
02
b10 6
#674130000000
1!
1%
1-
12
#674140000000
0!
0%
b11 *
0-
02
b11 6
#674150000000
1!
1%
1-
12
15
#674160000000
0!
0%
b100 *
0-
02
b100 6
#674170000000
1!
1%
1-
12
#674180000000
0!
0%
b101 *
0-
02
b101 6
#674190000000
1!
1%
1-
12
#674200000000
0!
0%
b110 *
0-
02
b110 6
#674210000000
1!
1%
1-
12
#674220000000
0!
0%
b111 *
0-
02
b111 6
#674230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#674240000000
0!
0%
b0 *
0-
02
b0 6
#674250000000
1!
1%
1-
12
#674260000000
0!
0%
b1 *
0-
02
b1 6
#674270000000
1!
1%
1-
12
#674280000000
0!
0%
b10 *
0-
02
b10 6
#674290000000
1!
1%
1-
12
#674300000000
0!
0%
b11 *
0-
02
b11 6
#674310000000
1!
1%
1-
12
15
#674320000000
0!
0%
b100 *
0-
02
b100 6
#674330000000
1!
1%
1-
12
#674340000000
0!
0%
b101 *
0-
02
b101 6
#674350000000
1!
1%
1-
12
#674360000000
0!
0%
b110 *
0-
02
b110 6
#674370000000
1!
1%
1-
12
#674380000000
0!
0%
b111 *
0-
02
b111 6
#674390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#674400000000
0!
0%
b0 *
0-
02
b0 6
#674410000000
1!
1%
1-
12
#674420000000
0!
0%
b1 *
0-
02
b1 6
#674430000000
1!
1%
1-
12
#674440000000
0!
0%
b10 *
0-
02
b10 6
#674450000000
1!
1%
1-
12
#674460000000
0!
0%
b11 *
0-
02
b11 6
#674470000000
1!
1%
1-
12
15
#674480000000
0!
0%
b100 *
0-
02
b100 6
#674490000000
1!
1%
1-
12
#674500000000
0!
0%
b101 *
0-
02
b101 6
#674510000000
1!
1%
1-
12
#674520000000
0!
0%
b110 *
0-
02
b110 6
#674530000000
1!
1%
1-
12
#674540000000
0!
0%
b111 *
0-
02
b111 6
#674550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#674560000000
0!
0%
b0 *
0-
02
b0 6
#674570000000
1!
1%
1-
12
#674580000000
0!
0%
b1 *
0-
02
b1 6
#674590000000
1!
1%
1-
12
#674600000000
0!
0%
b10 *
0-
02
b10 6
#674610000000
1!
1%
1-
12
#674620000000
0!
0%
b11 *
0-
02
b11 6
#674630000000
1!
1%
1-
12
15
#674640000000
0!
0%
b100 *
0-
02
b100 6
#674650000000
1!
1%
1-
12
#674660000000
0!
0%
b101 *
0-
02
b101 6
#674670000000
1!
1%
1-
12
#674680000000
0!
0%
b110 *
0-
02
b110 6
#674690000000
1!
1%
1-
12
#674700000000
0!
0%
b111 *
0-
02
b111 6
#674710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#674720000000
0!
0%
b0 *
0-
02
b0 6
#674730000000
1!
1%
1-
12
#674740000000
0!
0%
b1 *
0-
02
b1 6
#674750000000
1!
1%
1-
12
#674760000000
0!
0%
b10 *
0-
02
b10 6
#674770000000
1!
1%
1-
12
#674780000000
0!
0%
b11 *
0-
02
b11 6
#674790000000
1!
1%
1-
12
15
#674800000000
0!
0%
b100 *
0-
02
b100 6
#674810000000
1!
1%
1-
12
#674820000000
0!
0%
b101 *
0-
02
b101 6
#674830000000
1!
1%
1-
12
#674840000000
0!
0%
b110 *
0-
02
b110 6
#674850000000
1!
1%
1-
12
#674860000000
0!
0%
b111 *
0-
02
b111 6
#674870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#674880000000
0!
0%
b0 *
0-
02
b0 6
#674890000000
1!
1%
1-
12
#674900000000
0!
0%
b1 *
0-
02
b1 6
#674910000000
1!
1%
1-
12
#674920000000
0!
0%
b10 *
0-
02
b10 6
#674930000000
1!
1%
1-
12
#674940000000
0!
0%
b11 *
0-
02
b11 6
#674950000000
1!
1%
1-
12
15
#674960000000
0!
0%
b100 *
0-
02
b100 6
#674970000000
1!
1%
1-
12
#674980000000
0!
0%
b101 *
0-
02
b101 6
#674990000000
1!
1%
1-
12
#675000000000
0!
0%
b110 *
0-
02
b110 6
#675010000000
1!
1%
1-
12
#675020000000
0!
0%
b111 *
0-
02
b111 6
#675030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#675040000000
0!
0%
b0 *
0-
02
b0 6
#675050000000
1!
1%
1-
12
#675060000000
0!
0%
b1 *
0-
02
b1 6
#675070000000
1!
1%
1-
12
#675080000000
0!
0%
b10 *
0-
02
b10 6
#675090000000
1!
1%
1-
12
#675100000000
0!
0%
b11 *
0-
02
b11 6
#675110000000
1!
1%
1-
12
15
#675120000000
0!
0%
b100 *
0-
02
b100 6
#675130000000
1!
1%
1-
12
#675140000000
0!
0%
b101 *
0-
02
b101 6
#675150000000
1!
1%
1-
12
#675160000000
0!
0%
b110 *
0-
02
b110 6
#675170000000
1!
1%
1-
12
#675180000000
0!
0%
b111 *
0-
02
b111 6
#675190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#675200000000
0!
0%
b0 *
0-
02
b0 6
#675210000000
1!
1%
1-
12
#675220000000
0!
0%
b1 *
0-
02
b1 6
#675230000000
1!
1%
1-
12
#675240000000
0!
0%
b10 *
0-
02
b10 6
#675250000000
1!
1%
1-
12
#675260000000
0!
0%
b11 *
0-
02
b11 6
#675270000000
1!
1%
1-
12
15
#675280000000
0!
0%
b100 *
0-
02
b100 6
#675290000000
1!
1%
1-
12
#675300000000
0!
0%
b101 *
0-
02
b101 6
#675310000000
1!
1%
1-
12
#675320000000
0!
0%
b110 *
0-
02
b110 6
#675330000000
1!
1%
1-
12
#675340000000
0!
0%
b111 *
0-
02
b111 6
#675350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#675360000000
0!
0%
b0 *
0-
02
b0 6
#675370000000
1!
1%
1-
12
#675380000000
0!
0%
b1 *
0-
02
b1 6
#675390000000
1!
1%
1-
12
#675400000000
0!
0%
b10 *
0-
02
b10 6
#675410000000
1!
1%
1-
12
#675420000000
0!
0%
b11 *
0-
02
b11 6
#675430000000
1!
1%
1-
12
15
#675440000000
0!
0%
b100 *
0-
02
b100 6
#675450000000
1!
1%
1-
12
#675460000000
0!
0%
b101 *
0-
02
b101 6
#675470000000
1!
1%
1-
12
#675480000000
0!
0%
b110 *
0-
02
b110 6
#675490000000
1!
1%
1-
12
#675500000000
0!
0%
b111 *
0-
02
b111 6
#675510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#675520000000
0!
0%
b0 *
0-
02
b0 6
#675530000000
1!
1%
1-
12
#675540000000
0!
0%
b1 *
0-
02
b1 6
#675550000000
1!
1%
1-
12
#675560000000
0!
0%
b10 *
0-
02
b10 6
#675570000000
1!
1%
1-
12
#675580000000
0!
0%
b11 *
0-
02
b11 6
#675590000000
1!
1%
1-
12
15
#675600000000
0!
0%
b100 *
0-
02
b100 6
#675610000000
1!
1%
1-
12
#675620000000
0!
0%
b101 *
0-
02
b101 6
#675630000000
1!
1%
1-
12
#675640000000
0!
0%
b110 *
0-
02
b110 6
#675650000000
1!
1%
1-
12
#675660000000
0!
0%
b111 *
0-
02
b111 6
#675670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#675680000000
0!
0%
b0 *
0-
02
b0 6
#675690000000
1!
1%
1-
12
#675700000000
0!
0%
b1 *
0-
02
b1 6
#675710000000
1!
1%
1-
12
#675720000000
0!
0%
b10 *
0-
02
b10 6
#675730000000
1!
1%
1-
12
#675740000000
0!
0%
b11 *
0-
02
b11 6
#675750000000
1!
1%
1-
12
15
#675760000000
0!
0%
b100 *
0-
02
b100 6
#675770000000
1!
1%
1-
12
#675780000000
0!
0%
b101 *
0-
02
b101 6
#675790000000
1!
1%
1-
12
#675800000000
0!
0%
b110 *
0-
02
b110 6
#675810000000
1!
1%
1-
12
#675820000000
0!
0%
b111 *
0-
02
b111 6
#675830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#675840000000
0!
0%
b0 *
0-
02
b0 6
#675850000000
1!
1%
1-
12
#675860000000
0!
0%
b1 *
0-
02
b1 6
#675870000000
1!
1%
1-
12
#675880000000
0!
0%
b10 *
0-
02
b10 6
#675890000000
1!
1%
1-
12
#675900000000
0!
0%
b11 *
0-
02
b11 6
#675910000000
1!
1%
1-
12
15
#675920000000
0!
0%
b100 *
0-
02
b100 6
#675930000000
1!
1%
1-
12
#675940000000
0!
0%
b101 *
0-
02
b101 6
#675950000000
1!
1%
1-
12
#675960000000
0!
0%
b110 *
0-
02
b110 6
#675970000000
1!
1%
1-
12
#675980000000
0!
0%
b111 *
0-
02
b111 6
#675990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#676000000000
0!
0%
b0 *
0-
02
b0 6
#676010000000
1!
1%
1-
12
#676020000000
0!
0%
b1 *
0-
02
b1 6
#676030000000
1!
1%
1-
12
#676040000000
0!
0%
b10 *
0-
02
b10 6
#676050000000
1!
1%
1-
12
#676060000000
0!
0%
b11 *
0-
02
b11 6
#676070000000
1!
1%
1-
12
15
#676080000000
0!
0%
b100 *
0-
02
b100 6
#676090000000
1!
1%
1-
12
#676100000000
0!
0%
b101 *
0-
02
b101 6
#676110000000
1!
1%
1-
12
#676120000000
0!
0%
b110 *
0-
02
b110 6
#676130000000
1!
1%
1-
12
#676140000000
0!
0%
b111 *
0-
02
b111 6
#676150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#676160000000
0!
0%
b0 *
0-
02
b0 6
#676170000000
1!
1%
1-
12
#676180000000
0!
0%
b1 *
0-
02
b1 6
#676190000000
1!
1%
1-
12
#676200000000
0!
0%
b10 *
0-
02
b10 6
#676210000000
1!
1%
1-
12
#676220000000
0!
0%
b11 *
0-
02
b11 6
#676230000000
1!
1%
1-
12
15
#676240000000
0!
0%
b100 *
0-
02
b100 6
#676250000000
1!
1%
1-
12
#676260000000
0!
0%
b101 *
0-
02
b101 6
#676270000000
1!
1%
1-
12
#676280000000
0!
0%
b110 *
0-
02
b110 6
#676290000000
1!
1%
1-
12
#676300000000
0!
0%
b111 *
0-
02
b111 6
#676310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#676320000000
0!
0%
b0 *
0-
02
b0 6
#676330000000
1!
1%
1-
12
#676340000000
0!
0%
b1 *
0-
02
b1 6
#676350000000
1!
1%
1-
12
#676360000000
0!
0%
b10 *
0-
02
b10 6
#676370000000
1!
1%
1-
12
#676380000000
0!
0%
b11 *
0-
02
b11 6
#676390000000
1!
1%
1-
12
15
#676400000000
0!
0%
b100 *
0-
02
b100 6
#676410000000
1!
1%
1-
12
#676420000000
0!
0%
b101 *
0-
02
b101 6
#676430000000
1!
1%
1-
12
#676440000000
0!
0%
b110 *
0-
02
b110 6
#676450000000
1!
1%
1-
12
#676460000000
0!
0%
b111 *
0-
02
b111 6
#676470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#676480000000
0!
0%
b0 *
0-
02
b0 6
#676490000000
1!
1%
1-
12
#676500000000
0!
0%
b1 *
0-
02
b1 6
#676510000000
1!
1%
1-
12
#676520000000
0!
0%
b10 *
0-
02
b10 6
#676530000000
1!
1%
1-
12
#676540000000
0!
0%
b11 *
0-
02
b11 6
#676550000000
1!
1%
1-
12
15
#676560000000
0!
0%
b100 *
0-
02
b100 6
#676570000000
1!
1%
1-
12
#676580000000
0!
0%
b101 *
0-
02
b101 6
#676590000000
1!
1%
1-
12
#676600000000
0!
0%
b110 *
0-
02
b110 6
#676610000000
1!
1%
1-
12
#676620000000
0!
0%
b111 *
0-
02
b111 6
#676630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#676640000000
0!
0%
b0 *
0-
02
b0 6
#676650000000
1!
1%
1-
12
#676660000000
0!
0%
b1 *
0-
02
b1 6
#676670000000
1!
1%
1-
12
#676680000000
0!
0%
b10 *
0-
02
b10 6
#676690000000
1!
1%
1-
12
#676700000000
0!
0%
b11 *
0-
02
b11 6
#676710000000
1!
1%
1-
12
15
#676720000000
0!
0%
b100 *
0-
02
b100 6
#676730000000
1!
1%
1-
12
#676740000000
0!
0%
b101 *
0-
02
b101 6
#676750000000
1!
1%
1-
12
#676760000000
0!
0%
b110 *
0-
02
b110 6
#676770000000
1!
1%
1-
12
#676780000000
0!
0%
b111 *
0-
02
b111 6
#676790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#676800000000
0!
0%
b0 *
0-
02
b0 6
#676810000000
1!
1%
1-
12
#676820000000
0!
0%
b1 *
0-
02
b1 6
#676830000000
1!
1%
1-
12
#676840000000
0!
0%
b10 *
0-
02
b10 6
#676850000000
1!
1%
1-
12
#676860000000
0!
0%
b11 *
0-
02
b11 6
#676870000000
1!
1%
1-
12
15
#676880000000
0!
0%
b100 *
0-
02
b100 6
#676890000000
1!
1%
1-
12
#676900000000
0!
0%
b101 *
0-
02
b101 6
#676910000000
1!
1%
1-
12
#676920000000
0!
0%
b110 *
0-
02
b110 6
#676930000000
1!
1%
1-
12
#676940000000
0!
0%
b111 *
0-
02
b111 6
#676950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#676960000000
0!
0%
b0 *
0-
02
b0 6
#676970000000
1!
1%
1-
12
#676980000000
0!
0%
b1 *
0-
02
b1 6
#676990000000
1!
1%
1-
12
#677000000000
0!
0%
b10 *
0-
02
b10 6
#677010000000
1!
1%
1-
12
#677020000000
0!
0%
b11 *
0-
02
b11 6
#677030000000
1!
1%
1-
12
15
#677040000000
0!
0%
b100 *
0-
02
b100 6
#677050000000
1!
1%
1-
12
#677060000000
0!
0%
b101 *
0-
02
b101 6
#677070000000
1!
1%
1-
12
#677080000000
0!
0%
b110 *
0-
02
b110 6
#677090000000
1!
1%
1-
12
#677100000000
0!
0%
b111 *
0-
02
b111 6
#677110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#677120000000
0!
0%
b0 *
0-
02
b0 6
#677130000000
1!
1%
1-
12
#677140000000
0!
0%
b1 *
0-
02
b1 6
#677150000000
1!
1%
1-
12
#677160000000
0!
0%
b10 *
0-
02
b10 6
#677170000000
1!
1%
1-
12
#677180000000
0!
0%
b11 *
0-
02
b11 6
#677190000000
1!
1%
1-
12
15
#677200000000
0!
0%
b100 *
0-
02
b100 6
#677210000000
1!
1%
1-
12
#677220000000
0!
0%
b101 *
0-
02
b101 6
#677230000000
1!
1%
1-
12
#677240000000
0!
0%
b110 *
0-
02
b110 6
#677250000000
1!
1%
1-
12
#677260000000
0!
0%
b111 *
0-
02
b111 6
#677270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#677280000000
0!
0%
b0 *
0-
02
b0 6
#677290000000
1!
1%
1-
12
#677300000000
0!
0%
b1 *
0-
02
b1 6
#677310000000
1!
1%
1-
12
#677320000000
0!
0%
b10 *
0-
02
b10 6
#677330000000
1!
1%
1-
12
#677340000000
0!
0%
b11 *
0-
02
b11 6
#677350000000
1!
1%
1-
12
15
#677360000000
0!
0%
b100 *
0-
02
b100 6
#677370000000
1!
1%
1-
12
#677380000000
0!
0%
b101 *
0-
02
b101 6
#677390000000
1!
1%
1-
12
#677400000000
0!
0%
b110 *
0-
02
b110 6
#677410000000
1!
1%
1-
12
#677420000000
0!
0%
b111 *
0-
02
b111 6
#677430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#677440000000
0!
0%
b0 *
0-
02
b0 6
#677450000000
1!
1%
1-
12
#677460000000
0!
0%
b1 *
0-
02
b1 6
#677470000000
1!
1%
1-
12
#677480000000
0!
0%
b10 *
0-
02
b10 6
#677490000000
1!
1%
1-
12
#677500000000
0!
0%
b11 *
0-
02
b11 6
#677510000000
1!
1%
1-
12
15
#677520000000
0!
0%
b100 *
0-
02
b100 6
#677530000000
1!
1%
1-
12
#677540000000
0!
0%
b101 *
0-
02
b101 6
#677550000000
1!
1%
1-
12
#677560000000
0!
0%
b110 *
0-
02
b110 6
#677570000000
1!
1%
1-
12
#677580000000
0!
0%
b111 *
0-
02
b111 6
#677590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#677600000000
0!
0%
b0 *
0-
02
b0 6
#677610000000
1!
1%
1-
12
#677620000000
0!
0%
b1 *
0-
02
b1 6
#677630000000
1!
1%
1-
12
#677640000000
0!
0%
b10 *
0-
02
b10 6
#677650000000
1!
1%
1-
12
#677660000000
0!
0%
b11 *
0-
02
b11 6
#677670000000
1!
1%
1-
12
15
#677680000000
0!
0%
b100 *
0-
02
b100 6
#677690000000
1!
1%
1-
12
#677700000000
0!
0%
b101 *
0-
02
b101 6
#677710000000
1!
1%
1-
12
#677720000000
0!
0%
b110 *
0-
02
b110 6
#677730000000
1!
1%
1-
12
#677740000000
0!
0%
b111 *
0-
02
b111 6
#677750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#677760000000
0!
0%
b0 *
0-
02
b0 6
#677770000000
1!
1%
1-
12
#677780000000
0!
0%
b1 *
0-
02
b1 6
#677790000000
1!
1%
1-
12
#677800000000
0!
0%
b10 *
0-
02
b10 6
#677810000000
1!
1%
1-
12
#677820000000
0!
0%
b11 *
0-
02
b11 6
#677830000000
1!
1%
1-
12
15
#677840000000
0!
0%
b100 *
0-
02
b100 6
#677850000000
1!
1%
1-
12
#677860000000
0!
0%
b101 *
0-
02
b101 6
#677870000000
1!
1%
1-
12
#677880000000
0!
0%
b110 *
0-
02
b110 6
#677890000000
1!
1%
1-
12
#677900000000
0!
0%
b111 *
0-
02
b111 6
#677910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#677920000000
0!
0%
b0 *
0-
02
b0 6
#677930000000
1!
1%
1-
12
#677940000000
0!
0%
b1 *
0-
02
b1 6
#677950000000
1!
1%
1-
12
#677960000000
0!
0%
b10 *
0-
02
b10 6
#677970000000
1!
1%
1-
12
#677980000000
0!
0%
b11 *
0-
02
b11 6
#677990000000
1!
1%
1-
12
15
#678000000000
0!
0%
b100 *
0-
02
b100 6
#678010000000
1!
1%
1-
12
#678020000000
0!
0%
b101 *
0-
02
b101 6
#678030000000
1!
1%
1-
12
#678040000000
0!
0%
b110 *
0-
02
b110 6
#678050000000
1!
1%
1-
12
#678060000000
0!
0%
b111 *
0-
02
b111 6
#678070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#678080000000
0!
0%
b0 *
0-
02
b0 6
#678090000000
1!
1%
1-
12
#678100000000
0!
0%
b1 *
0-
02
b1 6
#678110000000
1!
1%
1-
12
#678120000000
0!
0%
b10 *
0-
02
b10 6
#678130000000
1!
1%
1-
12
#678140000000
0!
0%
b11 *
0-
02
b11 6
#678150000000
1!
1%
1-
12
15
#678160000000
0!
0%
b100 *
0-
02
b100 6
#678170000000
1!
1%
1-
12
#678180000000
0!
0%
b101 *
0-
02
b101 6
#678190000000
1!
1%
1-
12
#678200000000
0!
0%
b110 *
0-
02
b110 6
#678210000000
1!
1%
1-
12
#678220000000
0!
0%
b111 *
0-
02
b111 6
#678230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#678240000000
0!
0%
b0 *
0-
02
b0 6
#678250000000
1!
1%
1-
12
#678260000000
0!
0%
b1 *
0-
02
b1 6
#678270000000
1!
1%
1-
12
#678280000000
0!
0%
b10 *
0-
02
b10 6
#678290000000
1!
1%
1-
12
#678300000000
0!
0%
b11 *
0-
02
b11 6
#678310000000
1!
1%
1-
12
15
#678320000000
0!
0%
b100 *
0-
02
b100 6
#678330000000
1!
1%
1-
12
#678340000000
0!
0%
b101 *
0-
02
b101 6
#678350000000
1!
1%
1-
12
#678360000000
0!
0%
b110 *
0-
02
b110 6
#678370000000
1!
1%
1-
12
#678380000000
0!
0%
b111 *
0-
02
b111 6
#678390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#678400000000
0!
0%
b0 *
0-
02
b0 6
#678410000000
1!
1%
1-
12
#678420000000
0!
0%
b1 *
0-
02
b1 6
#678430000000
1!
1%
1-
12
#678440000000
0!
0%
b10 *
0-
02
b10 6
#678450000000
1!
1%
1-
12
#678460000000
0!
0%
b11 *
0-
02
b11 6
#678470000000
1!
1%
1-
12
15
#678480000000
0!
0%
b100 *
0-
02
b100 6
#678490000000
1!
1%
1-
12
#678500000000
0!
0%
b101 *
0-
02
b101 6
#678510000000
1!
1%
1-
12
#678520000000
0!
0%
b110 *
0-
02
b110 6
#678530000000
1!
1%
1-
12
#678540000000
0!
0%
b111 *
0-
02
b111 6
#678550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#678560000000
0!
0%
b0 *
0-
02
b0 6
#678570000000
1!
1%
1-
12
#678580000000
0!
0%
b1 *
0-
02
b1 6
#678590000000
1!
1%
1-
12
#678600000000
0!
0%
b10 *
0-
02
b10 6
#678610000000
1!
1%
1-
12
#678620000000
0!
0%
b11 *
0-
02
b11 6
#678630000000
1!
1%
1-
12
15
#678640000000
0!
0%
b100 *
0-
02
b100 6
#678650000000
1!
1%
1-
12
#678660000000
0!
0%
b101 *
0-
02
b101 6
#678670000000
1!
1%
1-
12
#678680000000
0!
0%
b110 *
0-
02
b110 6
#678690000000
1!
1%
1-
12
#678700000000
0!
0%
b111 *
0-
02
b111 6
#678710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#678720000000
0!
0%
b0 *
0-
02
b0 6
#678730000000
1!
1%
1-
12
#678740000000
0!
0%
b1 *
0-
02
b1 6
#678750000000
1!
1%
1-
12
#678760000000
0!
0%
b10 *
0-
02
b10 6
#678770000000
1!
1%
1-
12
#678780000000
0!
0%
b11 *
0-
02
b11 6
#678790000000
1!
1%
1-
12
15
#678800000000
0!
0%
b100 *
0-
02
b100 6
#678810000000
1!
1%
1-
12
#678820000000
0!
0%
b101 *
0-
02
b101 6
#678830000000
1!
1%
1-
12
#678840000000
0!
0%
b110 *
0-
02
b110 6
#678850000000
1!
1%
1-
12
#678860000000
0!
0%
b111 *
0-
02
b111 6
#678870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#678880000000
0!
0%
b0 *
0-
02
b0 6
#678890000000
1!
1%
1-
12
#678900000000
0!
0%
b1 *
0-
02
b1 6
#678910000000
1!
1%
1-
12
#678920000000
0!
0%
b10 *
0-
02
b10 6
#678930000000
1!
1%
1-
12
#678940000000
0!
0%
b11 *
0-
02
b11 6
#678950000000
1!
1%
1-
12
15
#678960000000
0!
0%
b100 *
0-
02
b100 6
#678970000000
1!
1%
1-
12
#678980000000
0!
0%
b101 *
0-
02
b101 6
#678990000000
1!
1%
1-
12
#679000000000
0!
0%
b110 *
0-
02
b110 6
#679010000000
1!
1%
1-
12
#679020000000
0!
0%
b111 *
0-
02
b111 6
#679030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#679040000000
0!
0%
b0 *
0-
02
b0 6
#679050000000
1!
1%
1-
12
#679060000000
0!
0%
b1 *
0-
02
b1 6
#679070000000
1!
1%
1-
12
#679080000000
0!
0%
b10 *
0-
02
b10 6
#679090000000
1!
1%
1-
12
#679100000000
0!
0%
b11 *
0-
02
b11 6
#679110000000
1!
1%
1-
12
15
#679120000000
0!
0%
b100 *
0-
02
b100 6
#679130000000
1!
1%
1-
12
#679140000000
0!
0%
b101 *
0-
02
b101 6
#679150000000
1!
1%
1-
12
#679160000000
0!
0%
b110 *
0-
02
b110 6
#679170000000
1!
1%
1-
12
#679180000000
0!
0%
b111 *
0-
02
b111 6
#679190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#679200000000
0!
0%
b0 *
0-
02
b0 6
#679210000000
1!
1%
1-
12
#679220000000
0!
0%
b1 *
0-
02
b1 6
#679230000000
1!
1%
1-
12
#679240000000
0!
0%
b10 *
0-
02
b10 6
#679250000000
1!
1%
1-
12
#679260000000
0!
0%
b11 *
0-
02
b11 6
#679270000000
1!
1%
1-
12
15
#679280000000
0!
0%
b100 *
0-
02
b100 6
#679290000000
1!
1%
1-
12
#679300000000
0!
0%
b101 *
0-
02
b101 6
#679310000000
1!
1%
1-
12
#679320000000
0!
0%
b110 *
0-
02
b110 6
#679330000000
1!
1%
1-
12
#679340000000
0!
0%
b111 *
0-
02
b111 6
#679350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#679360000000
0!
0%
b0 *
0-
02
b0 6
#679370000000
1!
1%
1-
12
#679380000000
0!
0%
b1 *
0-
02
b1 6
#679390000000
1!
1%
1-
12
#679400000000
0!
0%
b10 *
0-
02
b10 6
#679410000000
1!
1%
1-
12
#679420000000
0!
0%
b11 *
0-
02
b11 6
#679430000000
1!
1%
1-
12
15
#679440000000
0!
0%
b100 *
0-
02
b100 6
#679450000000
1!
1%
1-
12
#679460000000
0!
0%
b101 *
0-
02
b101 6
#679470000000
1!
1%
1-
12
#679480000000
0!
0%
b110 *
0-
02
b110 6
#679490000000
1!
1%
1-
12
#679500000000
0!
0%
b111 *
0-
02
b111 6
#679510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#679520000000
0!
0%
b0 *
0-
02
b0 6
#679530000000
1!
1%
1-
12
#679540000000
0!
0%
b1 *
0-
02
b1 6
#679550000000
1!
1%
1-
12
#679560000000
0!
0%
b10 *
0-
02
b10 6
#679570000000
1!
1%
1-
12
#679580000000
0!
0%
b11 *
0-
02
b11 6
#679590000000
1!
1%
1-
12
15
#679600000000
0!
0%
b100 *
0-
02
b100 6
#679610000000
1!
1%
1-
12
#679620000000
0!
0%
b101 *
0-
02
b101 6
#679630000000
1!
1%
1-
12
#679640000000
0!
0%
b110 *
0-
02
b110 6
#679650000000
1!
1%
1-
12
#679660000000
0!
0%
b111 *
0-
02
b111 6
#679670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#679680000000
0!
0%
b0 *
0-
02
b0 6
#679690000000
1!
1%
1-
12
#679700000000
0!
0%
b1 *
0-
02
b1 6
#679710000000
1!
1%
1-
12
#679720000000
0!
0%
b10 *
0-
02
b10 6
#679730000000
1!
1%
1-
12
#679740000000
0!
0%
b11 *
0-
02
b11 6
#679750000000
1!
1%
1-
12
15
#679760000000
0!
0%
b100 *
0-
02
b100 6
#679770000000
1!
1%
1-
12
#679780000000
0!
0%
b101 *
0-
02
b101 6
#679790000000
1!
1%
1-
12
#679800000000
0!
0%
b110 *
0-
02
b110 6
#679810000000
1!
1%
1-
12
#679820000000
0!
0%
b111 *
0-
02
b111 6
#679830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#679840000000
0!
0%
b0 *
0-
02
b0 6
#679850000000
1!
1%
1-
12
#679860000000
0!
0%
b1 *
0-
02
b1 6
#679870000000
1!
1%
1-
12
#679880000000
0!
0%
b10 *
0-
02
b10 6
#679890000000
1!
1%
1-
12
#679900000000
0!
0%
b11 *
0-
02
b11 6
#679910000000
1!
1%
1-
12
15
#679920000000
0!
0%
b100 *
0-
02
b100 6
#679930000000
1!
1%
1-
12
#679940000000
0!
0%
b101 *
0-
02
b101 6
#679950000000
1!
1%
1-
12
#679960000000
0!
0%
b110 *
0-
02
b110 6
#679970000000
1!
1%
1-
12
#679980000000
0!
0%
b111 *
0-
02
b111 6
#679990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#680000000000
0!
0%
b0 *
0-
02
b0 6
#680010000000
1!
1%
1-
12
#680020000000
0!
0%
b1 *
0-
02
b1 6
#680030000000
1!
1%
1-
12
#680040000000
0!
0%
b10 *
0-
02
b10 6
#680050000000
1!
1%
1-
12
#680060000000
0!
0%
b11 *
0-
02
b11 6
#680070000000
1!
1%
1-
12
15
#680080000000
0!
0%
b100 *
0-
02
b100 6
#680090000000
1!
1%
1-
12
#680100000000
0!
0%
b101 *
0-
02
b101 6
#680110000000
1!
1%
1-
12
#680120000000
0!
0%
b110 *
0-
02
b110 6
#680130000000
1!
1%
1-
12
#680140000000
0!
0%
b111 *
0-
02
b111 6
#680150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#680160000000
0!
0%
b0 *
0-
02
b0 6
#680170000000
1!
1%
1-
12
#680180000000
0!
0%
b1 *
0-
02
b1 6
#680190000000
1!
1%
1-
12
#680200000000
0!
0%
b10 *
0-
02
b10 6
#680210000000
1!
1%
1-
12
#680220000000
0!
0%
b11 *
0-
02
b11 6
#680230000000
1!
1%
1-
12
15
#680240000000
0!
0%
b100 *
0-
02
b100 6
#680250000000
1!
1%
1-
12
#680260000000
0!
0%
b101 *
0-
02
b101 6
#680270000000
1!
1%
1-
12
#680280000000
0!
0%
b110 *
0-
02
b110 6
#680290000000
1!
1%
1-
12
#680300000000
0!
0%
b111 *
0-
02
b111 6
#680310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#680320000000
0!
0%
b0 *
0-
02
b0 6
#680330000000
1!
1%
1-
12
#680340000000
0!
0%
b1 *
0-
02
b1 6
#680350000000
1!
1%
1-
12
#680360000000
0!
0%
b10 *
0-
02
b10 6
#680370000000
1!
1%
1-
12
#680380000000
0!
0%
b11 *
0-
02
b11 6
#680390000000
1!
1%
1-
12
15
#680400000000
0!
0%
b100 *
0-
02
b100 6
#680410000000
1!
1%
1-
12
#680420000000
0!
0%
b101 *
0-
02
b101 6
#680430000000
1!
1%
1-
12
#680440000000
0!
0%
b110 *
0-
02
b110 6
#680450000000
1!
1%
1-
12
#680460000000
0!
0%
b111 *
0-
02
b111 6
#680470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#680480000000
0!
0%
b0 *
0-
02
b0 6
#680490000000
1!
1%
1-
12
#680500000000
0!
0%
b1 *
0-
02
b1 6
#680510000000
1!
1%
1-
12
#680520000000
0!
0%
b10 *
0-
02
b10 6
#680530000000
1!
1%
1-
12
#680540000000
0!
0%
b11 *
0-
02
b11 6
#680550000000
1!
1%
1-
12
15
#680560000000
0!
0%
b100 *
0-
02
b100 6
#680570000000
1!
1%
1-
12
#680580000000
0!
0%
b101 *
0-
02
b101 6
#680590000000
1!
1%
1-
12
#680600000000
0!
0%
b110 *
0-
02
b110 6
#680610000000
1!
1%
1-
12
#680620000000
0!
0%
b111 *
0-
02
b111 6
#680630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#680640000000
0!
0%
b0 *
0-
02
b0 6
#680650000000
1!
1%
1-
12
#680660000000
0!
0%
b1 *
0-
02
b1 6
#680670000000
1!
1%
1-
12
#680680000000
0!
0%
b10 *
0-
02
b10 6
#680690000000
1!
1%
1-
12
#680700000000
0!
0%
b11 *
0-
02
b11 6
#680710000000
1!
1%
1-
12
15
#680720000000
0!
0%
b100 *
0-
02
b100 6
#680730000000
1!
1%
1-
12
#680740000000
0!
0%
b101 *
0-
02
b101 6
#680750000000
1!
1%
1-
12
#680760000000
0!
0%
b110 *
0-
02
b110 6
#680770000000
1!
1%
1-
12
#680780000000
0!
0%
b111 *
0-
02
b111 6
#680790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#680800000000
0!
0%
b0 *
0-
02
b0 6
#680810000000
1!
1%
1-
12
#680820000000
0!
0%
b1 *
0-
02
b1 6
#680830000000
1!
1%
1-
12
#680840000000
0!
0%
b10 *
0-
02
b10 6
#680850000000
1!
1%
1-
12
#680860000000
0!
0%
b11 *
0-
02
b11 6
#680870000000
1!
1%
1-
12
15
#680880000000
0!
0%
b100 *
0-
02
b100 6
#680890000000
1!
1%
1-
12
#680900000000
0!
0%
b101 *
0-
02
b101 6
#680910000000
1!
1%
1-
12
#680920000000
0!
0%
b110 *
0-
02
b110 6
#680930000000
1!
1%
1-
12
#680940000000
0!
0%
b111 *
0-
02
b111 6
#680950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#680960000000
0!
0%
b0 *
0-
02
b0 6
#680970000000
1!
1%
1-
12
#680980000000
0!
0%
b1 *
0-
02
b1 6
#680990000000
1!
1%
1-
12
#681000000000
0!
0%
b10 *
0-
02
b10 6
#681010000000
1!
1%
1-
12
#681020000000
0!
0%
b11 *
0-
02
b11 6
#681030000000
1!
1%
1-
12
15
#681040000000
0!
0%
b100 *
0-
02
b100 6
#681050000000
1!
1%
1-
12
#681060000000
0!
0%
b101 *
0-
02
b101 6
#681070000000
1!
1%
1-
12
#681080000000
0!
0%
b110 *
0-
02
b110 6
#681090000000
1!
1%
1-
12
#681100000000
0!
0%
b111 *
0-
02
b111 6
#681110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#681120000000
0!
0%
b0 *
0-
02
b0 6
#681130000000
1!
1%
1-
12
#681140000000
0!
0%
b1 *
0-
02
b1 6
#681150000000
1!
1%
1-
12
#681160000000
0!
0%
b10 *
0-
02
b10 6
#681170000000
1!
1%
1-
12
#681180000000
0!
0%
b11 *
0-
02
b11 6
#681190000000
1!
1%
1-
12
15
#681200000000
0!
0%
b100 *
0-
02
b100 6
#681210000000
1!
1%
1-
12
#681220000000
0!
0%
b101 *
0-
02
b101 6
#681230000000
1!
1%
1-
12
#681240000000
0!
0%
b110 *
0-
02
b110 6
#681250000000
1!
1%
1-
12
#681260000000
0!
0%
b111 *
0-
02
b111 6
#681270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#681280000000
0!
0%
b0 *
0-
02
b0 6
#681290000000
1!
1%
1-
12
#681300000000
0!
0%
b1 *
0-
02
b1 6
#681310000000
1!
1%
1-
12
#681320000000
0!
0%
b10 *
0-
02
b10 6
#681330000000
1!
1%
1-
12
#681340000000
0!
0%
b11 *
0-
02
b11 6
#681350000000
1!
1%
1-
12
15
#681360000000
0!
0%
b100 *
0-
02
b100 6
#681370000000
1!
1%
1-
12
#681380000000
0!
0%
b101 *
0-
02
b101 6
#681390000000
1!
1%
1-
12
#681400000000
0!
0%
b110 *
0-
02
b110 6
#681410000000
1!
1%
1-
12
#681420000000
0!
0%
b111 *
0-
02
b111 6
#681430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#681440000000
0!
0%
b0 *
0-
02
b0 6
#681450000000
1!
1%
1-
12
#681460000000
0!
0%
b1 *
0-
02
b1 6
#681470000000
1!
1%
1-
12
#681480000000
0!
0%
b10 *
0-
02
b10 6
#681490000000
1!
1%
1-
12
#681500000000
0!
0%
b11 *
0-
02
b11 6
#681510000000
1!
1%
1-
12
15
#681520000000
0!
0%
b100 *
0-
02
b100 6
#681530000000
1!
1%
1-
12
#681540000000
0!
0%
b101 *
0-
02
b101 6
#681550000000
1!
1%
1-
12
#681560000000
0!
0%
b110 *
0-
02
b110 6
#681570000000
1!
1%
1-
12
#681580000000
0!
0%
b111 *
0-
02
b111 6
#681590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#681600000000
0!
0%
b0 *
0-
02
b0 6
#681610000000
1!
1%
1-
12
#681620000000
0!
0%
b1 *
0-
02
b1 6
#681630000000
1!
1%
1-
12
#681640000000
0!
0%
b10 *
0-
02
b10 6
#681650000000
1!
1%
1-
12
#681660000000
0!
0%
b11 *
0-
02
b11 6
#681670000000
1!
1%
1-
12
15
#681680000000
0!
0%
b100 *
0-
02
b100 6
#681690000000
1!
1%
1-
12
#681700000000
0!
0%
b101 *
0-
02
b101 6
#681710000000
1!
1%
1-
12
#681720000000
0!
0%
b110 *
0-
02
b110 6
#681730000000
1!
1%
1-
12
#681740000000
0!
0%
b111 *
0-
02
b111 6
#681750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#681760000000
0!
0%
b0 *
0-
02
b0 6
#681770000000
1!
1%
1-
12
#681780000000
0!
0%
b1 *
0-
02
b1 6
#681790000000
1!
1%
1-
12
#681800000000
0!
0%
b10 *
0-
02
b10 6
#681810000000
1!
1%
1-
12
#681820000000
0!
0%
b11 *
0-
02
b11 6
#681830000000
1!
1%
1-
12
15
#681840000000
0!
0%
b100 *
0-
02
b100 6
#681850000000
1!
1%
1-
12
#681860000000
0!
0%
b101 *
0-
02
b101 6
#681870000000
1!
1%
1-
12
#681880000000
0!
0%
b110 *
0-
02
b110 6
#681890000000
1!
1%
1-
12
#681900000000
0!
0%
b111 *
0-
02
b111 6
#681910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#681920000000
0!
0%
b0 *
0-
02
b0 6
#681930000000
1!
1%
1-
12
#681940000000
0!
0%
b1 *
0-
02
b1 6
#681950000000
1!
1%
1-
12
#681960000000
0!
0%
b10 *
0-
02
b10 6
#681970000000
1!
1%
1-
12
#681980000000
0!
0%
b11 *
0-
02
b11 6
#681990000000
1!
1%
1-
12
15
#682000000000
0!
0%
b100 *
0-
02
b100 6
#682010000000
1!
1%
1-
12
#682020000000
0!
0%
b101 *
0-
02
b101 6
#682030000000
1!
1%
1-
12
#682040000000
0!
0%
b110 *
0-
02
b110 6
#682050000000
1!
1%
1-
12
#682060000000
0!
0%
b111 *
0-
02
b111 6
#682070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#682080000000
0!
0%
b0 *
0-
02
b0 6
#682090000000
1!
1%
1-
12
#682100000000
0!
0%
b1 *
0-
02
b1 6
#682110000000
1!
1%
1-
12
#682120000000
0!
0%
b10 *
0-
02
b10 6
#682130000000
1!
1%
1-
12
#682140000000
0!
0%
b11 *
0-
02
b11 6
#682150000000
1!
1%
1-
12
15
#682160000000
0!
0%
b100 *
0-
02
b100 6
#682170000000
1!
1%
1-
12
#682180000000
0!
0%
b101 *
0-
02
b101 6
#682190000000
1!
1%
1-
12
#682200000000
0!
0%
b110 *
0-
02
b110 6
#682210000000
1!
1%
1-
12
#682220000000
0!
0%
b111 *
0-
02
b111 6
#682230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#682240000000
0!
0%
b0 *
0-
02
b0 6
#682250000000
1!
1%
1-
12
#682260000000
0!
0%
b1 *
0-
02
b1 6
#682270000000
1!
1%
1-
12
#682280000000
0!
0%
b10 *
0-
02
b10 6
#682290000000
1!
1%
1-
12
#682300000000
0!
0%
b11 *
0-
02
b11 6
#682310000000
1!
1%
1-
12
15
#682320000000
0!
0%
b100 *
0-
02
b100 6
#682330000000
1!
1%
1-
12
#682340000000
0!
0%
b101 *
0-
02
b101 6
#682350000000
1!
1%
1-
12
#682360000000
0!
0%
b110 *
0-
02
b110 6
#682370000000
1!
1%
1-
12
#682380000000
0!
0%
b111 *
0-
02
b111 6
#682390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#682400000000
0!
0%
b0 *
0-
02
b0 6
#682410000000
1!
1%
1-
12
#682420000000
0!
0%
b1 *
0-
02
b1 6
#682430000000
1!
1%
1-
12
#682440000000
0!
0%
b10 *
0-
02
b10 6
#682450000000
1!
1%
1-
12
#682460000000
0!
0%
b11 *
0-
02
b11 6
#682470000000
1!
1%
1-
12
15
#682480000000
0!
0%
b100 *
0-
02
b100 6
#682490000000
1!
1%
1-
12
#682500000000
0!
0%
b101 *
0-
02
b101 6
#682510000000
1!
1%
1-
12
#682520000000
0!
0%
b110 *
0-
02
b110 6
#682530000000
1!
1%
1-
12
#682540000000
0!
0%
b111 *
0-
02
b111 6
#682550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#682560000000
0!
0%
b0 *
0-
02
b0 6
#682570000000
1!
1%
1-
12
#682580000000
0!
0%
b1 *
0-
02
b1 6
#682590000000
1!
1%
1-
12
#682600000000
0!
0%
b10 *
0-
02
b10 6
#682610000000
1!
1%
1-
12
#682620000000
0!
0%
b11 *
0-
02
b11 6
#682630000000
1!
1%
1-
12
15
#682640000000
0!
0%
b100 *
0-
02
b100 6
#682650000000
1!
1%
1-
12
#682660000000
0!
0%
b101 *
0-
02
b101 6
#682670000000
1!
1%
1-
12
#682680000000
0!
0%
b110 *
0-
02
b110 6
#682690000000
1!
1%
1-
12
#682700000000
0!
0%
b111 *
0-
02
b111 6
#682710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#682720000000
0!
0%
b0 *
0-
02
b0 6
#682730000000
1!
1%
1-
12
#682740000000
0!
0%
b1 *
0-
02
b1 6
#682750000000
1!
1%
1-
12
#682760000000
0!
0%
b10 *
0-
02
b10 6
#682770000000
1!
1%
1-
12
#682780000000
0!
0%
b11 *
0-
02
b11 6
#682790000000
1!
1%
1-
12
15
#682800000000
0!
0%
b100 *
0-
02
b100 6
#682810000000
1!
1%
1-
12
#682820000000
0!
0%
b101 *
0-
02
b101 6
#682830000000
1!
1%
1-
12
#682840000000
0!
0%
b110 *
0-
02
b110 6
#682850000000
1!
1%
1-
12
#682860000000
0!
0%
b111 *
0-
02
b111 6
#682870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#682880000000
0!
0%
b0 *
0-
02
b0 6
#682890000000
1!
1%
1-
12
#682900000000
0!
0%
b1 *
0-
02
b1 6
#682910000000
1!
1%
1-
12
#682920000000
0!
0%
b10 *
0-
02
b10 6
#682930000000
1!
1%
1-
12
#682940000000
0!
0%
b11 *
0-
02
b11 6
#682950000000
1!
1%
1-
12
15
#682960000000
0!
0%
b100 *
0-
02
b100 6
#682970000000
1!
1%
1-
12
#682980000000
0!
0%
b101 *
0-
02
b101 6
#682990000000
1!
1%
1-
12
#683000000000
0!
0%
b110 *
0-
02
b110 6
#683010000000
1!
1%
1-
12
#683020000000
0!
0%
b111 *
0-
02
b111 6
#683030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#683040000000
0!
0%
b0 *
0-
02
b0 6
#683050000000
1!
1%
1-
12
#683060000000
0!
0%
b1 *
0-
02
b1 6
#683070000000
1!
1%
1-
12
#683080000000
0!
0%
b10 *
0-
02
b10 6
#683090000000
1!
1%
1-
12
#683100000000
0!
0%
b11 *
0-
02
b11 6
#683110000000
1!
1%
1-
12
15
#683120000000
0!
0%
b100 *
0-
02
b100 6
#683130000000
1!
1%
1-
12
#683140000000
0!
0%
b101 *
0-
02
b101 6
#683150000000
1!
1%
1-
12
#683160000000
0!
0%
b110 *
0-
02
b110 6
#683170000000
1!
1%
1-
12
#683180000000
0!
0%
b111 *
0-
02
b111 6
#683190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#683200000000
0!
0%
b0 *
0-
02
b0 6
#683210000000
1!
1%
1-
12
#683220000000
0!
0%
b1 *
0-
02
b1 6
#683230000000
1!
1%
1-
12
#683240000000
0!
0%
b10 *
0-
02
b10 6
#683250000000
1!
1%
1-
12
#683260000000
0!
0%
b11 *
0-
02
b11 6
#683270000000
1!
1%
1-
12
15
#683280000000
0!
0%
b100 *
0-
02
b100 6
#683290000000
1!
1%
1-
12
#683300000000
0!
0%
b101 *
0-
02
b101 6
#683310000000
1!
1%
1-
12
#683320000000
0!
0%
b110 *
0-
02
b110 6
#683330000000
1!
1%
1-
12
#683340000000
0!
0%
b111 *
0-
02
b111 6
#683350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#683360000000
0!
0%
b0 *
0-
02
b0 6
#683370000000
1!
1%
1-
12
#683380000000
0!
0%
b1 *
0-
02
b1 6
#683390000000
1!
1%
1-
12
#683400000000
0!
0%
b10 *
0-
02
b10 6
#683410000000
1!
1%
1-
12
#683420000000
0!
0%
b11 *
0-
02
b11 6
#683430000000
1!
1%
1-
12
15
#683440000000
0!
0%
b100 *
0-
02
b100 6
#683450000000
1!
1%
1-
12
#683460000000
0!
0%
b101 *
0-
02
b101 6
#683470000000
1!
1%
1-
12
#683480000000
0!
0%
b110 *
0-
02
b110 6
#683490000000
1!
1%
1-
12
#683500000000
0!
0%
b111 *
0-
02
b111 6
#683510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#683520000000
0!
0%
b0 *
0-
02
b0 6
#683530000000
1!
1%
1-
12
#683540000000
0!
0%
b1 *
0-
02
b1 6
#683550000000
1!
1%
1-
12
#683560000000
0!
0%
b10 *
0-
02
b10 6
#683570000000
1!
1%
1-
12
#683580000000
0!
0%
b11 *
0-
02
b11 6
#683590000000
1!
1%
1-
12
15
#683600000000
0!
0%
b100 *
0-
02
b100 6
#683610000000
1!
1%
1-
12
#683620000000
0!
0%
b101 *
0-
02
b101 6
#683630000000
1!
1%
1-
12
#683640000000
0!
0%
b110 *
0-
02
b110 6
#683650000000
1!
1%
1-
12
#683660000000
0!
0%
b111 *
0-
02
b111 6
#683670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#683680000000
0!
0%
b0 *
0-
02
b0 6
#683690000000
1!
1%
1-
12
#683700000000
0!
0%
b1 *
0-
02
b1 6
#683710000000
1!
1%
1-
12
#683720000000
0!
0%
b10 *
0-
02
b10 6
#683730000000
1!
1%
1-
12
#683740000000
0!
0%
b11 *
0-
02
b11 6
#683750000000
1!
1%
1-
12
15
#683760000000
0!
0%
b100 *
0-
02
b100 6
#683770000000
1!
1%
1-
12
#683780000000
0!
0%
b101 *
0-
02
b101 6
#683790000000
1!
1%
1-
12
#683800000000
0!
0%
b110 *
0-
02
b110 6
#683810000000
1!
1%
1-
12
#683820000000
0!
0%
b111 *
0-
02
b111 6
#683830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#683840000000
0!
0%
b0 *
0-
02
b0 6
#683850000000
1!
1%
1-
12
#683860000000
0!
0%
b1 *
0-
02
b1 6
#683870000000
1!
1%
1-
12
#683880000000
0!
0%
b10 *
0-
02
b10 6
#683890000000
1!
1%
1-
12
#683900000000
0!
0%
b11 *
0-
02
b11 6
#683910000000
1!
1%
1-
12
15
#683920000000
0!
0%
b100 *
0-
02
b100 6
#683930000000
1!
1%
1-
12
#683940000000
0!
0%
b101 *
0-
02
b101 6
#683950000000
1!
1%
1-
12
#683960000000
0!
0%
b110 *
0-
02
b110 6
#683970000000
1!
1%
1-
12
#683980000000
0!
0%
b111 *
0-
02
b111 6
#683990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#684000000000
0!
0%
b0 *
0-
02
b0 6
#684010000000
1!
1%
1-
12
#684020000000
0!
0%
b1 *
0-
02
b1 6
#684030000000
1!
1%
1-
12
#684040000000
0!
0%
b10 *
0-
02
b10 6
#684050000000
1!
1%
1-
12
#684060000000
0!
0%
b11 *
0-
02
b11 6
#684070000000
1!
1%
1-
12
15
#684080000000
0!
0%
b100 *
0-
02
b100 6
#684090000000
1!
1%
1-
12
#684100000000
0!
0%
b101 *
0-
02
b101 6
#684110000000
1!
1%
1-
12
#684120000000
0!
0%
b110 *
0-
02
b110 6
#684130000000
1!
1%
1-
12
#684140000000
0!
0%
b111 *
0-
02
b111 6
#684150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#684160000000
0!
0%
b0 *
0-
02
b0 6
#684170000000
1!
1%
1-
12
#684180000000
0!
0%
b1 *
0-
02
b1 6
#684190000000
1!
1%
1-
12
#684200000000
0!
0%
b10 *
0-
02
b10 6
#684210000000
1!
1%
1-
12
#684220000000
0!
0%
b11 *
0-
02
b11 6
#684230000000
1!
1%
1-
12
15
#684240000000
0!
0%
b100 *
0-
02
b100 6
#684250000000
1!
1%
1-
12
#684260000000
0!
0%
b101 *
0-
02
b101 6
#684270000000
1!
1%
1-
12
#684280000000
0!
0%
b110 *
0-
02
b110 6
#684290000000
1!
1%
1-
12
#684300000000
0!
0%
b111 *
0-
02
b111 6
#684310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#684320000000
0!
0%
b0 *
0-
02
b0 6
#684330000000
1!
1%
1-
12
#684340000000
0!
0%
b1 *
0-
02
b1 6
#684350000000
1!
1%
1-
12
#684360000000
0!
0%
b10 *
0-
02
b10 6
#684370000000
1!
1%
1-
12
#684380000000
0!
0%
b11 *
0-
02
b11 6
#684390000000
1!
1%
1-
12
15
#684400000000
0!
0%
b100 *
0-
02
b100 6
#684410000000
1!
1%
1-
12
#684420000000
0!
0%
b101 *
0-
02
b101 6
#684430000000
1!
1%
1-
12
#684440000000
0!
0%
b110 *
0-
02
b110 6
#684450000000
1!
1%
1-
12
#684460000000
0!
0%
b111 *
0-
02
b111 6
#684470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#684480000000
0!
0%
b0 *
0-
02
b0 6
#684490000000
1!
1%
1-
12
#684500000000
0!
0%
b1 *
0-
02
b1 6
#684510000000
1!
1%
1-
12
#684520000000
0!
0%
b10 *
0-
02
b10 6
#684530000000
1!
1%
1-
12
#684540000000
0!
0%
b11 *
0-
02
b11 6
#684550000000
1!
1%
1-
12
15
#684560000000
0!
0%
b100 *
0-
02
b100 6
#684570000000
1!
1%
1-
12
#684580000000
0!
0%
b101 *
0-
02
b101 6
#684590000000
1!
1%
1-
12
#684600000000
0!
0%
b110 *
0-
02
b110 6
#684610000000
1!
1%
1-
12
#684620000000
0!
0%
b111 *
0-
02
b111 6
#684630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#684640000000
0!
0%
b0 *
0-
02
b0 6
#684650000000
1!
1%
1-
12
#684660000000
0!
0%
b1 *
0-
02
b1 6
#684670000000
1!
1%
1-
12
#684680000000
0!
0%
b10 *
0-
02
b10 6
#684690000000
1!
1%
1-
12
#684700000000
0!
0%
b11 *
0-
02
b11 6
#684710000000
1!
1%
1-
12
15
#684720000000
0!
0%
b100 *
0-
02
b100 6
#684730000000
1!
1%
1-
12
#684740000000
0!
0%
b101 *
0-
02
b101 6
#684750000000
1!
1%
1-
12
#684760000000
0!
0%
b110 *
0-
02
b110 6
#684770000000
1!
1%
1-
12
#684780000000
0!
0%
b111 *
0-
02
b111 6
#684790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#684800000000
0!
0%
b0 *
0-
02
b0 6
#684810000000
1!
1%
1-
12
#684820000000
0!
0%
b1 *
0-
02
b1 6
#684830000000
1!
1%
1-
12
#684840000000
0!
0%
b10 *
0-
02
b10 6
#684850000000
1!
1%
1-
12
#684860000000
0!
0%
b11 *
0-
02
b11 6
#684870000000
1!
1%
1-
12
15
#684880000000
0!
0%
b100 *
0-
02
b100 6
#684890000000
1!
1%
1-
12
#684900000000
0!
0%
b101 *
0-
02
b101 6
#684910000000
1!
1%
1-
12
#684920000000
0!
0%
b110 *
0-
02
b110 6
#684930000000
1!
1%
1-
12
#684940000000
0!
0%
b111 *
0-
02
b111 6
#684950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#684960000000
0!
0%
b0 *
0-
02
b0 6
#684970000000
1!
1%
1-
12
#684980000000
0!
0%
b1 *
0-
02
b1 6
#684990000000
1!
1%
1-
12
#685000000000
0!
0%
b10 *
0-
02
b10 6
#685010000000
1!
1%
1-
12
#685020000000
0!
0%
b11 *
0-
02
b11 6
#685030000000
1!
1%
1-
12
15
#685040000000
0!
0%
b100 *
0-
02
b100 6
#685050000000
1!
1%
1-
12
#685060000000
0!
0%
b101 *
0-
02
b101 6
#685070000000
1!
1%
1-
12
#685080000000
0!
0%
b110 *
0-
02
b110 6
#685090000000
1!
1%
1-
12
#685100000000
0!
0%
b111 *
0-
02
b111 6
#685110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#685120000000
0!
0%
b0 *
0-
02
b0 6
#685130000000
1!
1%
1-
12
#685140000000
0!
0%
b1 *
0-
02
b1 6
#685150000000
1!
1%
1-
12
#685160000000
0!
0%
b10 *
0-
02
b10 6
#685170000000
1!
1%
1-
12
#685180000000
0!
0%
b11 *
0-
02
b11 6
#685190000000
1!
1%
1-
12
15
#685200000000
0!
0%
b100 *
0-
02
b100 6
#685210000000
1!
1%
1-
12
#685220000000
0!
0%
b101 *
0-
02
b101 6
#685230000000
1!
1%
1-
12
#685240000000
0!
0%
b110 *
0-
02
b110 6
#685250000000
1!
1%
1-
12
#685260000000
0!
0%
b111 *
0-
02
b111 6
#685270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#685280000000
0!
0%
b0 *
0-
02
b0 6
#685290000000
1!
1%
1-
12
#685300000000
0!
0%
b1 *
0-
02
b1 6
#685310000000
1!
1%
1-
12
#685320000000
0!
0%
b10 *
0-
02
b10 6
#685330000000
1!
1%
1-
12
#685340000000
0!
0%
b11 *
0-
02
b11 6
#685350000000
1!
1%
1-
12
15
#685360000000
0!
0%
b100 *
0-
02
b100 6
#685370000000
1!
1%
1-
12
#685380000000
0!
0%
b101 *
0-
02
b101 6
#685390000000
1!
1%
1-
12
#685400000000
0!
0%
b110 *
0-
02
b110 6
#685410000000
1!
1%
1-
12
#685420000000
0!
0%
b111 *
0-
02
b111 6
#685430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#685440000000
0!
0%
b0 *
0-
02
b0 6
#685450000000
1!
1%
1-
12
#685460000000
0!
0%
b1 *
0-
02
b1 6
#685470000000
1!
1%
1-
12
#685480000000
0!
0%
b10 *
0-
02
b10 6
#685490000000
1!
1%
1-
12
#685500000000
0!
0%
b11 *
0-
02
b11 6
#685510000000
1!
1%
1-
12
15
#685520000000
0!
0%
b100 *
0-
02
b100 6
#685530000000
1!
1%
1-
12
#685540000000
0!
0%
b101 *
0-
02
b101 6
#685550000000
1!
1%
1-
12
#685560000000
0!
0%
b110 *
0-
02
b110 6
#685570000000
1!
1%
1-
12
#685580000000
0!
0%
b111 *
0-
02
b111 6
#685590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#685600000000
0!
0%
b0 *
0-
02
b0 6
#685610000000
1!
1%
1-
12
#685620000000
0!
0%
b1 *
0-
02
b1 6
#685630000000
1!
1%
1-
12
#685640000000
0!
0%
b10 *
0-
02
b10 6
#685650000000
1!
1%
1-
12
#685660000000
0!
0%
b11 *
0-
02
b11 6
#685670000000
1!
1%
1-
12
15
#685680000000
0!
0%
b100 *
0-
02
b100 6
#685690000000
1!
1%
1-
12
#685700000000
0!
0%
b101 *
0-
02
b101 6
#685710000000
1!
1%
1-
12
#685720000000
0!
0%
b110 *
0-
02
b110 6
#685730000000
1!
1%
1-
12
#685740000000
0!
0%
b111 *
0-
02
b111 6
#685750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#685760000000
0!
0%
b0 *
0-
02
b0 6
#685770000000
1!
1%
1-
12
#685780000000
0!
0%
b1 *
0-
02
b1 6
#685790000000
1!
1%
1-
12
#685800000000
0!
0%
b10 *
0-
02
b10 6
#685810000000
1!
1%
1-
12
#685820000000
0!
0%
b11 *
0-
02
b11 6
#685830000000
1!
1%
1-
12
15
#685840000000
0!
0%
b100 *
0-
02
b100 6
#685850000000
1!
1%
1-
12
#685860000000
0!
0%
b101 *
0-
02
b101 6
#685870000000
1!
1%
1-
12
#685880000000
0!
0%
b110 *
0-
02
b110 6
#685890000000
1!
1%
1-
12
#685900000000
0!
0%
b111 *
0-
02
b111 6
#685910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#685920000000
0!
0%
b0 *
0-
02
b0 6
#685930000000
1!
1%
1-
12
#685940000000
0!
0%
b1 *
0-
02
b1 6
#685950000000
1!
1%
1-
12
#685960000000
0!
0%
b10 *
0-
02
b10 6
#685970000000
1!
1%
1-
12
#685980000000
0!
0%
b11 *
0-
02
b11 6
#685990000000
1!
1%
1-
12
15
#686000000000
0!
0%
b100 *
0-
02
b100 6
#686010000000
1!
1%
1-
12
#686020000000
0!
0%
b101 *
0-
02
b101 6
#686030000000
1!
1%
1-
12
#686040000000
0!
0%
b110 *
0-
02
b110 6
#686050000000
1!
1%
1-
12
#686060000000
0!
0%
b111 *
0-
02
b111 6
#686070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#686080000000
0!
0%
b0 *
0-
02
b0 6
#686090000000
1!
1%
1-
12
#686100000000
0!
0%
b1 *
0-
02
b1 6
#686110000000
1!
1%
1-
12
#686120000000
0!
0%
b10 *
0-
02
b10 6
#686130000000
1!
1%
1-
12
#686140000000
0!
0%
b11 *
0-
02
b11 6
#686150000000
1!
1%
1-
12
15
#686160000000
0!
0%
b100 *
0-
02
b100 6
#686170000000
1!
1%
1-
12
#686180000000
0!
0%
b101 *
0-
02
b101 6
#686190000000
1!
1%
1-
12
#686200000000
0!
0%
b110 *
0-
02
b110 6
#686210000000
1!
1%
1-
12
#686220000000
0!
0%
b111 *
0-
02
b111 6
#686230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#686240000000
0!
0%
b0 *
0-
02
b0 6
#686250000000
1!
1%
1-
12
#686260000000
0!
0%
b1 *
0-
02
b1 6
#686270000000
1!
1%
1-
12
#686280000000
0!
0%
b10 *
0-
02
b10 6
#686290000000
1!
1%
1-
12
#686300000000
0!
0%
b11 *
0-
02
b11 6
#686310000000
1!
1%
1-
12
15
#686320000000
0!
0%
b100 *
0-
02
b100 6
#686330000000
1!
1%
1-
12
#686340000000
0!
0%
b101 *
0-
02
b101 6
#686350000000
1!
1%
1-
12
#686360000000
0!
0%
b110 *
0-
02
b110 6
#686370000000
1!
1%
1-
12
#686380000000
0!
0%
b111 *
0-
02
b111 6
#686390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#686400000000
0!
0%
b0 *
0-
02
b0 6
#686410000000
1!
1%
1-
12
#686420000000
0!
0%
b1 *
0-
02
b1 6
#686430000000
1!
1%
1-
12
#686440000000
0!
0%
b10 *
0-
02
b10 6
#686450000000
1!
1%
1-
12
#686460000000
0!
0%
b11 *
0-
02
b11 6
#686470000000
1!
1%
1-
12
15
#686480000000
0!
0%
b100 *
0-
02
b100 6
#686490000000
1!
1%
1-
12
#686500000000
0!
0%
b101 *
0-
02
b101 6
#686510000000
1!
1%
1-
12
#686520000000
0!
0%
b110 *
0-
02
b110 6
#686530000000
1!
1%
1-
12
#686540000000
0!
0%
b111 *
0-
02
b111 6
#686550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#686560000000
0!
0%
b0 *
0-
02
b0 6
#686570000000
1!
1%
1-
12
#686580000000
0!
0%
b1 *
0-
02
b1 6
#686590000000
1!
1%
1-
12
#686600000000
0!
0%
b10 *
0-
02
b10 6
#686610000000
1!
1%
1-
12
#686620000000
0!
0%
b11 *
0-
02
b11 6
#686630000000
1!
1%
1-
12
15
#686640000000
0!
0%
b100 *
0-
02
b100 6
#686650000000
1!
1%
1-
12
#686660000000
0!
0%
b101 *
0-
02
b101 6
#686670000000
1!
1%
1-
12
#686680000000
0!
0%
b110 *
0-
02
b110 6
#686690000000
1!
1%
1-
12
#686700000000
0!
0%
b111 *
0-
02
b111 6
#686710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#686720000000
0!
0%
b0 *
0-
02
b0 6
#686730000000
1!
1%
1-
12
#686740000000
0!
0%
b1 *
0-
02
b1 6
#686750000000
1!
1%
1-
12
#686760000000
0!
0%
b10 *
0-
02
b10 6
#686770000000
1!
1%
1-
12
#686780000000
0!
0%
b11 *
0-
02
b11 6
#686790000000
1!
1%
1-
12
15
#686800000000
0!
0%
b100 *
0-
02
b100 6
#686810000000
1!
1%
1-
12
#686820000000
0!
0%
b101 *
0-
02
b101 6
#686830000000
1!
1%
1-
12
#686840000000
0!
0%
b110 *
0-
02
b110 6
#686850000000
1!
1%
1-
12
#686860000000
0!
0%
b111 *
0-
02
b111 6
#686870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#686880000000
0!
0%
b0 *
0-
02
b0 6
#686890000000
1!
1%
1-
12
#686900000000
0!
0%
b1 *
0-
02
b1 6
#686910000000
1!
1%
1-
12
#686920000000
0!
0%
b10 *
0-
02
b10 6
#686930000000
1!
1%
1-
12
#686940000000
0!
0%
b11 *
0-
02
b11 6
#686950000000
1!
1%
1-
12
15
#686960000000
0!
0%
b100 *
0-
02
b100 6
#686970000000
1!
1%
1-
12
#686980000000
0!
0%
b101 *
0-
02
b101 6
#686990000000
1!
1%
1-
12
#687000000000
0!
0%
b110 *
0-
02
b110 6
#687010000000
1!
1%
1-
12
#687020000000
0!
0%
b111 *
0-
02
b111 6
#687030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#687040000000
0!
0%
b0 *
0-
02
b0 6
#687050000000
1!
1%
1-
12
#687060000000
0!
0%
b1 *
0-
02
b1 6
#687070000000
1!
1%
1-
12
#687080000000
0!
0%
b10 *
0-
02
b10 6
#687090000000
1!
1%
1-
12
#687100000000
0!
0%
b11 *
0-
02
b11 6
#687110000000
1!
1%
1-
12
15
#687120000000
0!
0%
b100 *
0-
02
b100 6
#687130000000
1!
1%
1-
12
#687140000000
0!
0%
b101 *
0-
02
b101 6
#687150000000
1!
1%
1-
12
#687160000000
0!
0%
b110 *
0-
02
b110 6
#687170000000
1!
1%
1-
12
#687180000000
0!
0%
b111 *
0-
02
b111 6
#687190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#687200000000
0!
0%
b0 *
0-
02
b0 6
#687210000000
1!
1%
1-
12
#687220000000
0!
0%
b1 *
0-
02
b1 6
#687230000000
1!
1%
1-
12
#687240000000
0!
0%
b10 *
0-
02
b10 6
#687250000000
1!
1%
1-
12
#687260000000
0!
0%
b11 *
0-
02
b11 6
#687270000000
1!
1%
1-
12
15
#687280000000
0!
0%
b100 *
0-
02
b100 6
#687290000000
1!
1%
1-
12
#687300000000
0!
0%
b101 *
0-
02
b101 6
#687310000000
1!
1%
1-
12
#687320000000
0!
0%
b110 *
0-
02
b110 6
#687330000000
1!
1%
1-
12
#687340000000
0!
0%
b111 *
0-
02
b111 6
#687350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#687360000000
0!
0%
b0 *
0-
02
b0 6
#687370000000
1!
1%
1-
12
#687380000000
0!
0%
b1 *
0-
02
b1 6
#687390000000
1!
1%
1-
12
#687400000000
0!
0%
b10 *
0-
02
b10 6
#687410000000
1!
1%
1-
12
#687420000000
0!
0%
b11 *
0-
02
b11 6
#687430000000
1!
1%
1-
12
15
#687440000000
0!
0%
b100 *
0-
02
b100 6
#687450000000
1!
1%
1-
12
#687460000000
0!
0%
b101 *
0-
02
b101 6
#687470000000
1!
1%
1-
12
#687480000000
0!
0%
b110 *
0-
02
b110 6
#687490000000
1!
1%
1-
12
#687500000000
0!
0%
b111 *
0-
02
b111 6
#687510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#687520000000
0!
0%
b0 *
0-
02
b0 6
#687530000000
1!
1%
1-
12
#687540000000
0!
0%
b1 *
0-
02
b1 6
#687550000000
1!
1%
1-
12
#687560000000
0!
0%
b10 *
0-
02
b10 6
#687570000000
1!
1%
1-
12
#687580000000
0!
0%
b11 *
0-
02
b11 6
#687590000000
1!
1%
1-
12
15
#687600000000
0!
0%
b100 *
0-
02
b100 6
#687610000000
1!
1%
1-
12
#687620000000
0!
0%
b101 *
0-
02
b101 6
#687630000000
1!
1%
1-
12
#687640000000
0!
0%
b110 *
0-
02
b110 6
#687650000000
1!
1%
1-
12
#687660000000
0!
0%
b111 *
0-
02
b111 6
#687670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#687680000000
0!
0%
b0 *
0-
02
b0 6
#687690000000
1!
1%
1-
12
#687700000000
0!
0%
b1 *
0-
02
b1 6
#687710000000
1!
1%
1-
12
#687720000000
0!
0%
b10 *
0-
02
b10 6
#687730000000
1!
1%
1-
12
#687740000000
0!
0%
b11 *
0-
02
b11 6
#687750000000
1!
1%
1-
12
15
#687760000000
0!
0%
b100 *
0-
02
b100 6
#687770000000
1!
1%
1-
12
#687780000000
0!
0%
b101 *
0-
02
b101 6
#687790000000
1!
1%
1-
12
#687800000000
0!
0%
b110 *
0-
02
b110 6
#687810000000
1!
1%
1-
12
#687820000000
0!
0%
b111 *
0-
02
b111 6
#687830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#687840000000
0!
0%
b0 *
0-
02
b0 6
#687850000000
1!
1%
1-
12
#687860000000
0!
0%
b1 *
0-
02
b1 6
#687870000000
1!
1%
1-
12
#687880000000
0!
0%
b10 *
0-
02
b10 6
#687890000000
1!
1%
1-
12
#687900000000
0!
0%
b11 *
0-
02
b11 6
#687910000000
1!
1%
1-
12
15
#687920000000
0!
0%
b100 *
0-
02
b100 6
#687930000000
1!
1%
1-
12
#687940000000
0!
0%
b101 *
0-
02
b101 6
#687950000000
1!
1%
1-
12
#687960000000
0!
0%
b110 *
0-
02
b110 6
#687970000000
1!
1%
1-
12
#687980000000
0!
0%
b111 *
0-
02
b111 6
#687990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#688000000000
0!
0%
b0 *
0-
02
b0 6
#688010000000
1!
1%
1-
12
#688020000000
0!
0%
b1 *
0-
02
b1 6
#688030000000
1!
1%
1-
12
#688040000000
0!
0%
b10 *
0-
02
b10 6
#688050000000
1!
1%
1-
12
#688060000000
0!
0%
b11 *
0-
02
b11 6
#688070000000
1!
1%
1-
12
15
#688080000000
0!
0%
b100 *
0-
02
b100 6
#688090000000
1!
1%
1-
12
#688100000000
0!
0%
b101 *
0-
02
b101 6
#688110000000
1!
1%
1-
12
#688120000000
0!
0%
b110 *
0-
02
b110 6
#688130000000
1!
1%
1-
12
#688140000000
0!
0%
b111 *
0-
02
b111 6
#688150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#688160000000
0!
0%
b0 *
0-
02
b0 6
#688170000000
1!
1%
1-
12
#688180000000
0!
0%
b1 *
0-
02
b1 6
#688190000000
1!
1%
1-
12
#688200000000
0!
0%
b10 *
0-
02
b10 6
#688210000000
1!
1%
1-
12
#688220000000
0!
0%
b11 *
0-
02
b11 6
#688230000000
1!
1%
1-
12
15
#688240000000
0!
0%
b100 *
0-
02
b100 6
#688250000000
1!
1%
1-
12
#688260000000
0!
0%
b101 *
0-
02
b101 6
#688270000000
1!
1%
1-
12
#688280000000
0!
0%
b110 *
0-
02
b110 6
#688290000000
1!
1%
1-
12
#688300000000
0!
0%
b111 *
0-
02
b111 6
#688310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#688320000000
0!
0%
b0 *
0-
02
b0 6
#688330000000
1!
1%
1-
12
#688340000000
0!
0%
b1 *
0-
02
b1 6
#688350000000
1!
1%
1-
12
#688360000000
0!
0%
b10 *
0-
02
b10 6
#688370000000
1!
1%
1-
12
#688380000000
0!
0%
b11 *
0-
02
b11 6
#688390000000
1!
1%
1-
12
15
#688400000000
0!
0%
b100 *
0-
02
b100 6
#688410000000
1!
1%
1-
12
#688420000000
0!
0%
b101 *
0-
02
b101 6
#688430000000
1!
1%
1-
12
#688440000000
0!
0%
b110 *
0-
02
b110 6
#688450000000
1!
1%
1-
12
#688460000000
0!
0%
b111 *
0-
02
b111 6
#688470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#688480000000
0!
0%
b0 *
0-
02
b0 6
#688490000000
1!
1%
1-
12
#688500000000
0!
0%
b1 *
0-
02
b1 6
#688510000000
1!
1%
1-
12
#688520000000
0!
0%
b10 *
0-
02
b10 6
#688530000000
1!
1%
1-
12
#688540000000
0!
0%
b11 *
0-
02
b11 6
#688550000000
1!
1%
1-
12
15
#688560000000
0!
0%
b100 *
0-
02
b100 6
#688570000000
1!
1%
1-
12
#688580000000
0!
0%
b101 *
0-
02
b101 6
#688590000000
1!
1%
1-
12
#688600000000
0!
0%
b110 *
0-
02
b110 6
#688610000000
1!
1%
1-
12
#688620000000
0!
0%
b111 *
0-
02
b111 6
#688630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#688640000000
0!
0%
b0 *
0-
02
b0 6
#688650000000
1!
1%
1-
12
#688660000000
0!
0%
b1 *
0-
02
b1 6
#688670000000
1!
1%
1-
12
#688680000000
0!
0%
b10 *
0-
02
b10 6
#688690000000
1!
1%
1-
12
#688700000000
0!
0%
b11 *
0-
02
b11 6
#688710000000
1!
1%
1-
12
15
#688720000000
0!
0%
b100 *
0-
02
b100 6
#688730000000
1!
1%
1-
12
#688740000000
0!
0%
b101 *
0-
02
b101 6
#688750000000
1!
1%
1-
12
#688760000000
0!
0%
b110 *
0-
02
b110 6
#688770000000
1!
1%
1-
12
#688780000000
0!
0%
b111 *
0-
02
b111 6
#688790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#688800000000
0!
0%
b0 *
0-
02
b0 6
#688810000000
1!
1%
1-
12
#688820000000
0!
0%
b1 *
0-
02
b1 6
#688830000000
1!
1%
1-
12
#688840000000
0!
0%
b10 *
0-
02
b10 6
#688850000000
1!
1%
1-
12
#688860000000
0!
0%
b11 *
0-
02
b11 6
#688870000000
1!
1%
1-
12
15
#688880000000
0!
0%
b100 *
0-
02
b100 6
#688890000000
1!
1%
1-
12
#688900000000
0!
0%
b101 *
0-
02
b101 6
#688910000000
1!
1%
1-
12
#688920000000
0!
0%
b110 *
0-
02
b110 6
#688930000000
1!
1%
1-
12
#688940000000
0!
0%
b111 *
0-
02
b111 6
#688950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#688960000000
0!
0%
b0 *
0-
02
b0 6
#688970000000
1!
1%
1-
12
#688980000000
0!
0%
b1 *
0-
02
b1 6
#688990000000
1!
1%
1-
12
#689000000000
0!
0%
b10 *
0-
02
b10 6
#689010000000
1!
1%
1-
12
#689020000000
0!
0%
b11 *
0-
02
b11 6
#689030000000
1!
1%
1-
12
15
#689040000000
0!
0%
b100 *
0-
02
b100 6
#689050000000
1!
1%
1-
12
#689060000000
0!
0%
b101 *
0-
02
b101 6
#689070000000
1!
1%
1-
12
#689080000000
0!
0%
b110 *
0-
02
b110 6
#689090000000
1!
1%
1-
12
#689100000000
0!
0%
b111 *
0-
02
b111 6
#689110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#689120000000
0!
0%
b0 *
0-
02
b0 6
#689130000000
1!
1%
1-
12
#689140000000
0!
0%
b1 *
0-
02
b1 6
#689150000000
1!
1%
1-
12
#689160000000
0!
0%
b10 *
0-
02
b10 6
#689170000000
1!
1%
1-
12
#689180000000
0!
0%
b11 *
0-
02
b11 6
#689190000000
1!
1%
1-
12
15
#689200000000
0!
0%
b100 *
0-
02
b100 6
#689210000000
1!
1%
1-
12
#689220000000
0!
0%
b101 *
0-
02
b101 6
#689230000000
1!
1%
1-
12
#689240000000
0!
0%
b110 *
0-
02
b110 6
#689250000000
1!
1%
1-
12
#689260000000
0!
0%
b111 *
0-
02
b111 6
#689270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#689280000000
0!
0%
b0 *
0-
02
b0 6
#689290000000
1!
1%
1-
12
#689300000000
0!
0%
b1 *
0-
02
b1 6
#689310000000
1!
1%
1-
12
#689320000000
0!
0%
b10 *
0-
02
b10 6
#689330000000
1!
1%
1-
12
#689340000000
0!
0%
b11 *
0-
02
b11 6
#689350000000
1!
1%
1-
12
15
#689360000000
0!
0%
b100 *
0-
02
b100 6
#689370000000
1!
1%
1-
12
#689380000000
0!
0%
b101 *
0-
02
b101 6
#689390000000
1!
1%
1-
12
#689400000000
0!
0%
b110 *
0-
02
b110 6
#689410000000
1!
1%
1-
12
#689420000000
0!
0%
b111 *
0-
02
b111 6
#689430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#689440000000
0!
0%
b0 *
0-
02
b0 6
#689450000000
1!
1%
1-
12
#689460000000
0!
0%
b1 *
0-
02
b1 6
#689470000000
1!
1%
1-
12
#689480000000
0!
0%
b10 *
0-
02
b10 6
#689490000000
1!
1%
1-
12
#689500000000
0!
0%
b11 *
0-
02
b11 6
#689510000000
1!
1%
1-
12
15
#689520000000
0!
0%
b100 *
0-
02
b100 6
#689530000000
1!
1%
1-
12
#689540000000
0!
0%
b101 *
0-
02
b101 6
#689550000000
1!
1%
1-
12
#689560000000
0!
0%
b110 *
0-
02
b110 6
#689570000000
1!
1%
1-
12
#689580000000
0!
0%
b111 *
0-
02
b111 6
#689590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#689600000000
0!
0%
b0 *
0-
02
b0 6
#689610000000
1!
1%
1-
12
#689620000000
0!
0%
b1 *
0-
02
b1 6
#689630000000
1!
1%
1-
12
#689640000000
0!
0%
b10 *
0-
02
b10 6
#689650000000
1!
1%
1-
12
#689660000000
0!
0%
b11 *
0-
02
b11 6
#689670000000
1!
1%
1-
12
15
#689680000000
0!
0%
b100 *
0-
02
b100 6
#689690000000
1!
1%
1-
12
#689700000000
0!
0%
b101 *
0-
02
b101 6
#689710000000
1!
1%
1-
12
#689720000000
0!
0%
b110 *
0-
02
b110 6
#689730000000
1!
1%
1-
12
#689740000000
0!
0%
b111 *
0-
02
b111 6
#689750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#689760000000
0!
0%
b0 *
0-
02
b0 6
#689770000000
1!
1%
1-
12
#689780000000
0!
0%
b1 *
0-
02
b1 6
#689790000000
1!
1%
1-
12
#689800000000
0!
0%
b10 *
0-
02
b10 6
#689810000000
1!
1%
1-
12
#689820000000
0!
0%
b11 *
0-
02
b11 6
#689830000000
1!
1%
1-
12
15
#689840000000
0!
0%
b100 *
0-
02
b100 6
#689850000000
1!
1%
1-
12
#689860000000
0!
0%
b101 *
0-
02
b101 6
#689870000000
1!
1%
1-
12
#689880000000
0!
0%
b110 *
0-
02
b110 6
#689890000000
1!
1%
1-
12
#689900000000
0!
0%
b111 *
0-
02
b111 6
#689910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#689920000000
0!
0%
b0 *
0-
02
b0 6
#689930000000
1!
1%
1-
12
#689940000000
0!
0%
b1 *
0-
02
b1 6
#689950000000
1!
1%
1-
12
#689960000000
0!
0%
b10 *
0-
02
b10 6
#689970000000
1!
1%
1-
12
#689980000000
0!
0%
b11 *
0-
02
b11 6
#689990000000
1!
1%
1-
12
15
#690000000000
0!
0%
b100 *
0-
02
b100 6
#690010000000
1!
1%
1-
12
#690020000000
0!
0%
b101 *
0-
02
b101 6
#690030000000
1!
1%
1-
12
#690040000000
0!
0%
b110 *
0-
02
b110 6
#690050000000
1!
1%
1-
12
#690060000000
0!
0%
b111 *
0-
02
b111 6
#690070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#690080000000
0!
0%
b0 *
0-
02
b0 6
#690090000000
1!
1%
1-
12
#690100000000
0!
0%
b1 *
0-
02
b1 6
#690110000000
1!
1%
1-
12
#690120000000
0!
0%
b10 *
0-
02
b10 6
#690130000000
1!
1%
1-
12
#690140000000
0!
0%
b11 *
0-
02
b11 6
#690150000000
1!
1%
1-
12
15
#690160000000
0!
0%
b100 *
0-
02
b100 6
#690170000000
1!
1%
1-
12
#690180000000
0!
0%
b101 *
0-
02
b101 6
#690190000000
1!
1%
1-
12
#690200000000
0!
0%
b110 *
0-
02
b110 6
#690210000000
1!
1%
1-
12
#690220000000
0!
0%
b111 *
0-
02
b111 6
#690230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#690240000000
0!
0%
b0 *
0-
02
b0 6
#690250000000
1!
1%
1-
12
#690260000000
0!
0%
b1 *
0-
02
b1 6
#690270000000
1!
1%
1-
12
#690280000000
0!
0%
b10 *
0-
02
b10 6
#690290000000
1!
1%
1-
12
#690300000000
0!
0%
b11 *
0-
02
b11 6
#690310000000
1!
1%
1-
12
15
#690320000000
0!
0%
b100 *
0-
02
b100 6
#690330000000
1!
1%
1-
12
#690340000000
0!
0%
b101 *
0-
02
b101 6
#690350000000
1!
1%
1-
12
#690360000000
0!
0%
b110 *
0-
02
b110 6
#690370000000
1!
1%
1-
12
#690380000000
0!
0%
b111 *
0-
02
b111 6
#690390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#690400000000
0!
0%
b0 *
0-
02
b0 6
#690410000000
1!
1%
1-
12
#690420000000
0!
0%
b1 *
0-
02
b1 6
#690430000000
1!
1%
1-
12
#690440000000
0!
0%
b10 *
0-
02
b10 6
#690450000000
1!
1%
1-
12
#690460000000
0!
0%
b11 *
0-
02
b11 6
#690470000000
1!
1%
1-
12
15
#690480000000
0!
0%
b100 *
0-
02
b100 6
#690490000000
1!
1%
1-
12
#690500000000
0!
0%
b101 *
0-
02
b101 6
#690510000000
1!
1%
1-
12
#690520000000
0!
0%
b110 *
0-
02
b110 6
#690530000000
1!
1%
1-
12
#690540000000
0!
0%
b111 *
0-
02
b111 6
#690550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#690560000000
0!
0%
b0 *
0-
02
b0 6
#690570000000
1!
1%
1-
12
#690580000000
0!
0%
b1 *
0-
02
b1 6
#690590000000
1!
1%
1-
12
#690600000000
0!
0%
b10 *
0-
02
b10 6
#690610000000
1!
1%
1-
12
#690620000000
0!
0%
b11 *
0-
02
b11 6
#690630000000
1!
1%
1-
12
15
#690640000000
0!
0%
b100 *
0-
02
b100 6
#690650000000
1!
1%
1-
12
#690660000000
0!
0%
b101 *
0-
02
b101 6
#690670000000
1!
1%
1-
12
#690680000000
0!
0%
b110 *
0-
02
b110 6
#690690000000
1!
1%
1-
12
#690700000000
0!
0%
b111 *
0-
02
b111 6
#690710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#690720000000
0!
0%
b0 *
0-
02
b0 6
#690730000000
1!
1%
1-
12
#690740000000
0!
0%
b1 *
0-
02
b1 6
#690750000000
1!
1%
1-
12
#690760000000
0!
0%
b10 *
0-
02
b10 6
#690770000000
1!
1%
1-
12
#690780000000
0!
0%
b11 *
0-
02
b11 6
#690790000000
1!
1%
1-
12
15
#690800000000
0!
0%
b100 *
0-
02
b100 6
#690810000000
1!
1%
1-
12
#690820000000
0!
0%
b101 *
0-
02
b101 6
#690830000000
1!
1%
1-
12
#690840000000
0!
0%
b110 *
0-
02
b110 6
#690850000000
1!
1%
1-
12
#690860000000
0!
0%
b111 *
0-
02
b111 6
#690870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#690880000000
0!
0%
b0 *
0-
02
b0 6
#690890000000
1!
1%
1-
12
#690900000000
0!
0%
b1 *
0-
02
b1 6
#690910000000
1!
1%
1-
12
#690920000000
0!
0%
b10 *
0-
02
b10 6
#690930000000
1!
1%
1-
12
#690940000000
0!
0%
b11 *
0-
02
b11 6
#690950000000
1!
1%
1-
12
15
#690960000000
0!
0%
b100 *
0-
02
b100 6
#690970000000
1!
1%
1-
12
#690980000000
0!
0%
b101 *
0-
02
b101 6
#690990000000
1!
1%
1-
12
#691000000000
0!
0%
b110 *
0-
02
b110 6
#691010000000
1!
1%
1-
12
#691020000000
0!
0%
b111 *
0-
02
b111 6
#691030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#691040000000
0!
0%
b0 *
0-
02
b0 6
#691050000000
1!
1%
1-
12
#691060000000
0!
0%
b1 *
0-
02
b1 6
#691070000000
1!
1%
1-
12
#691080000000
0!
0%
b10 *
0-
02
b10 6
#691090000000
1!
1%
1-
12
#691100000000
0!
0%
b11 *
0-
02
b11 6
#691110000000
1!
1%
1-
12
15
#691120000000
0!
0%
b100 *
0-
02
b100 6
#691130000000
1!
1%
1-
12
#691140000000
0!
0%
b101 *
0-
02
b101 6
#691150000000
1!
1%
1-
12
#691160000000
0!
0%
b110 *
0-
02
b110 6
#691170000000
1!
1%
1-
12
#691180000000
0!
0%
b111 *
0-
02
b111 6
#691190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#691200000000
0!
0%
b0 *
0-
02
b0 6
#691210000000
1!
1%
1-
12
#691220000000
0!
0%
b1 *
0-
02
b1 6
#691230000000
1!
1%
1-
12
#691240000000
0!
0%
b10 *
0-
02
b10 6
#691250000000
1!
1%
1-
12
#691260000000
0!
0%
b11 *
0-
02
b11 6
#691270000000
1!
1%
1-
12
15
#691280000000
0!
0%
b100 *
0-
02
b100 6
#691290000000
1!
1%
1-
12
#691300000000
0!
0%
b101 *
0-
02
b101 6
#691310000000
1!
1%
1-
12
#691320000000
0!
0%
b110 *
0-
02
b110 6
#691330000000
1!
1%
1-
12
#691340000000
0!
0%
b111 *
0-
02
b111 6
#691350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#691360000000
0!
0%
b0 *
0-
02
b0 6
#691370000000
1!
1%
1-
12
#691380000000
0!
0%
b1 *
0-
02
b1 6
#691390000000
1!
1%
1-
12
#691400000000
0!
0%
b10 *
0-
02
b10 6
#691410000000
1!
1%
1-
12
#691420000000
0!
0%
b11 *
0-
02
b11 6
#691430000000
1!
1%
1-
12
15
#691440000000
0!
0%
b100 *
0-
02
b100 6
#691450000000
1!
1%
1-
12
#691460000000
0!
0%
b101 *
0-
02
b101 6
#691470000000
1!
1%
1-
12
#691480000000
0!
0%
b110 *
0-
02
b110 6
#691490000000
1!
1%
1-
12
#691500000000
0!
0%
b111 *
0-
02
b111 6
#691510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#691520000000
0!
0%
b0 *
0-
02
b0 6
#691530000000
1!
1%
1-
12
#691540000000
0!
0%
b1 *
0-
02
b1 6
#691550000000
1!
1%
1-
12
#691560000000
0!
0%
b10 *
0-
02
b10 6
#691570000000
1!
1%
1-
12
#691580000000
0!
0%
b11 *
0-
02
b11 6
#691590000000
1!
1%
1-
12
15
#691600000000
0!
0%
b100 *
0-
02
b100 6
#691610000000
1!
1%
1-
12
#691620000000
0!
0%
b101 *
0-
02
b101 6
#691630000000
1!
1%
1-
12
#691640000000
0!
0%
b110 *
0-
02
b110 6
#691650000000
1!
1%
1-
12
#691660000000
0!
0%
b111 *
0-
02
b111 6
#691670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#691680000000
0!
0%
b0 *
0-
02
b0 6
#691690000000
1!
1%
1-
12
#691700000000
0!
0%
b1 *
0-
02
b1 6
#691710000000
1!
1%
1-
12
#691720000000
0!
0%
b10 *
0-
02
b10 6
#691730000000
1!
1%
1-
12
#691740000000
0!
0%
b11 *
0-
02
b11 6
#691750000000
1!
1%
1-
12
15
#691760000000
0!
0%
b100 *
0-
02
b100 6
#691770000000
1!
1%
1-
12
#691780000000
0!
0%
b101 *
0-
02
b101 6
#691790000000
1!
1%
1-
12
#691800000000
0!
0%
b110 *
0-
02
b110 6
#691810000000
1!
1%
1-
12
#691820000000
0!
0%
b111 *
0-
02
b111 6
#691830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#691840000000
0!
0%
b0 *
0-
02
b0 6
#691850000000
1!
1%
1-
12
#691860000000
0!
0%
b1 *
0-
02
b1 6
#691870000000
1!
1%
1-
12
#691880000000
0!
0%
b10 *
0-
02
b10 6
#691890000000
1!
1%
1-
12
#691900000000
0!
0%
b11 *
0-
02
b11 6
#691910000000
1!
1%
1-
12
15
#691920000000
0!
0%
b100 *
0-
02
b100 6
#691930000000
1!
1%
1-
12
#691940000000
0!
0%
b101 *
0-
02
b101 6
#691950000000
1!
1%
1-
12
#691960000000
0!
0%
b110 *
0-
02
b110 6
#691970000000
1!
1%
1-
12
#691980000000
0!
0%
b111 *
0-
02
b111 6
#691990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#692000000000
0!
0%
b0 *
0-
02
b0 6
#692010000000
1!
1%
1-
12
#692020000000
0!
0%
b1 *
0-
02
b1 6
#692030000000
1!
1%
1-
12
#692040000000
0!
0%
b10 *
0-
02
b10 6
#692050000000
1!
1%
1-
12
#692060000000
0!
0%
b11 *
0-
02
b11 6
#692070000000
1!
1%
1-
12
15
#692080000000
0!
0%
b100 *
0-
02
b100 6
#692090000000
1!
1%
1-
12
#692100000000
0!
0%
b101 *
0-
02
b101 6
#692110000000
1!
1%
1-
12
#692120000000
0!
0%
b110 *
0-
02
b110 6
#692130000000
1!
1%
1-
12
#692140000000
0!
0%
b111 *
0-
02
b111 6
#692150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#692160000000
0!
0%
b0 *
0-
02
b0 6
#692170000000
1!
1%
1-
12
#692180000000
0!
0%
b1 *
0-
02
b1 6
#692190000000
1!
1%
1-
12
#692200000000
0!
0%
b10 *
0-
02
b10 6
#692210000000
1!
1%
1-
12
#692220000000
0!
0%
b11 *
0-
02
b11 6
#692230000000
1!
1%
1-
12
15
#692240000000
0!
0%
b100 *
0-
02
b100 6
#692250000000
1!
1%
1-
12
#692260000000
0!
0%
b101 *
0-
02
b101 6
#692270000000
1!
1%
1-
12
#692280000000
0!
0%
b110 *
0-
02
b110 6
#692290000000
1!
1%
1-
12
#692300000000
0!
0%
b111 *
0-
02
b111 6
#692310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#692320000000
0!
0%
b0 *
0-
02
b0 6
#692330000000
1!
1%
1-
12
#692340000000
0!
0%
b1 *
0-
02
b1 6
#692350000000
1!
1%
1-
12
#692360000000
0!
0%
b10 *
0-
02
b10 6
#692370000000
1!
1%
1-
12
#692380000000
0!
0%
b11 *
0-
02
b11 6
#692390000000
1!
1%
1-
12
15
#692400000000
0!
0%
b100 *
0-
02
b100 6
#692410000000
1!
1%
1-
12
#692420000000
0!
0%
b101 *
0-
02
b101 6
#692430000000
1!
1%
1-
12
#692440000000
0!
0%
b110 *
0-
02
b110 6
#692450000000
1!
1%
1-
12
#692460000000
0!
0%
b111 *
0-
02
b111 6
#692470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#692480000000
0!
0%
b0 *
0-
02
b0 6
#692490000000
1!
1%
1-
12
#692500000000
0!
0%
b1 *
0-
02
b1 6
#692510000000
1!
1%
1-
12
#692520000000
0!
0%
b10 *
0-
02
b10 6
#692530000000
1!
1%
1-
12
#692540000000
0!
0%
b11 *
0-
02
b11 6
#692550000000
1!
1%
1-
12
15
#692560000000
0!
0%
b100 *
0-
02
b100 6
#692570000000
1!
1%
1-
12
#692580000000
0!
0%
b101 *
0-
02
b101 6
#692590000000
1!
1%
1-
12
#692600000000
0!
0%
b110 *
0-
02
b110 6
#692610000000
1!
1%
1-
12
#692620000000
0!
0%
b111 *
0-
02
b111 6
#692630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#692640000000
0!
0%
b0 *
0-
02
b0 6
#692650000000
1!
1%
1-
12
#692660000000
0!
0%
b1 *
0-
02
b1 6
#692670000000
1!
1%
1-
12
#692680000000
0!
0%
b10 *
0-
02
b10 6
#692690000000
1!
1%
1-
12
#692700000000
0!
0%
b11 *
0-
02
b11 6
#692710000000
1!
1%
1-
12
15
#692720000000
0!
0%
b100 *
0-
02
b100 6
#692730000000
1!
1%
1-
12
#692740000000
0!
0%
b101 *
0-
02
b101 6
#692750000000
1!
1%
1-
12
#692760000000
0!
0%
b110 *
0-
02
b110 6
#692770000000
1!
1%
1-
12
#692780000000
0!
0%
b111 *
0-
02
b111 6
#692790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#692800000000
0!
0%
b0 *
0-
02
b0 6
#692810000000
1!
1%
1-
12
#692820000000
0!
0%
b1 *
0-
02
b1 6
#692830000000
1!
1%
1-
12
#692840000000
0!
0%
b10 *
0-
02
b10 6
#692850000000
1!
1%
1-
12
#692860000000
0!
0%
b11 *
0-
02
b11 6
#692870000000
1!
1%
1-
12
15
#692880000000
0!
0%
b100 *
0-
02
b100 6
#692890000000
1!
1%
1-
12
#692900000000
0!
0%
b101 *
0-
02
b101 6
#692910000000
1!
1%
1-
12
#692920000000
0!
0%
b110 *
0-
02
b110 6
#692930000000
1!
1%
1-
12
#692940000000
0!
0%
b111 *
0-
02
b111 6
#692950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#692960000000
0!
0%
b0 *
0-
02
b0 6
#692970000000
1!
1%
1-
12
#692980000000
0!
0%
b1 *
0-
02
b1 6
#692990000000
1!
1%
1-
12
#693000000000
0!
0%
b10 *
0-
02
b10 6
#693010000000
1!
1%
1-
12
#693020000000
0!
0%
b11 *
0-
02
b11 6
#693030000000
1!
1%
1-
12
15
#693040000000
0!
0%
b100 *
0-
02
b100 6
#693050000000
1!
1%
1-
12
#693060000000
0!
0%
b101 *
0-
02
b101 6
#693070000000
1!
1%
1-
12
#693080000000
0!
0%
b110 *
0-
02
b110 6
#693090000000
1!
1%
1-
12
#693100000000
0!
0%
b111 *
0-
02
b111 6
#693110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#693120000000
0!
0%
b0 *
0-
02
b0 6
#693130000000
1!
1%
1-
12
#693140000000
0!
0%
b1 *
0-
02
b1 6
#693150000000
1!
1%
1-
12
#693160000000
0!
0%
b10 *
0-
02
b10 6
#693170000000
1!
1%
1-
12
#693180000000
0!
0%
b11 *
0-
02
b11 6
#693190000000
1!
1%
1-
12
15
#693200000000
0!
0%
b100 *
0-
02
b100 6
#693210000000
1!
1%
1-
12
#693220000000
0!
0%
b101 *
0-
02
b101 6
#693230000000
1!
1%
1-
12
#693240000000
0!
0%
b110 *
0-
02
b110 6
#693250000000
1!
1%
1-
12
#693260000000
0!
0%
b111 *
0-
02
b111 6
#693270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#693280000000
0!
0%
b0 *
0-
02
b0 6
#693290000000
1!
1%
1-
12
#693300000000
0!
0%
b1 *
0-
02
b1 6
#693310000000
1!
1%
1-
12
#693320000000
0!
0%
b10 *
0-
02
b10 6
#693330000000
1!
1%
1-
12
#693340000000
0!
0%
b11 *
0-
02
b11 6
#693350000000
1!
1%
1-
12
15
#693360000000
0!
0%
b100 *
0-
02
b100 6
#693370000000
1!
1%
1-
12
#693380000000
0!
0%
b101 *
0-
02
b101 6
#693390000000
1!
1%
1-
12
#693400000000
0!
0%
b110 *
0-
02
b110 6
#693410000000
1!
1%
1-
12
#693420000000
0!
0%
b111 *
0-
02
b111 6
#693430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#693440000000
0!
0%
b0 *
0-
02
b0 6
#693450000000
1!
1%
1-
12
#693460000000
0!
0%
b1 *
0-
02
b1 6
#693470000000
1!
1%
1-
12
#693480000000
0!
0%
b10 *
0-
02
b10 6
#693490000000
1!
1%
1-
12
#693500000000
0!
0%
b11 *
0-
02
b11 6
#693510000000
1!
1%
1-
12
15
#693520000000
0!
0%
b100 *
0-
02
b100 6
#693530000000
1!
1%
1-
12
#693540000000
0!
0%
b101 *
0-
02
b101 6
#693550000000
1!
1%
1-
12
#693560000000
0!
0%
b110 *
0-
02
b110 6
#693570000000
1!
1%
1-
12
#693580000000
0!
0%
b111 *
0-
02
b111 6
#693590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#693600000000
0!
0%
b0 *
0-
02
b0 6
#693610000000
1!
1%
1-
12
#693620000000
0!
0%
b1 *
0-
02
b1 6
#693630000000
1!
1%
1-
12
#693640000000
0!
0%
b10 *
0-
02
b10 6
#693650000000
1!
1%
1-
12
#693660000000
0!
0%
b11 *
0-
02
b11 6
#693670000000
1!
1%
1-
12
15
#693680000000
0!
0%
b100 *
0-
02
b100 6
#693690000000
1!
1%
1-
12
#693700000000
0!
0%
b101 *
0-
02
b101 6
#693710000000
1!
1%
1-
12
#693720000000
0!
0%
b110 *
0-
02
b110 6
#693730000000
1!
1%
1-
12
#693740000000
0!
0%
b111 *
0-
02
b111 6
#693750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#693760000000
0!
0%
b0 *
0-
02
b0 6
#693770000000
1!
1%
1-
12
#693780000000
0!
0%
b1 *
0-
02
b1 6
#693790000000
1!
1%
1-
12
#693800000000
0!
0%
b10 *
0-
02
b10 6
#693810000000
1!
1%
1-
12
#693820000000
0!
0%
b11 *
0-
02
b11 6
#693830000000
1!
1%
1-
12
15
#693840000000
0!
0%
b100 *
0-
02
b100 6
#693850000000
1!
1%
1-
12
#693860000000
0!
0%
b101 *
0-
02
b101 6
#693870000000
1!
1%
1-
12
#693880000000
0!
0%
b110 *
0-
02
b110 6
#693890000000
1!
1%
1-
12
#693900000000
0!
0%
b111 *
0-
02
b111 6
#693910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#693920000000
0!
0%
b0 *
0-
02
b0 6
#693930000000
1!
1%
1-
12
#693940000000
0!
0%
b1 *
0-
02
b1 6
#693950000000
1!
1%
1-
12
#693960000000
0!
0%
b10 *
0-
02
b10 6
#693970000000
1!
1%
1-
12
#693980000000
0!
0%
b11 *
0-
02
b11 6
#693990000000
1!
1%
1-
12
15
#694000000000
0!
0%
b100 *
0-
02
b100 6
#694010000000
1!
1%
1-
12
#694020000000
0!
0%
b101 *
0-
02
b101 6
#694030000000
1!
1%
1-
12
#694040000000
0!
0%
b110 *
0-
02
b110 6
#694050000000
1!
1%
1-
12
#694060000000
0!
0%
b111 *
0-
02
b111 6
#694070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#694080000000
0!
0%
b0 *
0-
02
b0 6
#694090000000
1!
1%
1-
12
#694100000000
0!
0%
b1 *
0-
02
b1 6
#694110000000
1!
1%
1-
12
#694120000000
0!
0%
b10 *
0-
02
b10 6
#694130000000
1!
1%
1-
12
#694140000000
0!
0%
b11 *
0-
02
b11 6
#694150000000
1!
1%
1-
12
15
#694160000000
0!
0%
b100 *
0-
02
b100 6
#694170000000
1!
1%
1-
12
#694180000000
0!
0%
b101 *
0-
02
b101 6
#694190000000
1!
1%
1-
12
#694200000000
0!
0%
b110 *
0-
02
b110 6
#694210000000
1!
1%
1-
12
#694220000000
0!
0%
b111 *
0-
02
b111 6
#694230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#694240000000
0!
0%
b0 *
0-
02
b0 6
#694250000000
1!
1%
1-
12
#694260000000
0!
0%
b1 *
0-
02
b1 6
#694270000000
1!
1%
1-
12
#694280000000
0!
0%
b10 *
0-
02
b10 6
#694290000000
1!
1%
1-
12
#694300000000
0!
0%
b11 *
0-
02
b11 6
#694310000000
1!
1%
1-
12
15
#694320000000
0!
0%
b100 *
0-
02
b100 6
#694330000000
1!
1%
1-
12
#694340000000
0!
0%
b101 *
0-
02
b101 6
#694350000000
1!
1%
1-
12
#694360000000
0!
0%
b110 *
0-
02
b110 6
#694370000000
1!
1%
1-
12
#694380000000
0!
0%
b111 *
0-
02
b111 6
#694390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#694400000000
0!
0%
b0 *
0-
02
b0 6
#694410000000
1!
1%
1-
12
#694420000000
0!
0%
b1 *
0-
02
b1 6
#694430000000
1!
1%
1-
12
#694440000000
0!
0%
b10 *
0-
02
b10 6
#694450000000
1!
1%
1-
12
#694460000000
0!
0%
b11 *
0-
02
b11 6
#694470000000
1!
1%
1-
12
15
#694480000000
0!
0%
b100 *
0-
02
b100 6
#694490000000
1!
1%
1-
12
#694500000000
0!
0%
b101 *
0-
02
b101 6
#694510000000
1!
1%
1-
12
#694520000000
0!
0%
b110 *
0-
02
b110 6
#694530000000
1!
1%
1-
12
#694540000000
0!
0%
b111 *
0-
02
b111 6
#694550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#694560000000
0!
0%
b0 *
0-
02
b0 6
#694570000000
1!
1%
1-
12
#694580000000
0!
0%
b1 *
0-
02
b1 6
#694590000000
1!
1%
1-
12
#694600000000
0!
0%
b10 *
0-
02
b10 6
#694610000000
1!
1%
1-
12
#694620000000
0!
0%
b11 *
0-
02
b11 6
#694630000000
1!
1%
1-
12
15
#694640000000
0!
0%
b100 *
0-
02
b100 6
#694650000000
1!
1%
1-
12
#694660000000
0!
0%
b101 *
0-
02
b101 6
#694670000000
1!
1%
1-
12
#694680000000
0!
0%
b110 *
0-
02
b110 6
#694690000000
1!
1%
1-
12
#694700000000
0!
0%
b111 *
0-
02
b111 6
#694710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#694720000000
0!
0%
b0 *
0-
02
b0 6
#694730000000
1!
1%
1-
12
#694740000000
0!
0%
b1 *
0-
02
b1 6
#694750000000
1!
1%
1-
12
#694760000000
0!
0%
b10 *
0-
02
b10 6
#694770000000
1!
1%
1-
12
#694780000000
0!
0%
b11 *
0-
02
b11 6
#694790000000
1!
1%
1-
12
15
#694800000000
0!
0%
b100 *
0-
02
b100 6
#694810000000
1!
1%
1-
12
#694820000000
0!
0%
b101 *
0-
02
b101 6
#694830000000
1!
1%
1-
12
#694840000000
0!
0%
b110 *
0-
02
b110 6
#694850000000
1!
1%
1-
12
#694860000000
0!
0%
b111 *
0-
02
b111 6
#694870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#694880000000
0!
0%
b0 *
0-
02
b0 6
#694890000000
1!
1%
1-
12
#694900000000
0!
0%
b1 *
0-
02
b1 6
#694910000000
1!
1%
1-
12
#694920000000
0!
0%
b10 *
0-
02
b10 6
#694930000000
1!
1%
1-
12
#694940000000
0!
0%
b11 *
0-
02
b11 6
#694950000000
1!
1%
1-
12
15
#694960000000
0!
0%
b100 *
0-
02
b100 6
#694970000000
1!
1%
1-
12
#694980000000
0!
0%
b101 *
0-
02
b101 6
#694990000000
1!
1%
1-
12
#695000000000
0!
0%
b110 *
0-
02
b110 6
#695010000000
1!
1%
1-
12
#695020000000
0!
0%
b111 *
0-
02
b111 6
#695030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#695040000000
0!
0%
b0 *
0-
02
b0 6
#695050000000
1!
1%
1-
12
#695060000000
0!
0%
b1 *
0-
02
b1 6
#695070000000
1!
1%
1-
12
#695080000000
0!
0%
b10 *
0-
02
b10 6
#695090000000
1!
1%
1-
12
#695100000000
0!
0%
b11 *
0-
02
b11 6
#695110000000
1!
1%
1-
12
15
#695120000000
0!
0%
b100 *
0-
02
b100 6
#695130000000
1!
1%
1-
12
#695140000000
0!
0%
b101 *
0-
02
b101 6
#695150000000
1!
1%
1-
12
#695160000000
0!
0%
b110 *
0-
02
b110 6
#695170000000
1!
1%
1-
12
#695180000000
0!
0%
b111 *
0-
02
b111 6
#695190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#695200000000
0!
0%
b0 *
0-
02
b0 6
#695210000000
1!
1%
1-
12
#695220000000
0!
0%
b1 *
0-
02
b1 6
#695230000000
1!
1%
1-
12
#695240000000
0!
0%
b10 *
0-
02
b10 6
#695250000000
1!
1%
1-
12
#695260000000
0!
0%
b11 *
0-
02
b11 6
#695270000000
1!
1%
1-
12
15
#695280000000
0!
0%
b100 *
0-
02
b100 6
#695290000000
1!
1%
1-
12
#695300000000
0!
0%
b101 *
0-
02
b101 6
#695310000000
1!
1%
1-
12
#695320000000
0!
0%
b110 *
0-
02
b110 6
#695330000000
1!
1%
1-
12
#695340000000
0!
0%
b111 *
0-
02
b111 6
#695350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#695360000000
0!
0%
b0 *
0-
02
b0 6
#695370000000
1!
1%
1-
12
#695380000000
0!
0%
b1 *
0-
02
b1 6
#695390000000
1!
1%
1-
12
#695400000000
0!
0%
b10 *
0-
02
b10 6
#695410000000
1!
1%
1-
12
#695420000000
0!
0%
b11 *
0-
02
b11 6
#695430000000
1!
1%
1-
12
15
#695440000000
0!
0%
b100 *
0-
02
b100 6
#695450000000
1!
1%
1-
12
#695460000000
0!
0%
b101 *
0-
02
b101 6
#695470000000
1!
1%
1-
12
#695480000000
0!
0%
b110 *
0-
02
b110 6
#695490000000
1!
1%
1-
12
#695500000000
0!
0%
b111 *
0-
02
b111 6
#695510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#695520000000
0!
0%
b0 *
0-
02
b0 6
#695530000000
1!
1%
1-
12
#695540000000
0!
0%
b1 *
0-
02
b1 6
#695550000000
1!
1%
1-
12
#695560000000
0!
0%
b10 *
0-
02
b10 6
#695570000000
1!
1%
1-
12
#695580000000
0!
0%
b11 *
0-
02
b11 6
#695590000000
1!
1%
1-
12
15
#695600000000
0!
0%
b100 *
0-
02
b100 6
#695610000000
1!
1%
1-
12
#695620000000
0!
0%
b101 *
0-
02
b101 6
#695630000000
1!
1%
1-
12
#695640000000
0!
0%
b110 *
0-
02
b110 6
#695650000000
1!
1%
1-
12
#695660000000
0!
0%
b111 *
0-
02
b111 6
#695670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#695680000000
0!
0%
b0 *
0-
02
b0 6
#695690000000
1!
1%
1-
12
#695700000000
0!
0%
b1 *
0-
02
b1 6
#695710000000
1!
1%
1-
12
#695720000000
0!
0%
b10 *
0-
02
b10 6
#695730000000
1!
1%
1-
12
#695740000000
0!
0%
b11 *
0-
02
b11 6
#695750000000
1!
1%
1-
12
15
#695760000000
0!
0%
b100 *
0-
02
b100 6
#695770000000
1!
1%
1-
12
#695780000000
0!
0%
b101 *
0-
02
b101 6
#695790000000
1!
1%
1-
12
#695800000000
0!
0%
b110 *
0-
02
b110 6
#695810000000
1!
1%
1-
12
#695820000000
0!
0%
b111 *
0-
02
b111 6
#695830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#695840000000
0!
0%
b0 *
0-
02
b0 6
#695850000000
1!
1%
1-
12
#695860000000
0!
0%
b1 *
0-
02
b1 6
#695870000000
1!
1%
1-
12
#695880000000
0!
0%
b10 *
0-
02
b10 6
#695890000000
1!
1%
1-
12
#695900000000
0!
0%
b11 *
0-
02
b11 6
#695910000000
1!
1%
1-
12
15
#695920000000
0!
0%
b100 *
0-
02
b100 6
#695930000000
1!
1%
1-
12
#695940000000
0!
0%
b101 *
0-
02
b101 6
#695950000000
1!
1%
1-
12
#695960000000
0!
0%
b110 *
0-
02
b110 6
#695970000000
1!
1%
1-
12
#695980000000
0!
0%
b111 *
0-
02
b111 6
#695990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#696000000000
0!
0%
b0 *
0-
02
b0 6
#696010000000
1!
1%
1-
12
#696020000000
0!
0%
b1 *
0-
02
b1 6
#696030000000
1!
1%
1-
12
#696040000000
0!
0%
b10 *
0-
02
b10 6
#696050000000
1!
1%
1-
12
#696060000000
0!
0%
b11 *
0-
02
b11 6
#696070000000
1!
1%
1-
12
15
#696080000000
0!
0%
b100 *
0-
02
b100 6
#696090000000
1!
1%
1-
12
#696100000000
0!
0%
b101 *
0-
02
b101 6
#696110000000
1!
1%
1-
12
#696120000000
0!
0%
b110 *
0-
02
b110 6
#696130000000
1!
1%
1-
12
#696140000000
0!
0%
b111 *
0-
02
b111 6
#696150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#696160000000
0!
0%
b0 *
0-
02
b0 6
#696170000000
1!
1%
1-
12
#696180000000
0!
0%
b1 *
0-
02
b1 6
#696190000000
1!
1%
1-
12
#696200000000
0!
0%
b10 *
0-
02
b10 6
#696210000000
1!
1%
1-
12
#696220000000
0!
0%
b11 *
0-
02
b11 6
#696230000000
1!
1%
1-
12
15
#696240000000
0!
0%
b100 *
0-
02
b100 6
#696250000000
1!
1%
1-
12
#696260000000
0!
0%
b101 *
0-
02
b101 6
#696270000000
1!
1%
1-
12
#696280000000
0!
0%
b110 *
0-
02
b110 6
#696290000000
1!
1%
1-
12
#696300000000
0!
0%
b111 *
0-
02
b111 6
#696310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#696320000000
0!
0%
b0 *
0-
02
b0 6
#696330000000
1!
1%
1-
12
#696340000000
0!
0%
b1 *
0-
02
b1 6
#696350000000
1!
1%
1-
12
#696360000000
0!
0%
b10 *
0-
02
b10 6
#696370000000
1!
1%
1-
12
#696380000000
0!
0%
b11 *
0-
02
b11 6
#696390000000
1!
1%
1-
12
15
#696400000000
0!
0%
b100 *
0-
02
b100 6
#696410000000
1!
1%
1-
12
#696420000000
0!
0%
b101 *
0-
02
b101 6
#696430000000
1!
1%
1-
12
#696440000000
0!
0%
b110 *
0-
02
b110 6
#696450000000
1!
1%
1-
12
#696460000000
0!
0%
b111 *
0-
02
b111 6
#696470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#696480000000
0!
0%
b0 *
0-
02
b0 6
#696490000000
1!
1%
1-
12
#696500000000
0!
0%
b1 *
0-
02
b1 6
#696510000000
1!
1%
1-
12
#696520000000
0!
0%
b10 *
0-
02
b10 6
#696530000000
1!
1%
1-
12
#696540000000
0!
0%
b11 *
0-
02
b11 6
#696550000000
1!
1%
1-
12
15
#696560000000
0!
0%
b100 *
0-
02
b100 6
#696570000000
1!
1%
1-
12
#696580000000
0!
0%
b101 *
0-
02
b101 6
#696590000000
1!
1%
1-
12
#696600000000
0!
0%
b110 *
0-
02
b110 6
#696610000000
1!
1%
1-
12
#696620000000
0!
0%
b111 *
0-
02
b111 6
#696630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#696640000000
0!
0%
b0 *
0-
02
b0 6
#696650000000
1!
1%
1-
12
#696660000000
0!
0%
b1 *
0-
02
b1 6
#696670000000
1!
1%
1-
12
#696680000000
0!
0%
b10 *
0-
02
b10 6
#696690000000
1!
1%
1-
12
#696700000000
0!
0%
b11 *
0-
02
b11 6
#696710000000
1!
1%
1-
12
15
#696720000000
0!
0%
b100 *
0-
02
b100 6
#696730000000
1!
1%
1-
12
#696740000000
0!
0%
b101 *
0-
02
b101 6
#696750000000
1!
1%
1-
12
#696760000000
0!
0%
b110 *
0-
02
b110 6
#696770000000
1!
1%
1-
12
#696780000000
0!
0%
b111 *
0-
02
b111 6
#696790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#696800000000
0!
0%
b0 *
0-
02
b0 6
#696810000000
1!
1%
1-
12
#696820000000
0!
0%
b1 *
0-
02
b1 6
#696830000000
1!
1%
1-
12
#696840000000
0!
0%
b10 *
0-
02
b10 6
#696850000000
1!
1%
1-
12
#696860000000
0!
0%
b11 *
0-
02
b11 6
#696870000000
1!
1%
1-
12
15
#696880000000
0!
0%
b100 *
0-
02
b100 6
#696890000000
1!
1%
1-
12
#696900000000
0!
0%
b101 *
0-
02
b101 6
#696910000000
1!
1%
1-
12
#696920000000
0!
0%
b110 *
0-
02
b110 6
#696930000000
1!
1%
1-
12
#696940000000
0!
0%
b111 *
0-
02
b111 6
#696950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#696960000000
0!
0%
b0 *
0-
02
b0 6
#696970000000
1!
1%
1-
12
#696980000000
0!
0%
b1 *
0-
02
b1 6
#696990000000
1!
1%
1-
12
#697000000000
0!
0%
b10 *
0-
02
b10 6
#697010000000
1!
1%
1-
12
#697020000000
0!
0%
b11 *
0-
02
b11 6
#697030000000
1!
1%
1-
12
15
#697040000000
0!
0%
b100 *
0-
02
b100 6
#697050000000
1!
1%
1-
12
#697060000000
0!
0%
b101 *
0-
02
b101 6
#697070000000
1!
1%
1-
12
#697080000000
0!
0%
b110 *
0-
02
b110 6
#697090000000
1!
1%
1-
12
#697100000000
0!
0%
b111 *
0-
02
b111 6
#697110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#697120000000
0!
0%
b0 *
0-
02
b0 6
#697130000000
1!
1%
1-
12
#697140000000
0!
0%
b1 *
0-
02
b1 6
#697150000000
1!
1%
1-
12
#697160000000
0!
0%
b10 *
0-
02
b10 6
#697170000000
1!
1%
1-
12
#697180000000
0!
0%
b11 *
0-
02
b11 6
#697190000000
1!
1%
1-
12
15
#697200000000
0!
0%
b100 *
0-
02
b100 6
#697210000000
1!
1%
1-
12
#697220000000
0!
0%
b101 *
0-
02
b101 6
#697230000000
1!
1%
1-
12
#697240000000
0!
0%
b110 *
0-
02
b110 6
#697250000000
1!
1%
1-
12
#697260000000
0!
0%
b111 *
0-
02
b111 6
#697270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#697280000000
0!
0%
b0 *
0-
02
b0 6
#697290000000
1!
1%
1-
12
#697300000000
0!
0%
b1 *
0-
02
b1 6
#697310000000
1!
1%
1-
12
#697320000000
0!
0%
b10 *
0-
02
b10 6
#697330000000
1!
1%
1-
12
#697340000000
0!
0%
b11 *
0-
02
b11 6
#697350000000
1!
1%
1-
12
15
#697360000000
0!
0%
b100 *
0-
02
b100 6
#697370000000
1!
1%
1-
12
#697380000000
0!
0%
b101 *
0-
02
b101 6
#697390000000
1!
1%
1-
12
#697400000000
0!
0%
b110 *
0-
02
b110 6
#697410000000
1!
1%
1-
12
#697420000000
0!
0%
b111 *
0-
02
b111 6
#697430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#697440000000
0!
0%
b0 *
0-
02
b0 6
#697450000000
1!
1%
1-
12
#697460000000
0!
0%
b1 *
0-
02
b1 6
#697470000000
1!
1%
1-
12
#697480000000
0!
0%
b10 *
0-
02
b10 6
#697490000000
1!
1%
1-
12
#697500000000
0!
0%
b11 *
0-
02
b11 6
#697510000000
1!
1%
1-
12
15
#697520000000
0!
0%
b100 *
0-
02
b100 6
#697530000000
1!
1%
1-
12
#697540000000
0!
0%
b101 *
0-
02
b101 6
#697550000000
1!
1%
1-
12
#697560000000
0!
0%
b110 *
0-
02
b110 6
#697570000000
1!
1%
1-
12
#697580000000
0!
0%
b111 *
0-
02
b111 6
#697590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#697600000000
0!
0%
b0 *
0-
02
b0 6
#697610000000
1!
1%
1-
12
#697620000000
0!
0%
b1 *
0-
02
b1 6
#697630000000
1!
1%
1-
12
#697640000000
0!
0%
b10 *
0-
02
b10 6
#697650000000
1!
1%
1-
12
#697660000000
0!
0%
b11 *
0-
02
b11 6
#697670000000
1!
1%
1-
12
15
#697680000000
0!
0%
b100 *
0-
02
b100 6
#697690000000
1!
1%
1-
12
#697700000000
0!
0%
b101 *
0-
02
b101 6
#697710000000
1!
1%
1-
12
#697720000000
0!
0%
b110 *
0-
02
b110 6
#697730000000
1!
1%
1-
12
#697740000000
0!
0%
b111 *
0-
02
b111 6
#697750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#697760000000
0!
0%
b0 *
0-
02
b0 6
#697770000000
1!
1%
1-
12
#697780000000
0!
0%
b1 *
0-
02
b1 6
#697790000000
1!
1%
1-
12
#697800000000
0!
0%
b10 *
0-
02
b10 6
#697810000000
1!
1%
1-
12
#697820000000
0!
0%
b11 *
0-
02
b11 6
#697830000000
1!
1%
1-
12
15
#697840000000
0!
0%
b100 *
0-
02
b100 6
#697850000000
1!
1%
1-
12
#697860000000
0!
0%
b101 *
0-
02
b101 6
#697870000000
1!
1%
1-
12
#697880000000
0!
0%
b110 *
0-
02
b110 6
#697890000000
1!
1%
1-
12
#697900000000
0!
0%
b111 *
0-
02
b111 6
#697910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#697920000000
0!
0%
b0 *
0-
02
b0 6
#697930000000
1!
1%
1-
12
#697940000000
0!
0%
b1 *
0-
02
b1 6
#697950000000
1!
1%
1-
12
#697960000000
0!
0%
b10 *
0-
02
b10 6
#697970000000
1!
1%
1-
12
#697980000000
0!
0%
b11 *
0-
02
b11 6
#697990000000
1!
1%
1-
12
15
#698000000000
0!
0%
b100 *
0-
02
b100 6
#698010000000
1!
1%
1-
12
#698020000000
0!
0%
b101 *
0-
02
b101 6
#698030000000
1!
1%
1-
12
#698040000000
0!
0%
b110 *
0-
02
b110 6
#698050000000
1!
1%
1-
12
#698060000000
0!
0%
b111 *
0-
02
b111 6
#698070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#698080000000
0!
0%
b0 *
0-
02
b0 6
#698090000000
1!
1%
1-
12
#698100000000
0!
0%
b1 *
0-
02
b1 6
#698110000000
1!
1%
1-
12
#698120000000
0!
0%
b10 *
0-
02
b10 6
#698130000000
1!
1%
1-
12
#698140000000
0!
0%
b11 *
0-
02
b11 6
#698150000000
1!
1%
1-
12
15
#698160000000
0!
0%
b100 *
0-
02
b100 6
#698170000000
1!
1%
1-
12
#698180000000
0!
0%
b101 *
0-
02
b101 6
#698190000000
1!
1%
1-
12
#698200000000
0!
0%
b110 *
0-
02
b110 6
#698210000000
1!
1%
1-
12
#698220000000
0!
0%
b111 *
0-
02
b111 6
#698230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#698240000000
0!
0%
b0 *
0-
02
b0 6
#698250000000
1!
1%
1-
12
#698260000000
0!
0%
b1 *
0-
02
b1 6
#698270000000
1!
1%
1-
12
#698280000000
0!
0%
b10 *
0-
02
b10 6
#698290000000
1!
1%
1-
12
#698300000000
0!
0%
b11 *
0-
02
b11 6
#698310000000
1!
1%
1-
12
15
#698320000000
0!
0%
b100 *
0-
02
b100 6
#698330000000
1!
1%
1-
12
#698340000000
0!
0%
b101 *
0-
02
b101 6
#698350000000
1!
1%
1-
12
#698360000000
0!
0%
b110 *
0-
02
b110 6
#698370000000
1!
1%
1-
12
#698380000000
0!
0%
b111 *
0-
02
b111 6
#698390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#698400000000
0!
0%
b0 *
0-
02
b0 6
#698410000000
1!
1%
1-
12
#698420000000
0!
0%
b1 *
0-
02
b1 6
#698430000000
1!
1%
1-
12
#698440000000
0!
0%
b10 *
0-
02
b10 6
#698450000000
1!
1%
1-
12
#698460000000
0!
0%
b11 *
0-
02
b11 6
#698470000000
1!
1%
1-
12
15
#698480000000
0!
0%
b100 *
0-
02
b100 6
#698490000000
1!
1%
1-
12
#698500000000
0!
0%
b101 *
0-
02
b101 6
#698510000000
1!
1%
1-
12
#698520000000
0!
0%
b110 *
0-
02
b110 6
#698530000000
1!
1%
1-
12
#698540000000
0!
0%
b111 *
0-
02
b111 6
#698550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#698560000000
0!
0%
b0 *
0-
02
b0 6
#698570000000
1!
1%
1-
12
#698580000000
0!
0%
b1 *
0-
02
b1 6
#698590000000
1!
1%
1-
12
#698600000000
0!
0%
b10 *
0-
02
b10 6
#698610000000
1!
1%
1-
12
#698620000000
0!
0%
b11 *
0-
02
b11 6
#698630000000
1!
1%
1-
12
15
#698640000000
0!
0%
b100 *
0-
02
b100 6
#698650000000
1!
1%
1-
12
#698660000000
0!
0%
b101 *
0-
02
b101 6
#698670000000
1!
1%
1-
12
#698680000000
0!
0%
b110 *
0-
02
b110 6
#698690000000
1!
1%
1-
12
#698700000000
0!
0%
b111 *
0-
02
b111 6
#698710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#698720000000
0!
0%
b0 *
0-
02
b0 6
#698730000000
1!
1%
1-
12
#698740000000
0!
0%
b1 *
0-
02
b1 6
#698750000000
1!
1%
1-
12
#698760000000
0!
0%
b10 *
0-
02
b10 6
#698770000000
1!
1%
1-
12
#698780000000
0!
0%
b11 *
0-
02
b11 6
#698790000000
1!
1%
1-
12
15
#698800000000
0!
0%
b100 *
0-
02
b100 6
#698810000000
1!
1%
1-
12
#698820000000
0!
0%
b101 *
0-
02
b101 6
#698830000000
1!
1%
1-
12
#698840000000
0!
0%
b110 *
0-
02
b110 6
#698850000000
1!
1%
1-
12
#698860000000
0!
0%
b111 *
0-
02
b111 6
#698870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#698880000000
0!
0%
b0 *
0-
02
b0 6
#698890000000
1!
1%
1-
12
#698900000000
0!
0%
b1 *
0-
02
b1 6
#698910000000
1!
1%
1-
12
#698920000000
0!
0%
b10 *
0-
02
b10 6
#698930000000
1!
1%
1-
12
#698940000000
0!
0%
b11 *
0-
02
b11 6
#698950000000
1!
1%
1-
12
15
#698960000000
0!
0%
b100 *
0-
02
b100 6
#698970000000
1!
1%
1-
12
#698980000000
0!
0%
b101 *
0-
02
b101 6
#698990000000
1!
1%
1-
12
#699000000000
0!
0%
b110 *
0-
02
b110 6
#699010000000
1!
1%
1-
12
#699020000000
0!
0%
b111 *
0-
02
b111 6
#699030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#699040000000
0!
0%
b0 *
0-
02
b0 6
#699050000000
1!
1%
1-
12
#699060000000
0!
0%
b1 *
0-
02
b1 6
#699070000000
1!
1%
1-
12
#699080000000
0!
0%
b10 *
0-
02
b10 6
#699090000000
1!
1%
1-
12
#699100000000
0!
0%
b11 *
0-
02
b11 6
#699110000000
1!
1%
1-
12
15
#699120000000
0!
0%
b100 *
0-
02
b100 6
#699130000000
1!
1%
1-
12
#699140000000
0!
0%
b101 *
0-
02
b101 6
#699150000000
1!
1%
1-
12
#699160000000
0!
0%
b110 *
0-
02
b110 6
#699170000000
1!
1%
1-
12
#699180000000
0!
0%
b111 *
0-
02
b111 6
#699190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#699200000000
0!
0%
b0 *
0-
02
b0 6
#699210000000
1!
1%
1-
12
#699220000000
0!
0%
b1 *
0-
02
b1 6
#699230000000
1!
1%
1-
12
#699240000000
0!
0%
b10 *
0-
02
b10 6
#699250000000
1!
1%
1-
12
#699260000000
0!
0%
b11 *
0-
02
b11 6
#699270000000
1!
1%
1-
12
15
#699280000000
0!
0%
b100 *
0-
02
b100 6
#699290000000
1!
1%
1-
12
#699300000000
0!
0%
b101 *
0-
02
b101 6
#699310000000
1!
1%
1-
12
#699320000000
0!
0%
b110 *
0-
02
b110 6
#699330000000
1!
1%
1-
12
#699340000000
0!
0%
b111 *
0-
02
b111 6
#699350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#699360000000
0!
0%
b0 *
0-
02
b0 6
#699370000000
1!
1%
1-
12
#699380000000
0!
0%
b1 *
0-
02
b1 6
#699390000000
1!
1%
1-
12
#699400000000
0!
0%
b10 *
0-
02
b10 6
#699410000000
1!
1%
1-
12
#699420000000
0!
0%
b11 *
0-
02
b11 6
#699430000000
1!
1%
1-
12
15
#699440000000
0!
0%
b100 *
0-
02
b100 6
#699450000000
1!
1%
1-
12
#699460000000
0!
0%
b101 *
0-
02
b101 6
#699470000000
1!
1%
1-
12
#699480000000
0!
0%
b110 *
0-
02
b110 6
#699490000000
1!
1%
1-
12
#699500000000
0!
0%
b111 *
0-
02
b111 6
#699510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#699520000000
0!
0%
b0 *
0-
02
b0 6
#699530000000
1!
1%
1-
12
#699540000000
0!
0%
b1 *
0-
02
b1 6
#699550000000
1!
1%
1-
12
#699560000000
0!
0%
b10 *
0-
02
b10 6
#699570000000
1!
1%
1-
12
#699580000000
0!
0%
b11 *
0-
02
b11 6
#699590000000
1!
1%
1-
12
15
#699600000000
0!
0%
b100 *
0-
02
b100 6
#699610000000
1!
1%
1-
12
#699620000000
0!
0%
b101 *
0-
02
b101 6
#699630000000
1!
1%
1-
12
#699640000000
0!
0%
b110 *
0-
02
b110 6
#699650000000
1!
1%
1-
12
#699660000000
0!
0%
b111 *
0-
02
b111 6
#699670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#699680000000
0!
0%
b0 *
0-
02
b0 6
#699690000000
1!
1%
1-
12
#699700000000
0!
0%
b1 *
0-
02
b1 6
#699710000000
1!
1%
1-
12
#699720000000
0!
0%
b10 *
0-
02
b10 6
#699730000000
1!
1%
1-
12
#699740000000
0!
0%
b11 *
0-
02
b11 6
#699750000000
1!
1%
1-
12
15
#699760000000
0!
0%
b100 *
0-
02
b100 6
#699770000000
1!
1%
1-
12
#699780000000
0!
0%
b101 *
0-
02
b101 6
#699790000000
1!
1%
1-
12
#699800000000
0!
0%
b110 *
0-
02
b110 6
#699810000000
1!
1%
1-
12
#699820000000
0!
0%
b111 *
0-
02
b111 6
#699830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#699840000000
0!
0%
b0 *
0-
02
b0 6
#699850000000
1!
1%
1-
12
#699860000000
0!
0%
b1 *
0-
02
b1 6
#699870000000
1!
1%
1-
12
#699880000000
0!
0%
b10 *
0-
02
b10 6
#699890000000
1!
1%
1-
12
#699900000000
0!
0%
b11 *
0-
02
b11 6
#699910000000
1!
1%
1-
12
15
#699920000000
0!
0%
b100 *
0-
02
b100 6
#699930000000
1!
1%
1-
12
#699940000000
0!
0%
b101 *
0-
02
b101 6
#699950000000
1!
1%
1-
12
#699960000000
0!
0%
b110 *
0-
02
b110 6
#699970000000
1!
1%
1-
12
#699980000000
0!
0%
b111 *
0-
02
b111 6
#699990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#700000000000
0!
0%
b0 *
0-
02
b0 6
#700010000000
1!
1%
1-
12
#700020000000
0!
0%
b1 *
0-
02
b1 6
#700030000000
1!
1%
1-
12
#700040000000
0!
0%
b10 *
0-
02
b10 6
#700050000000
1!
1%
1-
12
#700060000000
0!
0%
b11 *
0-
02
b11 6
#700070000000
1!
1%
1-
12
15
#700080000000
0!
0%
b100 *
0-
02
b100 6
#700090000000
1!
1%
1-
12
#700100000000
0!
0%
b101 *
0-
02
b101 6
#700110000000
1!
1%
1-
12
#700120000000
0!
0%
b110 *
0-
02
b110 6
#700130000000
1!
1%
1-
12
#700140000000
0!
0%
b111 *
0-
02
b111 6
#700150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#700160000000
0!
0%
b0 *
0-
02
b0 6
#700170000000
1!
1%
1-
12
#700180000000
0!
0%
b1 *
0-
02
b1 6
#700190000000
1!
1%
1-
12
#700200000000
0!
0%
b10 *
0-
02
b10 6
#700210000000
1!
1%
1-
12
#700220000000
0!
0%
b11 *
0-
02
b11 6
#700230000000
1!
1%
1-
12
15
#700240000000
0!
0%
b100 *
0-
02
b100 6
#700250000000
1!
1%
1-
12
#700260000000
0!
0%
b101 *
0-
02
b101 6
#700270000000
1!
1%
1-
12
#700280000000
0!
0%
b110 *
0-
02
b110 6
#700290000000
1!
1%
1-
12
#700300000000
0!
0%
b111 *
0-
02
b111 6
#700310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#700320000000
0!
0%
b0 *
0-
02
b0 6
#700330000000
1!
1%
1-
12
#700340000000
0!
0%
b1 *
0-
02
b1 6
#700350000000
1!
1%
1-
12
#700360000000
0!
0%
b10 *
0-
02
b10 6
#700370000000
1!
1%
1-
12
#700380000000
0!
0%
b11 *
0-
02
b11 6
#700390000000
1!
1%
1-
12
15
#700400000000
0!
0%
b100 *
0-
02
b100 6
#700410000000
1!
1%
1-
12
#700420000000
0!
0%
b101 *
0-
02
b101 6
#700430000000
1!
1%
1-
12
#700440000000
0!
0%
b110 *
0-
02
b110 6
#700450000000
1!
1%
1-
12
#700460000000
0!
0%
b111 *
0-
02
b111 6
#700470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#700480000000
0!
0%
b0 *
0-
02
b0 6
#700490000000
1!
1%
1-
12
#700500000000
0!
0%
b1 *
0-
02
b1 6
#700510000000
1!
1%
1-
12
#700520000000
0!
0%
b10 *
0-
02
b10 6
#700530000000
1!
1%
1-
12
#700540000000
0!
0%
b11 *
0-
02
b11 6
#700550000000
1!
1%
1-
12
15
#700560000000
0!
0%
b100 *
0-
02
b100 6
#700570000000
1!
1%
1-
12
#700580000000
0!
0%
b101 *
0-
02
b101 6
#700590000000
1!
1%
1-
12
#700600000000
0!
0%
b110 *
0-
02
b110 6
#700610000000
1!
1%
1-
12
#700620000000
0!
0%
b111 *
0-
02
b111 6
#700630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#700640000000
0!
0%
b0 *
0-
02
b0 6
#700650000000
1!
1%
1-
12
#700660000000
0!
0%
b1 *
0-
02
b1 6
#700670000000
1!
1%
1-
12
#700680000000
0!
0%
b10 *
0-
02
b10 6
#700690000000
1!
1%
1-
12
#700700000000
0!
0%
b11 *
0-
02
b11 6
#700710000000
1!
1%
1-
12
15
#700720000000
0!
0%
b100 *
0-
02
b100 6
#700730000000
1!
1%
1-
12
#700740000000
0!
0%
b101 *
0-
02
b101 6
#700750000000
1!
1%
1-
12
#700760000000
0!
0%
b110 *
0-
02
b110 6
#700770000000
1!
1%
1-
12
#700780000000
0!
0%
b111 *
0-
02
b111 6
#700790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#700800000000
0!
0%
b0 *
0-
02
b0 6
#700810000000
1!
1%
1-
12
#700820000000
0!
0%
b1 *
0-
02
b1 6
#700830000000
1!
1%
1-
12
#700840000000
0!
0%
b10 *
0-
02
b10 6
#700850000000
1!
1%
1-
12
#700860000000
0!
0%
b11 *
0-
02
b11 6
#700870000000
1!
1%
1-
12
15
#700880000000
0!
0%
b100 *
0-
02
b100 6
#700890000000
1!
1%
1-
12
#700900000000
0!
0%
b101 *
0-
02
b101 6
#700910000000
1!
1%
1-
12
#700920000000
0!
0%
b110 *
0-
02
b110 6
#700930000000
1!
1%
1-
12
#700940000000
0!
0%
b111 *
0-
02
b111 6
#700950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#700960000000
0!
0%
b0 *
0-
02
b0 6
#700970000000
1!
1%
1-
12
#700980000000
0!
0%
b1 *
0-
02
b1 6
#700990000000
1!
1%
1-
12
#701000000000
0!
0%
b10 *
0-
02
b10 6
#701010000000
1!
1%
1-
12
#701020000000
0!
0%
b11 *
0-
02
b11 6
#701030000000
1!
1%
1-
12
15
#701040000000
0!
0%
b100 *
0-
02
b100 6
#701050000000
1!
1%
1-
12
#701060000000
0!
0%
b101 *
0-
02
b101 6
#701070000000
1!
1%
1-
12
#701080000000
0!
0%
b110 *
0-
02
b110 6
#701090000000
1!
1%
1-
12
#701100000000
0!
0%
b111 *
0-
02
b111 6
#701110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#701120000000
0!
0%
b0 *
0-
02
b0 6
#701130000000
1!
1%
1-
12
#701140000000
0!
0%
b1 *
0-
02
b1 6
#701150000000
1!
1%
1-
12
#701160000000
0!
0%
b10 *
0-
02
b10 6
#701170000000
1!
1%
1-
12
#701180000000
0!
0%
b11 *
0-
02
b11 6
#701190000000
1!
1%
1-
12
15
#701200000000
0!
0%
b100 *
0-
02
b100 6
#701210000000
1!
1%
1-
12
#701220000000
0!
0%
b101 *
0-
02
b101 6
#701230000000
1!
1%
1-
12
#701240000000
0!
0%
b110 *
0-
02
b110 6
#701250000000
1!
1%
1-
12
#701260000000
0!
0%
b111 *
0-
02
b111 6
#701270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#701280000000
0!
0%
b0 *
0-
02
b0 6
#701290000000
1!
1%
1-
12
#701300000000
0!
0%
b1 *
0-
02
b1 6
#701310000000
1!
1%
1-
12
#701320000000
0!
0%
b10 *
0-
02
b10 6
#701330000000
1!
1%
1-
12
#701340000000
0!
0%
b11 *
0-
02
b11 6
#701350000000
1!
1%
1-
12
15
#701360000000
0!
0%
b100 *
0-
02
b100 6
#701370000000
1!
1%
1-
12
#701380000000
0!
0%
b101 *
0-
02
b101 6
#701390000000
1!
1%
1-
12
#701400000000
0!
0%
b110 *
0-
02
b110 6
#701410000000
1!
1%
1-
12
#701420000000
0!
0%
b111 *
0-
02
b111 6
#701430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#701440000000
0!
0%
b0 *
0-
02
b0 6
#701450000000
1!
1%
1-
12
#701460000000
0!
0%
b1 *
0-
02
b1 6
#701470000000
1!
1%
1-
12
#701480000000
0!
0%
b10 *
0-
02
b10 6
#701490000000
1!
1%
1-
12
#701500000000
0!
0%
b11 *
0-
02
b11 6
#701510000000
1!
1%
1-
12
15
#701520000000
0!
0%
b100 *
0-
02
b100 6
#701530000000
1!
1%
1-
12
#701540000000
0!
0%
b101 *
0-
02
b101 6
#701550000000
1!
1%
1-
12
#701560000000
0!
0%
b110 *
0-
02
b110 6
#701570000000
1!
1%
1-
12
#701580000000
0!
0%
b111 *
0-
02
b111 6
#701590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#701600000000
0!
0%
b0 *
0-
02
b0 6
#701610000000
1!
1%
1-
12
#701620000000
0!
0%
b1 *
0-
02
b1 6
#701630000000
1!
1%
1-
12
#701640000000
0!
0%
b10 *
0-
02
b10 6
#701650000000
1!
1%
1-
12
#701660000000
0!
0%
b11 *
0-
02
b11 6
#701670000000
1!
1%
1-
12
15
#701680000000
0!
0%
b100 *
0-
02
b100 6
#701690000000
1!
1%
1-
12
#701700000000
0!
0%
b101 *
0-
02
b101 6
#701710000000
1!
1%
1-
12
#701720000000
0!
0%
b110 *
0-
02
b110 6
#701730000000
1!
1%
1-
12
#701740000000
0!
0%
b111 *
0-
02
b111 6
#701750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#701760000000
0!
0%
b0 *
0-
02
b0 6
#701770000000
1!
1%
1-
12
#701780000000
0!
0%
b1 *
0-
02
b1 6
#701790000000
1!
1%
1-
12
#701800000000
0!
0%
b10 *
0-
02
b10 6
#701810000000
1!
1%
1-
12
#701820000000
0!
0%
b11 *
0-
02
b11 6
#701830000000
1!
1%
1-
12
15
#701840000000
0!
0%
b100 *
0-
02
b100 6
#701850000000
1!
1%
1-
12
#701860000000
0!
0%
b101 *
0-
02
b101 6
#701870000000
1!
1%
1-
12
#701880000000
0!
0%
b110 *
0-
02
b110 6
#701890000000
1!
1%
1-
12
#701900000000
0!
0%
b111 *
0-
02
b111 6
#701910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#701920000000
0!
0%
b0 *
0-
02
b0 6
#701930000000
1!
1%
1-
12
#701940000000
0!
0%
b1 *
0-
02
b1 6
#701950000000
1!
1%
1-
12
#701960000000
0!
0%
b10 *
0-
02
b10 6
#701970000000
1!
1%
1-
12
#701980000000
0!
0%
b11 *
0-
02
b11 6
#701990000000
1!
1%
1-
12
15
#702000000000
0!
0%
b100 *
0-
02
b100 6
#702010000000
1!
1%
1-
12
#702020000000
0!
0%
b101 *
0-
02
b101 6
#702030000000
1!
1%
1-
12
#702040000000
0!
0%
b110 *
0-
02
b110 6
#702050000000
1!
1%
1-
12
#702060000000
0!
0%
b111 *
0-
02
b111 6
#702070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#702080000000
0!
0%
b0 *
0-
02
b0 6
#702090000000
1!
1%
1-
12
#702100000000
0!
0%
b1 *
0-
02
b1 6
#702110000000
1!
1%
1-
12
#702120000000
0!
0%
b10 *
0-
02
b10 6
#702130000000
1!
1%
1-
12
#702140000000
0!
0%
b11 *
0-
02
b11 6
#702150000000
1!
1%
1-
12
15
#702160000000
0!
0%
b100 *
0-
02
b100 6
#702170000000
1!
1%
1-
12
#702180000000
0!
0%
b101 *
0-
02
b101 6
#702190000000
1!
1%
1-
12
#702200000000
0!
0%
b110 *
0-
02
b110 6
#702210000000
1!
1%
1-
12
#702220000000
0!
0%
b111 *
0-
02
b111 6
#702230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#702240000000
0!
0%
b0 *
0-
02
b0 6
#702250000000
1!
1%
1-
12
#702260000000
0!
0%
b1 *
0-
02
b1 6
#702270000000
1!
1%
1-
12
#702280000000
0!
0%
b10 *
0-
02
b10 6
#702290000000
1!
1%
1-
12
#702300000000
0!
0%
b11 *
0-
02
b11 6
#702310000000
1!
1%
1-
12
15
#702320000000
0!
0%
b100 *
0-
02
b100 6
#702330000000
1!
1%
1-
12
#702340000000
0!
0%
b101 *
0-
02
b101 6
#702350000000
1!
1%
1-
12
#702360000000
0!
0%
b110 *
0-
02
b110 6
#702370000000
1!
1%
1-
12
#702380000000
0!
0%
b111 *
0-
02
b111 6
#702390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#702400000000
0!
0%
b0 *
0-
02
b0 6
#702410000000
1!
1%
1-
12
#702420000000
0!
0%
b1 *
0-
02
b1 6
#702430000000
1!
1%
1-
12
#702440000000
0!
0%
b10 *
0-
02
b10 6
#702450000000
1!
1%
1-
12
#702460000000
0!
0%
b11 *
0-
02
b11 6
#702470000000
1!
1%
1-
12
15
#702480000000
0!
0%
b100 *
0-
02
b100 6
#702490000000
1!
1%
1-
12
#702500000000
0!
0%
b101 *
0-
02
b101 6
#702510000000
1!
1%
1-
12
#702520000000
0!
0%
b110 *
0-
02
b110 6
#702530000000
1!
1%
1-
12
#702540000000
0!
0%
b111 *
0-
02
b111 6
#702550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#702560000000
0!
0%
b0 *
0-
02
b0 6
#702570000000
1!
1%
1-
12
#702580000000
0!
0%
b1 *
0-
02
b1 6
#702590000000
1!
1%
1-
12
#702600000000
0!
0%
b10 *
0-
02
b10 6
#702610000000
1!
1%
1-
12
#702620000000
0!
0%
b11 *
0-
02
b11 6
#702630000000
1!
1%
1-
12
15
#702640000000
0!
0%
b100 *
0-
02
b100 6
#702650000000
1!
1%
1-
12
#702660000000
0!
0%
b101 *
0-
02
b101 6
#702670000000
1!
1%
1-
12
#702680000000
0!
0%
b110 *
0-
02
b110 6
#702690000000
1!
1%
1-
12
#702700000000
0!
0%
b111 *
0-
02
b111 6
#702710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#702720000000
0!
0%
b0 *
0-
02
b0 6
#702730000000
1!
1%
1-
12
#702740000000
0!
0%
b1 *
0-
02
b1 6
#702750000000
1!
1%
1-
12
#702760000000
0!
0%
b10 *
0-
02
b10 6
#702770000000
1!
1%
1-
12
#702780000000
0!
0%
b11 *
0-
02
b11 6
#702790000000
1!
1%
1-
12
15
#702800000000
0!
0%
b100 *
0-
02
b100 6
#702810000000
1!
1%
1-
12
#702820000000
0!
0%
b101 *
0-
02
b101 6
#702830000000
1!
1%
1-
12
#702840000000
0!
0%
b110 *
0-
02
b110 6
#702850000000
1!
1%
1-
12
#702860000000
0!
0%
b111 *
0-
02
b111 6
#702870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#702880000000
0!
0%
b0 *
0-
02
b0 6
#702890000000
1!
1%
1-
12
#702900000000
0!
0%
b1 *
0-
02
b1 6
#702910000000
1!
1%
1-
12
#702920000000
0!
0%
b10 *
0-
02
b10 6
#702930000000
1!
1%
1-
12
#702940000000
0!
0%
b11 *
0-
02
b11 6
#702950000000
1!
1%
1-
12
15
#702960000000
0!
0%
b100 *
0-
02
b100 6
#702970000000
1!
1%
1-
12
#702980000000
0!
0%
b101 *
0-
02
b101 6
#702990000000
1!
1%
1-
12
#703000000000
0!
0%
b110 *
0-
02
b110 6
#703010000000
1!
1%
1-
12
#703020000000
0!
0%
b111 *
0-
02
b111 6
#703030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#703040000000
0!
0%
b0 *
0-
02
b0 6
#703050000000
1!
1%
1-
12
#703060000000
0!
0%
b1 *
0-
02
b1 6
#703070000000
1!
1%
1-
12
#703080000000
0!
0%
b10 *
0-
02
b10 6
#703090000000
1!
1%
1-
12
#703100000000
0!
0%
b11 *
0-
02
b11 6
#703110000000
1!
1%
1-
12
15
#703120000000
0!
0%
b100 *
0-
02
b100 6
#703130000000
1!
1%
1-
12
#703140000000
0!
0%
b101 *
0-
02
b101 6
#703150000000
1!
1%
1-
12
#703160000000
0!
0%
b110 *
0-
02
b110 6
#703170000000
1!
1%
1-
12
#703180000000
0!
0%
b111 *
0-
02
b111 6
#703190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#703200000000
0!
0%
b0 *
0-
02
b0 6
#703210000000
1!
1%
1-
12
#703220000000
0!
0%
b1 *
0-
02
b1 6
#703230000000
1!
1%
1-
12
#703240000000
0!
0%
b10 *
0-
02
b10 6
#703250000000
1!
1%
1-
12
#703260000000
0!
0%
b11 *
0-
02
b11 6
#703270000000
1!
1%
1-
12
15
#703280000000
0!
0%
b100 *
0-
02
b100 6
#703290000000
1!
1%
1-
12
#703300000000
0!
0%
b101 *
0-
02
b101 6
#703310000000
1!
1%
1-
12
#703320000000
0!
0%
b110 *
0-
02
b110 6
#703330000000
1!
1%
1-
12
#703340000000
0!
0%
b111 *
0-
02
b111 6
#703350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#703360000000
0!
0%
b0 *
0-
02
b0 6
#703370000000
1!
1%
1-
12
#703380000000
0!
0%
b1 *
0-
02
b1 6
#703390000000
1!
1%
1-
12
#703400000000
0!
0%
b10 *
0-
02
b10 6
#703410000000
1!
1%
1-
12
#703420000000
0!
0%
b11 *
0-
02
b11 6
#703430000000
1!
1%
1-
12
15
#703440000000
0!
0%
b100 *
0-
02
b100 6
#703450000000
1!
1%
1-
12
#703460000000
0!
0%
b101 *
0-
02
b101 6
#703470000000
1!
1%
1-
12
#703480000000
0!
0%
b110 *
0-
02
b110 6
#703490000000
1!
1%
1-
12
#703500000000
0!
0%
b111 *
0-
02
b111 6
#703510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#703520000000
0!
0%
b0 *
0-
02
b0 6
#703530000000
1!
1%
1-
12
#703540000000
0!
0%
b1 *
0-
02
b1 6
#703550000000
1!
1%
1-
12
#703560000000
0!
0%
b10 *
0-
02
b10 6
#703570000000
1!
1%
1-
12
#703580000000
0!
0%
b11 *
0-
02
b11 6
#703590000000
1!
1%
1-
12
15
#703600000000
0!
0%
b100 *
0-
02
b100 6
#703610000000
1!
1%
1-
12
#703620000000
0!
0%
b101 *
0-
02
b101 6
#703630000000
1!
1%
1-
12
#703640000000
0!
0%
b110 *
0-
02
b110 6
#703650000000
1!
1%
1-
12
#703660000000
0!
0%
b111 *
0-
02
b111 6
#703670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#703680000000
0!
0%
b0 *
0-
02
b0 6
#703690000000
1!
1%
1-
12
#703700000000
0!
0%
b1 *
0-
02
b1 6
#703710000000
1!
1%
1-
12
#703720000000
0!
0%
b10 *
0-
02
b10 6
#703730000000
1!
1%
1-
12
#703740000000
0!
0%
b11 *
0-
02
b11 6
#703750000000
1!
1%
1-
12
15
#703760000000
0!
0%
b100 *
0-
02
b100 6
#703770000000
1!
1%
1-
12
#703780000000
0!
0%
b101 *
0-
02
b101 6
#703790000000
1!
1%
1-
12
#703800000000
0!
0%
b110 *
0-
02
b110 6
#703810000000
1!
1%
1-
12
#703820000000
0!
0%
b111 *
0-
02
b111 6
#703830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#703840000000
0!
0%
b0 *
0-
02
b0 6
#703850000000
1!
1%
1-
12
#703860000000
0!
0%
b1 *
0-
02
b1 6
#703870000000
1!
1%
1-
12
#703880000000
0!
0%
b10 *
0-
02
b10 6
#703890000000
1!
1%
1-
12
#703900000000
0!
0%
b11 *
0-
02
b11 6
#703910000000
1!
1%
1-
12
15
#703920000000
0!
0%
b100 *
0-
02
b100 6
#703930000000
1!
1%
1-
12
#703940000000
0!
0%
b101 *
0-
02
b101 6
#703950000000
1!
1%
1-
12
#703960000000
0!
0%
b110 *
0-
02
b110 6
#703970000000
1!
1%
1-
12
#703980000000
0!
0%
b111 *
0-
02
b111 6
#703990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#704000000000
0!
0%
b0 *
0-
02
b0 6
#704010000000
1!
1%
1-
12
#704020000000
0!
0%
b1 *
0-
02
b1 6
#704030000000
1!
1%
1-
12
#704040000000
0!
0%
b10 *
0-
02
b10 6
#704050000000
1!
1%
1-
12
#704060000000
0!
0%
b11 *
0-
02
b11 6
#704070000000
1!
1%
1-
12
15
#704080000000
0!
0%
b100 *
0-
02
b100 6
#704090000000
1!
1%
1-
12
#704100000000
0!
0%
b101 *
0-
02
b101 6
#704110000000
1!
1%
1-
12
#704120000000
0!
0%
b110 *
0-
02
b110 6
#704130000000
1!
1%
1-
12
#704140000000
0!
0%
b111 *
0-
02
b111 6
#704150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#704160000000
0!
0%
b0 *
0-
02
b0 6
#704170000000
1!
1%
1-
12
#704180000000
0!
0%
b1 *
0-
02
b1 6
#704190000000
1!
1%
1-
12
#704200000000
0!
0%
b10 *
0-
02
b10 6
#704210000000
1!
1%
1-
12
#704220000000
0!
0%
b11 *
0-
02
b11 6
#704230000000
1!
1%
1-
12
15
#704240000000
0!
0%
b100 *
0-
02
b100 6
#704250000000
1!
1%
1-
12
#704260000000
0!
0%
b101 *
0-
02
b101 6
#704270000000
1!
1%
1-
12
#704280000000
0!
0%
b110 *
0-
02
b110 6
#704290000000
1!
1%
1-
12
#704300000000
0!
0%
b111 *
0-
02
b111 6
#704310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#704320000000
0!
0%
b0 *
0-
02
b0 6
#704330000000
1!
1%
1-
12
#704340000000
0!
0%
b1 *
0-
02
b1 6
#704350000000
1!
1%
1-
12
#704360000000
0!
0%
b10 *
0-
02
b10 6
#704370000000
1!
1%
1-
12
#704380000000
0!
0%
b11 *
0-
02
b11 6
#704390000000
1!
1%
1-
12
15
#704400000000
0!
0%
b100 *
0-
02
b100 6
#704410000000
1!
1%
1-
12
#704420000000
0!
0%
b101 *
0-
02
b101 6
#704430000000
1!
1%
1-
12
#704440000000
0!
0%
b110 *
0-
02
b110 6
#704450000000
1!
1%
1-
12
#704460000000
0!
0%
b111 *
0-
02
b111 6
#704470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#704480000000
0!
0%
b0 *
0-
02
b0 6
#704490000000
1!
1%
1-
12
#704500000000
0!
0%
b1 *
0-
02
b1 6
#704510000000
1!
1%
1-
12
#704520000000
0!
0%
b10 *
0-
02
b10 6
#704530000000
1!
1%
1-
12
#704540000000
0!
0%
b11 *
0-
02
b11 6
#704550000000
1!
1%
1-
12
15
#704560000000
0!
0%
b100 *
0-
02
b100 6
#704570000000
1!
1%
1-
12
#704580000000
0!
0%
b101 *
0-
02
b101 6
#704590000000
1!
1%
1-
12
#704600000000
0!
0%
b110 *
0-
02
b110 6
#704610000000
1!
1%
1-
12
#704620000000
0!
0%
b111 *
0-
02
b111 6
#704630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#704640000000
0!
0%
b0 *
0-
02
b0 6
#704650000000
1!
1%
1-
12
#704660000000
0!
0%
b1 *
0-
02
b1 6
#704670000000
1!
1%
1-
12
#704680000000
0!
0%
b10 *
0-
02
b10 6
#704690000000
1!
1%
1-
12
#704700000000
0!
0%
b11 *
0-
02
b11 6
#704710000000
1!
1%
1-
12
15
#704720000000
0!
0%
b100 *
0-
02
b100 6
#704730000000
1!
1%
1-
12
#704740000000
0!
0%
b101 *
0-
02
b101 6
#704750000000
1!
1%
1-
12
#704760000000
0!
0%
b110 *
0-
02
b110 6
#704770000000
1!
1%
1-
12
#704780000000
0!
0%
b111 *
0-
02
b111 6
#704790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#704800000000
0!
0%
b0 *
0-
02
b0 6
#704810000000
1!
1%
1-
12
#704820000000
0!
0%
b1 *
0-
02
b1 6
#704830000000
1!
1%
1-
12
#704840000000
0!
0%
b10 *
0-
02
b10 6
#704850000000
1!
1%
1-
12
#704860000000
0!
0%
b11 *
0-
02
b11 6
#704870000000
1!
1%
1-
12
15
#704880000000
0!
0%
b100 *
0-
02
b100 6
#704890000000
1!
1%
1-
12
#704900000000
0!
0%
b101 *
0-
02
b101 6
#704910000000
1!
1%
1-
12
#704920000000
0!
0%
b110 *
0-
02
b110 6
#704930000000
1!
1%
1-
12
#704940000000
0!
0%
b111 *
0-
02
b111 6
#704950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#704960000000
0!
0%
b0 *
0-
02
b0 6
#704970000000
1!
1%
1-
12
#704980000000
0!
0%
b1 *
0-
02
b1 6
#704990000000
1!
1%
1-
12
#705000000000
0!
0%
b10 *
0-
02
b10 6
#705010000000
1!
1%
1-
12
#705020000000
0!
0%
b11 *
0-
02
b11 6
#705030000000
1!
1%
1-
12
15
#705040000000
0!
0%
b100 *
0-
02
b100 6
#705050000000
1!
1%
1-
12
#705060000000
0!
0%
b101 *
0-
02
b101 6
#705070000000
1!
1%
1-
12
#705080000000
0!
0%
b110 *
0-
02
b110 6
#705090000000
1!
1%
1-
12
#705100000000
0!
0%
b111 *
0-
02
b111 6
#705110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#705120000000
0!
0%
b0 *
0-
02
b0 6
#705130000000
1!
1%
1-
12
#705140000000
0!
0%
b1 *
0-
02
b1 6
#705150000000
1!
1%
1-
12
#705160000000
0!
0%
b10 *
0-
02
b10 6
#705170000000
1!
1%
1-
12
#705180000000
0!
0%
b11 *
0-
02
b11 6
#705190000000
1!
1%
1-
12
15
#705200000000
0!
0%
b100 *
0-
02
b100 6
#705210000000
1!
1%
1-
12
#705220000000
0!
0%
b101 *
0-
02
b101 6
#705230000000
1!
1%
1-
12
#705240000000
0!
0%
b110 *
0-
02
b110 6
#705250000000
1!
1%
1-
12
#705260000000
0!
0%
b111 *
0-
02
b111 6
#705270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#705280000000
0!
0%
b0 *
0-
02
b0 6
#705290000000
1!
1%
1-
12
#705300000000
0!
0%
b1 *
0-
02
b1 6
#705310000000
1!
1%
1-
12
#705320000000
0!
0%
b10 *
0-
02
b10 6
#705330000000
1!
1%
1-
12
#705340000000
0!
0%
b11 *
0-
02
b11 6
#705350000000
1!
1%
1-
12
15
#705360000000
0!
0%
b100 *
0-
02
b100 6
#705370000000
1!
1%
1-
12
#705380000000
0!
0%
b101 *
0-
02
b101 6
#705390000000
1!
1%
1-
12
#705400000000
0!
0%
b110 *
0-
02
b110 6
#705410000000
1!
1%
1-
12
#705420000000
0!
0%
b111 *
0-
02
b111 6
#705430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#705440000000
0!
0%
b0 *
0-
02
b0 6
#705450000000
1!
1%
1-
12
#705460000000
0!
0%
b1 *
0-
02
b1 6
#705470000000
1!
1%
1-
12
#705480000000
0!
0%
b10 *
0-
02
b10 6
#705490000000
1!
1%
1-
12
#705500000000
0!
0%
b11 *
0-
02
b11 6
#705510000000
1!
1%
1-
12
15
#705520000000
0!
0%
b100 *
0-
02
b100 6
#705530000000
1!
1%
1-
12
#705540000000
0!
0%
b101 *
0-
02
b101 6
#705550000000
1!
1%
1-
12
#705560000000
0!
0%
b110 *
0-
02
b110 6
#705570000000
1!
1%
1-
12
#705580000000
0!
0%
b111 *
0-
02
b111 6
#705590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#705600000000
0!
0%
b0 *
0-
02
b0 6
#705610000000
1!
1%
1-
12
#705620000000
0!
0%
b1 *
0-
02
b1 6
#705630000000
1!
1%
1-
12
#705640000000
0!
0%
b10 *
0-
02
b10 6
#705650000000
1!
1%
1-
12
#705660000000
0!
0%
b11 *
0-
02
b11 6
#705670000000
1!
1%
1-
12
15
#705680000000
0!
0%
b100 *
0-
02
b100 6
#705690000000
1!
1%
1-
12
#705700000000
0!
0%
b101 *
0-
02
b101 6
#705710000000
1!
1%
1-
12
#705720000000
0!
0%
b110 *
0-
02
b110 6
#705730000000
1!
1%
1-
12
#705740000000
0!
0%
b111 *
0-
02
b111 6
#705750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#705760000000
0!
0%
b0 *
0-
02
b0 6
#705770000000
1!
1%
1-
12
#705780000000
0!
0%
b1 *
0-
02
b1 6
#705790000000
1!
1%
1-
12
#705800000000
0!
0%
b10 *
0-
02
b10 6
#705810000000
1!
1%
1-
12
#705820000000
0!
0%
b11 *
0-
02
b11 6
#705830000000
1!
1%
1-
12
15
#705840000000
0!
0%
b100 *
0-
02
b100 6
#705850000000
1!
1%
1-
12
#705860000000
0!
0%
b101 *
0-
02
b101 6
#705870000000
1!
1%
1-
12
#705880000000
0!
0%
b110 *
0-
02
b110 6
#705890000000
1!
1%
1-
12
#705900000000
0!
0%
b111 *
0-
02
b111 6
#705910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#705920000000
0!
0%
b0 *
0-
02
b0 6
#705930000000
1!
1%
1-
12
#705940000000
0!
0%
b1 *
0-
02
b1 6
#705950000000
1!
1%
1-
12
#705960000000
0!
0%
b10 *
0-
02
b10 6
#705970000000
1!
1%
1-
12
#705980000000
0!
0%
b11 *
0-
02
b11 6
#705990000000
1!
1%
1-
12
15
#706000000000
0!
0%
b100 *
0-
02
b100 6
#706010000000
1!
1%
1-
12
#706020000000
0!
0%
b101 *
0-
02
b101 6
#706030000000
1!
1%
1-
12
#706040000000
0!
0%
b110 *
0-
02
b110 6
#706050000000
1!
1%
1-
12
#706060000000
0!
0%
b111 *
0-
02
b111 6
#706070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#706080000000
0!
0%
b0 *
0-
02
b0 6
#706090000000
1!
1%
1-
12
#706100000000
0!
0%
b1 *
0-
02
b1 6
#706110000000
1!
1%
1-
12
#706120000000
0!
0%
b10 *
0-
02
b10 6
#706130000000
1!
1%
1-
12
#706140000000
0!
0%
b11 *
0-
02
b11 6
#706150000000
1!
1%
1-
12
15
#706160000000
0!
0%
b100 *
0-
02
b100 6
#706170000000
1!
1%
1-
12
#706180000000
0!
0%
b101 *
0-
02
b101 6
#706190000000
1!
1%
1-
12
#706200000000
0!
0%
b110 *
0-
02
b110 6
#706210000000
1!
1%
1-
12
#706220000000
0!
0%
b111 *
0-
02
b111 6
#706230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#706240000000
0!
0%
b0 *
0-
02
b0 6
#706250000000
1!
1%
1-
12
#706260000000
0!
0%
b1 *
0-
02
b1 6
#706270000000
1!
1%
1-
12
#706280000000
0!
0%
b10 *
0-
02
b10 6
#706290000000
1!
1%
1-
12
#706300000000
0!
0%
b11 *
0-
02
b11 6
#706310000000
1!
1%
1-
12
15
#706320000000
0!
0%
b100 *
0-
02
b100 6
#706330000000
1!
1%
1-
12
#706340000000
0!
0%
b101 *
0-
02
b101 6
#706350000000
1!
1%
1-
12
#706360000000
0!
0%
b110 *
0-
02
b110 6
#706370000000
1!
1%
1-
12
#706380000000
0!
0%
b111 *
0-
02
b111 6
#706390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#706400000000
0!
0%
b0 *
0-
02
b0 6
#706410000000
1!
1%
1-
12
#706420000000
0!
0%
b1 *
0-
02
b1 6
#706430000000
1!
1%
1-
12
#706440000000
0!
0%
b10 *
0-
02
b10 6
#706450000000
1!
1%
1-
12
#706460000000
0!
0%
b11 *
0-
02
b11 6
#706470000000
1!
1%
1-
12
15
#706480000000
0!
0%
b100 *
0-
02
b100 6
#706490000000
1!
1%
1-
12
#706500000000
0!
0%
b101 *
0-
02
b101 6
#706510000000
1!
1%
1-
12
#706520000000
0!
0%
b110 *
0-
02
b110 6
#706530000000
1!
1%
1-
12
#706540000000
0!
0%
b111 *
0-
02
b111 6
#706550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#706560000000
0!
0%
b0 *
0-
02
b0 6
#706570000000
1!
1%
1-
12
#706580000000
0!
0%
b1 *
0-
02
b1 6
#706590000000
1!
1%
1-
12
#706600000000
0!
0%
b10 *
0-
02
b10 6
#706610000000
1!
1%
1-
12
#706620000000
0!
0%
b11 *
0-
02
b11 6
#706630000000
1!
1%
1-
12
15
#706640000000
0!
0%
b100 *
0-
02
b100 6
#706650000000
1!
1%
1-
12
#706660000000
0!
0%
b101 *
0-
02
b101 6
#706670000000
1!
1%
1-
12
#706680000000
0!
0%
b110 *
0-
02
b110 6
#706690000000
1!
1%
1-
12
#706700000000
0!
0%
b111 *
0-
02
b111 6
#706710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#706720000000
0!
0%
b0 *
0-
02
b0 6
#706730000000
1!
1%
1-
12
#706740000000
0!
0%
b1 *
0-
02
b1 6
#706750000000
1!
1%
1-
12
#706760000000
0!
0%
b10 *
0-
02
b10 6
#706770000000
1!
1%
1-
12
#706780000000
0!
0%
b11 *
0-
02
b11 6
#706790000000
1!
1%
1-
12
15
#706800000000
0!
0%
b100 *
0-
02
b100 6
#706810000000
1!
1%
1-
12
#706820000000
0!
0%
b101 *
0-
02
b101 6
#706830000000
1!
1%
1-
12
#706840000000
0!
0%
b110 *
0-
02
b110 6
#706850000000
1!
1%
1-
12
#706860000000
0!
0%
b111 *
0-
02
b111 6
#706870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#706880000000
0!
0%
b0 *
0-
02
b0 6
#706890000000
1!
1%
1-
12
#706900000000
0!
0%
b1 *
0-
02
b1 6
#706910000000
1!
1%
1-
12
#706920000000
0!
0%
b10 *
0-
02
b10 6
#706930000000
1!
1%
1-
12
#706940000000
0!
0%
b11 *
0-
02
b11 6
#706950000000
1!
1%
1-
12
15
#706960000000
0!
0%
b100 *
0-
02
b100 6
#706970000000
1!
1%
1-
12
#706980000000
0!
0%
b101 *
0-
02
b101 6
#706990000000
1!
1%
1-
12
#707000000000
0!
0%
b110 *
0-
02
b110 6
#707010000000
1!
1%
1-
12
#707020000000
0!
0%
b111 *
0-
02
b111 6
#707030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#707040000000
0!
0%
b0 *
0-
02
b0 6
#707050000000
1!
1%
1-
12
#707060000000
0!
0%
b1 *
0-
02
b1 6
#707070000000
1!
1%
1-
12
#707080000000
0!
0%
b10 *
0-
02
b10 6
#707090000000
1!
1%
1-
12
#707100000000
0!
0%
b11 *
0-
02
b11 6
#707110000000
1!
1%
1-
12
15
#707120000000
0!
0%
b100 *
0-
02
b100 6
#707130000000
1!
1%
1-
12
#707140000000
0!
0%
b101 *
0-
02
b101 6
#707150000000
1!
1%
1-
12
#707160000000
0!
0%
b110 *
0-
02
b110 6
#707170000000
1!
1%
1-
12
#707180000000
0!
0%
b111 *
0-
02
b111 6
#707190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#707200000000
0!
0%
b0 *
0-
02
b0 6
#707210000000
1!
1%
1-
12
#707220000000
0!
0%
b1 *
0-
02
b1 6
#707230000000
1!
1%
1-
12
#707240000000
0!
0%
b10 *
0-
02
b10 6
#707250000000
1!
1%
1-
12
#707260000000
0!
0%
b11 *
0-
02
b11 6
#707270000000
1!
1%
1-
12
15
#707280000000
0!
0%
b100 *
0-
02
b100 6
#707290000000
1!
1%
1-
12
#707300000000
0!
0%
b101 *
0-
02
b101 6
#707310000000
1!
1%
1-
12
#707320000000
0!
0%
b110 *
0-
02
b110 6
#707330000000
1!
1%
1-
12
#707340000000
0!
0%
b111 *
0-
02
b111 6
#707350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#707360000000
0!
0%
b0 *
0-
02
b0 6
#707370000000
1!
1%
1-
12
#707380000000
0!
0%
b1 *
0-
02
b1 6
#707390000000
1!
1%
1-
12
#707400000000
0!
0%
b10 *
0-
02
b10 6
#707410000000
1!
1%
1-
12
#707420000000
0!
0%
b11 *
0-
02
b11 6
#707430000000
1!
1%
1-
12
15
#707440000000
0!
0%
b100 *
0-
02
b100 6
#707450000000
1!
1%
1-
12
#707460000000
0!
0%
b101 *
0-
02
b101 6
#707470000000
1!
1%
1-
12
#707480000000
0!
0%
b110 *
0-
02
b110 6
#707490000000
1!
1%
1-
12
#707500000000
0!
0%
b111 *
0-
02
b111 6
#707510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#707520000000
0!
0%
b0 *
0-
02
b0 6
#707530000000
1!
1%
1-
12
#707540000000
0!
0%
b1 *
0-
02
b1 6
#707550000000
1!
1%
1-
12
#707560000000
0!
0%
b10 *
0-
02
b10 6
#707570000000
1!
1%
1-
12
#707580000000
0!
0%
b11 *
0-
02
b11 6
#707590000000
1!
1%
1-
12
15
#707600000000
0!
0%
b100 *
0-
02
b100 6
#707610000000
1!
1%
1-
12
#707620000000
0!
0%
b101 *
0-
02
b101 6
#707630000000
1!
1%
1-
12
#707640000000
0!
0%
b110 *
0-
02
b110 6
#707650000000
1!
1%
1-
12
#707660000000
0!
0%
b111 *
0-
02
b111 6
#707670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#707680000000
0!
0%
b0 *
0-
02
b0 6
#707690000000
1!
1%
1-
12
#707700000000
0!
0%
b1 *
0-
02
b1 6
#707710000000
1!
1%
1-
12
#707720000000
0!
0%
b10 *
0-
02
b10 6
#707730000000
1!
1%
1-
12
#707740000000
0!
0%
b11 *
0-
02
b11 6
#707750000000
1!
1%
1-
12
15
#707760000000
0!
0%
b100 *
0-
02
b100 6
#707770000000
1!
1%
1-
12
#707780000000
0!
0%
b101 *
0-
02
b101 6
#707790000000
1!
1%
1-
12
#707800000000
0!
0%
b110 *
0-
02
b110 6
#707810000000
1!
1%
1-
12
#707820000000
0!
0%
b111 *
0-
02
b111 6
#707830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#707840000000
0!
0%
b0 *
0-
02
b0 6
#707850000000
1!
1%
1-
12
#707860000000
0!
0%
b1 *
0-
02
b1 6
#707870000000
1!
1%
1-
12
#707880000000
0!
0%
b10 *
0-
02
b10 6
#707890000000
1!
1%
1-
12
#707900000000
0!
0%
b11 *
0-
02
b11 6
#707910000000
1!
1%
1-
12
15
#707920000000
0!
0%
b100 *
0-
02
b100 6
#707930000000
1!
1%
1-
12
#707940000000
0!
0%
b101 *
0-
02
b101 6
#707950000000
1!
1%
1-
12
#707960000000
0!
0%
b110 *
0-
02
b110 6
#707970000000
1!
1%
1-
12
#707980000000
0!
0%
b111 *
0-
02
b111 6
#707990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#708000000000
0!
0%
b0 *
0-
02
b0 6
#708010000000
1!
1%
1-
12
#708020000000
0!
0%
b1 *
0-
02
b1 6
#708030000000
1!
1%
1-
12
#708040000000
0!
0%
b10 *
0-
02
b10 6
#708050000000
1!
1%
1-
12
#708060000000
0!
0%
b11 *
0-
02
b11 6
#708070000000
1!
1%
1-
12
15
#708080000000
0!
0%
b100 *
0-
02
b100 6
#708090000000
1!
1%
1-
12
#708100000000
0!
0%
b101 *
0-
02
b101 6
#708110000000
1!
1%
1-
12
#708120000000
0!
0%
b110 *
0-
02
b110 6
#708130000000
1!
1%
1-
12
#708140000000
0!
0%
b111 *
0-
02
b111 6
#708150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#708160000000
0!
0%
b0 *
0-
02
b0 6
#708170000000
1!
1%
1-
12
#708180000000
0!
0%
b1 *
0-
02
b1 6
#708190000000
1!
1%
1-
12
#708200000000
0!
0%
b10 *
0-
02
b10 6
#708210000000
1!
1%
1-
12
#708220000000
0!
0%
b11 *
0-
02
b11 6
#708230000000
1!
1%
1-
12
15
#708240000000
0!
0%
b100 *
0-
02
b100 6
#708250000000
1!
1%
1-
12
#708260000000
0!
0%
b101 *
0-
02
b101 6
#708270000000
1!
1%
1-
12
#708280000000
0!
0%
b110 *
0-
02
b110 6
#708290000000
1!
1%
1-
12
#708300000000
0!
0%
b111 *
0-
02
b111 6
#708310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#708320000000
0!
0%
b0 *
0-
02
b0 6
#708330000000
1!
1%
1-
12
#708340000000
0!
0%
b1 *
0-
02
b1 6
#708350000000
1!
1%
1-
12
#708360000000
0!
0%
b10 *
0-
02
b10 6
#708370000000
1!
1%
1-
12
#708380000000
0!
0%
b11 *
0-
02
b11 6
#708390000000
1!
1%
1-
12
15
#708400000000
0!
0%
b100 *
0-
02
b100 6
#708410000000
1!
1%
1-
12
#708420000000
0!
0%
b101 *
0-
02
b101 6
#708430000000
1!
1%
1-
12
#708440000000
0!
0%
b110 *
0-
02
b110 6
#708450000000
1!
1%
1-
12
#708460000000
0!
0%
b111 *
0-
02
b111 6
#708470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#708480000000
0!
0%
b0 *
0-
02
b0 6
#708490000000
1!
1%
1-
12
#708500000000
0!
0%
b1 *
0-
02
b1 6
#708510000000
1!
1%
1-
12
#708520000000
0!
0%
b10 *
0-
02
b10 6
#708530000000
1!
1%
1-
12
#708540000000
0!
0%
b11 *
0-
02
b11 6
#708550000000
1!
1%
1-
12
15
#708560000000
0!
0%
b100 *
0-
02
b100 6
#708570000000
1!
1%
1-
12
#708580000000
0!
0%
b101 *
0-
02
b101 6
#708590000000
1!
1%
1-
12
#708600000000
0!
0%
b110 *
0-
02
b110 6
#708610000000
1!
1%
1-
12
#708620000000
0!
0%
b111 *
0-
02
b111 6
#708630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#708640000000
0!
0%
b0 *
0-
02
b0 6
#708650000000
1!
1%
1-
12
#708660000000
0!
0%
b1 *
0-
02
b1 6
#708670000000
1!
1%
1-
12
#708680000000
0!
0%
b10 *
0-
02
b10 6
#708690000000
1!
1%
1-
12
#708700000000
0!
0%
b11 *
0-
02
b11 6
#708710000000
1!
1%
1-
12
15
#708720000000
0!
0%
b100 *
0-
02
b100 6
#708730000000
1!
1%
1-
12
#708740000000
0!
0%
b101 *
0-
02
b101 6
#708750000000
1!
1%
1-
12
#708760000000
0!
0%
b110 *
0-
02
b110 6
#708770000000
1!
1%
1-
12
#708780000000
0!
0%
b111 *
0-
02
b111 6
#708790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#708800000000
0!
0%
b0 *
0-
02
b0 6
#708810000000
1!
1%
1-
12
#708820000000
0!
0%
b1 *
0-
02
b1 6
#708830000000
1!
1%
1-
12
#708840000000
0!
0%
b10 *
0-
02
b10 6
#708850000000
1!
1%
1-
12
#708860000000
0!
0%
b11 *
0-
02
b11 6
#708870000000
1!
1%
1-
12
15
#708880000000
0!
0%
b100 *
0-
02
b100 6
#708890000000
1!
1%
1-
12
#708900000000
0!
0%
b101 *
0-
02
b101 6
#708910000000
1!
1%
1-
12
#708920000000
0!
0%
b110 *
0-
02
b110 6
#708930000000
1!
1%
1-
12
#708940000000
0!
0%
b111 *
0-
02
b111 6
#708950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#708960000000
0!
0%
b0 *
0-
02
b0 6
#708970000000
1!
1%
1-
12
#708980000000
0!
0%
b1 *
0-
02
b1 6
#708990000000
1!
1%
1-
12
#709000000000
0!
0%
b10 *
0-
02
b10 6
#709010000000
1!
1%
1-
12
#709020000000
0!
0%
b11 *
0-
02
b11 6
#709030000000
1!
1%
1-
12
15
#709040000000
0!
0%
b100 *
0-
02
b100 6
#709050000000
1!
1%
1-
12
#709060000000
0!
0%
b101 *
0-
02
b101 6
#709070000000
1!
1%
1-
12
#709080000000
0!
0%
b110 *
0-
02
b110 6
#709090000000
1!
1%
1-
12
#709100000000
0!
0%
b111 *
0-
02
b111 6
#709110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#709120000000
0!
0%
b0 *
0-
02
b0 6
#709130000000
1!
1%
1-
12
#709140000000
0!
0%
b1 *
0-
02
b1 6
#709150000000
1!
1%
1-
12
#709160000000
0!
0%
b10 *
0-
02
b10 6
#709170000000
1!
1%
1-
12
#709180000000
0!
0%
b11 *
0-
02
b11 6
#709190000000
1!
1%
1-
12
15
#709200000000
0!
0%
b100 *
0-
02
b100 6
#709210000000
1!
1%
1-
12
#709220000000
0!
0%
b101 *
0-
02
b101 6
#709230000000
1!
1%
1-
12
#709240000000
0!
0%
b110 *
0-
02
b110 6
#709250000000
1!
1%
1-
12
#709260000000
0!
0%
b111 *
0-
02
b111 6
#709270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#709280000000
0!
0%
b0 *
0-
02
b0 6
#709290000000
1!
1%
1-
12
#709300000000
0!
0%
b1 *
0-
02
b1 6
#709310000000
1!
1%
1-
12
#709320000000
0!
0%
b10 *
0-
02
b10 6
#709330000000
1!
1%
1-
12
#709340000000
0!
0%
b11 *
0-
02
b11 6
#709350000000
1!
1%
1-
12
15
#709360000000
0!
0%
b100 *
0-
02
b100 6
#709370000000
1!
1%
1-
12
#709380000000
0!
0%
b101 *
0-
02
b101 6
#709390000000
1!
1%
1-
12
#709400000000
0!
0%
b110 *
0-
02
b110 6
#709410000000
1!
1%
1-
12
#709420000000
0!
0%
b111 *
0-
02
b111 6
#709430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#709440000000
0!
0%
b0 *
0-
02
b0 6
#709450000000
1!
1%
1-
12
#709460000000
0!
0%
b1 *
0-
02
b1 6
#709470000000
1!
1%
1-
12
#709480000000
0!
0%
b10 *
0-
02
b10 6
#709490000000
1!
1%
1-
12
#709500000000
0!
0%
b11 *
0-
02
b11 6
#709510000000
1!
1%
1-
12
15
#709520000000
0!
0%
b100 *
0-
02
b100 6
#709530000000
1!
1%
1-
12
#709540000000
0!
0%
b101 *
0-
02
b101 6
#709550000000
1!
1%
1-
12
#709560000000
0!
0%
b110 *
0-
02
b110 6
#709570000000
1!
1%
1-
12
#709580000000
0!
0%
b111 *
0-
02
b111 6
#709590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#709600000000
0!
0%
b0 *
0-
02
b0 6
#709610000000
1!
1%
1-
12
#709620000000
0!
0%
b1 *
0-
02
b1 6
#709630000000
1!
1%
1-
12
#709640000000
0!
0%
b10 *
0-
02
b10 6
#709650000000
1!
1%
1-
12
#709660000000
0!
0%
b11 *
0-
02
b11 6
#709670000000
1!
1%
1-
12
15
#709680000000
0!
0%
b100 *
0-
02
b100 6
#709690000000
1!
1%
1-
12
#709700000000
0!
0%
b101 *
0-
02
b101 6
#709710000000
1!
1%
1-
12
#709720000000
0!
0%
b110 *
0-
02
b110 6
#709730000000
1!
1%
1-
12
#709740000000
0!
0%
b111 *
0-
02
b111 6
#709750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#709760000000
0!
0%
b0 *
0-
02
b0 6
#709770000000
1!
1%
1-
12
#709780000000
0!
0%
b1 *
0-
02
b1 6
#709790000000
1!
1%
1-
12
#709800000000
0!
0%
b10 *
0-
02
b10 6
#709810000000
1!
1%
1-
12
#709820000000
0!
0%
b11 *
0-
02
b11 6
#709830000000
1!
1%
1-
12
15
#709840000000
0!
0%
b100 *
0-
02
b100 6
#709850000000
1!
1%
1-
12
#709860000000
0!
0%
b101 *
0-
02
b101 6
#709870000000
1!
1%
1-
12
#709880000000
0!
0%
b110 *
0-
02
b110 6
#709890000000
1!
1%
1-
12
#709900000000
0!
0%
b111 *
0-
02
b111 6
#709910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#709920000000
0!
0%
b0 *
0-
02
b0 6
#709930000000
1!
1%
1-
12
#709940000000
0!
0%
b1 *
0-
02
b1 6
#709950000000
1!
1%
1-
12
#709960000000
0!
0%
b10 *
0-
02
b10 6
#709970000000
1!
1%
1-
12
#709980000000
0!
0%
b11 *
0-
02
b11 6
#709990000000
1!
1%
1-
12
15
#710000000000
0!
0%
b100 *
0-
02
b100 6
#710010000000
1!
1%
1-
12
#710020000000
0!
0%
b101 *
0-
02
b101 6
#710030000000
1!
1%
1-
12
#710040000000
0!
0%
b110 *
0-
02
b110 6
#710050000000
1!
1%
1-
12
#710060000000
0!
0%
b111 *
0-
02
b111 6
#710070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#710080000000
0!
0%
b0 *
0-
02
b0 6
#710090000000
1!
1%
1-
12
#710100000000
0!
0%
b1 *
0-
02
b1 6
#710110000000
1!
1%
1-
12
#710120000000
0!
0%
b10 *
0-
02
b10 6
#710130000000
1!
1%
1-
12
#710140000000
0!
0%
b11 *
0-
02
b11 6
#710150000000
1!
1%
1-
12
15
#710160000000
0!
0%
b100 *
0-
02
b100 6
#710170000000
1!
1%
1-
12
#710180000000
0!
0%
b101 *
0-
02
b101 6
#710190000000
1!
1%
1-
12
#710200000000
0!
0%
b110 *
0-
02
b110 6
#710210000000
1!
1%
1-
12
#710220000000
0!
0%
b111 *
0-
02
b111 6
#710230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#710240000000
0!
0%
b0 *
0-
02
b0 6
#710250000000
1!
1%
1-
12
#710260000000
0!
0%
b1 *
0-
02
b1 6
#710270000000
1!
1%
1-
12
#710280000000
0!
0%
b10 *
0-
02
b10 6
#710290000000
1!
1%
1-
12
#710300000000
0!
0%
b11 *
0-
02
b11 6
#710310000000
1!
1%
1-
12
15
#710320000000
0!
0%
b100 *
0-
02
b100 6
#710330000000
1!
1%
1-
12
#710340000000
0!
0%
b101 *
0-
02
b101 6
#710350000000
1!
1%
1-
12
#710360000000
0!
0%
b110 *
0-
02
b110 6
#710370000000
1!
1%
1-
12
#710380000000
0!
0%
b111 *
0-
02
b111 6
#710390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#710400000000
0!
0%
b0 *
0-
02
b0 6
#710410000000
1!
1%
1-
12
#710420000000
0!
0%
b1 *
0-
02
b1 6
#710430000000
1!
1%
1-
12
#710440000000
0!
0%
b10 *
0-
02
b10 6
#710450000000
1!
1%
1-
12
#710460000000
0!
0%
b11 *
0-
02
b11 6
#710470000000
1!
1%
1-
12
15
#710480000000
0!
0%
b100 *
0-
02
b100 6
#710490000000
1!
1%
1-
12
#710500000000
0!
0%
b101 *
0-
02
b101 6
#710510000000
1!
1%
1-
12
#710520000000
0!
0%
b110 *
0-
02
b110 6
#710530000000
1!
1%
1-
12
#710540000000
0!
0%
b111 *
0-
02
b111 6
#710550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#710560000000
0!
0%
b0 *
0-
02
b0 6
#710570000000
1!
1%
1-
12
#710580000000
0!
0%
b1 *
0-
02
b1 6
#710590000000
1!
1%
1-
12
#710600000000
0!
0%
b10 *
0-
02
b10 6
#710610000000
1!
1%
1-
12
#710620000000
0!
0%
b11 *
0-
02
b11 6
#710630000000
1!
1%
1-
12
15
#710640000000
0!
0%
b100 *
0-
02
b100 6
#710650000000
1!
1%
1-
12
#710660000000
0!
0%
b101 *
0-
02
b101 6
#710670000000
1!
1%
1-
12
#710680000000
0!
0%
b110 *
0-
02
b110 6
#710690000000
1!
1%
1-
12
#710700000000
0!
0%
b111 *
0-
02
b111 6
#710710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#710720000000
0!
0%
b0 *
0-
02
b0 6
#710730000000
1!
1%
1-
12
#710740000000
0!
0%
b1 *
0-
02
b1 6
#710750000000
1!
1%
1-
12
#710760000000
0!
0%
b10 *
0-
02
b10 6
#710770000000
1!
1%
1-
12
#710780000000
0!
0%
b11 *
0-
02
b11 6
#710790000000
1!
1%
1-
12
15
#710800000000
0!
0%
b100 *
0-
02
b100 6
#710810000000
1!
1%
1-
12
#710820000000
0!
0%
b101 *
0-
02
b101 6
#710830000000
1!
1%
1-
12
#710840000000
0!
0%
b110 *
0-
02
b110 6
#710850000000
1!
1%
1-
12
#710860000000
0!
0%
b111 *
0-
02
b111 6
#710870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#710880000000
0!
0%
b0 *
0-
02
b0 6
#710890000000
1!
1%
1-
12
#710900000000
0!
0%
b1 *
0-
02
b1 6
#710910000000
1!
1%
1-
12
#710920000000
0!
0%
b10 *
0-
02
b10 6
#710930000000
1!
1%
1-
12
#710940000000
0!
0%
b11 *
0-
02
b11 6
#710950000000
1!
1%
1-
12
15
#710960000000
0!
0%
b100 *
0-
02
b100 6
#710970000000
1!
1%
1-
12
#710980000000
0!
0%
b101 *
0-
02
b101 6
#710990000000
1!
1%
1-
12
#711000000000
0!
0%
b110 *
0-
02
b110 6
#711010000000
1!
1%
1-
12
#711020000000
0!
0%
b111 *
0-
02
b111 6
#711030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#711040000000
0!
0%
b0 *
0-
02
b0 6
#711050000000
1!
1%
1-
12
#711060000000
0!
0%
b1 *
0-
02
b1 6
#711070000000
1!
1%
1-
12
#711080000000
0!
0%
b10 *
0-
02
b10 6
#711090000000
1!
1%
1-
12
#711100000000
0!
0%
b11 *
0-
02
b11 6
#711110000000
1!
1%
1-
12
15
#711120000000
0!
0%
b100 *
0-
02
b100 6
#711130000000
1!
1%
1-
12
#711140000000
0!
0%
b101 *
0-
02
b101 6
#711150000000
1!
1%
1-
12
#711160000000
0!
0%
b110 *
0-
02
b110 6
#711170000000
1!
1%
1-
12
#711180000000
0!
0%
b111 *
0-
02
b111 6
#711190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#711200000000
0!
0%
b0 *
0-
02
b0 6
#711210000000
1!
1%
1-
12
#711220000000
0!
0%
b1 *
0-
02
b1 6
#711230000000
1!
1%
1-
12
#711240000000
0!
0%
b10 *
0-
02
b10 6
#711250000000
1!
1%
1-
12
#711260000000
0!
0%
b11 *
0-
02
b11 6
#711270000000
1!
1%
1-
12
15
#711280000000
0!
0%
b100 *
0-
02
b100 6
#711290000000
1!
1%
1-
12
#711300000000
0!
0%
b101 *
0-
02
b101 6
#711310000000
1!
1%
1-
12
#711320000000
0!
0%
b110 *
0-
02
b110 6
#711330000000
1!
1%
1-
12
#711340000000
0!
0%
b111 *
0-
02
b111 6
#711350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#711360000000
0!
0%
b0 *
0-
02
b0 6
#711370000000
1!
1%
1-
12
#711380000000
0!
0%
b1 *
0-
02
b1 6
#711390000000
1!
1%
1-
12
#711400000000
0!
0%
b10 *
0-
02
b10 6
#711410000000
1!
1%
1-
12
#711420000000
0!
0%
b11 *
0-
02
b11 6
#711430000000
1!
1%
1-
12
15
#711440000000
0!
0%
b100 *
0-
02
b100 6
#711450000000
1!
1%
1-
12
#711460000000
0!
0%
b101 *
0-
02
b101 6
#711470000000
1!
1%
1-
12
#711480000000
0!
0%
b110 *
0-
02
b110 6
#711490000000
1!
1%
1-
12
#711500000000
0!
0%
b111 *
0-
02
b111 6
#711510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#711520000000
0!
0%
b0 *
0-
02
b0 6
#711530000000
1!
1%
1-
12
#711540000000
0!
0%
b1 *
0-
02
b1 6
#711550000000
1!
1%
1-
12
#711560000000
0!
0%
b10 *
0-
02
b10 6
#711570000000
1!
1%
1-
12
#711580000000
0!
0%
b11 *
0-
02
b11 6
#711590000000
1!
1%
1-
12
15
#711600000000
0!
0%
b100 *
0-
02
b100 6
#711610000000
1!
1%
1-
12
#711620000000
0!
0%
b101 *
0-
02
b101 6
#711630000000
1!
1%
1-
12
#711640000000
0!
0%
b110 *
0-
02
b110 6
#711650000000
1!
1%
1-
12
#711660000000
0!
0%
b111 *
0-
02
b111 6
#711670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#711680000000
0!
0%
b0 *
0-
02
b0 6
#711690000000
1!
1%
1-
12
#711700000000
0!
0%
b1 *
0-
02
b1 6
#711710000000
1!
1%
1-
12
#711720000000
0!
0%
b10 *
0-
02
b10 6
#711730000000
1!
1%
1-
12
#711740000000
0!
0%
b11 *
0-
02
b11 6
#711750000000
1!
1%
1-
12
15
#711760000000
0!
0%
b100 *
0-
02
b100 6
#711770000000
1!
1%
1-
12
#711780000000
0!
0%
b101 *
0-
02
b101 6
#711790000000
1!
1%
1-
12
#711800000000
0!
0%
b110 *
0-
02
b110 6
#711810000000
1!
1%
1-
12
#711820000000
0!
0%
b111 *
0-
02
b111 6
#711830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#711840000000
0!
0%
b0 *
0-
02
b0 6
#711850000000
1!
1%
1-
12
#711860000000
0!
0%
b1 *
0-
02
b1 6
#711870000000
1!
1%
1-
12
#711880000000
0!
0%
b10 *
0-
02
b10 6
#711890000000
1!
1%
1-
12
#711900000000
0!
0%
b11 *
0-
02
b11 6
#711910000000
1!
1%
1-
12
15
#711920000000
0!
0%
b100 *
0-
02
b100 6
#711930000000
1!
1%
1-
12
#711940000000
0!
0%
b101 *
0-
02
b101 6
#711950000000
1!
1%
1-
12
#711960000000
0!
0%
b110 *
0-
02
b110 6
#711970000000
1!
1%
1-
12
#711980000000
0!
0%
b111 *
0-
02
b111 6
#711990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#712000000000
0!
0%
b0 *
0-
02
b0 6
#712010000000
1!
1%
1-
12
#712020000000
0!
0%
b1 *
0-
02
b1 6
#712030000000
1!
1%
1-
12
#712040000000
0!
0%
b10 *
0-
02
b10 6
#712050000000
1!
1%
1-
12
#712060000000
0!
0%
b11 *
0-
02
b11 6
#712070000000
1!
1%
1-
12
15
#712080000000
0!
0%
b100 *
0-
02
b100 6
#712090000000
1!
1%
1-
12
#712100000000
0!
0%
b101 *
0-
02
b101 6
#712110000000
1!
1%
1-
12
#712120000000
0!
0%
b110 *
0-
02
b110 6
#712130000000
1!
1%
1-
12
#712140000000
0!
0%
b111 *
0-
02
b111 6
#712150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#712160000000
0!
0%
b0 *
0-
02
b0 6
#712170000000
1!
1%
1-
12
#712180000000
0!
0%
b1 *
0-
02
b1 6
#712190000000
1!
1%
1-
12
#712200000000
0!
0%
b10 *
0-
02
b10 6
#712210000000
1!
1%
1-
12
#712220000000
0!
0%
b11 *
0-
02
b11 6
#712230000000
1!
1%
1-
12
15
#712240000000
0!
0%
b100 *
0-
02
b100 6
#712250000000
1!
1%
1-
12
#712260000000
0!
0%
b101 *
0-
02
b101 6
#712270000000
1!
1%
1-
12
#712280000000
0!
0%
b110 *
0-
02
b110 6
#712290000000
1!
1%
1-
12
#712300000000
0!
0%
b111 *
0-
02
b111 6
#712310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#712320000000
0!
0%
b0 *
0-
02
b0 6
#712330000000
1!
1%
1-
12
#712340000000
0!
0%
b1 *
0-
02
b1 6
#712350000000
1!
1%
1-
12
#712360000000
0!
0%
b10 *
0-
02
b10 6
#712370000000
1!
1%
1-
12
#712380000000
0!
0%
b11 *
0-
02
b11 6
#712390000000
1!
1%
1-
12
15
#712400000000
0!
0%
b100 *
0-
02
b100 6
#712410000000
1!
1%
1-
12
#712420000000
0!
0%
b101 *
0-
02
b101 6
#712430000000
1!
1%
1-
12
#712440000000
0!
0%
b110 *
0-
02
b110 6
#712450000000
1!
1%
1-
12
#712460000000
0!
0%
b111 *
0-
02
b111 6
#712470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#712480000000
0!
0%
b0 *
0-
02
b0 6
#712490000000
1!
1%
1-
12
#712500000000
0!
0%
b1 *
0-
02
b1 6
#712510000000
1!
1%
1-
12
#712520000000
0!
0%
b10 *
0-
02
b10 6
#712530000000
1!
1%
1-
12
#712540000000
0!
0%
b11 *
0-
02
b11 6
#712550000000
1!
1%
1-
12
15
#712560000000
0!
0%
b100 *
0-
02
b100 6
#712570000000
1!
1%
1-
12
#712580000000
0!
0%
b101 *
0-
02
b101 6
#712590000000
1!
1%
1-
12
#712600000000
0!
0%
b110 *
0-
02
b110 6
#712610000000
1!
1%
1-
12
#712620000000
0!
0%
b111 *
0-
02
b111 6
#712630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#712640000000
0!
0%
b0 *
0-
02
b0 6
#712650000000
1!
1%
1-
12
#712660000000
0!
0%
b1 *
0-
02
b1 6
#712670000000
1!
1%
1-
12
#712680000000
0!
0%
b10 *
0-
02
b10 6
#712690000000
1!
1%
1-
12
#712700000000
0!
0%
b11 *
0-
02
b11 6
#712710000000
1!
1%
1-
12
15
#712720000000
0!
0%
b100 *
0-
02
b100 6
#712730000000
1!
1%
1-
12
#712740000000
0!
0%
b101 *
0-
02
b101 6
#712750000000
1!
1%
1-
12
#712760000000
0!
0%
b110 *
0-
02
b110 6
#712770000000
1!
1%
1-
12
#712780000000
0!
0%
b111 *
0-
02
b111 6
#712790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#712800000000
0!
0%
b0 *
0-
02
b0 6
#712810000000
1!
1%
1-
12
#712820000000
0!
0%
b1 *
0-
02
b1 6
#712830000000
1!
1%
1-
12
#712840000000
0!
0%
b10 *
0-
02
b10 6
#712850000000
1!
1%
1-
12
#712860000000
0!
0%
b11 *
0-
02
b11 6
#712870000000
1!
1%
1-
12
15
#712880000000
0!
0%
b100 *
0-
02
b100 6
#712890000000
1!
1%
1-
12
#712900000000
0!
0%
b101 *
0-
02
b101 6
#712910000000
1!
1%
1-
12
#712920000000
0!
0%
b110 *
0-
02
b110 6
#712930000000
1!
1%
1-
12
#712940000000
0!
0%
b111 *
0-
02
b111 6
#712950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#712960000000
0!
0%
b0 *
0-
02
b0 6
#712970000000
1!
1%
1-
12
#712980000000
0!
0%
b1 *
0-
02
b1 6
#712990000000
1!
1%
1-
12
#713000000000
0!
0%
b10 *
0-
02
b10 6
#713010000000
1!
1%
1-
12
#713020000000
0!
0%
b11 *
0-
02
b11 6
#713030000000
1!
1%
1-
12
15
#713040000000
0!
0%
b100 *
0-
02
b100 6
#713050000000
1!
1%
1-
12
#713060000000
0!
0%
b101 *
0-
02
b101 6
#713070000000
1!
1%
1-
12
#713080000000
0!
0%
b110 *
0-
02
b110 6
#713090000000
1!
1%
1-
12
#713100000000
0!
0%
b111 *
0-
02
b111 6
#713110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#713120000000
0!
0%
b0 *
0-
02
b0 6
#713130000000
1!
1%
1-
12
#713140000000
0!
0%
b1 *
0-
02
b1 6
#713150000000
1!
1%
1-
12
#713160000000
0!
0%
b10 *
0-
02
b10 6
#713170000000
1!
1%
1-
12
#713180000000
0!
0%
b11 *
0-
02
b11 6
#713190000000
1!
1%
1-
12
15
#713200000000
0!
0%
b100 *
0-
02
b100 6
#713210000000
1!
1%
1-
12
#713220000000
0!
0%
b101 *
0-
02
b101 6
#713230000000
1!
1%
1-
12
#713240000000
0!
0%
b110 *
0-
02
b110 6
#713250000000
1!
1%
1-
12
#713260000000
0!
0%
b111 *
0-
02
b111 6
#713270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#713280000000
0!
0%
b0 *
0-
02
b0 6
#713290000000
1!
1%
1-
12
#713300000000
0!
0%
b1 *
0-
02
b1 6
#713310000000
1!
1%
1-
12
#713320000000
0!
0%
b10 *
0-
02
b10 6
#713330000000
1!
1%
1-
12
#713340000000
0!
0%
b11 *
0-
02
b11 6
#713350000000
1!
1%
1-
12
15
#713360000000
0!
0%
b100 *
0-
02
b100 6
#713370000000
1!
1%
1-
12
#713380000000
0!
0%
b101 *
0-
02
b101 6
#713390000000
1!
1%
1-
12
#713400000000
0!
0%
b110 *
0-
02
b110 6
#713410000000
1!
1%
1-
12
#713420000000
0!
0%
b111 *
0-
02
b111 6
#713430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#713440000000
0!
0%
b0 *
0-
02
b0 6
#713450000000
1!
1%
1-
12
#713460000000
0!
0%
b1 *
0-
02
b1 6
#713470000000
1!
1%
1-
12
#713480000000
0!
0%
b10 *
0-
02
b10 6
#713490000000
1!
1%
1-
12
#713500000000
0!
0%
b11 *
0-
02
b11 6
#713510000000
1!
1%
1-
12
15
#713520000000
0!
0%
b100 *
0-
02
b100 6
#713530000000
1!
1%
1-
12
#713540000000
0!
0%
b101 *
0-
02
b101 6
#713550000000
1!
1%
1-
12
#713560000000
0!
0%
b110 *
0-
02
b110 6
#713570000000
1!
1%
1-
12
#713580000000
0!
0%
b111 *
0-
02
b111 6
#713590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#713600000000
0!
0%
b0 *
0-
02
b0 6
#713610000000
1!
1%
1-
12
#713620000000
0!
0%
b1 *
0-
02
b1 6
#713630000000
1!
1%
1-
12
#713640000000
0!
0%
b10 *
0-
02
b10 6
#713650000000
1!
1%
1-
12
#713660000000
0!
0%
b11 *
0-
02
b11 6
#713670000000
1!
1%
1-
12
15
#713680000000
0!
0%
b100 *
0-
02
b100 6
#713690000000
1!
1%
1-
12
#713700000000
0!
0%
b101 *
0-
02
b101 6
#713710000000
1!
1%
1-
12
#713720000000
0!
0%
b110 *
0-
02
b110 6
#713730000000
1!
1%
1-
12
#713740000000
0!
0%
b111 *
0-
02
b111 6
#713750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#713760000000
0!
0%
b0 *
0-
02
b0 6
#713770000000
1!
1%
1-
12
#713780000000
0!
0%
b1 *
0-
02
b1 6
#713790000000
1!
1%
1-
12
#713800000000
0!
0%
b10 *
0-
02
b10 6
#713810000000
1!
1%
1-
12
#713820000000
0!
0%
b11 *
0-
02
b11 6
#713830000000
1!
1%
1-
12
15
#713840000000
0!
0%
b100 *
0-
02
b100 6
#713850000000
1!
1%
1-
12
#713860000000
0!
0%
b101 *
0-
02
b101 6
#713870000000
1!
1%
1-
12
#713880000000
0!
0%
b110 *
0-
02
b110 6
#713890000000
1!
1%
1-
12
#713900000000
0!
0%
b111 *
0-
02
b111 6
#713910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#713920000000
0!
0%
b0 *
0-
02
b0 6
#713930000000
1!
1%
1-
12
#713940000000
0!
0%
b1 *
0-
02
b1 6
#713950000000
1!
1%
1-
12
#713960000000
0!
0%
b10 *
0-
02
b10 6
#713970000000
1!
1%
1-
12
#713980000000
0!
0%
b11 *
0-
02
b11 6
#713990000000
1!
1%
1-
12
15
#714000000000
0!
0%
b100 *
0-
02
b100 6
#714010000000
1!
1%
1-
12
#714020000000
0!
0%
b101 *
0-
02
b101 6
#714030000000
1!
1%
1-
12
#714040000000
0!
0%
b110 *
0-
02
b110 6
#714050000000
1!
1%
1-
12
#714060000000
0!
0%
b111 *
0-
02
b111 6
#714070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#714080000000
0!
0%
b0 *
0-
02
b0 6
#714090000000
1!
1%
1-
12
#714100000000
0!
0%
b1 *
0-
02
b1 6
#714110000000
1!
1%
1-
12
#714120000000
0!
0%
b10 *
0-
02
b10 6
#714130000000
1!
1%
1-
12
#714140000000
0!
0%
b11 *
0-
02
b11 6
#714150000000
1!
1%
1-
12
15
#714160000000
0!
0%
b100 *
0-
02
b100 6
#714170000000
1!
1%
1-
12
#714180000000
0!
0%
b101 *
0-
02
b101 6
#714190000000
1!
1%
1-
12
#714200000000
0!
0%
b110 *
0-
02
b110 6
#714210000000
1!
1%
1-
12
#714220000000
0!
0%
b111 *
0-
02
b111 6
#714230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#714240000000
0!
0%
b0 *
0-
02
b0 6
#714250000000
1!
1%
1-
12
#714260000000
0!
0%
b1 *
0-
02
b1 6
#714270000000
1!
1%
1-
12
#714280000000
0!
0%
b10 *
0-
02
b10 6
#714290000000
1!
1%
1-
12
#714300000000
0!
0%
b11 *
0-
02
b11 6
#714310000000
1!
1%
1-
12
15
#714320000000
0!
0%
b100 *
0-
02
b100 6
#714330000000
1!
1%
1-
12
#714340000000
0!
0%
b101 *
0-
02
b101 6
#714350000000
1!
1%
1-
12
#714360000000
0!
0%
b110 *
0-
02
b110 6
#714370000000
1!
1%
1-
12
#714380000000
0!
0%
b111 *
0-
02
b111 6
#714390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#714400000000
0!
0%
b0 *
0-
02
b0 6
#714410000000
1!
1%
1-
12
#714420000000
0!
0%
b1 *
0-
02
b1 6
#714430000000
1!
1%
1-
12
#714440000000
0!
0%
b10 *
0-
02
b10 6
#714450000000
1!
1%
1-
12
#714460000000
0!
0%
b11 *
0-
02
b11 6
#714470000000
1!
1%
1-
12
15
#714480000000
0!
0%
b100 *
0-
02
b100 6
#714490000000
1!
1%
1-
12
#714500000000
0!
0%
b101 *
0-
02
b101 6
#714510000000
1!
1%
1-
12
#714520000000
0!
0%
b110 *
0-
02
b110 6
#714530000000
1!
1%
1-
12
#714540000000
0!
0%
b111 *
0-
02
b111 6
#714550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#714560000000
0!
0%
b0 *
0-
02
b0 6
#714570000000
1!
1%
1-
12
#714580000000
0!
0%
b1 *
0-
02
b1 6
#714590000000
1!
1%
1-
12
#714600000000
0!
0%
b10 *
0-
02
b10 6
#714610000000
1!
1%
1-
12
#714620000000
0!
0%
b11 *
0-
02
b11 6
#714630000000
1!
1%
1-
12
15
#714640000000
0!
0%
b100 *
0-
02
b100 6
#714650000000
1!
1%
1-
12
#714660000000
0!
0%
b101 *
0-
02
b101 6
#714670000000
1!
1%
1-
12
#714680000000
0!
0%
b110 *
0-
02
b110 6
#714690000000
1!
1%
1-
12
#714700000000
0!
0%
b111 *
0-
02
b111 6
#714710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#714720000000
0!
0%
b0 *
0-
02
b0 6
#714730000000
1!
1%
1-
12
#714740000000
0!
0%
b1 *
0-
02
b1 6
#714750000000
1!
1%
1-
12
#714760000000
0!
0%
b10 *
0-
02
b10 6
#714770000000
1!
1%
1-
12
#714780000000
0!
0%
b11 *
0-
02
b11 6
#714790000000
1!
1%
1-
12
15
#714800000000
0!
0%
b100 *
0-
02
b100 6
#714810000000
1!
1%
1-
12
#714820000000
0!
0%
b101 *
0-
02
b101 6
#714830000000
1!
1%
1-
12
#714840000000
0!
0%
b110 *
0-
02
b110 6
#714850000000
1!
1%
1-
12
#714860000000
0!
0%
b111 *
0-
02
b111 6
#714870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#714880000000
0!
0%
b0 *
0-
02
b0 6
#714890000000
1!
1%
1-
12
#714900000000
0!
0%
b1 *
0-
02
b1 6
#714910000000
1!
1%
1-
12
#714920000000
0!
0%
b10 *
0-
02
b10 6
#714930000000
1!
1%
1-
12
#714940000000
0!
0%
b11 *
0-
02
b11 6
#714950000000
1!
1%
1-
12
15
#714960000000
0!
0%
b100 *
0-
02
b100 6
#714970000000
1!
1%
1-
12
#714980000000
0!
0%
b101 *
0-
02
b101 6
#714990000000
1!
1%
1-
12
#715000000000
0!
0%
b110 *
0-
02
b110 6
#715010000000
1!
1%
1-
12
#715020000000
0!
0%
b111 *
0-
02
b111 6
#715030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#715040000000
0!
0%
b0 *
0-
02
b0 6
#715050000000
1!
1%
1-
12
#715060000000
0!
0%
b1 *
0-
02
b1 6
#715070000000
1!
1%
1-
12
#715080000000
0!
0%
b10 *
0-
02
b10 6
#715090000000
1!
1%
1-
12
#715100000000
0!
0%
b11 *
0-
02
b11 6
#715110000000
1!
1%
1-
12
15
#715120000000
0!
0%
b100 *
0-
02
b100 6
#715130000000
1!
1%
1-
12
#715140000000
0!
0%
b101 *
0-
02
b101 6
#715150000000
1!
1%
1-
12
#715160000000
0!
0%
b110 *
0-
02
b110 6
#715170000000
1!
1%
1-
12
#715180000000
0!
0%
b111 *
0-
02
b111 6
#715190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#715200000000
0!
0%
b0 *
0-
02
b0 6
#715210000000
1!
1%
1-
12
#715220000000
0!
0%
b1 *
0-
02
b1 6
#715230000000
1!
1%
1-
12
#715240000000
0!
0%
b10 *
0-
02
b10 6
#715250000000
1!
1%
1-
12
#715260000000
0!
0%
b11 *
0-
02
b11 6
#715270000000
1!
1%
1-
12
15
#715280000000
0!
0%
b100 *
0-
02
b100 6
#715290000000
1!
1%
1-
12
#715300000000
0!
0%
b101 *
0-
02
b101 6
#715310000000
1!
1%
1-
12
#715320000000
0!
0%
b110 *
0-
02
b110 6
#715330000000
1!
1%
1-
12
#715340000000
0!
0%
b111 *
0-
02
b111 6
#715350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#715360000000
0!
0%
b0 *
0-
02
b0 6
#715370000000
1!
1%
1-
12
#715380000000
0!
0%
b1 *
0-
02
b1 6
#715390000000
1!
1%
1-
12
#715400000000
0!
0%
b10 *
0-
02
b10 6
#715410000000
1!
1%
1-
12
#715420000000
0!
0%
b11 *
0-
02
b11 6
#715430000000
1!
1%
1-
12
15
#715440000000
0!
0%
b100 *
0-
02
b100 6
#715450000000
1!
1%
1-
12
#715460000000
0!
0%
b101 *
0-
02
b101 6
#715470000000
1!
1%
1-
12
#715480000000
0!
0%
b110 *
0-
02
b110 6
#715490000000
1!
1%
1-
12
#715500000000
0!
0%
b111 *
0-
02
b111 6
#715510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#715520000000
0!
0%
b0 *
0-
02
b0 6
#715530000000
1!
1%
1-
12
#715540000000
0!
0%
b1 *
0-
02
b1 6
#715550000000
1!
1%
1-
12
#715560000000
0!
0%
b10 *
0-
02
b10 6
#715570000000
1!
1%
1-
12
#715580000000
0!
0%
b11 *
0-
02
b11 6
#715590000000
1!
1%
1-
12
15
#715600000000
0!
0%
b100 *
0-
02
b100 6
#715610000000
1!
1%
1-
12
#715620000000
0!
0%
b101 *
0-
02
b101 6
#715630000000
1!
1%
1-
12
#715640000000
0!
0%
b110 *
0-
02
b110 6
#715650000000
1!
1%
1-
12
#715660000000
0!
0%
b111 *
0-
02
b111 6
#715670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#715680000000
0!
0%
b0 *
0-
02
b0 6
#715690000000
1!
1%
1-
12
#715700000000
0!
0%
b1 *
0-
02
b1 6
#715710000000
1!
1%
1-
12
#715720000000
0!
0%
b10 *
0-
02
b10 6
#715730000000
1!
1%
1-
12
#715740000000
0!
0%
b11 *
0-
02
b11 6
#715750000000
1!
1%
1-
12
15
#715760000000
0!
0%
b100 *
0-
02
b100 6
#715770000000
1!
1%
1-
12
#715780000000
0!
0%
b101 *
0-
02
b101 6
#715790000000
1!
1%
1-
12
#715800000000
0!
0%
b110 *
0-
02
b110 6
#715810000000
1!
1%
1-
12
#715820000000
0!
0%
b111 *
0-
02
b111 6
#715830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#715840000000
0!
0%
b0 *
0-
02
b0 6
#715850000000
1!
1%
1-
12
#715860000000
0!
0%
b1 *
0-
02
b1 6
#715870000000
1!
1%
1-
12
#715880000000
0!
0%
b10 *
0-
02
b10 6
#715890000000
1!
1%
1-
12
#715900000000
0!
0%
b11 *
0-
02
b11 6
#715910000000
1!
1%
1-
12
15
#715920000000
0!
0%
b100 *
0-
02
b100 6
#715930000000
1!
1%
1-
12
#715940000000
0!
0%
b101 *
0-
02
b101 6
#715950000000
1!
1%
1-
12
#715960000000
0!
0%
b110 *
0-
02
b110 6
#715970000000
1!
1%
1-
12
#715980000000
0!
0%
b111 *
0-
02
b111 6
#715990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#716000000000
0!
0%
b0 *
0-
02
b0 6
#716010000000
1!
1%
1-
12
#716020000000
0!
0%
b1 *
0-
02
b1 6
#716030000000
1!
1%
1-
12
#716040000000
0!
0%
b10 *
0-
02
b10 6
#716050000000
1!
1%
1-
12
#716060000000
0!
0%
b11 *
0-
02
b11 6
#716070000000
1!
1%
1-
12
15
#716080000000
0!
0%
b100 *
0-
02
b100 6
#716090000000
1!
1%
1-
12
#716100000000
0!
0%
b101 *
0-
02
b101 6
#716110000000
1!
1%
1-
12
#716120000000
0!
0%
b110 *
0-
02
b110 6
#716130000000
1!
1%
1-
12
#716140000000
0!
0%
b111 *
0-
02
b111 6
#716150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#716160000000
0!
0%
b0 *
0-
02
b0 6
#716170000000
1!
1%
1-
12
#716180000000
0!
0%
b1 *
0-
02
b1 6
#716190000000
1!
1%
1-
12
#716200000000
0!
0%
b10 *
0-
02
b10 6
#716210000000
1!
1%
1-
12
#716220000000
0!
0%
b11 *
0-
02
b11 6
#716230000000
1!
1%
1-
12
15
#716240000000
0!
0%
b100 *
0-
02
b100 6
#716250000000
1!
1%
1-
12
#716260000000
0!
0%
b101 *
0-
02
b101 6
#716270000000
1!
1%
1-
12
#716280000000
0!
0%
b110 *
0-
02
b110 6
#716290000000
1!
1%
1-
12
#716300000000
0!
0%
b111 *
0-
02
b111 6
#716310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#716320000000
0!
0%
b0 *
0-
02
b0 6
#716330000000
1!
1%
1-
12
#716340000000
0!
0%
b1 *
0-
02
b1 6
#716350000000
1!
1%
1-
12
#716360000000
0!
0%
b10 *
0-
02
b10 6
#716370000000
1!
1%
1-
12
#716380000000
0!
0%
b11 *
0-
02
b11 6
#716390000000
1!
1%
1-
12
15
#716400000000
0!
0%
b100 *
0-
02
b100 6
#716410000000
1!
1%
1-
12
#716420000000
0!
0%
b101 *
0-
02
b101 6
#716430000000
1!
1%
1-
12
#716440000000
0!
0%
b110 *
0-
02
b110 6
#716450000000
1!
1%
1-
12
#716460000000
0!
0%
b111 *
0-
02
b111 6
#716470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#716480000000
0!
0%
b0 *
0-
02
b0 6
#716490000000
1!
1%
1-
12
#716500000000
0!
0%
b1 *
0-
02
b1 6
#716510000000
1!
1%
1-
12
#716520000000
0!
0%
b10 *
0-
02
b10 6
#716530000000
1!
1%
1-
12
#716540000000
0!
0%
b11 *
0-
02
b11 6
#716550000000
1!
1%
1-
12
15
#716560000000
0!
0%
b100 *
0-
02
b100 6
#716570000000
1!
1%
1-
12
#716580000000
0!
0%
b101 *
0-
02
b101 6
#716590000000
1!
1%
1-
12
#716600000000
0!
0%
b110 *
0-
02
b110 6
#716610000000
1!
1%
1-
12
#716620000000
0!
0%
b111 *
0-
02
b111 6
#716630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#716640000000
0!
0%
b0 *
0-
02
b0 6
#716650000000
1!
1%
1-
12
#716660000000
0!
0%
b1 *
0-
02
b1 6
#716670000000
1!
1%
1-
12
#716680000000
0!
0%
b10 *
0-
02
b10 6
#716690000000
1!
1%
1-
12
#716700000000
0!
0%
b11 *
0-
02
b11 6
#716710000000
1!
1%
1-
12
15
#716720000000
0!
0%
b100 *
0-
02
b100 6
#716730000000
1!
1%
1-
12
#716740000000
0!
0%
b101 *
0-
02
b101 6
#716750000000
1!
1%
1-
12
#716760000000
0!
0%
b110 *
0-
02
b110 6
#716770000000
1!
1%
1-
12
#716780000000
0!
0%
b111 *
0-
02
b111 6
#716790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#716800000000
0!
0%
b0 *
0-
02
b0 6
#716810000000
1!
1%
1-
12
#716820000000
0!
0%
b1 *
0-
02
b1 6
#716830000000
1!
1%
1-
12
#716840000000
0!
0%
b10 *
0-
02
b10 6
#716850000000
1!
1%
1-
12
#716860000000
0!
0%
b11 *
0-
02
b11 6
#716870000000
1!
1%
1-
12
15
#716880000000
0!
0%
b100 *
0-
02
b100 6
#716890000000
1!
1%
1-
12
#716900000000
0!
0%
b101 *
0-
02
b101 6
#716910000000
1!
1%
1-
12
#716920000000
0!
0%
b110 *
0-
02
b110 6
#716930000000
1!
1%
1-
12
#716940000000
0!
0%
b111 *
0-
02
b111 6
#716950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#716960000000
0!
0%
b0 *
0-
02
b0 6
#716970000000
1!
1%
1-
12
#716980000000
0!
0%
b1 *
0-
02
b1 6
#716990000000
1!
1%
1-
12
#717000000000
0!
0%
b10 *
0-
02
b10 6
#717010000000
1!
1%
1-
12
#717020000000
0!
0%
b11 *
0-
02
b11 6
#717030000000
1!
1%
1-
12
15
#717040000000
0!
0%
b100 *
0-
02
b100 6
#717050000000
1!
1%
1-
12
#717060000000
0!
0%
b101 *
0-
02
b101 6
#717070000000
1!
1%
1-
12
#717080000000
0!
0%
b110 *
0-
02
b110 6
#717090000000
1!
1%
1-
12
#717100000000
0!
0%
b111 *
0-
02
b111 6
#717110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#717120000000
0!
0%
b0 *
0-
02
b0 6
#717130000000
1!
1%
1-
12
#717140000000
0!
0%
b1 *
0-
02
b1 6
#717150000000
1!
1%
1-
12
#717160000000
0!
0%
b10 *
0-
02
b10 6
#717170000000
1!
1%
1-
12
#717180000000
0!
0%
b11 *
0-
02
b11 6
#717190000000
1!
1%
1-
12
15
#717200000000
0!
0%
b100 *
0-
02
b100 6
#717210000000
1!
1%
1-
12
#717220000000
0!
0%
b101 *
0-
02
b101 6
#717230000000
1!
1%
1-
12
#717240000000
0!
0%
b110 *
0-
02
b110 6
#717250000000
1!
1%
1-
12
#717260000000
0!
0%
b111 *
0-
02
b111 6
#717270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#717280000000
0!
0%
b0 *
0-
02
b0 6
#717290000000
1!
1%
1-
12
#717300000000
0!
0%
b1 *
0-
02
b1 6
#717310000000
1!
1%
1-
12
#717320000000
0!
0%
b10 *
0-
02
b10 6
#717330000000
1!
1%
1-
12
#717340000000
0!
0%
b11 *
0-
02
b11 6
#717350000000
1!
1%
1-
12
15
#717360000000
0!
0%
b100 *
0-
02
b100 6
#717370000000
1!
1%
1-
12
#717380000000
0!
0%
b101 *
0-
02
b101 6
#717390000000
1!
1%
1-
12
#717400000000
0!
0%
b110 *
0-
02
b110 6
#717410000000
1!
1%
1-
12
#717420000000
0!
0%
b111 *
0-
02
b111 6
#717430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#717440000000
0!
0%
b0 *
0-
02
b0 6
#717450000000
1!
1%
1-
12
#717460000000
0!
0%
b1 *
0-
02
b1 6
#717470000000
1!
1%
1-
12
#717480000000
0!
0%
b10 *
0-
02
b10 6
#717490000000
1!
1%
1-
12
#717500000000
0!
0%
b11 *
0-
02
b11 6
#717510000000
1!
1%
1-
12
15
#717520000000
0!
0%
b100 *
0-
02
b100 6
#717530000000
1!
1%
1-
12
#717540000000
0!
0%
b101 *
0-
02
b101 6
#717550000000
1!
1%
1-
12
#717560000000
0!
0%
b110 *
0-
02
b110 6
#717570000000
1!
1%
1-
12
#717580000000
0!
0%
b111 *
0-
02
b111 6
#717590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#717600000000
0!
0%
b0 *
0-
02
b0 6
#717610000000
1!
1%
1-
12
#717620000000
0!
0%
b1 *
0-
02
b1 6
#717630000000
1!
1%
1-
12
#717640000000
0!
0%
b10 *
0-
02
b10 6
#717650000000
1!
1%
1-
12
#717660000000
0!
0%
b11 *
0-
02
b11 6
#717670000000
1!
1%
1-
12
15
#717680000000
0!
0%
b100 *
0-
02
b100 6
#717690000000
1!
1%
1-
12
#717700000000
0!
0%
b101 *
0-
02
b101 6
#717710000000
1!
1%
1-
12
#717720000000
0!
0%
b110 *
0-
02
b110 6
#717730000000
1!
1%
1-
12
#717740000000
0!
0%
b111 *
0-
02
b111 6
#717750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#717760000000
0!
0%
b0 *
0-
02
b0 6
#717770000000
1!
1%
1-
12
#717780000000
0!
0%
b1 *
0-
02
b1 6
#717790000000
1!
1%
1-
12
#717800000000
0!
0%
b10 *
0-
02
b10 6
#717810000000
1!
1%
1-
12
#717820000000
0!
0%
b11 *
0-
02
b11 6
#717830000000
1!
1%
1-
12
15
#717840000000
0!
0%
b100 *
0-
02
b100 6
#717850000000
1!
1%
1-
12
#717860000000
0!
0%
b101 *
0-
02
b101 6
#717870000000
1!
1%
1-
12
#717880000000
0!
0%
b110 *
0-
02
b110 6
#717890000000
1!
1%
1-
12
#717900000000
0!
0%
b111 *
0-
02
b111 6
#717910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#717920000000
0!
0%
b0 *
0-
02
b0 6
#717930000000
1!
1%
1-
12
#717940000000
0!
0%
b1 *
0-
02
b1 6
#717950000000
1!
1%
1-
12
#717960000000
0!
0%
b10 *
0-
02
b10 6
#717970000000
1!
1%
1-
12
#717980000000
0!
0%
b11 *
0-
02
b11 6
#717990000000
1!
1%
1-
12
15
#718000000000
0!
0%
b100 *
0-
02
b100 6
#718010000000
1!
1%
1-
12
#718020000000
0!
0%
b101 *
0-
02
b101 6
#718030000000
1!
1%
1-
12
#718040000000
0!
0%
b110 *
0-
02
b110 6
#718050000000
1!
1%
1-
12
#718060000000
0!
0%
b111 *
0-
02
b111 6
#718070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#718080000000
0!
0%
b0 *
0-
02
b0 6
#718090000000
1!
1%
1-
12
#718100000000
0!
0%
b1 *
0-
02
b1 6
#718110000000
1!
1%
1-
12
#718120000000
0!
0%
b10 *
0-
02
b10 6
#718130000000
1!
1%
1-
12
#718140000000
0!
0%
b11 *
0-
02
b11 6
#718150000000
1!
1%
1-
12
15
#718160000000
0!
0%
b100 *
0-
02
b100 6
#718170000000
1!
1%
1-
12
#718180000000
0!
0%
b101 *
0-
02
b101 6
#718190000000
1!
1%
1-
12
#718200000000
0!
0%
b110 *
0-
02
b110 6
#718210000000
1!
1%
1-
12
#718220000000
0!
0%
b111 *
0-
02
b111 6
#718230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#718240000000
0!
0%
b0 *
0-
02
b0 6
#718250000000
1!
1%
1-
12
#718260000000
0!
0%
b1 *
0-
02
b1 6
#718270000000
1!
1%
1-
12
#718280000000
0!
0%
b10 *
0-
02
b10 6
#718290000000
1!
1%
1-
12
#718300000000
0!
0%
b11 *
0-
02
b11 6
#718310000000
1!
1%
1-
12
15
#718320000000
0!
0%
b100 *
0-
02
b100 6
#718330000000
1!
1%
1-
12
#718340000000
0!
0%
b101 *
0-
02
b101 6
#718350000000
1!
1%
1-
12
#718360000000
0!
0%
b110 *
0-
02
b110 6
#718370000000
1!
1%
1-
12
#718380000000
0!
0%
b111 *
0-
02
b111 6
#718390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#718400000000
0!
0%
b0 *
0-
02
b0 6
#718410000000
1!
1%
1-
12
#718420000000
0!
0%
b1 *
0-
02
b1 6
#718430000000
1!
1%
1-
12
#718440000000
0!
0%
b10 *
0-
02
b10 6
#718450000000
1!
1%
1-
12
#718460000000
0!
0%
b11 *
0-
02
b11 6
#718470000000
1!
1%
1-
12
15
#718480000000
0!
0%
b100 *
0-
02
b100 6
#718490000000
1!
1%
1-
12
#718500000000
0!
0%
b101 *
0-
02
b101 6
#718510000000
1!
1%
1-
12
#718520000000
0!
0%
b110 *
0-
02
b110 6
#718530000000
1!
1%
1-
12
#718540000000
0!
0%
b111 *
0-
02
b111 6
#718550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#718560000000
0!
0%
b0 *
0-
02
b0 6
#718570000000
1!
1%
1-
12
#718580000000
0!
0%
b1 *
0-
02
b1 6
#718590000000
1!
1%
1-
12
#718600000000
0!
0%
b10 *
0-
02
b10 6
#718610000000
1!
1%
1-
12
#718620000000
0!
0%
b11 *
0-
02
b11 6
#718630000000
1!
1%
1-
12
15
#718640000000
0!
0%
b100 *
0-
02
b100 6
#718650000000
1!
1%
1-
12
#718660000000
0!
0%
b101 *
0-
02
b101 6
#718670000000
1!
1%
1-
12
#718680000000
0!
0%
b110 *
0-
02
b110 6
#718690000000
1!
1%
1-
12
#718700000000
0!
0%
b111 *
0-
02
b111 6
#718710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#718720000000
0!
0%
b0 *
0-
02
b0 6
#718730000000
1!
1%
1-
12
#718740000000
0!
0%
b1 *
0-
02
b1 6
#718750000000
1!
1%
1-
12
#718760000000
0!
0%
b10 *
0-
02
b10 6
#718770000000
1!
1%
1-
12
#718780000000
0!
0%
b11 *
0-
02
b11 6
#718790000000
1!
1%
1-
12
15
#718800000000
0!
0%
b100 *
0-
02
b100 6
#718810000000
1!
1%
1-
12
#718820000000
0!
0%
b101 *
0-
02
b101 6
#718830000000
1!
1%
1-
12
#718840000000
0!
0%
b110 *
0-
02
b110 6
#718850000000
1!
1%
1-
12
#718860000000
0!
0%
b111 *
0-
02
b111 6
#718870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#718880000000
0!
0%
b0 *
0-
02
b0 6
#718890000000
1!
1%
1-
12
#718900000000
0!
0%
b1 *
0-
02
b1 6
#718910000000
1!
1%
1-
12
#718920000000
0!
0%
b10 *
0-
02
b10 6
#718930000000
1!
1%
1-
12
#718940000000
0!
0%
b11 *
0-
02
b11 6
#718950000000
1!
1%
1-
12
15
#718960000000
0!
0%
b100 *
0-
02
b100 6
#718970000000
1!
1%
1-
12
#718980000000
0!
0%
b101 *
0-
02
b101 6
#718990000000
1!
1%
1-
12
#719000000000
0!
0%
b110 *
0-
02
b110 6
#719010000000
1!
1%
1-
12
#719020000000
0!
0%
b111 *
0-
02
b111 6
#719030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#719040000000
0!
0%
b0 *
0-
02
b0 6
#719050000000
1!
1%
1-
12
#719060000000
0!
0%
b1 *
0-
02
b1 6
#719070000000
1!
1%
1-
12
#719080000000
0!
0%
b10 *
0-
02
b10 6
#719090000000
1!
1%
1-
12
#719100000000
0!
0%
b11 *
0-
02
b11 6
#719110000000
1!
1%
1-
12
15
#719120000000
0!
0%
b100 *
0-
02
b100 6
#719130000000
1!
1%
1-
12
#719140000000
0!
0%
b101 *
0-
02
b101 6
#719150000000
1!
1%
1-
12
#719160000000
0!
0%
b110 *
0-
02
b110 6
#719170000000
1!
1%
1-
12
#719180000000
0!
0%
b111 *
0-
02
b111 6
#719190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#719200000000
0!
0%
b0 *
0-
02
b0 6
#719210000000
1!
1%
1-
12
#719220000000
0!
0%
b1 *
0-
02
b1 6
#719230000000
1!
1%
1-
12
#719240000000
0!
0%
b10 *
0-
02
b10 6
#719250000000
1!
1%
1-
12
#719260000000
0!
0%
b11 *
0-
02
b11 6
#719270000000
1!
1%
1-
12
15
#719280000000
0!
0%
b100 *
0-
02
b100 6
#719290000000
1!
1%
1-
12
#719300000000
0!
0%
b101 *
0-
02
b101 6
#719310000000
1!
1%
1-
12
#719320000000
0!
0%
b110 *
0-
02
b110 6
#719330000000
1!
1%
1-
12
#719340000000
0!
0%
b111 *
0-
02
b111 6
#719350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#719360000000
0!
0%
b0 *
0-
02
b0 6
#719370000000
1!
1%
1-
12
#719380000000
0!
0%
b1 *
0-
02
b1 6
#719390000000
1!
1%
1-
12
#719400000000
0!
0%
b10 *
0-
02
b10 6
#719410000000
1!
1%
1-
12
#719420000000
0!
0%
b11 *
0-
02
b11 6
#719430000000
1!
1%
1-
12
15
#719440000000
0!
0%
b100 *
0-
02
b100 6
#719450000000
1!
1%
1-
12
#719460000000
0!
0%
b101 *
0-
02
b101 6
#719470000000
1!
1%
1-
12
#719480000000
0!
0%
b110 *
0-
02
b110 6
#719490000000
1!
1%
1-
12
#719500000000
0!
0%
b111 *
0-
02
b111 6
#719510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#719520000000
0!
0%
b0 *
0-
02
b0 6
#719530000000
1!
1%
1-
12
#719540000000
0!
0%
b1 *
0-
02
b1 6
#719550000000
1!
1%
1-
12
#719560000000
0!
0%
b10 *
0-
02
b10 6
#719570000000
1!
1%
1-
12
#719580000000
0!
0%
b11 *
0-
02
b11 6
#719590000000
1!
1%
1-
12
15
#719600000000
0!
0%
b100 *
0-
02
b100 6
#719610000000
1!
1%
1-
12
#719620000000
0!
0%
b101 *
0-
02
b101 6
#719630000000
1!
1%
1-
12
#719640000000
0!
0%
b110 *
0-
02
b110 6
#719650000000
1!
1%
1-
12
#719660000000
0!
0%
b111 *
0-
02
b111 6
#719670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#719680000000
0!
0%
b0 *
0-
02
b0 6
#719690000000
1!
1%
1-
12
#719700000000
0!
0%
b1 *
0-
02
b1 6
#719710000000
1!
1%
1-
12
#719720000000
0!
0%
b10 *
0-
02
b10 6
#719730000000
1!
1%
1-
12
#719740000000
0!
0%
b11 *
0-
02
b11 6
#719750000000
1!
1%
1-
12
15
#719760000000
0!
0%
b100 *
0-
02
b100 6
#719770000000
1!
1%
1-
12
#719780000000
0!
0%
b101 *
0-
02
b101 6
#719790000000
1!
1%
1-
12
#719800000000
0!
0%
b110 *
0-
02
b110 6
#719810000000
1!
1%
1-
12
#719820000000
0!
0%
b111 *
0-
02
b111 6
#719830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#719840000000
0!
0%
b0 *
0-
02
b0 6
#719850000000
1!
1%
1-
12
#719860000000
0!
0%
b1 *
0-
02
b1 6
#719870000000
1!
1%
1-
12
#719880000000
0!
0%
b10 *
0-
02
b10 6
#719890000000
1!
1%
1-
12
#719900000000
0!
0%
b11 *
0-
02
b11 6
#719910000000
1!
1%
1-
12
15
#719920000000
0!
0%
b100 *
0-
02
b100 6
#719930000000
1!
1%
1-
12
#719940000000
0!
0%
b101 *
0-
02
b101 6
#719950000000
1!
1%
1-
12
#719960000000
0!
0%
b110 *
0-
02
b110 6
#719970000000
1!
1%
1-
12
#719980000000
0!
0%
b111 *
0-
02
b111 6
#719990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#720000000000
0!
0%
b0 *
0-
02
b0 6
#720010000000
1!
1%
1-
12
#720020000000
0!
0%
b1 *
0-
02
b1 6
#720030000000
1!
1%
1-
12
#720040000000
0!
0%
b10 *
0-
02
b10 6
#720050000000
1!
1%
1-
12
#720060000000
0!
0%
b11 *
0-
02
b11 6
#720070000000
1!
1%
1-
12
15
#720080000000
0!
0%
b100 *
0-
02
b100 6
#720090000000
1!
1%
1-
12
#720100000000
0!
0%
b101 *
0-
02
b101 6
#720110000000
1!
1%
1-
12
#720120000000
0!
0%
b110 *
0-
02
b110 6
#720130000000
1!
1%
1-
12
#720140000000
0!
0%
b111 *
0-
02
b111 6
#720150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#720160000000
0!
0%
b0 *
0-
02
b0 6
#720170000000
1!
1%
1-
12
#720180000000
0!
0%
b1 *
0-
02
b1 6
#720190000000
1!
1%
1-
12
#720200000000
0!
0%
b10 *
0-
02
b10 6
#720210000000
1!
1%
1-
12
#720220000000
0!
0%
b11 *
0-
02
b11 6
#720230000000
1!
1%
1-
12
15
#720240000000
0!
0%
b100 *
0-
02
b100 6
#720250000000
1!
1%
1-
12
#720260000000
0!
0%
b101 *
0-
02
b101 6
#720270000000
1!
1%
1-
12
#720280000000
0!
0%
b110 *
0-
02
b110 6
#720290000000
1!
1%
1-
12
#720300000000
0!
0%
b111 *
0-
02
b111 6
#720310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#720320000000
0!
0%
b0 *
0-
02
b0 6
#720330000000
1!
1%
1-
12
#720340000000
0!
0%
b1 *
0-
02
b1 6
#720350000000
1!
1%
1-
12
#720360000000
0!
0%
b10 *
0-
02
b10 6
#720370000000
1!
1%
1-
12
#720380000000
0!
0%
b11 *
0-
02
b11 6
#720390000000
1!
1%
1-
12
15
#720400000000
0!
0%
b100 *
0-
02
b100 6
#720410000000
1!
1%
1-
12
#720420000000
0!
0%
b101 *
0-
02
b101 6
#720430000000
1!
1%
1-
12
#720440000000
0!
0%
b110 *
0-
02
b110 6
#720450000000
1!
1%
1-
12
#720460000000
0!
0%
b111 *
0-
02
b111 6
#720470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#720480000000
0!
0%
b0 *
0-
02
b0 6
#720490000000
1!
1%
1-
12
#720500000000
0!
0%
b1 *
0-
02
b1 6
#720510000000
1!
1%
1-
12
#720520000000
0!
0%
b10 *
0-
02
b10 6
#720530000000
1!
1%
1-
12
#720540000000
0!
0%
b11 *
0-
02
b11 6
#720550000000
1!
1%
1-
12
15
#720560000000
0!
0%
b100 *
0-
02
b100 6
#720570000000
1!
1%
1-
12
#720580000000
0!
0%
b101 *
0-
02
b101 6
#720590000000
1!
1%
1-
12
#720600000000
0!
0%
b110 *
0-
02
b110 6
#720610000000
1!
1%
1-
12
#720620000000
0!
0%
b111 *
0-
02
b111 6
#720630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#720640000000
0!
0%
b0 *
0-
02
b0 6
#720650000000
1!
1%
1-
12
#720660000000
0!
0%
b1 *
0-
02
b1 6
#720670000000
1!
1%
1-
12
#720680000000
0!
0%
b10 *
0-
02
b10 6
#720690000000
1!
1%
1-
12
#720700000000
0!
0%
b11 *
0-
02
b11 6
#720710000000
1!
1%
1-
12
15
#720720000000
0!
0%
b100 *
0-
02
b100 6
#720730000000
1!
1%
1-
12
#720740000000
0!
0%
b101 *
0-
02
b101 6
#720750000000
1!
1%
1-
12
#720760000000
0!
0%
b110 *
0-
02
b110 6
#720770000000
1!
1%
1-
12
#720780000000
0!
0%
b111 *
0-
02
b111 6
#720790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#720800000000
0!
0%
b0 *
0-
02
b0 6
#720810000000
1!
1%
1-
12
#720820000000
0!
0%
b1 *
0-
02
b1 6
#720830000000
1!
1%
1-
12
#720840000000
0!
0%
b10 *
0-
02
b10 6
#720850000000
1!
1%
1-
12
#720860000000
0!
0%
b11 *
0-
02
b11 6
#720870000000
1!
1%
1-
12
15
#720880000000
0!
0%
b100 *
0-
02
b100 6
#720890000000
1!
1%
1-
12
#720900000000
0!
0%
b101 *
0-
02
b101 6
#720910000000
1!
1%
1-
12
#720920000000
0!
0%
b110 *
0-
02
b110 6
#720930000000
1!
1%
1-
12
#720940000000
0!
0%
b111 *
0-
02
b111 6
#720950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#720960000000
0!
0%
b0 *
0-
02
b0 6
#720970000000
1!
1%
1-
12
#720980000000
0!
0%
b1 *
0-
02
b1 6
#720990000000
1!
1%
1-
12
#721000000000
0!
0%
b10 *
0-
02
b10 6
#721010000000
1!
1%
1-
12
#721020000000
0!
0%
b11 *
0-
02
b11 6
#721030000000
1!
1%
1-
12
15
#721040000000
0!
0%
b100 *
0-
02
b100 6
#721050000000
1!
1%
1-
12
#721060000000
0!
0%
b101 *
0-
02
b101 6
#721070000000
1!
1%
1-
12
#721080000000
0!
0%
b110 *
0-
02
b110 6
#721090000000
1!
1%
1-
12
#721100000000
0!
0%
b111 *
0-
02
b111 6
#721110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#721120000000
0!
0%
b0 *
0-
02
b0 6
#721130000000
1!
1%
1-
12
#721140000000
0!
0%
b1 *
0-
02
b1 6
#721150000000
1!
1%
1-
12
#721160000000
0!
0%
b10 *
0-
02
b10 6
#721170000000
1!
1%
1-
12
#721180000000
0!
0%
b11 *
0-
02
b11 6
#721190000000
1!
1%
1-
12
15
#721200000000
0!
0%
b100 *
0-
02
b100 6
#721210000000
1!
1%
1-
12
#721220000000
0!
0%
b101 *
0-
02
b101 6
#721230000000
1!
1%
1-
12
#721240000000
0!
0%
b110 *
0-
02
b110 6
#721250000000
1!
1%
1-
12
#721260000000
0!
0%
b111 *
0-
02
b111 6
#721270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#721280000000
0!
0%
b0 *
0-
02
b0 6
#721290000000
1!
1%
1-
12
#721300000000
0!
0%
b1 *
0-
02
b1 6
#721310000000
1!
1%
1-
12
#721320000000
0!
0%
b10 *
0-
02
b10 6
#721330000000
1!
1%
1-
12
#721340000000
0!
0%
b11 *
0-
02
b11 6
#721350000000
1!
1%
1-
12
15
#721360000000
0!
0%
b100 *
0-
02
b100 6
#721370000000
1!
1%
1-
12
#721380000000
0!
0%
b101 *
0-
02
b101 6
#721390000000
1!
1%
1-
12
#721400000000
0!
0%
b110 *
0-
02
b110 6
#721410000000
1!
1%
1-
12
#721420000000
0!
0%
b111 *
0-
02
b111 6
#721430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#721440000000
0!
0%
b0 *
0-
02
b0 6
#721450000000
1!
1%
1-
12
#721460000000
0!
0%
b1 *
0-
02
b1 6
#721470000000
1!
1%
1-
12
#721480000000
0!
0%
b10 *
0-
02
b10 6
#721490000000
1!
1%
1-
12
#721500000000
0!
0%
b11 *
0-
02
b11 6
#721510000000
1!
1%
1-
12
15
#721520000000
0!
0%
b100 *
0-
02
b100 6
#721530000000
1!
1%
1-
12
#721540000000
0!
0%
b101 *
0-
02
b101 6
#721550000000
1!
1%
1-
12
#721560000000
0!
0%
b110 *
0-
02
b110 6
#721570000000
1!
1%
1-
12
#721580000000
0!
0%
b111 *
0-
02
b111 6
#721590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#721600000000
0!
0%
b0 *
0-
02
b0 6
#721610000000
1!
1%
1-
12
#721620000000
0!
0%
b1 *
0-
02
b1 6
#721630000000
1!
1%
1-
12
#721640000000
0!
0%
b10 *
0-
02
b10 6
#721650000000
1!
1%
1-
12
#721660000000
0!
0%
b11 *
0-
02
b11 6
#721670000000
1!
1%
1-
12
15
#721680000000
0!
0%
b100 *
0-
02
b100 6
#721690000000
1!
1%
1-
12
#721700000000
0!
0%
b101 *
0-
02
b101 6
#721710000000
1!
1%
1-
12
#721720000000
0!
0%
b110 *
0-
02
b110 6
#721730000000
1!
1%
1-
12
#721740000000
0!
0%
b111 *
0-
02
b111 6
#721750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#721760000000
0!
0%
b0 *
0-
02
b0 6
#721770000000
1!
1%
1-
12
#721780000000
0!
0%
b1 *
0-
02
b1 6
#721790000000
1!
1%
1-
12
#721800000000
0!
0%
b10 *
0-
02
b10 6
#721810000000
1!
1%
1-
12
#721820000000
0!
0%
b11 *
0-
02
b11 6
#721830000000
1!
1%
1-
12
15
#721840000000
0!
0%
b100 *
0-
02
b100 6
#721850000000
1!
1%
1-
12
#721860000000
0!
0%
b101 *
0-
02
b101 6
#721870000000
1!
1%
1-
12
#721880000000
0!
0%
b110 *
0-
02
b110 6
#721890000000
1!
1%
1-
12
#721900000000
0!
0%
b111 *
0-
02
b111 6
#721910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#721920000000
0!
0%
b0 *
0-
02
b0 6
#721930000000
1!
1%
1-
12
#721940000000
0!
0%
b1 *
0-
02
b1 6
#721950000000
1!
1%
1-
12
#721960000000
0!
0%
b10 *
0-
02
b10 6
#721970000000
1!
1%
1-
12
#721980000000
0!
0%
b11 *
0-
02
b11 6
#721990000000
1!
1%
1-
12
15
#722000000000
0!
0%
b100 *
0-
02
b100 6
#722010000000
1!
1%
1-
12
#722020000000
0!
0%
b101 *
0-
02
b101 6
#722030000000
1!
1%
1-
12
#722040000000
0!
0%
b110 *
0-
02
b110 6
#722050000000
1!
1%
1-
12
#722060000000
0!
0%
b111 *
0-
02
b111 6
#722070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#722080000000
0!
0%
b0 *
0-
02
b0 6
#722090000000
1!
1%
1-
12
#722100000000
0!
0%
b1 *
0-
02
b1 6
#722110000000
1!
1%
1-
12
#722120000000
0!
0%
b10 *
0-
02
b10 6
#722130000000
1!
1%
1-
12
#722140000000
0!
0%
b11 *
0-
02
b11 6
#722150000000
1!
1%
1-
12
15
#722160000000
0!
0%
b100 *
0-
02
b100 6
#722170000000
1!
1%
1-
12
#722180000000
0!
0%
b101 *
0-
02
b101 6
#722190000000
1!
1%
1-
12
#722200000000
0!
0%
b110 *
0-
02
b110 6
#722210000000
1!
1%
1-
12
#722220000000
0!
0%
b111 *
0-
02
b111 6
#722230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#722240000000
0!
0%
b0 *
0-
02
b0 6
#722250000000
1!
1%
1-
12
#722260000000
0!
0%
b1 *
0-
02
b1 6
#722270000000
1!
1%
1-
12
#722280000000
0!
0%
b10 *
0-
02
b10 6
#722290000000
1!
1%
1-
12
#722300000000
0!
0%
b11 *
0-
02
b11 6
#722310000000
1!
1%
1-
12
15
#722320000000
0!
0%
b100 *
0-
02
b100 6
#722330000000
1!
1%
1-
12
#722340000000
0!
0%
b101 *
0-
02
b101 6
#722350000000
1!
1%
1-
12
#722360000000
0!
0%
b110 *
0-
02
b110 6
#722370000000
1!
1%
1-
12
#722380000000
0!
0%
b111 *
0-
02
b111 6
#722390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#722400000000
0!
0%
b0 *
0-
02
b0 6
#722410000000
1!
1%
1-
12
#722420000000
0!
0%
b1 *
0-
02
b1 6
#722430000000
1!
1%
1-
12
#722440000000
0!
0%
b10 *
0-
02
b10 6
#722450000000
1!
1%
1-
12
#722460000000
0!
0%
b11 *
0-
02
b11 6
#722470000000
1!
1%
1-
12
15
#722480000000
0!
0%
b100 *
0-
02
b100 6
#722490000000
1!
1%
1-
12
#722500000000
0!
0%
b101 *
0-
02
b101 6
#722510000000
1!
1%
1-
12
#722520000000
0!
0%
b110 *
0-
02
b110 6
#722530000000
1!
1%
1-
12
#722540000000
0!
0%
b111 *
0-
02
b111 6
#722550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#722560000000
0!
0%
b0 *
0-
02
b0 6
#722570000000
1!
1%
1-
12
#722580000000
0!
0%
b1 *
0-
02
b1 6
#722590000000
1!
1%
1-
12
#722600000000
0!
0%
b10 *
0-
02
b10 6
#722610000000
1!
1%
1-
12
#722620000000
0!
0%
b11 *
0-
02
b11 6
#722630000000
1!
1%
1-
12
15
#722640000000
0!
0%
b100 *
0-
02
b100 6
#722650000000
1!
1%
1-
12
#722660000000
0!
0%
b101 *
0-
02
b101 6
#722670000000
1!
1%
1-
12
#722680000000
0!
0%
b110 *
0-
02
b110 6
#722690000000
1!
1%
1-
12
#722700000000
0!
0%
b111 *
0-
02
b111 6
#722710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#722720000000
0!
0%
b0 *
0-
02
b0 6
#722730000000
1!
1%
1-
12
#722740000000
0!
0%
b1 *
0-
02
b1 6
#722750000000
1!
1%
1-
12
#722760000000
0!
0%
b10 *
0-
02
b10 6
#722770000000
1!
1%
1-
12
#722780000000
0!
0%
b11 *
0-
02
b11 6
#722790000000
1!
1%
1-
12
15
#722800000000
0!
0%
b100 *
0-
02
b100 6
#722810000000
1!
1%
1-
12
#722820000000
0!
0%
b101 *
0-
02
b101 6
#722830000000
1!
1%
1-
12
#722840000000
0!
0%
b110 *
0-
02
b110 6
#722850000000
1!
1%
1-
12
#722860000000
0!
0%
b111 *
0-
02
b111 6
#722870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#722880000000
0!
0%
b0 *
0-
02
b0 6
#722890000000
1!
1%
1-
12
#722900000000
0!
0%
b1 *
0-
02
b1 6
#722910000000
1!
1%
1-
12
#722920000000
0!
0%
b10 *
0-
02
b10 6
#722930000000
1!
1%
1-
12
#722940000000
0!
0%
b11 *
0-
02
b11 6
#722950000000
1!
1%
1-
12
15
#722960000000
0!
0%
b100 *
0-
02
b100 6
#722970000000
1!
1%
1-
12
#722980000000
0!
0%
b101 *
0-
02
b101 6
#722990000000
1!
1%
1-
12
#723000000000
0!
0%
b110 *
0-
02
b110 6
#723010000000
1!
1%
1-
12
#723020000000
0!
0%
b111 *
0-
02
b111 6
#723030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#723040000000
0!
0%
b0 *
0-
02
b0 6
#723050000000
1!
1%
1-
12
#723060000000
0!
0%
b1 *
0-
02
b1 6
#723070000000
1!
1%
1-
12
#723080000000
0!
0%
b10 *
0-
02
b10 6
#723090000000
1!
1%
1-
12
#723100000000
0!
0%
b11 *
0-
02
b11 6
#723110000000
1!
1%
1-
12
15
#723120000000
0!
0%
b100 *
0-
02
b100 6
#723130000000
1!
1%
1-
12
#723140000000
0!
0%
b101 *
0-
02
b101 6
#723150000000
1!
1%
1-
12
#723160000000
0!
0%
b110 *
0-
02
b110 6
#723170000000
1!
1%
1-
12
#723180000000
0!
0%
b111 *
0-
02
b111 6
#723190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#723200000000
0!
0%
b0 *
0-
02
b0 6
#723210000000
1!
1%
1-
12
#723220000000
0!
0%
b1 *
0-
02
b1 6
#723230000000
1!
1%
1-
12
#723240000000
0!
0%
b10 *
0-
02
b10 6
#723250000000
1!
1%
1-
12
#723260000000
0!
0%
b11 *
0-
02
b11 6
#723270000000
1!
1%
1-
12
15
#723280000000
0!
0%
b100 *
0-
02
b100 6
#723290000000
1!
1%
1-
12
#723300000000
0!
0%
b101 *
0-
02
b101 6
#723310000000
1!
1%
1-
12
#723320000000
0!
0%
b110 *
0-
02
b110 6
#723330000000
1!
1%
1-
12
#723340000000
0!
0%
b111 *
0-
02
b111 6
#723350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#723360000000
0!
0%
b0 *
0-
02
b0 6
#723370000000
1!
1%
1-
12
#723380000000
0!
0%
b1 *
0-
02
b1 6
#723390000000
1!
1%
1-
12
#723400000000
0!
0%
b10 *
0-
02
b10 6
#723410000000
1!
1%
1-
12
#723420000000
0!
0%
b11 *
0-
02
b11 6
#723430000000
1!
1%
1-
12
15
#723440000000
0!
0%
b100 *
0-
02
b100 6
#723450000000
1!
1%
1-
12
#723460000000
0!
0%
b101 *
0-
02
b101 6
#723470000000
1!
1%
1-
12
#723480000000
0!
0%
b110 *
0-
02
b110 6
#723490000000
1!
1%
1-
12
#723500000000
0!
0%
b111 *
0-
02
b111 6
#723510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#723520000000
0!
0%
b0 *
0-
02
b0 6
#723530000000
1!
1%
1-
12
#723540000000
0!
0%
b1 *
0-
02
b1 6
#723550000000
1!
1%
1-
12
#723560000000
0!
0%
b10 *
0-
02
b10 6
#723570000000
1!
1%
1-
12
#723580000000
0!
0%
b11 *
0-
02
b11 6
#723590000000
1!
1%
1-
12
15
#723600000000
0!
0%
b100 *
0-
02
b100 6
#723610000000
1!
1%
1-
12
#723620000000
0!
0%
b101 *
0-
02
b101 6
#723630000000
1!
1%
1-
12
#723640000000
0!
0%
b110 *
0-
02
b110 6
#723650000000
1!
1%
1-
12
#723660000000
0!
0%
b111 *
0-
02
b111 6
#723670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#723680000000
0!
0%
b0 *
0-
02
b0 6
#723690000000
1!
1%
1-
12
#723700000000
0!
0%
b1 *
0-
02
b1 6
#723710000000
1!
1%
1-
12
#723720000000
0!
0%
b10 *
0-
02
b10 6
#723730000000
1!
1%
1-
12
#723740000000
0!
0%
b11 *
0-
02
b11 6
#723750000000
1!
1%
1-
12
15
#723760000000
0!
0%
b100 *
0-
02
b100 6
#723770000000
1!
1%
1-
12
#723780000000
0!
0%
b101 *
0-
02
b101 6
#723790000000
1!
1%
1-
12
#723800000000
0!
0%
b110 *
0-
02
b110 6
#723810000000
1!
1%
1-
12
#723820000000
0!
0%
b111 *
0-
02
b111 6
#723830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#723840000000
0!
0%
b0 *
0-
02
b0 6
#723850000000
1!
1%
1-
12
#723860000000
0!
0%
b1 *
0-
02
b1 6
#723870000000
1!
1%
1-
12
#723880000000
0!
0%
b10 *
0-
02
b10 6
#723890000000
1!
1%
1-
12
#723900000000
0!
0%
b11 *
0-
02
b11 6
#723910000000
1!
1%
1-
12
15
#723920000000
0!
0%
b100 *
0-
02
b100 6
#723930000000
1!
1%
1-
12
#723940000000
0!
0%
b101 *
0-
02
b101 6
#723950000000
1!
1%
1-
12
#723960000000
0!
0%
b110 *
0-
02
b110 6
#723970000000
1!
1%
1-
12
#723980000000
0!
0%
b111 *
0-
02
b111 6
#723990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#724000000000
0!
0%
b0 *
0-
02
b0 6
#724010000000
1!
1%
1-
12
#724020000000
0!
0%
b1 *
0-
02
b1 6
#724030000000
1!
1%
1-
12
#724040000000
0!
0%
b10 *
0-
02
b10 6
#724050000000
1!
1%
1-
12
#724060000000
0!
0%
b11 *
0-
02
b11 6
#724070000000
1!
1%
1-
12
15
#724080000000
0!
0%
b100 *
0-
02
b100 6
#724090000000
1!
1%
1-
12
#724100000000
0!
0%
b101 *
0-
02
b101 6
#724110000000
1!
1%
1-
12
#724120000000
0!
0%
b110 *
0-
02
b110 6
#724130000000
1!
1%
1-
12
#724140000000
0!
0%
b111 *
0-
02
b111 6
#724150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#724160000000
0!
0%
b0 *
0-
02
b0 6
#724170000000
1!
1%
1-
12
#724180000000
0!
0%
b1 *
0-
02
b1 6
#724190000000
1!
1%
1-
12
#724200000000
0!
0%
b10 *
0-
02
b10 6
#724210000000
1!
1%
1-
12
#724220000000
0!
0%
b11 *
0-
02
b11 6
#724230000000
1!
1%
1-
12
15
#724240000000
0!
0%
b100 *
0-
02
b100 6
#724250000000
1!
1%
1-
12
#724260000000
0!
0%
b101 *
0-
02
b101 6
#724270000000
1!
1%
1-
12
#724280000000
0!
0%
b110 *
0-
02
b110 6
#724290000000
1!
1%
1-
12
#724300000000
0!
0%
b111 *
0-
02
b111 6
#724310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#724320000000
0!
0%
b0 *
0-
02
b0 6
#724330000000
1!
1%
1-
12
#724340000000
0!
0%
b1 *
0-
02
b1 6
#724350000000
1!
1%
1-
12
#724360000000
0!
0%
b10 *
0-
02
b10 6
#724370000000
1!
1%
1-
12
#724380000000
0!
0%
b11 *
0-
02
b11 6
#724390000000
1!
1%
1-
12
15
#724400000000
0!
0%
b100 *
0-
02
b100 6
#724410000000
1!
1%
1-
12
#724420000000
0!
0%
b101 *
0-
02
b101 6
#724430000000
1!
1%
1-
12
#724440000000
0!
0%
b110 *
0-
02
b110 6
#724450000000
1!
1%
1-
12
#724460000000
0!
0%
b111 *
0-
02
b111 6
#724470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#724480000000
0!
0%
b0 *
0-
02
b0 6
#724490000000
1!
1%
1-
12
#724500000000
0!
0%
b1 *
0-
02
b1 6
#724510000000
1!
1%
1-
12
#724520000000
0!
0%
b10 *
0-
02
b10 6
#724530000000
1!
1%
1-
12
#724540000000
0!
0%
b11 *
0-
02
b11 6
#724550000000
1!
1%
1-
12
15
#724560000000
0!
0%
b100 *
0-
02
b100 6
#724570000000
1!
1%
1-
12
#724580000000
0!
0%
b101 *
0-
02
b101 6
#724590000000
1!
1%
1-
12
#724600000000
0!
0%
b110 *
0-
02
b110 6
#724610000000
1!
1%
1-
12
#724620000000
0!
0%
b111 *
0-
02
b111 6
#724630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#724640000000
0!
0%
b0 *
0-
02
b0 6
#724650000000
1!
1%
1-
12
#724660000000
0!
0%
b1 *
0-
02
b1 6
#724670000000
1!
1%
1-
12
#724680000000
0!
0%
b10 *
0-
02
b10 6
#724690000000
1!
1%
1-
12
#724700000000
0!
0%
b11 *
0-
02
b11 6
#724710000000
1!
1%
1-
12
15
#724720000000
0!
0%
b100 *
0-
02
b100 6
#724730000000
1!
1%
1-
12
#724740000000
0!
0%
b101 *
0-
02
b101 6
#724750000000
1!
1%
1-
12
#724760000000
0!
0%
b110 *
0-
02
b110 6
#724770000000
1!
1%
1-
12
#724780000000
0!
0%
b111 *
0-
02
b111 6
#724790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#724800000000
0!
0%
b0 *
0-
02
b0 6
#724810000000
1!
1%
1-
12
#724820000000
0!
0%
b1 *
0-
02
b1 6
#724830000000
1!
1%
1-
12
#724840000000
0!
0%
b10 *
0-
02
b10 6
#724850000000
1!
1%
1-
12
#724860000000
0!
0%
b11 *
0-
02
b11 6
#724870000000
1!
1%
1-
12
15
#724880000000
0!
0%
b100 *
0-
02
b100 6
#724890000000
1!
1%
1-
12
#724900000000
0!
0%
b101 *
0-
02
b101 6
#724910000000
1!
1%
1-
12
#724920000000
0!
0%
b110 *
0-
02
b110 6
#724930000000
1!
1%
1-
12
#724940000000
0!
0%
b111 *
0-
02
b111 6
#724950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#724960000000
0!
0%
b0 *
0-
02
b0 6
#724970000000
1!
1%
1-
12
#724980000000
0!
0%
b1 *
0-
02
b1 6
#724990000000
1!
1%
1-
12
#725000000000
0!
0%
b10 *
0-
02
b10 6
#725010000000
1!
1%
1-
12
#725020000000
0!
0%
b11 *
0-
02
b11 6
#725030000000
1!
1%
1-
12
15
#725040000000
0!
0%
b100 *
0-
02
b100 6
#725050000000
1!
1%
1-
12
#725060000000
0!
0%
b101 *
0-
02
b101 6
#725070000000
1!
1%
1-
12
#725080000000
0!
0%
b110 *
0-
02
b110 6
#725090000000
1!
1%
1-
12
#725100000000
0!
0%
b111 *
0-
02
b111 6
#725110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#725120000000
0!
0%
b0 *
0-
02
b0 6
#725130000000
1!
1%
1-
12
#725140000000
0!
0%
b1 *
0-
02
b1 6
#725150000000
1!
1%
1-
12
#725160000000
0!
0%
b10 *
0-
02
b10 6
#725170000000
1!
1%
1-
12
#725180000000
0!
0%
b11 *
0-
02
b11 6
#725190000000
1!
1%
1-
12
15
#725200000000
0!
0%
b100 *
0-
02
b100 6
#725210000000
1!
1%
1-
12
#725220000000
0!
0%
b101 *
0-
02
b101 6
#725230000000
1!
1%
1-
12
#725240000000
0!
0%
b110 *
0-
02
b110 6
#725250000000
1!
1%
1-
12
#725260000000
0!
0%
b111 *
0-
02
b111 6
#725270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#725280000000
0!
0%
b0 *
0-
02
b0 6
#725290000000
1!
1%
1-
12
#725300000000
0!
0%
b1 *
0-
02
b1 6
#725310000000
1!
1%
1-
12
#725320000000
0!
0%
b10 *
0-
02
b10 6
#725330000000
1!
1%
1-
12
#725340000000
0!
0%
b11 *
0-
02
b11 6
#725350000000
1!
1%
1-
12
15
#725360000000
0!
0%
b100 *
0-
02
b100 6
#725370000000
1!
1%
1-
12
#725380000000
0!
0%
b101 *
0-
02
b101 6
#725390000000
1!
1%
1-
12
#725400000000
0!
0%
b110 *
0-
02
b110 6
#725410000000
1!
1%
1-
12
#725420000000
0!
0%
b111 *
0-
02
b111 6
#725430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#725440000000
0!
0%
b0 *
0-
02
b0 6
#725450000000
1!
1%
1-
12
#725460000000
0!
0%
b1 *
0-
02
b1 6
#725470000000
1!
1%
1-
12
#725480000000
0!
0%
b10 *
0-
02
b10 6
#725490000000
1!
1%
1-
12
#725500000000
0!
0%
b11 *
0-
02
b11 6
#725510000000
1!
1%
1-
12
15
#725520000000
0!
0%
b100 *
0-
02
b100 6
#725530000000
1!
1%
1-
12
#725540000000
0!
0%
b101 *
0-
02
b101 6
#725550000000
1!
1%
1-
12
#725560000000
0!
0%
b110 *
0-
02
b110 6
#725570000000
1!
1%
1-
12
#725580000000
0!
0%
b111 *
0-
02
b111 6
#725590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#725600000000
0!
0%
b0 *
0-
02
b0 6
#725610000000
1!
1%
1-
12
#725620000000
0!
0%
b1 *
0-
02
b1 6
#725630000000
1!
1%
1-
12
#725640000000
0!
0%
b10 *
0-
02
b10 6
#725650000000
1!
1%
1-
12
#725660000000
0!
0%
b11 *
0-
02
b11 6
#725670000000
1!
1%
1-
12
15
#725680000000
0!
0%
b100 *
0-
02
b100 6
#725690000000
1!
1%
1-
12
#725700000000
0!
0%
b101 *
0-
02
b101 6
#725710000000
1!
1%
1-
12
#725720000000
0!
0%
b110 *
0-
02
b110 6
#725730000000
1!
1%
1-
12
#725740000000
0!
0%
b111 *
0-
02
b111 6
#725750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#725760000000
0!
0%
b0 *
0-
02
b0 6
#725770000000
1!
1%
1-
12
#725780000000
0!
0%
b1 *
0-
02
b1 6
#725790000000
1!
1%
1-
12
#725800000000
0!
0%
b10 *
0-
02
b10 6
#725810000000
1!
1%
1-
12
#725820000000
0!
0%
b11 *
0-
02
b11 6
#725830000000
1!
1%
1-
12
15
#725840000000
0!
0%
b100 *
0-
02
b100 6
#725850000000
1!
1%
1-
12
#725860000000
0!
0%
b101 *
0-
02
b101 6
#725870000000
1!
1%
1-
12
#725880000000
0!
0%
b110 *
0-
02
b110 6
#725890000000
1!
1%
1-
12
#725900000000
0!
0%
b111 *
0-
02
b111 6
#725910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#725920000000
0!
0%
b0 *
0-
02
b0 6
#725930000000
1!
1%
1-
12
#725940000000
0!
0%
b1 *
0-
02
b1 6
#725950000000
1!
1%
1-
12
#725960000000
0!
0%
b10 *
0-
02
b10 6
#725970000000
1!
1%
1-
12
#725980000000
0!
0%
b11 *
0-
02
b11 6
#725990000000
1!
1%
1-
12
15
#726000000000
0!
0%
b100 *
0-
02
b100 6
#726010000000
1!
1%
1-
12
#726020000000
0!
0%
b101 *
0-
02
b101 6
#726030000000
1!
1%
1-
12
#726040000000
0!
0%
b110 *
0-
02
b110 6
#726050000000
1!
1%
1-
12
#726060000000
0!
0%
b111 *
0-
02
b111 6
#726070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#726080000000
0!
0%
b0 *
0-
02
b0 6
#726090000000
1!
1%
1-
12
#726100000000
0!
0%
b1 *
0-
02
b1 6
#726110000000
1!
1%
1-
12
#726120000000
0!
0%
b10 *
0-
02
b10 6
#726130000000
1!
1%
1-
12
#726140000000
0!
0%
b11 *
0-
02
b11 6
#726150000000
1!
1%
1-
12
15
#726160000000
0!
0%
b100 *
0-
02
b100 6
#726170000000
1!
1%
1-
12
#726180000000
0!
0%
b101 *
0-
02
b101 6
#726190000000
1!
1%
1-
12
#726200000000
0!
0%
b110 *
0-
02
b110 6
#726210000000
1!
1%
1-
12
#726220000000
0!
0%
b111 *
0-
02
b111 6
#726230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#726240000000
0!
0%
b0 *
0-
02
b0 6
#726250000000
1!
1%
1-
12
#726260000000
0!
0%
b1 *
0-
02
b1 6
#726270000000
1!
1%
1-
12
#726280000000
0!
0%
b10 *
0-
02
b10 6
#726290000000
1!
1%
1-
12
#726300000000
0!
0%
b11 *
0-
02
b11 6
#726310000000
1!
1%
1-
12
15
#726320000000
0!
0%
b100 *
0-
02
b100 6
#726330000000
1!
1%
1-
12
#726340000000
0!
0%
b101 *
0-
02
b101 6
#726350000000
1!
1%
1-
12
#726360000000
0!
0%
b110 *
0-
02
b110 6
#726370000000
1!
1%
1-
12
#726380000000
0!
0%
b111 *
0-
02
b111 6
#726390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#726400000000
0!
0%
b0 *
0-
02
b0 6
#726410000000
1!
1%
1-
12
#726420000000
0!
0%
b1 *
0-
02
b1 6
#726430000000
1!
1%
1-
12
#726440000000
0!
0%
b10 *
0-
02
b10 6
#726450000000
1!
1%
1-
12
#726460000000
0!
0%
b11 *
0-
02
b11 6
#726470000000
1!
1%
1-
12
15
#726480000000
0!
0%
b100 *
0-
02
b100 6
#726490000000
1!
1%
1-
12
#726500000000
0!
0%
b101 *
0-
02
b101 6
#726510000000
1!
1%
1-
12
#726520000000
0!
0%
b110 *
0-
02
b110 6
#726530000000
1!
1%
1-
12
#726540000000
0!
0%
b111 *
0-
02
b111 6
#726550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#726560000000
0!
0%
b0 *
0-
02
b0 6
#726570000000
1!
1%
1-
12
#726580000000
0!
0%
b1 *
0-
02
b1 6
#726590000000
1!
1%
1-
12
#726600000000
0!
0%
b10 *
0-
02
b10 6
#726610000000
1!
1%
1-
12
#726620000000
0!
0%
b11 *
0-
02
b11 6
#726630000000
1!
1%
1-
12
15
#726640000000
0!
0%
b100 *
0-
02
b100 6
#726650000000
1!
1%
1-
12
#726660000000
0!
0%
b101 *
0-
02
b101 6
#726670000000
1!
1%
1-
12
#726680000000
0!
0%
b110 *
0-
02
b110 6
#726690000000
1!
1%
1-
12
#726700000000
0!
0%
b111 *
0-
02
b111 6
#726710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#726720000000
0!
0%
b0 *
0-
02
b0 6
#726730000000
1!
1%
1-
12
#726740000000
0!
0%
b1 *
0-
02
b1 6
#726750000000
1!
1%
1-
12
#726760000000
0!
0%
b10 *
0-
02
b10 6
#726770000000
1!
1%
1-
12
#726780000000
0!
0%
b11 *
0-
02
b11 6
#726790000000
1!
1%
1-
12
15
#726800000000
0!
0%
b100 *
0-
02
b100 6
#726810000000
1!
1%
1-
12
#726820000000
0!
0%
b101 *
0-
02
b101 6
#726830000000
1!
1%
1-
12
#726840000000
0!
0%
b110 *
0-
02
b110 6
#726850000000
1!
1%
1-
12
#726860000000
0!
0%
b111 *
0-
02
b111 6
#726870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#726880000000
0!
0%
b0 *
0-
02
b0 6
#726890000000
1!
1%
1-
12
#726900000000
0!
0%
b1 *
0-
02
b1 6
#726910000000
1!
1%
1-
12
#726920000000
0!
0%
b10 *
0-
02
b10 6
#726930000000
1!
1%
1-
12
#726940000000
0!
0%
b11 *
0-
02
b11 6
#726950000000
1!
1%
1-
12
15
#726960000000
0!
0%
b100 *
0-
02
b100 6
#726970000000
1!
1%
1-
12
#726980000000
0!
0%
b101 *
0-
02
b101 6
#726990000000
1!
1%
1-
12
#727000000000
0!
0%
b110 *
0-
02
b110 6
#727010000000
1!
1%
1-
12
#727020000000
0!
0%
b111 *
0-
02
b111 6
#727030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#727040000000
0!
0%
b0 *
0-
02
b0 6
#727050000000
1!
1%
1-
12
#727060000000
0!
0%
b1 *
0-
02
b1 6
#727070000000
1!
1%
1-
12
#727080000000
0!
0%
b10 *
0-
02
b10 6
#727090000000
1!
1%
1-
12
#727100000000
0!
0%
b11 *
0-
02
b11 6
#727110000000
1!
1%
1-
12
15
#727120000000
0!
0%
b100 *
0-
02
b100 6
#727130000000
1!
1%
1-
12
#727140000000
0!
0%
b101 *
0-
02
b101 6
#727150000000
1!
1%
1-
12
#727160000000
0!
0%
b110 *
0-
02
b110 6
#727170000000
1!
1%
1-
12
#727180000000
0!
0%
b111 *
0-
02
b111 6
#727190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#727200000000
0!
0%
b0 *
0-
02
b0 6
#727210000000
1!
1%
1-
12
#727220000000
0!
0%
b1 *
0-
02
b1 6
#727230000000
1!
1%
1-
12
#727240000000
0!
0%
b10 *
0-
02
b10 6
#727250000000
1!
1%
1-
12
#727260000000
0!
0%
b11 *
0-
02
b11 6
#727270000000
1!
1%
1-
12
15
#727280000000
0!
0%
b100 *
0-
02
b100 6
#727290000000
1!
1%
1-
12
#727300000000
0!
0%
b101 *
0-
02
b101 6
#727310000000
1!
1%
1-
12
#727320000000
0!
0%
b110 *
0-
02
b110 6
#727330000000
1!
1%
1-
12
#727340000000
0!
0%
b111 *
0-
02
b111 6
#727350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#727360000000
0!
0%
b0 *
0-
02
b0 6
#727370000000
1!
1%
1-
12
#727380000000
0!
0%
b1 *
0-
02
b1 6
#727390000000
1!
1%
1-
12
#727400000000
0!
0%
b10 *
0-
02
b10 6
#727410000000
1!
1%
1-
12
#727420000000
0!
0%
b11 *
0-
02
b11 6
#727430000000
1!
1%
1-
12
15
#727440000000
0!
0%
b100 *
0-
02
b100 6
#727450000000
1!
1%
1-
12
#727460000000
0!
0%
b101 *
0-
02
b101 6
#727470000000
1!
1%
1-
12
#727480000000
0!
0%
b110 *
0-
02
b110 6
#727490000000
1!
1%
1-
12
#727500000000
0!
0%
b111 *
0-
02
b111 6
#727510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#727520000000
0!
0%
b0 *
0-
02
b0 6
#727530000000
1!
1%
1-
12
#727540000000
0!
0%
b1 *
0-
02
b1 6
#727550000000
1!
1%
1-
12
#727560000000
0!
0%
b10 *
0-
02
b10 6
#727570000000
1!
1%
1-
12
#727580000000
0!
0%
b11 *
0-
02
b11 6
#727590000000
1!
1%
1-
12
15
#727600000000
0!
0%
b100 *
0-
02
b100 6
#727610000000
1!
1%
1-
12
#727620000000
0!
0%
b101 *
0-
02
b101 6
#727630000000
1!
1%
1-
12
#727640000000
0!
0%
b110 *
0-
02
b110 6
#727650000000
1!
1%
1-
12
#727660000000
0!
0%
b111 *
0-
02
b111 6
#727670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#727680000000
0!
0%
b0 *
0-
02
b0 6
#727690000000
1!
1%
1-
12
#727700000000
0!
0%
b1 *
0-
02
b1 6
#727710000000
1!
1%
1-
12
#727720000000
0!
0%
b10 *
0-
02
b10 6
#727730000000
1!
1%
1-
12
#727740000000
0!
0%
b11 *
0-
02
b11 6
#727750000000
1!
1%
1-
12
15
#727760000000
0!
0%
b100 *
0-
02
b100 6
#727770000000
1!
1%
1-
12
#727780000000
0!
0%
b101 *
0-
02
b101 6
#727790000000
1!
1%
1-
12
#727800000000
0!
0%
b110 *
0-
02
b110 6
#727810000000
1!
1%
1-
12
#727820000000
0!
0%
b111 *
0-
02
b111 6
#727830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#727840000000
0!
0%
b0 *
0-
02
b0 6
#727850000000
1!
1%
1-
12
#727860000000
0!
0%
b1 *
0-
02
b1 6
#727870000000
1!
1%
1-
12
#727880000000
0!
0%
b10 *
0-
02
b10 6
#727890000000
1!
1%
1-
12
#727900000000
0!
0%
b11 *
0-
02
b11 6
#727910000000
1!
1%
1-
12
15
#727920000000
0!
0%
b100 *
0-
02
b100 6
#727930000000
1!
1%
1-
12
#727940000000
0!
0%
b101 *
0-
02
b101 6
#727950000000
1!
1%
1-
12
#727960000000
0!
0%
b110 *
0-
02
b110 6
#727970000000
1!
1%
1-
12
#727980000000
0!
0%
b111 *
0-
02
b111 6
#727990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#728000000000
0!
0%
b0 *
0-
02
b0 6
#728010000000
1!
1%
1-
12
#728020000000
0!
0%
b1 *
0-
02
b1 6
#728030000000
1!
1%
1-
12
#728040000000
0!
0%
b10 *
0-
02
b10 6
#728050000000
1!
1%
1-
12
#728060000000
0!
0%
b11 *
0-
02
b11 6
#728070000000
1!
1%
1-
12
15
#728080000000
0!
0%
b100 *
0-
02
b100 6
#728090000000
1!
1%
1-
12
#728100000000
0!
0%
b101 *
0-
02
b101 6
#728110000000
1!
1%
1-
12
#728120000000
0!
0%
b110 *
0-
02
b110 6
#728130000000
1!
1%
1-
12
#728140000000
0!
0%
b111 *
0-
02
b111 6
#728150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#728160000000
0!
0%
b0 *
0-
02
b0 6
#728170000000
1!
1%
1-
12
#728180000000
0!
0%
b1 *
0-
02
b1 6
#728190000000
1!
1%
1-
12
#728200000000
0!
0%
b10 *
0-
02
b10 6
#728210000000
1!
1%
1-
12
#728220000000
0!
0%
b11 *
0-
02
b11 6
#728230000000
1!
1%
1-
12
15
#728240000000
0!
0%
b100 *
0-
02
b100 6
#728250000000
1!
1%
1-
12
#728260000000
0!
0%
b101 *
0-
02
b101 6
#728270000000
1!
1%
1-
12
#728280000000
0!
0%
b110 *
0-
02
b110 6
#728290000000
1!
1%
1-
12
#728300000000
0!
0%
b111 *
0-
02
b111 6
#728310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#728320000000
0!
0%
b0 *
0-
02
b0 6
#728330000000
1!
1%
1-
12
#728340000000
0!
0%
b1 *
0-
02
b1 6
#728350000000
1!
1%
1-
12
#728360000000
0!
0%
b10 *
0-
02
b10 6
#728370000000
1!
1%
1-
12
#728380000000
0!
0%
b11 *
0-
02
b11 6
#728390000000
1!
1%
1-
12
15
#728400000000
0!
0%
b100 *
0-
02
b100 6
#728410000000
1!
1%
1-
12
#728420000000
0!
0%
b101 *
0-
02
b101 6
#728430000000
1!
1%
1-
12
#728440000000
0!
0%
b110 *
0-
02
b110 6
#728450000000
1!
1%
1-
12
#728460000000
0!
0%
b111 *
0-
02
b111 6
#728470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#728480000000
0!
0%
b0 *
0-
02
b0 6
#728490000000
1!
1%
1-
12
#728500000000
0!
0%
b1 *
0-
02
b1 6
#728510000000
1!
1%
1-
12
#728520000000
0!
0%
b10 *
0-
02
b10 6
#728530000000
1!
1%
1-
12
#728540000000
0!
0%
b11 *
0-
02
b11 6
#728550000000
1!
1%
1-
12
15
#728560000000
0!
0%
b100 *
0-
02
b100 6
#728570000000
1!
1%
1-
12
#728580000000
0!
0%
b101 *
0-
02
b101 6
#728590000000
1!
1%
1-
12
#728600000000
0!
0%
b110 *
0-
02
b110 6
#728610000000
1!
1%
1-
12
#728620000000
0!
0%
b111 *
0-
02
b111 6
#728630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#728640000000
0!
0%
b0 *
0-
02
b0 6
#728650000000
1!
1%
1-
12
#728660000000
0!
0%
b1 *
0-
02
b1 6
#728670000000
1!
1%
1-
12
#728680000000
0!
0%
b10 *
0-
02
b10 6
#728690000000
1!
1%
1-
12
#728700000000
0!
0%
b11 *
0-
02
b11 6
#728710000000
1!
1%
1-
12
15
#728720000000
0!
0%
b100 *
0-
02
b100 6
#728730000000
1!
1%
1-
12
#728740000000
0!
0%
b101 *
0-
02
b101 6
#728750000000
1!
1%
1-
12
#728760000000
0!
0%
b110 *
0-
02
b110 6
#728770000000
1!
1%
1-
12
#728780000000
0!
0%
b111 *
0-
02
b111 6
#728790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#728800000000
0!
0%
b0 *
0-
02
b0 6
#728810000000
1!
1%
1-
12
#728820000000
0!
0%
b1 *
0-
02
b1 6
#728830000000
1!
1%
1-
12
#728840000000
0!
0%
b10 *
0-
02
b10 6
#728850000000
1!
1%
1-
12
#728860000000
0!
0%
b11 *
0-
02
b11 6
#728870000000
1!
1%
1-
12
15
#728880000000
0!
0%
b100 *
0-
02
b100 6
#728890000000
1!
1%
1-
12
#728900000000
0!
0%
b101 *
0-
02
b101 6
#728910000000
1!
1%
1-
12
#728920000000
0!
0%
b110 *
0-
02
b110 6
#728930000000
1!
1%
1-
12
#728940000000
0!
0%
b111 *
0-
02
b111 6
#728950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#728960000000
0!
0%
b0 *
0-
02
b0 6
#728970000000
1!
1%
1-
12
#728980000000
0!
0%
b1 *
0-
02
b1 6
#728990000000
1!
1%
1-
12
#729000000000
0!
0%
b10 *
0-
02
b10 6
#729010000000
1!
1%
1-
12
#729020000000
0!
0%
b11 *
0-
02
b11 6
#729030000000
1!
1%
1-
12
15
#729040000000
0!
0%
b100 *
0-
02
b100 6
#729050000000
1!
1%
1-
12
#729060000000
0!
0%
b101 *
0-
02
b101 6
#729070000000
1!
1%
1-
12
#729080000000
0!
0%
b110 *
0-
02
b110 6
#729090000000
1!
1%
1-
12
#729100000000
0!
0%
b111 *
0-
02
b111 6
#729110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#729120000000
0!
0%
b0 *
0-
02
b0 6
#729130000000
1!
1%
1-
12
#729140000000
0!
0%
b1 *
0-
02
b1 6
#729150000000
1!
1%
1-
12
#729160000000
0!
0%
b10 *
0-
02
b10 6
#729170000000
1!
1%
1-
12
#729180000000
0!
0%
b11 *
0-
02
b11 6
#729190000000
1!
1%
1-
12
15
#729200000000
0!
0%
b100 *
0-
02
b100 6
#729210000000
1!
1%
1-
12
#729220000000
0!
0%
b101 *
0-
02
b101 6
#729230000000
1!
1%
1-
12
#729240000000
0!
0%
b110 *
0-
02
b110 6
#729250000000
1!
1%
1-
12
#729260000000
0!
0%
b111 *
0-
02
b111 6
#729270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#729280000000
0!
0%
b0 *
0-
02
b0 6
#729290000000
1!
1%
1-
12
#729300000000
0!
0%
b1 *
0-
02
b1 6
#729310000000
1!
1%
1-
12
#729320000000
0!
0%
b10 *
0-
02
b10 6
#729330000000
1!
1%
1-
12
#729340000000
0!
0%
b11 *
0-
02
b11 6
#729350000000
1!
1%
1-
12
15
#729360000000
0!
0%
b100 *
0-
02
b100 6
#729370000000
1!
1%
1-
12
#729380000000
0!
0%
b101 *
0-
02
b101 6
#729390000000
1!
1%
1-
12
#729400000000
0!
0%
b110 *
0-
02
b110 6
#729410000000
1!
1%
1-
12
#729420000000
0!
0%
b111 *
0-
02
b111 6
#729430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#729440000000
0!
0%
b0 *
0-
02
b0 6
#729450000000
1!
1%
1-
12
#729460000000
0!
0%
b1 *
0-
02
b1 6
#729470000000
1!
1%
1-
12
#729480000000
0!
0%
b10 *
0-
02
b10 6
#729490000000
1!
1%
1-
12
#729500000000
0!
0%
b11 *
0-
02
b11 6
#729510000000
1!
1%
1-
12
15
#729520000000
0!
0%
b100 *
0-
02
b100 6
#729530000000
1!
1%
1-
12
#729540000000
0!
0%
b101 *
0-
02
b101 6
#729550000000
1!
1%
1-
12
#729560000000
0!
0%
b110 *
0-
02
b110 6
#729570000000
1!
1%
1-
12
#729580000000
0!
0%
b111 *
0-
02
b111 6
#729590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#729600000000
0!
0%
b0 *
0-
02
b0 6
#729610000000
1!
1%
1-
12
#729620000000
0!
0%
b1 *
0-
02
b1 6
#729630000000
1!
1%
1-
12
#729640000000
0!
0%
b10 *
0-
02
b10 6
#729650000000
1!
1%
1-
12
#729660000000
0!
0%
b11 *
0-
02
b11 6
#729670000000
1!
1%
1-
12
15
#729680000000
0!
0%
b100 *
0-
02
b100 6
#729690000000
1!
1%
1-
12
#729700000000
0!
0%
b101 *
0-
02
b101 6
#729710000000
1!
1%
1-
12
#729720000000
0!
0%
b110 *
0-
02
b110 6
#729730000000
1!
1%
1-
12
#729740000000
0!
0%
b111 *
0-
02
b111 6
#729750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#729760000000
0!
0%
b0 *
0-
02
b0 6
#729770000000
1!
1%
1-
12
#729780000000
0!
0%
b1 *
0-
02
b1 6
#729790000000
1!
1%
1-
12
#729800000000
0!
0%
b10 *
0-
02
b10 6
#729810000000
1!
1%
1-
12
#729820000000
0!
0%
b11 *
0-
02
b11 6
#729830000000
1!
1%
1-
12
15
#729840000000
0!
0%
b100 *
0-
02
b100 6
#729850000000
1!
1%
1-
12
#729860000000
0!
0%
b101 *
0-
02
b101 6
#729870000000
1!
1%
1-
12
#729880000000
0!
0%
b110 *
0-
02
b110 6
#729890000000
1!
1%
1-
12
#729900000000
0!
0%
b111 *
0-
02
b111 6
#729910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#729920000000
0!
0%
b0 *
0-
02
b0 6
#729930000000
1!
1%
1-
12
#729940000000
0!
0%
b1 *
0-
02
b1 6
#729950000000
1!
1%
1-
12
#729960000000
0!
0%
b10 *
0-
02
b10 6
#729970000000
1!
1%
1-
12
#729980000000
0!
0%
b11 *
0-
02
b11 6
#729990000000
1!
1%
1-
12
15
#730000000000
0!
0%
b100 *
0-
02
b100 6
#730010000000
1!
1%
1-
12
#730020000000
0!
0%
b101 *
0-
02
b101 6
#730030000000
1!
1%
1-
12
#730040000000
0!
0%
b110 *
0-
02
b110 6
#730050000000
1!
1%
1-
12
#730060000000
0!
0%
b111 *
0-
02
b111 6
#730070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#730080000000
0!
0%
b0 *
0-
02
b0 6
#730090000000
1!
1%
1-
12
#730100000000
0!
0%
b1 *
0-
02
b1 6
#730110000000
1!
1%
1-
12
#730120000000
0!
0%
b10 *
0-
02
b10 6
#730130000000
1!
1%
1-
12
#730140000000
0!
0%
b11 *
0-
02
b11 6
#730150000000
1!
1%
1-
12
15
#730160000000
0!
0%
b100 *
0-
02
b100 6
#730170000000
1!
1%
1-
12
#730180000000
0!
0%
b101 *
0-
02
b101 6
#730190000000
1!
1%
1-
12
#730200000000
0!
0%
b110 *
0-
02
b110 6
#730210000000
1!
1%
1-
12
#730220000000
0!
0%
b111 *
0-
02
b111 6
#730230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#730240000000
0!
0%
b0 *
0-
02
b0 6
#730250000000
1!
1%
1-
12
#730260000000
0!
0%
b1 *
0-
02
b1 6
#730270000000
1!
1%
1-
12
#730280000000
0!
0%
b10 *
0-
02
b10 6
#730290000000
1!
1%
1-
12
#730300000000
0!
0%
b11 *
0-
02
b11 6
#730310000000
1!
1%
1-
12
15
#730320000000
0!
0%
b100 *
0-
02
b100 6
#730330000000
1!
1%
1-
12
#730340000000
0!
0%
b101 *
0-
02
b101 6
#730350000000
1!
1%
1-
12
#730360000000
0!
0%
b110 *
0-
02
b110 6
#730370000000
1!
1%
1-
12
#730380000000
0!
0%
b111 *
0-
02
b111 6
#730390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#730400000000
0!
0%
b0 *
0-
02
b0 6
#730410000000
1!
1%
1-
12
#730420000000
0!
0%
b1 *
0-
02
b1 6
#730430000000
1!
1%
1-
12
#730440000000
0!
0%
b10 *
0-
02
b10 6
#730450000000
1!
1%
1-
12
#730460000000
0!
0%
b11 *
0-
02
b11 6
#730470000000
1!
1%
1-
12
15
#730480000000
0!
0%
b100 *
0-
02
b100 6
#730490000000
1!
1%
1-
12
#730500000000
0!
0%
b101 *
0-
02
b101 6
#730510000000
1!
1%
1-
12
#730520000000
0!
0%
b110 *
0-
02
b110 6
#730530000000
1!
1%
1-
12
#730540000000
0!
0%
b111 *
0-
02
b111 6
#730550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#730560000000
0!
0%
b0 *
0-
02
b0 6
#730570000000
1!
1%
1-
12
#730580000000
0!
0%
b1 *
0-
02
b1 6
#730590000000
1!
1%
1-
12
#730600000000
0!
0%
b10 *
0-
02
b10 6
#730610000000
1!
1%
1-
12
#730620000000
0!
0%
b11 *
0-
02
b11 6
#730630000000
1!
1%
1-
12
15
#730640000000
0!
0%
b100 *
0-
02
b100 6
#730650000000
1!
1%
1-
12
#730660000000
0!
0%
b101 *
0-
02
b101 6
#730670000000
1!
1%
1-
12
#730680000000
0!
0%
b110 *
0-
02
b110 6
#730690000000
1!
1%
1-
12
#730700000000
0!
0%
b111 *
0-
02
b111 6
#730710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#730720000000
0!
0%
b0 *
0-
02
b0 6
#730730000000
1!
1%
1-
12
#730740000000
0!
0%
b1 *
0-
02
b1 6
#730750000000
1!
1%
1-
12
#730760000000
0!
0%
b10 *
0-
02
b10 6
#730770000000
1!
1%
1-
12
#730780000000
0!
0%
b11 *
0-
02
b11 6
#730790000000
1!
1%
1-
12
15
#730800000000
0!
0%
b100 *
0-
02
b100 6
#730810000000
1!
1%
1-
12
#730820000000
0!
0%
b101 *
0-
02
b101 6
#730830000000
1!
1%
1-
12
#730840000000
0!
0%
b110 *
0-
02
b110 6
#730850000000
1!
1%
1-
12
#730860000000
0!
0%
b111 *
0-
02
b111 6
#730870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#730880000000
0!
0%
b0 *
0-
02
b0 6
#730890000000
1!
1%
1-
12
#730900000000
0!
0%
b1 *
0-
02
b1 6
#730910000000
1!
1%
1-
12
#730920000000
0!
0%
b10 *
0-
02
b10 6
#730930000000
1!
1%
1-
12
#730940000000
0!
0%
b11 *
0-
02
b11 6
#730950000000
1!
1%
1-
12
15
#730960000000
0!
0%
b100 *
0-
02
b100 6
#730970000000
1!
1%
1-
12
#730980000000
0!
0%
b101 *
0-
02
b101 6
#730990000000
1!
1%
1-
12
#731000000000
0!
0%
b110 *
0-
02
b110 6
#731010000000
1!
1%
1-
12
#731020000000
0!
0%
b111 *
0-
02
b111 6
#731030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#731040000000
0!
0%
b0 *
0-
02
b0 6
#731050000000
1!
1%
1-
12
#731060000000
0!
0%
b1 *
0-
02
b1 6
#731070000000
1!
1%
1-
12
#731080000000
0!
0%
b10 *
0-
02
b10 6
#731090000000
1!
1%
1-
12
#731100000000
0!
0%
b11 *
0-
02
b11 6
#731110000000
1!
1%
1-
12
15
#731120000000
0!
0%
b100 *
0-
02
b100 6
#731130000000
1!
1%
1-
12
#731140000000
0!
0%
b101 *
0-
02
b101 6
#731150000000
1!
1%
1-
12
#731160000000
0!
0%
b110 *
0-
02
b110 6
#731170000000
1!
1%
1-
12
#731180000000
0!
0%
b111 *
0-
02
b111 6
#731190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#731200000000
0!
0%
b0 *
0-
02
b0 6
#731210000000
1!
1%
1-
12
#731220000000
0!
0%
b1 *
0-
02
b1 6
#731230000000
1!
1%
1-
12
#731240000000
0!
0%
b10 *
0-
02
b10 6
#731250000000
1!
1%
1-
12
#731260000000
0!
0%
b11 *
0-
02
b11 6
#731270000000
1!
1%
1-
12
15
#731280000000
0!
0%
b100 *
0-
02
b100 6
#731290000000
1!
1%
1-
12
#731300000000
0!
0%
b101 *
0-
02
b101 6
#731310000000
1!
1%
1-
12
#731320000000
0!
0%
b110 *
0-
02
b110 6
#731330000000
1!
1%
1-
12
#731340000000
0!
0%
b111 *
0-
02
b111 6
#731350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#731360000000
0!
0%
b0 *
0-
02
b0 6
#731370000000
1!
1%
1-
12
#731380000000
0!
0%
b1 *
0-
02
b1 6
#731390000000
1!
1%
1-
12
#731400000000
0!
0%
b10 *
0-
02
b10 6
#731410000000
1!
1%
1-
12
#731420000000
0!
0%
b11 *
0-
02
b11 6
#731430000000
1!
1%
1-
12
15
#731440000000
0!
0%
b100 *
0-
02
b100 6
#731450000000
1!
1%
1-
12
#731460000000
0!
0%
b101 *
0-
02
b101 6
#731470000000
1!
1%
1-
12
#731480000000
0!
0%
b110 *
0-
02
b110 6
#731490000000
1!
1%
1-
12
#731500000000
0!
0%
b111 *
0-
02
b111 6
#731510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#731520000000
0!
0%
b0 *
0-
02
b0 6
#731530000000
1!
1%
1-
12
#731540000000
0!
0%
b1 *
0-
02
b1 6
#731550000000
1!
1%
1-
12
#731560000000
0!
0%
b10 *
0-
02
b10 6
#731570000000
1!
1%
1-
12
#731580000000
0!
0%
b11 *
0-
02
b11 6
#731590000000
1!
1%
1-
12
15
#731600000000
0!
0%
b100 *
0-
02
b100 6
#731610000000
1!
1%
1-
12
#731620000000
0!
0%
b101 *
0-
02
b101 6
#731630000000
1!
1%
1-
12
#731640000000
0!
0%
b110 *
0-
02
b110 6
#731650000000
1!
1%
1-
12
#731660000000
0!
0%
b111 *
0-
02
b111 6
#731670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#731680000000
0!
0%
b0 *
0-
02
b0 6
#731690000000
1!
1%
1-
12
#731700000000
0!
0%
b1 *
0-
02
b1 6
#731710000000
1!
1%
1-
12
#731720000000
0!
0%
b10 *
0-
02
b10 6
#731730000000
1!
1%
1-
12
#731740000000
0!
0%
b11 *
0-
02
b11 6
#731750000000
1!
1%
1-
12
15
#731760000000
0!
0%
b100 *
0-
02
b100 6
#731770000000
1!
1%
1-
12
#731780000000
0!
0%
b101 *
0-
02
b101 6
#731790000000
1!
1%
1-
12
#731800000000
0!
0%
b110 *
0-
02
b110 6
#731810000000
1!
1%
1-
12
#731820000000
0!
0%
b111 *
0-
02
b111 6
#731830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#731840000000
0!
0%
b0 *
0-
02
b0 6
#731850000000
1!
1%
1-
12
#731860000000
0!
0%
b1 *
0-
02
b1 6
#731870000000
1!
1%
1-
12
#731880000000
0!
0%
b10 *
0-
02
b10 6
#731890000000
1!
1%
1-
12
#731900000000
0!
0%
b11 *
0-
02
b11 6
#731910000000
1!
1%
1-
12
15
#731920000000
0!
0%
b100 *
0-
02
b100 6
#731930000000
1!
1%
1-
12
#731940000000
0!
0%
b101 *
0-
02
b101 6
#731950000000
1!
1%
1-
12
#731960000000
0!
0%
b110 *
0-
02
b110 6
#731970000000
1!
1%
1-
12
#731980000000
0!
0%
b111 *
0-
02
b111 6
#731990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#732000000000
0!
0%
b0 *
0-
02
b0 6
#732010000000
1!
1%
1-
12
#732020000000
0!
0%
b1 *
0-
02
b1 6
#732030000000
1!
1%
1-
12
#732040000000
0!
0%
b10 *
0-
02
b10 6
#732050000000
1!
1%
1-
12
#732060000000
0!
0%
b11 *
0-
02
b11 6
#732070000000
1!
1%
1-
12
15
#732080000000
0!
0%
b100 *
0-
02
b100 6
#732090000000
1!
1%
1-
12
#732100000000
0!
0%
b101 *
0-
02
b101 6
#732110000000
1!
1%
1-
12
#732120000000
0!
0%
b110 *
0-
02
b110 6
#732130000000
1!
1%
1-
12
#732140000000
0!
0%
b111 *
0-
02
b111 6
#732150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#732160000000
0!
0%
b0 *
0-
02
b0 6
#732170000000
1!
1%
1-
12
#732180000000
0!
0%
b1 *
0-
02
b1 6
#732190000000
1!
1%
1-
12
#732200000000
0!
0%
b10 *
0-
02
b10 6
#732210000000
1!
1%
1-
12
#732220000000
0!
0%
b11 *
0-
02
b11 6
#732230000000
1!
1%
1-
12
15
#732240000000
0!
0%
b100 *
0-
02
b100 6
#732250000000
1!
1%
1-
12
#732260000000
0!
0%
b101 *
0-
02
b101 6
#732270000000
1!
1%
1-
12
#732280000000
0!
0%
b110 *
0-
02
b110 6
#732290000000
1!
1%
1-
12
#732300000000
0!
0%
b111 *
0-
02
b111 6
#732310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#732320000000
0!
0%
b0 *
0-
02
b0 6
#732330000000
1!
1%
1-
12
#732340000000
0!
0%
b1 *
0-
02
b1 6
#732350000000
1!
1%
1-
12
#732360000000
0!
0%
b10 *
0-
02
b10 6
#732370000000
1!
1%
1-
12
#732380000000
0!
0%
b11 *
0-
02
b11 6
#732390000000
1!
1%
1-
12
15
#732400000000
0!
0%
b100 *
0-
02
b100 6
#732410000000
1!
1%
1-
12
#732420000000
0!
0%
b101 *
0-
02
b101 6
#732430000000
1!
1%
1-
12
#732440000000
0!
0%
b110 *
0-
02
b110 6
#732450000000
1!
1%
1-
12
#732460000000
0!
0%
b111 *
0-
02
b111 6
#732470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#732480000000
0!
0%
b0 *
0-
02
b0 6
#732490000000
1!
1%
1-
12
#732500000000
0!
0%
b1 *
0-
02
b1 6
#732510000000
1!
1%
1-
12
#732520000000
0!
0%
b10 *
0-
02
b10 6
#732530000000
1!
1%
1-
12
#732540000000
0!
0%
b11 *
0-
02
b11 6
#732550000000
1!
1%
1-
12
15
#732560000000
0!
0%
b100 *
0-
02
b100 6
#732570000000
1!
1%
1-
12
#732580000000
0!
0%
b101 *
0-
02
b101 6
#732590000000
1!
1%
1-
12
#732600000000
0!
0%
b110 *
0-
02
b110 6
#732610000000
1!
1%
1-
12
#732620000000
0!
0%
b111 *
0-
02
b111 6
#732630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#732640000000
0!
0%
b0 *
0-
02
b0 6
#732650000000
1!
1%
1-
12
#732660000000
0!
0%
b1 *
0-
02
b1 6
#732670000000
1!
1%
1-
12
#732680000000
0!
0%
b10 *
0-
02
b10 6
#732690000000
1!
1%
1-
12
#732700000000
0!
0%
b11 *
0-
02
b11 6
#732710000000
1!
1%
1-
12
15
#732720000000
0!
0%
b100 *
0-
02
b100 6
#732730000000
1!
1%
1-
12
#732740000000
0!
0%
b101 *
0-
02
b101 6
#732750000000
1!
1%
1-
12
#732760000000
0!
0%
b110 *
0-
02
b110 6
#732770000000
1!
1%
1-
12
#732780000000
0!
0%
b111 *
0-
02
b111 6
#732790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#732800000000
0!
0%
b0 *
0-
02
b0 6
#732810000000
1!
1%
1-
12
#732820000000
0!
0%
b1 *
0-
02
b1 6
#732830000000
1!
1%
1-
12
#732840000000
0!
0%
b10 *
0-
02
b10 6
#732850000000
1!
1%
1-
12
#732860000000
0!
0%
b11 *
0-
02
b11 6
#732870000000
1!
1%
1-
12
15
#732880000000
0!
0%
b100 *
0-
02
b100 6
#732890000000
1!
1%
1-
12
#732900000000
0!
0%
b101 *
0-
02
b101 6
#732910000000
1!
1%
1-
12
#732920000000
0!
0%
b110 *
0-
02
b110 6
#732930000000
1!
1%
1-
12
#732940000000
0!
0%
b111 *
0-
02
b111 6
#732950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#732960000000
0!
0%
b0 *
0-
02
b0 6
#732970000000
1!
1%
1-
12
#732980000000
0!
0%
b1 *
0-
02
b1 6
#732990000000
1!
1%
1-
12
#733000000000
0!
0%
b10 *
0-
02
b10 6
#733010000000
1!
1%
1-
12
#733020000000
0!
0%
b11 *
0-
02
b11 6
#733030000000
1!
1%
1-
12
15
#733040000000
0!
0%
b100 *
0-
02
b100 6
#733050000000
1!
1%
1-
12
#733060000000
0!
0%
b101 *
0-
02
b101 6
#733070000000
1!
1%
1-
12
#733080000000
0!
0%
b110 *
0-
02
b110 6
#733090000000
1!
1%
1-
12
#733100000000
0!
0%
b111 *
0-
02
b111 6
#733110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#733120000000
0!
0%
b0 *
0-
02
b0 6
#733130000000
1!
1%
1-
12
#733140000000
0!
0%
b1 *
0-
02
b1 6
#733150000000
1!
1%
1-
12
#733160000000
0!
0%
b10 *
0-
02
b10 6
#733170000000
1!
1%
1-
12
#733180000000
0!
0%
b11 *
0-
02
b11 6
#733190000000
1!
1%
1-
12
15
#733200000000
0!
0%
b100 *
0-
02
b100 6
#733210000000
1!
1%
1-
12
#733220000000
0!
0%
b101 *
0-
02
b101 6
#733230000000
1!
1%
1-
12
#733240000000
0!
0%
b110 *
0-
02
b110 6
#733250000000
1!
1%
1-
12
#733260000000
0!
0%
b111 *
0-
02
b111 6
#733270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#733280000000
0!
0%
b0 *
0-
02
b0 6
#733290000000
1!
1%
1-
12
#733300000000
0!
0%
b1 *
0-
02
b1 6
#733310000000
1!
1%
1-
12
#733320000000
0!
0%
b10 *
0-
02
b10 6
#733330000000
1!
1%
1-
12
#733340000000
0!
0%
b11 *
0-
02
b11 6
#733350000000
1!
1%
1-
12
15
#733360000000
0!
0%
b100 *
0-
02
b100 6
#733370000000
1!
1%
1-
12
#733380000000
0!
0%
b101 *
0-
02
b101 6
#733390000000
1!
1%
1-
12
#733400000000
0!
0%
b110 *
0-
02
b110 6
#733410000000
1!
1%
1-
12
#733420000000
0!
0%
b111 *
0-
02
b111 6
#733430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#733440000000
0!
0%
b0 *
0-
02
b0 6
#733450000000
1!
1%
1-
12
#733460000000
0!
0%
b1 *
0-
02
b1 6
#733470000000
1!
1%
1-
12
#733480000000
0!
0%
b10 *
0-
02
b10 6
#733490000000
1!
1%
1-
12
#733500000000
0!
0%
b11 *
0-
02
b11 6
#733510000000
1!
1%
1-
12
15
#733520000000
0!
0%
b100 *
0-
02
b100 6
#733530000000
1!
1%
1-
12
#733540000000
0!
0%
b101 *
0-
02
b101 6
#733550000000
1!
1%
1-
12
#733560000000
0!
0%
b110 *
0-
02
b110 6
#733570000000
1!
1%
1-
12
#733580000000
0!
0%
b111 *
0-
02
b111 6
#733590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#733600000000
0!
0%
b0 *
0-
02
b0 6
#733610000000
1!
1%
1-
12
#733620000000
0!
0%
b1 *
0-
02
b1 6
#733630000000
1!
1%
1-
12
#733640000000
0!
0%
b10 *
0-
02
b10 6
#733650000000
1!
1%
1-
12
#733660000000
0!
0%
b11 *
0-
02
b11 6
#733670000000
1!
1%
1-
12
15
#733680000000
0!
0%
b100 *
0-
02
b100 6
#733690000000
1!
1%
1-
12
#733700000000
0!
0%
b101 *
0-
02
b101 6
#733710000000
1!
1%
1-
12
#733720000000
0!
0%
b110 *
0-
02
b110 6
#733730000000
1!
1%
1-
12
#733740000000
0!
0%
b111 *
0-
02
b111 6
#733750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#733760000000
0!
0%
b0 *
0-
02
b0 6
#733770000000
1!
1%
1-
12
#733780000000
0!
0%
b1 *
0-
02
b1 6
#733790000000
1!
1%
1-
12
#733800000000
0!
0%
b10 *
0-
02
b10 6
#733810000000
1!
1%
1-
12
#733820000000
0!
0%
b11 *
0-
02
b11 6
#733830000000
1!
1%
1-
12
15
#733840000000
0!
0%
b100 *
0-
02
b100 6
#733850000000
1!
1%
1-
12
#733860000000
0!
0%
b101 *
0-
02
b101 6
#733870000000
1!
1%
1-
12
#733880000000
0!
0%
b110 *
0-
02
b110 6
#733890000000
1!
1%
1-
12
#733900000000
0!
0%
b111 *
0-
02
b111 6
#733910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#733920000000
0!
0%
b0 *
0-
02
b0 6
#733930000000
1!
1%
1-
12
#733940000000
0!
0%
b1 *
0-
02
b1 6
#733950000000
1!
1%
1-
12
#733960000000
0!
0%
b10 *
0-
02
b10 6
#733970000000
1!
1%
1-
12
#733980000000
0!
0%
b11 *
0-
02
b11 6
#733990000000
1!
1%
1-
12
15
#734000000000
0!
0%
b100 *
0-
02
b100 6
#734010000000
1!
1%
1-
12
#734020000000
0!
0%
b101 *
0-
02
b101 6
#734030000000
1!
1%
1-
12
#734040000000
0!
0%
b110 *
0-
02
b110 6
#734050000000
1!
1%
1-
12
#734060000000
0!
0%
b111 *
0-
02
b111 6
#734070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#734080000000
0!
0%
b0 *
0-
02
b0 6
#734090000000
1!
1%
1-
12
#734100000000
0!
0%
b1 *
0-
02
b1 6
#734110000000
1!
1%
1-
12
#734120000000
0!
0%
b10 *
0-
02
b10 6
#734130000000
1!
1%
1-
12
#734140000000
0!
0%
b11 *
0-
02
b11 6
#734150000000
1!
1%
1-
12
15
#734160000000
0!
0%
b100 *
0-
02
b100 6
#734170000000
1!
1%
1-
12
#734180000000
0!
0%
b101 *
0-
02
b101 6
#734190000000
1!
1%
1-
12
#734200000000
0!
0%
b110 *
0-
02
b110 6
#734210000000
1!
1%
1-
12
#734220000000
0!
0%
b111 *
0-
02
b111 6
#734230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#734240000000
0!
0%
b0 *
0-
02
b0 6
#734250000000
1!
1%
1-
12
#734260000000
0!
0%
b1 *
0-
02
b1 6
#734270000000
1!
1%
1-
12
#734280000000
0!
0%
b10 *
0-
02
b10 6
#734290000000
1!
1%
1-
12
#734300000000
0!
0%
b11 *
0-
02
b11 6
#734310000000
1!
1%
1-
12
15
#734320000000
0!
0%
b100 *
0-
02
b100 6
#734330000000
1!
1%
1-
12
#734340000000
0!
0%
b101 *
0-
02
b101 6
#734350000000
1!
1%
1-
12
#734360000000
0!
0%
b110 *
0-
02
b110 6
#734370000000
1!
1%
1-
12
#734380000000
0!
0%
b111 *
0-
02
b111 6
#734390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#734400000000
0!
0%
b0 *
0-
02
b0 6
#734410000000
1!
1%
1-
12
#734420000000
0!
0%
b1 *
0-
02
b1 6
#734430000000
1!
1%
1-
12
#734440000000
0!
0%
b10 *
0-
02
b10 6
#734450000000
1!
1%
1-
12
#734460000000
0!
0%
b11 *
0-
02
b11 6
#734470000000
1!
1%
1-
12
15
#734480000000
0!
0%
b100 *
0-
02
b100 6
#734490000000
1!
1%
1-
12
#734500000000
0!
0%
b101 *
0-
02
b101 6
#734510000000
1!
1%
1-
12
#734520000000
0!
0%
b110 *
0-
02
b110 6
#734530000000
1!
1%
1-
12
#734540000000
0!
0%
b111 *
0-
02
b111 6
#734550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#734560000000
0!
0%
b0 *
0-
02
b0 6
#734570000000
1!
1%
1-
12
#734580000000
0!
0%
b1 *
0-
02
b1 6
#734590000000
1!
1%
1-
12
#734600000000
0!
0%
b10 *
0-
02
b10 6
#734610000000
1!
1%
1-
12
#734620000000
0!
0%
b11 *
0-
02
b11 6
#734630000000
1!
1%
1-
12
15
#734640000000
0!
0%
b100 *
0-
02
b100 6
#734650000000
1!
1%
1-
12
#734660000000
0!
0%
b101 *
0-
02
b101 6
#734670000000
1!
1%
1-
12
#734680000000
0!
0%
b110 *
0-
02
b110 6
#734690000000
1!
1%
1-
12
#734700000000
0!
0%
b111 *
0-
02
b111 6
#734710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#734720000000
0!
0%
b0 *
0-
02
b0 6
#734730000000
1!
1%
1-
12
#734740000000
0!
0%
b1 *
0-
02
b1 6
#734750000000
1!
1%
1-
12
#734760000000
0!
0%
b10 *
0-
02
b10 6
#734770000000
1!
1%
1-
12
#734780000000
0!
0%
b11 *
0-
02
b11 6
#734790000000
1!
1%
1-
12
15
#734800000000
0!
0%
b100 *
0-
02
b100 6
#734810000000
1!
1%
1-
12
#734820000000
0!
0%
b101 *
0-
02
b101 6
#734830000000
1!
1%
1-
12
#734840000000
0!
0%
b110 *
0-
02
b110 6
#734850000000
1!
1%
1-
12
#734860000000
0!
0%
b111 *
0-
02
b111 6
#734870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#734880000000
0!
0%
b0 *
0-
02
b0 6
#734890000000
1!
1%
1-
12
#734900000000
0!
0%
b1 *
0-
02
b1 6
#734910000000
1!
1%
1-
12
#734920000000
0!
0%
b10 *
0-
02
b10 6
#734930000000
1!
1%
1-
12
#734940000000
0!
0%
b11 *
0-
02
b11 6
#734950000000
1!
1%
1-
12
15
#734960000000
0!
0%
b100 *
0-
02
b100 6
#734970000000
1!
1%
1-
12
#734980000000
0!
0%
b101 *
0-
02
b101 6
#734990000000
1!
1%
1-
12
#735000000000
0!
0%
b110 *
0-
02
b110 6
#735010000000
1!
1%
1-
12
#735020000000
0!
0%
b111 *
0-
02
b111 6
#735030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#735040000000
0!
0%
b0 *
0-
02
b0 6
#735050000000
1!
1%
1-
12
#735060000000
0!
0%
b1 *
0-
02
b1 6
#735070000000
1!
1%
1-
12
#735080000000
0!
0%
b10 *
0-
02
b10 6
#735090000000
1!
1%
1-
12
#735100000000
0!
0%
b11 *
0-
02
b11 6
#735110000000
1!
1%
1-
12
15
#735120000000
0!
0%
b100 *
0-
02
b100 6
#735130000000
1!
1%
1-
12
#735140000000
0!
0%
b101 *
0-
02
b101 6
#735150000000
1!
1%
1-
12
#735160000000
0!
0%
b110 *
0-
02
b110 6
#735170000000
1!
1%
1-
12
#735180000000
0!
0%
b111 *
0-
02
b111 6
#735190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#735200000000
0!
0%
b0 *
0-
02
b0 6
#735210000000
1!
1%
1-
12
#735220000000
0!
0%
b1 *
0-
02
b1 6
#735230000000
1!
1%
1-
12
#735240000000
0!
0%
b10 *
0-
02
b10 6
#735250000000
1!
1%
1-
12
#735260000000
0!
0%
b11 *
0-
02
b11 6
#735270000000
1!
1%
1-
12
15
#735280000000
0!
0%
b100 *
0-
02
b100 6
#735290000000
1!
1%
1-
12
#735300000000
0!
0%
b101 *
0-
02
b101 6
#735310000000
1!
1%
1-
12
#735320000000
0!
0%
b110 *
0-
02
b110 6
#735330000000
1!
1%
1-
12
#735340000000
0!
0%
b111 *
0-
02
b111 6
#735350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#735360000000
0!
0%
b0 *
0-
02
b0 6
#735370000000
1!
1%
1-
12
#735380000000
0!
0%
b1 *
0-
02
b1 6
#735390000000
1!
1%
1-
12
#735400000000
0!
0%
b10 *
0-
02
b10 6
#735410000000
1!
1%
1-
12
#735420000000
0!
0%
b11 *
0-
02
b11 6
#735430000000
1!
1%
1-
12
15
#735440000000
0!
0%
b100 *
0-
02
b100 6
#735450000000
1!
1%
1-
12
#735460000000
0!
0%
b101 *
0-
02
b101 6
#735470000000
1!
1%
1-
12
#735480000000
0!
0%
b110 *
0-
02
b110 6
#735490000000
1!
1%
1-
12
#735500000000
0!
0%
b111 *
0-
02
b111 6
#735510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#735520000000
0!
0%
b0 *
0-
02
b0 6
#735530000000
1!
1%
1-
12
#735540000000
0!
0%
b1 *
0-
02
b1 6
#735550000000
1!
1%
1-
12
#735560000000
0!
0%
b10 *
0-
02
b10 6
#735570000000
1!
1%
1-
12
#735580000000
0!
0%
b11 *
0-
02
b11 6
#735590000000
1!
1%
1-
12
15
#735600000000
0!
0%
b100 *
0-
02
b100 6
#735610000000
1!
1%
1-
12
#735620000000
0!
0%
b101 *
0-
02
b101 6
#735630000000
1!
1%
1-
12
#735640000000
0!
0%
b110 *
0-
02
b110 6
#735650000000
1!
1%
1-
12
#735660000000
0!
0%
b111 *
0-
02
b111 6
#735670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#735680000000
0!
0%
b0 *
0-
02
b0 6
#735690000000
1!
1%
1-
12
#735700000000
0!
0%
b1 *
0-
02
b1 6
#735710000000
1!
1%
1-
12
#735720000000
0!
0%
b10 *
0-
02
b10 6
#735730000000
1!
1%
1-
12
#735740000000
0!
0%
b11 *
0-
02
b11 6
#735750000000
1!
1%
1-
12
15
#735760000000
0!
0%
b100 *
0-
02
b100 6
#735770000000
1!
1%
1-
12
#735780000000
0!
0%
b101 *
0-
02
b101 6
#735790000000
1!
1%
1-
12
#735800000000
0!
0%
b110 *
0-
02
b110 6
#735810000000
1!
1%
1-
12
#735820000000
0!
0%
b111 *
0-
02
b111 6
#735830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#735840000000
0!
0%
b0 *
0-
02
b0 6
#735850000000
1!
1%
1-
12
#735860000000
0!
0%
b1 *
0-
02
b1 6
#735870000000
1!
1%
1-
12
#735880000000
0!
0%
b10 *
0-
02
b10 6
#735890000000
1!
1%
1-
12
#735900000000
0!
0%
b11 *
0-
02
b11 6
#735910000000
1!
1%
1-
12
15
#735920000000
0!
0%
b100 *
0-
02
b100 6
#735930000000
1!
1%
1-
12
#735940000000
0!
0%
b101 *
0-
02
b101 6
#735950000000
1!
1%
1-
12
#735960000000
0!
0%
b110 *
0-
02
b110 6
#735970000000
1!
1%
1-
12
#735980000000
0!
0%
b111 *
0-
02
b111 6
#735990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#736000000000
0!
0%
b0 *
0-
02
b0 6
#736010000000
1!
1%
1-
12
#736020000000
0!
0%
b1 *
0-
02
b1 6
#736030000000
1!
1%
1-
12
#736040000000
0!
0%
b10 *
0-
02
b10 6
#736050000000
1!
1%
1-
12
#736060000000
0!
0%
b11 *
0-
02
b11 6
#736070000000
1!
1%
1-
12
15
#736080000000
0!
0%
b100 *
0-
02
b100 6
#736090000000
1!
1%
1-
12
#736100000000
0!
0%
b101 *
0-
02
b101 6
#736110000000
1!
1%
1-
12
#736120000000
0!
0%
b110 *
0-
02
b110 6
#736130000000
1!
1%
1-
12
#736140000000
0!
0%
b111 *
0-
02
b111 6
#736150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#736160000000
0!
0%
b0 *
0-
02
b0 6
#736170000000
1!
1%
1-
12
#736180000000
0!
0%
b1 *
0-
02
b1 6
#736190000000
1!
1%
1-
12
#736200000000
0!
0%
b10 *
0-
02
b10 6
#736210000000
1!
1%
1-
12
#736220000000
0!
0%
b11 *
0-
02
b11 6
#736230000000
1!
1%
1-
12
15
#736240000000
0!
0%
b100 *
0-
02
b100 6
#736250000000
1!
1%
1-
12
#736260000000
0!
0%
b101 *
0-
02
b101 6
#736270000000
1!
1%
1-
12
#736280000000
0!
0%
b110 *
0-
02
b110 6
#736290000000
1!
1%
1-
12
#736300000000
0!
0%
b111 *
0-
02
b111 6
#736310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#736320000000
0!
0%
b0 *
0-
02
b0 6
#736330000000
1!
1%
1-
12
#736340000000
0!
0%
b1 *
0-
02
b1 6
#736350000000
1!
1%
1-
12
#736360000000
0!
0%
b10 *
0-
02
b10 6
#736370000000
1!
1%
1-
12
#736380000000
0!
0%
b11 *
0-
02
b11 6
#736390000000
1!
1%
1-
12
15
#736400000000
0!
0%
b100 *
0-
02
b100 6
#736410000000
1!
1%
1-
12
#736420000000
0!
0%
b101 *
0-
02
b101 6
#736430000000
1!
1%
1-
12
#736440000000
0!
0%
b110 *
0-
02
b110 6
#736450000000
1!
1%
1-
12
#736460000000
0!
0%
b111 *
0-
02
b111 6
#736470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#736480000000
0!
0%
b0 *
0-
02
b0 6
#736490000000
1!
1%
1-
12
#736500000000
0!
0%
b1 *
0-
02
b1 6
#736510000000
1!
1%
1-
12
#736520000000
0!
0%
b10 *
0-
02
b10 6
#736530000000
1!
1%
1-
12
#736540000000
0!
0%
b11 *
0-
02
b11 6
#736550000000
1!
1%
1-
12
15
#736560000000
0!
0%
b100 *
0-
02
b100 6
#736570000000
1!
1%
1-
12
#736580000000
0!
0%
b101 *
0-
02
b101 6
#736590000000
1!
1%
1-
12
#736600000000
0!
0%
b110 *
0-
02
b110 6
#736610000000
1!
1%
1-
12
#736620000000
0!
0%
b111 *
0-
02
b111 6
#736630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#736640000000
0!
0%
b0 *
0-
02
b0 6
#736650000000
1!
1%
1-
12
#736660000000
0!
0%
b1 *
0-
02
b1 6
#736670000000
1!
1%
1-
12
#736680000000
0!
0%
b10 *
0-
02
b10 6
#736690000000
1!
1%
1-
12
#736700000000
0!
0%
b11 *
0-
02
b11 6
#736710000000
1!
1%
1-
12
15
#736720000000
0!
0%
b100 *
0-
02
b100 6
#736730000000
1!
1%
1-
12
#736740000000
0!
0%
b101 *
0-
02
b101 6
#736750000000
1!
1%
1-
12
#736760000000
0!
0%
b110 *
0-
02
b110 6
#736770000000
1!
1%
1-
12
#736780000000
0!
0%
b111 *
0-
02
b111 6
#736790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#736800000000
0!
0%
b0 *
0-
02
b0 6
#736810000000
1!
1%
1-
12
#736820000000
0!
0%
b1 *
0-
02
b1 6
#736830000000
1!
1%
1-
12
#736840000000
0!
0%
b10 *
0-
02
b10 6
#736850000000
1!
1%
1-
12
#736860000000
0!
0%
b11 *
0-
02
b11 6
#736870000000
1!
1%
1-
12
15
#736880000000
0!
0%
b100 *
0-
02
b100 6
#736890000000
1!
1%
1-
12
#736900000000
0!
0%
b101 *
0-
02
b101 6
#736910000000
1!
1%
1-
12
#736920000000
0!
0%
b110 *
0-
02
b110 6
#736930000000
1!
1%
1-
12
#736940000000
0!
0%
b111 *
0-
02
b111 6
#736950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#736960000000
0!
0%
b0 *
0-
02
b0 6
#736970000000
1!
1%
1-
12
#736980000000
0!
0%
b1 *
0-
02
b1 6
#736990000000
1!
1%
1-
12
#737000000000
0!
0%
b10 *
0-
02
b10 6
#737010000000
1!
1%
1-
12
#737020000000
0!
0%
b11 *
0-
02
b11 6
#737030000000
1!
1%
1-
12
15
#737040000000
0!
0%
b100 *
0-
02
b100 6
#737050000000
1!
1%
1-
12
#737060000000
0!
0%
b101 *
0-
02
b101 6
#737070000000
1!
1%
1-
12
#737080000000
0!
0%
b110 *
0-
02
b110 6
#737090000000
1!
1%
1-
12
#737100000000
0!
0%
b111 *
0-
02
b111 6
#737110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#737120000000
0!
0%
b0 *
0-
02
b0 6
#737130000000
1!
1%
1-
12
#737140000000
0!
0%
b1 *
0-
02
b1 6
#737150000000
1!
1%
1-
12
#737160000000
0!
0%
b10 *
0-
02
b10 6
#737170000000
1!
1%
1-
12
#737180000000
0!
0%
b11 *
0-
02
b11 6
#737190000000
1!
1%
1-
12
15
#737200000000
0!
0%
b100 *
0-
02
b100 6
#737210000000
1!
1%
1-
12
#737220000000
0!
0%
b101 *
0-
02
b101 6
#737230000000
1!
1%
1-
12
#737240000000
0!
0%
b110 *
0-
02
b110 6
#737250000000
1!
1%
1-
12
#737260000000
0!
0%
b111 *
0-
02
b111 6
#737270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#737280000000
0!
0%
b0 *
0-
02
b0 6
#737290000000
1!
1%
1-
12
#737300000000
0!
0%
b1 *
0-
02
b1 6
#737310000000
1!
1%
1-
12
#737320000000
0!
0%
b10 *
0-
02
b10 6
#737330000000
1!
1%
1-
12
#737340000000
0!
0%
b11 *
0-
02
b11 6
#737350000000
1!
1%
1-
12
15
#737360000000
0!
0%
b100 *
0-
02
b100 6
#737370000000
1!
1%
1-
12
#737380000000
0!
0%
b101 *
0-
02
b101 6
#737390000000
1!
1%
1-
12
#737400000000
0!
0%
b110 *
0-
02
b110 6
#737410000000
1!
1%
1-
12
#737420000000
0!
0%
b111 *
0-
02
b111 6
#737430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#737440000000
0!
0%
b0 *
0-
02
b0 6
#737450000000
1!
1%
1-
12
#737460000000
0!
0%
b1 *
0-
02
b1 6
#737470000000
1!
1%
1-
12
#737480000000
0!
0%
b10 *
0-
02
b10 6
#737490000000
1!
1%
1-
12
#737500000000
0!
0%
b11 *
0-
02
b11 6
#737510000000
1!
1%
1-
12
15
#737520000000
0!
0%
b100 *
0-
02
b100 6
#737530000000
1!
1%
1-
12
#737540000000
0!
0%
b101 *
0-
02
b101 6
#737550000000
1!
1%
1-
12
#737560000000
0!
0%
b110 *
0-
02
b110 6
#737570000000
1!
1%
1-
12
#737580000000
0!
0%
b111 *
0-
02
b111 6
#737590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#737600000000
0!
0%
b0 *
0-
02
b0 6
#737610000000
1!
1%
1-
12
#737620000000
0!
0%
b1 *
0-
02
b1 6
#737630000000
1!
1%
1-
12
#737640000000
0!
0%
b10 *
0-
02
b10 6
#737650000000
1!
1%
1-
12
#737660000000
0!
0%
b11 *
0-
02
b11 6
#737670000000
1!
1%
1-
12
15
#737680000000
0!
0%
b100 *
0-
02
b100 6
#737690000000
1!
1%
1-
12
#737700000000
0!
0%
b101 *
0-
02
b101 6
#737710000000
1!
1%
1-
12
#737720000000
0!
0%
b110 *
0-
02
b110 6
#737730000000
1!
1%
1-
12
#737740000000
0!
0%
b111 *
0-
02
b111 6
#737750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#737760000000
0!
0%
b0 *
0-
02
b0 6
#737770000000
1!
1%
1-
12
#737780000000
0!
0%
b1 *
0-
02
b1 6
#737790000000
1!
1%
1-
12
#737800000000
0!
0%
b10 *
0-
02
b10 6
#737810000000
1!
1%
1-
12
#737820000000
0!
0%
b11 *
0-
02
b11 6
#737830000000
1!
1%
1-
12
15
#737840000000
0!
0%
b100 *
0-
02
b100 6
#737850000000
1!
1%
1-
12
#737860000000
0!
0%
b101 *
0-
02
b101 6
#737870000000
1!
1%
1-
12
#737880000000
0!
0%
b110 *
0-
02
b110 6
#737890000000
1!
1%
1-
12
#737900000000
0!
0%
b111 *
0-
02
b111 6
#737910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#737920000000
0!
0%
b0 *
0-
02
b0 6
#737930000000
1!
1%
1-
12
#737940000000
0!
0%
b1 *
0-
02
b1 6
#737950000000
1!
1%
1-
12
#737960000000
0!
0%
b10 *
0-
02
b10 6
#737970000000
1!
1%
1-
12
#737980000000
0!
0%
b11 *
0-
02
b11 6
#737990000000
1!
1%
1-
12
15
#738000000000
0!
0%
b100 *
0-
02
b100 6
#738010000000
1!
1%
1-
12
#738020000000
0!
0%
b101 *
0-
02
b101 6
#738030000000
1!
1%
1-
12
#738040000000
0!
0%
b110 *
0-
02
b110 6
#738050000000
1!
1%
1-
12
#738060000000
0!
0%
b111 *
0-
02
b111 6
#738070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#738080000000
0!
0%
b0 *
0-
02
b0 6
#738090000000
1!
1%
1-
12
#738100000000
0!
0%
b1 *
0-
02
b1 6
#738110000000
1!
1%
1-
12
#738120000000
0!
0%
b10 *
0-
02
b10 6
#738130000000
1!
1%
1-
12
#738140000000
0!
0%
b11 *
0-
02
b11 6
#738150000000
1!
1%
1-
12
15
#738160000000
0!
0%
b100 *
0-
02
b100 6
#738170000000
1!
1%
1-
12
#738180000000
0!
0%
b101 *
0-
02
b101 6
#738190000000
1!
1%
1-
12
#738200000000
0!
0%
b110 *
0-
02
b110 6
#738210000000
1!
1%
1-
12
#738220000000
0!
0%
b111 *
0-
02
b111 6
#738230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#738240000000
0!
0%
b0 *
0-
02
b0 6
#738250000000
1!
1%
1-
12
#738260000000
0!
0%
b1 *
0-
02
b1 6
#738270000000
1!
1%
1-
12
#738280000000
0!
0%
b10 *
0-
02
b10 6
#738290000000
1!
1%
1-
12
#738300000000
0!
0%
b11 *
0-
02
b11 6
#738310000000
1!
1%
1-
12
15
#738320000000
0!
0%
b100 *
0-
02
b100 6
#738330000000
1!
1%
1-
12
#738340000000
0!
0%
b101 *
0-
02
b101 6
#738350000000
1!
1%
1-
12
#738360000000
0!
0%
b110 *
0-
02
b110 6
#738370000000
1!
1%
1-
12
#738380000000
0!
0%
b111 *
0-
02
b111 6
#738390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#738400000000
0!
0%
b0 *
0-
02
b0 6
#738410000000
1!
1%
1-
12
#738420000000
0!
0%
b1 *
0-
02
b1 6
#738430000000
1!
1%
1-
12
#738440000000
0!
0%
b10 *
0-
02
b10 6
#738450000000
1!
1%
1-
12
#738460000000
0!
0%
b11 *
0-
02
b11 6
#738470000000
1!
1%
1-
12
15
#738480000000
0!
0%
b100 *
0-
02
b100 6
#738490000000
1!
1%
1-
12
#738500000000
0!
0%
b101 *
0-
02
b101 6
#738510000000
1!
1%
1-
12
#738520000000
0!
0%
b110 *
0-
02
b110 6
#738530000000
1!
1%
1-
12
#738540000000
0!
0%
b111 *
0-
02
b111 6
#738550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#738560000000
0!
0%
b0 *
0-
02
b0 6
#738570000000
1!
1%
1-
12
#738580000000
0!
0%
b1 *
0-
02
b1 6
#738590000000
1!
1%
1-
12
#738600000000
0!
0%
b10 *
0-
02
b10 6
#738610000000
1!
1%
1-
12
#738620000000
0!
0%
b11 *
0-
02
b11 6
#738630000000
1!
1%
1-
12
15
#738640000000
0!
0%
b100 *
0-
02
b100 6
#738650000000
1!
1%
1-
12
#738660000000
0!
0%
b101 *
0-
02
b101 6
#738670000000
1!
1%
1-
12
#738680000000
0!
0%
b110 *
0-
02
b110 6
#738690000000
1!
1%
1-
12
#738700000000
0!
0%
b111 *
0-
02
b111 6
#738710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#738720000000
0!
0%
b0 *
0-
02
b0 6
#738730000000
1!
1%
1-
12
#738740000000
0!
0%
b1 *
0-
02
b1 6
#738750000000
1!
1%
1-
12
#738760000000
0!
0%
b10 *
0-
02
b10 6
#738770000000
1!
1%
1-
12
#738780000000
0!
0%
b11 *
0-
02
b11 6
#738790000000
1!
1%
1-
12
15
#738800000000
0!
0%
b100 *
0-
02
b100 6
#738810000000
1!
1%
1-
12
#738820000000
0!
0%
b101 *
0-
02
b101 6
#738830000000
1!
1%
1-
12
#738840000000
0!
0%
b110 *
0-
02
b110 6
#738850000000
1!
1%
1-
12
#738860000000
0!
0%
b111 *
0-
02
b111 6
#738870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#738880000000
0!
0%
b0 *
0-
02
b0 6
#738890000000
1!
1%
1-
12
#738900000000
0!
0%
b1 *
0-
02
b1 6
#738910000000
1!
1%
1-
12
#738920000000
0!
0%
b10 *
0-
02
b10 6
#738930000000
1!
1%
1-
12
#738940000000
0!
0%
b11 *
0-
02
b11 6
#738950000000
1!
1%
1-
12
15
#738960000000
0!
0%
b100 *
0-
02
b100 6
#738970000000
1!
1%
1-
12
#738980000000
0!
0%
b101 *
0-
02
b101 6
#738990000000
1!
1%
1-
12
#739000000000
0!
0%
b110 *
0-
02
b110 6
#739010000000
1!
1%
1-
12
#739020000000
0!
0%
b111 *
0-
02
b111 6
#739030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#739040000000
0!
0%
b0 *
0-
02
b0 6
#739050000000
1!
1%
1-
12
#739060000000
0!
0%
b1 *
0-
02
b1 6
#739070000000
1!
1%
1-
12
#739080000000
0!
0%
b10 *
0-
02
b10 6
#739090000000
1!
1%
1-
12
#739100000000
0!
0%
b11 *
0-
02
b11 6
#739110000000
1!
1%
1-
12
15
#739120000000
0!
0%
b100 *
0-
02
b100 6
#739130000000
1!
1%
1-
12
#739140000000
0!
0%
b101 *
0-
02
b101 6
#739150000000
1!
1%
1-
12
#739160000000
0!
0%
b110 *
0-
02
b110 6
#739170000000
1!
1%
1-
12
#739180000000
0!
0%
b111 *
0-
02
b111 6
#739190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#739200000000
0!
0%
b0 *
0-
02
b0 6
#739210000000
1!
1%
1-
12
#739220000000
0!
0%
b1 *
0-
02
b1 6
#739230000000
1!
1%
1-
12
#739240000000
0!
0%
b10 *
0-
02
b10 6
#739250000000
1!
1%
1-
12
#739260000000
0!
0%
b11 *
0-
02
b11 6
#739270000000
1!
1%
1-
12
15
#739280000000
0!
0%
b100 *
0-
02
b100 6
#739290000000
1!
1%
1-
12
#739300000000
0!
0%
b101 *
0-
02
b101 6
#739310000000
1!
1%
1-
12
#739320000000
0!
0%
b110 *
0-
02
b110 6
#739330000000
1!
1%
1-
12
#739340000000
0!
0%
b111 *
0-
02
b111 6
#739350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#739360000000
0!
0%
b0 *
0-
02
b0 6
#739370000000
1!
1%
1-
12
#739380000000
0!
0%
b1 *
0-
02
b1 6
#739390000000
1!
1%
1-
12
#739400000000
0!
0%
b10 *
0-
02
b10 6
#739410000000
1!
1%
1-
12
#739420000000
0!
0%
b11 *
0-
02
b11 6
#739430000000
1!
1%
1-
12
15
#739440000000
0!
0%
b100 *
0-
02
b100 6
#739450000000
1!
1%
1-
12
#739460000000
0!
0%
b101 *
0-
02
b101 6
#739470000000
1!
1%
1-
12
#739480000000
0!
0%
b110 *
0-
02
b110 6
#739490000000
1!
1%
1-
12
#739500000000
0!
0%
b111 *
0-
02
b111 6
#739510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#739520000000
0!
0%
b0 *
0-
02
b0 6
#739530000000
1!
1%
1-
12
#739540000000
0!
0%
b1 *
0-
02
b1 6
#739550000000
1!
1%
1-
12
#739560000000
0!
0%
b10 *
0-
02
b10 6
#739570000000
1!
1%
1-
12
#739580000000
0!
0%
b11 *
0-
02
b11 6
#739590000000
1!
1%
1-
12
15
#739600000000
0!
0%
b100 *
0-
02
b100 6
#739610000000
1!
1%
1-
12
#739620000000
0!
0%
b101 *
0-
02
b101 6
#739630000000
1!
1%
1-
12
#739640000000
0!
0%
b110 *
0-
02
b110 6
#739650000000
1!
1%
1-
12
#739660000000
0!
0%
b111 *
0-
02
b111 6
#739670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#739680000000
0!
0%
b0 *
0-
02
b0 6
#739690000000
1!
1%
1-
12
#739700000000
0!
0%
b1 *
0-
02
b1 6
#739710000000
1!
1%
1-
12
#739720000000
0!
0%
b10 *
0-
02
b10 6
#739730000000
1!
1%
1-
12
#739740000000
0!
0%
b11 *
0-
02
b11 6
#739750000000
1!
1%
1-
12
15
#739760000000
0!
0%
b100 *
0-
02
b100 6
#739770000000
1!
1%
1-
12
#739780000000
0!
0%
b101 *
0-
02
b101 6
#739790000000
1!
1%
1-
12
#739800000000
0!
0%
b110 *
0-
02
b110 6
#739810000000
1!
1%
1-
12
#739820000000
0!
0%
b111 *
0-
02
b111 6
#739830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#739840000000
0!
0%
b0 *
0-
02
b0 6
#739850000000
1!
1%
1-
12
#739860000000
0!
0%
b1 *
0-
02
b1 6
#739870000000
1!
1%
1-
12
#739880000000
0!
0%
b10 *
0-
02
b10 6
#739890000000
1!
1%
1-
12
#739900000000
0!
0%
b11 *
0-
02
b11 6
#739910000000
1!
1%
1-
12
15
#739920000000
0!
0%
b100 *
0-
02
b100 6
#739930000000
1!
1%
1-
12
#739940000000
0!
0%
b101 *
0-
02
b101 6
#739950000000
1!
1%
1-
12
#739960000000
0!
0%
b110 *
0-
02
b110 6
#739970000000
1!
1%
1-
12
#739980000000
0!
0%
b111 *
0-
02
b111 6
#739990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#740000000000
0!
0%
b0 *
0-
02
b0 6
#740010000000
1!
1%
1-
12
#740020000000
0!
0%
b1 *
0-
02
b1 6
#740030000000
1!
1%
1-
12
#740040000000
0!
0%
b10 *
0-
02
b10 6
#740050000000
1!
1%
1-
12
#740060000000
0!
0%
b11 *
0-
02
b11 6
#740070000000
1!
1%
1-
12
15
#740080000000
0!
0%
b100 *
0-
02
b100 6
#740090000000
1!
1%
1-
12
#740100000000
0!
0%
b101 *
0-
02
b101 6
#740110000000
1!
1%
1-
12
#740120000000
0!
0%
b110 *
0-
02
b110 6
#740130000000
1!
1%
1-
12
#740140000000
0!
0%
b111 *
0-
02
b111 6
#740150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#740160000000
0!
0%
b0 *
0-
02
b0 6
#740170000000
1!
1%
1-
12
#740180000000
0!
0%
b1 *
0-
02
b1 6
#740190000000
1!
1%
1-
12
#740200000000
0!
0%
b10 *
0-
02
b10 6
#740210000000
1!
1%
1-
12
#740220000000
0!
0%
b11 *
0-
02
b11 6
#740230000000
1!
1%
1-
12
15
#740240000000
0!
0%
b100 *
0-
02
b100 6
#740250000000
1!
1%
1-
12
#740260000000
0!
0%
b101 *
0-
02
b101 6
#740270000000
1!
1%
1-
12
#740280000000
0!
0%
b110 *
0-
02
b110 6
#740290000000
1!
1%
1-
12
#740300000000
0!
0%
b111 *
0-
02
b111 6
#740310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#740320000000
0!
0%
b0 *
0-
02
b0 6
#740330000000
1!
1%
1-
12
#740340000000
0!
0%
b1 *
0-
02
b1 6
#740350000000
1!
1%
1-
12
#740360000000
0!
0%
b10 *
0-
02
b10 6
#740370000000
1!
1%
1-
12
#740380000000
0!
0%
b11 *
0-
02
b11 6
#740390000000
1!
1%
1-
12
15
#740400000000
0!
0%
b100 *
0-
02
b100 6
#740410000000
1!
1%
1-
12
#740420000000
0!
0%
b101 *
0-
02
b101 6
#740430000000
1!
1%
1-
12
#740440000000
0!
0%
b110 *
0-
02
b110 6
#740450000000
1!
1%
1-
12
#740460000000
0!
0%
b111 *
0-
02
b111 6
#740470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#740480000000
0!
0%
b0 *
0-
02
b0 6
#740490000000
1!
1%
1-
12
#740500000000
0!
0%
b1 *
0-
02
b1 6
#740510000000
1!
1%
1-
12
#740520000000
0!
0%
b10 *
0-
02
b10 6
#740530000000
1!
1%
1-
12
#740540000000
0!
0%
b11 *
0-
02
b11 6
#740550000000
1!
1%
1-
12
15
#740560000000
0!
0%
b100 *
0-
02
b100 6
#740570000000
1!
1%
1-
12
#740580000000
0!
0%
b101 *
0-
02
b101 6
#740590000000
1!
1%
1-
12
#740600000000
0!
0%
b110 *
0-
02
b110 6
#740610000000
1!
1%
1-
12
#740620000000
0!
0%
b111 *
0-
02
b111 6
#740630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#740640000000
0!
0%
b0 *
0-
02
b0 6
#740650000000
1!
1%
1-
12
#740660000000
0!
0%
b1 *
0-
02
b1 6
#740670000000
1!
1%
1-
12
#740680000000
0!
0%
b10 *
0-
02
b10 6
#740690000000
1!
1%
1-
12
#740700000000
0!
0%
b11 *
0-
02
b11 6
#740710000000
1!
1%
1-
12
15
#740720000000
0!
0%
b100 *
0-
02
b100 6
#740730000000
1!
1%
1-
12
#740740000000
0!
0%
b101 *
0-
02
b101 6
#740750000000
1!
1%
1-
12
#740760000000
0!
0%
b110 *
0-
02
b110 6
#740770000000
1!
1%
1-
12
#740780000000
0!
0%
b111 *
0-
02
b111 6
#740790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#740800000000
0!
0%
b0 *
0-
02
b0 6
#740810000000
1!
1%
1-
12
#740820000000
0!
0%
b1 *
0-
02
b1 6
#740830000000
1!
1%
1-
12
#740840000000
0!
0%
b10 *
0-
02
b10 6
#740850000000
1!
1%
1-
12
#740860000000
0!
0%
b11 *
0-
02
b11 6
#740870000000
1!
1%
1-
12
15
#740880000000
0!
0%
b100 *
0-
02
b100 6
#740890000000
1!
1%
1-
12
#740900000000
0!
0%
b101 *
0-
02
b101 6
#740910000000
1!
1%
1-
12
#740920000000
0!
0%
b110 *
0-
02
b110 6
#740930000000
1!
1%
1-
12
#740940000000
0!
0%
b111 *
0-
02
b111 6
#740950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#740960000000
0!
0%
b0 *
0-
02
b0 6
#740970000000
1!
1%
1-
12
#740980000000
0!
0%
b1 *
0-
02
b1 6
#740990000000
1!
1%
1-
12
#741000000000
0!
0%
b10 *
0-
02
b10 6
#741010000000
1!
1%
1-
12
#741020000000
0!
0%
b11 *
0-
02
b11 6
#741030000000
1!
1%
1-
12
15
#741040000000
0!
0%
b100 *
0-
02
b100 6
#741050000000
1!
1%
1-
12
#741060000000
0!
0%
b101 *
0-
02
b101 6
#741070000000
1!
1%
1-
12
#741080000000
0!
0%
b110 *
0-
02
b110 6
#741090000000
1!
1%
1-
12
#741100000000
0!
0%
b111 *
0-
02
b111 6
#741110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#741120000000
0!
0%
b0 *
0-
02
b0 6
#741130000000
1!
1%
1-
12
#741140000000
0!
0%
b1 *
0-
02
b1 6
#741150000000
1!
1%
1-
12
#741160000000
0!
0%
b10 *
0-
02
b10 6
#741170000000
1!
1%
1-
12
#741180000000
0!
0%
b11 *
0-
02
b11 6
#741190000000
1!
1%
1-
12
15
#741200000000
0!
0%
b100 *
0-
02
b100 6
#741210000000
1!
1%
1-
12
#741220000000
0!
0%
b101 *
0-
02
b101 6
#741230000000
1!
1%
1-
12
#741240000000
0!
0%
b110 *
0-
02
b110 6
#741250000000
1!
1%
1-
12
#741260000000
0!
0%
b111 *
0-
02
b111 6
#741270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#741280000000
0!
0%
b0 *
0-
02
b0 6
#741290000000
1!
1%
1-
12
#741300000000
0!
0%
b1 *
0-
02
b1 6
#741310000000
1!
1%
1-
12
#741320000000
0!
0%
b10 *
0-
02
b10 6
#741330000000
1!
1%
1-
12
#741340000000
0!
0%
b11 *
0-
02
b11 6
#741350000000
1!
1%
1-
12
15
#741360000000
0!
0%
b100 *
0-
02
b100 6
#741370000000
1!
1%
1-
12
#741380000000
0!
0%
b101 *
0-
02
b101 6
#741390000000
1!
1%
1-
12
#741400000000
0!
0%
b110 *
0-
02
b110 6
#741410000000
1!
1%
1-
12
#741420000000
0!
0%
b111 *
0-
02
b111 6
#741430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#741440000000
0!
0%
b0 *
0-
02
b0 6
#741450000000
1!
1%
1-
12
#741460000000
0!
0%
b1 *
0-
02
b1 6
#741470000000
1!
1%
1-
12
#741480000000
0!
0%
b10 *
0-
02
b10 6
#741490000000
1!
1%
1-
12
#741500000000
0!
0%
b11 *
0-
02
b11 6
#741510000000
1!
1%
1-
12
15
#741520000000
0!
0%
b100 *
0-
02
b100 6
#741530000000
1!
1%
1-
12
#741540000000
0!
0%
b101 *
0-
02
b101 6
#741550000000
1!
1%
1-
12
#741560000000
0!
0%
b110 *
0-
02
b110 6
#741570000000
1!
1%
1-
12
#741580000000
0!
0%
b111 *
0-
02
b111 6
#741590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#741600000000
0!
0%
b0 *
0-
02
b0 6
#741610000000
1!
1%
1-
12
#741620000000
0!
0%
b1 *
0-
02
b1 6
#741630000000
1!
1%
1-
12
#741640000000
0!
0%
b10 *
0-
02
b10 6
#741650000000
1!
1%
1-
12
#741660000000
0!
0%
b11 *
0-
02
b11 6
#741670000000
1!
1%
1-
12
15
#741680000000
0!
0%
b100 *
0-
02
b100 6
#741690000000
1!
1%
1-
12
#741700000000
0!
0%
b101 *
0-
02
b101 6
#741710000000
1!
1%
1-
12
#741720000000
0!
0%
b110 *
0-
02
b110 6
#741730000000
1!
1%
1-
12
#741740000000
0!
0%
b111 *
0-
02
b111 6
#741750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#741760000000
0!
0%
b0 *
0-
02
b0 6
#741770000000
1!
1%
1-
12
#741780000000
0!
0%
b1 *
0-
02
b1 6
#741790000000
1!
1%
1-
12
#741800000000
0!
0%
b10 *
0-
02
b10 6
#741810000000
1!
1%
1-
12
#741820000000
0!
0%
b11 *
0-
02
b11 6
#741830000000
1!
1%
1-
12
15
#741840000000
0!
0%
b100 *
0-
02
b100 6
#741850000000
1!
1%
1-
12
#741860000000
0!
0%
b101 *
0-
02
b101 6
#741870000000
1!
1%
1-
12
#741880000000
0!
0%
b110 *
0-
02
b110 6
#741890000000
1!
1%
1-
12
#741900000000
0!
0%
b111 *
0-
02
b111 6
#741910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#741920000000
0!
0%
b0 *
0-
02
b0 6
#741930000000
1!
1%
1-
12
#741940000000
0!
0%
b1 *
0-
02
b1 6
#741950000000
1!
1%
1-
12
#741960000000
0!
0%
b10 *
0-
02
b10 6
#741970000000
1!
1%
1-
12
#741980000000
0!
0%
b11 *
0-
02
b11 6
#741990000000
1!
1%
1-
12
15
#742000000000
0!
0%
b100 *
0-
02
b100 6
#742010000000
1!
1%
1-
12
#742020000000
0!
0%
b101 *
0-
02
b101 6
#742030000000
1!
1%
1-
12
#742040000000
0!
0%
b110 *
0-
02
b110 6
#742050000000
1!
1%
1-
12
#742060000000
0!
0%
b111 *
0-
02
b111 6
#742070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#742080000000
0!
0%
b0 *
0-
02
b0 6
#742090000000
1!
1%
1-
12
#742100000000
0!
0%
b1 *
0-
02
b1 6
#742110000000
1!
1%
1-
12
#742120000000
0!
0%
b10 *
0-
02
b10 6
#742130000000
1!
1%
1-
12
#742140000000
0!
0%
b11 *
0-
02
b11 6
#742150000000
1!
1%
1-
12
15
#742160000000
0!
0%
b100 *
0-
02
b100 6
#742170000000
1!
1%
1-
12
#742180000000
0!
0%
b101 *
0-
02
b101 6
#742190000000
1!
1%
1-
12
#742200000000
0!
0%
b110 *
0-
02
b110 6
#742210000000
1!
1%
1-
12
#742220000000
0!
0%
b111 *
0-
02
b111 6
#742230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#742240000000
0!
0%
b0 *
0-
02
b0 6
#742250000000
1!
1%
1-
12
#742260000000
0!
0%
b1 *
0-
02
b1 6
#742270000000
1!
1%
1-
12
#742280000000
0!
0%
b10 *
0-
02
b10 6
#742290000000
1!
1%
1-
12
#742300000000
0!
0%
b11 *
0-
02
b11 6
#742310000000
1!
1%
1-
12
15
#742320000000
0!
0%
b100 *
0-
02
b100 6
#742330000000
1!
1%
1-
12
#742340000000
0!
0%
b101 *
0-
02
b101 6
#742350000000
1!
1%
1-
12
#742360000000
0!
0%
b110 *
0-
02
b110 6
#742370000000
1!
1%
1-
12
#742380000000
0!
0%
b111 *
0-
02
b111 6
#742390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#742400000000
0!
0%
b0 *
0-
02
b0 6
#742410000000
1!
1%
1-
12
#742420000000
0!
0%
b1 *
0-
02
b1 6
#742430000000
1!
1%
1-
12
#742440000000
0!
0%
b10 *
0-
02
b10 6
#742450000000
1!
1%
1-
12
#742460000000
0!
0%
b11 *
0-
02
b11 6
#742470000000
1!
1%
1-
12
15
#742480000000
0!
0%
b100 *
0-
02
b100 6
#742490000000
1!
1%
1-
12
#742500000000
0!
0%
b101 *
0-
02
b101 6
#742510000000
1!
1%
1-
12
#742520000000
0!
0%
b110 *
0-
02
b110 6
#742530000000
1!
1%
1-
12
#742540000000
0!
0%
b111 *
0-
02
b111 6
#742550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#742560000000
0!
0%
b0 *
0-
02
b0 6
#742570000000
1!
1%
1-
12
#742580000000
0!
0%
b1 *
0-
02
b1 6
#742590000000
1!
1%
1-
12
#742600000000
0!
0%
b10 *
0-
02
b10 6
#742610000000
1!
1%
1-
12
#742620000000
0!
0%
b11 *
0-
02
b11 6
#742630000000
1!
1%
1-
12
15
#742640000000
0!
0%
b100 *
0-
02
b100 6
#742650000000
1!
1%
1-
12
#742660000000
0!
0%
b101 *
0-
02
b101 6
#742670000000
1!
1%
1-
12
#742680000000
0!
0%
b110 *
0-
02
b110 6
#742690000000
1!
1%
1-
12
#742700000000
0!
0%
b111 *
0-
02
b111 6
#742710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#742720000000
0!
0%
b0 *
0-
02
b0 6
#742730000000
1!
1%
1-
12
#742740000000
0!
0%
b1 *
0-
02
b1 6
#742750000000
1!
1%
1-
12
#742760000000
0!
0%
b10 *
0-
02
b10 6
#742770000000
1!
1%
1-
12
#742780000000
0!
0%
b11 *
0-
02
b11 6
#742790000000
1!
1%
1-
12
15
#742800000000
0!
0%
b100 *
0-
02
b100 6
#742810000000
1!
1%
1-
12
#742820000000
0!
0%
b101 *
0-
02
b101 6
#742830000000
1!
1%
1-
12
#742840000000
0!
0%
b110 *
0-
02
b110 6
#742850000000
1!
1%
1-
12
#742860000000
0!
0%
b111 *
0-
02
b111 6
#742870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#742880000000
0!
0%
b0 *
0-
02
b0 6
#742890000000
1!
1%
1-
12
#742900000000
0!
0%
b1 *
0-
02
b1 6
#742910000000
1!
1%
1-
12
#742920000000
0!
0%
b10 *
0-
02
b10 6
#742930000000
1!
1%
1-
12
#742940000000
0!
0%
b11 *
0-
02
b11 6
#742950000000
1!
1%
1-
12
15
#742960000000
0!
0%
b100 *
0-
02
b100 6
#742970000000
1!
1%
1-
12
#742980000000
0!
0%
b101 *
0-
02
b101 6
#742990000000
1!
1%
1-
12
#743000000000
0!
0%
b110 *
0-
02
b110 6
#743010000000
1!
1%
1-
12
#743020000000
0!
0%
b111 *
0-
02
b111 6
#743030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#743040000000
0!
0%
b0 *
0-
02
b0 6
#743050000000
1!
1%
1-
12
#743060000000
0!
0%
b1 *
0-
02
b1 6
#743070000000
1!
1%
1-
12
#743080000000
0!
0%
b10 *
0-
02
b10 6
#743090000000
1!
1%
1-
12
#743100000000
0!
0%
b11 *
0-
02
b11 6
#743110000000
1!
1%
1-
12
15
#743120000000
0!
0%
b100 *
0-
02
b100 6
#743130000000
1!
1%
1-
12
#743140000000
0!
0%
b101 *
0-
02
b101 6
#743150000000
1!
1%
1-
12
#743160000000
0!
0%
b110 *
0-
02
b110 6
#743170000000
1!
1%
1-
12
#743180000000
0!
0%
b111 *
0-
02
b111 6
#743190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#743200000000
0!
0%
b0 *
0-
02
b0 6
#743210000000
1!
1%
1-
12
#743220000000
0!
0%
b1 *
0-
02
b1 6
#743230000000
1!
1%
1-
12
#743240000000
0!
0%
b10 *
0-
02
b10 6
#743250000000
1!
1%
1-
12
#743260000000
0!
0%
b11 *
0-
02
b11 6
#743270000000
1!
1%
1-
12
15
#743280000000
0!
0%
b100 *
0-
02
b100 6
#743290000000
1!
1%
1-
12
#743300000000
0!
0%
b101 *
0-
02
b101 6
#743310000000
1!
1%
1-
12
#743320000000
0!
0%
b110 *
0-
02
b110 6
#743330000000
1!
1%
1-
12
#743340000000
0!
0%
b111 *
0-
02
b111 6
#743350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#743360000000
0!
0%
b0 *
0-
02
b0 6
#743370000000
1!
1%
1-
12
#743380000000
0!
0%
b1 *
0-
02
b1 6
#743390000000
1!
1%
1-
12
#743400000000
0!
0%
b10 *
0-
02
b10 6
#743410000000
1!
1%
1-
12
#743420000000
0!
0%
b11 *
0-
02
b11 6
#743430000000
1!
1%
1-
12
15
#743440000000
0!
0%
b100 *
0-
02
b100 6
#743450000000
1!
1%
1-
12
#743460000000
0!
0%
b101 *
0-
02
b101 6
#743470000000
1!
1%
1-
12
#743480000000
0!
0%
b110 *
0-
02
b110 6
#743490000000
1!
1%
1-
12
#743500000000
0!
0%
b111 *
0-
02
b111 6
#743510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#743520000000
0!
0%
b0 *
0-
02
b0 6
#743530000000
1!
1%
1-
12
#743540000000
0!
0%
b1 *
0-
02
b1 6
#743550000000
1!
1%
1-
12
#743560000000
0!
0%
b10 *
0-
02
b10 6
#743570000000
1!
1%
1-
12
#743580000000
0!
0%
b11 *
0-
02
b11 6
#743590000000
1!
1%
1-
12
15
#743600000000
0!
0%
b100 *
0-
02
b100 6
#743610000000
1!
1%
1-
12
#743620000000
0!
0%
b101 *
0-
02
b101 6
#743630000000
1!
1%
1-
12
#743640000000
0!
0%
b110 *
0-
02
b110 6
#743650000000
1!
1%
1-
12
#743660000000
0!
0%
b111 *
0-
02
b111 6
#743670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#743680000000
0!
0%
b0 *
0-
02
b0 6
#743690000000
1!
1%
1-
12
#743700000000
0!
0%
b1 *
0-
02
b1 6
#743710000000
1!
1%
1-
12
#743720000000
0!
0%
b10 *
0-
02
b10 6
#743730000000
1!
1%
1-
12
#743740000000
0!
0%
b11 *
0-
02
b11 6
#743750000000
1!
1%
1-
12
15
#743760000000
0!
0%
b100 *
0-
02
b100 6
#743770000000
1!
1%
1-
12
#743780000000
0!
0%
b101 *
0-
02
b101 6
#743790000000
1!
1%
1-
12
#743800000000
0!
0%
b110 *
0-
02
b110 6
#743810000000
1!
1%
1-
12
#743820000000
0!
0%
b111 *
0-
02
b111 6
#743830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#743840000000
0!
0%
b0 *
0-
02
b0 6
#743850000000
1!
1%
1-
12
#743860000000
0!
0%
b1 *
0-
02
b1 6
#743870000000
1!
1%
1-
12
#743880000000
0!
0%
b10 *
0-
02
b10 6
#743890000000
1!
1%
1-
12
#743900000000
0!
0%
b11 *
0-
02
b11 6
#743910000000
1!
1%
1-
12
15
#743920000000
0!
0%
b100 *
0-
02
b100 6
#743930000000
1!
1%
1-
12
#743940000000
0!
0%
b101 *
0-
02
b101 6
#743950000000
1!
1%
1-
12
#743960000000
0!
0%
b110 *
0-
02
b110 6
#743970000000
1!
1%
1-
12
#743980000000
0!
0%
b111 *
0-
02
b111 6
#743990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#744000000000
0!
0%
b0 *
0-
02
b0 6
#744010000000
1!
1%
1-
12
#744020000000
0!
0%
b1 *
0-
02
b1 6
#744030000000
1!
1%
1-
12
#744040000000
0!
0%
b10 *
0-
02
b10 6
#744050000000
1!
1%
1-
12
#744060000000
0!
0%
b11 *
0-
02
b11 6
#744070000000
1!
1%
1-
12
15
#744080000000
0!
0%
b100 *
0-
02
b100 6
#744090000000
1!
1%
1-
12
#744100000000
0!
0%
b101 *
0-
02
b101 6
#744110000000
1!
1%
1-
12
#744120000000
0!
0%
b110 *
0-
02
b110 6
#744130000000
1!
1%
1-
12
#744140000000
0!
0%
b111 *
0-
02
b111 6
#744150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#744160000000
0!
0%
b0 *
0-
02
b0 6
#744170000000
1!
1%
1-
12
#744180000000
0!
0%
b1 *
0-
02
b1 6
#744190000000
1!
1%
1-
12
#744200000000
0!
0%
b10 *
0-
02
b10 6
#744210000000
1!
1%
1-
12
#744220000000
0!
0%
b11 *
0-
02
b11 6
#744230000000
1!
1%
1-
12
15
#744240000000
0!
0%
b100 *
0-
02
b100 6
#744250000000
1!
1%
1-
12
#744260000000
0!
0%
b101 *
0-
02
b101 6
#744270000000
1!
1%
1-
12
#744280000000
0!
0%
b110 *
0-
02
b110 6
#744290000000
1!
1%
1-
12
#744300000000
0!
0%
b111 *
0-
02
b111 6
#744310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#744320000000
0!
0%
b0 *
0-
02
b0 6
#744330000000
1!
1%
1-
12
#744340000000
0!
0%
b1 *
0-
02
b1 6
#744350000000
1!
1%
1-
12
#744360000000
0!
0%
b10 *
0-
02
b10 6
#744370000000
1!
1%
1-
12
#744380000000
0!
0%
b11 *
0-
02
b11 6
#744390000000
1!
1%
1-
12
15
#744400000000
0!
0%
b100 *
0-
02
b100 6
#744410000000
1!
1%
1-
12
#744420000000
0!
0%
b101 *
0-
02
b101 6
#744430000000
1!
1%
1-
12
#744440000000
0!
0%
b110 *
0-
02
b110 6
#744450000000
1!
1%
1-
12
#744460000000
0!
0%
b111 *
0-
02
b111 6
#744470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#744480000000
0!
0%
b0 *
0-
02
b0 6
#744490000000
1!
1%
1-
12
#744500000000
0!
0%
b1 *
0-
02
b1 6
#744510000000
1!
1%
1-
12
#744520000000
0!
0%
b10 *
0-
02
b10 6
#744530000000
1!
1%
1-
12
#744540000000
0!
0%
b11 *
0-
02
b11 6
#744550000000
1!
1%
1-
12
15
#744560000000
0!
0%
b100 *
0-
02
b100 6
#744570000000
1!
1%
1-
12
#744580000000
0!
0%
b101 *
0-
02
b101 6
#744590000000
1!
1%
1-
12
#744600000000
0!
0%
b110 *
0-
02
b110 6
#744610000000
1!
1%
1-
12
#744620000000
0!
0%
b111 *
0-
02
b111 6
#744630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#744640000000
0!
0%
b0 *
0-
02
b0 6
#744650000000
1!
1%
1-
12
#744660000000
0!
0%
b1 *
0-
02
b1 6
#744670000000
1!
1%
1-
12
#744680000000
0!
0%
b10 *
0-
02
b10 6
#744690000000
1!
1%
1-
12
#744700000000
0!
0%
b11 *
0-
02
b11 6
#744710000000
1!
1%
1-
12
15
#744720000000
0!
0%
b100 *
0-
02
b100 6
#744730000000
1!
1%
1-
12
#744740000000
0!
0%
b101 *
0-
02
b101 6
#744750000000
1!
1%
1-
12
#744760000000
0!
0%
b110 *
0-
02
b110 6
#744770000000
1!
1%
1-
12
#744780000000
0!
0%
b111 *
0-
02
b111 6
#744790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#744800000000
0!
0%
b0 *
0-
02
b0 6
#744810000000
1!
1%
1-
12
#744820000000
0!
0%
b1 *
0-
02
b1 6
#744830000000
1!
1%
1-
12
#744840000000
0!
0%
b10 *
0-
02
b10 6
#744850000000
1!
1%
1-
12
#744860000000
0!
0%
b11 *
0-
02
b11 6
#744870000000
1!
1%
1-
12
15
#744880000000
0!
0%
b100 *
0-
02
b100 6
#744890000000
1!
1%
1-
12
#744900000000
0!
0%
b101 *
0-
02
b101 6
#744910000000
1!
1%
1-
12
#744920000000
0!
0%
b110 *
0-
02
b110 6
#744930000000
1!
1%
1-
12
#744940000000
0!
0%
b111 *
0-
02
b111 6
#744950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#744960000000
0!
0%
b0 *
0-
02
b0 6
#744970000000
1!
1%
1-
12
#744980000000
0!
0%
b1 *
0-
02
b1 6
#744990000000
1!
1%
1-
12
#745000000000
0!
0%
b10 *
0-
02
b10 6
#745010000000
1!
1%
1-
12
#745020000000
0!
0%
b11 *
0-
02
b11 6
#745030000000
1!
1%
1-
12
15
#745040000000
0!
0%
b100 *
0-
02
b100 6
#745050000000
1!
1%
1-
12
#745060000000
0!
0%
b101 *
0-
02
b101 6
#745070000000
1!
1%
1-
12
#745080000000
0!
0%
b110 *
0-
02
b110 6
#745090000000
1!
1%
1-
12
#745100000000
0!
0%
b111 *
0-
02
b111 6
#745110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#745120000000
0!
0%
b0 *
0-
02
b0 6
#745130000000
1!
1%
1-
12
#745140000000
0!
0%
b1 *
0-
02
b1 6
#745150000000
1!
1%
1-
12
#745160000000
0!
0%
b10 *
0-
02
b10 6
#745170000000
1!
1%
1-
12
#745180000000
0!
0%
b11 *
0-
02
b11 6
#745190000000
1!
1%
1-
12
15
#745200000000
0!
0%
b100 *
0-
02
b100 6
#745210000000
1!
1%
1-
12
#745220000000
0!
0%
b101 *
0-
02
b101 6
#745230000000
1!
1%
1-
12
#745240000000
0!
0%
b110 *
0-
02
b110 6
#745250000000
1!
1%
1-
12
#745260000000
0!
0%
b111 *
0-
02
b111 6
#745270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#745280000000
0!
0%
b0 *
0-
02
b0 6
#745290000000
1!
1%
1-
12
#745300000000
0!
0%
b1 *
0-
02
b1 6
#745310000000
1!
1%
1-
12
#745320000000
0!
0%
b10 *
0-
02
b10 6
#745330000000
1!
1%
1-
12
#745340000000
0!
0%
b11 *
0-
02
b11 6
#745350000000
1!
1%
1-
12
15
#745360000000
0!
0%
b100 *
0-
02
b100 6
#745370000000
1!
1%
1-
12
#745380000000
0!
0%
b101 *
0-
02
b101 6
#745390000000
1!
1%
1-
12
#745400000000
0!
0%
b110 *
0-
02
b110 6
#745410000000
1!
1%
1-
12
#745420000000
0!
0%
b111 *
0-
02
b111 6
#745430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#745440000000
0!
0%
b0 *
0-
02
b0 6
#745450000000
1!
1%
1-
12
#745460000000
0!
0%
b1 *
0-
02
b1 6
#745470000000
1!
1%
1-
12
#745480000000
0!
0%
b10 *
0-
02
b10 6
#745490000000
1!
1%
1-
12
#745500000000
0!
0%
b11 *
0-
02
b11 6
#745510000000
1!
1%
1-
12
15
#745520000000
0!
0%
b100 *
0-
02
b100 6
#745530000000
1!
1%
1-
12
#745540000000
0!
0%
b101 *
0-
02
b101 6
#745550000000
1!
1%
1-
12
#745560000000
0!
0%
b110 *
0-
02
b110 6
#745570000000
1!
1%
1-
12
#745580000000
0!
0%
b111 *
0-
02
b111 6
#745590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#745600000000
0!
0%
b0 *
0-
02
b0 6
#745610000000
1!
1%
1-
12
#745620000000
0!
0%
b1 *
0-
02
b1 6
#745630000000
1!
1%
1-
12
#745640000000
0!
0%
b10 *
0-
02
b10 6
#745650000000
1!
1%
1-
12
#745660000000
0!
0%
b11 *
0-
02
b11 6
#745670000000
1!
1%
1-
12
15
#745680000000
0!
0%
b100 *
0-
02
b100 6
#745690000000
1!
1%
1-
12
#745700000000
0!
0%
b101 *
0-
02
b101 6
#745710000000
1!
1%
1-
12
#745720000000
0!
0%
b110 *
0-
02
b110 6
#745730000000
1!
1%
1-
12
#745740000000
0!
0%
b111 *
0-
02
b111 6
#745750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#745760000000
0!
0%
b0 *
0-
02
b0 6
#745770000000
1!
1%
1-
12
#745780000000
0!
0%
b1 *
0-
02
b1 6
#745790000000
1!
1%
1-
12
#745800000000
0!
0%
b10 *
0-
02
b10 6
#745810000000
1!
1%
1-
12
#745820000000
0!
0%
b11 *
0-
02
b11 6
#745830000000
1!
1%
1-
12
15
#745840000000
0!
0%
b100 *
0-
02
b100 6
#745850000000
1!
1%
1-
12
#745860000000
0!
0%
b101 *
0-
02
b101 6
#745870000000
1!
1%
1-
12
#745880000000
0!
0%
b110 *
0-
02
b110 6
#745890000000
1!
1%
1-
12
#745900000000
0!
0%
b111 *
0-
02
b111 6
#745910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#745920000000
0!
0%
b0 *
0-
02
b0 6
#745930000000
1!
1%
1-
12
#745940000000
0!
0%
b1 *
0-
02
b1 6
#745950000000
1!
1%
1-
12
#745960000000
0!
0%
b10 *
0-
02
b10 6
#745970000000
1!
1%
1-
12
#745980000000
0!
0%
b11 *
0-
02
b11 6
#745990000000
1!
1%
1-
12
15
#746000000000
0!
0%
b100 *
0-
02
b100 6
#746010000000
1!
1%
1-
12
#746020000000
0!
0%
b101 *
0-
02
b101 6
#746030000000
1!
1%
1-
12
#746040000000
0!
0%
b110 *
0-
02
b110 6
#746050000000
1!
1%
1-
12
#746060000000
0!
0%
b111 *
0-
02
b111 6
#746070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#746080000000
0!
0%
b0 *
0-
02
b0 6
#746090000000
1!
1%
1-
12
#746100000000
0!
0%
b1 *
0-
02
b1 6
#746110000000
1!
1%
1-
12
#746120000000
0!
0%
b10 *
0-
02
b10 6
#746130000000
1!
1%
1-
12
#746140000000
0!
0%
b11 *
0-
02
b11 6
#746150000000
1!
1%
1-
12
15
#746160000000
0!
0%
b100 *
0-
02
b100 6
#746170000000
1!
1%
1-
12
#746180000000
0!
0%
b101 *
0-
02
b101 6
#746190000000
1!
1%
1-
12
#746200000000
0!
0%
b110 *
0-
02
b110 6
#746210000000
1!
1%
1-
12
#746220000000
0!
0%
b111 *
0-
02
b111 6
#746230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#746240000000
0!
0%
b0 *
0-
02
b0 6
#746250000000
1!
1%
1-
12
#746260000000
0!
0%
b1 *
0-
02
b1 6
#746270000000
1!
1%
1-
12
#746280000000
0!
0%
b10 *
0-
02
b10 6
#746290000000
1!
1%
1-
12
#746300000000
0!
0%
b11 *
0-
02
b11 6
#746310000000
1!
1%
1-
12
15
#746320000000
0!
0%
b100 *
0-
02
b100 6
#746330000000
1!
1%
1-
12
#746340000000
0!
0%
b101 *
0-
02
b101 6
#746350000000
1!
1%
1-
12
#746360000000
0!
0%
b110 *
0-
02
b110 6
#746370000000
1!
1%
1-
12
#746380000000
0!
0%
b111 *
0-
02
b111 6
#746390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#746400000000
0!
0%
b0 *
0-
02
b0 6
#746410000000
1!
1%
1-
12
#746420000000
0!
0%
b1 *
0-
02
b1 6
#746430000000
1!
1%
1-
12
#746440000000
0!
0%
b10 *
0-
02
b10 6
#746450000000
1!
1%
1-
12
#746460000000
0!
0%
b11 *
0-
02
b11 6
#746470000000
1!
1%
1-
12
15
#746480000000
0!
0%
b100 *
0-
02
b100 6
#746490000000
1!
1%
1-
12
#746500000000
0!
0%
b101 *
0-
02
b101 6
#746510000000
1!
1%
1-
12
#746520000000
0!
0%
b110 *
0-
02
b110 6
#746530000000
1!
1%
1-
12
#746540000000
0!
0%
b111 *
0-
02
b111 6
#746550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#746560000000
0!
0%
b0 *
0-
02
b0 6
#746570000000
1!
1%
1-
12
#746580000000
0!
0%
b1 *
0-
02
b1 6
#746590000000
1!
1%
1-
12
#746600000000
0!
0%
b10 *
0-
02
b10 6
#746610000000
1!
1%
1-
12
#746620000000
0!
0%
b11 *
0-
02
b11 6
#746630000000
1!
1%
1-
12
15
#746640000000
0!
0%
b100 *
0-
02
b100 6
#746650000000
1!
1%
1-
12
#746660000000
0!
0%
b101 *
0-
02
b101 6
#746670000000
1!
1%
1-
12
#746680000000
0!
0%
b110 *
0-
02
b110 6
#746690000000
1!
1%
1-
12
#746700000000
0!
0%
b111 *
0-
02
b111 6
#746710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#746720000000
0!
0%
b0 *
0-
02
b0 6
#746730000000
1!
1%
1-
12
#746740000000
0!
0%
b1 *
0-
02
b1 6
#746750000000
1!
1%
1-
12
#746760000000
0!
0%
b10 *
0-
02
b10 6
#746770000000
1!
1%
1-
12
#746780000000
0!
0%
b11 *
0-
02
b11 6
#746790000000
1!
1%
1-
12
15
#746800000000
0!
0%
b100 *
0-
02
b100 6
#746810000000
1!
1%
1-
12
#746820000000
0!
0%
b101 *
0-
02
b101 6
#746830000000
1!
1%
1-
12
#746840000000
0!
0%
b110 *
0-
02
b110 6
#746850000000
1!
1%
1-
12
#746860000000
0!
0%
b111 *
0-
02
b111 6
#746870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#746880000000
0!
0%
b0 *
0-
02
b0 6
#746890000000
1!
1%
1-
12
#746900000000
0!
0%
b1 *
0-
02
b1 6
#746910000000
1!
1%
1-
12
#746920000000
0!
0%
b10 *
0-
02
b10 6
#746930000000
1!
1%
1-
12
#746940000000
0!
0%
b11 *
0-
02
b11 6
#746950000000
1!
1%
1-
12
15
#746960000000
0!
0%
b100 *
0-
02
b100 6
#746970000000
1!
1%
1-
12
#746980000000
0!
0%
b101 *
0-
02
b101 6
#746990000000
1!
1%
1-
12
#747000000000
0!
0%
b110 *
0-
02
b110 6
#747010000000
1!
1%
1-
12
#747020000000
0!
0%
b111 *
0-
02
b111 6
#747030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#747040000000
0!
0%
b0 *
0-
02
b0 6
#747050000000
1!
1%
1-
12
#747060000000
0!
0%
b1 *
0-
02
b1 6
#747070000000
1!
1%
1-
12
#747080000000
0!
0%
b10 *
0-
02
b10 6
#747090000000
1!
1%
1-
12
#747100000000
0!
0%
b11 *
0-
02
b11 6
#747110000000
1!
1%
1-
12
15
#747120000000
0!
0%
b100 *
0-
02
b100 6
#747130000000
1!
1%
1-
12
#747140000000
0!
0%
b101 *
0-
02
b101 6
#747150000000
1!
1%
1-
12
#747160000000
0!
0%
b110 *
0-
02
b110 6
#747170000000
1!
1%
1-
12
#747180000000
0!
0%
b111 *
0-
02
b111 6
#747190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#747200000000
0!
0%
b0 *
0-
02
b0 6
#747210000000
1!
1%
1-
12
#747220000000
0!
0%
b1 *
0-
02
b1 6
#747230000000
1!
1%
1-
12
#747240000000
0!
0%
b10 *
0-
02
b10 6
#747250000000
1!
1%
1-
12
#747260000000
0!
0%
b11 *
0-
02
b11 6
#747270000000
1!
1%
1-
12
15
#747280000000
0!
0%
b100 *
0-
02
b100 6
#747290000000
1!
1%
1-
12
#747300000000
0!
0%
b101 *
0-
02
b101 6
#747310000000
1!
1%
1-
12
#747320000000
0!
0%
b110 *
0-
02
b110 6
#747330000000
1!
1%
1-
12
#747340000000
0!
0%
b111 *
0-
02
b111 6
#747350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#747360000000
0!
0%
b0 *
0-
02
b0 6
#747370000000
1!
1%
1-
12
#747380000000
0!
0%
b1 *
0-
02
b1 6
#747390000000
1!
1%
1-
12
#747400000000
0!
0%
b10 *
0-
02
b10 6
#747410000000
1!
1%
1-
12
#747420000000
0!
0%
b11 *
0-
02
b11 6
#747430000000
1!
1%
1-
12
15
#747440000000
0!
0%
b100 *
0-
02
b100 6
#747450000000
1!
1%
1-
12
#747460000000
0!
0%
b101 *
0-
02
b101 6
#747470000000
1!
1%
1-
12
#747480000000
0!
0%
b110 *
0-
02
b110 6
#747490000000
1!
1%
1-
12
#747500000000
0!
0%
b111 *
0-
02
b111 6
#747510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#747520000000
0!
0%
b0 *
0-
02
b0 6
#747530000000
1!
1%
1-
12
#747540000000
0!
0%
b1 *
0-
02
b1 6
#747550000000
1!
1%
1-
12
#747560000000
0!
0%
b10 *
0-
02
b10 6
#747570000000
1!
1%
1-
12
#747580000000
0!
0%
b11 *
0-
02
b11 6
#747590000000
1!
1%
1-
12
15
#747600000000
0!
0%
b100 *
0-
02
b100 6
#747610000000
1!
1%
1-
12
#747620000000
0!
0%
b101 *
0-
02
b101 6
#747630000000
1!
1%
1-
12
#747640000000
0!
0%
b110 *
0-
02
b110 6
#747650000000
1!
1%
1-
12
#747660000000
0!
0%
b111 *
0-
02
b111 6
#747670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#747680000000
0!
0%
b0 *
0-
02
b0 6
#747690000000
1!
1%
1-
12
#747700000000
0!
0%
b1 *
0-
02
b1 6
#747710000000
1!
1%
1-
12
#747720000000
0!
0%
b10 *
0-
02
b10 6
#747730000000
1!
1%
1-
12
#747740000000
0!
0%
b11 *
0-
02
b11 6
#747750000000
1!
1%
1-
12
15
#747760000000
0!
0%
b100 *
0-
02
b100 6
#747770000000
1!
1%
1-
12
#747780000000
0!
0%
b101 *
0-
02
b101 6
#747790000000
1!
1%
1-
12
#747800000000
0!
0%
b110 *
0-
02
b110 6
#747810000000
1!
1%
1-
12
#747820000000
0!
0%
b111 *
0-
02
b111 6
#747830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#747840000000
0!
0%
b0 *
0-
02
b0 6
#747850000000
1!
1%
1-
12
#747860000000
0!
0%
b1 *
0-
02
b1 6
#747870000000
1!
1%
1-
12
#747880000000
0!
0%
b10 *
0-
02
b10 6
#747890000000
1!
1%
1-
12
#747900000000
0!
0%
b11 *
0-
02
b11 6
#747910000000
1!
1%
1-
12
15
#747920000000
0!
0%
b100 *
0-
02
b100 6
#747930000000
1!
1%
1-
12
#747940000000
0!
0%
b101 *
0-
02
b101 6
#747950000000
1!
1%
1-
12
#747960000000
0!
0%
b110 *
0-
02
b110 6
#747970000000
1!
1%
1-
12
#747980000000
0!
0%
b111 *
0-
02
b111 6
#747990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#748000000000
0!
0%
b0 *
0-
02
b0 6
#748010000000
1!
1%
1-
12
#748020000000
0!
0%
b1 *
0-
02
b1 6
#748030000000
1!
1%
1-
12
#748040000000
0!
0%
b10 *
0-
02
b10 6
#748050000000
1!
1%
1-
12
#748060000000
0!
0%
b11 *
0-
02
b11 6
#748070000000
1!
1%
1-
12
15
#748080000000
0!
0%
b100 *
0-
02
b100 6
#748090000000
1!
1%
1-
12
#748100000000
0!
0%
b101 *
0-
02
b101 6
#748110000000
1!
1%
1-
12
#748120000000
0!
0%
b110 *
0-
02
b110 6
#748130000000
1!
1%
1-
12
#748140000000
0!
0%
b111 *
0-
02
b111 6
#748150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#748160000000
0!
0%
b0 *
0-
02
b0 6
#748170000000
1!
1%
1-
12
#748180000000
0!
0%
b1 *
0-
02
b1 6
#748190000000
1!
1%
1-
12
#748200000000
0!
0%
b10 *
0-
02
b10 6
#748210000000
1!
1%
1-
12
#748220000000
0!
0%
b11 *
0-
02
b11 6
#748230000000
1!
1%
1-
12
15
#748240000000
0!
0%
b100 *
0-
02
b100 6
#748250000000
1!
1%
1-
12
#748260000000
0!
0%
b101 *
0-
02
b101 6
#748270000000
1!
1%
1-
12
#748280000000
0!
0%
b110 *
0-
02
b110 6
#748290000000
1!
1%
1-
12
#748300000000
0!
0%
b111 *
0-
02
b111 6
#748310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#748320000000
0!
0%
b0 *
0-
02
b0 6
#748330000000
1!
1%
1-
12
#748340000000
0!
0%
b1 *
0-
02
b1 6
#748350000000
1!
1%
1-
12
#748360000000
0!
0%
b10 *
0-
02
b10 6
#748370000000
1!
1%
1-
12
#748380000000
0!
0%
b11 *
0-
02
b11 6
#748390000000
1!
1%
1-
12
15
#748400000000
0!
0%
b100 *
0-
02
b100 6
#748410000000
1!
1%
1-
12
#748420000000
0!
0%
b101 *
0-
02
b101 6
#748430000000
1!
1%
1-
12
#748440000000
0!
0%
b110 *
0-
02
b110 6
#748450000000
1!
1%
1-
12
#748460000000
0!
0%
b111 *
0-
02
b111 6
#748470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#748480000000
0!
0%
b0 *
0-
02
b0 6
#748490000000
1!
1%
1-
12
#748500000000
0!
0%
b1 *
0-
02
b1 6
#748510000000
1!
1%
1-
12
#748520000000
0!
0%
b10 *
0-
02
b10 6
#748530000000
1!
1%
1-
12
#748540000000
0!
0%
b11 *
0-
02
b11 6
#748550000000
1!
1%
1-
12
15
#748560000000
0!
0%
b100 *
0-
02
b100 6
#748570000000
1!
1%
1-
12
#748580000000
0!
0%
b101 *
0-
02
b101 6
#748590000000
1!
1%
1-
12
#748600000000
0!
0%
b110 *
0-
02
b110 6
#748610000000
1!
1%
1-
12
#748620000000
0!
0%
b111 *
0-
02
b111 6
#748630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#748640000000
0!
0%
b0 *
0-
02
b0 6
#748650000000
1!
1%
1-
12
#748660000000
0!
0%
b1 *
0-
02
b1 6
#748670000000
1!
1%
1-
12
#748680000000
0!
0%
b10 *
0-
02
b10 6
#748690000000
1!
1%
1-
12
#748700000000
0!
0%
b11 *
0-
02
b11 6
#748710000000
1!
1%
1-
12
15
#748720000000
0!
0%
b100 *
0-
02
b100 6
#748730000000
1!
1%
1-
12
#748740000000
0!
0%
b101 *
0-
02
b101 6
#748750000000
1!
1%
1-
12
#748760000000
0!
0%
b110 *
0-
02
b110 6
#748770000000
1!
1%
1-
12
#748780000000
0!
0%
b111 *
0-
02
b111 6
#748790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#748800000000
0!
0%
b0 *
0-
02
b0 6
#748810000000
1!
1%
1-
12
#748820000000
0!
0%
b1 *
0-
02
b1 6
#748830000000
1!
1%
1-
12
#748840000000
0!
0%
b10 *
0-
02
b10 6
#748850000000
1!
1%
1-
12
#748860000000
0!
0%
b11 *
0-
02
b11 6
#748870000000
1!
1%
1-
12
15
#748880000000
0!
0%
b100 *
0-
02
b100 6
#748890000000
1!
1%
1-
12
#748900000000
0!
0%
b101 *
0-
02
b101 6
#748910000000
1!
1%
1-
12
#748920000000
0!
0%
b110 *
0-
02
b110 6
#748930000000
1!
1%
1-
12
#748940000000
0!
0%
b111 *
0-
02
b111 6
#748950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#748960000000
0!
0%
b0 *
0-
02
b0 6
#748970000000
1!
1%
1-
12
#748980000000
0!
0%
b1 *
0-
02
b1 6
#748990000000
1!
1%
1-
12
#749000000000
0!
0%
b10 *
0-
02
b10 6
#749010000000
1!
1%
1-
12
#749020000000
0!
0%
b11 *
0-
02
b11 6
#749030000000
1!
1%
1-
12
15
#749040000000
0!
0%
b100 *
0-
02
b100 6
#749050000000
1!
1%
1-
12
#749060000000
0!
0%
b101 *
0-
02
b101 6
#749070000000
1!
1%
1-
12
#749080000000
0!
0%
b110 *
0-
02
b110 6
#749090000000
1!
1%
1-
12
#749100000000
0!
0%
b111 *
0-
02
b111 6
#749110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#749120000000
0!
0%
b0 *
0-
02
b0 6
#749130000000
1!
1%
1-
12
#749140000000
0!
0%
b1 *
0-
02
b1 6
#749150000000
1!
1%
1-
12
#749160000000
0!
0%
b10 *
0-
02
b10 6
#749170000000
1!
1%
1-
12
#749180000000
0!
0%
b11 *
0-
02
b11 6
#749190000000
1!
1%
1-
12
15
#749200000000
0!
0%
b100 *
0-
02
b100 6
#749210000000
1!
1%
1-
12
#749220000000
0!
0%
b101 *
0-
02
b101 6
#749230000000
1!
1%
1-
12
#749240000000
0!
0%
b110 *
0-
02
b110 6
#749250000000
1!
1%
1-
12
#749260000000
0!
0%
b111 *
0-
02
b111 6
#749270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#749280000000
0!
0%
b0 *
0-
02
b0 6
#749290000000
1!
1%
1-
12
#749300000000
0!
0%
b1 *
0-
02
b1 6
#749310000000
1!
1%
1-
12
#749320000000
0!
0%
b10 *
0-
02
b10 6
#749330000000
1!
1%
1-
12
#749340000000
0!
0%
b11 *
0-
02
b11 6
#749350000000
1!
1%
1-
12
15
#749360000000
0!
0%
b100 *
0-
02
b100 6
#749370000000
1!
1%
1-
12
#749380000000
0!
0%
b101 *
0-
02
b101 6
#749390000000
1!
1%
1-
12
#749400000000
0!
0%
b110 *
0-
02
b110 6
#749410000000
1!
1%
1-
12
#749420000000
0!
0%
b111 *
0-
02
b111 6
#749430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#749440000000
0!
0%
b0 *
0-
02
b0 6
#749450000000
1!
1%
1-
12
#749460000000
0!
0%
b1 *
0-
02
b1 6
#749470000000
1!
1%
1-
12
#749480000000
0!
0%
b10 *
0-
02
b10 6
#749490000000
1!
1%
1-
12
#749500000000
0!
0%
b11 *
0-
02
b11 6
#749510000000
1!
1%
1-
12
15
#749520000000
0!
0%
b100 *
0-
02
b100 6
#749530000000
1!
1%
1-
12
#749540000000
0!
0%
b101 *
0-
02
b101 6
#749550000000
1!
1%
1-
12
#749560000000
0!
0%
b110 *
0-
02
b110 6
#749570000000
1!
1%
1-
12
#749580000000
0!
0%
b111 *
0-
02
b111 6
#749590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#749600000000
0!
0%
b0 *
0-
02
b0 6
#749610000000
1!
1%
1-
12
#749620000000
0!
0%
b1 *
0-
02
b1 6
#749630000000
1!
1%
1-
12
#749640000000
0!
0%
b10 *
0-
02
b10 6
#749650000000
1!
1%
1-
12
#749660000000
0!
0%
b11 *
0-
02
b11 6
#749670000000
1!
1%
1-
12
15
#749680000000
0!
0%
b100 *
0-
02
b100 6
#749690000000
1!
1%
1-
12
#749700000000
0!
0%
b101 *
0-
02
b101 6
#749710000000
1!
1%
1-
12
#749720000000
0!
0%
b110 *
0-
02
b110 6
#749730000000
1!
1%
1-
12
#749740000000
0!
0%
b111 *
0-
02
b111 6
#749750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#749760000000
0!
0%
b0 *
0-
02
b0 6
#749770000000
1!
1%
1-
12
#749780000000
0!
0%
b1 *
0-
02
b1 6
#749790000000
1!
1%
1-
12
#749800000000
0!
0%
b10 *
0-
02
b10 6
#749810000000
1!
1%
1-
12
#749820000000
0!
0%
b11 *
0-
02
b11 6
#749830000000
1!
1%
1-
12
15
#749840000000
0!
0%
b100 *
0-
02
b100 6
#749850000000
1!
1%
1-
12
#749860000000
0!
0%
b101 *
0-
02
b101 6
#749870000000
1!
1%
1-
12
#749880000000
0!
0%
b110 *
0-
02
b110 6
#749890000000
1!
1%
1-
12
#749900000000
0!
0%
b111 *
0-
02
b111 6
#749910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#749920000000
0!
0%
b0 *
0-
02
b0 6
#749930000000
1!
1%
1-
12
#749940000000
0!
0%
b1 *
0-
02
b1 6
#749950000000
1!
1%
1-
12
#749960000000
0!
0%
b10 *
0-
02
b10 6
#749970000000
1!
1%
1-
12
#749980000000
0!
0%
b11 *
0-
02
b11 6
#749990000000
1!
1%
1-
12
15
#750000000000
0!
0%
b100 *
0-
02
b100 6
#750010000000
1!
1%
1-
12
#750020000000
0!
0%
b101 *
0-
02
b101 6
#750030000000
1!
1%
1-
12
#750040000000
0!
0%
b110 *
0-
02
b110 6
#750050000000
1!
1%
1-
12
#750060000000
0!
0%
b111 *
0-
02
b111 6
#750070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#750080000000
0!
0%
b0 *
0-
02
b0 6
#750090000000
1!
1%
1-
12
#750100000000
0!
0%
b1 *
0-
02
b1 6
#750110000000
1!
1%
1-
12
#750120000000
0!
0%
b10 *
0-
02
b10 6
#750130000000
1!
1%
1-
12
#750140000000
0!
0%
b11 *
0-
02
b11 6
#750150000000
1!
1%
1-
12
15
#750160000000
0!
0%
b100 *
0-
02
b100 6
#750170000000
1!
1%
1-
12
#750180000000
0!
0%
b101 *
0-
02
b101 6
#750190000000
1!
1%
1-
12
#750200000000
0!
0%
b110 *
0-
02
b110 6
#750210000000
1!
1%
1-
12
#750220000000
0!
0%
b111 *
0-
02
b111 6
#750230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#750240000000
0!
0%
b0 *
0-
02
b0 6
#750250000000
1!
1%
1-
12
#750260000000
0!
0%
b1 *
0-
02
b1 6
#750270000000
1!
1%
1-
12
#750280000000
0!
0%
b10 *
0-
02
b10 6
#750290000000
1!
1%
1-
12
#750300000000
0!
0%
b11 *
0-
02
b11 6
#750310000000
1!
1%
1-
12
15
#750320000000
0!
0%
b100 *
0-
02
b100 6
#750330000000
1!
1%
1-
12
#750340000000
0!
0%
b101 *
0-
02
b101 6
#750350000000
1!
1%
1-
12
#750360000000
0!
0%
b110 *
0-
02
b110 6
#750370000000
1!
1%
1-
12
#750380000000
0!
0%
b111 *
0-
02
b111 6
#750390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#750400000000
0!
0%
b0 *
0-
02
b0 6
#750410000000
1!
1%
1-
12
#750420000000
0!
0%
b1 *
0-
02
b1 6
#750430000000
1!
1%
1-
12
#750440000000
0!
0%
b10 *
0-
02
b10 6
#750450000000
1!
1%
1-
12
#750460000000
0!
0%
b11 *
0-
02
b11 6
#750470000000
1!
1%
1-
12
15
#750480000000
0!
0%
b100 *
0-
02
b100 6
#750490000000
1!
1%
1-
12
#750500000000
0!
0%
b101 *
0-
02
b101 6
#750510000000
1!
1%
1-
12
#750520000000
0!
0%
b110 *
0-
02
b110 6
#750530000000
1!
1%
1-
12
#750540000000
0!
0%
b111 *
0-
02
b111 6
#750550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#750560000000
0!
0%
b0 *
0-
02
b0 6
#750570000000
1!
1%
1-
12
#750580000000
0!
0%
b1 *
0-
02
b1 6
#750590000000
1!
1%
1-
12
#750600000000
0!
0%
b10 *
0-
02
b10 6
#750610000000
1!
1%
1-
12
#750620000000
0!
0%
b11 *
0-
02
b11 6
#750630000000
1!
1%
1-
12
15
#750640000000
0!
0%
b100 *
0-
02
b100 6
#750650000000
1!
1%
1-
12
#750660000000
0!
0%
b101 *
0-
02
b101 6
#750670000000
1!
1%
1-
12
#750680000000
0!
0%
b110 *
0-
02
b110 6
#750690000000
1!
1%
1-
12
#750700000000
0!
0%
b111 *
0-
02
b111 6
#750710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#750720000000
0!
0%
b0 *
0-
02
b0 6
#750730000000
1!
1%
1-
12
#750740000000
0!
0%
b1 *
0-
02
b1 6
#750750000000
1!
1%
1-
12
#750760000000
0!
0%
b10 *
0-
02
b10 6
#750770000000
1!
1%
1-
12
#750780000000
0!
0%
b11 *
0-
02
b11 6
#750790000000
1!
1%
1-
12
15
#750800000000
0!
0%
b100 *
0-
02
b100 6
#750810000000
1!
1%
1-
12
#750820000000
0!
0%
b101 *
0-
02
b101 6
#750830000000
1!
1%
1-
12
#750840000000
0!
0%
b110 *
0-
02
b110 6
#750850000000
1!
1%
1-
12
#750860000000
0!
0%
b111 *
0-
02
b111 6
#750870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#750880000000
0!
0%
b0 *
0-
02
b0 6
#750890000000
1!
1%
1-
12
#750900000000
0!
0%
b1 *
0-
02
b1 6
#750910000000
1!
1%
1-
12
#750920000000
0!
0%
b10 *
0-
02
b10 6
#750930000000
1!
1%
1-
12
#750940000000
0!
0%
b11 *
0-
02
b11 6
#750950000000
1!
1%
1-
12
15
#750960000000
0!
0%
b100 *
0-
02
b100 6
#750970000000
1!
1%
1-
12
#750980000000
0!
0%
b101 *
0-
02
b101 6
#750990000000
1!
1%
1-
12
#751000000000
0!
0%
b110 *
0-
02
b110 6
#751010000000
1!
1%
1-
12
#751020000000
0!
0%
b111 *
0-
02
b111 6
#751030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#751040000000
0!
0%
b0 *
0-
02
b0 6
#751050000000
1!
1%
1-
12
#751060000000
0!
0%
b1 *
0-
02
b1 6
#751070000000
1!
1%
1-
12
#751080000000
0!
0%
b10 *
0-
02
b10 6
#751090000000
1!
1%
1-
12
#751100000000
0!
0%
b11 *
0-
02
b11 6
#751110000000
1!
1%
1-
12
15
#751120000000
0!
0%
b100 *
0-
02
b100 6
#751130000000
1!
1%
1-
12
#751140000000
0!
0%
b101 *
0-
02
b101 6
#751150000000
1!
1%
1-
12
#751160000000
0!
0%
b110 *
0-
02
b110 6
#751170000000
1!
1%
1-
12
#751180000000
0!
0%
b111 *
0-
02
b111 6
#751190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#751200000000
0!
0%
b0 *
0-
02
b0 6
#751210000000
1!
1%
1-
12
#751220000000
0!
0%
b1 *
0-
02
b1 6
#751230000000
1!
1%
1-
12
#751240000000
0!
0%
b10 *
0-
02
b10 6
#751250000000
1!
1%
1-
12
#751260000000
0!
0%
b11 *
0-
02
b11 6
#751270000000
1!
1%
1-
12
15
#751280000000
0!
0%
b100 *
0-
02
b100 6
#751290000000
1!
1%
1-
12
#751300000000
0!
0%
b101 *
0-
02
b101 6
#751310000000
1!
1%
1-
12
#751320000000
0!
0%
b110 *
0-
02
b110 6
#751330000000
1!
1%
1-
12
#751340000000
0!
0%
b111 *
0-
02
b111 6
#751350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#751360000000
0!
0%
b0 *
0-
02
b0 6
#751370000000
1!
1%
1-
12
#751380000000
0!
0%
b1 *
0-
02
b1 6
#751390000000
1!
1%
1-
12
#751400000000
0!
0%
b10 *
0-
02
b10 6
#751410000000
1!
1%
1-
12
#751420000000
0!
0%
b11 *
0-
02
b11 6
#751430000000
1!
1%
1-
12
15
#751440000000
0!
0%
b100 *
0-
02
b100 6
#751450000000
1!
1%
1-
12
#751460000000
0!
0%
b101 *
0-
02
b101 6
#751470000000
1!
1%
1-
12
#751480000000
0!
0%
b110 *
0-
02
b110 6
#751490000000
1!
1%
1-
12
#751500000000
0!
0%
b111 *
0-
02
b111 6
#751510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#751520000000
0!
0%
b0 *
0-
02
b0 6
#751530000000
1!
1%
1-
12
#751540000000
0!
0%
b1 *
0-
02
b1 6
#751550000000
1!
1%
1-
12
#751560000000
0!
0%
b10 *
0-
02
b10 6
#751570000000
1!
1%
1-
12
#751580000000
0!
0%
b11 *
0-
02
b11 6
#751590000000
1!
1%
1-
12
15
#751600000000
0!
0%
b100 *
0-
02
b100 6
#751610000000
1!
1%
1-
12
#751620000000
0!
0%
b101 *
0-
02
b101 6
#751630000000
1!
1%
1-
12
#751640000000
0!
0%
b110 *
0-
02
b110 6
#751650000000
1!
1%
1-
12
#751660000000
0!
0%
b111 *
0-
02
b111 6
#751670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#751680000000
0!
0%
b0 *
0-
02
b0 6
#751690000000
1!
1%
1-
12
#751700000000
0!
0%
b1 *
0-
02
b1 6
#751710000000
1!
1%
1-
12
#751720000000
0!
0%
b10 *
0-
02
b10 6
#751730000000
1!
1%
1-
12
#751740000000
0!
0%
b11 *
0-
02
b11 6
#751750000000
1!
1%
1-
12
15
#751760000000
0!
0%
b100 *
0-
02
b100 6
#751770000000
1!
1%
1-
12
#751780000000
0!
0%
b101 *
0-
02
b101 6
#751790000000
1!
1%
1-
12
#751800000000
0!
0%
b110 *
0-
02
b110 6
#751810000000
1!
1%
1-
12
#751820000000
0!
0%
b111 *
0-
02
b111 6
#751830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#751840000000
0!
0%
b0 *
0-
02
b0 6
#751850000000
1!
1%
1-
12
#751860000000
0!
0%
b1 *
0-
02
b1 6
#751870000000
1!
1%
1-
12
#751880000000
0!
0%
b10 *
0-
02
b10 6
#751890000000
1!
1%
1-
12
#751900000000
0!
0%
b11 *
0-
02
b11 6
#751910000000
1!
1%
1-
12
15
#751920000000
0!
0%
b100 *
0-
02
b100 6
#751930000000
1!
1%
1-
12
#751940000000
0!
0%
b101 *
0-
02
b101 6
#751950000000
1!
1%
1-
12
#751960000000
0!
0%
b110 *
0-
02
b110 6
#751970000000
1!
1%
1-
12
#751980000000
0!
0%
b111 *
0-
02
b111 6
#751990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#752000000000
0!
0%
b0 *
0-
02
b0 6
#752010000000
1!
1%
1-
12
#752020000000
0!
0%
b1 *
0-
02
b1 6
#752030000000
1!
1%
1-
12
#752040000000
0!
0%
b10 *
0-
02
b10 6
#752050000000
1!
1%
1-
12
#752060000000
0!
0%
b11 *
0-
02
b11 6
#752070000000
1!
1%
1-
12
15
#752080000000
0!
0%
b100 *
0-
02
b100 6
#752090000000
1!
1%
1-
12
#752100000000
0!
0%
b101 *
0-
02
b101 6
#752110000000
1!
1%
1-
12
#752120000000
0!
0%
b110 *
0-
02
b110 6
#752130000000
1!
1%
1-
12
#752140000000
0!
0%
b111 *
0-
02
b111 6
#752150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#752160000000
0!
0%
b0 *
0-
02
b0 6
#752170000000
1!
1%
1-
12
#752180000000
0!
0%
b1 *
0-
02
b1 6
#752190000000
1!
1%
1-
12
#752200000000
0!
0%
b10 *
0-
02
b10 6
#752210000000
1!
1%
1-
12
#752220000000
0!
0%
b11 *
0-
02
b11 6
#752230000000
1!
1%
1-
12
15
#752240000000
0!
0%
b100 *
0-
02
b100 6
#752250000000
1!
1%
1-
12
#752260000000
0!
0%
b101 *
0-
02
b101 6
#752270000000
1!
1%
1-
12
#752280000000
0!
0%
b110 *
0-
02
b110 6
#752290000000
1!
1%
1-
12
#752300000000
0!
0%
b111 *
0-
02
b111 6
#752310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#752320000000
0!
0%
b0 *
0-
02
b0 6
#752330000000
1!
1%
1-
12
#752340000000
0!
0%
b1 *
0-
02
b1 6
#752350000000
1!
1%
1-
12
#752360000000
0!
0%
b10 *
0-
02
b10 6
#752370000000
1!
1%
1-
12
#752380000000
0!
0%
b11 *
0-
02
b11 6
#752390000000
1!
1%
1-
12
15
#752400000000
0!
0%
b100 *
0-
02
b100 6
#752410000000
1!
1%
1-
12
#752420000000
0!
0%
b101 *
0-
02
b101 6
#752430000000
1!
1%
1-
12
#752440000000
0!
0%
b110 *
0-
02
b110 6
#752450000000
1!
1%
1-
12
#752460000000
0!
0%
b111 *
0-
02
b111 6
#752470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#752480000000
0!
0%
b0 *
0-
02
b0 6
#752490000000
1!
1%
1-
12
#752500000000
0!
0%
b1 *
0-
02
b1 6
#752510000000
1!
1%
1-
12
#752520000000
0!
0%
b10 *
0-
02
b10 6
#752530000000
1!
1%
1-
12
#752540000000
0!
0%
b11 *
0-
02
b11 6
#752550000000
1!
1%
1-
12
15
#752560000000
0!
0%
b100 *
0-
02
b100 6
#752570000000
1!
1%
1-
12
#752580000000
0!
0%
b101 *
0-
02
b101 6
#752590000000
1!
1%
1-
12
#752600000000
0!
0%
b110 *
0-
02
b110 6
#752610000000
1!
1%
1-
12
#752620000000
0!
0%
b111 *
0-
02
b111 6
#752630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#752640000000
0!
0%
b0 *
0-
02
b0 6
#752650000000
1!
1%
1-
12
#752660000000
0!
0%
b1 *
0-
02
b1 6
#752670000000
1!
1%
1-
12
#752680000000
0!
0%
b10 *
0-
02
b10 6
#752690000000
1!
1%
1-
12
#752700000000
0!
0%
b11 *
0-
02
b11 6
#752710000000
1!
1%
1-
12
15
#752720000000
0!
0%
b100 *
0-
02
b100 6
#752730000000
1!
1%
1-
12
#752740000000
0!
0%
b101 *
0-
02
b101 6
#752750000000
1!
1%
1-
12
#752760000000
0!
0%
b110 *
0-
02
b110 6
#752770000000
1!
1%
1-
12
#752780000000
0!
0%
b111 *
0-
02
b111 6
#752790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#752800000000
0!
0%
b0 *
0-
02
b0 6
#752810000000
1!
1%
1-
12
#752820000000
0!
0%
b1 *
0-
02
b1 6
#752830000000
1!
1%
1-
12
#752840000000
0!
0%
b10 *
0-
02
b10 6
#752850000000
1!
1%
1-
12
#752860000000
0!
0%
b11 *
0-
02
b11 6
#752870000000
1!
1%
1-
12
15
#752880000000
0!
0%
b100 *
0-
02
b100 6
#752890000000
1!
1%
1-
12
#752900000000
0!
0%
b101 *
0-
02
b101 6
#752910000000
1!
1%
1-
12
#752920000000
0!
0%
b110 *
0-
02
b110 6
#752930000000
1!
1%
1-
12
#752940000000
0!
0%
b111 *
0-
02
b111 6
#752950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#752960000000
0!
0%
b0 *
0-
02
b0 6
#752970000000
1!
1%
1-
12
#752980000000
0!
0%
b1 *
0-
02
b1 6
#752990000000
1!
1%
1-
12
#753000000000
0!
0%
b10 *
0-
02
b10 6
#753010000000
1!
1%
1-
12
#753020000000
0!
0%
b11 *
0-
02
b11 6
#753030000000
1!
1%
1-
12
15
#753040000000
0!
0%
b100 *
0-
02
b100 6
#753050000000
1!
1%
1-
12
#753060000000
0!
0%
b101 *
0-
02
b101 6
#753070000000
1!
1%
1-
12
#753080000000
0!
0%
b110 *
0-
02
b110 6
#753090000000
1!
1%
1-
12
#753100000000
0!
0%
b111 *
0-
02
b111 6
#753110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#753120000000
0!
0%
b0 *
0-
02
b0 6
#753130000000
1!
1%
1-
12
#753140000000
0!
0%
b1 *
0-
02
b1 6
#753150000000
1!
1%
1-
12
#753160000000
0!
0%
b10 *
0-
02
b10 6
#753170000000
1!
1%
1-
12
#753180000000
0!
0%
b11 *
0-
02
b11 6
#753190000000
1!
1%
1-
12
15
#753200000000
0!
0%
b100 *
0-
02
b100 6
#753210000000
1!
1%
1-
12
#753220000000
0!
0%
b101 *
0-
02
b101 6
#753230000000
1!
1%
1-
12
#753240000000
0!
0%
b110 *
0-
02
b110 6
#753250000000
1!
1%
1-
12
#753260000000
0!
0%
b111 *
0-
02
b111 6
#753270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#753280000000
0!
0%
b0 *
0-
02
b0 6
#753290000000
1!
1%
1-
12
#753300000000
0!
0%
b1 *
0-
02
b1 6
#753310000000
1!
1%
1-
12
#753320000000
0!
0%
b10 *
0-
02
b10 6
#753330000000
1!
1%
1-
12
#753340000000
0!
0%
b11 *
0-
02
b11 6
#753350000000
1!
1%
1-
12
15
#753360000000
0!
0%
b100 *
0-
02
b100 6
#753370000000
1!
1%
1-
12
#753380000000
0!
0%
b101 *
0-
02
b101 6
#753390000000
1!
1%
1-
12
#753400000000
0!
0%
b110 *
0-
02
b110 6
#753410000000
1!
1%
1-
12
#753420000000
0!
0%
b111 *
0-
02
b111 6
#753430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#753440000000
0!
0%
b0 *
0-
02
b0 6
#753450000000
1!
1%
1-
12
#753460000000
0!
0%
b1 *
0-
02
b1 6
#753470000000
1!
1%
1-
12
#753480000000
0!
0%
b10 *
0-
02
b10 6
#753490000000
1!
1%
1-
12
#753500000000
0!
0%
b11 *
0-
02
b11 6
#753510000000
1!
1%
1-
12
15
#753520000000
0!
0%
b100 *
0-
02
b100 6
#753530000000
1!
1%
1-
12
#753540000000
0!
0%
b101 *
0-
02
b101 6
#753550000000
1!
1%
1-
12
#753560000000
0!
0%
b110 *
0-
02
b110 6
#753570000000
1!
1%
1-
12
#753580000000
0!
0%
b111 *
0-
02
b111 6
#753590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#753600000000
0!
0%
b0 *
0-
02
b0 6
#753610000000
1!
1%
1-
12
#753620000000
0!
0%
b1 *
0-
02
b1 6
#753630000000
1!
1%
1-
12
#753640000000
0!
0%
b10 *
0-
02
b10 6
#753650000000
1!
1%
1-
12
#753660000000
0!
0%
b11 *
0-
02
b11 6
#753670000000
1!
1%
1-
12
15
#753680000000
0!
0%
b100 *
0-
02
b100 6
#753690000000
1!
1%
1-
12
#753700000000
0!
0%
b101 *
0-
02
b101 6
#753710000000
1!
1%
1-
12
#753720000000
0!
0%
b110 *
0-
02
b110 6
#753730000000
1!
1%
1-
12
#753740000000
0!
0%
b111 *
0-
02
b111 6
#753750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#753760000000
0!
0%
b0 *
0-
02
b0 6
#753770000000
1!
1%
1-
12
#753780000000
0!
0%
b1 *
0-
02
b1 6
#753790000000
1!
1%
1-
12
#753800000000
0!
0%
b10 *
0-
02
b10 6
#753810000000
1!
1%
1-
12
#753820000000
0!
0%
b11 *
0-
02
b11 6
#753830000000
1!
1%
1-
12
15
#753840000000
0!
0%
b100 *
0-
02
b100 6
#753850000000
1!
1%
1-
12
#753860000000
0!
0%
b101 *
0-
02
b101 6
#753870000000
1!
1%
1-
12
#753880000000
0!
0%
b110 *
0-
02
b110 6
#753890000000
1!
1%
1-
12
#753900000000
0!
0%
b111 *
0-
02
b111 6
#753910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#753920000000
0!
0%
b0 *
0-
02
b0 6
#753930000000
1!
1%
1-
12
#753940000000
0!
0%
b1 *
0-
02
b1 6
#753950000000
1!
1%
1-
12
#753960000000
0!
0%
b10 *
0-
02
b10 6
#753970000000
1!
1%
1-
12
#753980000000
0!
0%
b11 *
0-
02
b11 6
#753990000000
1!
1%
1-
12
15
#754000000000
0!
0%
b100 *
0-
02
b100 6
#754010000000
1!
1%
1-
12
#754020000000
0!
0%
b101 *
0-
02
b101 6
#754030000000
1!
1%
1-
12
#754040000000
0!
0%
b110 *
0-
02
b110 6
#754050000000
1!
1%
1-
12
#754060000000
0!
0%
b111 *
0-
02
b111 6
#754070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#754080000000
0!
0%
b0 *
0-
02
b0 6
#754090000000
1!
1%
1-
12
#754100000000
0!
0%
b1 *
0-
02
b1 6
#754110000000
1!
1%
1-
12
#754120000000
0!
0%
b10 *
0-
02
b10 6
#754130000000
1!
1%
1-
12
#754140000000
0!
0%
b11 *
0-
02
b11 6
#754150000000
1!
1%
1-
12
15
#754160000000
0!
0%
b100 *
0-
02
b100 6
#754170000000
1!
1%
1-
12
#754180000000
0!
0%
b101 *
0-
02
b101 6
#754190000000
1!
1%
1-
12
#754200000000
0!
0%
b110 *
0-
02
b110 6
#754210000000
1!
1%
1-
12
#754220000000
0!
0%
b111 *
0-
02
b111 6
#754230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#754240000000
0!
0%
b0 *
0-
02
b0 6
#754250000000
1!
1%
1-
12
#754260000000
0!
0%
b1 *
0-
02
b1 6
#754270000000
1!
1%
1-
12
#754280000000
0!
0%
b10 *
0-
02
b10 6
#754290000000
1!
1%
1-
12
#754300000000
0!
0%
b11 *
0-
02
b11 6
#754310000000
1!
1%
1-
12
15
#754320000000
0!
0%
b100 *
0-
02
b100 6
#754330000000
1!
1%
1-
12
#754340000000
0!
0%
b101 *
0-
02
b101 6
#754350000000
1!
1%
1-
12
#754360000000
0!
0%
b110 *
0-
02
b110 6
#754370000000
1!
1%
1-
12
#754380000000
0!
0%
b111 *
0-
02
b111 6
#754390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#754400000000
0!
0%
b0 *
0-
02
b0 6
#754410000000
1!
1%
1-
12
#754420000000
0!
0%
b1 *
0-
02
b1 6
#754430000000
1!
1%
1-
12
#754440000000
0!
0%
b10 *
0-
02
b10 6
#754450000000
1!
1%
1-
12
#754460000000
0!
0%
b11 *
0-
02
b11 6
#754470000000
1!
1%
1-
12
15
#754480000000
0!
0%
b100 *
0-
02
b100 6
#754490000000
1!
1%
1-
12
#754500000000
0!
0%
b101 *
0-
02
b101 6
#754510000000
1!
1%
1-
12
#754520000000
0!
0%
b110 *
0-
02
b110 6
#754530000000
1!
1%
1-
12
#754540000000
0!
0%
b111 *
0-
02
b111 6
#754550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#754560000000
0!
0%
b0 *
0-
02
b0 6
#754570000000
1!
1%
1-
12
#754580000000
0!
0%
b1 *
0-
02
b1 6
#754590000000
1!
1%
1-
12
#754600000000
0!
0%
b10 *
0-
02
b10 6
#754610000000
1!
1%
1-
12
#754620000000
0!
0%
b11 *
0-
02
b11 6
#754630000000
1!
1%
1-
12
15
#754640000000
0!
0%
b100 *
0-
02
b100 6
#754650000000
1!
1%
1-
12
#754660000000
0!
0%
b101 *
0-
02
b101 6
#754670000000
1!
1%
1-
12
#754680000000
0!
0%
b110 *
0-
02
b110 6
#754690000000
1!
1%
1-
12
#754700000000
0!
0%
b111 *
0-
02
b111 6
#754710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#754720000000
0!
0%
b0 *
0-
02
b0 6
#754730000000
1!
1%
1-
12
#754740000000
0!
0%
b1 *
0-
02
b1 6
#754750000000
1!
1%
1-
12
#754760000000
0!
0%
b10 *
0-
02
b10 6
#754770000000
1!
1%
1-
12
#754780000000
0!
0%
b11 *
0-
02
b11 6
#754790000000
1!
1%
1-
12
15
#754800000000
0!
0%
b100 *
0-
02
b100 6
#754810000000
1!
1%
1-
12
#754820000000
0!
0%
b101 *
0-
02
b101 6
#754830000000
1!
1%
1-
12
#754840000000
0!
0%
b110 *
0-
02
b110 6
#754850000000
1!
1%
1-
12
#754860000000
0!
0%
b111 *
0-
02
b111 6
#754870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#754880000000
0!
0%
b0 *
0-
02
b0 6
#754890000000
1!
1%
1-
12
#754900000000
0!
0%
b1 *
0-
02
b1 6
#754910000000
1!
1%
1-
12
#754920000000
0!
0%
b10 *
0-
02
b10 6
#754930000000
1!
1%
1-
12
#754940000000
0!
0%
b11 *
0-
02
b11 6
#754950000000
1!
1%
1-
12
15
#754960000000
0!
0%
b100 *
0-
02
b100 6
#754970000000
1!
1%
1-
12
#754980000000
0!
0%
b101 *
0-
02
b101 6
#754990000000
1!
1%
1-
12
#755000000000
0!
0%
b110 *
0-
02
b110 6
#755010000000
1!
1%
1-
12
#755020000000
0!
0%
b111 *
0-
02
b111 6
#755030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#755040000000
0!
0%
b0 *
0-
02
b0 6
#755050000000
1!
1%
1-
12
#755060000000
0!
0%
b1 *
0-
02
b1 6
#755070000000
1!
1%
1-
12
#755080000000
0!
0%
b10 *
0-
02
b10 6
#755090000000
1!
1%
1-
12
#755100000000
0!
0%
b11 *
0-
02
b11 6
#755110000000
1!
1%
1-
12
15
#755120000000
0!
0%
b100 *
0-
02
b100 6
#755130000000
1!
1%
1-
12
#755140000000
0!
0%
b101 *
0-
02
b101 6
#755150000000
1!
1%
1-
12
#755160000000
0!
0%
b110 *
0-
02
b110 6
#755170000000
1!
1%
1-
12
#755180000000
0!
0%
b111 *
0-
02
b111 6
#755190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#755200000000
0!
0%
b0 *
0-
02
b0 6
#755210000000
1!
1%
1-
12
#755220000000
0!
0%
b1 *
0-
02
b1 6
#755230000000
1!
1%
1-
12
#755240000000
0!
0%
b10 *
0-
02
b10 6
#755250000000
1!
1%
1-
12
#755260000000
0!
0%
b11 *
0-
02
b11 6
#755270000000
1!
1%
1-
12
15
#755280000000
0!
0%
b100 *
0-
02
b100 6
#755290000000
1!
1%
1-
12
#755300000000
0!
0%
b101 *
0-
02
b101 6
#755310000000
1!
1%
1-
12
#755320000000
0!
0%
b110 *
0-
02
b110 6
#755330000000
1!
1%
1-
12
#755340000000
0!
0%
b111 *
0-
02
b111 6
#755350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#755360000000
0!
0%
b0 *
0-
02
b0 6
#755370000000
1!
1%
1-
12
#755380000000
0!
0%
b1 *
0-
02
b1 6
#755390000000
1!
1%
1-
12
#755400000000
0!
0%
b10 *
0-
02
b10 6
#755410000000
1!
1%
1-
12
#755420000000
0!
0%
b11 *
0-
02
b11 6
#755430000000
1!
1%
1-
12
15
#755440000000
0!
0%
b100 *
0-
02
b100 6
#755450000000
1!
1%
1-
12
#755460000000
0!
0%
b101 *
0-
02
b101 6
#755470000000
1!
1%
1-
12
#755480000000
0!
0%
b110 *
0-
02
b110 6
#755490000000
1!
1%
1-
12
#755500000000
0!
0%
b111 *
0-
02
b111 6
#755510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#755520000000
0!
0%
b0 *
0-
02
b0 6
#755530000000
1!
1%
1-
12
#755540000000
0!
0%
b1 *
0-
02
b1 6
#755550000000
1!
1%
1-
12
#755560000000
0!
0%
b10 *
0-
02
b10 6
#755570000000
1!
1%
1-
12
#755580000000
0!
0%
b11 *
0-
02
b11 6
#755590000000
1!
1%
1-
12
15
#755600000000
0!
0%
b100 *
0-
02
b100 6
#755610000000
1!
1%
1-
12
#755620000000
0!
0%
b101 *
0-
02
b101 6
#755630000000
1!
1%
1-
12
#755640000000
0!
0%
b110 *
0-
02
b110 6
#755650000000
1!
1%
1-
12
#755660000000
0!
0%
b111 *
0-
02
b111 6
#755670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#755680000000
0!
0%
b0 *
0-
02
b0 6
#755690000000
1!
1%
1-
12
#755700000000
0!
0%
b1 *
0-
02
b1 6
#755710000000
1!
1%
1-
12
#755720000000
0!
0%
b10 *
0-
02
b10 6
#755730000000
1!
1%
1-
12
#755740000000
0!
0%
b11 *
0-
02
b11 6
#755750000000
1!
1%
1-
12
15
#755760000000
0!
0%
b100 *
0-
02
b100 6
#755770000000
1!
1%
1-
12
#755780000000
0!
0%
b101 *
0-
02
b101 6
#755790000000
1!
1%
1-
12
#755800000000
0!
0%
b110 *
0-
02
b110 6
#755810000000
1!
1%
1-
12
#755820000000
0!
0%
b111 *
0-
02
b111 6
#755830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#755840000000
0!
0%
b0 *
0-
02
b0 6
#755850000000
1!
1%
1-
12
#755860000000
0!
0%
b1 *
0-
02
b1 6
#755870000000
1!
1%
1-
12
#755880000000
0!
0%
b10 *
0-
02
b10 6
#755890000000
1!
1%
1-
12
#755900000000
0!
0%
b11 *
0-
02
b11 6
#755910000000
1!
1%
1-
12
15
#755920000000
0!
0%
b100 *
0-
02
b100 6
#755930000000
1!
1%
1-
12
#755940000000
0!
0%
b101 *
0-
02
b101 6
#755950000000
1!
1%
1-
12
#755960000000
0!
0%
b110 *
0-
02
b110 6
#755970000000
1!
1%
1-
12
#755980000000
0!
0%
b111 *
0-
02
b111 6
#755990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#756000000000
0!
0%
b0 *
0-
02
b0 6
#756010000000
1!
1%
1-
12
#756020000000
0!
0%
b1 *
0-
02
b1 6
#756030000000
1!
1%
1-
12
#756040000000
0!
0%
b10 *
0-
02
b10 6
#756050000000
1!
1%
1-
12
#756060000000
0!
0%
b11 *
0-
02
b11 6
#756070000000
1!
1%
1-
12
15
#756080000000
0!
0%
b100 *
0-
02
b100 6
#756090000000
1!
1%
1-
12
#756100000000
0!
0%
b101 *
0-
02
b101 6
#756110000000
1!
1%
1-
12
#756120000000
0!
0%
b110 *
0-
02
b110 6
#756130000000
1!
1%
1-
12
#756140000000
0!
0%
b111 *
0-
02
b111 6
#756150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#756160000000
0!
0%
b0 *
0-
02
b0 6
#756170000000
1!
1%
1-
12
#756180000000
0!
0%
b1 *
0-
02
b1 6
#756190000000
1!
1%
1-
12
#756200000000
0!
0%
b10 *
0-
02
b10 6
#756210000000
1!
1%
1-
12
#756220000000
0!
0%
b11 *
0-
02
b11 6
#756230000000
1!
1%
1-
12
15
#756240000000
0!
0%
b100 *
0-
02
b100 6
#756250000000
1!
1%
1-
12
#756260000000
0!
0%
b101 *
0-
02
b101 6
#756270000000
1!
1%
1-
12
#756280000000
0!
0%
b110 *
0-
02
b110 6
#756290000000
1!
1%
1-
12
#756300000000
0!
0%
b111 *
0-
02
b111 6
#756310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#756320000000
0!
0%
b0 *
0-
02
b0 6
#756330000000
1!
1%
1-
12
#756340000000
0!
0%
b1 *
0-
02
b1 6
#756350000000
1!
1%
1-
12
#756360000000
0!
0%
b10 *
0-
02
b10 6
#756370000000
1!
1%
1-
12
#756380000000
0!
0%
b11 *
0-
02
b11 6
#756390000000
1!
1%
1-
12
15
#756400000000
0!
0%
b100 *
0-
02
b100 6
#756410000000
1!
1%
1-
12
#756420000000
0!
0%
b101 *
0-
02
b101 6
#756430000000
1!
1%
1-
12
#756440000000
0!
0%
b110 *
0-
02
b110 6
#756450000000
1!
1%
1-
12
#756460000000
0!
0%
b111 *
0-
02
b111 6
#756470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#756480000000
0!
0%
b0 *
0-
02
b0 6
#756490000000
1!
1%
1-
12
#756500000000
0!
0%
b1 *
0-
02
b1 6
#756510000000
1!
1%
1-
12
#756520000000
0!
0%
b10 *
0-
02
b10 6
#756530000000
1!
1%
1-
12
#756540000000
0!
0%
b11 *
0-
02
b11 6
#756550000000
1!
1%
1-
12
15
#756560000000
0!
0%
b100 *
0-
02
b100 6
#756570000000
1!
1%
1-
12
#756580000000
0!
0%
b101 *
0-
02
b101 6
#756590000000
1!
1%
1-
12
#756600000000
0!
0%
b110 *
0-
02
b110 6
#756610000000
1!
1%
1-
12
#756620000000
0!
0%
b111 *
0-
02
b111 6
#756630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#756640000000
0!
0%
b0 *
0-
02
b0 6
#756650000000
1!
1%
1-
12
#756660000000
0!
0%
b1 *
0-
02
b1 6
#756670000000
1!
1%
1-
12
#756680000000
0!
0%
b10 *
0-
02
b10 6
#756690000000
1!
1%
1-
12
#756700000000
0!
0%
b11 *
0-
02
b11 6
#756710000000
1!
1%
1-
12
15
#756720000000
0!
0%
b100 *
0-
02
b100 6
#756730000000
1!
1%
1-
12
#756740000000
0!
0%
b101 *
0-
02
b101 6
#756750000000
1!
1%
1-
12
#756760000000
0!
0%
b110 *
0-
02
b110 6
#756770000000
1!
1%
1-
12
#756780000000
0!
0%
b111 *
0-
02
b111 6
#756790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#756800000000
0!
0%
b0 *
0-
02
b0 6
#756810000000
1!
1%
1-
12
#756820000000
0!
0%
b1 *
0-
02
b1 6
#756830000000
1!
1%
1-
12
#756840000000
0!
0%
b10 *
0-
02
b10 6
#756850000000
1!
1%
1-
12
#756860000000
0!
0%
b11 *
0-
02
b11 6
#756870000000
1!
1%
1-
12
15
#756880000000
0!
0%
b100 *
0-
02
b100 6
#756890000000
1!
1%
1-
12
#756900000000
0!
0%
b101 *
0-
02
b101 6
#756910000000
1!
1%
1-
12
#756920000000
0!
0%
b110 *
0-
02
b110 6
#756930000000
1!
1%
1-
12
#756940000000
0!
0%
b111 *
0-
02
b111 6
#756950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#756960000000
0!
0%
b0 *
0-
02
b0 6
#756970000000
1!
1%
1-
12
#756980000000
0!
0%
b1 *
0-
02
b1 6
#756990000000
1!
1%
1-
12
#757000000000
0!
0%
b10 *
0-
02
b10 6
#757010000000
1!
1%
1-
12
#757020000000
0!
0%
b11 *
0-
02
b11 6
#757030000000
1!
1%
1-
12
15
#757040000000
0!
0%
b100 *
0-
02
b100 6
#757050000000
1!
1%
1-
12
#757060000000
0!
0%
b101 *
0-
02
b101 6
#757070000000
1!
1%
1-
12
#757080000000
0!
0%
b110 *
0-
02
b110 6
#757090000000
1!
1%
1-
12
#757100000000
0!
0%
b111 *
0-
02
b111 6
#757110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#757120000000
0!
0%
b0 *
0-
02
b0 6
#757130000000
1!
1%
1-
12
#757140000000
0!
0%
b1 *
0-
02
b1 6
#757150000000
1!
1%
1-
12
#757160000000
0!
0%
b10 *
0-
02
b10 6
#757170000000
1!
1%
1-
12
#757180000000
0!
0%
b11 *
0-
02
b11 6
#757190000000
1!
1%
1-
12
15
#757200000000
0!
0%
b100 *
0-
02
b100 6
#757210000000
1!
1%
1-
12
#757220000000
0!
0%
b101 *
0-
02
b101 6
#757230000000
1!
1%
1-
12
#757240000000
0!
0%
b110 *
0-
02
b110 6
#757250000000
1!
1%
1-
12
#757260000000
0!
0%
b111 *
0-
02
b111 6
#757270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#757280000000
0!
0%
b0 *
0-
02
b0 6
#757290000000
1!
1%
1-
12
#757300000000
0!
0%
b1 *
0-
02
b1 6
#757310000000
1!
1%
1-
12
#757320000000
0!
0%
b10 *
0-
02
b10 6
#757330000000
1!
1%
1-
12
#757340000000
0!
0%
b11 *
0-
02
b11 6
#757350000000
1!
1%
1-
12
15
#757360000000
0!
0%
b100 *
0-
02
b100 6
#757370000000
1!
1%
1-
12
#757380000000
0!
0%
b101 *
0-
02
b101 6
#757390000000
1!
1%
1-
12
#757400000000
0!
0%
b110 *
0-
02
b110 6
#757410000000
1!
1%
1-
12
#757420000000
0!
0%
b111 *
0-
02
b111 6
#757430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#757440000000
0!
0%
b0 *
0-
02
b0 6
#757450000000
1!
1%
1-
12
#757460000000
0!
0%
b1 *
0-
02
b1 6
#757470000000
1!
1%
1-
12
#757480000000
0!
0%
b10 *
0-
02
b10 6
#757490000000
1!
1%
1-
12
#757500000000
0!
0%
b11 *
0-
02
b11 6
#757510000000
1!
1%
1-
12
15
#757520000000
0!
0%
b100 *
0-
02
b100 6
#757530000000
1!
1%
1-
12
#757540000000
0!
0%
b101 *
0-
02
b101 6
#757550000000
1!
1%
1-
12
#757560000000
0!
0%
b110 *
0-
02
b110 6
#757570000000
1!
1%
1-
12
#757580000000
0!
0%
b111 *
0-
02
b111 6
#757590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#757600000000
0!
0%
b0 *
0-
02
b0 6
#757610000000
1!
1%
1-
12
#757620000000
0!
0%
b1 *
0-
02
b1 6
#757630000000
1!
1%
1-
12
#757640000000
0!
0%
b10 *
0-
02
b10 6
#757650000000
1!
1%
1-
12
#757660000000
0!
0%
b11 *
0-
02
b11 6
#757670000000
1!
1%
1-
12
15
#757680000000
0!
0%
b100 *
0-
02
b100 6
#757690000000
1!
1%
1-
12
#757700000000
0!
0%
b101 *
0-
02
b101 6
#757710000000
1!
1%
1-
12
#757720000000
0!
0%
b110 *
0-
02
b110 6
#757730000000
1!
1%
1-
12
#757740000000
0!
0%
b111 *
0-
02
b111 6
#757750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#757760000000
0!
0%
b0 *
0-
02
b0 6
#757770000000
1!
1%
1-
12
#757780000000
0!
0%
b1 *
0-
02
b1 6
#757790000000
1!
1%
1-
12
#757800000000
0!
0%
b10 *
0-
02
b10 6
#757810000000
1!
1%
1-
12
#757820000000
0!
0%
b11 *
0-
02
b11 6
#757830000000
1!
1%
1-
12
15
#757840000000
0!
0%
b100 *
0-
02
b100 6
#757850000000
1!
1%
1-
12
#757860000000
0!
0%
b101 *
0-
02
b101 6
#757870000000
1!
1%
1-
12
#757880000000
0!
0%
b110 *
0-
02
b110 6
#757890000000
1!
1%
1-
12
#757900000000
0!
0%
b111 *
0-
02
b111 6
#757910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#757920000000
0!
0%
b0 *
0-
02
b0 6
#757930000000
1!
1%
1-
12
#757940000000
0!
0%
b1 *
0-
02
b1 6
#757950000000
1!
1%
1-
12
#757960000000
0!
0%
b10 *
0-
02
b10 6
#757970000000
1!
1%
1-
12
#757980000000
0!
0%
b11 *
0-
02
b11 6
#757990000000
1!
1%
1-
12
15
#758000000000
0!
0%
b100 *
0-
02
b100 6
#758010000000
1!
1%
1-
12
#758020000000
0!
0%
b101 *
0-
02
b101 6
#758030000000
1!
1%
1-
12
#758040000000
0!
0%
b110 *
0-
02
b110 6
#758050000000
1!
1%
1-
12
#758060000000
0!
0%
b111 *
0-
02
b111 6
#758070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#758080000000
0!
0%
b0 *
0-
02
b0 6
#758090000000
1!
1%
1-
12
#758100000000
0!
0%
b1 *
0-
02
b1 6
#758110000000
1!
1%
1-
12
#758120000000
0!
0%
b10 *
0-
02
b10 6
#758130000000
1!
1%
1-
12
#758140000000
0!
0%
b11 *
0-
02
b11 6
#758150000000
1!
1%
1-
12
15
#758160000000
0!
0%
b100 *
0-
02
b100 6
#758170000000
1!
1%
1-
12
#758180000000
0!
0%
b101 *
0-
02
b101 6
#758190000000
1!
1%
1-
12
#758200000000
0!
0%
b110 *
0-
02
b110 6
#758210000000
1!
1%
1-
12
#758220000000
0!
0%
b111 *
0-
02
b111 6
#758230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#758240000000
0!
0%
b0 *
0-
02
b0 6
#758250000000
1!
1%
1-
12
#758260000000
0!
0%
b1 *
0-
02
b1 6
#758270000000
1!
1%
1-
12
#758280000000
0!
0%
b10 *
0-
02
b10 6
#758290000000
1!
1%
1-
12
#758300000000
0!
0%
b11 *
0-
02
b11 6
#758310000000
1!
1%
1-
12
15
#758320000000
0!
0%
b100 *
0-
02
b100 6
#758330000000
1!
1%
1-
12
#758340000000
0!
0%
b101 *
0-
02
b101 6
#758350000000
1!
1%
1-
12
#758360000000
0!
0%
b110 *
0-
02
b110 6
#758370000000
1!
1%
1-
12
#758380000000
0!
0%
b111 *
0-
02
b111 6
#758390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#758400000000
0!
0%
b0 *
0-
02
b0 6
#758410000000
1!
1%
1-
12
#758420000000
0!
0%
b1 *
0-
02
b1 6
#758430000000
1!
1%
1-
12
#758440000000
0!
0%
b10 *
0-
02
b10 6
#758450000000
1!
1%
1-
12
#758460000000
0!
0%
b11 *
0-
02
b11 6
#758470000000
1!
1%
1-
12
15
#758480000000
0!
0%
b100 *
0-
02
b100 6
#758490000000
1!
1%
1-
12
#758500000000
0!
0%
b101 *
0-
02
b101 6
#758510000000
1!
1%
1-
12
#758520000000
0!
0%
b110 *
0-
02
b110 6
#758530000000
1!
1%
1-
12
#758540000000
0!
0%
b111 *
0-
02
b111 6
#758550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#758560000000
0!
0%
b0 *
0-
02
b0 6
#758570000000
1!
1%
1-
12
#758580000000
0!
0%
b1 *
0-
02
b1 6
#758590000000
1!
1%
1-
12
#758600000000
0!
0%
b10 *
0-
02
b10 6
#758610000000
1!
1%
1-
12
#758620000000
0!
0%
b11 *
0-
02
b11 6
#758630000000
1!
1%
1-
12
15
#758640000000
0!
0%
b100 *
0-
02
b100 6
#758650000000
1!
1%
1-
12
#758660000000
0!
0%
b101 *
0-
02
b101 6
#758670000000
1!
1%
1-
12
#758680000000
0!
0%
b110 *
0-
02
b110 6
#758690000000
1!
1%
1-
12
#758700000000
0!
0%
b111 *
0-
02
b111 6
#758710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#758720000000
0!
0%
b0 *
0-
02
b0 6
#758730000000
1!
1%
1-
12
#758740000000
0!
0%
b1 *
0-
02
b1 6
#758750000000
1!
1%
1-
12
#758760000000
0!
0%
b10 *
0-
02
b10 6
#758770000000
1!
1%
1-
12
#758780000000
0!
0%
b11 *
0-
02
b11 6
#758790000000
1!
1%
1-
12
15
#758800000000
0!
0%
b100 *
0-
02
b100 6
#758810000000
1!
1%
1-
12
#758820000000
0!
0%
b101 *
0-
02
b101 6
#758830000000
1!
1%
1-
12
#758840000000
0!
0%
b110 *
0-
02
b110 6
#758850000000
1!
1%
1-
12
#758860000000
0!
0%
b111 *
0-
02
b111 6
#758870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#758880000000
0!
0%
b0 *
0-
02
b0 6
#758890000000
1!
1%
1-
12
#758900000000
0!
0%
b1 *
0-
02
b1 6
#758910000000
1!
1%
1-
12
#758920000000
0!
0%
b10 *
0-
02
b10 6
#758930000000
1!
1%
1-
12
#758940000000
0!
0%
b11 *
0-
02
b11 6
#758950000000
1!
1%
1-
12
15
#758960000000
0!
0%
b100 *
0-
02
b100 6
#758970000000
1!
1%
1-
12
#758980000000
0!
0%
b101 *
0-
02
b101 6
#758990000000
1!
1%
1-
12
#759000000000
0!
0%
b110 *
0-
02
b110 6
#759010000000
1!
1%
1-
12
#759020000000
0!
0%
b111 *
0-
02
b111 6
#759030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#759040000000
0!
0%
b0 *
0-
02
b0 6
#759050000000
1!
1%
1-
12
#759060000000
0!
0%
b1 *
0-
02
b1 6
#759070000000
1!
1%
1-
12
#759080000000
0!
0%
b10 *
0-
02
b10 6
#759090000000
1!
1%
1-
12
#759100000000
0!
0%
b11 *
0-
02
b11 6
#759110000000
1!
1%
1-
12
15
#759120000000
0!
0%
b100 *
0-
02
b100 6
#759130000000
1!
1%
1-
12
#759140000000
0!
0%
b101 *
0-
02
b101 6
#759150000000
1!
1%
1-
12
#759160000000
0!
0%
b110 *
0-
02
b110 6
#759170000000
1!
1%
1-
12
#759180000000
0!
0%
b111 *
0-
02
b111 6
#759190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#759200000000
0!
0%
b0 *
0-
02
b0 6
#759210000000
1!
1%
1-
12
#759220000000
0!
0%
b1 *
0-
02
b1 6
#759230000000
1!
1%
1-
12
#759240000000
0!
0%
b10 *
0-
02
b10 6
#759250000000
1!
1%
1-
12
#759260000000
0!
0%
b11 *
0-
02
b11 6
#759270000000
1!
1%
1-
12
15
#759280000000
0!
0%
b100 *
0-
02
b100 6
#759290000000
1!
1%
1-
12
#759300000000
0!
0%
b101 *
0-
02
b101 6
#759310000000
1!
1%
1-
12
#759320000000
0!
0%
b110 *
0-
02
b110 6
#759330000000
1!
1%
1-
12
#759340000000
0!
0%
b111 *
0-
02
b111 6
#759350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#759360000000
0!
0%
b0 *
0-
02
b0 6
#759370000000
1!
1%
1-
12
#759380000000
0!
0%
b1 *
0-
02
b1 6
#759390000000
1!
1%
1-
12
#759400000000
0!
0%
b10 *
0-
02
b10 6
#759410000000
1!
1%
1-
12
#759420000000
0!
0%
b11 *
0-
02
b11 6
#759430000000
1!
1%
1-
12
15
#759440000000
0!
0%
b100 *
0-
02
b100 6
#759450000000
1!
1%
1-
12
#759460000000
0!
0%
b101 *
0-
02
b101 6
#759470000000
1!
1%
1-
12
#759480000000
0!
0%
b110 *
0-
02
b110 6
#759490000000
1!
1%
1-
12
#759500000000
0!
0%
b111 *
0-
02
b111 6
#759510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#759520000000
0!
0%
b0 *
0-
02
b0 6
#759530000000
1!
1%
1-
12
#759540000000
0!
0%
b1 *
0-
02
b1 6
#759550000000
1!
1%
1-
12
#759560000000
0!
0%
b10 *
0-
02
b10 6
#759570000000
1!
1%
1-
12
#759580000000
0!
0%
b11 *
0-
02
b11 6
#759590000000
1!
1%
1-
12
15
#759600000000
0!
0%
b100 *
0-
02
b100 6
#759610000000
1!
1%
1-
12
#759620000000
0!
0%
b101 *
0-
02
b101 6
#759630000000
1!
1%
1-
12
#759640000000
0!
0%
b110 *
0-
02
b110 6
#759650000000
1!
1%
1-
12
#759660000000
0!
0%
b111 *
0-
02
b111 6
#759670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#759680000000
0!
0%
b0 *
0-
02
b0 6
#759690000000
1!
1%
1-
12
#759700000000
0!
0%
b1 *
0-
02
b1 6
#759710000000
1!
1%
1-
12
#759720000000
0!
0%
b10 *
0-
02
b10 6
#759730000000
1!
1%
1-
12
#759740000000
0!
0%
b11 *
0-
02
b11 6
#759750000000
1!
1%
1-
12
15
#759760000000
0!
0%
b100 *
0-
02
b100 6
#759770000000
1!
1%
1-
12
#759780000000
0!
0%
b101 *
0-
02
b101 6
#759790000000
1!
1%
1-
12
#759800000000
0!
0%
b110 *
0-
02
b110 6
#759810000000
1!
1%
1-
12
#759820000000
0!
0%
b111 *
0-
02
b111 6
#759830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#759840000000
0!
0%
b0 *
0-
02
b0 6
#759850000000
1!
1%
1-
12
#759860000000
0!
0%
b1 *
0-
02
b1 6
#759870000000
1!
1%
1-
12
#759880000000
0!
0%
b10 *
0-
02
b10 6
#759890000000
1!
1%
1-
12
#759900000000
0!
0%
b11 *
0-
02
b11 6
#759910000000
1!
1%
1-
12
15
#759920000000
0!
0%
b100 *
0-
02
b100 6
#759930000000
1!
1%
1-
12
#759940000000
0!
0%
b101 *
0-
02
b101 6
#759950000000
1!
1%
1-
12
#759960000000
0!
0%
b110 *
0-
02
b110 6
#759970000000
1!
1%
1-
12
#759980000000
0!
0%
b111 *
0-
02
b111 6
#759990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#760000000000
0!
0%
b0 *
0-
02
b0 6
#760010000000
1!
1%
1-
12
#760020000000
0!
0%
b1 *
0-
02
b1 6
#760030000000
1!
1%
1-
12
#760040000000
0!
0%
b10 *
0-
02
b10 6
#760050000000
1!
1%
1-
12
#760060000000
0!
0%
b11 *
0-
02
b11 6
#760070000000
1!
1%
1-
12
15
#760080000000
0!
0%
b100 *
0-
02
b100 6
#760090000000
1!
1%
1-
12
#760100000000
0!
0%
b101 *
0-
02
b101 6
#760110000000
1!
1%
1-
12
#760120000000
0!
0%
b110 *
0-
02
b110 6
#760130000000
1!
1%
1-
12
#760140000000
0!
0%
b111 *
0-
02
b111 6
#760150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#760160000000
0!
0%
b0 *
0-
02
b0 6
#760170000000
1!
1%
1-
12
#760180000000
0!
0%
b1 *
0-
02
b1 6
#760190000000
1!
1%
1-
12
#760200000000
0!
0%
b10 *
0-
02
b10 6
#760210000000
1!
1%
1-
12
#760220000000
0!
0%
b11 *
0-
02
b11 6
#760230000000
1!
1%
1-
12
15
#760240000000
0!
0%
b100 *
0-
02
b100 6
#760250000000
1!
1%
1-
12
#760260000000
0!
0%
b101 *
0-
02
b101 6
#760270000000
1!
1%
1-
12
#760280000000
0!
0%
b110 *
0-
02
b110 6
#760290000000
1!
1%
1-
12
#760300000000
0!
0%
b111 *
0-
02
b111 6
#760310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#760320000000
0!
0%
b0 *
0-
02
b0 6
#760330000000
1!
1%
1-
12
#760340000000
0!
0%
b1 *
0-
02
b1 6
#760350000000
1!
1%
1-
12
#760360000000
0!
0%
b10 *
0-
02
b10 6
#760370000000
1!
1%
1-
12
#760380000000
0!
0%
b11 *
0-
02
b11 6
#760390000000
1!
1%
1-
12
15
#760400000000
0!
0%
b100 *
0-
02
b100 6
#760410000000
1!
1%
1-
12
#760420000000
0!
0%
b101 *
0-
02
b101 6
#760430000000
1!
1%
1-
12
#760440000000
0!
0%
b110 *
0-
02
b110 6
#760450000000
1!
1%
1-
12
#760460000000
0!
0%
b111 *
0-
02
b111 6
#760470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#760480000000
0!
0%
b0 *
0-
02
b0 6
#760490000000
1!
1%
1-
12
#760500000000
0!
0%
b1 *
0-
02
b1 6
#760510000000
1!
1%
1-
12
#760520000000
0!
0%
b10 *
0-
02
b10 6
#760530000000
1!
1%
1-
12
#760540000000
0!
0%
b11 *
0-
02
b11 6
#760550000000
1!
1%
1-
12
15
#760560000000
0!
0%
b100 *
0-
02
b100 6
#760570000000
1!
1%
1-
12
#760580000000
0!
0%
b101 *
0-
02
b101 6
#760590000000
1!
1%
1-
12
#760600000000
0!
0%
b110 *
0-
02
b110 6
#760610000000
1!
1%
1-
12
#760620000000
0!
0%
b111 *
0-
02
b111 6
#760630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#760640000000
0!
0%
b0 *
0-
02
b0 6
#760650000000
1!
1%
1-
12
#760660000000
0!
0%
b1 *
0-
02
b1 6
#760670000000
1!
1%
1-
12
#760680000000
0!
0%
b10 *
0-
02
b10 6
#760690000000
1!
1%
1-
12
#760700000000
0!
0%
b11 *
0-
02
b11 6
#760710000000
1!
1%
1-
12
15
#760720000000
0!
0%
b100 *
0-
02
b100 6
#760730000000
1!
1%
1-
12
#760740000000
0!
0%
b101 *
0-
02
b101 6
#760750000000
1!
1%
1-
12
#760760000000
0!
0%
b110 *
0-
02
b110 6
#760770000000
1!
1%
1-
12
#760780000000
0!
0%
b111 *
0-
02
b111 6
#760790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#760800000000
0!
0%
b0 *
0-
02
b0 6
#760810000000
1!
1%
1-
12
#760820000000
0!
0%
b1 *
0-
02
b1 6
#760830000000
1!
1%
1-
12
#760840000000
0!
0%
b10 *
0-
02
b10 6
#760850000000
1!
1%
1-
12
#760860000000
0!
0%
b11 *
0-
02
b11 6
#760870000000
1!
1%
1-
12
15
#760880000000
0!
0%
b100 *
0-
02
b100 6
#760890000000
1!
1%
1-
12
#760900000000
0!
0%
b101 *
0-
02
b101 6
#760910000000
1!
1%
1-
12
#760920000000
0!
0%
b110 *
0-
02
b110 6
#760930000000
1!
1%
1-
12
#760940000000
0!
0%
b111 *
0-
02
b111 6
#760950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#760960000000
0!
0%
b0 *
0-
02
b0 6
#760970000000
1!
1%
1-
12
#760980000000
0!
0%
b1 *
0-
02
b1 6
#760990000000
1!
1%
1-
12
#761000000000
0!
0%
b10 *
0-
02
b10 6
#761010000000
1!
1%
1-
12
#761020000000
0!
0%
b11 *
0-
02
b11 6
#761030000000
1!
1%
1-
12
15
#761040000000
0!
0%
b100 *
0-
02
b100 6
#761050000000
1!
1%
1-
12
#761060000000
0!
0%
b101 *
0-
02
b101 6
#761070000000
1!
1%
1-
12
#761080000000
0!
0%
b110 *
0-
02
b110 6
#761090000000
1!
1%
1-
12
#761100000000
0!
0%
b111 *
0-
02
b111 6
#761110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#761120000000
0!
0%
b0 *
0-
02
b0 6
#761130000000
1!
1%
1-
12
#761140000000
0!
0%
b1 *
0-
02
b1 6
#761150000000
1!
1%
1-
12
#761160000000
0!
0%
b10 *
0-
02
b10 6
#761170000000
1!
1%
1-
12
#761180000000
0!
0%
b11 *
0-
02
b11 6
#761190000000
1!
1%
1-
12
15
#761200000000
0!
0%
b100 *
0-
02
b100 6
#761210000000
1!
1%
1-
12
#761220000000
0!
0%
b101 *
0-
02
b101 6
#761230000000
1!
1%
1-
12
#761240000000
0!
0%
b110 *
0-
02
b110 6
#761250000000
1!
1%
1-
12
#761260000000
0!
0%
b111 *
0-
02
b111 6
#761270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#761280000000
0!
0%
b0 *
0-
02
b0 6
#761290000000
1!
1%
1-
12
#761300000000
0!
0%
b1 *
0-
02
b1 6
#761310000000
1!
1%
1-
12
#761320000000
0!
0%
b10 *
0-
02
b10 6
#761330000000
1!
1%
1-
12
#761340000000
0!
0%
b11 *
0-
02
b11 6
#761350000000
1!
1%
1-
12
15
#761360000000
0!
0%
b100 *
0-
02
b100 6
#761370000000
1!
1%
1-
12
#761380000000
0!
0%
b101 *
0-
02
b101 6
#761390000000
1!
1%
1-
12
#761400000000
0!
0%
b110 *
0-
02
b110 6
#761410000000
1!
1%
1-
12
#761420000000
0!
0%
b111 *
0-
02
b111 6
#761430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#761440000000
0!
0%
b0 *
0-
02
b0 6
#761450000000
1!
1%
1-
12
#761460000000
0!
0%
b1 *
0-
02
b1 6
#761470000000
1!
1%
1-
12
#761480000000
0!
0%
b10 *
0-
02
b10 6
#761490000000
1!
1%
1-
12
#761500000000
0!
0%
b11 *
0-
02
b11 6
#761510000000
1!
1%
1-
12
15
#761520000000
0!
0%
b100 *
0-
02
b100 6
#761530000000
1!
1%
1-
12
#761540000000
0!
0%
b101 *
0-
02
b101 6
#761550000000
1!
1%
1-
12
#761560000000
0!
0%
b110 *
0-
02
b110 6
#761570000000
1!
1%
1-
12
#761580000000
0!
0%
b111 *
0-
02
b111 6
#761590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#761600000000
0!
0%
b0 *
0-
02
b0 6
#761610000000
1!
1%
1-
12
#761620000000
0!
0%
b1 *
0-
02
b1 6
#761630000000
1!
1%
1-
12
#761640000000
0!
0%
b10 *
0-
02
b10 6
#761650000000
1!
1%
1-
12
#761660000000
0!
0%
b11 *
0-
02
b11 6
#761670000000
1!
1%
1-
12
15
#761680000000
0!
0%
b100 *
0-
02
b100 6
#761690000000
1!
1%
1-
12
#761700000000
0!
0%
b101 *
0-
02
b101 6
#761710000000
1!
1%
1-
12
#761720000000
0!
0%
b110 *
0-
02
b110 6
#761730000000
1!
1%
1-
12
#761740000000
0!
0%
b111 *
0-
02
b111 6
#761750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#761760000000
0!
0%
b0 *
0-
02
b0 6
#761770000000
1!
1%
1-
12
#761780000000
0!
0%
b1 *
0-
02
b1 6
#761790000000
1!
1%
1-
12
#761800000000
0!
0%
b10 *
0-
02
b10 6
#761810000000
1!
1%
1-
12
#761820000000
0!
0%
b11 *
0-
02
b11 6
#761830000000
1!
1%
1-
12
15
#761840000000
0!
0%
b100 *
0-
02
b100 6
#761850000000
1!
1%
1-
12
#761860000000
0!
0%
b101 *
0-
02
b101 6
#761870000000
1!
1%
1-
12
#761880000000
0!
0%
b110 *
0-
02
b110 6
#761890000000
1!
1%
1-
12
#761900000000
0!
0%
b111 *
0-
02
b111 6
#761910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#761920000000
0!
0%
b0 *
0-
02
b0 6
#761930000000
1!
1%
1-
12
#761940000000
0!
0%
b1 *
0-
02
b1 6
#761950000000
1!
1%
1-
12
#761960000000
0!
0%
b10 *
0-
02
b10 6
#761970000000
1!
1%
1-
12
#761980000000
0!
0%
b11 *
0-
02
b11 6
#761990000000
1!
1%
1-
12
15
#762000000000
0!
0%
b100 *
0-
02
b100 6
#762010000000
1!
1%
1-
12
#762020000000
0!
0%
b101 *
0-
02
b101 6
#762030000000
1!
1%
1-
12
#762040000000
0!
0%
b110 *
0-
02
b110 6
#762050000000
1!
1%
1-
12
#762060000000
0!
0%
b111 *
0-
02
b111 6
#762070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#762080000000
0!
0%
b0 *
0-
02
b0 6
#762090000000
1!
1%
1-
12
#762100000000
0!
0%
b1 *
0-
02
b1 6
#762110000000
1!
1%
1-
12
#762120000000
0!
0%
b10 *
0-
02
b10 6
#762130000000
1!
1%
1-
12
#762140000000
0!
0%
b11 *
0-
02
b11 6
#762150000000
1!
1%
1-
12
15
#762160000000
0!
0%
b100 *
0-
02
b100 6
#762170000000
1!
1%
1-
12
#762180000000
0!
0%
b101 *
0-
02
b101 6
#762190000000
1!
1%
1-
12
#762200000000
0!
0%
b110 *
0-
02
b110 6
#762210000000
1!
1%
1-
12
#762220000000
0!
0%
b111 *
0-
02
b111 6
#762230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#762240000000
0!
0%
b0 *
0-
02
b0 6
#762250000000
1!
1%
1-
12
#762260000000
0!
0%
b1 *
0-
02
b1 6
#762270000000
1!
1%
1-
12
#762280000000
0!
0%
b10 *
0-
02
b10 6
#762290000000
1!
1%
1-
12
#762300000000
0!
0%
b11 *
0-
02
b11 6
#762310000000
1!
1%
1-
12
15
#762320000000
0!
0%
b100 *
0-
02
b100 6
#762330000000
1!
1%
1-
12
#762340000000
0!
0%
b101 *
0-
02
b101 6
#762350000000
1!
1%
1-
12
#762360000000
0!
0%
b110 *
0-
02
b110 6
#762370000000
1!
1%
1-
12
#762380000000
0!
0%
b111 *
0-
02
b111 6
#762390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#762400000000
0!
0%
b0 *
0-
02
b0 6
#762410000000
1!
1%
1-
12
#762420000000
0!
0%
b1 *
0-
02
b1 6
#762430000000
1!
1%
1-
12
#762440000000
0!
0%
b10 *
0-
02
b10 6
#762450000000
1!
1%
1-
12
#762460000000
0!
0%
b11 *
0-
02
b11 6
#762470000000
1!
1%
1-
12
15
#762480000000
0!
0%
b100 *
0-
02
b100 6
#762490000000
1!
1%
1-
12
#762500000000
0!
0%
b101 *
0-
02
b101 6
#762510000000
1!
1%
1-
12
#762520000000
0!
0%
b110 *
0-
02
b110 6
#762530000000
1!
1%
1-
12
#762540000000
0!
0%
b111 *
0-
02
b111 6
#762550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#762560000000
0!
0%
b0 *
0-
02
b0 6
#762570000000
1!
1%
1-
12
#762580000000
0!
0%
b1 *
0-
02
b1 6
#762590000000
1!
1%
1-
12
#762600000000
0!
0%
b10 *
0-
02
b10 6
#762610000000
1!
1%
1-
12
#762620000000
0!
0%
b11 *
0-
02
b11 6
#762630000000
1!
1%
1-
12
15
#762640000000
0!
0%
b100 *
0-
02
b100 6
#762650000000
1!
1%
1-
12
#762660000000
0!
0%
b101 *
0-
02
b101 6
#762670000000
1!
1%
1-
12
#762680000000
0!
0%
b110 *
0-
02
b110 6
#762690000000
1!
1%
1-
12
#762700000000
0!
0%
b111 *
0-
02
b111 6
#762710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#762720000000
0!
0%
b0 *
0-
02
b0 6
#762730000000
1!
1%
1-
12
#762740000000
0!
0%
b1 *
0-
02
b1 6
#762750000000
1!
1%
1-
12
#762760000000
0!
0%
b10 *
0-
02
b10 6
#762770000000
1!
1%
1-
12
#762780000000
0!
0%
b11 *
0-
02
b11 6
#762790000000
1!
1%
1-
12
15
#762800000000
0!
0%
b100 *
0-
02
b100 6
#762810000000
1!
1%
1-
12
#762820000000
0!
0%
b101 *
0-
02
b101 6
#762830000000
1!
1%
1-
12
#762840000000
0!
0%
b110 *
0-
02
b110 6
#762850000000
1!
1%
1-
12
#762860000000
0!
0%
b111 *
0-
02
b111 6
#762870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#762880000000
0!
0%
b0 *
0-
02
b0 6
#762890000000
1!
1%
1-
12
#762900000000
0!
0%
b1 *
0-
02
b1 6
#762910000000
1!
1%
1-
12
#762920000000
0!
0%
b10 *
0-
02
b10 6
#762930000000
1!
1%
1-
12
#762940000000
0!
0%
b11 *
0-
02
b11 6
#762950000000
1!
1%
1-
12
15
#762960000000
0!
0%
b100 *
0-
02
b100 6
#762970000000
1!
1%
1-
12
#762980000000
0!
0%
b101 *
0-
02
b101 6
#762990000000
1!
1%
1-
12
#763000000000
0!
0%
b110 *
0-
02
b110 6
#763010000000
1!
1%
1-
12
#763020000000
0!
0%
b111 *
0-
02
b111 6
#763030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#763040000000
0!
0%
b0 *
0-
02
b0 6
#763050000000
1!
1%
1-
12
#763060000000
0!
0%
b1 *
0-
02
b1 6
#763070000000
1!
1%
1-
12
#763080000000
0!
0%
b10 *
0-
02
b10 6
#763090000000
1!
1%
1-
12
#763100000000
0!
0%
b11 *
0-
02
b11 6
#763110000000
1!
1%
1-
12
15
#763120000000
0!
0%
b100 *
0-
02
b100 6
#763130000000
1!
1%
1-
12
#763140000000
0!
0%
b101 *
0-
02
b101 6
#763150000000
1!
1%
1-
12
#763160000000
0!
0%
b110 *
0-
02
b110 6
#763170000000
1!
1%
1-
12
#763180000000
0!
0%
b111 *
0-
02
b111 6
#763190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#763200000000
0!
0%
b0 *
0-
02
b0 6
#763210000000
1!
1%
1-
12
#763220000000
0!
0%
b1 *
0-
02
b1 6
#763230000000
1!
1%
1-
12
#763240000000
0!
0%
b10 *
0-
02
b10 6
#763250000000
1!
1%
1-
12
#763260000000
0!
0%
b11 *
0-
02
b11 6
#763270000000
1!
1%
1-
12
15
#763280000000
0!
0%
b100 *
0-
02
b100 6
#763290000000
1!
1%
1-
12
#763300000000
0!
0%
b101 *
0-
02
b101 6
#763310000000
1!
1%
1-
12
#763320000000
0!
0%
b110 *
0-
02
b110 6
#763330000000
1!
1%
1-
12
#763340000000
0!
0%
b111 *
0-
02
b111 6
#763350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#763360000000
0!
0%
b0 *
0-
02
b0 6
#763370000000
1!
1%
1-
12
#763380000000
0!
0%
b1 *
0-
02
b1 6
#763390000000
1!
1%
1-
12
#763400000000
0!
0%
b10 *
0-
02
b10 6
#763410000000
1!
1%
1-
12
#763420000000
0!
0%
b11 *
0-
02
b11 6
#763430000000
1!
1%
1-
12
15
#763440000000
0!
0%
b100 *
0-
02
b100 6
#763450000000
1!
1%
1-
12
#763460000000
0!
0%
b101 *
0-
02
b101 6
#763470000000
1!
1%
1-
12
#763480000000
0!
0%
b110 *
0-
02
b110 6
#763490000000
1!
1%
1-
12
#763500000000
0!
0%
b111 *
0-
02
b111 6
#763510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#763520000000
0!
0%
b0 *
0-
02
b0 6
#763530000000
1!
1%
1-
12
#763540000000
0!
0%
b1 *
0-
02
b1 6
#763550000000
1!
1%
1-
12
#763560000000
0!
0%
b10 *
0-
02
b10 6
#763570000000
1!
1%
1-
12
#763580000000
0!
0%
b11 *
0-
02
b11 6
#763590000000
1!
1%
1-
12
15
#763600000000
0!
0%
b100 *
0-
02
b100 6
#763610000000
1!
1%
1-
12
#763620000000
0!
0%
b101 *
0-
02
b101 6
#763630000000
1!
1%
1-
12
#763640000000
0!
0%
b110 *
0-
02
b110 6
#763650000000
1!
1%
1-
12
#763660000000
0!
0%
b111 *
0-
02
b111 6
#763670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#763680000000
0!
0%
b0 *
0-
02
b0 6
#763690000000
1!
1%
1-
12
#763700000000
0!
0%
b1 *
0-
02
b1 6
#763710000000
1!
1%
1-
12
#763720000000
0!
0%
b10 *
0-
02
b10 6
#763730000000
1!
1%
1-
12
#763740000000
0!
0%
b11 *
0-
02
b11 6
#763750000000
1!
1%
1-
12
15
#763760000000
0!
0%
b100 *
0-
02
b100 6
#763770000000
1!
1%
1-
12
#763780000000
0!
0%
b101 *
0-
02
b101 6
#763790000000
1!
1%
1-
12
#763800000000
0!
0%
b110 *
0-
02
b110 6
#763810000000
1!
1%
1-
12
#763820000000
0!
0%
b111 *
0-
02
b111 6
#763830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#763840000000
0!
0%
b0 *
0-
02
b0 6
#763850000000
1!
1%
1-
12
#763860000000
0!
0%
b1 *
0-
02
b1 6
#763870000000
1!
1%
1-
12
#763880000000
0!
0%
b10 *
0-
02
b10 6
#763890000000
1!
1%
1-
12
#763900000000
0!
0%
b11 *
0-
02
b11 6
#763910000000
1!
1%
1-
12
15
#763920000000
0!
0%
b100 *
0-
02
b100 6
#763930000000
1!
1%
1-
12
#763940000000
0!
0%
b101 *
0-
02
b101 6
#763950000000
1!
1%
1-
12
#763960000000
0!
0%
b110 *
0-
02
b110 6
#763970000000
1!
1%
1-
12
#763980000000
0!
0%
b111 *
0-
02
b111 6
#763990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#764000000000
0!
0%
b0 *
0-
02
b0 6
#764010000000
1!
1%
1-
12
#764020000000
0!
0%
b1 *
0-
02
b1 6
#764030000000
1!
1%
1-
12
#764040000000
0!
0%
b10 *
0-
02
b10 6
#764050000000
1!
1%
1-
12
#764060000000
0!
0%
b11 *
0-
02
b11 6
#764070000000
1!
1%
1-
12
15
#764080000000
0!
0%
b100 *
0-
02
b100 6
#764090000000
1!
1%
1-
12
#764100000000
0!
0%
b101 *
0-
02
b101 6
#764110000000
1!
1%
1-
12
#764120000000
0!
0%
b110 *
0-
02
b110 6
#764130000000
1!
1%
1-
12
#764140000000
0!
0%
b111 *
0-
02
b111 6
#764150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#764160000000
0!
0%
b0 *
0-
02
b0 6
#764170000000
1!
1%
1-
12
#764180000000
0!
0%
b1 *
0-
02
b1 6
#764190000000
1!
1%
1-
12
#764200000000
0!
0%
b10 *
0-
02
b10 6
#764210000000
1!
1%
1-
12
#764220000000
0!
0%
b11 *
0-
02
b11 6
#764230000000
1!
1%
1-
12
15
#764240000000
0!
0%
b100 *
0-
02
b100 6
#764250000000
1!
1%
1-
12
#764260000000
0!
0%
b101 *
0-
02
b101 6
#764270000000
1!
1%
1-
12
#764280000000
0!
0%
b110 *
0-
02
b110 6
#764290000000
1!
1%
1-
12
#764300000000
0!
0%
b111 *
0-
02
b111 6
#764310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#764320000000
0!
0%
b0 *
0-
02
b0 6
#764330000000
1!
1%
1-
12
#764340000000
0!
0%
b1 *
0-
02
b1 6
#764350000000
1!
1%
1-
12
#764360000000
0!
0%
b10 *
0-
02
b10 6
#764370000000
1!
1%
1-
12
#764380000000
0!
0%
b11 *
0-
02
b11 6
#764390000000
1!
1%
1-
12
15
#764400000000
0!
0%
b100 *
0-
02
b100 6
#764410000000
1!
1%
1-
12
#764420000000
0!
0%
b101 *
0-
02
b101 6
#764430000000
1!
1%
1-
12
#764440000000
0!
0%
b110 *
0-
02
b110 6
#764450000000
1!
1%
1-
12
#764460000000
0!
0%
b111 *
0-
02
b111 6
#764470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#764480000000
0!
0%
b0 *
0-
02
b0 6
#764490000000
1!
1%
1-
12
#764500000000
0!
0%
b1 *
0-
02
b1 6
#764510000000
1!
1%
1-
12
#764520000000
0!
0%
b10 *
0-
02
b10 6
#764530000000
1!
1%
1-
12
#764540000000
0!
0%
b11 *
0-
02
b11 6
#764550000000
1!
1%
1-
12
15
#764560000000
0!
0%
b100 *
0-
02
b100 6
#764570000000
1!
1%
1-
12
#764580000000
0!
0%
b101 *
0-
02
b101 6
#764590000000
1!
1%
1-
12
#764600000000
0!
0%
b110 *
0-
02
b110 6
#764610000000
1!
1%
1-
12
#764620000000
0!
0%
b111 *
0-
02
b111 6
#764630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#764640000000
0!
0%
b0 *
0-
02
b0 6
#764650000000
1!
1%
1-
12
#764660000000
0!
0%
b1 *
0-
02
b1 6
#764670000000
1!
1%
1-
12
#764680000000
0!
0%
b10 *
0-
02
b10 6
#764690000000
1!
1%
1-
12
#764700000000
0!
0%
b11 *
0-
02
b11 6
#764710000000
1!
1%
1-
12
15
#764720000000
0!
0%
b100 *
0-
02
b100 6
#764730000000
1!
1%
1-
12
#764740000000
0!
0%
b101 *
0-
02
b101 6
#764750000000
1!
1%
1-
12
#764760000000
0!
0%
b110 *
0-
02
b110 6
#764770000000
1!
1%
1-
12
#764780000000
0!
0%
b111 *
0-
02
b111 6
#764790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#764800000000
0!
0%
b0 *
0-
02
b0 6
#764810000000
1!
1%
1-
12
#764820000000
0!
0%
b1 *
0-
02
b1 6
#764830000000
1!
1%
1-
12
#764840000000
0!
0%
b10 *
0-
02
b10 6
#764850000000
1!
1%
1-
12
#764860000000
0!
0%
b11 *
0-
02
b11 6
#764870000000
1!
1%
1-
12
15
#764880000000
0!
0%
b100 *
0-
02
b100 6
#764890000000
1!
1%
1-
12
#764900000000
0!
0%
b101 *
0-
02
b101 6
#764910000000
1!
1%
1-
12
#764920000000
0!
0%
b110 *
0-
02
b110 6
#764930000000
1!
1%
1-
12
#764940000000
0!
0%
b111 *
0-
02
b111 6
#764950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#764960000000
0!
0%
b0 *
0-
02
b0 6
#764970000000
1!
1%
1-
12
#764980000000
0!
0%
b1 *
0-
02
b1 6
#764990000000
1!
1%
1-
12
#765000000000
0!
0%
b10 *
0-
02
b10 6
#765010000000
1!
1%
1-
12
#765020000000
0!
0%
b11 *
0-
02
b11 6
#765030000000
1!
1%
1-
12
15
#765040000000
0!
0%
b100 *
0-
02
b100 6
#765050000000
1!
1%
1-
12
#765060000000
0!
0%
b101 *
0-
02
b101 6
#765070000000
1!
1%
1-
12
#765080000000
0!
0%
b110 *
0-
02
b110 6
#765090000000
1!
1%
1-
12
#765100000000
0!
0%
b111 *
0-
02
b111 6
#765110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#765120000000
0!
0%
b0 *
0-
02
b0 6
#765130000000
1!
1%
1-
12
#765140000000
0!
0%
b1 *
0-
02
b1 6
#765150000000
1!
1%
1-
12
#765160000000
0!
0%
b10 *
0-
02
b10 6
#765170000000
1!
1%
1-
12
#765180000000
0!
0%
b11 *
0-
02
b11 6
#765190000000
1!
1%
1-
12
15
#765200000000
0!
0%
b100 *
0-
02
b100 6
#765210000000
1!
1%
1-
12
#765220000000
0!
0%
b101 *
0-
02
b101 6
#765230000000
1!
1%
1-
12
#765240000000
0!
0%
b110 *
0-
02
b110 6
#765250000000
1!
1%
1-
12
#765260000000
0!
0%
b111 *
0-
02
b111 6
#765270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#765280000000
0!
0%
b0 *
0-
02
b0 6
#765290000000
1!
1%
1-
12
#765300000000
0!
0%
b1 *
0-
02
b1 6
#765310000000
1!
1%
1-
12
#765320000000
0!
0%
b10 *
0-
02
b10 6
#765330000000
1!
1%
1-
12
#765340000000
0!
0%
b11 *
0-
02
b11 6
#765350000000
1!
1%
1-
12
15
#765360000000
0!
0%
b100 *
0-
02
b100 6
#765370000000
1!
1%
1-
12
#765380000000
0!
0%
b101 *
0-
02
b101 6
#765390000000
1!
1%
1-
12
#765400000000
0!
0%
b110 *
0-
02
b110 6
#765410000000
1!
1%
1-
12
#765420000000
0!
0%
b111 *
0-
02
b111 6
#765430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#765440000000
0!
0%
b0 *
0-
02
b0 6
#765450000000
1!
1%
1-
12
#765460000000
0!
0%
b1 *
0-
02
b1 6
#765470000000
1!
1%
1-
12
#765480000000
0!
0%
b10 *
0-
02
b10 6
#765490000000
1!
1%
1-
12
#765500000000
0!
0%
b11 *
0-
02
b11 6
#765510000000
1!
1%
1-
12
15
#765520000000
0!
0%
b100 *
0-
02
b100 6
#765530000000
1!
1%
1-
12
#765540000000
0!
0%
b101 *
0-
02
b101 6
#765550000000
1!
1%
1-
12
#765560000000
0!
0%
b110 *
0-
02
b110 6
#765570000000
1!
1%
1-
12
#765580000000
0!
0%
b111 *
0-
02
b111 6
#765590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#765600000000
0!
0%
b0 *
0-
02
b0 6
#765610000000
1!
1%
1-
12
#765620000000
0!
0%
b1 *
0-
02
b1 6
#765630000000
1!
1%
1-
12
#765640000000
0!
0%
b10 *
0-
02
b10 6
#765650000000
1!
1%
1-
12
#765660000000
0!
0%
b11 *
0-
02
b11 6
#765670000000
1!
1%
1-
12
15
#765680000000
0!
0%
b100 *
0-
02
b100 6
#765690000000
1!
1%
1-
12
#765700000000
0!
0%
b101 *
0-
02
b101 6
#765710000000
1!
1%
1-
12
#765720000000
0!
0%
b110 *
0-
02
b110 6
#765730000000
1!
1%
1-
12
#765740000000
0!
0%
b111 *
0-
02
b111 6
#765750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#765760000000
0!
0%
b0 *
0-
02
b0 6
#765770000000
1!
1%
1-
12
#765780000000
0!
0%
b1 *
0-
02
b1 6
#765790000000
1!
1%
1-
12
#765800000000
0!
0%
b10 *
0-
02
b10 6
#765810000000
1!
1%
1-
12
#765820000000
0!
0%
b11 *
0-
02
b11 6
#765830000000
1!
1%
1-
12
15
#765840000000
0!
0%
b100 *
0-
02
b100 6
#765850000000
1!
1%
1-
12
#765860000000
0!
0%
b101 *
0-
02
b101 6
#765870000000
1!
1%
1-
12
#765880000000
0!
0%
b110 *
0-
02
b110 6
#765890000000
1!
1%
1-
12
#765900000000
0!
0%
b111 *
0-
02
b111 6
#765910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#765920000000
0!
0%
b0 *
0-
02
b0 6
#765930000000
1!
1%
1-
12
#765940000000
0!
0%
b1 *
0-
02
b1 6
#765950000000
1!
1%
1-
12
#765960000000
0!
0%
b10 *
0-
02
b10 6
#765970000000
1!
1%
1-
12
#765980000000
0!
0%
b11 *
0-
02
b11 6
#765990000000
1!
1%
1-
12
15
#766000000000
0!
0%
b100 *
0-
02
b100 6
#766010000000
1!
1%
1-
12
#766020000000
0!
0%
b101 *
0-
02
b101 6
#766030000000
1!
1%
1-
12
#766040000000
0!
0%
b110 *
0-
02
b110 6
#766050000000
1!
1%
1-
12
#766060000000
0!
0%
b111 *
0-
02
b111 6
#766070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#766080000000
0!
0%
b0 *
0-
02
b0 6
#766090000000
1!
1%
1-
12
#766100000000
0!
0%
b1 *
0-
02
b1 6
#766110000000
1!
1%
1-
12
#766120000000
0!
0%
b10 *
0-
02
b10 6
#766130000000
1!
1%
1-
12
#766140000000
0!
0%
b11 *
0-
02
b11 6
#766150000000
1!
1%
1-
12
15
#766160000000
0!
0%
b100 *
0-
02
b100 6
#766170000000
1!
1%
1-
12
#766180000000
0!
0%
b101 *
0-
02
b101 6
#766190000000
1!
1%
1-
12
#766200000000
0!
0%
b110 *
0-
02
b110 6
#766210000000
1!
1%
1-
12
#766220000000
0!
0%
b111 *
0-
02
b111 6
#766230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#766240000000
0!
0%
b0 *
0-
02
b0 6
#766250000000
1!
1%
1-
12
#766260000000
0!
0%
b1 *
0-
02
b1 6
#766270000000
1!
1%
1-
12
#766280000000
0!
0%
b10 *
0-
02
b10 6
#766290000000
1!
1%
1-
12
#766300000000
0!
0%
b11 *
0-
02
b11 6
#766310000000
1!
1%
1-
12
15
#766320000000
0!
0%
b100 *
0-
02
b100 6
#766330000000
1!
1%
1-
12
#766340000000
0!
0%
b101 *
0-
02
b101 6
#766350000000
1!
1%
1-
12
#766360000000
0!
0%
b110 *
0-
02
b110 6
#766370000000
1!
1%
1-
12
#766380000000
0!
0%
b111 *
0-
02
b111 6
#766390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#766400000000
0!
0%
b0 *
0-
02
b0 6
#766410000000
1!
1%
1-
12
#766420000000
0!
0%
b1 *
0-
02
b1 6
#766430000000
1!
1%
1-
12
#766440000000
0!
0%
b10 *
0-
02
b10 6
#766450000000
1!
1%
1-
12
#766460000000
0!
0%
b11 *
0-
02
b11 6
#766470000000
1!
1%
1-
12
15
#766480000000
0!
0%
b100 *
0-
02
b100 6
#766490000000
1!
1%
1-
12
#766500000000
0!
0%
b101 *
0-
02
b101 6
#766510000000
1!
1%
1-
12
#766520000000
0!
0%
b110 *
0-
02
b110 6
#766530000000
1!
1%
1-
12
#766540000000
0!
0%
b111 *
0-
02
b111 6
#766550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#766560000000
0!
0%
b0 *
0-
02
b0 6
#766570000000
1!
1%
1-
12
#766580000000
0!
0%
b1 *
0-
02
b1 6
#766590000000
1!
1%
1-
12
#766600000000
0!
0%
b10 *
0-
02
b10 6
#766610000000
1!
1%
1-
12
#766620000000
0!
0%
b11 *
0-
02
b11 6
#766630000000
1!
1%
1-
12
15
#766640000000
0!
0%
b100 *
0-
02
b100 6
#766650000000
1!
1%
1-
12
#766660000000
0!
0%
b101 *
0-
02
b101 6
#766670000000
1!
1%
1-
12
#766680000000
0!
0%
b110 *
0-
02
b110 6
#766690000000
1!
1%
1-
12
#766700000000
0!
0%
b111 *
0-
02
b111 6
#766710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#766720000000
0!
0%
b0 *
0-
02
b0 6
#766730000000
1!
1%
1-
12
#766740000000
0!
0%
b1 *
0-
02
b1 6
#766750000000
1!
1%
1-
12
#766760000000
0!
0%
b10 *
0-
02
b10 6
#766770000000
1!
1%
1-
12
#766780000000
0!
0%
b11 *
0-
02
b11 6
#766790000000
1!
1%
1-
12
15
#766800000000
0!
0%
b100 *
0-
02
b100 6
#766810000000
1!
1%
1-
12
#766820000000
0!
0%
b101 *
0-
02
b101 6
#766830000000
1!
1%
1-
12
#766840000000
0!
0%
b110 *
0-
02
b110 6
#766850000000
1!
1%
1-
12
#766860000000
0!
0%
b111 *
0-
02
b111 6
#766870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#766880000000
0!
0%
b0 *
0-
02
b0 6
#766890000000
1!
1%
1-
12
#766900000000
0!
0%
b1 *
0-
02
b1 6
#766910000000
1!
1%
1-
12
#766920000000
0!
0%
b10 *
0-
02
b10 6
#766930000000
1!
1%
1-
12
#766940000000
0!
0%
b11 *
0-
02
b11 6
#766950000000
1!
1%
1-
12
15
#766960000000
0!
0%
b100 *
0-
02
b100 6
#766970000000
1!
1%
1-
12
#766980000000
0!
0%
b101 *
0-
02
b101 6
#766990000000
1!
1%
1-
12
#767000000000
0!
0%
b110 *
0-
02
b110 6
#767010000000
1!
1%
1-
12
#767020000000
0!
0%
b111 *
0-
02
b111 6
#767030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#767040000000
0!
0%
b0 *
0-
02
b0 6
#767050000000
1!
1%
1-
12
#767060000000
0!
0%
b1 *
0-
02
b1 6
#767070000000
1!
1%
1-
12
#767080000000
0!
0%
b10 *
0-
02
b10 6
#767090000000
1!
1%
1-
12
#767100000000
0!
0%
b11 *
0-
02
b11 6
#767110000000
1!
1%
1-
12
15
#767120000000
0!
0%
b100 *
0-
02
b100 6
#767130000000
1!
1%
1-
12
#767140000000
0!
0%
b101 *
0-
02
b101 6
#767150000000
1!
1%
1-
12
#767160000000
0!
0%
b110 *
0-
02
b110 6
#767170000000
1!
1%
1-
12
#767180000000
0!
0%
b111 *
0-
02
b111 6
#767190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#767200000000
0!
0%
b0 *
0-
02
b0 6
#767210000000
1!
1%
1-
12
#767220000000
0!
0%
b1 *
0-
02
b1 6
#767230000000
1!
1%
1-
12
#767240000000
0!
0%
b10 *
0-
02
b10 6
#767250000000
1!
1%
1-
12
#767260000000
0!
0%
b11 *
0-
02
b11 6
#767270000000
1!
1%
1-
12
15
#767280000000
0!
0%
b100 *
0-
02
b100 6
#767290000000
1!
1%
1-
12
#767300000000
0!
0%
b101 *
0-
02
b101 6
#767310000000
1!
1%
1-
12
#767320000000
0!
0%
b110 *
0-
02
b110 6
#767330000000
1!
1%
1-
12
#767340000000
0!
0%
b111 *
0-
02
b111 6
#767350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#767360000000
0!
0%
b0 *
0-
02
b0 6
#767370000000
1!
1%
1-
12
#767380000000
0!
0%
b1 *
0-
02
b1 6
#767390000000
1!
1%
1-
12
#767400000000
0!
0%
b10 *
0-
02
b10 6
#767410000000
1!
1%
1-
12
#767420000000
0!
0%
b11 *
0-
02
b11 6
#767430000000
1!
1%
1-
12
15
#767440000000
0!
0%
b100 *
0-
02
b100 6
#767450000000
1!
1%
1-
12
#767460000000
0!
0%
b101 *
0-
02
b101 6
#767470000000
1!
1%
1-
12
#767480000000
0!
0%
b110 *
0-
02
b110 6
#767490000000
1!
1%
1-
12
#767500000000
0!
0%
b111 *
0-
02
b111 6
#767510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#767520000000
0!
0%
b0 *
0-
02
b0 6
#767530000000
1!
1%
1-
12
#767540000000
0!
0%
b1 *
0-
02
b1 6
#767550000000
1!
1%
1-
12
#767560000000
0!
0%
b10 *
0-
02
b10 6
#767570000000
1!
1%
1-
12
#767580000000
0!
0%
b11 *
0-
02
b11 6
#767590000000
1!
1%
1-
12
15
#767600000000
0!
0%
b100 *
0-
02
b100 6
#767610000000
1!
1%
1-
12
#767620000000
0!
0%
b101 *
0-
02
b101 6
#767630000000
1!
1%
1-
12
#767640000000
0!
0%
b110 *
0-
02
b110 6
#767650000000
1!
1%
1-
12
#767660000000
0!
0%
b111 *
0-
02
b111 6
#767670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#767680000000
0!
0%
b0 *
0-
02
b0 6
#767690000000
1!
1%
1-
12
#767700000000
0!
0%
b1 *
0-
02
b1 6
#767710000000
1!
1%
1-
12
#767720000000
0!
0%
b10 *
0-
02
b10 6
#767730000000
1!
1%
1-
12
#767740000000
0!
0%
b11 *
0-
02
b11 6
#767750000000
1!
1%
1-
12
15
#767760000000
0!
0%
b100 *
0-
02
b100 6
#767770000000
1!
1%
1-
12
#767780000000
0!
0%
b101 *
0-
02
b101 6
#767790000000
1!
1%
1-
12
#767800000000
0!
0%
b110 *
0-
02
b110 6
#767810000000
1!
1%
1-
12
#767820000000
0!
0%
b111 *
0-
02
b111 6
#767830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#767840000000
0!
0%
b0 *
0-
02
b0 6
#767850000000
1!
1%
1-
12
#767860000000
0!
0%
b1 *
0-
02
b1 6
#767870000000
1!
1%
1-
12
#767880000000
0!
0%
b10 *
0-
02
b10 6
#767890000000
1!
1%
1-
12
#767900000000
0!
0%
b11 *
0-
02
b11 6
#767910000000
1!
1%
1-
12
15
#767920000000
0!
0%
b100 *
0-
02
b100 6
#767930000000
1!
1%
1-
12
#767940000000
0!
0%
b101 *
0-
02
b101 6
#767950000000
1!
1%
1-
12
#767960000000
0!
0%
b110 *
0-
02
b110 6
#767970000000
1!
1%
1-
12
#767980000000
0!
0%
b111 *
0-
02
b111 6
#767990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#768000000000
0!
0%
b0 *
0-
02
b0 6
#768010000000
1!
1%
1-
12
#768020000000
0!
0%
b1 *
0-
02
b1 6
#768030000000
1!
1%
1-
12
#768040000000
0!
0%
b10 *
0-
02
b10 6
#768050000000
1!
1%
1-
12
#768060000000
0!
0%
b11 *
0-
02
b11 6
#768070000000
1!
1%
1-
12
15
#768080000000
0!
0%
b100 *
0-
02
b100 6
#768090000000
1!
1%
1-
12
#768100000000
0!
0%
b101 *
0-
02
b101 6
#768110000000
1!
1%
1-
12
#768120000000
0!
0%
b110 *
0-
02
b110 6
#768130000000
1!
1%
1-
12
#768140000000
0!
0%
b111 *
0-
02
b111 6
#768150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#768160000000
0!
0%
b0 *
0-
02
b0 6
#768170000000
1!
1%
1-
12
#768180000000
0!
0%
b1 *
0-
02
b1 6
#768190000000
1!
1%
1-
12
#768200000000
0!
0%
b10 *
0-
02
b10 6
#768210000000
1!
1%
1-
12
#768220000000
0!
0%
b11 *
0-
02
b11 6
#768230000000
1!
1%
1-
12
15
#768240000000
0!
0%
b100 *
0-
02
b100 6
#768250000000
1!
1%
1-
12
#768260000000
0!
0%
b101 *
0-
02
b101 6
#768270000000
1!
1%
1-
12
#768280000000
0!
0%
b110 *
0-
02
b110 6
#768290000000
1!
1%
1-
12
#768300000000
0!
0%
b111 *
0-
02
b111 6
#768310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#768320000000
0!
0%
b0 *
0-
02
b0 6
#768330000000
1!
1%
1-
12
#768340000000
0!
0%
b1 *
0-
02
b1 6
#768350000000
1!
1%
1-
12
#768360000000
0!
0%
b10 *
0-
02
b10 6
#768370000000
1!
1%
1-
12
#768380000000
0!
0%
b11 *
0-
02
b11 6
#768390000000
1!
1%
1-
12
15
#768400000000
0!
0%
b100 *
0-
02
b100 6
#768410000000
1!
1%
1-
12
#768420000000
0!
0%
b101 *
0-
02
b101 6
#768430000000
1!
1%
1-
12
#768440000000
0!
0%
b110 *
0-
02
b110 6
#768450000000
1!
1%
1-
12
#768460000000
0!
0%
b111 *
0-
02
b111 6
#768470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#768480000000
0!
0%
b0 *
0-
02
b0 6
#768490000000
1!
1%
1-
12
#768500000000
0!
0%
b1 *
0-
02
b1 6
#768510000000
1!
1%
1-
12
#768520000000
0!
0%
b10 *
0-
02
b10 6
#768530000000
1!
1%
1-
12
#768540000000
0!
0%
b11 *
0-
02
b11 6
#768550000000
1!
1%
1-
12
15
#768560000000
0!
0%
b100 *
0-
02
b100 6
#768570000000
1!
1%
1-
12
#768580000000
0!
0%
b101 *
0-
02
b101 6
#768590000000
1!
1%
1-
12
#768600000000
0!
0%
b110 *
0-
02
b110 6
#768610000000
1!
1%
1-
12
#768620000000
0!
0%
b111 *
0-
02
b111 6
#768630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#768640000000
0!
0%
b0 *
0-
02
b0 6
#768650000000
1!
1%
1-
12
#768660000000
0!
0%
b1 *
0-
02
b1 6
#768670000000
1!
1%
1-
12
#768680000000
0!
0%
b10 *
0-
02
b10 6
#768690000000
1!
1%
1-
12
#768700000000
0!
0%
b11 *
0-
02
b11 6
#768710000000
1!
1%
1-
12
15
#768720000000
0!
0%
b100 *
0-
02
b100 6
#768730000000
1!
1%
1-
12
#768740000000
0!
0%
b101 *
0-
02
b101 6
#768750000000
1!
1%
1-
12
#768760000000
0!
0%
b110 *
0-
02
b110 6
#768770000000
1!
1%
1-
12
#768780000000
0!
0%
b111 *
0-
02
b111 6
#768790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#768800000000
0!
0%
b0 *
0-
02
b0 6
#768810000000
1!
1%
1-
12
#768820000000
0!
0%
b1 *
0-
02
b1 6
#768830000000
1!
1%
1-
12
#768840000000
0!
0%
b10 *
0-
02
b10 6
#768850000000
1!
1%
1-
12
#768860000000
0!
0%
b11 *
0-
02
b11 6
#768870000000
1!
1%
1-
12
15
#768880000000
0!
0%
b100 *
0-
02
b100 6
#768890000000
1!
1%
1-
12
#768900000000
0!
0%
b101 *
0-
02
b101 6
#768910000000
1!
1%
1-
12
#768920000000
0!
0%
b110 *
0-
02
b110 6
#768930000000
1!
1%
1-
12
#768940000000
0!
0%
b111 *
0-
02
b111 6
#768950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#768960000000
0!
0%
b0 *
0-
02
b0 6
#768970000000
1!
1%
1-
12
#768980000000
0!
0%
b1 *
0-
02
b1 6
#768990000000
1!
1%
1-
12
#769000000000
0!
0%
b10 *
0-
02
b10 6
#769010000000
1!
1%
1-
12
#769020000000
0!
0%
b11 *
0-
02
b11 6
#769030000000
1!
1%
1-
12
15
#769040000000
0!
0%
b100 *
0-
02
b100 6
#769050000000
1!
1%
1-
12
#769060000000
0!
0%
b101 *
0-
02
b101 6
#769070000000
1!
1%
1-
12
#769080000000
0!
0%
b110 *
0-
02
b110 6
#769090000000
1!
1%
1-
12
#769100000000
0!
0%
b111 *
0-
02
b111 6
#769110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#769120000000
0!
0%
b0 *
0-
02
b0 6
#769130000000
1!
1%
1-
12
#769140000000
0!
0%
b1 *
0-
02
b1 6
#769150000000
1!
1%
1-
12
#769160000000
0!
0%
b10 *
0-
02
b10 6
#769170000000
1!
1%
1-
12
#769180000000
0!
0%
b11 *
0-
02
b11 6
#769190000000
1!
1%
1-
12
15
#769200000000
0!
0%
b100 *
0-
02
b100 6
#769210000000
1!
1%
1-
12
#769220000000
0!
0%
b101 *
0-
02
b101 6
#769230000000
1!
1%
1-
12
#769240000000
0!
0%
b110 *
0-
02
b110 6
#769250000000
1!
1%
1-
12
#769260000000
0!
0%
b111 *
0-
02
b111 6
#769270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#769280000000
0!
0%
b0 *
0-
02
b0 6
#769290000000
1!
1%
1-
12
#769300000000
0!
0%
b1 *
0-
02
b1 6
#769310000000
1!
1%
1-
12
#769320000000
0!
0%
b10 *
0-
02
b10 6
#769330000000
1!
1%
1-
12
#769340000000
0!
0%
b11 *
0-
02
b11 6
#769350000000
1!
1%
1-
12
15
#769360000000
0!
0%
b100 *
0-
02
b100 6
#769370000000
1!
1%
1-
12
#769380000000
0!
0%
b101 *
0-
02
b101 6
#769390000000
1!
1%
1-
12
#769400000000
0!
0%
b110 *
0-
02
b110 6
#769410000000
1!
1%
1-
12
#769420000000
0!
0%
b111 *
0-
02
b111 6
#769430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#769440000000
0!
0%
b0 *
0-
02
b0 6
#769450000000
1!
1%
1-
12
#769460000000
0!
0%
b1 *
0-
02
b1 6
#769470000000
1!
1%
1-
12
#769480000000
0!
0%
b10 *
0-
02
b10 6
#769490000000
1!
1%
1-
12
#769500000000
0!
0%
b11 *
0-
02
b11 6
#769510000000
1!
1%
1-
12
15
#769520000000
0!
0%
b100 *
0-
02
b100 6
#769530000000
1!
1%
1-
12
#769540000000
0!
0%
b101 *
0-
02
b101 6
#769550000000
1!
1%
1-
12
#769560000000
0!
0%
b110 *
0-
02
b110 6
#769570000000
1!
1%
1-
12
#769580000000
0!
0%
b111 *
0-
02
b111 6
#769590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#769600000000
0!
0%
b0 *
0-
02
b0 6
#769610000000
1!
1%
1-
12
#769620000000
0!
0%
b1 *
0-
02
b1 6
#769630000000
1!
1%
1-
12
#769640000000
0!
0%
b10 *
0-
02
b10 6
#769650000000
1!
1%
1-
12
#769660000000
0!
0%
b11 *
0-
02
b11 6
#769670000000
1!
1%
1-
12
15
#769680000000
0!
0%
b100 *
0-
02
b100 6
#769690000000
1!
1%
1-
12
#769700000000
0!
0%
b101 *
0-
02
b101 6
#769710000000
1!
1%
1-
12
#769720000000
0!
0%
b110 *
0-
02
b110 6
#769730000000
1!
1%
1-
12
#769740000000
0!
0%
b111 *
0-
02
b111 6
#769750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#769760000000
0!
0%
b0 *
0-
02
b0 6
#769770000000
1!
1%
1-
12
#769780000000
0!
0%
b1 *
0-
02
b1 6
#769790000000
1!
1%
1-
12
#769800000000
0!
0%
b10 *
0-
02
b10 6
#769810000000
1!
1%
1-
12
#769820000000
0!
0%
b11 *
0-
02
b11 6
#769830000000
1!
1%
1-
12
15
#769840000000
0!
0%
b100 *
0-
02
b100 6
#769850000000
1!
1%
1-
12
#769860000000
0!
0%
b101 *
0-
02
b101 6
#769870000000
1!
1%
1-
12
#769880000000
0!
0%
b110 *
0-
02
b110 6
#769890000000
1!
1%
1-
12
#769900000000
0!
0%
b111 *
0-
02
b111 6
#769910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#769920000000
0!
0%
b0 *
0-
02
b0 6
#769930000000
1!
1%
1-
12
#769940000000
0!
0%
b1 *
0-
02
b1 6
#769950000000
1!
1%
1-
12
#769960000000
0!
0%
b10 *
0-
02
b10 6
#769970000000
1!
1%
1-
12
#769980000000
0!
0%
b11 *
0-
02
b11 6
#769990000000
1!
1%
1-
12
15
#770000000000
0!
0%
b100 *
0-
02
b100 6
#770010000000
1!
1%
1-
12
#770020000000
0!
0%
b101 *
0-
02
b101 6
#770030000000
1!
1%
1-
12
#770040000000
0!
0%
b110 *
0-
02
b110 6
#770050000000
1!
1%
1-
12
#770060000000
0!
0%
b111 *
0-
02
b111 6
#770070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#770080000000
0!
0%
b0 *
0-
02
b0 6
#770090000000
1!
1%
1-
12
#770100000000
0!
0%
b1 *
0-
02
b1 6
#770110000000
1!
1%
1-
12
#770120000000
0!
0%
b10 *
0-
02
b10 6
#770130000000
1!
1%
1-
12
#770140000000
0!
0%
b11 *
0-
02
b11 6
#770150000000
1!
1%
1-
12
15
#770160000000
0!
0%
b100 *
0-
02
b100 6
#770170000000
1!
1%
1-
12
#770180000000
0!
0%
b101 *
0-
02
b101 6
#770190000000
1!
1%
1-
12
#770200000000
0!
0%
b110 *
0-
02
b110 6
#770210000000
1!
1%
1-
12
#770220000000
0!
0%
b111 *
0-
02
b111 6
#770230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#770240000000
0!
0%
b0 *
0-
02
b0 6
#770250000000
1!
1%
1-
12
#770260000000
0!
0%
b1 *
0-
02
b1 6
#770270000000
1!
1%
1-
12
#770280000000
0!
0%
b10 *
0-
02
b10 6
#770290000000
1!
1%
1-
12
#770300000000
0!
0%
b11 *
0-
02
b11 6
#770310000000
1!
1%
1-
12
15
#770320000000
0!
0%
b100 *
0-
02
b100 6
#770330000000
1!
1%
1-
12
#770340000000
0!
0%
b101 *
0-
02
b101 6
#770350000000
1!
1%
1-
12
#770360000000
0!
0%
b110 *
0-
02
b110 6
#770370000000
1!
1%
1-
12
#770380000000
0!
0%
b111 *
0-
02
b111 6
#770390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#770400000000
0!
0%
b0 *
0-
02
b0 6
#770410000000
1!
1%
1-
12
#770420000000
0!
0%
b1 *
0-
02
b1 6
#770430000000
1!
1%
1-
12
#770440000000
0!
0%
b10 *
0-
02
b10 6
#770450000000
1!
1%
1-
12
#770460000000
0!
0%
b11 *
0-
02
b11 6
#770470000000
1!
1%
1-
12
15
#770480000000
0!
0%
b100 *
0-
02
b100 6
#770490000000
1!
1%
1-
12
#770500000000
0!
0%
b101 *
0-
02
b101 6
#770510000000
1!
1%
1-
12
#770520000000
0!
0%
b110 *
0-
02
b110 6
#770530000000
1!
1%
1-
12
#770540000000
0!
0%
b111 *
0-
02
b111 6
#770550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#770560000000
0!
0%
b0 *
0-
02
b0 6
#770570000000
1!
1%
1-
12
#770580000000
0!
0%
b1 *
0-
02
b1 6
#770590000000
1!
1%
1-
12
#770600000000
0!
0%
b10 *
0-
02
b10 6
#770610000000
1!
1%
1-
12
#770620000000
0!
0%
b11 *
0-
02
b11 6
#770630000000
1!
1%
1-
12
15
#770640000000
0!
0%
b100 *
0-
02
b100 6
#770650000000
1!
1%
1-
12
#770660000000
0!
0%
b101 *
0-
02
b101 6
#770670000000
1!
1%
1-
12
#770680000000
0!
0%
b110 *
0-
02
b110 6
#770690000000
1!
1%
1-
12
#770700000000
0!
0%
b111 *
0-
02
b111 6
#770710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#770720000000
0!
0%
b0 *
0-
02
b0 6
#770730000000
1!
1%
1-
12
#770740000000
0!
0%
b1 *
0-
02
b1 6
#770750000000
1!
1%
1-
12
#770760000000
0!
0%
b10 *
0-
02
b10 6
#770770000000
1!
1%
1-
12
#770780000000
0!
0%
b11 *
0-
02
b11 6
#770790000000
1!
1%
1-
12
15
#770800000000
0!
0%
b100 *
0-
02
b100 6
#770810000000
1!
1%
1-
12
#770820000000
0!
0%
b101 *
0-
02
b101 6
#770830000000
1!
1%
1-
12
#770840000000
0!
0%
b110 *
0-
02
b110 6
#770850000000
1!
1%
1-
12
#770860000000
0!
0%
b111 *
0-
02
b111 6
#770870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#770880000000
0!
0%
b0 *
0-
02
b0 6
#770890000000
1!
1%
1-
12
#770900000000
0!
0%
b1 *
0-
02
b1 6
#770910000000
1!
1%
1-
12
#770920000000
0!
0%
b10 *
0-
02
b10 6
#770930000000
1!
1%
1-
12
#770940000000
0!
0%
b11 *
0-
02
b11 6
#770950000000
1!
1%
1-
12
15
#770960000000
0!
0%
b100 *
0-
02
b100 6
#770970000000
1!
1%
1-
12
#770980000000
0!
0%
b101 *
0-
02
b101 6
#770990000000
1!
1%
1-
12
#771000000000
0!
0%
b110 *
0-
02
b110 6
#771010000000
1!
1%
1-
12
#771020000000
0!
0%
b111 *
0-
02
b111 6
#771030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#771040000000
0!
0%
b0 *
0-
02
b0 6
#771050000000
1!
1%
1-
12
#771060000000
0!
0%
b1 *
0-
02
b1 6
#771070000000
1!
1%
1-
12
#771080000000
0!
0%
b10 *
0-
02
b10 6
#771090000000
1!
1%
1-
12
#771100000000
0!
0%
b11 *
0-
02
b11 6
#771110000000
1!
1%
1-
12
15
#771120000000
0!
0%
b100 *
0-
02
b100 6
#771130000000
1!
1%
1-
12
#771140000000
0!
0%
b101 *
0-
02
b101 6
#771150000000
1!
1%
1-
12
#771160000000
0!
0%
b110 *
0-
02
b110 6
#771170000000
1!
1%
1-
12
#771180000000
0!
0%
b111 *
0-
02
b111 6
#771190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#771200000000
0!
0%
b0 *
0-
02
b0 6
#771210000000
1!
1%
1-
12
#771220000000
0!
0%
b1 *
0-
02
b1 6
#771230000000
1!
1%
1-
12
#771240000000
0!
0%
b10 *
0-
02
b10 6
#771250000000
1!
1%
1-
12
#771260000000
0!
0%
b11 *
0-
02
b11 6
#771270000000
1!
1%
1-
12
15
#771280000000
0!
0%
b100 *
0-
02
b100 6
#771290000000
1!
1%
1-
12
#771300000000
0!
0%
b101 *
0-
02
b101 6
#771310000000
1!
1%
1-
12
#771320000000
0!
0%
b110 *
0-
02
b110 6
#771330000000
1!
1%
1-
12
#771340000000
0!
0%
b111 *
0-
02
b111 6
#771350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#771360000000
0!
0%
b0 *
0-
02
b0 6
#771370000000
1!
1%
1-
12
#771380000000
0!
0%
b1 *
0-
02
b1 6
#771390000000
1!
1%
1-
12
#771400000000
0!
0%
b10 *
0-
02
b10 6
#771410000000
1!
1%
1-
12
#771420000000
0!
0%
b11 *
0-
02
b11 6
#771430000000
1!
1%
1-
12
15
#771440000000
0!
0%
b100 *
0-
02
b100 6
#771450000000
1!
1%
1-
12
#771460000000
0!
0%
b101 *
0-
02
b101 6
#771470000000
1!
1%
1-
12
#771480000000
0!
0%
b110 *
0-
02
b110 6
#771490000000
1!
1%
1-
12
#771500000000
0!
0%
b111 *
0-
02
b111 6
#771510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#771520000000
0!
0%
b0 *
0-
02
b0 6
#771530000000
1!
1%
1-
12
#771540000000
0!
0%
b1 *
0-
02
b1 6
#771550000000
1!
1%
1-
12
#771560000000
0!
0%
b10 *
0-
02
b10 6
#771570000000
1!
1%
1-
12
#771580000000
0!
0%
b11 *
0-
02
b11 6
#771590000000
1!
1%
1-
12
15
#771600000000
0!
0%
b100 *
0-
02
b100 6
#771610000000
1!
1%
1-
12
#771620000000
0!
0%
b101 *
0-
02
b101 6
#771630000000
1!
1%
1-
12
#771640000000
0!
0%
b110 *
0-
02
b110 6
#771650000000
1!
1%
1-
12
#771660000000
0!
0%
b111 *
0-
02
b111 6
#771670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#771680000000
0!
0%
b0 *
0-
02
b0 6
#771690000000
1!
1%
1-
12
#771700000000
0!
0%
b1 *
0-
02
b1 6
#771710000000
1!
1%
1-
12
#771720000000
0!
0%
b10 *
0-
02
b10 6
#771730000000
1!
1%
1-
12
#771740000000
0!
0%
b11 *
0-
02
b11 6
#771750000000
1!
1%
1-
12
15
#771760000000
0!
0%
b100 *
0-
02
b100 6
#771770000000
1!
1%
1-
12
#771780000000
0!
0%
b101 *
0-
02
b101 6
#771790000000
1!
1%
1-
12
#771800000000
0!
0%
b110 *
0-
02
b110 6
#771810000000
1!
1%
1-
12
#771820000000
0!
0%
b111 *
0-
02
b111 6
#771830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#771840000000
0!
0%
b0 *
0-
02
b0 6
#771850000000
1!
1%
1-
12
#771860000000
0!
0%
b1 *
0-
02
b1 6
#771870000000
1!
1%
1-
12
#771880000000
0!
0%
b10 *
0-
02
b10 6
#771890000000
1!
1%
1-
12
#771900000000
0!
0%
b11 *
0-
02
b11 6
#771910000000
1!
1%
1-
12
15
#771920000000
0!
0%
b100 *
0-
02
b100 6
#771930000000
1!
1%
1-
12
#771940000000
0!
0%
b101 *
0-
02
b101 6
#771950000000
1!
1%
1-
12
#771960000000
0!
0%
b110 *
0-
02
b110 6
#771970000000
1!
1%
1-
12
#771980000000
0!
0%
b111 *
0-
02
b111 6
#771990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#772000000000
0!
0%
b0 *
0-
02
b0 6
#772010000000
1!
1%
1-
12
#772020000000
0!
0%
b1 *
0-
02
b1 6
#772030000000
1!
1%
1-
12
#772040000000
0!
0%
b10 *
0-
02
b10 6
#772050000000
1!
1%
1-
12
#772060000000
0!
0%
b11 *
0-
02
b11 6
#772070000000
1!
1%
1-
12
15
#772080000000
0!
0%
b100 *
0-
02
b100 6
#772090000000
1!
1%
1-
12
#772100000000
0!
0%
b101 *
0-
02
b101 6
#772110000000
1!
1%
1-
12
#772120000000
0!
0%
b110 *
0-
02
b110 6
#772130000000
1!
1%
1-
12
#772140000000
0!
0%
b111 *
0-
02
b111 6
#772150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#772160000000
0!
0%
b0 *
0-
02
b0 6
#772170000000
1!
1%
1-
12
#772180000000
0!
0%
b1 *
0-
02
b1 6
#772190000000
1!
1%
1-
12
#772200000000
0!
0%
b10 *
0-
02
b10 6
#772210000000
1!
1%
1-
12
#772220000000
0!
0%
b11 *
0-
02
b11 6
#772230000000
1!
1%
1-
12
15
#772240000000
0!
0%
b100 *
0-
02
b100 6
#772250000000
1!
1%
1-
12
#772260000000
0!
0%
b101 *
0-
02
b101 6
#772270000000
1!
1%
1-
12
#772280000000
0!
0%
b110 *
0-
02
b110 6
#772290000000
1!
1%
1-
12
#772300000000
0!
0%
b111 *
0-
02
b111 6
#772310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#772320000000
0!
0%
b0 *
0-
02
b0 6
#772330000000
1!
1%
1-
12
#772340000000
0!
0%
b1 *
0-
02
b1 6
#772350000000
1!
1%
1-
12
#772360000000
0!
0%
b10 *
0-
02
b10 6
#772370000000
1!
1%
1-
12
#772380000000
0!
0%
b11 *
0-
02
b11 6
#772390000000
1!
1%
1-
12
15
#772400000000
0!
0%
b100 *
0-
02
b100 6
#772410000000
1!
1%
1-
12
#772420000000
0!
0%
b101 *
0-
02
b101 6
#772430000000
1!
1%
1-
12
#772440000000
0!
0%
b110 *
0-
02
b110 6
#772450000000
1!
1%
1-
12
#772460000000
0!
0%
b111 *
0-
02
b111 6
#772470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#772480000000
0!
0%
b0 *
0-
02
b0 6
#772490000000
1!
1%
1-
12
#772500000000
0!
0%
b1 *
0-
02
b1 6
#772510000000
1!
1%
1-
12
#772520000000
0!
0%
b10 *
0-
02
b10 6
#772530000000
1!
1%
1-
12
#772540000000
0!
0%
b11 *
0-
02
b11 6
#772550000000
1!
1%
1-
12
15
#772560000000
0!
0%
b100 *
0-
02
b100 6
#772570000000
1!
1%
1-
12
#772580000000
0!
0%
b101 *
0-
02
b101 6
#772590000000
1!
1%
1-
12
#772600000000
0!
0%
b110 *
0-
02
b110 6
#772610000000
1!
1%
1-
12
#772620000000
0!
0%
b111 *
0-
02
b111 6
#772630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#772640000000
0!
0%
b0 *
0-
02
b0 6
#772650000000
1!
1%
1-
12
#772660000000
0!
0%
b1 *
0-
02
b1 6
#772670000000
1!
1%
1-
12
#772680000000
0!
0%
b10 *
0-
02
b10 6
#772690000000
1!
1%
1-
12
#772700000000
0!
0%
b11 *
0-
02
b11 6
#772710000000
1!
1%
1-
12
15
#772720000000
0!
0%
b100 *
0-
02
b100 6
#772730000000
1!
1%
1-
12
#772740000000
0!
0%
b101 *
0-
02
b101 6
#772750000000
1!
1%
1-
12
#772760000000
0!
0%
b110 *
0-
02
b110 6
#772770000000
1!
1%
1-
12
#772780000000
0!
0%
b111 *
0-
02
b111 6
#772790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#772800000000
0!
0%
b0 *
0-
02
b0 6
#772810000000
1!
1%
1-
12
#772820000000
0!
0%
b1 *
0-
02
b1 6
#772830000000
1!
1%
1-
12
#772840000000
0!
0%
b10 *
0-
02
b10 6
#772850000000
1!
1%
1-
12
#772860000000
0!
0%
b11 *
0-
02
b11 6
#772870000000
1!
1%
1-
12
15
#772880000000
0!
0%
b100 *
0-
02
b100 6
#772890000000
1!
1%
1-
12
#772900000000
0!
0%
b101 *
0-
02
b101 6
#772910000000
1!
1%
1-
12
#772920000000
0!
0%
b110 *
0-
02
b110 6
#772930000000
1!
1%
1-
12
#772940000000
0!
0%
b111 *
0-
02
b111 6
#772950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#772960000000
0!
0%
b0 *
0-
02
b0 6
#772970000000
1!
1%
1-
12
#772980000000
0!
0%
b1 *
0-
02
b1 6
#772990000000
1!
1%
1-
12
#773000000000
0!
0%
b10 *
0-
02
b10 6
#773010000000
1!
1%
1-
12
#773020000000
0!
0%
b11 *
0-
02
b11 6
#773030000000
1!
1%
1-
12
15
#773040000000
0!
0%
b100 *
0-
02
b100 6
#773050000000
1!
1%
1-
12
#773060000000
0!
0%
b101 *
0-
02
b101 6
#773070000000
1!
1%
1-
12
#773080000000
0!
0%
b110 *
0-
02
b110 6
#773090000000
1!
1%
1-
12
#773100000000
0!
0%
b111 *
0-
02
b111 6
#773110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#773120000000
0!
0%
b0 *
0-
02
b0 6
#773130000000
1!
1%
1-
12
#773140000000
0!
0%
b1 *
0-
02
b1 6
#773150000000
1!
1%
1-
12
#773160000000
0!
0%
b10 *
0-
02
b10 6
#773170000000
1!
1%
1-
12
#773180000000
0!
0%
b11 *
0-
02
b11 6
#773190000000
1!
1%
1-
12
15
#773200000000
0!
0%
b100 *
0-
02
b100 6
#773210000000
1!
1%
1-
12
#773220000000
0!
0%
b101 *
0-
02
b101 6
#773230000000
1!
1%
1-
12
#773240000000
0!
0%
b110 *
0-
02
b110 6
#773250000000
1!
1%
1-
12
#773260000000
0!
0%
b111 *
0-
02
b111 6
#773270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#773280000000
0!
0%
b0 *
0-
02
b0 6
#773290000000
1!
1%
1-
12
#773300000000
0!
0%
b1 *
0-
02
b1 6
#773310000000
1!
1%
1-
12
#773320000000
0!
0%
b10 *
0-
02
b10 6
#773330000000
1!
1%
1-
12
#773340000000
0!
0%
b11 *
0-
02
b11 6
#773350000000
1!
1%
1-
12
15
#773360000000
0!
0%
b100 *
0-
02
b100 6
#773370000000
1!
1%
1-
12
#773380000000
0!
0%
b101 *
0-
02
b101 6
#773390000000
1!
1%
1-
12
#773400000000
0!
0%
b110 *
0-
02
b110 6
#773410000000
1!
1%
1-
12
#773420000000
0!
0%
b111 *
0-
02
b111 6
#773430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#773440000000
0!
0%
b0 *
0-
02
b0 6
#773450000000
1!
1%
1-
12
#773460000000
0!
0%
b1 *
0-
02
b1 6
#773470000000
1!
1%
1-
12
#773480000000
0!
0%
b10 *
0-
02
b10 6
#773490000000
1!
1%
1-
12
#773500000000
0!
0%
b11 *
0-
02
b11 6
#773510000000
1!
1%
1-
12
15
#773520000000
0!
0%
b100 *
0-
02
b100 6
#773530000000
1!
1%
1-
12
#773540000000
0!
0%
b101 *
0-
02
b101 6
#773550000000
1!
1%
1-
12
#773560000000
0!
0%
b110 *
0-
02
b110 6
#773570000000
1!
1%
1-
12
#773580000000
0!
0%
b111 *
0-
02
b111 6
#773590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#773600000000
0!
0%
b0 *
0-
02
b0 6
#773610000000
1!
1%
1-
12
#773620000000
0!
0%
b1 *
0-
02
b1 6
#773630000000
1!
1%
1-
12
#773640000000
0!
0%
b10 *
0-
02
b10 6
#773650000000
1!
1%
1-
12
#773660000000
0!
0%
b11 *
0-
02
b11 6
#773670000000
1!
1%
1-
12
15
#773680000000
0!
0%
b100 *
0-
02
b100 6
#773690000000
1!
1%
1-
12
#773700000000
0!
0%
b101 *
0-
02
b101 6
#773710000000
1!
1%
1-
12
#773720000000
0!
0%
b110 *
0-
02
b110 6
#773730000000
1!
1%
1-
12
#773740000000
0!
0%
b111 *
0-
02
b111 6
#773750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#773760000000
0!
0%
b0 *
0-
02
b0 6
#773770000000
1!
1%
1-
12
#773780000000
0!
0%
b1 *
0-
02
b1 6
#773790000000
1!
1%
1-
12
#773800000000
0!
0%
b10 *
0-
02
b10 6
#773810000000
1!
1%
1-
12
#773820000000
0!
0%
b11 *
0-
02
b11 6
#773830000000
1!
1%
1-
12
15
#773840000000
0!
0%
b100 *
0-
02
b100 6
#773850000000
1!
1%
1-
12
#773860000000
0!
0%
b101 *
0-
02
b101 6
#773870000000
1!
1%
1-
12
#773880000000
0!
0%
b110 *
0-
02
b110 6
#773890000000
1!
1%
1-
12
#773900000000
0!
0%
b111 *
0-
02
b111 6
#773910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#773920000000
0!
0%
b0 *
0-
02
b0 6
#773930000000
1!
1%
1-
12
#773940000000
0!
0%
b1 *
0-
02
b1 6
#773950000000
1!
1%
1-
12
#773960000000
0!
0%
b10 *
0-
02
b10 6
#773970000000
1!
1%
1-
12
#773980000000
0!
0%
b11 *
0-
02
b11 6
#773990000000
1!
1%
1-
12
15
#774000000000
0!
0%
b100 *
0-
02
b100 6
#774010000000
1!
1%
1-
12
#774020000000
0!
0%
b101 *
0-
02
b101 6
#774030000000
1!
1%
1-
12
#774040000000
0!
0%
b110 *
0-
02
b110 6
#774050000000
1!
1%
1-
12
#774060000000
0!
0%
b111 *
0-
02
b111 6
#774070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#774080000000
0!
0%
b0 *
0-
02
b0 6
#774090000000
1!
1%
1-
12
#774100000000
0!
0%
b1 *
0-
02
b1 6
#774110000000
1!
1%
1-
12
#774120000000
0!
0%
b10 *
0-
02
b10 6
#774130000000
1!
1%
1-
12
#774140000000
0!
0%
b11 *
0-
02
b11 6
#774150000000
1!
1%
1-
12
15
#774160000000
0!
0%
b100 *
0-
02
b100 6
#774170000000
1!
1%
1-
12
#774180000000
0!
0%
b101 *
0-
02
b101 6
#774190000000
1!
1%
1-
12
#774200000000
0!
0%
b110 *
0-
02
b110 6
#774210000000
1!
1%
1-
12
#774220000000
0!
0%
b111 *
0-
02
b111 6
#774230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#774240000000
0!
0%
b0 *
0-
02
b0 6
#774250000000
1!
1%
1-
12
#774260000000
0!
0%
b1 *
0-
02
b1 6
#774270000000
1!
1%
1-
12
#774280000000
0!
0%
b10 *
0-
02
b10 6
#774290000000
1!
1%
1-
12
#774300000000
0!
0%
b11 *
0-
02
b11 6
#774310000000
1!
1%
1-
12
15
#774320000000
0!
0%
b100 *
0-
02
b100 6
#774330000000
1!
1%
1-
12
#774340000000
0!
0%
b101 *
0-
02
b101 6
#774350000000
1!
1%
1-
12
#774360000000
0!
0%
b110 *
0-
02
b110 6
#774370000000
1!
1%
1-
12
#774380000000
0!
0%
b111 *
0-
02
b111 6
#774390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#774400000000
0!
0%
b0 *
0-
02
b0 6
#774410000000
1!
1%
1-
12
#774420000000
0!
0%
b1 *
0-
02
b1 6
#774430000000
1!
1%
1-
12
#774440000000
0!
0%
b10 *
0-
02
b10 6
#774450000000
1!
1%
1-
12
#774460000000
0!
0%
b11 *
0-
02
b11 6
#774470000000
1!
1%
1-
12
15
#774480000000
0!
0%
b100 *
0-
02
b100 6
#774490000000
1!
1%
1-
12
#774500000000
0!
0%
b101 *
0-
02
b101 6
#774510000000
1!
1%
1-
12
#774520000000
0!
0%
b110 *
0-
02
b110 6
#774530000000
1!
1%
1-
12
#774540000000
0!
0%
b111 *
0-
02
b111 6
#774550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#774560000000
0!
0%
b0 *
0-
02
b0 6
#774570000000
1!
1%
1-
12
#774580000000
0!
0%
b1 *
0-
02
b1 6
#774590000000
1!
1%
1-
12
#774600000000
0!
0%
b10 *
0-
02
b10 6
#774610000000
1!
1%
1-
12
#774620000000
0!
0%
b11 *
0-
02
b11 6
#774630000000
1!
1%
1-
12
15
#774640000000
0!
0%
b100 *
0-
02
b100 6
#774650000000
1!
1%
1-
12
#774660000000
0!
0%
b101 *
0-
02
b101 6
#774670000000
1!
1%
1-
12
#774680000000
0!
0%
b110 *
0-
02
b110 6
#774690000000
1!
1%
1-
12
#774700000000
0!
0%
b111 *
0-
02
b111 6
#774710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#774720000000
0!
0%
b0 *
0-
02
b0 6
#774730000000
1!
1%
1-
12
#774740000000
0!
0%
b1 *
0-
02
b1 6
#774750000000
1!
1%
1-
12
#774760000000
0!
0%
b10 *
0-
02
b10 6
#774770000000
1!
1%
1-
12
#774780000000
0!
0%
b11 *
0-
02
b11 6
#774790000000
1!
1%
1-
12
15
#774800000000
0!
0%
b100 *
0-
02
b100 6
#774810000000
1!
1%
1-
12
#774820000000
0!
0%
b101 *
0-
02
b101 6
#774830000000
1!
1%
1-
12
#774840000000
0!
0%
b110 *
0-
02
b110 6
#774850000000
1!
1%
1-
12
#774860000000
0!
0%
b111 *
0-
02
b111 6
#774870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#774880000000
0!
0%
b0 *
0-
02
b0 6
#774890000000
1!
1%
1-
12
#774900000000
0!
0%
b1 *
0-
02
b1 6
#774910000000
1!
1%
1-
12
#774920000000
0!
0%
b10 *
0-
02
b10 6
#774930000000
1!
1%
1-
12
#774940000000
0!
0%
b11 *
0-
02
b11 6
#774950000000
1!
1%
1-
12
15
#774960000000
0!
0%
b100 *
0-
02
b100 6
#774970000000
1!
1%
1-
12
#774980000000
0!
0%
b101 *
0-
02
b101 6
#774990000000
1!
1%
1-
12
#775000000000
0!
0%
b110 *
0-
02
b110 6
#775010000000
1!
1%
1-
12
#775020000000
0!
0%
b111 *
0-
02
b111 6
#775030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#775040000000
0!
0%
b0 *
0-
02
b0 6
#775050000000
1!
1%
1-
12
#775060000000
0!
0%
b1 *
0-
02
b1 6
#775070000000
1!
1%
1-
12
#775080000000
0!
0%
b10 *
0-
02
b10 6
#775090000000
1!
1%
1-
12
#775100000000
0!
0%
b11 *
0-
02
b11 6
#775110000000
1!
1%
1-
12
15
#775120000000
0!
0%
b100 *
0-
02
b100 6
#775130000000
1!
1%
1-
12
#775140000000
0!
0%
b101 *
0-
02
b101 6
#775150000000
1!
1%
1-
12
#775160000000
0!
0%
b110 *
0-
02
b110 6
#775170000000
1!
1%
1-
12
#775180000000
0!
0%
b111 *
0-
02
b111 6
#775190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#775200000000
0!
0%
b0 *
0-
02
b0 6
#775210000000
1!
1%
1-
12
#775220000000
0!
0%
b1 *
0-
02
b1 6
#775230000000
1!
1%
1-
12
#775240000000
0!
0%
b10 *
0-
02
b10 6
#775250000000
1!
1%
1-
12
#775260000000
0!
0%
b11 *
0-
02
b11 6
#775270000000
1!
1%
1-
12
15
#775280000000
0!
0%
b100 *
0-
02
b100 6
#775290000000
1!
1%
1-
12
#775300000000
0!
0%
b101 *
0-
02
b101 6
#775310000000
1!
1%
1-
12
#775320000000
0!
0%
b110 *
0-
02
b110 6
#775330000000
1!
1%
1-
12
#775340000000
0!
0%
b111 *
0-
02
b111 6
#775350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#775360000000
0!
0%
b0 *
0-
02
b0 6
#775370000000
1!
1%
1-
12
#775380000000
0!
0%
b1 *
0-
02
b1 6
#775390000000
1!
1%
1-
12
#775400000000
0!
0%
b10 *
0-
02
b10 6
#775410000000
1!
1%
1-
12
#775420000000
0!
0%
b11 *
0-
02
b11 6
#775430000000
1!
1%
1-
12
15
#775440000000
0!
0%
b100 *
0-
02
b100 6
#775450000000
1!
1%
1-
12
#775460000000
0!
0%
b101 *
0-
02
b101 6
#775470000000
1!
1%
1-
12
#775480000000
0!
0%
b110 *
0-
02
b110 6
#775490000000
1!
1%
1-
12
#775500000000
0!
0%
b111 *
0-
02
b111 6
#775510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#775520000000
0!
0%
b0 *
0-
02
b0 6
#775530000000
1!
1%
1-
12
#775540000000
0!
0%
b1 *
0-
02
b1 6
#775550000000
1!
1%
1-
12
#775560000000
0!
0%
b10 *
0-
02
b10 6
#775570000000
1!
1%
1-
12
#775580000000
0!
0%
b11 *
0-
02
b11 6
#775590000000
1!
1%
1-
12
15
#775600000000
0!
0%
b100 *
0-
02
b100 6
#775610000000
1!
1%
1-
12
#775620000000
0!
0%
b101 *
0-
02
b101 6
#775630000000
1!
1%
1-
12
#775640000000
0!
0%
b110 *
0-
02
b110 6
#775650000000
1!
1%
1-
12
#775660000000
0!
0%
b111 *
0-
02
b111 6
#775670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#775680000000
0!
0%
b0 *
0-
02
b0 6
#775690000000
1!
1%
1-
12
#775700000000
0!
0%
b1 *
0-
02
b1 6
#775710000000
1!
1%
1-
12
#775720000000
0!
0%
b10 *
0-
02
b10 6
#775730000000
1!
1%
1-
12
#775740000000
0!
0%
b11 *
0-
02
b11 6
#775750000000
1!
1%
1-
12
15
#775760000000
0!
0%
b100 *
0-
02
b100 6
#775770000000
1!
1%
1-
12
#775780000000
0!
0%
b101 *
0-
02
b101 6
#775790000000
1!
1%
1-
12
#775800000000
0!
0%
b110 *
0-
02
b110 6
#775810000000
1!
1%
1-
12
#775820000000
0!
0%
b111 *
0-
02
b111 6
#775830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#775840000000
0!
0%
b0 *
0-
02
b0 6
#775850000000
1!
1%
1-
12
#775860000000
0!
0%
b1 *
0-
02
b1 6
#775870000000
1!
1%
1-
12
#775880000000
0!
0%
b10 *
0-
02
b10 6
#775890000000
1!
1%
1-
12
#775900000000
0!
0%
b11 *
0-
02
b11 6
#775910000000
1!
1%
1-
12
15
#775920000000
0!
0%
b100 *
0-
02
b100 6
#775930000000
1!
1%
1-
12
#775940000000
0!
0%
b101 *
0-
02
b101 6
#775950000000
1!
1%
1-
12
#775960000000
0!
0%
b110 *
0-
02
b110 6
#775970000000
1!
1%
1-
12
#775980000000
0!
0%
b111 *
0-
02
b111 6
#775990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#776000000000
0!
0%
b0 *
0-
02
b0 6
#776010000000
1!
1%
1-
12
#776020000000
0!
0%
b1 *
0-
02
b1 6
#776030000000
1!
1%
1-
12
#776040000000
0!
0%
b10 *
0-
02
b10 6
#776050000000
1!
1%
1-
12
#776060000000
0!
0%
b11 *
0-
02
b11 6
#776070000000
1!
1%
1-
12
15
#776080000000
0!
0%
b100 *
0-
02
b100 6
#776090000000
1!
1%
1-
12
#776100000000
0!
0%
b101 *
0-
02
b101 6
#776110000000
1!
1%
1-
12
#776120000000
0!
0%
b110 *
0-
02
b110 6
#776130000000
1!
1%
1-
12
#776140000000
0!
0%
b111 *
0-
02
b111 6
#776150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#776160000000
0!
0%
b0 *
0-
02
b0 6
#776170000000
1!
1%
1-
12
#776180000000
0!
0%
b1 *
0-
02
b1 6
#776190000000
1!
1%
1-
12
#776200000000
0!
0%
b10 *
0-
02
b10 6
#776210000000
1!
1%
1-
12
#776220000000
0!
0%
b11 *
0-
02
b11 6
#776230000000
1!
1%
1-
12
15
#776240000000
0!
0%
b100 *
0-
02
b100 6
#776250000000
1!
1%
1-
12
#776260000000
0!
0%
b101 *
0-
02
b101 6
#776270000000
1!
1%
1-
12
#776280000000
0!
0%
b110 *
0-
02
b110 6
#776290000000
1!
1%
1-
12
#776300000000
0!
0%
b111 *
0-
02
b111 6
#776310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#776320000000
0!
0%
b0 *
0-
02
b0 6
#776330000000
1!
1%
1-
12
#776340000000
0!
0%
b1 *
0-
02
b1 6
#776350000000
1!
1%
1-
12
#776360000000
0!
0%
b10 *
0-
02
b10 6
#776370000000
1!
1%
1-
12
#776380000000
0!
0%
b11 *
0-
02
b11 6
#776390000000
1!
1%
1-
12
15
#776400000000
0!
0%
b100 *
0-
02
b100 6
#776410000000
1!
1%
1-
12
#776420000000
0!
0%
b101 *
0-
02
b101 6
#776430000000
1!
1%
1-
12
#776440000000
0!
0%
b110 *
0-
02
b110 6
#776450000000
1!
1%
1-
12
#776460000000
0!
0%
b111 *
0-
02
b111 6
#776470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#776480000000
0!
0%
b0 *
0-
02
b0 6
#776490000000
1!
1%
1-
12
#776500000000
0!
0%
b1 *
0-
02
b1 6
#776510000000
1!
1%
1-
12
#776520000000
0!
0%
b10 *
0-
02
b10 6
#776530000000
1!
1%
1-
12
#776540000000
0!
0%
b11 *
0-
02
b11 6
#776550000000
1!
1%
1-
12
15
#776560000000
0!
0%
b100 *
0-
02
b100 6
#776570000000
1!
1%
1-
12
#776580000000
0!
0%
b101 *
0-
02
b101 6
#776590000000
1!
1%
1-
12
#776600000000
0!
0%
b110 *
0-
02
b110 6
#776610000000
1!
1%
1-
12
#776620000000
0!
0%
b111 *
0-
02
b111 6
#776630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#776640000000
0!
0%
b0 *
0-
02
b0 6
#776650000000
1!
1%
1-
12
#776660000000
0!
0%
b1 *
0-
02
b1 6
#776670000000
1!
1%
1-
12
#776680000000
0!
0%
b10 *
0-
02
b10 6
#776690000000
1!
1%
1-
12
#776700000000
0!
0%
b11 *
0-
02
b11 6
#776710000000
1!
1%
1-
12
15
#776720000000
0!
0%
b100 *
0-
02
b100 6
#776730000000
1!
1%
1-
12
#776740000000
0!
0%
b101 *
0-
02
b101 6
#776750000000
1!
1%
1-
12
#776760000000
0!
0%
b110 *
0-
02
b110 6
#776770000000
1!
1%
1-
12
#776780000000
0!
0%
b111 *
0-
02
b111 6
#776790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#776800000000
0!
0%
b0 *
0-
02
b0 6
#776810000000
1!
1%
1-
12
#776820000000
0!
0%
b1 *
0-
02
b1 6
#776830000000
1!
1%
1-
12
#776840000000
0!
0%
b10 *
0-
02
b10 6
#776850000000
1!
1%
1-
12
#776860000000
0!
0%
b11 *
0-
02
b11 6
#776870000000
1!
1%
1-
12
15
#776880000000
0!
0%
b100 *
0-
02
b100 6
#776890000000
1!
1%
1-
12
#776900000000
0!
0%
b101 *
0-
02
b101 6
#776910000000
1!
1%
1-
12
#776920000000
0!
0%
b110 *
0-
02
b110 6
#776930000000
1!
1%
1-
12
#776940000000
0!
0%
b111 *
0-
02
b111 6
#776950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#776960000000
0!
0%
b0 *
0-
02
b0 6
#776970000000
1!
1%
1-
12
#776980000000
0!
0%
b1 *
0-
02
b1 6
#776990000000
1!
1%
1-
12
#777000000000
0!
0%
b10 *
0-
02
b10 6
#777010000000
1!
1%
1-
12
#777020000000
0!
0%
b11 *
0-
02
b11 6
#777030000000
1!
1%
1-
12
15
#777040000000
0!
0%
b100 *
0-
02
b100 6
#777050000000
1!
1%
1-
12
#777060000000
0!
0%
b101 *
0-
02
b101 6
#777070000000
1!
1%
1-
12
#777080000000
0!
0%
b110 *
0-
02
b110 6
#777090000000
1!
1%
1-
12
#777100000000
0!
0%
b111 *
0-
02
b111 6
#777110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#777120000000
0!
0%
b0 *
0-
02
b0 6
#777130000000
1!
1%
1-
12
#777140000000
0!
0%
b1 *
0-
02
b1 6
#777150000000
1!
1%
1-
12
#777160000000
0!
0%
b10 *
0-
02
b10 6
#777170000000
1!
1%
1-
12
#777180000000
0!
0%
b11 *
0-
02
b11 6
#777190000000
1!
1%
1-
12
15
#777200000000
0!
0%
b100 *
0-
02
b100 6
#777210000000
1!
1%
1-
12
#777220000000
0!
0%
b101 *
0-
02
b101 6
#777230000000
1!
1%
1-
12
#777240000000
0!
0%
b110 *
0-
02
b110 6
#777250000000
1!
1%
1-
12
#777260000000
0!
0%
b111 *
0-
02
b111 6
#777270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#777280000000
0!
0%
b0 *
0-
02
b0 6
#777290000000
1!
1%
1-
12
#777300000000
0!
0%
b1 *
0-
02
b1 6
#777310000000
1!
1%
1-
12
#777320000000
0!
0%
b10 *
0-
02
b10 6
#777330000000
1!
1%
1-
12
#777340000000
0!
0%
b11 *
0-
02
b11 6
#777350000000
1!
1%
1-
12
15
#777360000000
0!
0%
b100 *
0-
02
b100 6
#777370000000
1!
1%
1-
12
#777380000000
0!
0%
b101 *
0-
02
b101 6
#777390000000
1!
1%
1-
12
#777400000000
0!
0%
b110 *
0-
02
b110 6
#777410000000
1!
1%
1-
12
#777420000000
0!
0%
b111 *
0-
02
b111 6
#777430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#777440000000
0!
0%
b0 *
0-
02
b0 6
#777450000000
1!
1%
1-
12
#777460000000
0!
0%
b1 *
0-
02
b1 6
#777470000000
1!
1%
1-
12
#777480000000
0!
0%
b10 *
0-
02
b10 6
#777490000000
1!
1%
1-
12
#777500000000
0!
0%
b11 *
0-
02
b11 6
#777510000000
1!
1%
1-
12
15
#777520000000
0!
0%
b100 *
0-
02
b100 6
#777530000000
1!
1%
1-
12
#777540000000
0!
0%
b101 *
0-
02
b101 6
#777550000000
1!
1%
1-
12
#777560000000
0!
0%
b110 *
0-
02
b110 6
#777570000000
1!
1%
1-
12
#777580000000
0!
0%
b111 *
0-
02
b111 6
#777590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#777600000000
0!
0%
b0 *
0-
02
b0 6
#777610000000
1!
1%
1-
12
#777620000000
0!
0%
b1 *
0-
02
b1 6
#777630000000
1!
1%
1-
12
#777640000000
0!
0%
b10 *
0-
02
b10 6
#777650000000
1!
1%
1-
12
#777660000000
0!
0%
b11 *
0-
02
b11 6
#777670000000
1!
1%
1-
12
15
#777680000000
0!
0%
b100 *
0-
02
b100 6
#777690000000
1!
1%
1-
12
#777700000000
0!
0%
b101 *
0-
02
b101 6
#777710000000
1!
1%
1-
12
#777720000000
0!
0%
b110 *
0-
02
b110 6
#777730000000
1!
1%
1-
12
#777740000000
0!
0%
b111 *
0-
02
b111 6
#777750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#777760000000
0!
0%
b0 *
0-
02
b0 6
#777770000000
1!
1%
1-
12
#777780000000
0!
0%
b1 *
0-
02
b1 6
#777790000000
1!
1%
1-
12
#777800000000
0!
0%
b10 *
0-
02
b10 6
#777810000000
1!
1%
1-
12
#777820000000
0!
0%
b11 *
0-
02
b11 6
#777830000000
1!
1%
1-
12
15
#777840000000
0!
0%
b100 *
0-
02
b100 6
#777850000000
1!
1%
1-
12
#777860000000
0!
0%
b101 *
0-
02
b101 6
#777870000000
1!
1%
1-
12
#777880000000
0!
0%
b110 *
0-
02
b110 6
#777890000000
1!
1%
1-
12
#777900000000
0!
0%
b111 *
0-
02
b111 6
#777910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#777920000000
0!
0%
b0 *
0-
02
b0 6
#777930000000
1!
1%
1-
12
#777940000000
0!
0%
b1 *
0-
02
b1 6
#777950000000
1!
1%
1-
12
#777960000000
0!
0%
b10 *
0-
02
b10 6
#777970000000
1!
1%
1-
12
#777980000000
0!
0%
b11 *
0-
02
b11 6
#777990000000
1!
1%
1-
12
15
#778000000000
0!
0%
b100 *
0-
02
b100 6
#778010000000
1!
1%
1-
12
#778020000000
0!
0%
b101 *
0-
02
b101 6
#778030000000
1!
1%
1-
12
#778040000000
0!
0%
b110 *
0-
02
b110 6
#778050000000
1!
1%
1-
12
#778060000000
0!
0%
b111 *
0-
02
b111 6
#778070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#778080000000
0!
0%
b0 *
0-
02
b0 6
#778090000000
1!
1%
1-
12
#778100000000
0!
0%
b1 *
0-
02
b1 6
#778110000000
1!
1%
1-
12
#778120000000
0!
0%
b10 *
0-
02
b10 6
#778130000000
1!
1%
1-
12
#778140000000
0!
0%
b11 *
0-
02
b11 6
#778150000000
1!
1%
1-
12
15
#778160000000
0!
0%
b100 *
0-
02
b100 6
#778170000000
1!
1%
1-
12
#778180000000
0!
0%
b101 *
0-
02
b101 6
#778190000000
1!
1%
1-
12
#778200000000
0!
0%
b110 *
0-
02
b110 6
#778210000000
1!
1%
1-
12
#778220000000
0!
0%
b111 *
0-
02
b111 6
#778230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#778240000000
0!
0%
b0 *
0-
02
b0 6
#778250000000
1!
1%
1-
12
#778260000000
0!
0%
b1 *
0-
02
b1 6
#778270000000
1!
1%
1-
12
#778280000000
0!
0%
b10 *
0-
02
b10 6
#778290000000
1!
1%
1-
12
#778300000000
0!
0%
b11 *
0-
02
b11 6
#778310000000
1!
1%
1-
12
15
#778320000000
0!
0%
b100 *
0-
02
b100 6
#778330000000
1!
1%
1-
12
#778340000000
0!
0%
b101 *
0-
02
b101 6
#778350000000
1!
1%
1-
12
#778360000000
0!
0%
b110 *
0-
02
b110 6
#778370000000
1!
1%
1-
12
#778380000000
0!
0%
b111 *
0-
02
b111 6
#778390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#778400000000
0!
0%
b0 *
0-
02
b0 6
#778410000000
1!
1%
1-
12
#778420000000
0!
0%
b1 *
0-
02
b1 6
#778430000000
1!
1%
1-
12
#778440000000
0!
0%
b10 *
0-
02
b10 6
#778450000000
1!
1%
1-
12
#778460000000
0!
0%
b11 *
0-
02
b11 6
#778470000000
1!
1%
1-
12
15
#778480000000
0!
0%
b100 *
0-
02
b100 6
#778490000000
1!
1%
1-
12
#778500000000
0!
0%
b101 *
0-
02
b101 6
#778510000000
1!
1%
1-
12
#778520000000
0!
0%
b110 *
0-
02
b110 6
#778530000000
1!
1%
1-
12
#778540000000
0!
0%
b111 *
0-
02
b111 6
#778550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#778560000000
0!
0%
b0 *
0-
02
b0 6
#778570000000
1!
1%
1-
12
#778580000000
0!
0%
b1 *
0-
02
b1 6
#778590000000
1!
1%
1-
12
#778600000000
0!
0%
b10 *
0-
02
b10 6
#778610000000
1!
1%
1-
12
#778620000000
0!
0%
b11 *
0-
02
b11 6
#778630000000
1!
1%
1-
12
15
#778640000000
0!
0%
b100 *
0-
02
b100 6
#778650000000
1!
1%
1-
12
#778660000000
0!
0%
b101 *
0-
02
b101 6
#778670000000
1!
1%
1-
12
#778680000000
0!
0%
b110 *
0-
02
b110 6
#778690000000
1!
1%
1-
12
#778700000000
0!
0%
b111 *
0-
02
b111 6
#778710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#778720000000
0!
0%
b0 *
0-
02
b0 6
#778730000000
1!
1%
1-
12
#778740000000
0!
0%
b1 *
0-
02
b1 6
#778750000000
1!
1%
1-
12
#778760000000
0!
0%
b10 *
0-
02
b10 6
#778770000000
1!
1%
1-
12
#778780000000
0!
0%
b11 *
0-
02
b11 6
#778790000000
1!
1%
1-
12
15
#778800000000
0!
0%
b100 *
0-
02
b100 6
#778810000000
1!
1%
1-
12
#778820000000
0!
0%
b101 *
0-
02
b101 6
#778830000000
1!
1%
1-
12
#778840000000
0!
0%
b110 *
0-
02
b110 6
#778850000000
1!
1%
1-
12
#778860000000
0!
0%
b111 *
0-
02
b111 6
#778870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#778880000000
0!
0%
b0 *
0-
02
b0 6
#778890000000
1!
1%
1-
12
#778900000000
0!
0%
b1 *
0-
02
b1 6
#778910000000
1!
1%
1-
12
#778920000000
0!
0%
b10 *
0-
02
b10 6
#778930000000
1!
1%
1-
12
#778940000000
0!
0%
b11 *
0-
02
b11 6
#778950000000
1!
1%
1-
12
15
#778960000000
0!
0%
b100 *
0-
02
b100 6
#778970000000
1!
1%
1-
12
#778980000000
0!
0%
b101 *
0-
02
b101 6
#778990000000
1!
1%
1-
12
#779000000000
0!
0%
b110 *
0-
02
b110 6
#779010000000
1!
1%
1-
12
#779020000000
0!
0%
b111 *
0-
02
b111 6
#779030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#779040000000
0!
0%
b0 *
0-
02
b0 6
#779050000000
1!
1%
1-
12
#779060000000
0!
0%
b1 *
0-
02
b1 6
#779070000000
1!
1%
1-
12
#779080000000
0!
0%
b10 *
0-
02
b10 6
#779090000000
1!
1%
1-
12
#779100000000
0!
0%
b11 *
0-
02
b11 6
#779110000000
1!
1%
1-
12
15
#779120000000
0!
0%
b100 *
0-
02
b100 6
#779130000000
1!
1%
1-
12
#779140000000
0!
0%
b101 *
0-
02
b101 6
#779150000000
1!
1%
1-
12
#779160000000
0!
0%
b110 *
0-
02
b110 6
#779170000000
1!
1%
1-
12
#779180000000
0!
0%
b111 *
0-
02
b111 6
#779190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#779200000000
0!
0%
b0 *
0-
02
b0 6
#779210000000
1!
1%
1-
12
#779220000000
0!
0%
b1 *
0-
02
b1 6
#779230000000
1!
1%
1-
12
#779240000000
0!
0%
b10 *
0-
02
b10 6
#779250000000
1!
1%
1-
12
#779260000000
0!
0%
b11 *
0-
02
b11 6
#779270000000
1!
1%
1-
12
15
#779280000000
0!
0%
b100 *
0-
02
b100 6
#779290000000
1!
1%
1-
12
#779300000000
0!
0%
b101 *
0-
02
b101 6
#779310000000
1!
1%
1-
12
#779320000000
0!
0%
b110 *
0-
02
b110 6
#779330000000
1!
1%
1-
12
#779340000000
0!
0%
b111 *
0-
02
b111 6
#779350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#779360000000
0!
0%
b0 *
0-
02
b0 6
#779370000000
1!
1%
1-
12
#779380000000
0!
0%
b1 *
0-
02
b1 6
#779390000000
1!
1%
1-
12
#779400000000
0!
0%
b10 *
0-
02
b10 6
#779410000000
1!
1%
1-
12
#779420000000
0!
0%
b11 *
0-
02
b11 6
#779430000000
1!
1%
1-
12
15
#779440000000
0!
0%
b100 *
0-
02
b100 6
#779450000000
1!
1%
1-
12
#779460000000
0!
0%
b101 *
0-
02
b101 6
#779470000000
1!
1%
1-
12
#779480000000
0!
0%
b110 *
0-
02
b110 6
#779490000000
1!
1%
1-
12
#779500000000
0!
0%
b111 *
0-
02
b111 6
#779510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#779520000000
0!
0%
b0 *
0-
02
b0 6
#779530000000
1!
1%
1-
12
#779540000000
0!
0%
b1 *
0-
02
b1 6
#779550000000
1!
1%
1-
12
#779560000000
0!
0%
b10 *
0-
02
b10 6
#779570000000
1!
1%
1-
12
#779580000000
0!
0%
b11 *
0-
02
b11 6
#779590000000
1!
1%
1-
12
15
#779600000000
0!
0%
b100 *
0-
02
b100 6
#779610000000
1!
1%
1-
12
#779620000000
0!
0%
b101 *
0-
02
b101 6
#779630000000
1!
1%
1-
12
#779640000000
0!
0%
b110 *
0-
02
b110 6
#779650000000
1!
1%
1-
12
#779660000000
0!
0%
b111 *
0-
02
b111 6
#779670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#779680000000
0!
0%
b0 *
0-
02
b0 6
#779690000000
1!
1%
1-
12
#779700000000
0!
0%
b1 *
0-
02
b1 6
#779710000000
1!
1%
1-
12
#779720000000
0!
0%
b10 *
0-
02
b10 6
#779730000000
1!
1%
1-
12
#779740000000
0!
0%
b11 *
0-
02
b11 6
#779750000000
1!
1%
1-
12
15
#779760000000
0!
0%
b100 *
0-
02
b100 6
#779770000000
1!
1%
1-
12
#779780000000
0!
0%
b101 *
0-
02
b101 6
#779790000000
1!
1%
1-
12
#779800000000
0!
0%
b110 *
0-
02
b110 6
#779810000000
1!
1%
1-
12
#779820000000
0!
0%
b111 *
0-
02
b111 6
#779830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#779840000000
0!
0%
b0 *
0-
02
b0 6
#779850000000
1!
1%
1-
12
#779860000000
0!
0%
b1 *
0-
02
b1 6
#779870000000
1!
1%
1-
12
#779880000000
0!
0%
b10 *
0-
02
b10 6
#779890000000
1!
1%
1-
12
#779900000000
0!
0%
b11 *
0-
02
b11 6
#779910000000
1!
1%
1-
12
15
#779920000000
0!
0%
b100 *
0-
02
b100 6
#779930000000
1!
1%
1-
12
#779940000000
0!
0%
b101 *
0-
02
b101 6
#779950000000
1!
1%
1-
12
#779960000000
0!
0%
b110 *
0-
02
b110 6
#779970000000
1!
1%
1-
12
#779980000000
0!
0%
b111 *
0-
02
b111 6
#779990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#780000000000
0!
0%
b0 *
0-
02
b0 6
#780010000000
1!
1%
1-
12
#780020000000
0!
0%
b1 *
0-
02
b1 6
#780030000000
1!
1%
1-
12
#780040000000
0!
0%
b10 *
0-
02
b10 6
#780050000000
1!
1%
1-
12
#780060000000
0!
0%
b11 *
0-
02
b11 6
#780070000000
1!
1%
1-
12
15
#780080000000
0!
0%
b100 *
0-
02
b100 6
#780090000000
1!
1%
1-
12
#780100000000
0!
0%
b101 *
0-
02
b101 6
#780110000000
1!
1%
1-
12
#780120000000
0!
0%
b110 *
0-
02
b110 6
#780130000000
1!
1%
1-
12
#780140000000
0!
0%
b111 *
0-
02
b111 6
#780150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#780160000000
0!
0%
b0 *
0-
02
b0 6
#780170000000
1!
1%
1-
12
#780180000000
0!
0%
b1 *
0-
02
b1 6
#780190000000
1!
1%
1-
12
#780200000000
0!
0%
b10 *
0-
02
b10 6
#780210000000
1!
1%
1-
12
#780220000000
0!
0%
b11 *
0-
02
b11 6
#780230000000
1!
1%
1-
12
15
#780240000000
0!
0%
b100 *
0-
02
b100 6
#780250000000
1!
1%
1-
12
#780260000000
0!
0%
b101 *
0-
02
b101 6
#780270000000
1!
1%
1-
12
#780280000000
0!
0%
b110 *
0-
02
b110 6
#780290000000
1!
1%
1-
12
#780300000000
0!
0%
b111 *
0-
02
b111 6
#780310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#780320000000
0!
0%
b0 *
0-
02
b0 6
#780330000000
1!
1%
1-
12
#780340000000
0!
0%
b1 *
0-
02
b1 6
#780350000000
1!
1%
1-
12
#780360000000
0!
0%
b10 *
0-
02
b10 6
#780370000000
1!
1%
1-
12
#780380000000
0!
0%
b11 *
0-
02
b11 6
#780390000000
1!
1%
1-
12
15
#780400000000
0!
0%
b100 *
0-
02
b100 6
#780410000000
1!
1%
1-
12
#780420000000
0!
0%
b101 *
0-
02
b101 6
#780430000000
1!
1%
1-
12
#780440000000
0!
0%
b110 *
0-
02
b110 6
#780450000000
1!
1%
1-
12
#780460000000
0!
0%
b111 *
0-
02
b111 6
#780470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#780480000000
0!
0%
b0 *
0-
02
b0 6
#780490000000
1!
1%
1-
12
#780500000000
0!
0%
b1 *
0-
02
b1 6
#780510000000
1!
1%
1-
12
#780520000000
0!
0%
b10 *
0-
02
b10 6
#780530000000
1!
1%
1-
12
#780540000000
0!
0%
b11 *
0-
02
b11 6
#780550000000
1!
1%
1-
12
15
#780560000000
0!
0%
b100 *
0-
02
b100 6
#780570000000
1!
1%
1-
12
#780580000000
0!
0%
b101 *
0-
02
b101 6
#780590000000
1!
1%
1-
12
#780600000000
0!
0%
b110 *
0-
02
b110 6
#780610000000
1!
1%
1-
12
#780620000000
0!
0%
b111 *
0-
02
b111 6
#780630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#780640000000
0!
0%
b0 *
0-
02
b0 6
#780650000000
1!
1%
1-
12
#780660000000
0!
0%
b1 *
0-
02
b1 6
#780670000000
1!
1%
1-
12
#780680000000
0!
0%
b10 *
0-
02
b10 6
#780690000000
1!
1%
1-
12
#780700000000
0!
0%
b11 *
0-
02
b11 6
#780710000000
1!
1%
1-
12
15
#780720000000
0!
0%
b100 *
0-
02
b100 6
#780730000000
1!
1%
1-
12
#780740000000
0!
0%
b101 *
0-
02
b101 6
#780750000000
1!
1%
1-
12
#780760000000
0!
0%
b110 *
0-
02
b110 6
#780770000000
1!
1%
1-
12
#780780000000
0!
0%
b111 *
0-
02
b111 6
#780790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#780800000000
0!
0%
b0 *
0-
02
b0 6
#780810000000
1!
1%
1-
12
#780820000000
0!
0%
b1 *
0-
02
b1 6
#780830000000
1!
1%
1-
12
#780840000000
0!
0%
b10 *
0-
02
b10 6
#780850000000
1!
1%
1-
12
#780860000000
0!
0%
b11 *
0-
02
b11 6
#780870000000
1!
1%
1-
12
15
#780880000000
0!
0%
b100 *
0-
02
b100 6
#780890000000
1!
1%
1-
12
#780900000000
0!
0%
b101 *
0-
02
b101 6
#780910000000
1!
1%
1-
12
#780920000000
0!
0%
b110 *
0-
02
b110 6
#780930000000
1!
1%
1-
12
#780940000000
0!
0%
b111 *
0-
02
b111 6
#780950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#780960000000
0!
0%
b0 *
0-
02
b0 6
#780970000000
1!
1%
1-
12
#780980000000
0!
0%
b1 *
0-
02
b1 6
#780990000000
1!
1%
1-
12
#781000000000
0!
0%
b10 *
0-
02
b10 6
#781010000000
1!
1%
1-
12
#781020000000
0!
0%
b11 *
0-
02
b11 6
#781030000000
1!
1%
1-
12
15
#781040000000
0!
0%
b100 *
0-
02
b100 6
#781050000000
1!
1%
1-
12
#781060000000
0!
0%
b101 *
0-
02
b101 6
#781070000000
1!
1%
1-
12
#781080000000
0!
0%
b110 *
0-
02
b110 6
#781090000000
1!
1%
1-
12
#781100000000
0!
0%
b111 *
0-
02
b111 6
#781110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#781120000000
0!
0%
b0 *
0-
02
b0 6
#781130000000
1!
1%
1-
12
#781140000000
0!
0%
b1 *
0-
02
b1 6
#781150000000
1!
1%
1-
12
#781160000000
0!
0%
b10 *
0-
02
b10 6
#781170000000
1!
1%
1-
12
#781180000000
0!
0%
b11 *
0-
02
b11 6
#781190000000
1!
1%
1-
12
15
#781200000000
0!
0%
b100 *
0-
02
b100 6
#781210000000
1!
1%
1-
12
#781220000000
0!
0%
b101 *
0-
02
b101 6
#781230000000
1!
1%
1-
12
#781240000000
0!
0%
b110 *
0-
02
b110 6
#781250000000
1!
1%
1-
12
#781260000000
0!
0%
b111 *
0-
02
b111 6
#781270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#781280000000
0!
0%
b0 *
0-
02
b0 6
#781290000000
1!
1%
1-
12
#781300000000
0!
0%
b1 *
0-
02
b1 6
#781310000000
1!
1%
1-
12
#781320000000
0!
0%
b10 *
0-
02
b10 6
#781330000000
1!
1%
1-
12
#781340000000
0!
0%
b11 *
0-
02
b11 6
#781350000000
1!
1%
1-
12
15
#781360000000
0!
0%
b100 *
0-
02
b100 6
#781370000000
1!
1%
1-
12
#781380000000
0!
0%
b101 *
0-
02
b101 6
#781390000000
1!
1%
1-
12
#781400000000
0!
0%
b110 *
0-
02
b110 6
#781410000000
1!
1%
1-
12
#781420000000
0!
0%
b111 *
0-
02
b111 6
#781430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#781440000000
0!
0%
b0 *
0-
02
b0 6
#781450000000
1!
1%
1-
12
#781460000000
0!
0%
b1 *
0-
02
b1 6
#781470000000
1!
1%
1-
12
#781480000000
0!
0%
b10 *
0-
02
b10 6
#781490000000
1!
1%
1-
12
#781500000000
0!
0%
b11 *
0-
02
b11 6
#781510000000
1!
1%
1-
12
15
#781520000000
0!
0%
b100 *
0-
02
b100 6
#781530000000
1!
1%
1-
12
#781540000000
0!
0%
b101 *
0-
02
b101 6
#781550000000
1!
1%
1-
12
#781560000000
0!
0%
b110 *
0-
02
b110 6
#781570000000
1!
1%
1-
12
#781580000000
0!
0%
b111 *
0-
02
b111 6
#781590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#781600000000
0!
0%
b0 *
0-
02
b0 6
#781610000000
1!
1%
1-
12
#781620000000
0!
0%
b1 *
0-
02
b1 6
#781630000000
1!
1%
1-
12
#781640000000
0!
0%
b10 *
0-
02
b10 6
#781650000000
1!
1%
1-
12
#781660000000
0!
0%
b11 *
0-
02
b11 6
#781670000000
1!
1%
1-
12
15
#781680000000
0!
0%
b100 *
0-
02
b100 6
#781690000000
1!
1%
1-
12
#781700000000
0!
0%
b101 *
0-
02
b101 6
#781710000000
1!
1%
1-
12
#781720000000
0!
0%
b110 *
0-
02
b110 6
#781730000000
1!
1%
1-
12
#781740000000
0!
0%
b111 *
0-
02
b111 6
#781750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#781760000000
0!
0%
b0 *
0-
02
b0 6
#781770000000
1!
1%
1-
12
#781780000000
0!
0%
b1 *
0-
02
b1 6
#781790000000
1!
1%
1-
12
#781800000000
0!
0%
b10 *
0-
02
b10 6
#781810000000
1!
1%
1-
12
#781820000000
0!
0%
b11 *
0-
02
b11 6
#781830000000
1!
1%
1-
12
15
#781840000000
0!
0%
b100 *
0-
02
b100 6
#781850000000
1!
1%
1-
12
#781860000000
0!
0%
b101 *
0-
02
b101 6
#781870000000
1!
1%
1-
12
#781880000000
0!
0%
b110 *
0-
02
b110 6
#781890000000
1!
1%
1-
12
#781900000000
0!
0%
b111 *
0-
02
b111 6
#781910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#781920000000
0!
0%
b0 *
0-
02
b0 6
#781930000000
1!
1%
1-
12
#781940000000
0!
0%
b1 *
0-
02
b1 6
#781950000000
1!
1%
1-
12
#781960000000
0!
0%
b10 *
0-
02
b10 6
#781970000000
1!
1%
1-
12
#781980000000
0!
0%
b11 *
0-
02
b11 6
#781990000000
1!
1%
1-
12
15
#782000000000
0!
0%
b100 *
0-
02
b100 6
#782010000000
1!
1%
1-
12
#782020000000
0!
0%
b101 *
0-
02
b101 6
#782030000000
1!
1%
1-
12
#782040000000
0!
0%
b110 *
0-
02
b110 6
#782050000000
1!
1%
1-
12
#782060000000
0!
0%
b111 *
0-
02
b111 6
#782070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#782080000000
0!
0%
b0 *
0-
02
b0 6
#782090000000
1!
1%
1-
12
#782100000000
0!
0%
b1 *
0-
02
b1 6
#782110000000
1!
1%
1-
12
#782120000000
0!
0%
b10 *
0-
02
b10 6
#782130000000
1!
1%
1-
12
#782140000000
0!
0%
b11 *
0-
02
b11 6
#782150000000
1!
1%
1-
12
15
#782160000000
0!
0%
b100 *
0-
02
b100 6
#782170000000
1!
1%
1-
12
#782180000000
0!
0%
b101 *
0-
02
b101 6
#782190000000
1!
1%
1-
12
#782200000000
0!
0%
b110 *
0-
02
b110 6
#782210000000
1!
1%
1-
12
#782220000000
0!
0%
b111 *
0-
02
b111 6
#782230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#782240000000
0!
0%
b0 *
0-
02
b0 6
#782250000000
1!
1%
1-
12
#782260000000
0!
0%
b1 *
0-
02
b1 6
#782270000000
1!
1%
1-
12
#782280000000
0!
0%
b10 *
0-
02
b10 6
#782290000000
1!
1%
1-
12
#782300000000
0!
0%
b11 *
0-
02
b11 6
#782310000000
1!
1%
1-
12
15
#782320000000
0!
0%
b100 *
0-
02
b100 6
#782330000000
1!
1%
1-
12
#782340000000
0!
0%
b101 *
0-
02
b101 6
#782350000000
1!
1%
1-
12
#782360000000
0!
0%
b110 *
0-
02
b110 6
#782370000000
1!
1%
1-
12
#782380000000
0!
0%
b111 *
0-
02
b111 6
#782390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#782400000000
0!
0%
b0 *
0-
02
b0 6
#782410000000
1!
1%
1-
12
#782420000000
0!
0%
b1 *
0-
02
b1 6
#782430000000
1!
1%
1-
12
#782440000000
0!
0%
b10 *
0-
02
b10 6
#782450000000
1!
1%
1-
12
#782460000000
0!
0%
b11 *
0-
02
b11 6
#782470000000
1!
1%
1-
12
15
#782480000000
0!
0%
b100 *
0-
02
b100 6
#782490000000
1!
1%
1-
12
#782500000000
0!
0%
b101 *
0-
02
b101 6
#782510000000
1!
1%
1-
12
#782520000000
0!
0%
b110 *
0-
02
b110 6
#782530000000
1!
1%
1-
12
#782540000000
0!
0%
b111 *
0-
02
b111 6
#782550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#782560000000
0!
0%
b0 *
0-
02
b0 6
#782570000000
1!
1%
1-
12
#782580000000
0!
0%
b1 *
0-
02
b1 6
#782590000000
1!
1%
1-
12
#782600000000
0!
0%
b10 *
0-
02
b10 6
#782610000000
1!
1%
1-
12
#782620000000
0!
0%
b11 *
0-
02
b11 6
#782630000000
1!
1%
1-
12
15
#782640000000
0!
0%
b100 *
0-
02
b100 6
#782650000000
1!
1%
1-
12
#782660000000
0!
0%
b101 *
0-
02
b101 6
#782670000000
1!
1%
1-
12
#782680000000
0!
0%
b110 *
0-
02
b110 6
#782690000000
1!
1%
1-
12
#782700000000
0!
0%
b111 *
0-
02
b111 6
#782710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#782720000000
0!
0%
b0 *
0-
02
b0 6
#782730000000
1!
1%
1-
12
#782740000000
0!
0%
b1 *
0-
02
b1 6
#782750000000
1!
1%
1-
12
#782760000000
0!
0%
b10 *
0-
02
b10 6
#782770000000
1!
1%
1-
12
#782780000000
0!
0%
b11 *
0-
02
b11 6
#782790000000
1!
1%
1-
12
15
#782800000000
0!
0%
b100 *
0-
02
b100 6
#782810000000
1!
1%
1-
12
#782820000000
0!
0%
b101 *
0-
02
b101 6
#782830000000
1!
1%
1-
12
#782840000000
0!
0%
b110 *
0-
02
b110 6
#782850000000
1!
1%
1-
12
#782860000000
0!
0%
b111 *
0-
02
b111 6
#782870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#782880000000
0!
0%
b0 *
0-
02
b0 6
#782890000000
1!
1%
1-
12
#782900000000
0!
0%
b1 *
0-
02
b1 6
#782910000000
1!
1%
1-
12
#782920000000
0!
0%
b10 *
0-
02
b10 6
#782930000000
1!
1%
1-
12
#782940000000
0!
0%
b11 *
0-
02
b11 6
#782950000000
1!
1%
1-
12
15
#782960000000
0!
0%
b100 *
0-
02
b100 6
#782970000000
1!
1%
1-
12
#782980000000
0!
0%
b101 *
0-
02
b101 6
#782990000000
1!
1%
1-
12
#783000000000
0!
0%
b110 *
0-
02
b110 6
#783010000000
1!
1%
1-
12
#783020000000
0!
0%
b111 *
0-
02
b111 6
#783030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#783040000000
0!
0%
b0 *
0-
02
b0 6
#783050000000
1!
1%
1-
12
#783060000000
0!
0%
b1 *
0-
02
b1 6
#783070000000
1!
1%
1-
12
#783080000000
0!
0%
b10 *
0-
02
b10 6
#783090000000
1!
1%
1-
12
#783100000000
0!
0%
b11 *
0-
02
b11 6
#783110000000
1!
1%
1-
12
15
#783120000000
0!
0%
b100 *
0-
02
b100 6
#783130000000
1!
1%
1-
12
#783140000000
0!
0%
b101 *
0-
02
b101 6
#783150000000
1!
1%
1-
12
#783160000000
0!
0%
b110 *
0-
02
b110 6
#783170000000
1!
1%
1-
12
#783180000000
0!
0%
b111 *
0-
02
b111 6
#783190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#783200000000
0!
0%
b0 *
0-
02
b0 6
#783210000000
1!
1%
1-
12
#783220000000
0!
0%
b1 *
0-
02
b1 6
#783230000000
1!
1%
1-
12
#783240000000
0!
0%
b10 *
0-
02
b10 6
#783250000000
1!
1%
1-
12
#783260000000
0!
0%
b11 *
0-
02
b11 6
#783270000000
1!
1%
1-
12
15
#783280000000
0!
0%
b100 *
0-
02
b100 6
#783290000000
1!
1%
1-
12
#783300000000
0!
0%
b101 *
0-
02
b101 6
#783310000000
1!
1%
1-
12
#783320000000
0!
0%
b110 *
0-
02
b110 6
#783330000000
1!
1%
1-
12
#783340000000
0!
0%
b111 *
0-
02
b111 6
#783350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#783360000000
0!
0%
b0 *
0-
02
b0 6
#783370000000
1!
1%
1-
12
#783380000000
0!
0%
b1 *
0-
02
b1 6
#783390000000
1!
1%
1-
12
#783400000000
0!
0%
b10 *
0-
02
b10 6
#783410000000
1!
1%
1-
12
#783420000000
0!
0%
b11 *
0-
02
b11 6
#783430000000
1!
1%
1-
12
15
#783440000000
0!
0%
b100 *
0-
02
b100 6
#783450000000
1!
1%
1-
12
#783460000000
0!
0%
b101 *
0-
02
b101 6
#783470000000
1!
1%
1-
12
#783480000000
0!
0%
b110 *
0-
02
b110 6
#783490000000
1!
1%
1-
12
#783500000000
0!
0%
b111 *
0-
02
b111 6
#783510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#783520000000
0!
0%
b0 *
0-
02
b0 6
#783530000000
1!
1%
1-
12
#783540000000
0!
0%
b1 *
0-
02
b1 6
#783550000000
1!
1%
1-
12
#783560000000
0!
0%
b10 *
0-
02
b10 6
#783570000000
1!
1%
1-
12
#783580000000
0!
0%
b11 *
0-
02
b11 6
#783590000000
1!
1%
1-
12
15
#783600000000
0!
0%
b100 *
0-
02
b100 6
#783610000000
1!
1%
1-
12
#783620000000
0!
0%
b101 *
0-
02
b101 6
#783630000000
1!
1%
1-
12
#783640000000
0!
0%
b110 *
0-
02
b110 6
#783650000000
1!
1%
1-
12
#783660000000
0!
0%
b111 *
0-
02
b111 6
#783670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#783680000000
0!
0%
b0 *
0-
02
b0 6
#783690000000
1!
1%
1-
12
#783700000000
0!
0%
b1 *
0-
02
b1 6
#783710000000
1!
1%
1-
12
#783720000000
0!
0%
b10 *
0-
02
b10 6
#783730000000
1!
1%
1-
12
#783740000000
0!
0%
b11 *
0-
02
b11 6
#783750000000
1!
1%
1-
12
15
#783760000000
0!
0%
b100 *
0-
02
b100 6
#783770000000
1!
1%
1-
12
#783780000000
0!
0%
b101 *
0-
02
b101 6
#783790000000
1!
1%
1-
12
#783800000000
0!
0%
b110 *
0-
02
b110 6
#783810000000
1!
1%
1-
12
#783820000000
0!
0%
b111 *
0-
02
b111 6
#783830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#783840000000
0!
0%
b0 *
0-
02
b0 6
#783850000000
1!
1%
1-
12
#783860000000
0!
0%
b1 *
0-
02
b1 6
#783870000000
1!
1%
1-
12
#783880000000
0!
0%
b10 *
0-
02
b10 6
#783890000000
1!
1%
1-
12
#783900000000
0!
0%
b11 *
0-
02
b11 6
#783910000000
1!
1%
1-
12
15
#783920000000
0!
0%
b100 *
0-
02
b100 6
#783930000000
1!
1%
1-
12
#783940000000
0!
0%
b101 *
0-
02
b101 6
#783950000000
1!
1%
1-
12
#783960000000
0!
0%
b110 *
0-
02
b110 6
#783970000000
1!
1%
1-
12
#783980000000
0!
0%
b111 *
0-
02
b111 6
#783990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#784000000000
0!
0%
b0 *
0-
02
b0 6
#784010000000
1!
1%
1-
12
#784020000000
0!
0%
b1 *
0-
02
b1 6
#784030000000
1!
1%
1-
12
#784040000000
0!
0%
b10 *
0-
02
b10 6
#784050000000
1!
1%
1-
12
#784060000000
0!
0%
b11 *
0-
02
b11 6
#784070000000
1!
1%
1-
12
15
#784080000000
0!
0%
b100 *
0-
02
b100 6
#784090000000
1!
1%
1-
12
#784100000000
0!
0%
b101 *
0-
02
b101 6
#784110000000
1!
1%
1-
12
#784120000000
0!
0%
b110 *
0-
02
b110 6
#784130000000
1!
1%
1-
12
#784140000000
0!
0%
b111 *
0-
02
b111 6
#784150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#784160000000
0!
0%
b0 *
0-
02
b0 6
#784170000000
1!
1%
1-
12
#784180000000
0!
0%
b1 *
0-
02
b1 6
#784190000000
1!
1%
1-
12
#784200000000
0!
0%
b10 *
0-
02
b10 6
#784210000000
1!
1%
1-
12
#784220000000
0!
0%
b11 *
0-
02
b11 6
#784230000000
1!
1%
1-
12
15
#784240000000
0!
0%
b100 *
0-
02
b100 6
#784250000000
1!
1%
1-
12
#784260000000
0!
0%
b101 *
0-
02
b101 6
#784270000000
1!
1%
1-
12
#784280000000
0!
0%
b110 *
0-
02
b110 6
#784290000000
1!
1%
1-
12
#784300000000
0!
0%
b111 *
0-
02
b111 6
#784310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#784320000000
0!
0%
b0 *
0-
02
b0 6
#784330000000
1!
1%
1-
12
#784340000000
0!
0%
b1 *
0-
02
b1 6
#784350000000
1!
1%
1-
12
#784360000000
0!
0%
b10 *
0-
02
b10 6
#784370000000
1!
1%
1-
12
#784380000000
0!
0%
b11 *
0-
02
b11 6
#784390000000
1!
1%
1-
12
15
#784400000000
0!
0%
b100 *
0-
02
b100 6
#784410000000
1!
1%
1-
12
#784420000000
0!
0%
b101 *
0-
02
b101 6
#784430000000
1!
1%
1-
12
#784440000000
0!
0%
b110 *
0-
02
b110 6
#784450000000
1!
1%
1-
12
#784460000000
0!
0%
b111 *
0-
02
b111 6
#784470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#784480000000
0!
0%
b0 *
0-
02
b0 6
#784490000000
1!
1%
1-
12
#784500000000
0!
0%
b1 *
0-
02
b1 6
#784510000000
1!
1%
1-
12
#784520000000
0!
0%
b10 *
0-
02
b10 6
#784530000000
1!
1%
1-
12
#784540000000
0!
0%
b11 *
0-
02
b11 6
#784550000000
1!
1%
1-
12
15
#784560000000
0!
0%
b100 *
0-
02
b100 6
#784570000000
1!
1%
1-
12
#784580000000
0!
0%
b101 *
0-
02
b101 6
#784590000000
1!
1%
1-
12
#784600000000
0!
0%
b110 *
0-
02
b110 6
#784610000000
1!
1%
1-
12
#784620000000
0!
0%
b111 *
0-
02
b111 6
#784630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#784640000000
0!
0%
b0 *
0-
02
b0 6
#784650000000
1!
1%
1-
12
#784660000000
0!
0%
b1 *
0-
02
b1 6
#784670000000
1!
1%
1-
12
#784680000000
0!
0%
b10 *
0-
02
b10 6
#784690000000
1!
1%
1-
12
#784700000000
0!
0%
b11 *
0-
02
b11 6
#784710000000
1!
1%
1-
12
15
#784720000000
0!
0%
b100 *
0-
02
b100 6
#784730000000
1!
1%
1-
12
#784740000000
0!
0%
b101 *
0-
02
b101 6
#784750000000
1!
1%
1-
12
#784760000000
0!
0%
b110 *
0-
02
b110 6
#784770000000
1!
1%
1-
12
#784780000000
0!
0%
b111 *
0-
02
b111 6
#784790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#784800000000
0!
0%
b0 *
0-
02
b0 6
#784810000000
1!
1%
1-
12
#784820000000
0!
0%
b1 *
0-
02
b1 6
#784830000000
1!
1%
1-
12
#784840000000
0!
0%
b10 *
0-
02
b10 6
#784850000000
1!
1%
1-
12
#784860000000
0!
0%
b11 *
0-
02
b11 6
#784870000000
1!
1%
1-
12
15
#784880000000
0!
0%
b100 *
0-
02
b100 6
#784890000000
1!
1%
1-
12
#784900000000
0!
0%
b101 *
0-
02
b101 6
#784910000000
1!
1%
1-
12
#784920000000
0!
0%
b110 *
0-
02
b110 6
#784930000000
1!
1%
1-
12
#784940000000
0!
0%
b111 *
0-
02
b111 6
#784950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#784960000000
0!
0%
b0 *
0-
02
b0 6
#784970000000
1!
1%
1-
12
#784980000000
0!
0%
b1 *
0-
02
b1 6
#784990000000
1!
1%
1-
12
#785000000000
0!
0%
b10 *
0-
02
b10 6
#785010000000
1!
1%
1-
12
#785020000000
0!
0%
b11 *
0-
02
b11 6
#785030000000
1!
1%
1-
12
15
#785040000000
0!
0%
b100 *
0-
02
b100 6
#785050000000
1!
1%
1-
12
#785060000000
0!
0%
b101 *
0-
02
b101 6
#785070000000
1!
1%
1-
12
#785080000000
0!
0%
b110 *
0-
02
b110 6
#785090000000
1!
1%
1-
12
#785100000000
0!
0%
b111 *
0-
02
b111 6
#785110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#785120000000
0!
0%
b0 *
0-
02
b0 6
#785130000000
1!
1%
1-
12
#785140000000
0!
0%
b1 *
0-
02
b1 6
#785150000000
1!
1%
1-
12
#785160000000
0!
0%
b10 *
0-
02
b10 6
#785170000000
1!
1%
1-
12
#785180000000
0!
0%
b11 *
0-
02
b11 6
#785190000000
1!
1%
1-
12
15
#785200000000
0!
0%
b100 *
0-
02
b100 6
#785210000000
1!
1%
1-
12
#785220000000
0!
0%
b101 *
0-
02
b101 6
#785230000000
1!
1%
1-
12
#785240000000
0!
0%
b110 *
0-
02
b110 6
#785250000000
1!
1%
1-
12
#785260000000
0!
0%
b111 *
0-
02
b111 6
#785270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#785280000000
0!
0%
b0 *
0-
02
b0 6
#785290000000
1!
1%
1-
12
#785300000000
0!
0%
b1 *
0-
02
b1 6
#785310000000
1!
1%
1-
12
#785320000000
0!
0%
b10 *
0-
02
b10 6
#785330000000
1!
1%
1-
12
#785340000000
0!
0%
b11 *
0-
02
b11 6
#785350000000
1!
1%
1-
12
15
#785360000000
0!
0%
b100 *
0-
02
b100 6
#785370000000
1!
1%
1-
12
#785380000000
0!
0%
b101 *
0-
02
b101 6
#785390000000
1!
1%
1-
12
#785400000000
0!
0%
b110 *
0-
02
b110 6
#785410000000
1!
1%
1-
12
#785420000000
0!
0%
b111 *
0-
02
b111 6
#785430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#785440000000
0!
0%
b0 *
0-
02
b0 6
#785450000000
1!
1%
1-
12
#785460000000
0!
0%
b1 *
0-
02
b1 6
#785470000000
1!
1%
1-
12
#785480000000
0!
0%
b10 *
0-
02
b10 6
#785490000000
1!
1%
1-
12
#785500000000
0!
0%
b11 *
0-
02
b11 6
#785510000000
1!
1%
1-
12
15
#785520000000
0!
0%
b100 *
0-
02
b100 6
#785530000000
1!
1%
1-
12
#785540000000
0!
0%
b101 *
0-
02
b101 6
#785550000000
1!
1%
1-
12
#785560000000
0!
0%
b110 *
0-
02
b110 6
#785570000000
1!
1%
1-
12
#785580000000
0!
0%
b111 *
0-
02
b111 6
#785590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#785600000000
0!
0%
b0 *
0-
02
b0 6
#785610000000
1!
1%
1-
12
#785620000000
0!
0%
b1 *
0-
02
b1 6
#785630000000
1!
1%
1-
12
#785640000000
0!
0%
b10 *
0-
02
b10 6
#785650000000
1!
1%
1-
12
#785660000000
0!
0%
b11 *
0-
02
b11 6
#785670000000
1!
1%
1-
12
15
#785680000000
0!
0%
b100 *
0-
02
b100 6
#785690000000
1!
1%
1-
12
#785700000000
0!
0%
b101 *
0-
02
b101 6
#785710000000
1!
1%
1-
12
#785720000000
0!
0%
b110 *
0-
02
b110 6
#785730000000
1!
1%
1-
12
#785740000000
0!
0%
b111 *
0-
02
b111 6
#785750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#785760000000
0!
0%
b0 *
0-
02
b0 6
#785770000000
1!
1%
1-
12
#785780000000
0!
0%
b1 *
0-
02
b1 6
#785790000000
1!
1%
1-
12
#785800000000
0!
0%
b10 *
0-
02
b10 6
#785810000000
1!
1%
1-
12
#785820000000
0!
0%
b11 *
0-
02
b11 6
#785830000000
1!
1%
1-
12
15
#785840000000
0!
0%
b100 *
0-
02
b100 6
#785850000000
1!
1%
1-
12
#785860000000
0!
0%
b101 *
0-
02
b101 6
#785870000000
1!
1%
1-
12
#785880000000
0!
0%
b110 *
0-
02
b110 6
#785890000000
1!
1%
1-
12
#785900000000
0!
0%
b111 *
0-
02
b111 6
#785910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#785920000000
0!
0%
b0 *
0-
02
b0 6
#785930000000
1!
1%
1-
12
#785940000000
0!
0%
b1 *
0-
02
b1 6
#785950000000
1!
1%
1-
12
#785960000000
0!
0%
b10 *
0-
02
b10 6
#785970000000
1!
1%
1-
12
#785980000000
0!
0%
b11 *
0-
02
b11 6
#785990000000
1!
1%
1-
12
15
#786000000000
0!
0%
b100 *
0-
02
b100 6
#786010000000
1!
1%
1-
12
#786020000000
0!
0%
b101 *
0-
02
b101 6
#786030000000
1!
1%
1-
12
#786040000000
0!
0%
b110 *
0-
02
b110 6
#786050000000
1!
1%
1-
12
#786060000000
0!
0%
b111 *
0-
02
b111 6
#786070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#786080000000
0!
0%
b0 *
0-
02
b0 6
#786090000000
1!
1%
1-
12
#786100000000
0!
0%
b1 *
0-
02
b1 6
#786110000000
1!
1%
1-
12
#786120000000
0!
0%
b10 *
0-
02
b10 6
#786130000000
1!
1%
1-
12
#786140000000
0!
0%
b11 *
0-
02
b11 6
#786150000000
1!
1%
1-
12
15
#786160000000
0!
0%
b100 *
0-
02
b100 6
#786170000000
1!
1%
1-
12
#786180000000
0!
0%
b101 *
0-
02
b101 6
#786190000000
1!
1%
1-
12
#786200000000
0!
0%
b110 *
0-
02
b110 6
#786210000000
1!
1%
1-
12
#786220000000
0!
0%
b111 *
0-
02
b111 6
#786230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#786240000000
0!
0%
b0 *
0-
02
b0 6
#786250000000
1!
1%
1-
12
#786260000000
0!
0%
b1 *
0-
02
b1 6
#786270000000
1!
1%
1-
12
#786280000000
0!
0%
b10 *
0-
02
b10 6
#786290000000
1!
1%
1-
12
#786300000000
0!
0%
b11 *
0-
02
b11 6
#786310000000
1!
1%
1-
12
15
#786320000000
0!
0%
b100 *
0-
02
b100 6
#786330000000
1!
1%
1-
12
#786340000000
0!
0%
b101 *
0-
02
b101 6
#786350000000
1!
1%
1-
12
#786360000000
0!
0%
b110 *
0-
02
b110 6
#786370000000
1!
1%
1-
12
#786380000000
0!
0%
b111 *
0-
02
b111 6
#786390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#786400000000
0!
0%
b0 *
0-
02
b0 6
#786410000000
1!
1%
1-
12
#786420000000
0!
0%
b1 *
0-
02
b1 6
#786430000000
1!
1%
1-
12
#786440000000
0!
0%
b10 *
0-
02
b10 6
#786450000000
1!
1%
1-
12
#786460000000
0!
0%
b11 *
0-
02
b11 6
#786470000000
1!
1%
1-
12
15
#786480000000
0!
0%
b100 *
0-
02
b100 6
#786490000000
1!
1%
1-
12
#786500000000
0!
0%
b101 *
0-
02
b101 6
#786510000000
1!
1%
1-
12
#786520000000
0!
0%
b110 *
0-
02
b110 6
#786530000000
1!
1%
1-
12
#786540000000
0!
0%
b111 *
0-
02
b111 6
#786550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#786560000000
0!
0%
b0 *
0-
02
b0 6
#786570000000
1!
1%
1-
12
#786580000000
0!
0%
b1 *
0-
02
b1 6
#786590000000
1!
1%
1-
12
#786600000000
0!
0%
b10 *
0-
02
b10 6
#786610000000
1!
1%
1-
12
#786620000000
0!
0%
b11 *
0-
02
b11 6
#786630000000
1!
1%
1-
12
15
#786640000000
0!
0%
b100 *
0-
02
b100 6
#786650000000
1!
1%
1-
12
#786660000000
0!
0%
b101 *
0-
02
b101 6
#786670000000
1!
1%
1-
12
#786680000000
0!
0%
b110 *
0-
02
b110 6
#786690000000
1!
1%
1-
12
#786700000000
0!
0%
b111 *
0-
02
b111 6
#786710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#786720000000
0!
0%
b0 *
0-
02
b0 6
#786730000000
1!
1%
1-
12
#786740000000
0!
0%
b1 *
0-
02
b1 6
#786750000000
1!
1%
1-
12
#786760000000
0!
0%
b10 *
0-
02
b10 6
#786770000000
1!
1%
1-
12
#786780000000
0!
0%
b11 *
0-
02
b11 6
#786790000000
1!
1%
1-
12
15
#786800000000
0!
0%
b100 *
0-
02
b100 6
#786810000000
1!
1%
1-
12
#786820000000
0!
0%
b101 *
0-
02
b101 6
#786830000000
1!
1%
1-
12
#786840000000
0!
0%
b110 *
0-
02
b110 6
#786850000000
1!
1%
1-
12
#786860000000
0!
0%
b111 *
0-
02
b111 6
#786870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#786880000000
0!
0%
b0 *
0-
02
b0 6
#786890000000
1!
1%
1-
12
#786900000000
0!
0%
b1 *
0-
02
b1 6
#786910000000
1!
1%
1-
12
#786920000000
0!
0%
b10 *
0-
02
b10 6
#786930000000
1!
1%
1-
12
#786940000000
0!
0%
b11 *
0-
02
b11 6
#786950000000
1!
1%
1-
12
15
#786960000000
0!
0%
b100 *
0-
02
b100 6
#786970000000
1!
1%
1-
12
#786980000000
0!
0%
b101 *
0-
02
b101 6
#786990000000
1!
1%
1-
12
#787000000000
0!
0%
b110 *
0-
02
b110 6
#787010000000
1!
1%
1-
12
#787020000000
0!
0%
b111 *
0-
02
b111 6
#787030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#787040000000
0!
0%
b0 *
0-
02
b0 6
#787050000000
1!
1%
1-
12
#787060000000
0!
0%
b1 *
0-
02
b1 6
#787070000000
1!
1%
1-
12
#787080000000
0!
0%
b10 *
0-
02
b10 6
#787090000000
1!
1%
1-
12
#787100000000
0!
0%
b11 *
0-
02
b11 6
#787110000000
1!
1%
1-
12
15
#787120000000
0!
0%
b100 *
0-
02
b100 6
#787130000000
1!
1%
1-
12
#787140000000
0!
0%
b101 *
0-
02
b101 6
#787150000000
1!
1%
1-
12
#787160000000
0!
0%
b110 *
0-
02
b110 6
#787170000000
1!
1%
1-
12
#787180000000
0!
0%
b111 *
0-
02
b111 6
#787190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#787200000000
0!
0%
b0 *
0-
02
b0 6
#787210000000
1!
1%
1-
12
#787220000000
0!
0%
b1 *
0-
02
b1 6
#787230000000
1!
1%
1-
12
#787240000000
0!
0%
b10 *
0-
02
b10 6
#787250000000
1!
1%
1-
12
#787260000000
0!
0%
b11 *
0-
02
b11 6
#787270000000
1!
1%
1-
12
15
#787280000000
0!
0%
b100 *
0-
02
b100 6
#787290000000
1!
1%
1-
12
#787300000000
0!
0%
b101 *
0-
02
b101 6
#787310000000
1!
1%
1-
12
#787320000000
0!
0%
b110 *
0-
02
b110 6
#787330000000
1!
1%
1-
12
#787340000000
0!
0%
b111 *
0-
02
b111 6
#787350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#787360000000
0!
0%
b0 *
0-
02
b0 6
#787370000000
1!
1%
1-
12
#787380000000
0!
0%
b1 *
0-
02
b1 6
#787390000000
1!
1%
1-
12
#787400000000
0!
0%
b10 *
0-
02
b10 6
#787410000000
1!
1%
1-
12
#787420000000
0!
0%
b11 *
0-
02
b11 6
#787430000000
1!
1%
1-
12
15
#787440000000
0!
0%
b100 *
0-
02
b100 6
#787450000000
1!
1%
1-
12
#787460000000
0!
0%
b101 *
0-
02
b101 6
#787470000000
1!
1%
1-
12
#787480000000
0!
0%
b110 *
0-
02
b110 6
#787490000000
1!
1%
1-
12
#787500000000
0!
0%
b111 *
0-
02
b111 6
#787510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#787520000000
0!
0%
b0 *
0-
02
b0 6
#787530000000
1!
1%
1-
12
#787540000000
0!
0%
b1 *
0-
02
b1 6
#787550000000
1!
1%
1-
12
#787560000000
0!
0%
b10 *
0-
02
b10 6
#787570000000
1!
1%
1-
12
#787580000000
0!
0%
b11 *
0-
02
b11 6
#787590000000
1!
1%
1-
12
15
#787600000000
0!
0%
b100 *
0-
02
b100 6
#787610000000
1!
1%
1-
12
#787620000000
0!
0%
b101 *
0-
02
b101 6
#787630000000
1!
1%
1-
12
#787640000000
0!
0%
b110 *
0-
02
b110 6
#787650000000
1!
1%
1-
12
#787660000000
0!
0%
b111 *
0-
02
b111 6
#787670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#787680000000
0!
0%
b0 *
0-
02
b0 6
#787690000000
1!
1%
1-
12
#787700000000
0!
0%
b1 *
0-
02
b1 6
#787710000000
1!
1%
1-
12
#787720000000
0!
0%
b10 *
0-
02
b10 6
#787730000000
1!
1%
1-
12
#787740000000
0!
0%
b11 *
0-
02
b11 6
#787750000000
1!
1%
1-
12
15
#787760000000
0!
0%
b100 *
0-
02
b100 6
#787770000000
1!
1%
1-
12
#787780000000
0!
0%
b101 *
0-
02
b101 6
#787790000000
1!
1%
1-
12
#787800000000
0!
0%
b110 *
0-
02
b110 6
#787810000000
1!
1%
1-
12
#787820000000
0!
0%
b111 *
0-
02
b111 6
#787830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#787840000000
0!
0%
b0 *
0-
02
b0 6
#787850000000
1!
1%
1-
12
#787860000000
0!
0%
b1 *
0-
02
b1 6
#787870000000
1!
1%
1-
12
#787880000000
0!
0%
b10 *
0-
02
b10 6
#787890000000
1!
1%
1-
12
#787900000000
0!
0%
b11 *
0-
02
b11 6
#787910000000
1!
1%
1-
12
15
#787920000000
0!
0%
b100 *
0-
02
b100 6
#787930000000
1!
1%
1-
12
#787940000000
0!
0%
b101 *
0-
02
b101 6
#787950000000
1!
1%
1-
12
#787960000000
0!
0%
b110 *
0-
02
b110 6
#787970000000
1!
1%
1-
12
#787980000000
0!
0%
b111 *
0-
02
b111 6
#787990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#788000000000
0!
0%
b0 *
0-
02
b0 6
#788010000000
1!
1%
1-
12
#788020000000
0!
0%
b1 *
0-
02
b1 6
#788030000000
1!
1%
1-
12
#788040000000
0!
0%
b10 *
0-
02
b10 6
#788050000000
1!
1%
1-
12
#788060000000
0!
0%
b11 *
0-
02
b11 6
#788070000000
1!
1%
1-
12
15
#788080000000
0!
0%
b100 *
0-
02
b100 6
#788090000000
1!
1%
1-
12
#788100000000
0!
0%
b101 *
0-
02
b101 6
#788110000000
1!
1%
1-
12
#788120000000
0!
0%
b110 *
0-
02
b110 6
#788130000000
1!
1%
1-
12
#788140000000
0!
0%
b111 *
0-
02
b111 6
#788150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#788160000000
0!
0%
b0 *
0-
02
b0 6
#788170000000
1!
1%
1-
12
#788180000000
0!
0%
b1 *
0-
02
b1 6
#788190000000
1!
1%
1-
12
#788200000000
0!
0%
b10 *
0-
02
b10 6
#788210000000
1!
1%
1-
12
#788220000000
0!
0%
b11 *
0-
02
b11 6
#788230000000
1!
1%
1-
12
15
#788240000000
0!
0%
b100 *
0-
02
b100 6
#788250000000
1!
1%
1-
12
#788260000000
0!
0%
b101 *
0-
02
b101 6
#788270000000
1!
1%
1-
12
#788280000000
0!
0%
b110 *
0-
02
b110 6
#788290000000
1!
1%
1-
12
#788300000000
0!
0%
b111 *
0-
02
b111 6
#788310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#788320000000
0!
0%
b0 *
0-
02
b0 6
#788330000000
1!
1%
1-
12
#788340000000
0!
0%
b1 *
0-
02
b1 6
#788350000000
1!
1%
1-
12
#788360000000
0!
0%
b10 *
0-
02
b10 6
#788370000000
1!
1%
1-
12
#788380000000
0!
0%
b11 *
0-
02
b11 6
#788390000000
1!
1%
1-
12
15
#788400000000
0!
0%
b100 *
0-
02
b100 6
#788410000000
1!
1%
1-
12
#788420000000
0!
0%
b101 *
0-
02
b101 6
#788430000000
1!
1%
1-
12
#788440000000
0!
0%
b110 *
0-
02
b110 6
#788450000000
1!
1%
1-
12
#788460000000
0!
0%
b111 *
0-
02
b111 6
#788470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#788480000000
0!
0%
b0 *
0-
02
b0 6
#788490000000
1!
1%
1-
12
#788500000000
0!
0%
b1 *
0-
02
b1 6
#788510000000
1!
1%
1-
12
#788520000000
0!
0%
b10 *
0-
02
b10 6
#788530000000
1!
1%
1-
12
#788540000000
0!
0%
b11 *
0-
02
b11 6
#788550000000
1!
1%
1-
12
15
#788560000000
0!
0%
b100 *
0-
02
b100 6
#788570000000
1!
1%
1-
12
#788580000000
0!
0%
b101 *
0-
02
b101 6
#788590000000
1!
1%
1-
12
#788600000000
0!
0%
b110 *
0-
02
b110 6
#788610000000
1!
1%
1-
12
#788620000000
0!
0%
b111 *
0-
02
b111 6
#788630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#788640000000
0!
0%
b0 *
0-
02
b0 6
#788650000000
1!
1%
1-
12
#788660000000
0!
0%
b1 *
0-
02
b1 6
#788670000000
1!
1%
1-
12
#788680000000
0!
0%
b10 *
0-
02
b10 6
#788690000000
1!
1%
1-
12
#788700000000
0!
0%
b11 *
0-
02
b11 6
#788710000000
1!
1%
1-
12
15
#788720000000
0!
0%
b100 *
0-
02
b100 6
#788730000000
1!
1%
1-
12
#788740000000
0!
0%
b101 *
0-
02
b101 6
#788750000000
1!
1%
1-
12
#788760000000
0!
0%
b110 *
0-
02
b110 6
#788770000000
1!
1%
1-
12
#788780000000
0!
0%
b111 *
0-
02
b111 6
#788790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#788800000000
0!
0%
b0 *
0-
02
b0 6
#788810000000
1!
1%
1-
12
#788820000000
0!
0%
b1 *
0-
02
b1 6
#788830000000
1!
1%
1-
12
#788840000000
0!
0%
b10 *
0-
02
b10 6
#788850000000
1!
1%
1-
12
#788860000000
0!
0%
b11 *
0-
02
b11 6
#788870000000
1!
1%
1-
12
15
#788880000000
0!
0%
b100 *
0-
02
b100 6
#788890000000
1!
1%
1-
12
#788900000000
0!
0%
b101 *
0-
02
b101 6
#788910000000
1!
1%
1-
12
#788920000000
0!
0%
b110 *
0-
02
b110 6
#788930000000
1!
1%
1-
12
#788940000000
0!
0%
b111 *
0-
02
b111 6
#788950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#788960000000
0!
0%
b0 *
0-
02
b0 6
#788970000000
1!
1%
1-
12
#788980000000
0!
0%
b1 *
0-
02
b1 6
#788990000000
1!
1%
1-
12
#789000000000
0!
0%
b10 *
0-
02
b10 6
#789010000000
1!
1%
1-
12
#789020000000
0!
0%
b11 *
0-
02
b11 6
#789030000000
1!
1%
1-
12
15
#789040000000
0!
0%
b100 *
0-
02
b100 6
#789050000000
1!
1%
1-
12
#789060000000
0!
0%
b101 *
0-
02
b101 6
#789070000000
1!
1%
1-
12
#789080000000
0!
0%
b110 *
0-
02
b110 6
#789090000000
1!
1%
1-
12
#789100000000
0!
0%
b111 *
0-
02
b111 6
#789110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#789120000000
0!
0%
b0 *
0-
02
b0 6
#789130000000
1!
1%
1-
12
#789140000000
0!
0%
b1 *
0-
02
b1 6
#789150000000
1!
1%
1-
12
#789160000000
0!
0%
b10 *
0-
02
b10 6
#789170000000
1!
1%
1-
12
#789180000000
0!
0%
b11 *
0-
02
b11 6
#789190000000
1!
1%
1-
12
15
#789200000000
0!
0%
b100 *
0-
02
b100 6
#789210000000
1!
1%
1-
12
#789220000000
0!
0%
b101 *
0-
02
b101 6
#789230000000
1!
1%
1-
12
#789240000000
0!
0%
b110 *
0-
02
b110 6
#789250000000
1!
1%
1-
12
#789260000000
0!
0%
b111 *
0-
02
b111 6
#789270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#789280000000
0!
0%
b0 *
0-
02
b0 6
#789290000000
1!
1%
1-
12
#789300000000
0!
0%
b1 *
0-
02
b1 6
#789310000000
1!
1%
1-
12
#789320000000
0!
0%
b10 *
0-
02
b10 6
#789330000000
1!
1%
1-
12
#789340000000
0!
0%
b11 *
0-
02
b11 6
#789350000000
1!
1%
1-
12
15
#789360000000
0!
0%
b100 *
0-
02
b100 6
#789370000000
1!
1%
1-
12
#789380000000
0!
0%
b101 *
0-
02
b101 6
#789390000000
1!
1%
1-
12
#789400000000
0!
0%
b110 *
0-
02
b110 6
#789410000000
1!
1%
1-
12
#789420000000
0!
0%
b111 *
0-
02
b111 6
#789430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#789440000000
0!
0%
b0 *
0-
02
b0 6
#789450000000
1!
1%
1-
12
#789460000000
0!
0%
b1 *
0-
02
b1 6
#789470000000
1!
1%
1-
12
#789480000000
0!
0%
b10 *
0-
02
b10 6
#789490000000
1!
1%
1-
12
#789500000000
0!
0%
b11 *
0-
02
b11 6
#789510000000
1!
1%
1-
12
15
#789520000000
0!
0%
b100 *
0-
02
b100 6
#789530000000
1!
1%
1-
12
#789540000000
0!
0%
b101 *
0-
02
b101 6
#789550000000
1!
1%
1-
12
#789560000000
0!
0%
b110 *
0-
02
b110 6
#789570000000
1!
1%
1-
12
#789580000000
0!
0%
b111 *
0-
02
b111 6
#789590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#789600000000
0!
0%
b0 *
0-
02
b0 6
#789610000000
1!
1%
1-
12
#789620000000
0!
0%
b1 *
0-
02
b1 6
#789630000000
1!
1%
1-
12
#789640000000
0!
0%
b10 *
0-
02
b10 6
#789650000000
1!
1%
1-
12
#789660000000
0!
0%
b11 *
0-
02
b11 6
#789670000000
1!
1%
1-
12
15
#789680000000
0!
0%
b100 *
0-
02
b100 6
#789690000000
1!
1%
1-
12
#789700000000
0!
0%
b101 *
0-
02
b101 6
#789710000000
1!
1%
1-
12
#789720000000
0!
0%
b110 *
0-
02
b110 6
#789730000000
1!
1%
1-
12
#789740000000
0!
0%
b111 *
0-
02
b111 6
#789750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#789760000000
0!
0%
b0 *
0-
02
b0 6
#789770000000
1!
1%
1-
12
#789780000000
0!
0%
b1 *
0-
02
b1 6
#789790000000
1!
1%
1-
12
#789800000000
0!
0%
b10 *
0-
02
b10 6
#789810000000
1!
1%
1-
12
#789820000000
0!
0%
b11 *
0-
02
b11 6
#789830000000
1!
1%
1-
12
15
#789840000000
0!
0%
b100 *
0-
02
b100 6
#789850000000
1!
1%
1-
12
#789860000000
0!
0%
b101 *
0-
02
b101 6
#789870000000
1!
1%
1-
12
#789880000000
0!
0%
b110 *
0-
02
b110 6
#789890000000
1!
1%
1-
12
#789900000000
0!
0%
b111 *
0-
02
b111 6
#789910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#789920000000
0!
0%
b0 *
0-
02
b0 6
#789930000000
1!
1%
1-
12
#789940000000
0!
0%
b1 *
0-
02
b1 6
#789950000000
1!
1%
1-
12
#789960000000
0!
0%
b10 *
0-
02
b10 6
#789970000000
1!
1%
1-
12
#789980000000
0!
0%
b11 *
0-
02
b11 6
#789990000000
1!
1%
1-
12
15
#790000000000
0!
0%
b100 *
0-
02
b100 6
#790010000000
1!
1%
1-
12
#790020000000
0!
0%
b101 *
0-
02
b101 6
#790030000000
1!
1%
1-
12
#790040000000
0!
0%
b110 *
0-
02
b110 6
#790050000000
1!
1%
1-
12
#790060000000
0!
0%
b111 *
0-
02
b111 6
#790070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#790080000000
0!
0%
b0 *
0-
02
b0 6
#790090000000
1!
1%
1-
12
#790100000000
0!
0%
b1 *
0-
02
b1 6
#790110000000
1!
1%
1-
12
#790120000000
0!
0%
b10 *
0-
02
b10 6
#790130000000
1!
1%
1-
12
#790140000000
0!
0%
b11 *
0-
02
b11 6
#790150000000
1!
1%
1-
12
15
#790160000000
0!
0%
b100 *
0-
02
b100 6
#790170000000
1!
1%
1-
12
#790180000000
0!
0%
b101 *
0-
02
b101 6
#790190000000
1!
1%
1-
12
#790200000000
0!
0%
b110 *
0-
02
b110 6
#790210000000
1!
1%
1-
12
#790220000000
0!
0%
b111 *
0-
02
b111 6
#790230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#790240000000
0!
0%
b0 *
0-
02
b0 6
#790250000000
1!
1%
1-
12
#790260000000
0!
0%
b1 *
0-
02
b1 6
#790270000000
1!
1%
1-
12
#790280000000
0!
0%
b10 *
0-
02
b10 6
#790290000000
1!
1%
1-
12
#790300000000
0!
0%
b11 *
0-
02
b11 6
#790310000000
1!
1%
1-
12
15
#790320000000
0!
0%
b100 *
0-
02
b100 6
#790330000000
1!
1%
1-
12
#790340000000
0!
0%
b101 *
0-
02
b101 6
#790350000000
1!
1%
1-
12
#790360000000
0!
0%
b110 *
0-
02
b110 6
#790370000000
1!
1%
1-
12
#790380000000
0!
0%
b111 *
0-
02
b111 6
#790390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#790400000000
0!
0%
b0 *
0-
02
b0 6
#790410000000
1!
1%
1-
12
#790420000000
0!
0%
b1 *
0-
02
b1 6
#790430000000
1!
1%
1-
12
#790440000000
0!
0%
b10 *
0-
02
b10 6
#790450000000
1!
1%
1-
12
#790460000000
0!
0%
b11 *
0-
02
b11 6
#790470000000
1!
1%
1-
12
15
#790480000000
0!
0%
b100 *
0-
02
b100 6
#790490000000
1!
1%
1-
12
#790500000000
0!
0%
b101 *
0-
02
b101 6
#790510000000
1!
1%
1-
12
#790520000000
0!
0%
b110 *
0-
02
b110 6
#790530000000
1!
1%
1-
12
#790540000000
0!
0%
b111 *
0-
02
b111 6
#790550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#790560000000
0!
0%
b0 *
0-
02
b0 6
#790570000000
1!
1%
1-
12
#790580000000
0!
0%
b1 *
0-
02
b1 6
#790590000000
1!
1%
1-
12
#790600000000
0!
0%
b10 *
0-
02
b10 6
#790610000000
1!
1%
1-
12
#790620000000
0!
0%
b11 *
0-
02
b11 6
#790630000000
1!
1%
1-
12
15
#790640000000
0!
0%
b100 *
0-
02
b100 6
#790650000000
1!
1%
1-
12
#790660000000
0!
0%
b101 *
0-
02
b101 6
#790670000000
1!
1%
1-
12
#790680000000
0!
0%
b110 *
0-
02
b110 6
#790690000000
1!
1%
1-
12
#790700000000
0!
0%
b111 *
0-
02
b111 6
#790710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#790720000000
0!
0%
b0 *
0-
02
b0 6
#790730000000
1!
1%
1-
12
#790740000000
0!
0%
b1 *
0-
02
b1 6
#790750000000
1!
1%
1-
12
#790760000000
0!
0%
b10 *
0-
02
b10 6
#790770000000
1!
1%
1-
12
#790780000000
0!
0%
b11 *
0-
02
b11 6
#790790000000
1!
1%
1-
12
15
#790800000000
0!
0%
b100 *
0-
02
b100 6
#790810000000
1!
1%
1-
12
#790820000000
0!
0%
b101 *
0-
02
b101 6
#790830000000
1!
1%
1-
12
#790840000000
0!
0%
b110 *
0-
02
b110 6
#790850000000
1!
1%
1-
12
#790860000000
0!
0%
b111 *
0-
02
b111 6
#790870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#790880000000
0!
0%
b0 *
0-
02
b0 6
#790890000000
1!
1%
1-
12
#790900000000
0!
0%
b1 *
0-
02
b1 6
#790910000000
1!
1%
1-
12
#790920000000
0!
0%
b10 *
0-
02
b10 6
#790930000000
1!
1%
1-
12
#790940000000
0!
0%
b11 *
0-
02
b11 6
#790950000000
1!
1%
1-
12
15
#790960000000
0!
0%
b100 *
0-
02
b100 6
#790970000000
1!
1%
1-
12
#790980000000
0!
0%
b101 *
0-
02
b101 6
#790990000000
1!
1%
1-
12
#791000000000
0!
0%
b110 *
0-
02
b110 6
#791010000000
1!
1%
1-
12
#791020000000
0!
0%
b111 *
0-
02
b111 6
#791030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#791040000000
0!
0%
b0 *
0-
02
b0 6
#791050000000
1!
1%
1-
12
#791060000000
0!
0%
b1 *
0-
02
b1 6
#791070000000
1!
1%
1-
12
#791080000000
0!
0%
b10 *
0-
02
b10 6
#791090000000
1!
1%
1-
12
#791100000000
0!
0%
b11 *
0-
02
b11 6
#791110000000
1!
1%
1-
12
15
#791120000000
0!
0%
b100 *
0-
02
b100 6
#791130000000
1!
1%
1-
12
#791140000000
0!
0%
b101 *
0-
02
b101 6
#791150000000
1!
1%
1-
12
#791160000000
0!
0%
b110 *
0-
02
b110 6
#791170000000
1!
1%
1-
12
#791180000000
0!
0%
b111 *
0-
02
b111 6
#791190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#791200000000
0!
0%
b0 *
0-
02
b0 6
#791210000000
1!
1%
1-
12
#791220000000
0!
0%
b1 *
0-
02
b1 6
#791230000000
1!
1%
1-
12
#791240000000
0!
0%
b10 *
0-
02
b10 6
#791250000000
1!
1%
1-
12
#791260000000
0!
0%
b11 *
0-
02
b11 6
#791270000000
1!
1%
1-
12
15
#791280000000
0!
0%
b100 *
0-
02
b100 6
#791290000000
1!
1%
1-
12
#791300000000
0!
0%
b101 *
0-
02
b101 6
#791310000000
1!
1%
1-
12
#791320000000
0!
0%
b110 *
0-
02
b110 6
#791330000000
1!
1%
1-
12
#791340000000
0!
0%
b111 *
0-
02
b111 6
#791350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#791360000000
0!
0%
b0 *
0-
02
b0 6
#791370000000
1!
1%
1-
12
#791380000000
0!
0%
b1 *
0-
02
b1 6
#791390000000
1!
1%
1-
12
#791400000000
0!
0%
b10 *
0-
02
b10 6
#791410000000
1!
1%
1-
12
#791420000000
0!
0%
b11 *
0-
02
b11 6
#791430000000
1!
1%
1-
12
15
#791440000000
0!
0%
b100 *
0-
02
b100 6
#791450000000
1!
1%
1-
12
#791460000000
0!
0%
b101 *
0-
02
b101 6
#791470000000
1!
1%
1-
12
#791480000000
0!
0%
b110 *
0-
02
b110 6
#791490000000
1!
1%
1-
12
#791500000000
0!
0%
b111 *
0-
02
b111 6
#791510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#791520000000
0!
0%
b0 *
0-
02
b0 6
#791530000000
1!
1%
1-
12
#791540000000
0!
0%
b1 *
0-
02
b1 6
#791550000000
1!
1%
1-
12
#791560000000
0!
0%
b10 *
0-
02
b10 6
#791570000000
1!
1%
1-
12
#791580000000
0!
0%
b11 *
0-
02
b11 6
#791590000000
1!
1%
1-
12
15
#791600000000
0!
0%
b100 *
0-
02
b100 6
#791610000000
1!
1%
1-
12
#791620000000
0!
0%
b101 *
0-
02
b101 6
#791630000000
1!
1%
1-
12
#791640000000
0!
0%
b110 *
0-
02
b110 6
#791650000000
1!
1%
1-
12
#791660000000
0!
0%
b111 *
0-
02
b111 6
#791670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#791680000000
0!
0%
b0 *
0-
02
b0 6
#791690000000
1!
1%
1-
12
#791700000000
0!
0%
b1 *
0-
02
b1 6
#791710000000
1!
1%
1-
12
#791720000000
0!
0%
b10 *
0-
02
b10 6
#791730000000
1!
1%
1-
12
#791740000000
0!
0%
b11 *
0-
02
b11 6
#791750000000
1!
1%
1-
12
15
#791760000000
0!
0%
b100 *
0-
02
b100 6
#791770000000
1!
1%
1-
12
#791780000000
0!
0%
b101 *
0-
02
b101 6
#791790000000
1!
1%
1-
12
#791800000000
0!
0%
b110 *
0-
02
b110 6
#791810000000
1!
1%
1-
12
#791820000000
0!
0%
b111 *
0-
02
b111 6
#791830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#791840000000
0!
0%
b0 *
0-
02
b0 6
#791850000000
1!
1%
1-
12
#791860000000
0!
0%
b1 *
0-
02
b1 6
#791870000000
1!
1%
1-
12
#791880000000
0!
0%
b10 *
0-
02
b10 6
#791890000000
1!
1%
1-
12
#791900000000
0!
0%
b11 *
0-
02
b11 6
#791910000000
1!
1%
1-
12
15
#791920000000
0!
0%
b100 *
0-
02
b100 6
#791930000000
1!
1%
1-
12
#791940000000
0!
0%
b101 *
0-
02
b101 6
#791950000000
1!
1%
1-
12
#791960000000
0!
0%
b110 *
0-
02
b110 6
#791970000000
1!
1%
1-
12
#791980000000
0!
0%
b111 *
0-
02
b111 6
#791990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#792000000000
0!
0%
b0 *
0-
02
b0 6
#792010000000
1!
1%
1-
12
#792020000000
0!
0%
b1 *
0-
02
b1 6
#792030000000
1!
1%
1-
12
#792040000000
0!
0%
b10 *
0-
02
b10 6
#792050000000
1!
1%
1-
12
#792060000000
0!
0%
b11 *
0-
02
b11 6
#792070000000
1!
1%
1-
12
15
#792080000000
0!
0%
b100 *
0-
02
b100 6
#792090000000
1!
1%
1-
12
#792100000000
0!
0%
b101 *
0-
02
b101 6
#792110000000
1!
1%
1-
12
#792120000000
0!
0%
b110 *
0-
02
b110 6
#792130000000
1!
1%
1-
12
#792140000000
0!
0%
b111 *
0-
02
b111 6
#792150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#792160000000
0!
0%
b0 *
0-
02
b0 6
#792170000000
1!
1%
1-
12
#792180000000
0!
0%
b1 *
0-
02
b1 6
#792190000000
1!
1%
1-
12
#792200000000
0!
0%
b10 *
0-
02
b10 6
#792210000000
1!
1%
1-
12
#792220000000
0!
0%
b11 *
0-
02
b11 6
#792230000000
1!
1%
1-
12
15
#792240000000
0!
0%
b100 *
0-
02
b100 6
#792250000000
1!
1%
1-
12
#792260000000
0!
0%
b101 *
0-
02
b101 6
#792270000000
1!
1%
1-
12
#792280000000
0!
0%
b110 *
0-
02
b110 6
#792290000000
1!
1%
1-
12
#792300000000
0!
0%
b111 *
0-
02
b111 6
#792310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#792320000000
0!
0%
b0 *
0-
02
b0 6
#792330000000
1!
1%
1-
12
#792340000000
0!
0%
b1 *
0-
02
b1 6
#792350000000
1!
1%
1-
12
#792360000000
0!
0%
b10 *
0-
02
b10 6
#792370000000
1!
1%
1-
12
#792380000000
0!
0%
b11 *
0-
02
b11 6
#792390000000
1!
1%
1-
12
15
#792400000000
0!
0%
b100 *
0-
02
b100 6
#792410000000
1!
1%
1-
12
#792420000000
0!
0%
b101 *
0-
02
b101 6
#792430000000
1!
1%
1-
12
#792440000000
0!
0%
b110 *
0-
02
b110 6
#792450000000
1!
1%
1-
12
#792460000000
0!
0%
b111 *
0-
02
b111 6
#792470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#792480000000
0!
0%
b0 *
0-
02
b0 6
#792490000000
1!
1%
1-
12
#792500000000
0!
0%
b1 *
0-
02
b1 6
#792510000000
1!
1%
1-
12
#792520000000
0!
0%
b10 *
0-
02
b10 6
#792530000000
1!
1%
1-
12
#792540000000
0!
0%
b11 *
0-
02
b11 6
#792550000000
1!
1%
1-
12
15
#792560000000
0!
0%
b100 *
0-
02
b100 6
#792570000000
1!
1%
1-
12
#792580000000
0!
0%
b101 *
0-
02
b101 6
#792590000000
1!
1%
1-
12
#792600000000
0!
0%
b110 *
0-
02
b110 6
#792610000000
1!
1%
1-
12
#792620000000
0!
0%
b111 *
0-
02
b111 6
#792630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#792640000000
0!
0%
b0 *
0-
02
b0 6
#792650000000
1!
1%
1-
12
#792660000000
0!
0%
b1 *
0-
02
b1 6
#792670000000
1!
1%
1-
12
#792680000000
0!
0%
b10 *
0-
02
b10 6
#792690000000
1!
1%
1-
12
#792700000000
0!
0%
b11 *
0-
02
b11 6
#792710000000
1!
1%
1-
12
15
#792720000000
0!
0%
b100 *
0-
02
b100 6
#792730000000
1!
1%
1-
12
#792740000000
0!
0%
b101 *
0-
02
b101 6
#792750000000
1!
1%
1-
12
#792760000000
0!
0%
b110 *
0-
02
b110 6
#792770000000
1!
1%
1-
12
#792780000000
0!
0%
b111 *
0-
02
b111 6
#792790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#792800000000
0!
0%
b0 *
0-
02
b0 6
#792810000000
1!
1%
1-
12
#792820000000
0!
0%
b1 *
0-
02
b1 6
#792830000000
1!
1%
1-
12
#792840000000
0!
0%
b10 *
0-
02
b10 6
#792850000000
1!
1%
1-
12
#792860000000
0!
0%
b11 *
0-
02
b11 6
#792870000000
1!
1%
1-
12
15
#792880000000
0!
0%
b100 *
0-
02
b100 6
#792890000000
1!
1%
1-
12
#792900000000
0!
0%
b101 *
0-
02
b101 6
#792910000000
1!
1%
1-
12
#792920000000
0!
0%
b110 *
0-
02
b110 6
#792930000000
1!
1%
1-
12
#792940000000
0!
0%
b111 *
0-
02
b111 6
#792950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#792960000000
0!
0%
b0 *
0-
02
b0 6
#792970000000
1!
1%
1-
12
#792980000000
0!
0%
b1 *
0-
02
b1 6
#792990000000
1!
1%
1-
12
#793000000000
0!
0%
b10 *
0-
02
b10 6
#793010000000
1!
1%
1-
12
#793020000000
0!
0%
b11 *
0-
02
b11 6
#793030000000
1!
1%
1-
12
15
#793040000000
0!
0%
b100 *
0-
02
b100 6
#793050000000
1!
1%
1-
12
#793060000000
0!
0%
b101 *
0-
02
b101 6
#793070000000
1!
1%
1-
12
#793080000000
0!
0%
b110 *
0-
02
b110 6
#793090000000
1!
1%
1-
12
#793100000000
0!
0%
b111 *
0-
02
b111 6
#793110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#793120000000
0!
0%
b0 *
0-
02
b0 6
#793130000000
1!
1%
1-
12
#793140000000
0!
0%
b1 *
0-
02
b1 6
#793150000000
1!
1%
1-
12
#793160000000
0!
0%
b10 *
0-
02
b10 6
#793170000000
1!
1%
1-
12
#793180000000
0!
0%
b11 *
0-
02
b11 6
#793190000000
1!
1%
1-
12
15
#793200000000
0!
0%
b100 *
0-
02
b100 6
#793210000000
1!
1%
1-
12
#793220000000
0!
0%
b101 *
0-
02
b101 6
#793230000000
1!
1%
1-
12
#793240000000
0!
0%
b110 *
0-
02
b110 6
#793250000000
1!
1%
1-
12
#793260000000
0!
0%
b111 *
0-
02
b111 6
#793270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#793280000000
0!
0%
b0 *
0-
02
b0 6
#793290000000
1!
1%
1-
12
#793300000000
0!
0%
b1 *
0-
02
b1 6
#793310000000
1!
1%
1-
12
#793320000000
0!
0%
b10 *
0-
02
b10 6
#793330000000
1!
1%
1-
12
#793340000000
0!
0%
b11 *
0-
02
b11 6
#793350000000
1!
1%
1-
12
15
#793360000000
0!
0%
b100 *
0-
02
b100 6
#793370000000
1!
1%
1-
12
#793380000000
0!
0%
b101 *
0-
02
b101 6
#793390000000
1!
1%
1-
12
#793400000000
0!
0%
b110 *
0-
02
b110 6
#793410000000
1!
1%
1-
12
#793420000000
0!
0%
b111 *
0-
02
b111 6
#793430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#793440000000
0!
0%
b0 *
0-
02
b0 6
#793450000000
1!
1%
1-
12
#793460000000
0!
0%
b1 *
0-
02
b1 6
#793470000000
1!
1%
1-
12
#793480000000
0!
0%
b10 *
0-
02
b10 6
#793490000000
1!
1%
1-
12
#793500000000
0!
0%
b11 *
0-
02
b11 6
#793510000000
1!
1%
1-
12
15
#793520000000
0!
0%
b100 *
0-
02
b100 6
#793530000000
1!
1%
1-
12
#793540000000
0!
0%
b101 *
0-
02
b101 6
#793550000000
1!
1%
1-
12
#793560000000
0!
0%
b110 *
0-
02
b110 6
#793570000000
1!
1%
1-
12
#793580000000
0!
0%
b111 *
0-
02
b111 6
#793590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#793600000000
0!
0%
b0 *
0-
02
b0 6
#793610000000
1!
1%
1-
12
#793620000000
0!
0%
b1 *
0-
02
b1 6
#793630000000
1!
1%
1-
12
#793640000000
0!
0%
b10 *
0-
02
b10 6
#793650000000
1!
1%
1-
12
#793660000000
0!
0%
b11 *
0-
02
b11 6
#793670000000
1!
1%
1-
12
15
#793680000000
0!
0%
b100 *
0-
02
b100 6
#793690000000
1!
1%
1-
12
#793700000000
0!
0%
b101 *
0-
02
b101 6
#793710000000
1!
1%
1-
12
#793720000000
0!
0%
b110 *
0-
02
b110 6
#793730000000
1!
1%
1-
12
#793740000000
0!
0%
b111 *
0-
02
b111 6
#793750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#793760000000
0!
0%
b0 *
0-
02
b0 6
#793770000000
1!
1%
1-
12
#793780000000
0!
0%
b1 *
0-
02
b1 6
#793790000000
1!
1%
1-
12
#793800000000
0!
0%
b10 *
0-
02
b10 6
#793810000000
1!
1%
1-
12
#793820000000
0!
0%
b11 *
0-
02
b11 6
#793830000000
1!
1%
1-
12
15
#793840000000
0!
0%
b100 *
0-
02
b100 6
#793850000000
1!
1%
1-
12
#793860000000
0!
0%
b101 *
0-
02
b101 6
#793870000000
1!
1%
1-
12
#793880000000
0!
0%
b110 *
0-
02
b110 6
#793890000000
1!
1%
1-
12
#793900000000
0!
0%
b111 *
0-
02
b111 6
#793910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#793920000000
0!
0%
b0 *
0-
02
b0 6
#793930000000
1!
1%
1-
12
#793940000000
0!
0%
b1 *
0-
02
b1 6
#793950000000
1!
1%
1-
12
#793960000000
0!
0%
b10 *
0-
02
b10 6
#793970000000
1!
1%
1-
12
#793980000000
0!
0%
b11 *
0-
02
b11 6
#793990000000
1!
1%
1-
12
15
#794000000000
0!
0%
b100 *
0-
02
b100 6
#794010000000
1!
1%
1-
12
#794020000000
0!
0%
b101 *
0-
02
b101 6
#794030000000
1!
1%
1-
12
#794040000000
0!
0%
b110 *
0-
02
b110 6
#794050000000
1!
1%
1-
12
#794060000000
0!
0%
b111 *
0-
02
b111 6
#794070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#794080000000
0!
0%
b0 *
0-
02
b0 6
#794090000000
1!
1%
1-
12
#794100000000
0!
0%
b1 *
0-
02
b1 6
#794110000000
1!
1%
1-
12
#794120000000
0!
0%
b10 *
0-
02
b10 6
#794130000000
1!
1%
1-
12
#794140000000
0!
0%
b11 *
0-
02
b11 6
#794150000000
1!
1%
1-
12
15
#794160000000
0!
0%
b100 *
0-
02
b100 6
#794170000000
1!
1%
1-
12
#794180000000
0!
0%
b101 *
0-
02
b101 6
#794190000000
1!
1%
1-
12
#794200000000
0!
0%
b110 *
0-
02
b110 6
#794210000000
1!
1%
1-
12
#794220000000
0!
0%
b111 *
0-
02
b111 6
#794230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#794240000000
0!
0%
b0 *
0-
02
b0 6
#794250000000
1!
1%
1-
12
#794260000000
0!
0%
b1 *
0-
02
b1 6
#794270000000
1!
1%
1-
12
#794280000000
0!
0%
b10 *
0-
02
b10 6
#794290000000
1!
1%
1-
12
#794300000000
0!
0%
b11 *
0-
02
b11 6
#794310000000
1!
1%
1-
12
15
#794320000000
0!
0%
b100 *
0-
02
b100 6
#794330000000
1!
1%
1-
12
#794340000000
0!
0%
b101 *
0-
02
b101 6
#794350000000
1!
1%
1-
12
#794360000000
0!
0%
b110 *
0-
02
b110 6
#794370000000
1!
1%
1-
12
#794380000000
0!
0%
b111 *
0-
02
b111 6
#794390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#794400000000
0!
0%
b0 *
0-
02
b0 6
#794410000000
1!
1%
1-
12
#794420000000
0!
0%
b1 *
0-
02
b1 6
#794430000000
1!
1%
1-
12
#794440000000
0!
0%
b10 *
0-
02
b10 6
#794450000000
1!
1%
1-
12
#794460000000
0!
0%
b11 *
0-
02
b11 6
#794470000000
1!
1%
1-
12
15
#794480000000
0!
0%
b100 *
0-
02
b100 6
#794490000000
1!
1%
1-
12
#794500000000
0!
0%
b101 *
0-
02
b101 6
#794510000000
1!
1%
1-
12
#794520000000
0!
0%
b110 *
0-
02
b110 6
#794530000000
1!
1%
1-
12
#794540000000
0!
0%
b111 *
0-
02
b111 6
#794550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#794560000000
0!
0%
b0 *
0-
02
b0 6
#794570000000
1!
1%
1-
12
#794580000000
0!
0%
b1 *
0-
02
b1 6
#794590000000
1!
1%
1-
12
#794600000000
0!
0%
b10 *
0-
02
b10 6
#794610000000
1!
1%
1-
12
#794620000000
0!
0%
b11 *
0-
02
b11 6
#794630000000
1!
1%
1-
12
15
#794640000000
0!
0%
b100 *
0-
02
b100 6
#794650000000
1!
1%
1-
12
#794660000000
0!
0%
b101 *
0-
02
b101 6
#794670000000
1!
1%
1-
12
#794680000000
0!
0%
b110 *
0-
02
b110 6
#794690000000
1!
1%
1-
12
#794700000000
0!
0%
b111 *
0-
02
b111 6
#794710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#794720000000
0!
0%
b0 *
0-
02
b0 6
#794730000000
1!
1%
1-
12
#794740000000
0!
0%
b1 *
0-
02
b1 6
#794750000000
1!
1%
1-
12
#794760000000
0!
0%
b10 *
0-
02
b10 6
#794770000000
1!
1%
1-
12
#794780000000
0!
0%
b11 *
0-
02
b11 6
#794790000000
1!
1%
1-
12
15
#794800000000
0!
0%
b100 *
0-
02
b100 6
#794810000000
1!
1%
1-
12
#794820000000
0!
0%
b101 *
0-
02
b101 6
#794830000000
1!
1%
1-
12
#794840000000
0!
0%
b110 *
0-
02
b110 6
#794850000000
1!
1%
1-
12
#794860000000
0!
0%
b111 *
0-
02
b111 6
#794870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#794880000000
0!
0%
b0 *
0-
02
b0 6
#794890000000
1!
1%
1-
12
#794900000000
0!
0%
b1 *
0-
02
b1 6
#794910000000
1!
1%
1-
12
#794920000000
0!
0%
b10 *
0-
02
b10 6
#794930000000
1!
1%
1-
12
#794940000000
0!
0%
b11 *
0-
02
b11 6
#794950000000
1!
1%
1-
12
15
#794960000000
0!
0%
b100 *
0-
02
b100 6
#794970000000
1!
1%
1-
12
#794980000000
0!
0%
b101 *
0-
02
b101 6
#794990000000
1!
1%
1-
12
#795000000000
0!
0%
b110 *
0-
02
b110 6
#795010000000
1!
1%
1-
12
#795020000000
0!
0%
b111 *
0-
02
b111 6
#795030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#795040000000
0!
0%
b0 *
0-
02
b0 6
#795050000000
1!
1%
1-
12
#795060000000
0!
0%
b1 *
0-
02
b1 6
#795070000000
1!
1%
1-
12
#795080000000
0!
0%
b10 *
0-
02
b10 6
#795090000000
1!
1%
1-
12
#795100000000
0!
0%
b11 *
0-
02
b11 6
#795110000000
1!
1%
1-
12
15
#795120000000
0!
0%
b100 *
0-
02
b100 6
#795130000000
1!
1%
1-
12
#795140000000
0!
0%
b101 *
0-
02
b101 6
#795150000000
1!
1%
1-
12
#795160000000
0!
0%
b110 *
0-
02
b110 6
#795170000000
1!
1%
1-
12
#795180000000
0!
0%
b111 *
0-
02
b111 6
#795190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#795200000000
0!
0%
b0 *
0-
02
b0 6
#795210000000
1!
1%
1-
12
#795220000000
0!
0%
b1 *
0-
02
b1 6
#795230000000
1!
1%
1-
12
#795240000000
0!
0%
b10 *
0-
02
b10 6
#795250000000
1!
1%
1-
12
#795260000000
0!
0%
b11 *
0-
02
b11 6
#795270000000
1!
1%
1-
12
15
#795280000000
0!
0%
b100 *
0-
02
b100 6
#795290000000
1!
1%
1-
12
#795300000000
0!
0%
b101 *
0-
02
b101 6
#795310000000
1!
1%
1-
12
#795320000000
0!
0%
b110 *
0-
02
b110 6
#795330000000
1!
1%
1-
12
#795340000000
0!
0%
b111 *
0-
02
b111 6
#795350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#795360000000
0!
0%
b0 *
0-
02
b0 6
#795370000000
1!
1%
1-
12
#795380000000
0!
0%
b1 *
0-
02
b1 6
#795390000000
1!
1%
1-
12
#795400000000
0!
0%
b10 *
0-
02
b10 6
#795410000000
1!
1%
1-
12
#795420000000
0!
0%
b11 *
0-
02
b11 6
#795430000000
1!
1%
1-
12
15
#795440000000
0!
0%
b100 *
0-
02
b100 6
#795450000000
1!
1%
1-
12
#795460000000
0!
0%
b101 *
0-
02
b101 6
#795470000000
1!
1%
1-
12
#795480000000
0!
0%
b110 *
0-
02
b110 6
#795490000000
1!
1%
1-
12
#795500000000
0!
0%
b111 *
0-
02
b111 6
#795510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#795520000000
0!
0%
b0 *
0-
02
b0 6
#795530000000
1!
1%
1-
12
#795540000000
0!
0%
b1 *
0-
02
b1 6
#795550000000
1!
1%
1-
12
#795560000000
0!
0%
b10 *
0-
02
b10 6
#795570000000
1!
1%
1-
12
#795580000000
0!
0%
b11 *
0-
02
b11 6
#795590000000
1!
1%
1-
12
15
#795600000000
0!
0%
b100 *
0-
02
b100 6
#795610000000
1!
1%
1-
12
#795620000000
0!
0%
b101 *
0-
02
b101 6
#795630000000
1!
1%
1-
12
#795640000000
0!
0%
b110 *
0-
02
b110 6
#795650000000
1!
1%
1-
12
#795660000000
0!
0%
b111 *
0-
02
b111 6
#795670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#795680000000
0!
0%
b0 *
0-
02
b0 6
#795690000000
1!
1%
1-
12
#795700000000
0!
0%
b1 *
0-
02
b1 6
#795710000000
1!
1%
1-
12
#795720000000
0!
0%
b10 *
0-
02
b10 6
#795730000000
1!
1%
1-
12
#795740000000
0!
0%
b11 *
0-
02
b11 6
#795750000000
1!
1%
1-
12
15
#795760000000
0!
0%
b100 *
0-
02
b100 6
#795770000000
1!
1%
1-
12
#795780000000
0!
0%
b101 *
0-
02
b101 6
#795790000000
1!
1%
1-
12
#795800000000
0!
0%
b110 *
0-
02
b110 6
#795810000000
1!
1%
1-
12
#795820000000
0!
0%
b111 *
0-
02
b111 6
#795830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#795840000000
0!
0%
b0 *
0-
02
b0 6
#795850000000
1!
1%
1-
12
#795860000000
0!
0%
b1 *
0-
02
b1 6
#795870000000
1!
1%
1-
12
#795880000000
0!
0%
b10 *
0-
02
b10 6
#795890000000
1!
1%
1-
12
#795900000000
0!
0%
b11 *
0-
02
b11 6
#795910000000
1!
1%
1-
12
15
#795920000000
0!
0%
b100 *
0-
02
b100 6
#795930000000
1!
1%
1-
12
#795940000000
0!
0%
b101 *
0-
02
b101 6
#795950000000
1!
1%
1-
12
#795960000000
0!
0%
b110 *
0-
02
b110 6
#795970000000
1!
1%
1-
12
#795980000000
0!
0%
b111 *
0-
02
b111 6
#795990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#796000000000
0!
0%
b0 *
0-
02
b0 6
#796010000000
1!
1%
1-
12
#796020000000
0!
0%
b1 *
0-
02
b1 6
#796030000000
1!
1%
1-
12
#796040000000
0!
0%
b10 *
0-
02
b10 6
#796050000000
1!
1%
1-
12
#796060000000
0!
0%
b11 *
0-
02
b11 6
#796070000000
1!
1%
1-
12
15
#796080000000
0!
0%
b100 *
0-
02
b100 6
#796090000000
1!
1%
1-
12
#796100000000
0!
0%
b101 *
0-
02
b101 6
#796110000000
1!
1%
1-
12
#796120000000
0!
0%
b110 *
0-
02
b110 6
#796130000000
1!
1%
1-
12
#796140000000
0!
0%
b111 *
0-
02
b111 6
#796150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#796160000000
0!
0%
b0 *
0-
02
b0 6
#796170000000
1!
1%
1-
12
#796180000000
0!
0%
b1 *
0-
02
b1 6
#796190000000
1!
1%
1-
12
#796200000000
0!
0%
b10 *
0-
02
b10 6
#796210000000
1!
1%
1-
12
#796220000000
0!
0%
b11 *
0-
02
b11 6
#796230000000
1!
1%
1-
12
15
#796240000000
0!
0%
b100 *
0-
02
b100 6
#796250000000
1!
1%
1-
12
#796260000000
0!
0%
b101 *
0-
02
b101 6
#796270000000
1!
1%
1-
12
#796280000000
0!
0%
b110 *
0-
02
b110 6
#796290000000
1!
1%
1-
12
#796300000000
0!
0%
b111 *
0-
02
b111 6
#796310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#796320000000
0!
0%
b0 *
0-
02
b0 6
#796330000000
1!
1%
1-
12
#796340000000
0!
0%
b1 *
0-
02
b1 6
#796350000000
1!
1%
1-
12
#796360000000
0!
0%
b10 *
0-
02
b10 6
#796370000000
1!
1%
1-
12
#796380000000
0!
0%
b11 *
0-
02
b11 6
#796390000000
1!
1%
1-
12
15
#796400000000
0!
0%
b100 *
0-
02
b100 6
#796410000000
1!
1%
1-
12
#796420000000
0!
0%
b101 *
0-
02
b101 6
#796430000000
1!
1%
1-
12
#796440000000
0!
0%
b110 *
0-
02
b110 6
#796450000000
1!
1%
1-
12
#796460000000
0!
0%
b111 *
0-
02
b111 6
#796470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#796480000000
0!
0%
b0 *
0-
02
b0 6
#796490000000
1!
1%
1-
12
#796500000000
0!
0%
b1 *
0-
02
b1 6
#796510000000
1!
1%
1-
12
#796520000000
0!
0%
b10 *
0-
02
b10 6
#796530000000
1!
1%
1-
12
#796540000000
0!
0%
b11 *
0-
02
b11 6
#796550000000
1!
1%
1-
12
15
#796560000000
0!
0%
b100 *
0-
02
b100 6
#796570000000
1!
1%
1-
12
#796580000000
0!
0%
b101 *
0-
02
b101 6
#796590000000
1!
1%
1-
12
#796600000000
0!
0%
b110 *
0-
02
b110 6
#796610000000
1!
1%
1-
12
#796620000000
0!
0%
b111 *
0-
02
b111 6
#796630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#796640000000
0!
0%
b0 *
0-
02
b0 6
#796650000000
1!
1%
1-
12
#796660000000
0!
0%
b1 *
0-
02
b1 6
#796670000000
1!
1%
1-
12
#796680000000
0!
0%
b10 *
0-
02
b10 6
#796690000000
1!
1%
1-
12
#796700000000
0!
0%
b11 *
0-
02
b11 6
#796710000000
1!
1%
1-
12
15
#796720000000
0!
0%
b100 *
0-
02
b100 6
#796730000000
1!
1%
1-
12
#796740000000
0!
0%
b101 *
0-
02
b101 6
#796750000000
1!
1%
1-
12
#796760000000
0!
0%
b110 *
0-
02
b110 6
#796770000000
1!
1%
1-
12
#796780000000
0!
0%
b111 *
0-
02
b111 6
#796790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#796800000000
0!
0%
b0 *
0-
02
b0 6
#796810000000
1!
1%
1-
12
#796820000000
0!
0%
b1 *
0-
02
b1 6
#796830000000
1!
1%
1-
12
#796840000000
0!
0%
b10 *
0-
02
b10 6
#796850000000
1!
1%
1-
12
#796860000000
0!
0%
b11 *
0-
02
b11 6
#796870000000
1!
1%
1-
12
15
#796880000000
0!
0%
b100 *
0-
02
b100 6
#796890000000
1!
1%
1-
12
#796900000000
0!
0%
b101 *
0-
02
b101 6
#796910000000
1!
1%
1-
12
#796920000000
0!
0%
b110 *
0-
02
b110 6
#796930000000
1!
1%
1-
12
#796940000000
0!
0%
b111 *
0-
02
b111 6
#796950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#796960000000
0!
0%
b0 *
0-
02
b0 6
#796970000000
1!
1%
1-
12
#796980000000
0!
0%
b1 *
0-
02
b1 6
#796990000000
1!
1%
1-
12
#797000000000
0!
0%
b10 *
0-
02
b10 6
#797010000000
1!
1%
1-
12
#797020000000
0!
0%
b11 *
0-
02
b11 6
#797030000000
1!
1%
1-
12
15
#797040000000
0!
0%
b100 *
0-
02
b100 6
#797050000000
1!
1%
1-
12
#797060000000
0!
0%
b101 *
0-
02
b101 6
#797070000000
1!
1%
1-
12
#797080000000
0!
0%
b110 *
0-
02
b110 6
#797090000000
1!
1%
1-
12
#797100000000
0!
0%
b111 *
0-
02
b111 6
#797110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#797120000000
0!
0%
b0 *
0-
02
b0 6
#797130000000
1!
1%
1-
12
#797140000000
0!
0%
b1 *
0-
02
b1 6
#797150000000
1!
1%
1-
12
#797160000000
0!
0%
b10 *
0-
02
b10 6
#797170000000
1!
1%
1-
12
#797180000000
0!
0%
b11 *
0-
02
b11 6
#797190000000
1!
1%
1-
12
15
#797200000000
0!
0%
b100 *
0-
02
b100 6
#797210000000
1!
1%
1-
12
#797220000000
0!
0%
b101 *
0-
02
b101 6
#797230000000
1!
1%
1-
12
#797240000000
0!
0%
b110 *
0-
02
b110 6
#797250000000
1!
1%
1-
12
#797260000000
0!
0%
b111 *
0-
02
b111 6
#797270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#797280000000
0!
0%
b0 *
0-
02
b0 6
#797290000000
1!
1%
1-
12
#797300000000
0!
0%
b1 *
0-
02
b1 6
#797310000000
1!
1%
1-
12
#797320000000
0!
0%
b10 *
0-
02
b10 6
#797330000000
1!
1%
1-
12
#797340000000
0!
0%
b11 *
0-
02
b11 6
#797350000000
1!
1%
1-
12
15
#797360000000
0!
0%
b100 *
0-
02
b100 6
#797370000000
1!
1%
1-
12
#797380000000
0!
0%
b101 *
0-
02
b101 6
#797390000000
1!
1%
1-
12
#797400000000
0!
0%
b110 *
0-
02
b110 6
#797410000000
1!
1%
1-
12
#797420000000
0!
0%
b111 *
0-
02
b111 6
#797430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#797440000000
0!
0%
b0 *
0-
02
b0 6
#797450000000
1!
1%
1-
12
#797460000000
0!
0%
b1 *
0-
02
b1 6
#797470000000
1!
1%
1-
12
#797480000000
0!
0%
b10 *
0-
02
b10 6
#797490000000
1!
1%
1-
12
#797500000000
0!
0%
b11 *
0-
02
b11 6
#797510000000
1!
1%
1-
12
15
#797520000000
0!
0%
b100 *
0-
02
b100 6
#797530000000
1!
1%
1-
12
#797540000000
0!
0%
b101 *
0-
02
b101 6
#797550000000
1!
1%
1-
12
#797560000000
0!
0%
b110 *
0-
02
b110 6
#797570000000
1!
1%
1-
12
#797580000000
0!
0%
b111 *
0-
02
b111 6
#797590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#797600000000
0!
0%
b0 *
0-
02
b0 6
#797610000000
1!
1%
1-
12
#797620000000
0!
0%
b1 *
0-
02
b1 6
#797630000000
1!
1%
1-
12
#797640000000
0!
0%
b10 *
0-
02
b10 6
#797650000000
1!
1%
1-
12
#797660000000
0!
0%
b11 *
0-
02
b11 6
#797670000000
1!
1%
1-
12
15
#797680000000
0!
0%
b100 *
0-
02
b100 6
#797690000000
1!
1%
1-
12
#797700000000
0!
0%
b101 *
0-
02
b101 6
#797710000000
1!
1%
1-
12
#797720000000
0!
0%
b110 *
0-
02
b110 6
#797730000000
1!
1%
1-
12
#797740000000
0!
0%
b111 *
0-
02
b111 6
#797750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#797760000000
0!
0%
b0 *
0-
02
b0 6
#797770000000
1!
1%
1-
12
#797780000000
0!
0%
b1 *
0-
02
b1 6
#797790000000
1!
1%
1-
12
#797800000000
0!
0%
b10 *
0-
02
b10 6
#797810000000
1!
1%
1-
12
#797820000000
0!
0%
b11 *
0-
02
b11 6
#797830000000
1!
1%
1-
12
15
#797840000000
0!
0%
b100 *
0-
02
b100 6
#797850000000
1!
1%
1-
12
#797860000000
0!
0%
b101 *
0-
02
b101 6
#797870000000
1!
1%
1-
12
#797880000000
0!
0%
b110 *
0-
02
b110 6
#797890000000
1!
1%
1-
12
#797900000000
0!
0%
b111 *
0-
02
b111 6
#797910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#797920000000
0!
0%
b0 *
0-
02
b0 6
#797930000000
1!
1%
1-
12
#797940000000
0!
0%
b1 *
0-
02
b1 6
#797950000000
1!
1%
1-
12
#797960000000
0!
0%
b10 *
0-
02
b10 6
#797970000000
1!
1%
1-
12
#797980000000
0!
0%
b11 *
0-
02
b11 6
#797990000000
1!
1%
1-
12
15
#798000000000
0!
0%
b100 *
0-
02
b100 6
#798010000000
1!
1%
1-
12
#798020000000
0!
0%
b101 *
0-
02
b101 6
#798030000000
1!
1%
1-
12
#798040000000
0!
0%
b110 *
0-
02
b110 6
#798050000000
1!
1%
1-
12
#798060000000
0!
0%
b111 *
0-
02
b111 6
#798070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#798080000000
0!
0%
b0 *
0-
02
b0 6
#798090000000
1!
1%
1-
12
#798100000000
0!
0%
b1 *
0-
02
b1 6
#798110000000
1!
1%
1-
12
#798120000000
0!
0%
b10 *
0-
02
b10 6
#798130000000
1!
1%
1-
12
#798140000000
0!
0%
b11 *
0-
02
b11 6
#798150000000
1!
1%
1-
12
15
#798160000000
0!
0%
b100 *
0-
02
b100 6
#798170000000
1!
1%
1-
12
#798180000000
0!
0%
b101 *
0-
02
b101 6
#798190000000
1!
1%
1-
12
#798200000000
0!
0%
b110 *
0-
02
b110 6
#798210000000
1!
1%
1-
12
#798220000000
0!
0%
b111 *
0-
02
b111 6
#798230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#798240000000
0!
0%
b0 *
0-
02
b0 6
#798250000000
1!
1%
1-
12
#798260000000
0!
0%
b1 *
0-
02
b1 6
#798270000000
1!
1%
1-
12
#798280000000
0!
0%
b10 *
0-
02
b10 6
#798290000000
1!
1%
1-
12
#798300000000
0!
0%
b11 *
0-
02
b11 6
#798310000000
1!
1%
1-
12
15
#798320000000
0!
0%
b100 *
0-
02
b100 6
#798330000000
1!
1%
1-
12
#798340000000
0!
0%
b101 *
0-
02
b101 6
#798350000000
1!
1%
1-
12
#798360000000
0!
0%
b110 *
0-
02
b110 6
#798370000000
1!
1%
1-
12
#798380000000
0!
0%
b111 *
0-
02
b111 6
#798390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#798400000000
0!
0%
b0 *
0-
02
b0 6
#798410000000
1!
1%
1-
12
#798420000000
0!
0%
b1 *
0-
02
b1 6
#798430000000
1!
1%
1-
12
#798440000000
0!
0%
b10 *
0-
02
b10 6
#798450000000
1!
1%
1-
12
#798460000000
0!
0%
b11 *
0-
02
b11 6
#798470000000
1!
1%
1-
12
15
#798480000000
0!
0%
b100 *
0-
02
b100 6
#798490000000
1!
1%
1-
12
#798500000000
0!
0%
b101 *
0-
02
b101 6
#798510000000
1!
1%
1-
12
#798520000000
0!
0%
b110 *
0-
02
b110 6
#798530000000
1!
1%
1-
12
#798540000000
0!
0%
b111 *
0-
02
b111 6
#798550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#798560000000
0!
0%
b0 *
0-
02
b0 6
#798570000000
1!
1%
1-
12
#798580000000
0!
0%
b1 *
0-
02
b1 6
#798590000000
1!
1%
1-
12
#798600000000
0!
0%
b10 *
0-
02
b10 6
#798610000000
1!
1%
1-
12
#798620000000
0!
0%
b11 *
0-
02
b11 6
#798630000000
1!
1%
1-
12
15
#798640000000
0!
0%
b100 *
0-
02
b100 6
#798650000000
1!
1%
1-
12
#798660000000
0!
0%
b101 *
0-
02
b101 6
#798670000000
1!
1%
1-
12
#798680000000
0!
0%
b110 *
0-
02
b110 6
#798690000000
1!
1%
1-
12
#798700000000
0!
0%
b111 *
0-
02
b111 6
#798710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#798720000000
0!
0%
b0 *
0-
02
b0 6
#798730000000
1!
1%
1-
12
#798740000000
0!
0%
b1 *
0-
02
b1 6
#798750000000
1!
1%
1-
12
#798760000000
0!
0%
b10 *
0-
02
b10 6
#798770000000
1!
1%
1-
12
#798780000000
0!
0%
b11 *
0-
02
b11 6
#798790000000
1!
1%
1-
12
15
#798800000000
0!
0%
b100 *
0-
02
b100 6
#798810000000
1!
1%
1-
12
#798820000000
0!
0%
b101 *
0-
02
b101 6
#798830000000
1!
1%
1-
12
#798840000000
0!
0%
b110 *
0-
02
b110 6
#798850000000
1!
1%
1-
12
#798860000000
0!
0%
b111 *
0-
02
b111 6
#798870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#798880000000
0!
0%
b0 *
0-
02
b0 6
#798890000000
1!
1%
1-
12
#798900000000
0!
0%
b1 *
0-
02
b1 6
#798910000000
1!
1%
1-
12
#798920000000
0!
0%
b10 *
0-
02
b10 6
#798930000000
1!
1%
1-
12
#798940000000
0!
0%
b11 *
0-
02
b11 6
#798950000000
1!
1%
1-
12
15
#798960000000
0!
0%
b100 *
0-
02
b100 6
#798970000000
1!
1%
1-
12
#798980000000
0!
0%
b101 *
0-
02
b101 6
#798990000000
1!
1%
1-
12
#799000000000
0!
0%
b110 *
0-
02
b110 6
#799010000000
1!
1%
1-
12
#799020000000
0!
0%
b111 *
0-
02
b111 6
#799030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#799040000000
0!
0%
b0 *
0-
02
b0 6
#799050000000
1!
1%
1-
12
#799060000000
0!
0%
b1 *
0-
02
b1 6
#799070000000
1!
1%
1-
12
#799080000000
0!
0%
b10 *
0-
02
b10 6
#799090000000
1!
1%
1-
12
#799100000000
0!
0%
b11 *
0-
02
b11 6
#799110000000
1!
1%
1-
12
15
#799120000000
0!
0%
b100 *
0-
02
b100 6
#799130000000
1!
1%
1-
12
#799140000000
0!
0%
b101 *
0-
02
b101 6
#799150000000
1!
1%
1-
12
#799160000000
0!
0%
b110 *
0-
02
b110 6
#799170000000
1!
1%
1-
12
#799180000000
0!
0%
b111 *
0-
02
b111 6
#799190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#799200000000
0!
0%
b0 *
0-
02
b0 6
#799210000000
1!
1%
1-
12
#799220000000
0!
0%
b1 *
0-
02
b1 6
#799230000000
1!
1%
1-
12
#799240000000
0!
0%
b10 *
0-
02
b10 6
#799250000000
1!
1%
1-
12
#799260000000
0!
0%
b11 *
0-
02
b11 6
#799270000000
1!
1%
1-
12
15
#799280000000
0!
0%
b100 *
0-
02
b100 6
#799290000000
1!
1%
1-
12
#799300000000
0!
0%
b101 *
0-
02
b101 6
#799310000000
1!
1%
1-
12
#799320000000
0!
0%
b110 *
0-
02
b110 6
#799330000000
1!
1%
1-
12
#799340000000
0!
0%
b111 *
0-
02
b111 6
#799350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#799360000000
0!
0%
b0 *
0-
02
b0 6
#799370000000
1!
1%
1-
12
#799380000000
0!
0%
b1 *
0-
02
b1 6
#799390000000
1!
1%
1-
12
#799400000000
0!
0%
b10 *
0-
02
b10 6
#799410000000
1!
1%
1-
12
#799420000000
0!
0%
b11 *
0-
02
b11 6
#799430000000
1!
1%
1-
12
15
#799440000000
0!
0%
b100 *
0-
02
b100 6
#799450000000
1!
1%
1-
12
#799460000000
0!
0%
b101 *
0-
02
b101 6
#799470000000
1!
1%
1-
12
#799480000000
0!
0%
b110 *
0-
02
b110 6
#799490000000
1!
1%
1-
12
#799500000000
0!
0%
b111 *
0-
02
b111 6
#799510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#799520000000
0!
0%
b0 *
0-
02
b0 6
#799530000000
1!
1%
1-
12
#799540000000
0!
0%
b1 *
0-
02
b1 6
#799550000000
1!
1%
1-
12
#799560000000
0!
0%
b10 *
0-
02
b10 6
#799570000000
1!
1%
1-
12
#799580000000
0!
0%
b11 *
0-
02
b11 6
#799590000000
1!
1%
1-
12
15
#799600000000
0!
0%
b100 *
0-
02
b100 6
#799610000000
1!
1%
1-
12
#799620000000
0!
0%
b101 *
0-
02
b101 6
#799630000000
1!
1%
1-
12
#799640000000
0!
0%
b110 *
0-
02
b110 6
#799650000000
1!
1%
1-
12
#799660000000
0!
0%
b111 *
0-
02
b111 6
#799670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#799680000000
0!
0%
b0 *
0-
02
b0 6
#799690000000
1!
1%
1-
12
#799700000000
0!
0%
b1 *
0-
02
b1 6
#799710000000
1!
1%
1-
12
#799720000000
0!
0%
b10 *
0-
02
b10 6
#799730000000
1!
1%
1-
12
#799740000000
0!
0%
b11 *
0-
02
b11 6
#799750000000
1!
1%
1-
12
15
#799760000000
0!
0%
b100 *
0-
02
b100 6
#799770000000
1!
1%
1-
12
#799780000000
0!
0%
b101 *
0-
02
b101 6
#799790000000
1!
1%
1-
12
#799800000000
0!
0%
b110 *
0-
02
b110 6
#799810000000
1!
1%
1-
12
#799820000000
0!
0%
b111 *
0-
02
b111 6
#799830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#799840000000
0!
0%
b0 *
0-
02
b0 6
#799850000000
1!
1%
1-
12
#799860000000
0!
0%
b1 *
0-
02
b1 6
#799870000000
1!
1%
1-
12
#799880000000
0!
0%
b10 *
0-
02
b10 6
#799890000000
1!
1%
1-
12
#799900000000
0!
0%
b11 *
0-
02
b11 6
#799910000000
1!
1%
1-
12
15
#799920000000
0!
0%
b100 *
0-
02
b100 6
#799930000000
1!
1%
1-
12
#799940000000
0!
0%
b101 *
0-
02
b101 6
#799950000000
1!
1%
1-
12
#799960000000
0!
0%
b110 *
0-
02
b110 6
#799970000000
1!
1%
1-
12
#799980000000
0!
0%
b111 *
0-
02
b111 6
#799990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#800000000000
0!
0%
b0 *
0-
02
b0 6
#800010000000
1!
1%
1-
12
#800020000000
0!
0%
b1 *
0-
02
b1 6
#800030000000
1!
1%
1-
12
#800040000000
0!
0%
b10 *
0-
02
b10 6
#800050000000
1!
1%
1-
12
#800060000000
0!
0%
b11 *
0-
02
b11 6
#800070000000
1!
1%
1-
12
15
#800080000000
0!
0%
b100 *
0-
02
b100 6
#800090000000
1!
1%
1-
12
#800100000000
0!
0%
b101 *
0-
02
b101 6
#800110000000
1!
1%
1-
12
#800120000000
0!
0%
b110 *
0-
02
b110 6
#800130000000
1!
1%
1-
12
#800140000000
0!
0%
b111 *
0-
02
b111 6
#800150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#800160000000
0!
0%
b0 *
0-
02
b0 6
#800170000000
1!
1%
1-
12
#800180000000
0!
0%
b1 *
0-
02
b1 6
#800190000000
1!
1%
1-
12
#800200000000
0!
0%
b10 *
0-
02
b10 6
#800210000000
1!
1%
1-
12
#800220000000
0!
0%
b11 *
0-
02
b11 6
#800230000000
1!
1%
1-
12
15
#800240000000
0!
0%
b100 *
0-
02
b100 6
#800250000000
1!
1%
1-
12
#800260000000
0!
0%
b101 *
0-
02
b101 6
#800270000000
1!
1%
1-
12
#800280000000
0!
0%
b110 *
0-
02
b110 6
#800290000000
1!
1%
1-
12
#800300000000
0!
0%
b111 *
0-
02
b111 6
#800310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#800320000000
0!
0%
b0 *
0-
02
b0 6
#800330000000
1!
1%
1-
12
#800340000000
0!
0%
b1 *
0-
02
b1 6
#800350000000
1!
1%
1-
12
#800360000000
0!
0%
b10 *
0-
02
b10 6
#800370000000
1!
1%
1-
12
#800380000000
0!
0%
b11 *
0-
02
b11 6
#800390000000
1!
1%
1-
12
15
#800400000000
0!
0%
b100 *
0-
02
b100 6
#800410000000
1!
1%
1-
12
#800420000000
0!
0%
b101 *
0-
02
b101 6
#800430000000
1!
1%
1-
12
#800440000000
0!
0%
b110 *
0-
02
b110 6
#800450000000
1!
1%
1-
12
#800460000000
0!
0%
b111 *
0-
02
b111 6
#800470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#800480000000
0!
0%
b0 *
0-
02
b0 6
#800490000000
1!
1%
1-
12
#800500000000
0!
0%
b1 *
0-
02
b1 6
#800510000000
1!
1%
1-
12
#800520000000
0!
0%
b10 *
0-
02
b10 6
#800530000000
1!
1%
1-
12
#800540000000
0!
0%
b11 *
0-
02
b11 6
#800550000000
1!
1%
1-
12
15
#800560000000
0!
0%
b100 *
0-
02
b100 6
#800570000000
1!
1%
1-
12
#800580000000
0!
0%
b101 *
0-
02
b101 6
#800590000000
1!
1%
1-
12
#800600000000
0!
0%
b110 *
0-
02
b110 6
#800610000000
1!
1%
1-
12
#800620000000
0!
0%
b111 *
0-
02
b111 6
#800630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#800640000000
0!
0%
b0 *
0-
02
b0 6
#800650000000
1!
1%
1-
12
#800660000000
0!
0%
b1 *
0-
02
b1 6
#800670000000
1!
1%
1-
12
#800680000000
0!
0%
b10 *
0-
02
b10 6
#800690000000
1!
1%
1-
12
#800700000000
0!
0%
b11 *
0-
02
b11 6
#800710000000
1!
1%
1-
12
15
#800720000000
0!
0%
b100 *
0-
02
b100 6
#800730000000
1!
1%
1-
12
#800740000000
0!
0%
b101 *
0-
02
b101 6
#800750000000
1!
1%
1-
12
#800760000000
0!
0%
b110 *
0-
02
b110 6
#800770000000
1!
1%
1-
12
#800780000000
0!
0%
b111 *
0-
02
b111 6
#800790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#800800000000
0!
0%
b0 *
0-
02
b0 6
#800810000000
1!
1%
1-
12
#800820000000
0!
0%
b1 *
0-
02
b1 6
#800830000000
1!
1%
1-
12
#800840000000
0!
0%
b10 *
0-
02
b10 6
#800850000000
1!
1%
1-
12
#800860000000
0!
0%
b11 *
0-
02
b11 6
#800870000000
1!
1%
1-
12
15
#800880000000
0!
0%
b100 *
0-
02
b100 6
#800890000000
1!
1%
1-
12
#800900000000
0!
0%
b101 *
0-
02
b101 6
#800910000000
1!
1%
1-
12
#800920000000
0!
0%
b110 *
0-
02
b110 6
#800930000000
1!
1%
1-
12
#800940000000
0!
0%
b111 *
0-
02
b111 6
#800950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#800960000000
0!
0%
b0 *
0-
02
b0 6
#800970000000
1!
1%
1-
12
#800980000000
0!
0%
b1 *
0-
02
b1 6
#800990000000
1!
1%
1-
12
#801000000000
0!
0%
b10 *
0-
02
b10 6
#801010000000
1!
1%
1-
12
#801020000000
0!
0%
b11 *
0-
02
b11 6
#801030000000
1!
1%
1-
12
15
#801040000000
0!
0%
b100 *
0-
02
b100 6
#801050000000
1!
1%
1-
12
#801060000000
0!
0%
b101 *
0-
02
b101 6
#801070000000
1!
1%
1-
12
#801080000000
0!
0%
b110 *
0-
02
b110 6
#801090000000
1!
1%
1-
12
#801100000000
0!
0%
b111 *
0-
02
b111 6
#801110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#801120000000
0!
0%
b0 *
0-
02
b0 6
#801130000000
1!
1%
1-
12
#801140000000
0!
0%
b1 *
0-
02
b1 6
#801150000000
1!
1%
1-
12
#801160000000
0!
0%
b10 *
0-
02
b10 6
#801170000000
1!
1%
1-
12
#801180000000
0!
0%
b11 *
0-
02
b11 6
#801190000000
1!
1%
1-
12
15
#801200000000
0!
0%
b100 *
0-
02
b100 6
#801210000000
1!
1%
1-
12
#801220000000
0!
0%
b101 *
0-
02
b101 6
#801230000000
1!
1%
1-
12
#801240000000
0!
0%
b110 *
0-
02
b110 6
#801250000000
1!
1%
1-
12
#801260000000
0!
0%
b111 *
0-
02
b111 6
#801270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#801280000000
0!
0%
b0 *
0-
02
b0 6
#801290000000
1!
1%
1-
12
#801300000000
0!
0%
b1 *
0-
02
b1 6
#801310000000
1!
1%
1-
12
#801320000000
0!
0%
b10 *
0-
02
b10 6
#801330000000
1!
1%
1-
12
#801340000000
0!
0%
b11 *
0-
02
b11 6
#801350000000
1!
1%
1-
12
15
#801360000000
0!
0%
b100 *
0-
02
b100 6
#801370000000
1!
1%
1-
12
#801380000000
0!
0%
b101 *
0-
02
b101 6
#801390000000
1!
1%
1-
12
#801400000000
0!
0%
b110 *
0-
02
b110 6
#801410000000
1!
1%
1-
12
#801420000000
0!
0%
b111 *
0-
02
b111 6
#801430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#801440000000
0!
0%
b0 *
0-
02
b0 6
#801450000000
1!
1%
1-
12
#801460000000
0!
0%
b1 *
0-
02
b1 6
#801470000000
1!
1%
1-
12
#801480000000
0!
0%
b10 *
0-
02
b10 6
#801490000000
1!
1%
1-
12
#801500000000
0!
0%
b11 *
0-
02
b11 6
#801510000000
1!
1%
1-
12
15
#801520000000
0!
0%
b100 *
0-
02
b100 6
#801530000000
1!
1%
1-
12
#801540000000
0!
0%
b101 *
0-
02
b101 6
#801550000000
1!
1%
1-
12
#801560000000
0!
0%
b110 *
0-
02
b110 6
#801570000000
1!
1%
1-
12
#801580000000
0!
0%
b111 *
0-
02
b111 6
#801590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#801600000000
0!
0%
b0 *
0-
02
b0 6
#801610000000
1!
1%
1-
12
#801620000000
0!
0%
b1 *
0-
02
b1 6
#801630000000
1!
1%
1-
12
#801640000000
0!
0%
b10 *
0-
02
b10 6
#801650000000
1!
1%
1-
12
#801660000000
0!
0%
b11 *
0-
02
b11 6
#801670000000
1!
1%
1-
12
15
#801680000000
0!
0%
b100 *
0-
02
b100 6
#801690000000
1!
1%
1-
12
#801700000000
0!
0%
b101 *
0-
02
b101 6
#801710000000
1!
1%
1-
12
#801720000000
0!
0%
b110 *
0-
02
b110 6
#801730000000
1!
1%
1-
12
#801740000000
0!
0%
b111 *
0-
02
b111 6
#801750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#801760000000
0!
0%
b0 *
0-
02
b0 6
#801770000000
1!
1%
1-
12
#801780000000
0!
0%
b1 *
0-
02
b1 6
#801790000000
1!
1%
1-
12
#801800000000
0!
0%
b10 *
0-
02
b10 6
#801810000000
1!
1%
1-
12
#801820000000
0!
0%
b11 *
0-
02
b11 6
#801830000000
1!
1%
1-
12
15
#801840000000
0!
0%
b100 *
0-
02
b100 6
#801850000000
1!
1%
1-
12
#801860000000
0!
0%
b101 *
0-
02
b101 6
#801870000000
1!
1%
1-
12
#801880000000
0!
0%
b110 *
0-
02
b110 6
#801890000000
1!
1%
1-
12
#801900000000
0!
0%
b111 *
0-
02
b111 6
#801910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#801920000000
0!
0%
b0 *
0-
02
b0 6
#801930000000
1!
1%
1-
12
#801940000000
0!
0%
b1 *
0-
02
b1 6
#801950000000
1!
1%
1-
12
#801960000000
0!
0%
b10 *
0-
02
b10 6
#801970000000
1!
1%
1-
12
#801980000000
0!
0%
b11 *
0-
02
b11 6
#801990000000
1!
1%
1-
12
15
#802000000000
0!
0%
b100 *
0-
02
b100 6
#802010000000
1!
1%
1-
12
#802020000000
0!
0%
b101 *
0-
02
b101 6
#802030000000
1!
1%
1-
12
#802040000000
0!
0%
b110 *
0-
02
b110 6
#802050000000
1!
1%
1-
12
#802060000000
0!
0%
b111 *
0-
02
b111 6
#802070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#802080000000
0!
0%
b0 *
0-
02
b0 6
#802090000000
1!
1%
1-
12
#802100000000
0!
0%
b1 *
0-
02
b1 6
#802110000000
1!
1%
1-
12
#802120000000
0!
0%
b10 *
0-
02
b10 6
#802130000000
1!
1%
1-
12
#802140000000
0!
0%
b11 *
0-
02
b11 6
#802150000000
1!
1%
1-
12
15
#802160000000
0!
0%
b100 *
0-
02
b100 6
#802170000000
1!
1%
1-
12
#802180000000
0!
0%
b101 *
0-
02
b101 6
#802190000000
1!
1%
1-
12
#802200000000
0!
0%
b110 *
0-
02
b110 6
#802210000000
1!
1%
1-
12
#802220000000
0!
0%
b111 *
0-
02
b111 6
#802230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#802240000000
0!
0%
b0 *
0-
02
b0 6
#802250000000
1!
1%
1-
12
#802260000000
0!
0%
b1 *
0-
02
b1 6
#802270000000
1!
1%
1-
12
#802280000000
0!
0%
b10 *
0-
02
b10 6
#802290000000
1!
1%
1-
12
#802300000000
0!
0%
b11 *
0-
02
b11 6
#802310000000
1!
1%
1-
12
15
#802320000000
0!
0%
b100 *
0-
02
b100 6
#802330000000
1!
1%
1-
12
#802340000000
0!
0%
b101 *
0-
02
b101 6
#802350000000
1!
1%
1-
12
#802360000000
0!
0%
b110 *
0-
02
b110 6
#802370000000
1!
1%
1-
12
#802380000000
0!
0%
b111 *
0-
02
b111 6
#802390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#802400000000
0!
0%
b0 *
0-
02
b0 6
#802410000000
1!
1%
1-
12
#802420000000
0!
0%
b1 *
0-
02
b1 6
#802430000000
1!
1%
1-
12
#802440000000
0!
0%
b10 *
0-
02
b10 6
#802450000000
1!
1%
1-
12
#802460000000
0!
0%
b11 *
0-
02
b11 6
#802470000000
1!
1%
1-
12
15
#802480000000
0!
0%
b100 *
0-
02
b100 6
#802490000000
1!
1%
1-
12
#802500000000
0!
0%
b101 *
0-
02
b101 6
#802510000000
1!
1%
1-
12
#802520000000
0!
0%
b110 *
0-
02
b110 6
#802530000000
1!
1%
1-
12
#802540000000
0!
0%
b111 *
0-
02
b111 6
#802550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#802560000000
0!
0%
b0 *
0-
02
b0 6
#802570000000
1!
1%
1-
12
#802580000000
0!
0%
b1 *
0-
02
b1 6
#802590000000
1!
1%
1-
12
#802600000000
0!
0%
b10 *
0-
02
b10 6
#802610000000
1!
1%
1-
12
#802620000000
0!
0%
b11 *
0-
02
b11 6
#802630000000
1!
1%
1-
12
15
#802640000000
0!
0%
b100 *
0-
02
b100 6
#802650000000
1!
1%
1-
12
#802660000000
0!
0%
b101 *
0-
02
b101 6
#802670000000
1!
1%
1-
12
#802680000000
0!
0%
b110 *
0-
02
b110 6
#802690000000
1!
1%
1-
12
#802700000000
0!
0%
b111 *
0-
02
b111 6
#802710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#802720000000
0!
0%
b0 *
0-
02
b0 6
#802730000000
1!
1%
1-
12
#802740000000
0!
0%
b1 *
0-
02
b1 6
#802750000000
1!
1%
1-
12
#802760000000
0!
0%
b10 *
0-
02
b10 6
#802770000000
1!
1%
1-
12
#802780000000
0!
0%
b11 *
0-
02
b11 6
#802790000000
1!
1%
1-
12
15
#802800000000
0!
0%
b100 *
0-
02
b100 6
#802810000000
1!
1%
1-
12
#802820000000
0!
0%
b101 *
0-
02
b101 6
#802830000000
1!
1%
1-
12
#802840000000
0!
0%
b110 *
0-
02
b110 6
#802850000000
1!
1%
1-
12
#802860000000
0!
0%
b111 *
0-
02
b111 6
#802870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#802880000000
0!
0%
b0 *
0-
02
b0 6
#802890000000
1!
1%
1-
12
#802900000000
0!
0%
b1 *
0-
02
b1 6
#802910000000
1!
1%
1-
12
#802920000000
0!
0%
b10 *
0-
02
b10 6
#802930000000
1!
1%
1-
12
#802940000000
0!
0%
b11 *
0-
02
b11 6
#802950000000
1!
1%
1-
12
15
#802960000000
0!
0%
b100 *
0-
02
b100 6
#802970000000
1!
1%
1-
12
#802980000000
0!
0%
b101 *
0-
02
b101 6
#802990000000
1!
1%
1-
12
#803000000000
0!
0%
b110 *
0-
02
b110 6
#803010000000
1!
1%
1-
12
#803020000000
0!
0%
b111 *
0-
02
b111 6
#803030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#803040000000
0!
0%
b0 *
0-
02
b0 6
#803050000000
1!
1%
1-
12
#803060000000
0!
0%
b1 *
0-
02
b1 6
#803070000000
1!
1%
1-
12
#803080000000
0!
0%
b10 *
0-
02
b10 6
#803090000000
1!
1%
1-
12
#803100000000
0!
0%
b11 *
0-
02
b11 6
#803110000000
1!
1%
1-
12
15
#803120000000
0!
0%
b100 *
0-
02
b100 6
#803130000000
1!
1%
1-
12
#803140000000
0!
0%
b101 *
0-
02
b101 6
#803150000000
1!
1%
1-
12
#803160000000
0!
0%
b110 *
0-
02
b110 6
#803170000000
1!
1%
1-
12
#803180000000
0!
0%
b111 *
0-
02
b111 6
#803190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#803200000000
0!
0%
b0 *
0-
02
b0 6
#803210000000
1!
1%
1-
12
#803220000000
0!
0%
b1 *
0-
02
b1 6
#803230000000
1!
1%
1-
12
#803240000000
0!
0%
b10 *
0-
02
b10 6
#803250000000
1!
1%
1-
12
#803260000000
0!
0%
b11 *
0-
02
b11 6
#803270000000
1!
1%
1-
12
15
#803280000000
0!
0%
b100 *
0-
02
b100 6
#803290000000
1!
1%
1-
12
#803300000000
0!
0%
b101 *
0-
02
b101 6
#803310000000
1!
1%
1-
12
#803320000000
0!
0%
b110 *
0-
02
b110 6
#803330000000
1!
1%
1-
12
#803340000000
0!
0%
b111 *
0-
02
b111 6
#803350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#803360000000
0!
0%
b0 *
0-
02
b0 6
#803370000000
1!
1%
1-
12
#803380000000
0!
0%
b1 *
0-
02
b1 6
#803390000000
1!
1%
1-
12
#803400000000
0!
0%
b10 *
0-
02
b10 6
#803410000000
1!
1%
1-
12
#803420000000
0!
0%
b11 *
0-
02
b11 6
#803430000000
1!
1%
1-
12
15
#803440000000
0!
0%
b100 *
0-
02
b100 6
#803450000000
1!
1%
1-
12
#803460000000
0!
0%
b101 *
0-
02
b101 6
#803470000000
1!
1%
1-
12
#803480000000
0!
0%
b110 *
0-
02
b110 6
#803490000000
1!
1%
1-
12
#803500000000
0!
0%
b111 *
0-
02
b111 6
#803510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#803520000000
0!
0%
b0 *
0-
02
b0 6
#803530000000
1!
1%
1-
12
#803540000000
0!
0%
b1 *
0-
02
b1 6
#803550000000
1!
1%
1-
12
#803560000000
0!
0%
b10 *
0-
02
b10 6
#803570000000
1!
1%
1-
12
#803580000000
0!
0%
b11 *
0-
02
b11 6
#803590000000
1!
1%
1-
12
15
#803600000000
0!
0%
b100 *
0-
02
b100 6
#803610000000
1!
1%
1-
12
#803620000000
0!
0%
b101 *
0-
02
b101 6
#803630000000
1!
1%
1-
12
#803640000000
0!
0%
b110 *
0-
02
b110 6
#803650000000
1!
1%
1-
12
#803660000000
0!
0%
b111 *
0-
02
b111 6
#803670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#803680000000
0!
0%
b0 *
0-
02
b0 6
#803690000000
1!
1%
1-
12
#803700000000
0!
0%
b1 *
0-
02
b1 6
#803710000000
1!
1%
1-
12
#803720000000
0!
0%
b10 *
0-
02
b10 6
#803730000000
1!
1%
1-
12
#803740000000
0!
0%
b11 *
0-
02
b11 6
#803750000000
1!
1%
1-
12
15
#803760000000
0!
0%
b100 *
0-
02
b100 6
#803770000000
1!
1%
1-
12
#803780000000
0!
0%
b101 *
0-
02
b101 6
#803790000000
1!
1%
1-
12
#803800000000
0!
0%
b110 *
0-
02
b110 6
#803810000000
1!
1%
1-
12
#803820000000
0!
0%
b111 *
0-
02
b111 6
#803830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#803840000000
0!
0%
b0 *
0-
02
b0 6
#803850000000
1!
1%
1-
12
#803860000000
0!
0%
b1 *
0-
02
b1 6
#803870000000
1!
1%
1-
12
#803880000000
0!
0%
b10 *
0-
02
b10 6
#803890000000
1!
1%
1-
12
#803900000000
0!
0%
b11 *
0-
02
b11 6
#803910000000
1!
1%
1-
12
15
#803920000000
0!
0%
b100 *
0-
02
b100 6
#803930000000
1!
1%
1-
12
#803940000000
0!
0%
b101 *
0-
02
b101 6
#803950000000
1!
1%
1-
12
#803960000000
0!
0%
b110 *
0-
02
b110 6
#803970000000
1!
1%
1-
12
#803980000000
0!
0%
b111 *
0-
02
b111 6
#803990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#804000000000
0!
0%
b0 *
0-
02
b0 6
#804010000000
1!
1%
1-
12
#804020000000
0!
0%
b1 *
0-
02
b1 6
#804030000000
1!
1%
1-
12
#804040000000
0!
0%
b10 *
0-
02
b10 6
#804050000000
1!
1%
1-
12
#804060000000
0!
0%
b11 *
0-
02
b11 6
#804070000000
1!
1%
1-
12
15
#804080000000
0!
0%
b100 *
0-
02
b100 6
#804090000000
1!
1%
1-
12
#804100000000
0!
0%
b101 *
0-
02
b101 6
#804110000000
1!
1%
1-
12
#804120000000
0!
0%
b110 *
0-
02
b110 6
#804130000000
1!
1%
1-
12
#804140000000
0!
0%
b111 *
0-
02
b111 6
#804150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#804160000000
0!
0%
b0 *
0-
02
b0 6
#804170000000
1!
1%
1-
12
#804180000000
0!
0%
b1 *
0-
02
b1 6
#804190000000
1!
1%
1-
12
#804200000000
0!
0%
b10 *
0-
02
b10 6
#804210000000
1!
1%
1-
12
#804220000000
0!
0%
b11 *
0-
02
b11 6
#804230000000
1!
1%
1-
12
15
#804240000000
0!
0%
b100 *
0-
02
b100 6
#804250000000
1!
1%
1-
12
#804260000000
0!
0%
b101 *
0-
02
b101 6
#804270000000
1!
1%
1-
12
#804280000000
0!
0%
b110 *
0-
02
b110 6
#804290000000
1!
1%
1-
12
#804300000000
0!
0%
b111 *
0-
02
b111 6
#804310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#804320000000
0!
0%
b0 *
0-
02
b0 6
#804330000000
1!
1%
1-
12
#804340000000
0!
0%
b1 *
0-
02
b1 6
#804350000000
1!
1%
1-
12
#804360000000
0!
0%
b10 *
0-
02
b10 6
#804370000000
1!
1%
1-
12
#804380000000
0!
0%
b11 *
0-
02
b11 6
#804390000000
1!
1%
1-
12
15
#804400000000
0!
0%
b100 *
0-
02
b100 6
#804410000000
1!
1%
1-
12
#804420000000
0!
0%
b101 *
0-
02
b101 6
#804430000000
1!
1%
1-
12
#804440000000
0!
0%
b110 *
0-
02
b110 6
#804450000000
1!
1%
1-
12
#804460000000
0!
0%
b111 *
0-
02
b111 6
#804470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#804480000000
0!
0%
b0 *
0-
02
b0 6
#804490000000
1!
1%
1-
12
#804500000000
0!
0%
b1 *
0-
02
b1 6
#804510000000
1!
1%
1-
12
#804520000000
0!
0%
b10 *
0-
02
b10 6
#804530000000
1!
1%
1-
12
#804540000000
0!
0%
b11 *
0-
02
b11 6
#804550000000
1!
1%
1-
12
15
#804560000000
0!
0%
b100 *
0-
02
b100 6
#804570000000
1!
1%
1-
12
#804580000000
0!
0%
b101 *
0-
02
b101 6
#804590000000
1!
1%
1-
12
#804600000000
0!
0%
b110 *
0-
02
b110 6
#804610000000
1!
1%
1-
12
#804620000000
0!
0%
b111 *
0-
02
b111 6
#804630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#804640000000
0!
0%
b0 *
0-
02
b0 6
#804650000000
1!
1%
1-
12
#804660000000
0!
0%
b1 *
0-
02
b1 6
#804670000000
1!
1%
1-
12
#804680000000
0!
0%
b10 *
0-
02
b10 6
#804690000000
1!
1%
1-
12
#804700000000
0!
0%
b11 *
0-
02
b11 6
#804710000000
1!
1%
1-
12
15
#804720000000
0!
0%
b100 *
0-
02
b100 6
#804730000000
1!
1%
1-
12
#804740000000
0!
0%
b101 *
0-
02
b101 6
#804750000000
1!
1%
1-
12
#804760000000
0!
0%
b110 *
0-
02
b110 6
#804770000000
1!
1%
1-
12
#804780000000
0!
0%
b111 *
0-
02
b111 6
#804790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#804800000000
0!
0%
b0 *
0-
02
b0 6
#804810000000
1!
1%
1-
12
#804820000000
0!
0%
b1 *
0-
02
b1 6
#804830000000
1!
1%
1-
12
#804840000000
0!
0%
b10 *
0-
02
b10 6
#804850000000
1!
1%
1-
12
#804860000000
0!
0%
b11 *
0-
02
b11 6
#804870000000
1!
1%
1-
12
15
#804880000000
0!
0%
b100 *
0-
02
b100 6
#804890000000
1!
1%
1-
12
#804900000000
0!
0%
b101 *
0-
02
b101 6
#804910000000
1!
1%
1-
12
#804920000000
0!
0%
b110 *
0-
02
b110 6
#804930000000
1!
1%
1-
12
#804940000000
0!
0%
b111 *
0-
02
b111 6
#804950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#804960000000
0!
0%
b0 *
0-
02
b0 6
#804970000000
1!
1%
1-
12
#804980000000
0!
0%
b1 *
0-
02
b1 6
#804990000000
1!
1%
1-
12
#805000000000
0!
0%
b10 *
0-
02
b10 6
#805010000000
1!
1%
1-
12
#805020000000
0!
0%
b11 *
0-
02
b11 6
#805030000000
1!
1%
1-
12
15
#805040000000
0!
0%
b100 *
0-
02
b100 6
#805050000000
1!
1%
1-
12
#805060000000
0!
0%
b101 *
0-
02
b101 6
#805070000000
1!
1%
1-
12
#805080000000
0!
0%
b110 *
0-
02
b110 6
#805090000000
1!
1%
1-
12
#805100000000
0!
0%
b111 *
0-
02
b111 6
#805110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#805120000000
0!
0%
b0 *
0-
02
b0 6
#805130000000
1!
1%
1-
12
#805140000000
0!
0%
b1 *
0-
02
b1 6
#805150000000
1!
1%
1-
12
#805160000000
0!
0%
b10 *
0-
02
b10 6
#805170000000
1!
1%
1-
12
#805180000000
0!
0%
b11 *
0-
02
b11 6
#805190000000
1!
1%
1-
12
15
#805200000000
0!
0%
b100 *
0-
02
b100 6
#805210000000
1!
1%
1-
12
#805220000000
0!
0%
b101 *
0-
02
b101 6
#805230000000
1!
1%
1-
12
#805240000000
0!
0%
b110 *
0-
02
b110 6
#805250000000
1!
1%
1-
12
#805260000000
0!
0%
b111 *
0-
02
b111 6
#805270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#805280000000
0!
0%
b0 *
0-
02
b0 6
#805290000000
1!
1%
1-
12
#805300000000
0!
0%
b1 *
0-
02
b1 6
#805310000000
1!
1%
1-
12
#805320000000
0!
0%
b10 *
0-
02
b10 6
#805330000000
1!
1%
1-
12
#805340000000
0!
0%
b11 *
0-
02
b11 6
#805350000000
1!
1%
1-
12
15
#805360000000
0!
0%
b100 *
0-
02
b100 6
#805370000000
1!
1%
1-
12
#805380000000
0!
0%
b101 *
0-
02
b101 6
#805390000000
1!
1%
1-
12
#805400000000
0!
0%
b110 *
0-
02
b110 6
#805410000000
1!
1%
1-
12
#805420000000
0!
0%
b111 *
0-
02
b111 6
#805430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#805440000000
0!
0%
b0 *
0-
02
b0 6
#805450000000
1!
1%
1-
12
#805460000000
0!
0%
b1 *
0-
02
b1 6
#805470000000
1!
1%
1-
12
#805480000000
0!
0%
b10 *
0-
02
b10 6
#805490000000
1!
1%
1-
12
#805500000000
0!
0%
b11 *
0-
02
b11 6
#805510000000
1!
1%
1-
12
15
#805520000000
0!
0%
b100 *
0-
02
b100 6
#805530000000
1!
1%
1-
12
#805540000000
0!
0%
b101 *
0-
02
b101 6
#805550000000
1!
1%
1-
12
#805560000000
0!
0%
b110 *
0-
02
b110 6
#805570000000
1!
1%
1-
12
#805580000000
0!
0%
b111 *
0-
02
b111 6
#805590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#805600000000
0!
0%
b0 *
0-
02
b0 6
#805610000000
1!
1%
1-
12
#805620000000
0!
0%
b1 *
0-
02
b1 6
#805630000000
1!
1%
1-
12
#805640000000
0!
0%
b10 *
0-
02
b10 6
#805650000000
1!
1%
1-
12
#805660000000
0!
0%
b11 *
0-
02
b11 6
#805670000000
1!
1%
1-
12
15
#805680000000
0!
0%
b100 *
0-
02
b100 6
#805690000000
1!
1%
1-
12
#805700000000
0!
0%
b101 *
0-
02
b101 6
#805710000000
1!
1%
1-
12
#805720000000
0!
0%
b110 *
0-
02
b110 6
#805730000000
1!
1%
1-
12
#805740000000
0!
0%
b111 *
0-
02
b111 6
#805750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#805760000000
0!
0%
b0 *
0-
02
b0 6
#805770000000
1!
1%
1-
12
#805780000000
0!
0%
b1 *
0-
02
b1 6
#805790000000
1!
1%
1-
12
#805800000000
0!
0%
b10 *
0-
02
b10 6
#805810000000
1!
1%
1-
12
#805820000000
0!
0%
b11 *
0-
02
b11 6
#805830000000
1!
1%
1-
12
15
#805840000000
0!
0%
b100 *
0-
02
b100 6
#805850000000
1!
1%
1-
12
#805860000000
0!
0%
b101 *
0-
02
b101 6
#805870000000
1!
1%
1-
12
#805880000000
0!
0%
b110 *
0-
02
b110 6
#805890000000
1!
1%
1-
12
#805900000000
0!
0%
b111 *
0-
02
b111 6
#805910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#805920000000
0!
0%
b0 *
0-
02
b0 6
#805930000000
1!
1%
1-
12
#805940000000
0!
0%
b1 *
0-
02
b1 6
#805950000000
1!
1%
1-
12
#805960000000
0!
0%
b10 *
0-
02
b10 6
#805970000000
1!
1%
1-
12
#805980000000
0!
0%
b11 *
0-
02
b11 6
#805990000000
1!
1%
1-
12
15
#806000000000
0!
0%
b100 *
0-
02
b100 6
#806010000000
1!
1%
1-
12
#806020000000
0!
0%
b101 *
0-
02
b101 6
#806030000000
1!
1%
1-
12
#806040000000
0!
0%
b110 *
0-
02
b110 6
#806050000000
1!
1%
1-
12
#806060000000
0!
0%
b111 *
0-
02
b111 6
#806070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#806080000000
0!
0%
b0 *
0-
02
b0 6
#806090000000
1!
1%
1-
12
#806100000000
0!
0%
b1 *
0-
02
b1 6
#806110000000
1!
1%
1-
12
#806120000000
0!
0%
b10 *
0-
02
b10 6
#806130000000
1!
1%
1-
12
#806140000000
0!
0%
b11 *
0-
02
b11 6
#806150000000
1!
1%
1-
12
15
#806160000000
0!
0%
b100 *
0-
02
b100 6
#806170000000
1!
1%
1-
12
#806180000000
0!
0%
b101 *
0-
02
b101 6
#806190000000
1!
1%
1-
12
#806200000000
0!
0%
b110 *
0-
02
b110 6
#806210000000
1!
1%
1-
12
#806220000000
0!
0%
b111 *
0-
02
b111 6
#806230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#806240000000
0!
0%
b0 *
0-
02
b0 6
#806250000000
1!
1%
1-
12
#806260000000
0!
0%
b1 *
0-
02
b1 6
#806270000000
1!
1%
1-
12
#806280000000
0!
0%
b10 *
0-
02
b10 6
#806290000000
1!
1%
1-
12
#806300000000
0!
0%
b11 *
0-
02
b11 6
#806310000000
1!
1%
1-
12
15
#806320000000
0!
0%
b100 *
0-
02
b100 6
#806330000000
1!
1%
1-
12
#806340000000
0!
0%
b101 *
0-
02
b101 6
#806350000000
1!
1%
1-
12
#806360000000
0!
0%
b110 *
0-
02
b110 6
#806370000000
1!
1%
1-
12
#806380000000
0!
0%
b111 *
0-
02
b111 6
#806390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#806400000000
0!
0%
b0 *
0-
02
b0 6
#806410000000
1!
1%
1-
12
#806420000000
0!
0%
b1 *
0-
02
b1 6
#806430000000
1!
1%
1-
12
#806440000000
0!
0%
b10 *
0-
02
b10 6
#806450000000
1!
1%
1-
12
#806460000000
0!
0%
b11 *
0-
02
b11 6
#806470000000
1!
1%
1-
12
15
#806480000000
0!
0%
b100 *
0-
02
b100 6
#806490000000
1!
1%
1-
12
#806500000000
0!
0%
b101 *
0-
02
b101 6
#806510000000
1!
1%
1-
12
#806520000000
0!
0%
b110 *
0-
02
b110 6
#806530000000
1!
1%
1-
12
#806540000000
0!
0%
b111 *
0-
02
b111 6
#806550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#806560000000
0!
0%
b0 *
0-
02
b0 6
#806570000000
1!
1%
1-
12
#806580000000
0!
0%
b1 *
0-
02
b1 6
#806590000000
1!
1%
1-
12
#806600000000
0!
0%
b10 *
0-
02
b10 6
#806610000000
1!
1%
1-
12
#806620000000
0!
0%
b11 *
0-
02
b11 6
#806630000000
1!
1%
1-
12
15
#806640000000
0!
0%
b100 *
0-
02
b100 6
#806650000000
1!
1%
1-
12
#806660000000
0!
0%
b101 *
0-
02
b101 6
#806670000000
1!
1%
1-
12
#806680000000
0!
0%
b110 *
0-
02
b110 6
#806690000000
1!
1%
1-
12
#806700000000
0!
0%
b111 *
0-
02
b111 6
#806710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#806720000000
0!
0%
b0 *
0-
02
b0 6
#806730000000
1!
1%
1-
12
#806740000000
0!
0%
b1 *
0-
02
b1 6
#806750000000
1!
1%
1-
12
#806760000000
0!
0%
b10 *
0-
02
b10 6
#806770000000
1!
1%
1-
12
#806780000000
0!
0%
b11 *
0-
02
b11 6
#806790000000
1!
1%
1-
12
15
#806800000000
0!
0%
b100 *
0-
02
b100 6
#806810000000
1!
1%
1-
12
#806820000000
0!
0%
b101 *
0-
02
b101 6
#806830000000
1!
1%
1-
12
#806840000000
0!
0%
b110 *
0-
02
b110 6
#806850000000
1!
1%
1-
12
#806860000000
0!
0%
b111 *
0-
02
b111 6
#806870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#806880000000
0!
0%
b0 *
0-
02
b0 6
#806890000000
1!
1%
1-
12
#806900000000
0!
0%
b1 *
0-
02
b1 6
#806910000000
1!
1%
1-
12
#806920000000
0!
0%
b10 *
0-
02
b10 6
#806930000000
1!
1%
1-
12
#806940000000
0!
0%
b11 *
0-
02
b11 6
#806950000000
1!
1%
1-
12
15
#806960000000
0!
0%
b100 *
0-
02
b100 6
#806970000000
1!
1%
1-
12
#806980000000
0!
0%
b101 *
0-
02
b101 6
#806990000000
1!
1%
1-
12
#807000000000
0!
0%
b110 *
0-
02
b110 6
#807010000000
1!
1%
1-
12
#807020000000
0!
0%
b111 *
0-
02
b111 6
#807030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#807040000000
0!
0%
b0 *
0-
02
b0 6
#807050000000
1!
1%
1-
12
#807060000000
0!
0%
b1 *
0-
02
b1 6
#807070000000
1!
1%
1-
12
#807080000000
0!
0%
b10 *
0-
02
b10 6
#807090000000
1!
1%
1-
12
#807100000000
0!
0%
b11 *
0-
02
b11 6
#807110000000
1!
1%
1-
12
15
#807120000000
0!
0%
b100 *
0-
02
b100 6
#807130000000
1!
1%
1-
12
#807140000000
0!
0%
b101 *
0-
02
b101 6
#807150000000
1!
1%
1-
12
#807160000000
0!
0%
b110 *
0-
02
b110 6
#807170000000
1!
1%
1-
12
#807180000000
0!
0%
b111 *
0-
02
b111 6
#807190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#807200000000
0!
0%
b0 *
0-
02
b0 6
#807210000000
1!
1%
1-
12
#807220000000
0!
0%
b1 *
0-
02
b1 6
#807230000000
1!
1%
1-
12
#807240000000
0!
0%
b10 *
0-
02
b10 6
#807250000000
1!
1%
1-
12
#807260000000
0!
0%
b11 *
0-
02
b11 6
#807270000000
1!
1%
1-
12
15
#807280000000
0!
0%
b100 *
0-
02
b100 6
#807290000000
1!
1%
1-
12
#807300000000
0!
0%
b101 *
0-
02
b101 6
#807310000000
1!
1%
1-
12
#807320000000
0!
0%
b110 *
0-
02
b110 6
#807330000000
1!
1%
1-
12
#807340000000
0!
0%
b111 *
0-
02
b111 6
#807350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#807360000000
0!
0%
b0 *
0-
02
b0 6
#807370000000
1!
1%
1-
12
#807380000000
0!
0%
b1 *
0-
02
b1 6
#807390000000
1!
1%
1-
12
#807400000000
0!
0%
b10 *
0-
02
b10 6
#807410000000
1!
1%
1-
12
#807420000000
0!
0%
b11 *
0-
02
b11 6
#807430000000
1!
1%
1-
12
15
#807440000000
0!
0%
b100 *
0-
02
b100 6
#807450000000
1!
1%
1-
12
#807460000000
0!
0%
b101 *
0-
02
b101 6
#807470000000
1!
1%
1-
12
#807480000000
0!
0%
b110 *
0-
02
b110 6
#807490000000
1!
1%
1-
12
#807500000000
0!
0%
b111 *
0-
02
b111 6
#807510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#807520000000
0!
0%
b0 *
0-
02
b0 6
#807530000000
1!
1%
1-
12
#807540000000
0!
0%
b1 *
0-
02
b1 6
#807550000000
1!
1%
1-
12
#807560000000
0!
0%
b10 *
0-
02
b10 6
#807570000000
1!
1%
1-
12
#807580000000
0!
0%
b11 *
0-
02
b11 6
#807590000000
1!
1%
1-
12
15
#807600000000
0!
0%
b100 *
0-
02
b100 6
#807610000000
1!
1%
1-
12
#807620000000
0!
0%
b101 *
0-
02
b101 6
#807630000000
1!
1%
1-
12
#807640000000
0!
0%
b110 *
0-
02
b110 6
#807650000000
1!
1%
1-
12
#807660000000
0!
0%
b111 *
0-
02
b111 6
#807670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#807680000000
0!
0%
b0 *
0-
02
b0 6
#807690000000
1!
1%
1-
12
#807700000000
0!
0%
b1 *
0-
02
b1 6
#807710000000
1!
1%
1-
12
#807720000000
0!
0%
b10 *
0-
02
b10 6
#807730000000
1!
1%
1-
12
#807740000000
0!
0%
b11 *
0-
02
b11 6
#807750000000
1!
1%
1-
12
15
#807760000000
0!
0%
b100 *
0-
02
b100 6
#807770000000
1!
1%
1-
12
#807780000000
0!
0%
b101 *
0-
02
b101 6
#807790000000
1!
1%
1-
12
#807800000000
0!
0%
b110 *
0-
02
b110 6
#807810000000
1!
1%
1-
12
#807820000000
0!
0%
b111 *
0-
02
b111 6
#807830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#807840000000
0!
0%
b0 *
0-
02
b0 6
#807850000000
1!
1%
1-
12
#807860000000
0!
0%
b1 *
0-
02
b1 6
#807870000000
1!
1%
1-
12
#807880000000
0!
0%
b10 *
0-
02
b10 6
#807890000000
1!
1%
1-
12
#807900000000
0!
0%
b11 *
0-
02
b11 6
#807910000000
1!
1%
1-
12
15
#807920000000
0!
0%
b100 *
0-
02
b100 6
#807930000000
1!
1%
1-
12
#807940000000
0!
0%
b101 *
0-
02
b101 6
#807950000000
1!
1%
1-
12
#807960000000
0!
0%
b110 *
0-
02
b110 6
#807970000000
1!
1%
1-
12
#807980000000
0!
0%
b111 *
0-
02
b111 6
#807990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#808000000000
0!
0%
b0 *
0-
02
b0 6
#808010000000
1!
1%
1-
12
#808020000000
0!
0%
b1 *
0-
02
b1 6
#808030000000
1!
1%
1-
12
#808040000000
0!
0%
b10 *
0-
02
b10 6
#808050000000
1!
1%
1-
12
#808060000000
0!
0%
b11 *
0-
02
b11 6
#808070000000
1!
1%
1-
12
15
#808080000000
0!
0%
b100 *
0-
02
b100 6
#808090000000
1!
1%
1-
12
#808100000000
0!
0%
b101 *
0-
02
b101 6
#808110000000
1!
1%
1-
12
#808120000000
0!
0%
b110 *
0-
02
b110 6
#808130000000
1!
1%
1-
12
#808140000000
0!
0%
b111 *
0-
02
b111 6
#808150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#808160000000
0!
0%
b0 *
0-
02
b0 6
#808170000000
1!
1%
1-
12
#808180000000
0!
0%
b1 *
0-
02
b1 6
#808190000000
1!
1%
1-
12
#808200000000
0!
0%
b10 *
0-
02
b10 6
#808210000000
1!
1%
1-
12
#808220000000
0!
0%
b11 *
0-
02
b11 6
#808230000000
1!
1%
1-
12
15
#808240000000
0!
0%
b100 *
0-
02
b100 6
#808250000000
1!
1%
1-
12
#808260000000
0!
0%
b101 *
0-
02
b101 6
#808270000000
1!
1%
1-
12
#808280000000
0!
0%
b110 *
0-
02
b110 6
#808290000000
1!
1%
1-
12
#808300000000
0!
0%
b111 *
0-
02
b111 6
#808310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#808320000000
0!
0%
b0 *
0-
02
b0 6
#808330000000
1!
1%
1-
12
#808340000000
0!
0%
b1 *
0-
02
b1 6
#808350000000
1!
1%
1-
12
#808360000000
0!
0%
b10 *
0-
02
b10 6
#808370000000
1!
1%
1-
12
#808380000000
0!
0%
b11 *
0-
02
b11 6
#808390000000
1!
1%
1-
12
15
#808400000000
0!
0%
b100 *
0-
02
b100 6
#808410000000
1!
1%
1-
12
#808420000000
0!
0%
b101 *
0-
02
b101 6
#808430000000
1!
1%
1-
12
#808440000000
0!
0%
b110 *
0-
02
b110 6
#808450000000
1!
1%
1-
12
#808460000000
0!
0%
b111 *
0-
02
b111 6
#808470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#808480000000
0!
0%
b0 *
0-
02
b0 6
#808490000000
1!
1%
1-
12
#808500000000
0!
0%
b1 *
0-
02
b1 6
#808510000000
1!
1%
1-
12
#808520000000
0!
0%
b10 *
0-
02
b10 6
#808530000000
1!
1%
1-
12
#808540000000
0!
0%
b11 *
0-
02
b11 6
#808550000000
1!
1%
1-
12
15
#808560000000
0!
0%
b100 *
0-
02
b100 6
#808570000000
1!
1%
1-
12
#808580000000
0!
0%
b101 *
0-
02
b101 6
#808590000000
1!
1%
1-
12
#808600000000
0!
0%
b110 *
0-
02
b110 6
#808610000000
1!
1%
1-
12
#808620000000
0!
0%
b111 *
0-
02
b111 6
#808630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#808640000000
0!
0%
b0 *
0-
02
b0 6
#808650000000
1!
1%
1-
12
#808660000000
0!
0%
b1 *
0-
02
b1 6
#808670000000
1!
1%
1-
12
#808680000000
0!
0%
b10 *
0-
02
b10 6
#808690000000
1!
1%
1-
12
#808700000000
0!
0%
b11 *
0-
02
b11 6
#808710000000
1!
1%
1-
12
15
#808720000000
0!
0%
b100 *
0-
02
b100 6
#808730000000
1!
1%
1-
12
#808740000000
0!
0%
b101 *
0-
02
b101 6
#808750000000
1!
1%
1-
12
#808760000000
0!
0%
b110 *
0-
02
b110 6
#808770000000
1!
1%
1-
12
#808780000000
0!
0%
b111 *
0-
02
b111 6
#808790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#808800000000
0!
0%
b0 *
0-
02
b0 6
#808810000000
1!
1%
1-
12
#808820000000
0!
0%
b1 *
0-
02
b1 6
#808830000000
1!
1%
1-
12
#808840000000
0!
0%
b10 *
0-
02
b10 6
#808850000000
1!
1%
1-
12
#808860000000
0!
0%
b11 *
0-
02
b11 6
#808870000000
1!
1%
1-
12
15
#808880000000
0!
0%
b100 *
0-
02
b100 6
#808890000000
1!
1%
1-
12
#808900000000
0!
0%
b101 *
0-
02
b101 6
#808910000000
1!
1%
1-
12
#808920000000
0!
0%
b110 *
0-
02
b110 6
#808930000000
1!
1%
1-
12
#808940000000
0!
0%
b111 *
0-
02
b111 6
#808950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#808960000000
0!
0%
b0 *
0-
02
b0 6
#808970000000
1!
1%
1-
12
#808980000000
0!
0%
b1 *
0-
02
b1 6
#808990000000
1!
1%
1-
12
#809000000000
0!
0%
b10 *
0-
02
b10 6
#809010000000
1!
1%
1-
12
#809020000000
0!
0%
b11 *
0-
02
b11 6
#809030000000
1!
1%
1-
12
15
#809040000000
0!
0%
b100 *
0-
02
b100 6
#809050000000
1!
1%
1-
12
#809060000000
0!
0%
b101 *
0-
02
b101 6
#809070000000
1!
1%
1-
12
#809080000000
0!
0%
b110 *
0-
02
b110 6
#809090000000
1!
1%
1-
12
#809100000000
0!
0%
b111 *
0-
02
b111 6
#809110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#809120000000
0!
0%
b0 *
0-
02
b0 6
#809130000000
1!
1%
1-
12
#809140000000
0!
0%
b1 *
0-
02
b1 6
#809150000000
1!
1%
1-
12
#809160000000
0!
0%
b10 *
0-
02
b10 6
#809170000000
1!
1%
1-
12
#809180000000
0!
0%
b11 *
0-
02
b11 6
#809190000000
1!
1%
1-
12
15
#809200000000
0!
0%
b100 *
0-
02
b100 6
#809210000000
1!
1%
1-
12
#809220000000
0!
0%
b101 *
0-
02
b101 6
#809230000000
1!
1%
1-
12
#809240000000
0!
0%
b110 *
0-
02
b110 6
#809250000000
1!
1%
1-
12
#809260000000
0!
0%
b111 *
0-
02
b111 6
#809270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#809280000000
0!
0%
b0 *
0-
02
b0 6
#809290000000
1!
1%
1-
12
#809300000000
0!
0%
b1 *
0-
02
b1 6
#809310000000
1!
1%
1-
12
#809320000000
0!
0%
b10 *
0-
02
b10 6
#809330000000
1!
1%
1-
12
#809340000000
0!
0%
b11 *
0-
02
b11 6
#809350000000
1!
1%
1-
12
15
#809360000000
0!
0%
b100 *
0-
02
b100 6
#809370000000
1!
1%
1-
12
#809380000000
0!
0%
b101 *
0-
02
b101 6
#809390000000
1!
1%
1-
12
#809400000000
0!
0%
b110 *
0-
02
b110 6
#809410000000
1!
1%
1-
12
#809420000000
0!
0%
b111 *
0-
02
b111 6
#809430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#809440000000
0!
0%
b0 *
0-
02
b0 6
#809450000000
1!
1%
1-
12
#809460000000
0!
0%
b1 *
0-
02
b1 6
#809470000000
1!
1%
1-
12
#809480000000
0!
0%
b10 *
0-
02
b10 6
#809490000000
1!
1%
1-
12
#809500000000
0!
0%
b11 *
0-
02
b11 6
#809510000000
1!
1%
1-
12
15
#809520000000
0!
0%
b100 *
0-
02
b100 6
#809530000000
1!
1%
1-
12
#809540000000
0!
0%
b101 *
0-
02
b101 6
#809550000000
1!
1%
1-
12
#809560000000
0!
0%
b110 *
0-
02
b110 6
#809570000000
1!
1%
1-
12
#809580000000
0!
0%
b111 *
0-
02
b111 6
#809590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#809600000000
0!
0%
b0 *
0-
02
b0 6
#809610000000
1!
1%
1-
12
#809620000000
0!
0%
b1 *
0-
02
b1 6
#809630000000
1!
1%
1-
12
#809640000000
0!
0%
b10 *
0-
02
b10 6
#809650000000
1!
1%
1-
12
#809660000000
0!
0%
b11 *
0-
02
b11 6
#809670000000
1!
1%
1-
12
15
#809680000000
0!
0%
b100 *
0-
02
b100 6
#809690000000
1!
1%
1-
12
#809700000000
0!
0%
b101 *
0-
02
b101 6
#809710000000
1!
1%
1-
12
#809720000000
0!
0%
b110 *
0-
02
b110 6
#809730000000
1!
1%
1-
12
#809740000000
0!
0%
b111 *
0-
02
b111 6
#809750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#809760000000
0!
0%
b0 *
0-
02
b0 6
#809770000000
1!
1%
1-
12
#809780000000
0!
0%
b1 *
0-
02
b1 6
#809790000000
1!
1%
1-
12
#809800000000
0!
0%
b10 *
0-
02
b10 6
#809810000000
1!
1%
1-
12
#809820000000
0!
0%
b11 *
0-
02
b11 6
#809830000000
1!
1%
1-
12
15
#809840000000
0!
0%
b100 *
0-
02
b100 6
#809850000000
1!
1%
1-
12
#809860000000
0!
0%
b101 *
0-
02
b101 6
#809870000000
1!
1%
1-
12
#809880000000
0!
0%
b110 *
0-
02
b110 6
#809890000000
1!
1%
1-
12
#809900000000
0!
0%
b111 *
0-
02
b111 6
#809910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#809920000000
0!
0%
b0 *
0-
02
b0 6
#809930000000
1!
1%
1-
12
#809940000000
0!
0%
b1 *
0-
02
b1 6
#809950000000
1!
1%
1-
12
#809960000000
0!
0%
b10 *
0-
02
b10 6
#809970000000
1!
1%
1-
12
#809980000000
0!
0%
b11 *
0-
02
b11 6
#809990000000
1!
1%
1-
12
15
#810000000000
0!
0%
b100 *
0-
02
b100 6
#810010000000
1!
1%
1-
12
#810020000000
0!
0%
b101 *
0-
02
b101 6
#810030000000
1!
1%
1-
12
#810040000000
0!
0%
b110 *
0-
02
b110 6
#810050000000
1!
1%
1-
12
#810060000000
0!
0%
b111 *
0-
02
b111 6
#810070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#810080000000
0!
0%
b0 *
0-
02
b0 6
#810090000000
1!
1%
1-
12
#810100000000
0!
0%
b1 *
0-
02
b1 6
#810110000000
1!
1%
1-
12
#810120000000
0!
0%
b10 *
0-
02
b10 6
#810130000000
1!
1%
1-
12
#810140000000
0!
0%
b11 *
0-
02
b11 6
#810150000000
1!
1%
1-
12
15
#810160000000
0!
0%
b100 *
0-
02
b100 6
#810170000000
1!
1%
1-
12
#810180000000
0!
0%
b101 *
0-
02
b101 6
#810190000000
1!
1%
1-
12
#810200000000
0!
0%
b110 *
0-
02
b110 6
#810210000000
1!
1%
1-
12
#810220000000
0!
0%
b111 *
0-
02
b111 6
#810230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#810240000000
0!
0%
b0 *
0-
02
b0 6
#810250000000
1!
1%
1-
12
#810260000000
0!
0%
b1 *
0-
02
b1 6
#810270000000
1!
1%
1-
12
#810280000000
0!
0%
b10 *
0-
02
b10 6
#810290000000
1!
1%
1-
12
#810300000000
0!
0%
b11 *
0-
02
b11 6
#810310000000
1!
1%
1-
12
15
#810320000000
0!
0%
b100 *
0-
02
b100 6
#810330000000
1!
1%
1-
12
#810340000000
0!
0%
b101 *
0-
02
b101 6
#810350000000
1!
1%
1-
12
#810360000000
0!
0%
b110 *
0-
02
b110 6
#810370000000
1!
1%
1-
12
#810380000000
0!
0%
b111 *
0-
02
b111 6
#810390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#810400000000
0!
0%
b0 *
0-
02
b0 6
#810410000000
1!
1%
1-
12
#810420000000
0!
0%
b1 *
0-
02
b1 6
#810430000000
1!
1%
1-
12
#810440000000
0!
0%
b10 *
0-
02
b10 6
#810450000000
1!
1%
1-
12
#810460000000
0!
0%
b11 *
0-
02
b11 6
#810470000000
1!
1%
1-
12
15
#810480000000
0!
0%
b100 *
0-
02
b100 6
#810490000000
1!
1%
1-
12
#810500000000
0!
0%
b101 *
0-
02
b101 6
#810510000000
1!
1%
1-
12
#810520000000
0!
0%
b110 *
0-
02
b110 6
#810530000000
1!
1%
1-
12
#810540000000
0!
0%
b111 *
0-
02
b111 6
#810550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#810560000000
0!
0%
b0 *
0-
02
b0 6
#810570000000
1!
1%
1-
12
#810580000000
0!
0%
b1 *
0-
02
b1 6
#810590000000
1!
1%
1-
12
#810600000000
0!
0%
b10 *
0-
02
b10 6
#810610000000
1!
1%
1-
12
#810620000000
0!
0%
b11 *
0-
02
b11 6
#810630000000
1!
1%
1-
12
15
#810640000000
0!
0%
b100 *
0-
02
b100 6
#810650000000
1!
1%
1-
12
#810660000000
0!
0%
b101 *
0-
02
b101 6
#810670000000
1!
1%
1-
12
#810680000000
0!
0%
b110 *
0-
02
b110 6
#810690000000
1!
1%
1-
12
#810700000000
0!
0%
b111 *
0-
02
b111 6
#810710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#810720000000
0!
0%
b0 *
0-
02
b0 6
#810730000000
1!
1%
1-
12
#810740000000
0!
0%
b1 *
0-
02
b1 6
#810750000000
1!
1%
1-
12
#810760000000
0!
0%
b10 *
0-
02
b10 6
#810770000000
1!
1%
1-
12
#810780000000
0!
0%
b11 *
0-
02
b11 6
#810790000000
1!
1%
1-
12
15
#810800000000
0!
0%
b100 *
0-
02
b100 6
#810810000000
1!
1%
1-
12
#810820000000
0!
0%
b101 *
0-
02
b101 6
#810830000000
1!
1%
1-
12
#810840000000
0!
0%
b110 *
0-
02
b110 6
#810850000000
1!
1%
1-
12
#810860000000
0!
0%
b111 *
0-
02
b111 6
#810870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#810880000000
0!
0%
b0 *
0-
02
b0 6
#810890000000
1!
1%
1-
12
#810900000000
0!
0%
b1 *
0-
02
b1 6
#810910000000
1!
1%
1-
12
#810920000000
0!
0%
b10 *
0-
02
b10 6
#810930000000
1!
1%
1-
12
#810940000000
0!
0%
b11 *
0-
02
b11 6
#810950000000
1!
1%
1-
12
15
#810960000000
0!
0%
b100 *
0-
02
b100 6
#810970000000
1!
1%
1-
12
#810980000000
0!
0%
b101 *
0-
02
b101 6
#810990000000
1!
1%
1-
12
#811000000000
0!
0%
b110 *
0-
02
b110 6
#811010000000
1!
1%
1-
12
#811020000000
0!
0%
b111 *
0-
02
b111 6
#811030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#811040000000
0!
0%
b0 *
0-
02
b0 6
#811050000000
1!
1%
1-
12
#811060000000
0!
0%
b1 *
0-
02
b1 6
#811070000000
1!
1%
1-
12
#811080000000
0!
0%
b10 *
0-
02
b10 6
#811090000000
1!
1%
1-
12
#811100000000
0!
0%
b11 *
0-
02
b11 6
#811110000000
1!
1%
1-
12
15
#811120000000
0!
0%
b100 *
0-
02
b100 6
#811130000000
1!
1%
1-
12
#811140000000
0!
0%
b101 *
0-
02
b101 6
#811150000000
1!
1%
1-
12
#811160000000
0!
0%
b110 *
0-
02
b110 6
#811170000000
1!
1%
1-
12
#811180000000
0!
0%
b111 *
0-
02
b111 6
#811190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#811200000000
0!
0%
b0 *
0-
02
b0 6
#811210000000
1!
1%
1-
12
#811220000000
0!
0%
b1 *
0-
02
b1 6
#811230000000
1!
1%
1-
12
#811240000000
0!
0%
b10 *
0-
02
b10 6
#811250000000
1!
1%
1-
12
#811260000000
0!
0%
b11 *
0-
02
b11 6
#811270000000
1!
1%
1-
12
15
#811280000000
0!
0%
b100 *
0-
02
b100 6
#811290000000
1!
1%
1-
12
#811300000000
0!
0%
b101 *
0-
02
b101 6
#811310000000
1!
1%
1-
12
#811320000000
0!
0%
b110 *
0-
02
b110 6
#811330000000
1!
1%
1-
12
#811340000000
0!
0%
b111 *
0-
02
b111 6
#811350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#811360000000
0!
0%
b0 *
0-
02
b0 6
#811370000000
1!
1%
1-
12
#811380000000
0!
0%
b1 *
0-
02
b1 6
#811390000000
1!
1%
1-
12
#811400000000
0!
0%
b10 *
0-
02
b10 6
#811410000000
1!
1%
1-
12
#811420000000
0!
0%
b11 *
0-
02
b11 6
#811430000000
1!
1%
1-
12
15
#811440000000
0!
0%
b100 *
0-
02
b100 6
#811450000000
1!
1%
1-
12
#811460000000
0!
0%
b101 *
0-
02
b101 6
#811470000000
1!
1%
1-
12
#811480000000
0!
0%
b110 *
0-
02
b110 6
#811490000000
1!
1%
1-
12
#811500000000
0!
0%
b111 *
0-
02
b111 6
#811510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#811520000000
0!
0%
b0 *
0-
02
b0 6
#811530000000
1!
1%
1-
12
#811540000000
0!
0%
b1 *
0-
02
b1 6
#811550000000
1!
1%
1-
12
#811560000000
0!
0%
b10 *
0-
02
b10 6
#811570000000
1!
1%
1-
12
#811580000000
0!
0%
b11 *
0-
02
b11 6
#811590000000
1!
1%
1-
12
15
#811600000000
0!
0%
b100 *
0-
02
b100 6
#811610000000
1!
1%
1-
12
#811620000000
0!
0%
b101 *
0-
02
b101 6
#811630000000
1!
1%
1-
12
#811640000000
0!
0%
b110 *
0-
02
b110 6
#811650000000
1!
1%
1-
12
#811660000000
0!
0%
b111 *
0-
02
b111 6
#811670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#811680000000
0!
0%
b0 *
0-
02
b0 6
#811690000000
1!
1%
1-
12
#811700000000
0!
0%
b1 *
0-
02
b1 6
#811710000000
1!
1%
1-
12
#811720000000
0!
0%
b10 *
0-
02
b10 6
#811730000000
1!
1%
1-
12
#811740000000
0!
0%
b11 *
0-
02
b11 6
#811750000000
1!
1%
1-
12
15
#811760000000
0!
0%
b100 *
0-
02
b100 6
#811770000000
1!
1%
1-
12
#811780000000
0!
0%
b101 *
0-
02
b101 6
#811790000000
1!
1%
1-
12
#811800000000
0!
0%
b110 *
0-
02
b110 6
#811810000000
1!
1%
1-
12
#811820000000
0!
0%
b111 *
0-
02
b111 6
#811830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#811840000000
0!
0%
b0 *
0-
02
b0 6
#811850000000
1!
1%
1-
12
#811860000000
0!
0%
b1 *
0-
02
b1 6
#811870000000
1!
1%
1-
12
#811880000000
0!
0%
b10 *
0-
02
b10 6
#811890000000
1!
1%
1-
12
#811900000000
0!
0%
b11 *
0-
02
b11 6
#811910000000
1!
1%
1-
12
15
#811920000000
0!
0%
b100 *
0-
02
b100 6
#811930000000
1!
1%
1-
12
#811940000000
0!
0%
b101 *
0-
02
b101 6
#811950000000
1!
1%
1-
12
#811960000000
0!
0%
b110 *
0-
02
b110 6
#811970000000
1!
1%
1-
12
#811980000000
0!
0%
b111 *
0-
02
b111 6
#811990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#812000000000
0!
0%
b0 *
0-
02
b0 6
#812010000000
1!
1%
1-
12
#812020000000
0!
0%
b1 *
0-
02
b1 6
#812030000000
1!
1%
1-
12
#812040000000
0!
0%
b10 *
0-
02
b10 6
#812050000000
1!
1%
1-
12
#812060000000
0!
0%
b11 *
0-
02
b11 6
#812070000000
1!
1%
1-
12
15
#812080000000
0!
0%
b100 *
0-
02
b100 6
#812090000000
1!
1%
1-
12
#812100000000
0!
0%
b101 *
0-
02
b101 6
#812110000000
1!
1%
1-
12
#812120000000
0!
0%
b110 *
0-
02
b110 6
#812130000000
1!
1%
1-
12
#812140000000
0!
0%
b111 *
0-
02
b111 6
#812150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#812160000000
0!
0%
b0 *
0-
02
b0 6
#812170000000
1!
1%
1-
12
#812180000000
0!
0%
b1 *
0-
02
b1 6
#812190000000
1!
1%
1-
12
#812200000000
0!
0%
b10 *
0-
02
b10 6
#812210000000
1!
1%
1-
12
#812220000000
0!
0%
b11 *
0-
02
b11 6
#812230000000
1!
1%
1-
12
15
#812240000000
0!
0%
b100 *
0-
02
b100 6
#812250000000
1!
1%
1-
12
#812260000000
0!
0%
b101 *
0-
02
b101 6
#812270000000
1!
1%
1-
12
#812280000000
0!
0%
b110 *
0-
02
b110 6
#812290000000
1!
1%
1-
12
#812300000000
0!
0%
b111 *
0-
02
b111 6
#812310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#812320000000
0!
0%
b0 *
0-
02
b0 6
#812330000000
1!
1%
1-
12
#812340000000
0!
0%
b1 *
0-
02
b1 6
#812350000000
1!
1%
1-
12
#812360000000
0!
0%
b10 *
0-
02
b10 6
#812370000000
1!
1%
1-
12
#812380000000
0!
0%
b11 *
0-
02
b11 6
#812390000000
1!
1%
1-
12
15
#812400000000
0!
0%
b100 *
0-
02
b100 6
#812410000000
1!
1%
1-
12
#812420000000
0!
0%
b101 *
0-
02
b101 6
#812430000000
1!
1%
1-
12
#812440000000
0!
0%
b110 *
0-
02
b110 6
#812450000000
1!
1%
1-
12
#812460000000
0!
0%
b111 *
0-
02
b111 6
#812470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#812480000000
0!
0%
b0 *
0-
02
b0 6
#812490000000
1!
1%
1-
12
#812500000000
0!
0%
b1 *
0-
02
b1 6
#812510000000
1!
1%
1-
12
#812520000000
0!
0%
b10 *
0-
02
b10 6
#812530000000
1!
1%
1-
12
#812540000000
0!
0%
b11 *
0-
02
b11 6
#812550000000
1!
1%
1-
12
15
#812560000000
0!
0%
b100 *
0-
02
b100 6
#812570000000
1!
1%
1-
12
#812580000000
0!
0%
b101 *
0-
02
b101 6
#812590000000
1!
1%
1-
12
#812600000000
0!
0%
b110 *
0-
02
b110 6
#812610000000
1!
1%
1-
12
#812620000000
0!
0%
b111 *
0-
02
b111 6
#812630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#812640000000
0!
0%
b0 *
0-
02
b0 6
#812650000000
1!
1%
1-
12
#812660000000
0!
0%
b1 *
0-
02
b1 6
#812670000000
1!
1%
1-
12
#812680000000
0!
0%
b10 *
0-
02
b10 6
#812690000000
1!
1%
1-
12
#812700000000
0!
0%
b11 *
0-
02
b11 6
#812710000000
1!
1%
1-
12
15
#812720000000
0!
0%
b100 *
0-
02
b100 6
#812730000000
1!
1%
1-
12
#812740000000
0!
0%
b101 *
0-
02
b101 6
#812750000000
1!
1%
1-
12
#812760000000
0!
0%
b110 *
0-
02
b110 6
#812770000000
1!
1%
1-
12
#812780000000
0!
0%
b111 *
0-
02
b111 6
#812790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#812800000000
0!
0%
b0 *
0-
02
b0 6
#812810000000
1!
1%
1-
12
#812820000000
0!
0%
b1 *
0-
02
b1 6
#812830000000
1!
1%
1-
12
#812840000000
0!
0%
b10 *
0-
02
b10 6
#812850000000
1!
1%
1-
12
#812860000000
0!
0%
b11 *
0-
02
b11 6
#812870000000
1!
1%
1-
12
15
#812880000000
0!
0%
b100 *
0-
02
b100 6
#812890000000
1!
1%
1-
12
#812900000000
0!
0%
b101 *
0-
02
b101 6
#812910000000
1!
1%
1-
12
#812920000000
0!
0%
b110 *
0-
02
b110 6
#812930000000
1!
1%
1-
12
#812940000000
0!
0%
b111 *
0-
02
b111 6
#812950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#812960000000
0!
0%
b0 *
0-
02
b0 6
#812970000000
1!
1%
1-
12
#812980000000
0!
0%
b1 *
0-
02
b1 6
#812990000000
1!
1%
1-
12
#813000000000
0!
0%
b10 *
0-
02
b10 6
#813010000000
1!
1%
1-
12
#813020000000
0!
0%
b11 *
0-
02
b11 6
#813030000000
1!
1%
1-
12
15
#813040000000
0!
0%
b100 *
0-
02
b100 6
#813050000000
1!
1%
1-
12
#813060000000
0!
0%
b101 *
0-
02
b101 6
#813070000000
1!
1%
1-
12
#813080000000
0!
0%
b110 *
0-
02
b110 6
#813090000000
1!
1%
1-
12
#813100000000
0!
0%
b111 *
0-
02
b111 6
#813110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#813120000000
0!
0%
b0 *
0-
02
b0 6
#813130000000
1!
1%
1-
12
#813140000000
0!
0%
b1 *
0-
02
b1 6
#813150000000
1!
1%
1-
12
#813160000000
0!
0%
b10 *
0-
02
b10 6
#813170000000
1!
1%
1-
12
#813180000000
0!
0%
b11 *
0-
02
b11 6
#813190000000
1!
1%
1-
12
15
#813200000000
0!
0%
b100 *
0-
02
b100 6
#813210000000
1!
1%
1-
12
#813220000000
0!
0%
b101 *
0-
02
b101 6
#813230000000
1!
1%
1-
12
#813240000000
0!
0%
b110 *
0-
02
b110 6
#813250000000
1!
1%
1-
12
#813260000000
0!
0%
b111 *
0-
02
b111 6
#813270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#813280000000
0!
0%
b0 *
0-
02
b0 6
#813290000000
1!
1%
1-
12
#813300000000
0!
0%
b1 *
0-
02
b1 6
#813310000000
1!
1%
1-
12
#813320000000
0!
0%
b10 *
0-
02
b10 6
#813330000000
1!
1%
1-
12
#813340000000
0!
0%
b11 *
0-
02
b11 6
#813350000000
1!
1%
1-
12
15
#813360000000
0!
0%
b100 *
0-
02
b100 6
#813370000000
1!
1%
1-
12
#813380000000
0!
0%
b101 *
0-
02
b101 6
#813390000000
1!
1%
1-
12
#813400000000
0!
0%
b110 *
0-
02
b110 6
#813410000000
1!
1%
1-
12
#813420000000
0!
0%
b111 *
0-
02
b111 6
#813430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#813440000000
0!
0%
b0 *
0-
02
b0 6
#813450000000
1!
1%
1-
12
#813460000000
0!
0%
b1 *
0-
02
b1 6
#813470000000
1!
1%
1-
12
#813480000000
0!
0%
b10 *
0-
02
b10 6
#813490000000
1!
1%
1-
12
#813500000000
0!
0%
b11 *
0-
02
b11 6
#813510000000
1!
1%
1-
12
15
#813520000000
0!
0%
b100 *
0-
02
b100 6
#813530000000
1!
1%
1-
12
#813540000000
0!
0%
b101 *
0-
02
b101 6
#813550000000
1!
1%
1-
12
#813560000000
0!
0%
b110 *
0-
02
b110 6
#813570000000
1!
1%
1-
12
#813580000000
0!
0%
b111 *
0-
02
b111 6
#813590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#813600000000
0!
0%
b0 *
0-
02
b0 6
#813610000000
1!
1%
1-
12
#813620000000
0!
0%
b1 *
0-
02
b1 6
#813630000000
1!
1%
1-
12
#813640000000
0!
0%
b10 *
0-
02
b10 6
#813650000000
1!
1%
1-
12
#813660000000
0!
0%
b11 *
0-
02
b11 6
#813670000000
1!
1%
1-
12
15
#813680000000
0!
0%
b100 *
0-
02
b100 6
#813690000000
1!
1%
1-
12
#813700000000
0!
0%
b101 *
0-
02
b101 6
#813710000000
1!
1%
1-
12
#813720000000
0!
0%
b110 *
0-
02
b110 6
#813730000000
1!
1%
1-
12
#813740000000
0!
0%
b111 *
0-
02
b111 6
#813750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#813760000000
0!
0%
b0 *
0-
02
b0 6
#813770000000
1!
1%
1-
12
#813780000000
0!
0%
b1 *
0-
02
b1 6
#813790000000
1!
1%
1-
12
#813800000000
0!
0%
b10 *
0-
02
b10 6
#813810000000
1!
1%
1-
12
#813820000000
0!
0%
b11 *
0-
02
b11 6
#813830000000
1!
1%
1-
12
15
#813840000000
0!
0%
b100 *
0-
02
b100 6
#813850000000
1!
1%
1-
12
#813860000000
0!
0%
b101 *
0-
02
b101 6
#813870000000
1!
1%
1-
12
#813880000000
0!
0%
b110 *
0-
02
b110 6
#813890000000
1!
1%
1-
12
#813900000000
0!
0%
b111 *
0-
02
b111 6
#813910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#813920000000
0!
0%
b0 *
0-
02
b0 6
#813930000000
1!
1%
1-
12
#813940000000
0!
0%
b1 *
0-
02
b1 6
#813950000000
1!
1%
1-
12
#813960000000
0!
0%
b10 *
0-
02
b10 6
#813970000000
1!
1%
1-
12
#813980000000
0!
0%
b11 *
0-
02
b11 6
#813990000000
1!
1%
1-
12
15
#814000000000
0!
0%
b100 *
0-
02
b100 6
#814010000000
1!
1%
1-
12
#814020000000
0!
0%
b101 *
0-
02
b101 6
#814030000000
1!
1%
1-
12
#814040000000
0!
0%
b110 *
0-
02
b110 6
#814050000000
1!
1%
1-
12
#814060000000
0!
0%
b111 *
0-
02
b111 6
#814070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#814080000000
0!
0%
b0 *
0-
02
b0 6
#814090000000
1!
1%
1-
12
#814100000000
0!
0%
b1 *
0-
02
b1 6
#814110000000
1!
1%
1-
12
#814120000000
0!
0%
b10 *
0-
02
b10 6
#814130000000
1!
1%
1-
12
#814140000000
0!
0%
b11 *
0-
02
b11 6
#814150000000
1!
1%
1-
12
15
#814160000000
0!
0%
b100 *
0-
02
b100 6
#814170000000
1!
1%
1-
12
#814180000000
0!
0%
b101 *
0-
02
b101 6
#814190000000
1!
1%
1-
12
#814200000000
0!
0%
b110 *
0-
02
b110 6
#814210000000
1!
1%
1-
12
#814220000000
0!
0%
b111 *
0-
02
b111 6
#814230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#814240000000
0!
0%
b0 *
0-
02
b0 6
#814250000000
1!
1%
1-
12
#814260000000
0!
0%
b1 *
0-
02
b1 6
#814270000000
1!
1%
1-
12
#814280000000
0!
0%
b10 *
0-
02
b10 6
#814290000000
1!
1%
1-
12
#814300000000
0!
0%
b11 *
0-
02
b11 6
#814310000000
1!
1%
1-
12
15
#814320000000
0!
0%
b100 *
0-
02
b100 6
#814330000000
1!
1%
1-
12
#814340000000
0!
0%
b101 *
0-
02
b101 6
#814350000000
1!
1%
1-
12
#814360000000
0!
0%
b110 *
0-
02
b110 6
#814370000000
1!
1%
1-
12
#814380000000
0!
0%
b111 *
0-
02
b111 6
#814390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#814400000000
0!
0%
b0 *
0-
02
b0 6
#814410000000
1!
1%
1-
12
#814420000000
0!
0%
b1 *
0-
02
b1 6
#814430000000
1!
1%
1-
12
#814440000000
0!
0%
b10 *
0-
02
b10 6
#814450000000
1!
1%
1-
12
#814460000000
0!
0%
b11 *
0-
02
b11 6
#814470000000
1!
1%
1-
12
15
#814480000000
0!
0%
b100 *
0-
02
b100 6
#814490000000
1!
1%
1-
12
#814500000000
0!
0%
b101 *
0-
02
b101 6
#814510000000
1!
1%
1-
12
#814520000000
0!
0%
b110 *
0-
02
b110 6
#814530000000
1!
1%
1-
12
#814540000000
0!
0%
b111 *
0-
02
b111 6
#814550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#814560000000
0!
0%
b0 *
0-
02
b0 6
#814570000000
1!
1%
1-
12
#814580000000
0!
0%
b1 *
0-
02
b1 6
#814590000000
1!
1%
1-
12
#814600000000
0!
0%
b10 *
0-
02
b10 6
#814610000000
1!
1%
1-
12
#814620000000
0!
0%
b11 *
0-
02
b11 6
#814630000000
1!
1%
1-
12
15
#814640000000
0!
0%
b100 *
0-
02
b100 6
#814650000000
1!
1%
1-
12
#814660000000
0!
0%
b101 *
0-
02
b101 6
#814670000000
1!
1%
1-
12
#814680000000
0!
0%
b110 *
0-
02
b110 6
#814690000000
1!
1%
1-
12
#814700000000
0!
0%
b111 *
0-
02
b111 6
#814710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#814720000000
0!
0%
b0 *
0-
02
b0 6
#814730000000
1!
1%
1-
12
#814740000000
0!
0%
b1 *
0-
02
b1 6
#814750000000
1!
1%
1-
12
#814760000000
0!
0%
b10 *
0-
02
b10 6
#814770000000
1!
1%
1-
12
#814780000000
0!
0%
b11 *
0-
02
b11 6
#814790000000
1!
1%
1-
12
15
#814800000000
0!
0%
b100 *
0-
02
b100 6
#814810000000
1!
1%
1-
12
#814820000000
0!
0%
b101 *
0-
02
b101 6
#814830000000
1!
1%
1-
12
#814840000000
0!
0%
b110 *
0-
02
b110 6
#814850000000
1!
1%
1-
12
#814860000000
0!
0%
b111 *
0-
02
b111 6
#814870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#814880000000
0!
0%
b0 *
0-
02
b0 6
#814890000000
1!
1%
1-
12
#814900000000
0!
0%
b1 *
0-
02
b1 6
#814910000000
1!
1%
1-
12
#814920000000
0!
0%
b10 *
0-
02
b10 6
#814930000000
1!
1%
1-
12
#814940000000
0!
0%
b11 *
0-
02
b11 6
#814950000000
1!
1%
1-
12
15
#814960000000
0!
0%
b100 *
0-
02
b100 6
#814970000000
1!
1%
1-
12
#814980000000
0!
0%
b101 *
0-
02
b101 6
#814990000000
1!
1%
1-
12
#815000000000
0!
0%
b110 *
0-
02
b110 6
#815010000000
1!
1%
1-
12
#815020000000
0!
0%
b111 *
0-
02
b111 6
#815030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#815040000000
0!
0%
b0 *
0-
02
b0 6
#815050000000
1!
1%
1-
12
#815060000000
0!
0%
b1 *
0-
02
b1 6
#815070000000
1!
1%
1-
12
#815080000000
0!
0%
b10 *
0-
02
b10 6
#815090000000
1!
1%
1-
12
#815100000000
0!
0%
b11 *
0-
02
b11 6
#815110000000
1!
1%
1-
12
15
#815120000000
0!
0%
b100 *
0-
02
b100 6
#815130000000
1!
1%
1-
12
#815140000000
0!
0%
b101 *
0-
02
b101 6
#815150000000
1!
1%
1-
12
#815160000000
0!
0%
b110 *
0-
02
b110 6
#815170000000
1!
1%
1-
12
#815180000000
0!
0%
b111 *
0-
02
b111 6
#815190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#815200000000
0!
0%
b0 *
0-
02
b0 6
#815210000000
1!
1%
1-
12
#815220000000
0!
0%
b1 *
0-
02
b1 6
#815230000000
1!
1%
1-
12
#815240000000
0!
0%
b10 *
0-
02
b10 6
#815250000000
1!
1%
1-
12
#815260000000
0!
0%
b11 *
0-
02
b11 6
#815270000000
1!
1%
1-
12
15
#815280000000
0!
0%
b100 *
0-
02
b100 6
#815290000000
1!
1%
1-
12
#815300000000
0!
0%
b101 *
0-
02
b101 6
#815310000000
1!
1%
1-
12
#815320000000
0!
0%
b110 *
0-
02
b110 6
#815330000000
1!
1%
1-
12
#815340000000
0!
0%
b111 *
0-
02
b111 6
#815350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#815360000000
0!
0%
b0 *
0-
02
b0 6
#815370000000
1!
1%
1-
12
#815380000000
0!
0%
b1 *
0-
02
b1 6
#815390000000
1!
1%
1-
12
#815400000000
0!
0%
b10 *
0-
02
b10 6
#815410000000
1!
1%
1-
12
#815420000000
0!
0%
b11 *
0-
02
b11 6
#815430000000
1!
1%
1-
12
15
#815440000000
0!
0%
b100 *
0-
02
b100 6
#815450000000
1!
1%
1-
12
#815460000000
0!
0%
b101 *
0-
02
b101 6
#815470000000
1!
1%
1-
12
#815480000000
0!
0%
b110 *
0-
02
b110 6
#815490000000
1!
1%
1-
12
#815500000000
0!
0%
b111 *
0-
02
b111 6
#815510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#815520000000
0!
0%
b0 *
0-
02
b0 6
#815530000000
1!
1%
1-
12
#815540000000
0!
0%
b1 *
0-
02
b1 6
#815550000000
1!
1%
1-
12
#815560000000
0!
0%
b10 *
0-
02
b10 6
#815570000000
1!
1%
1-
12
#815580000000
0!
0%
b11 *
0-
02
b11 6
#815590000000
1!
1%
1-
12
15
#815600000000
0!
0%
b100 *
0-
02
b100 6
#815610000000
1!
1%
1-
12
#815620000000
0!
0%
b101 *
0-
02
b101 6
#815630000000
1!
1%
1-
12
#815640000000
0!
0%
b110 *
0-
02
b110 6
#815650000000
1!
1%
1-
12
#815660000000
0!
0%
b111 *
0-
02
b111 6
#815670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#815680000000
0!
0%
b0 *
0-
02
b0 6
#815690000000
1!
1%
1-
12
#815700000000
0!
0%
b1 *
0-
02
b1 6
#815710000000
1!
1%
1-
12
#815720000000
0!
0%
b10 *
0-
02
b10 6
#815730000000
1!
1%
1-
12
#815740000000
0!
0%
b11 *
0-
02
b11 6
#815750000000
1!
1%
1-
12
15
#815760000000
0!
0%
b100 *
0-
02
b100 6
#815770000000
1!
1%
1-
12
#815780000000
0!
0%
b101 *
0-
02
b101 6
#815790000000
1!
1%
1-
12
#815800000000
0!
0%
b110 *
0-
02
b110 6
#815810000000
1!
1%
1-
12
#815820000000
0!
0%
b111 *
0-
02
b111 6
#815830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#815840000000
0!
0%
b0 *
0-
02
b0 6
#815850000000
1!
1%
1-
12
#815860000000
0!
0%
b1 *
0-
02
b1 6
#815870000000
1!
1%
1-
12
#815880000000
0!
0%
b10 *
0-
02
b10 6
#815890000000
1!
1%
1-
12
#815900000000
0!
0%
b11 *
0-
02
b11 6
#815910000000
1!
1%
1-
12
15
#815920000000
0!
0%
b100 *
0-
02
b100 6
#815930000000
1!
1%
1-
12
#815940000000
0!
0%
b101 *
0-
02
b101 6
#815950000000
1!
1%
1-
12
#815960000000
0!
0%
b110 *
0-
02
b110 6
#815970000000
1!
1%
1-
12
#815980000000
0!
0%
b111 *
0-
02
b111 6
#815990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#816000000000
0!
0%
b0 *
0-
02
b0 6
#816010000000
1!
1%
1-
12
#816020000000
0!
0%
b1 *
0-
02
b1 6
#816030000000
1!
1%
1-
12
#816040000000
0!
0%
b10 *
0-
02
b10 6
#816050000000
1!
1%
1-
12
#816060000000
0!
0%
b11 *
0-
02
b11 6
#816070000000
1!
1%
1-
12
15
#816080000000
0!
0%
b100 *
0-
02
b100 6
#816090000000
1!
1%
1-
12
#816100000000
0!
0%
b101 *
0-
02
b101 6
#816110000000
1!
1%
1-
12
#816120000000
0!
0%
b110 *
0-
02
b110 6
#816130000000
1!
1%
1-
12
#816140000000
0!
0%
b111 *
0-
02
b111 6
#816150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#816160000000
0!
0%
b0 *
0-
02
b0 6
#816170000000
1!
1%
1-
12
#816180000000
0!
0%
b1 *
0-
02
b1 6
#816190000000
1!
1%
1-
12
#816200000000
0!
0%
b10 *
0-
02
b10 6
#816210000000
1!
1%
1-
12
#816220000000
0!
0%
b11 *
0-
02
b11 6
#816230000000
1!
1%
1-
12
15
#816240000000
0!
0%
b100 *
0-
02
b100 6
#816250000000
1!
1%
1-
12
#816260000000
0!
0%
b101 *
0-
02
b101 6
#816270000000
1!
1%
1-
12
#816280000000
0!
0%
b110 *
0-
02
b110 6
#816290000000
1!
1%
1-
12
#816300000000
0!
0%
b111 *
0-
02
b111 6
#816310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#816320000000
0!
0%
b0 *
0-
02
b0 6
#816330000000
1!
1%
1-
12
#816340000000
0!
0%
b1 *
0-
02
b1 6
#816350000000
1!
1%
1-
12
#816360000000
0!
0%
b10 *
0-
02
b10 6
#816370000000
1!
1%
1-
12
#816380000000
0!
0%
b11 *
0-
02
b11 6
#816390000000
1!
1%
1-
12
15
#816400000000
0!
0%
b100 *
0-
02
b100 6
#816410000000
1!
1%
1-
12
#816420000000
0!
0%
b101 *
0-
02
b101 6
#816430000000
1!
1%
1-
12
#816440000000
0!
0%
b110 *
0-
02
b110 6
#816450000000
1!
1%
1-
12
#816460000000
0!
0%
b111 *
0-
02
b111 6
#816470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#816480000000
0!
0%
b0 *
0-
02
b0 6
#816490000000
1!
1%
1-
12
#816500000000
0!
0%
b1 *
0-
02
b1 6
#816510000000
1!
1%
1-
12
#816520000000
0!
0%
b10 *
0-
02
b10 6
#816530000000
1!
1%
1-
12
#816540000000
0!
0%
b11 *
0-
02
b11 6
#816550000000
1!
1%
1-
12
15
#816560000000
0!
0%
b100 *
0-
02
b100 6
#816570000000
1!
1%
1-
12
#816580000000
0!
0%
b101 *
0-
02
b101 6
#816590000000
1!
1%
1-
12
#816600000000
0!
0%
b110 *
0-
02
b110 6
#816610000000
1!
1%
1-
12
#816620000000
0!
0%
b111 *
0-
02
b111 6
#816630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#816640000000
0!
0%
b0 *
0-
02
b0 6
#816650000000
1!
1%
1-
12
#816660000000
0!
0%
b1 *
0-
02
b1 6
#816670000000
1!
1%
1-
12
#816680000000
0!
0%
b10 *
0-
02
b10 6
#816690000000
1!
1%
1-
12
#816700000000
0!
0%
b11 *
0-
02
b11 6
#816710000000
1!
1%
1-
12
15
#816720000000
0!
0%
b100 *
0-
02
b100 6
#816730000000
1!
1%
1-
12
#816740000000
0!
0%
b101 *
0-
02
b101 6
#816750000000
1!
1%
1-
12
#816760000000
0!
0%
b110 *
0-
02
b110 6
#816770000000
1!
1%
1-
12
#816780000000
0!
0%
b111 *
0-
02
b111 6
#816790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#816800000000
0!
0%
b0 *
0-
02
b0 6
#816810000000
1!
1%
1-
12
#816820000000
0!
0%
b1 *
0-
02
b1 6
#816830000000
1!
1%
1-
12
#816840000000
0!
0%
b10 *
0-
02
b10 6
#816850000000
1!
1%
1-
12
#816860000000
0!
0%
b11 *
0-
02
b11 6
#816870000000
1!
1%
1-
12
15
#816880000000
0!
0%
b100 *
0-
02
b100 6
#816890000000
1!
1%
1-
12
#816900000000
0!
0%
b101 *
0-
02
b101 6
#816910000000
1!
1%
1-
12
#816920000000
0!
0%
b110 *
0-
02
b110 6
#816930000000
1!
1%
1-
12
#816940000000
0!
0%
b111 *
0-
02
b111 6
#816950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#816960000000
0!
0%
b0 *
0-
02
b0 6
#816970000000
1!
1%
1-
12
#816980000000
0!
0%
b1 *
0-
02
b1 6
#816990000000
1!
1%
1-
12
#817000000000
0!
0%
b10 *
0-
02
b10 6
#817010000000
1!
1%
1-
12
#817020000000
0!
0%
b11 *
0-
02
b11 6
#817030000000
1!
1%
1-
12
15
#817040000000
0!
0%
b100 *
0-
02
b100 6
#817050000000
1!
1%
1-
12
#817060000000
0!
0%
b101 *
0-
02
b101 6
#817070000000
1!
1%
1-
12
#817080000000
0!
0%
b110 *
0-
02
b110 6
#817090000000
1!
1%
1-
12
#817100000000
0!
0%
b111 *
0-
02
b111 6
#817110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#817120000000
0!
0%
b0 *
0-
02
b0 6
#817130000000
1!
1%
1-
12
#817140000000
0!
0%
b1 *
0-
02
b1 6
#817150000000
1!
1%
1-
12
#817160000000
0!
0%
b10 *
0-
02
b10 6
#817170000000
1!
1%
1-
12
#817180000000
0!
0%
b11 *
0-
02
b11 6
#817190000000
1!
1%
1-
12
15
#817200000000
0!
0%
b100 *
0-
02
b100 6
#817210000000
1!
1%
1-
12
#817220000000
0!
0%
b101 *
0-
02
b101 6
#817230000000
1!
1%
1-
12
#817240000000
0!
0%
b110 *
0-
02
b110 6
#817250000000
1!
1%
1-
12
#817260000000
0!
0%
b111 *
0-
02
b111 6
#817270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#817280000000
0!
0%
b0 *
0-
02
b0 6
#817290000000
1!
1%
1-
12
#817300000000
0!
0%
b1 *
0-
02
b1 6
#817310000000
1!
1%
1-
12
#817320000000
0!
0%
b10 *
0-
02
b10 6
#817330000000
1!
1%
1-
12
#817340000000
0!
0%
b11 *
0-
02
b11 6
#817350000000
1!
1%
1-
12
15
#817360000000
0!
0%
b100 *
0-
02
b100 6
#817370000000
1!
1%
1-
12
#817380000000
0!
0%
b101 *
0-
02
b101 6
#817390000000
1!
1%
1-
12
#817400000000
0!
0%
b110 *
0-
02
b110 6
#817410000000
1!
1%
1-
12
#817420000000
0!
0%
b111 *
0-
02
b111 6
#817430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#817440000000
0!
0%
b0 *
0-
02
b0 6
#817450000000
1!
1%
1-
12
#817460000000
0!
0%
b1 *
0-
02
b1 6
#817470000000
1!
1%
1-
12
#817480000000
0!
0%
b10 *
0-
02
b10 6
#817490000000
1!
1%
1-
12
#817500000000
0!
0%
b11 *
0-
02
b11 6
#817510000000
1!
1%
1-
12
15
#817520000000
0!
0%
b100 *
0-
02
b100 6
#817530000000
1!
1%
1-
12
#817540000000
0!
0%
b101 *
0-
02
b101 6
#817550000000
1!
1%
1-
12
#817560000000
0!
0%
b110 *
0-
02
b110 6
#817570000000
1!
1%
1-
12
#817580000000
0!
0%
b111 *
0-
02
b111 6
#817590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#817600000000
0!
0%
b0 *
0-
02
b0 6
#817610000000
1!
1%
1-
12
#817620000000
0!
0%
b1 *
0-
02
b1 6
#817630000000
1!
1%
1-
12
#817640000000
0!
0%
b10 *
0-
02
b10 6
#817650000000
1!
1%
1-
12
#817660000000
0!
0%
b11 *
0-
02
b11 6
#817670000000
1!
1%
1-
12
15
#817680000000
0!
0%
b100 *
0-
02
b100 6
#817690000000
1!
1%
1-
12
#817700000000
0!
0%
b101 *
0-
02
b101 6
#817710000000
1!
1%
1-
12
#817720000000
0!
0%
b110 *
0-
02
b110 6
#817730000000
1!
1%
1-
12
#817740000000
0!
0%
b111 *
0-
02
b111 6
#817750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#817760000000
0!
0%
b0 *
0-
02
b0 6
#817770000000
1!
1%
1-
12
#817780000000
0!
0%
b1 *
0-
02
b1 6
#817790000000
1!
1%
1-
12
#817800000000
0!
0%
b10 *
0-
02
b10 6
#817810000000
1!
1%
1-
12
#817820000000
0!
0%
b11 *
0-
02
b11 6
#817830000000
1!
1%
1-
12
15
#817840000000
0!
0%
b100 *
0-
02
b100 6
#817850000000
1!
1%
1-
12
#817860000000
0!
0%
b101 *
0-
02
b101 6
#817870000000
1!
1%
1-
12
#817880000000
0!
0%
b110 *
0-
02
b110 6
#817890000000
1!
1%
1-
12
#817900000000
0!
0%
b111 *
0-
02
b111 6
#817910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#817920000000
0!
0%
b0 *
0-
02
b0 6
#817930000000
1!
1%
1-
12
#817940000000
0!
0%
b1 *
0-
02
b1 6
#817950000000
1!
1%
1-
12
#817960000000
0!
0%
b10 *
0-
02
b10 6
#817970000000
1!
1%
1-
12
#817980000000
0!
0%
b11 *
0-
02
b11 6
#817990000000
1!
1%
1-
12
15
#818000000000
0!
0%
b100 *
0-
02
b100 6
#818010000000
1!
1%
1-
12
#818020000000
0!
0%
b101 *
0-
02
b101 6
#818030000000
1!
1%
1-
12
#818040000000
0!
0%
b110 *
0-
02
b110 6
#818050000000
1!
1%
1-
12
#818060000000
0!
0%
b111 *
0-
02
b111 6
#818070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#818080000000
0!
0%
b0 *
0-
02
b0 6
#818090000000
1!
1%
1-
12
#818100000000
0!
0%
b1 *
0-
02
b1 6
#818110000000
1!
1%
1-
12
#818120000000
0!
0%
b10 *
0-
02
b10 6
#818130000000
1!
1%
1-
12
#818140000000
0!
0%
b11 *
0-
02
b11 6
#818150000000
1!
1%
1-
12
15
#818160000000
0!
0%
b100 *
0-
02
b100 6
#818170000000
1!
1%
1-
12
#818180000000
0!
0%
b101 *
0-
02
b101 6
#818190000000
1!
1%
1-
12
#818200000000
0!
0%
b110 *
0-
02
b110 6
#818210000000
1!
1%
1-
12
#818220000000
0!
0%
b111 *
0-
02
b111 6
#818230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#818240000000
0!
0%
b0 *
0-
02
b0 6
#818250000000
1!
1%
1-
12
#818260000000
0!
0%
b1 *
0-
02
b1 6
#818270000000
1!
1%
1-
12
#818280000000
0!
0%
b10 *
0-
02
b10 6
#818290000000
1!
1%
1-
12
#818300000000
0!
0%
b11 *
0-
02
b11 6
#818310000000
1!
1%
1-
12
15
#818320000000
0!
0%
b100 *
0-
02
b100 6
#818330000000
1!
1%
1-
12
#818340000000
0!
0%
b101 *
0-
02
b101 6
#818350000000
1!
1%
1-
12
#818360000000
0!
0%
b110 *
0-
02
b110 6
#818370000000
1!
1%
1-
12
#818380000000
0!
0%
b111 *
0-
02
b111 6
#818390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#818400000000
0!
0%
b0 *
0-
02
b0 6
#818410000000
1!
1%
1-
12
#818420000000
0!
0%
b1 *
0-
02
b1 6
#818430000000
1!
1%
1-
12
#818440000000
0!
0%
b10 *
0-
02
b10 6
#818450000000
1!
1%
1-
12
#818460000000
0!
0%
b11 *
0-
02
b11 6
#818470000000
1!
1%
1-
12
15
#818480000000
0!
0%
b100 *
0-
02
b100 6
#818490000000
1!
1%
1-
12
#818500000000
0!
0%
b101 *
0-
02
b101 6
#818510000000
1!
1%
1-
12
#818520000000
0!
0%
b110 *
0-
02
b110 6
#818530000000
1!
1%
1-
12
#818540000000
0!
0%
b111 *
0-
02
b111 6
#818550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#818560000000
0!
0%
b0 *
0-
02
b0 6
#818570000000
1!
1%
1-
12
#818580000000
0!
0%
b1 *
0-
02
b1 6
#818590000000
1!
1%
1-
12
#818600000000
0!
0%
b10 *
0-
02
b10 6
#818610000000
1!
1%
1-
12
#818620000000
0!
0%
b11 *
0-
02
b11 6
#818630000000
1!
1%
1-
12
15
#818640000000
0!
0%
b100 *
0-
02
b100 6
#818650000000
1!
1%
1-
12
#818660000000
0!
0%
b101 *
0-
02
b101 6
#818670000000
1!
1%
1-
12
#818680000000
0!
0%
b110 *
0-
02
b110 6
#818690000000
1!
1%
1-
12
#818700000000
0!
0%
b111 *
0-
02
b111 6
#818710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#818720000000
0!
0%
b0 *
0-
02
b0 6
#818730000000
1!
1%
1-
12
#818740000000
0!
0%
b1 *
0-
02
b1 6
#818750000000
1!
1%
1-
12
#818760000000
0!
0%
b10 *
0-
02
b10 6
#818770000000
1!
1%
1-
12
#818780000000
0!
0%
b11 *
0-
02
b11 6
#818790000000
1!
1%
1-
12
15
#818800000000
0!
0%
b100 *
0-
02
b100 6
#818810000000
1!
1%
1-
12
#818820000000
0!
0%
b101 *
0-
02
b101 6
#818830000000
1!
1%
1-
12
#818840000000
0!
0%
b110 *
0-
02
b110 6
#818850000000
1!
1%
1-
12
#818860000000
0!
0%
b111 *
0-
02
b111 6
#818870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#818880000000
0!
0%
b0 *
0-
02
b0 6
#818890000000
1!
1%
1-
12
#818900000000
0!
0%
b1 *
0-
02
b1 6
#818910000000
1!
1%
1-
12
#818920000000
0!
0%
b10 *
0-
02
b10 6
#818930000000
1!
1%
1-
12
#818940000000
0!
0%
b11 *
0-
02
b11 6
#818950000000
1!
1%
1-
12
15
#818960000000
0!
0%
b100 *
0-
02
b100 6
#818970000000
1!
1%
1-
12
#818980000000
0!
0%
b101 *
0-
02
b101 6
#818990000000
1!
1%
1-
12
#819000000000
0!
0%
b110 *
0-
02
b110 6
#819010000000
1!
1%
1-
12
#819020000000
0!
0%
b111 *
0-
02
b111 6
#819030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#819040000000
0!
0%
b0 *
0-
02
b0 6
#819050000000
1!
1%
1-
12
#819060000000
0!
0%
b1 *
0-
02
b1 6
#819070000000
1!
1%
1-
12
#819080000000
0!
0%
b10 *
0-
02
b10 6
#819090000000
1!
1%
1-
12
#819100000000
0!
0%
b11 *
0-
02
b11 6
#819110000000
1!
1%
1-
12
15
#819120000000
0!
0%
b100 *
0-
02
b100 6
#819130000000
1!
1%
1-
12
#819140000000
0!
0%
b101 *
0-
02
b101 6
#819150000000
1!
1%
1-
12
#819160000000
0!
0%
b110 *
0-
02
b110 6
#819170000000
1!
1%
1-
12
#819180000000
0!
0%
b111 *
0-
02
b111 6
#819190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#819200000000
0!
0%
b0 *
0-
02
b0 6
#819210000000
1!
1%
1-
12
#819220000000
0!
0%
b1 *
0-
02
b1 6
#819230000000
1!
1%
1-
12
#819240000000
0!
0%
b10 *
0-
02
b10 6
#819250000000
1!
1%
1-
12
#819260000000
0!
0%
b11 *
0-
02
b11 6
#819270000000
1!
1%
1-
12
15
#819280000000
0!
0%
b100 *
0-
02
b100 6
#819290000000
1!
1%
1-
12
#819300000000
0!
0%
b101 *
0-
02
b101 6
#819310000000
1!
1%
1-
12
#819320000000
0!
0%
b110 *
0-
02
b110 6
#819330000000
1!
1%
1-
12
#819340000000
0!
0%
b111 *
0-
02
b111 6
#819350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#819360000000
0!
0%
b0 *
0-
02
b0 6
#819370000000
1!
1%
1-
12
#819380000000
0!
0%
b1 *
0-
02
b1 6
#819390000000
1!
1%
1-
12
#819400000000
0!
0%
b10 *
0-
02
b10 6
#819410000000
1!
1%
1-
12
#819420000000
0!
0%
b11 *
0-
02
b11 6
#819430000000
1!
1%
1-
12
15
#819440000000
0!
0%
b100 *
0-
02
b100 6
#819450000000
1!
1%
1-
12
#819460000000
0!
0%
b101 *
0-
02
b101 6
#819470000000
1!
1%
1-
12
#819480000000
0!
0%
b110 *
0-
02
b110 6
#819490000000
1!
1%
1-
12
#819500000000
0!
0%
b111 *
0-
02
b111 6
#819510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#819520000000
0!
0%
b0 *
0-
02
b0 6
#819530000000
1!
1%
1-
12
#819540000000
0!
0%
b1 *
0-
02
b1 6
#819550000000
1!
1%
1-
12
#819560000000
0!
0%
b10 *
0-
02
b10 6
#819570000000
1!
1%
1-
12
#819580000000
0!
0%
b11 *
0-
02
b11 6
#819590000000
1!
1%
1-
12
15
#819600000000
0!
0%
b100 *
0-
02
b100 6
#819610000000
1!
1%
1-
12
#819620000000
0!
0%
b101 *
0-
02
b101 6
#819630000000
1!
1%
1-
12
#819640000000
0!
0%
b110 *
0-
02
b110 6
#819650000000
1!
1%
1-
12
#819660000000
0!
0%
b111 *
0-
02
b111 6
#819670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#819680000000
0!
0%
b0 *
0-
02
b0 6
#819690000000
1!
1%
1-
12
#819700000000
0!
0%
b1 *
0-
02
b1 6
#819710000000
1!
1%
1-
12
#819720000000
0!
0%
b10 *
0-
02
b10 6
#819730000000
1!
1%
1-
12
#819740000000
0!
0%
b11 *
0-
02
b11 6
#819750000000
1!
1%
1-
12
15
#819760000000
0!
0%
b100 *
0-
02
b100 6
#819770000000
1!
1%
1-
12
#819780000000
0!
0%
b101 *
0-
02
b101 6
#819790000000
1!
1%
1-
12
#819800000000
0!
0%
b110 *
0-
02
b110 6
#819810000000
1!
1%
1-
12
#819820000000
0!
0%
b111 *
0-
02
b111 6
#819830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#819840000000
0!
0%
b0 *
0-
02
b0 6
#819850000000
1!
1%
1-
12
#819860000000
0!
0%
b1 *
0-
02
b1 6
#819870000000
1!
1%
1-
12
#819880000000
0!
0%
b10 *
0-
02
b10 6
#819890000000
1!
1%
1-
12
#819900000000
0!
0%
b11 *
0-
02
b11 6
#819910000000
1!
1%
1-
12
15
#819920000000
0!
0%
b100 *
0-
02
b100 6
#819930000000
1!
1%
1-
12
#819940000000
0!
0%
b101 *
0-
02
b101 6
#819950000000
1!
1%
1-
12
#819960000000
0!
0%
b110 *
0-
02
b110 6
#819970000000
1!
1%
1-
12
#819980000000
0!
0%
b111 *
0-
02
b111 6
#819990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#820000000000
0!
0%
b0 *
0-
02
b0 6
#820010000000
1!
1%
1-
12
#820020000000
0!
0%
b1 *
0-
02
b1 6
#820030000000
1!
1%
1-
12
#820040000000
0!
0%
b10 *
0-
02
b10 6
#820050000000
1!
1%
1-
12
#820060000000
0!
0%
b11 *
0-
02
b11 6
#820070000000
1!
1%
1-
12
15
#820080000000
0!
0%
b100 *
0-
02
b100 6
#820090000000
1!
1%
1-
12
#820100000000
0!
0%
b101 *
0-
02
b101 6
#820110000000
1!
1%
1-
12
#820120000000
0!
0%
b110 *
0-
02
b110 6
#820130000000
1!
1%
1-
12
#820140000000
0!
0%
b111 *
0-
02
b111 6
#820150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#820160000000
0!
0%
b0 *
0-
02
b0 6
#820170000000
1!
1%
1-
12
#820180000000
0!
0%
b1 *
0-
02
b1 6
#820190000000
1!
1%
1-
12
#820200000000
0!
0%
b10 *
0-
02
b10 6
#820210000000
1!
1%
1-
12
#820220000000
0!
0%
b11 *
0-
02
b11 6
#820230000000
1!
1%
1-
12
15
#820240000000
0!
0%
b100 *
0-
02
b100 6
#820250000000
1!
1%
1-
12
#820260000000
0!
0%
b101 *
0-
02
b101 6
#820270000000
1!
1%
1-
12
#820280000000
0!
0%
b110 *
0-
02
b110 6
#820290000000
1!
1%
1-
12
#820300000000
0!
0%
b111 *
0-
02
b111 6
#820310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#820320000000
0!
0%
b0 *
0-
02
b0 6
#820330000000
1!
1%
1-
12
#820340000000
0!
0%
b1 *
0-
02
b1 6
#820350000000
1!
1%
1-
12
#820360000000
0!
0%
b10 *
0-
02
b10 6
#820370000000
1!
1%
1-
12
#820380000000
0!
0%
b11 *
0-
02
b11 6
#820390000000
1!
1%
1-
12
15
#820400000000
0!
0%
b100 *
0-
02
b100 6
#820410000000
1!
1%
1-
12
#820420000000
0!
0%
b101 *
0-
02
b101 6
#820430000000
1!
1%
1-
12
#820440000000
0!
0%
b110 *
0-
02
b110 6
#820450000000
1!
1%
1-
12
#820460000000
0!
0%
b111 *
0-
02
b111 6
#820470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#820480000000
0!
0%
b0 *
0-
02
b0 6
#820490000000
1!
1%
1-
12
#820500000000
0!
0%
b1 *
0-
02
b1 6
#820510000000
1!
1%
1-
12
#820520000000
0!
0%
b10 *
0-
02
b10 6
#820530000000
1!
1%
1-
12
#820540000000
0!
0%
b11 *
0-
02
b11 6
#820550000000
1!
1%
1-
12
15
#820560000000
0!
0%
b100 *
0-
02
b100 6
#820570000000
1!
1%
1-
12
#820580000000
0!
0%
b101 *
0-
02
b101 6
#820590000000
1!
1%
1-
12
#820600000000
0!
0%
b110 *
0-
02
b110 6
#820610000000
1!
1%
1-
12
#820620000000
0!
0%
b111 *
0-
02
b111 6
#820630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#820640000000
0!
0%
b0 *
0-
02
b0 6
#820650000000
1!
1%
1-
12
#820660000000
0!
0%
b1 *
0-
02
b1 6
#820670000000
1!
1%
1-
12
#820680000000
0!
0%
b10 *
0-
02
b10 6
#820690000000
1!
1%
1-
12
#820700000000
0!
0%
b11 *
0-
02
b11 6
#820710000000
1!
1%
1-
12
15
#820720000000
0!
0%
b100 *
0-
02
b100 6
#820730000000
1!
1%
1-
12
#820740000000
0!
0%
b101 *
0-
02
b101 6
#820750000000
1!
1%
1-
12
#820760000000
0!
0%
b110 *
0-
02
b110 6
#820770000000
1!
1%
1-
12
#820780000000
0!
0%
b111 *
0-
02
b111 6
#820790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#820800000000
0!
0%
b0 *
0-
02
b0 6
#820810000000
1!
1%
1-
12
#820820000000
0!
0%
b1 *
0-
02
b1 6
#820830000000
1!
1%
1-
12
#820840000000
0!
0%
b10 *
0-
02
b10 6
#820850000000
1!
1%
1-
12
#820860000000
0!
0%
b11 *
0-
02
b11 6
#820870000000
1!
1%
1-
12
15
#820880000000
0!
0%
b100 *
0-
02
b100 6
#820890000000
1!
1%
1-
12
#820900000000
0!
0%
b101 *
0-
02
b101 6
#820910000000
1!
1%
1-
12
#820920000000
0!
0%
b110 *
0-
02
b110 6
#820930000000
1!
1%
1-
12
#820940000000
0!
0%
b111 *
0-
02
b111 6
#820950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#820960000000
0!
0%
b0 *
0-
02
b0 6
#820970000000
1!
1%
1-
12
#820980000000
0!
0%
b1 *
0-
02
b1 6
#820990000000
1!
1%
1-
12
#821000000000
0!
0%
b10 *
0-
02
b10 6
#821010000000
1!
1%
1-
12
#821020000000
0!
0%
b11 *
0-
02
b11 6
#821030000000
1!
1%
1-
12
15
#821040000000
0!
0%
b100 *
0-
02
b100 6
#821050000000
1!
1%
1-
12
#821060000000
0!
0%
b101 *
0-
02
b101 6
#821070000000
1!
1%
1-
12
#821080000000
0!
0%
b110 *
0-
02
b110 6
#821090000000
1!
1%
1-
12
#821100000000
0!
0%
b111 *
0-
02
b111 6
#821110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#821120000000
0!
0%
b0 *
0-
02
b0 6
#821130000000
1!
1%
1-
12
#821140000000
0!
0%
b1 *
0-
02
b1 6
#821150000000
1!
1%
1-
12
#821160000000
0!
0%
b10 *
0-
02
b10 6
#821170000000
1!
1%
1-
12
#821180000000
0!
0%
b11 *
0-
02
b11 6
#821190000000
1!
1%
1-
12
15
#821200000000
0!
0%
b100 *
0-
02
b100 6
#821210000000
1!
1%
1-
12
#821220000000
0!
0%
b101 *
0-
02
b101 6
#821230000000
1!
1%
1-
12
#821240000000
0!
0%
b110 *
0-
02
b110 6
#821250000000
1!
1%
1-
12
#821260000000
0!
0%
b111 *
0-
02
b111 6
#821270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#821280000000
0!
0%
b0 *
0-
02
b0 6
#821290000000
1!
1%
1-
12
#821300000000
0!
0%
b1 *
0-
02
b1 6
#821310000000
1!
1%
1-
12
#821320000000
0!
0%
b10 *
0-
02
b10 6
#821330000000
1!
1%
1-
12
#821340000000
0!
0%
b11 *
0-
02
b11 6
#821350000000
1!
1%
1-
12
15
#821360000000
0!
0%
b100 *
0-
02
b100 6
#821370000000
1!
1%
1-
12
#821380000000
0!
0%
b101 *
0-
02
b101 6
#821390000000
1!
1%
1-
12
#821400000000
0!
0%
b110 *
0-
02
b110 6
#821410000000
1!
1%
1-
12
#821420000000
0!
0%
b111 *
0-
02
b111 6
#821430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#821440000000
0!
0%
b0 *
0-
02
b0 6
#821450000000
1!
1%
1-
12
#821460000000
0!
0%
b1 *
0-
02
b1 6
#821470000000
1!
1%
1-
12
#821480000000
0!
0%
b10 *
0-
02
b10 6
#821490000000
1!
1%
1-
12
#821500000000
0!
0%
b11 *
0-
02
b11 6
#821510000000
1!
1%
1-
12
15
#821520000000
0!
0%
b100 *
0-
02
b100 6
#821530000000
1!
1%
1-
12
#821540000000
0!
0%
b101 *
0-
02
b101 6
#821550000000
1!
1%
1-
12
#821560000000
0!
0%
b110 *
0-
02
b110 6
#821570000000
1!
1%
1-
12
#821580000000
0!
0%
b111 *
0-
02
b111 6
#821590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#821600000000
0!
0%
b0 *
0-
02
b0 6
#821610000000
1!
1%
1-
12
#821620000000
0!
0%
b1 *
0-
02
b1 6
#821630000000
1!
1%
1-
12
#821640000000
0!
0%
b10 *
0-
02
b10 6
#821650000000
1!
1%
1-
12
#821660000000
0!
0%
b11 *
0-
02
b11 6
#821670000000
1!
1%
1-
12
15
#821680000000
0!
0%
b100 *
0-
02
b100 6
#821690000000
1!
1%
1-
12
#821700000000
0!
0%
b101 *
0-
02
b101 6
#821710000000
1!
1%
1-
12
#821720000000
0!
0%
b110 *
0-
02
b110 6
#821730000000
1!
1%
1-
12
#821740000000
0!
0%
b111 *
0-
02
b111 6
#821750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#821760000000
0!
0%
b0 *
0-
02
b0 6
#821770000000
1!
1%
1-
12
#821780000000
0!
0%
b1 *
0-
02
b1 6
#821790000000
1!
1%
1-
12
#821800000000
0!
0%
b10 *
0-
02
b10 6
#821810000000
1!
1%
1-
12
#821820000000
0!
0%
b11 *
0-
02
b11 6
#821830000000
1!
1%
1-
12
15
#821840000000
0!
0%
b100 *
0-
02
b100 6
#821850000000
1!
1%
1-
12
#821860000000
0!
0%
b101 *
0-
02
b101 6
#821870000000
1!
1%
1-
12
#821880000000
0!
0%
b110 *
0-
02
b110 6
#821890000000
1!
1%
1-
12
#821900000000
0!
0%
b111 *
0-
02
b111 6
#821910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#821920000000
0!
0%
b0 *
0-
02
b0 6
#821930000000
1!
1%
1-
12
#821940000000
0!
0%
b1 *
0-
02
b1 6
#821950000000
1!
1%
1-
12
#821960000000
0!
0%
b10 *
0-
02
b10 6
#821970000000
1!
1%
1-
12
#821980000000
0!
0%
b11 *
0-
02
b11 6
#821990000000
1!
1%
1-
12
15
#822000000000
0!
0%
b100 *
0-
02
b100 6
#822010000000
1!
1%
1-
12
#822020000000
0!
0%
b101 *
0-
02
b101 6
#822030000000
1!
1%
1-
12
#822040000000
0!
0%
b110 *
0-
02
b110 6
#822050000000
1!
1%
1-
12
#822060000000
0!
0%
b111 *
0-
02
b111 6
#822070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#822080000000
0!
0%
b0 *
0-
02
b0 6
#822090000000
1!
1%
1-
12
#822100000000
0!
0%
b1 *
0-
02
b1 6
#822110000000
1!
1%
1-
12
#822120000000
0!
0%
b10 *
0-
02
b10 6
#822130000000
1!
1%
1-
12
#822140000000
0!
0%
b11 *
0-
02
b11 6
#822150000000
1!
1%
1-
12
15
#822160000000
0!
0%
b100 *
0-
02
b100 6
#822170000000
1!
1%
1-
12
#822180000000
0!
0%
b101 *
0-
02
b101 6
#822190000000
1!
1%
1-
12
#822200000000
0!
0%
b110 *
0-
02
b110 6
#822210000000
1!
1%
1-
12
#822220000000
0!
0%
b111 *
0-
02
b111 6
#822230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#822240000000
0!
0%
b0 *
0-
02
b0 6
#822250000000
1!
1%
1-
12
#822260000000
0!
0%
b1 *
0-
02
b1 6
#822270000000
1!
1%
1-
12
#822280000000
0!
0%
b10 *
0-
02
b10 6
#822290000000
1!
1%
1-
12
#822300000000
0!
0%
b11 *
0-
02
b11 6
#822310000000
1!
1%
1-
12
15
#822320000000
0!
0%
b100 *
0-
02
b100 6
#822330000000
1!
1%
1-
12
#822340000000
0!
0%
b101 *
0-
02
b101 6
#822350000000
1!
1%
1-
12
#822360000000
0!
0%
b110 *
0-
02
b110 6
#822370000000
1!
1%
1-
12
#822380000000
0!
0%
b111 *
0-
02
b111 6
#822390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#822400000000
0!
0%
b0 *
0-
02
b0 6
#822410000000
1!
1%
1-
12
#822420000000
0!
0%
b1 *
0-
02
b1 6
#822430000000
1!
1%
1-
12
#822440000000
0!
0%
b10 *
0-
02
b10 6
#822450000000
1!
1%
1-
12
#822460000000
0!
0%
b11 *
0-
02
b11 6
#822470000000
1!
1%
1-
12
15
#822480000000
0!
0%
b100 *
0-
02
b100 6
#822490000000
1!
1%
1-
12
#822500000000
0!
0%
b101 *
0-
02
b101 6
#822510000000
1!
1%
1-
12
#822520000000
0!
0%
b110 *
0-
02
b110 6
#822530000000
1!
1%
1-
12
#822540000000
0!
0%
b111 *
0-
02
b111 6
#822550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#822560000000
0!
0%
b0 *
0-
02
b0 6
#822570000000
1!
1%
1-
12
#822580000000
0!
0%
b1 *
0-
02
b1 6
#822590000000
1!
1%
1-
12
#822600000000
0!
0%
b10 *
0-
02
b10 6
#822610000000
1!
1%
1-
12
#822620000000
0!
0%
b11 *
0-
02
b11 6
#822630000000
1!
1%
1-
12
15
#822640000000
0!
0%
b100 *
0-
02
b100 6
#822650000000
1!
1%
1-
12
#822660000000
0!
0%
b101 *
0-
02
b101 6
#822670000000
1!
1%
1-
12
#822680000000
0!
0%
b110 *
0-
02
b110 6
#822690000000
1!
1%
1-
12
#822700000000
0!
0%
b111 *
0-
02
b111 6
#822710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#822720000000
0!
0%
b0 *
0-
02
b0 6
#822730000000
1!
1%
1-
12
#822740000000
0!
0%
b1 *
0-
02
b1 6
#822750000000
1!
1%
1-
12
#822760000000
0!
0%
b10 *
0-
02
b10 6
#822770000000
1!
1%
1-
12
#822780000000
0!
0%
b11 *
0-
02
b11 6
#822790000000
1!
1%
1-
12
15
#822800000000
0!
0%
b100 *
0-
02
b100 6
#822810000000
1!
1%
1-
12
#822820000000
0!
0%
b101 *
0-
02
b101 6
#822830000000
1!
1%
1-
12
#822840000000
0!
0%
b110 *
0-
02
b110 6
#822850000000
1!
1%
1-
12
#822860000000
0!
0%
b111 *
0-
02
b111 6
#822870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#822880000000
0!
0%
b0 *
0-
02
b0 6
#822890000000
1!
1%
1-
12
#822900000000
0!
0%
b1 *
0-
02
b1 6
#822910000000
1!
1%
1-
12
#822920000000
0!
0%
b10 *
0-
02
b10 6
#822930000000
1!
1%
1-
12
#822940000000
0!
0%
b11 *
0-
02
b11 6
#822950000000
1!
1%
1-
12
15
#822960000000
0!
0%
b100 *
0-
02
b100 6
#822970000000
1!
1%
1-
12
#822980000000
0!
0%
b101 *
0-
02
b101 6
#822990000000
1!
1%
1-
12
#823000000000
0!
0%
b110 *
0-
02
b110 6
#823010000000
1!
1%
1-
12
#823020000000
0!
0%
b111 *
0-
02
b111 6
#823030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#823040000000
0!
0%
b0 *
0-
02
b0 6
#823050000000
1!
1%
1-
12
#823060000000
0!
0%
b1 *
0-
02
b1 6
#823070000000
1!
1%
1-
12
#823080000000
0!
0%
b10 *
0-
02
b10 6
#823090000000
1!
1%
1-
12
#823100000000
0!
0%
b11 *
0-
02
b11 6
#823110000000
1!
1%
1-
12
15
#823120000000
0!
0%
b100 *
0-
02
b100 6
#823130000000
1!
1%
1-
12
#823140000000
0!
0%
b101 *
0-
02
b101 6
#823150000000
1!
1%
1-
12
#823160000000
0!
0%
b110 *
0-
02
b110 6
#823170000000
1!
1%
1-
12
#823180000000
0!
0%
b111 *
0-
02
b111 6
#823190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#823200000000
0!
0%
b0 *
0-
02
b0 6
#823210000000
1!
1%
1-
12
#823220000000
0!
0%
b1 *
0-
02
b1 6
#823230000000
1!
1%
1-
12
#823240000000
0!
0%
b10 *
0-
02
b10 6
#823250000000
1!
1%
1-
12
#823260000000
0!
0%
b11 *
0-
02
b11 6
#823270000000
1!
1%
1-
12
15
#823280000000
0!
0%
b100 *
0-
02
b100 6
#823290000000
1!
1%
1-
12
#823300000000
0!
0%
b101 *
0-
02
b101 6
#823310000000
1!
1%
1-
12
#823320000000
0!
0%
b110 *
0-
02
b110 6
#823330000000
1!
1%
1-
12
#823340000000
0!
0%
b111 *
0-
02
b111 6
#823350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#823360000000
0!
0%
b0 *
0-
02
b0 6
#823370000000
1!
1%
1-
12
#823380000000
0!
0%
b1 *
0-
02
b1 6
#823390000000
1!
1%
1-
12
#823400000000
0!
0%
b10 *
0-
02
b10 6
#823410000000
1!
1%
1-
12
#823420000000
0!
0%
b11 *
0-
02
b11 6
#823430000000
1!
1%
1-
12
15
#823440000000
0!
0%
b100 *
0-
02
b100 6
#823450000000
1!
1%
1-
12
#823460000000
0!
0%
b101 *
0-
02
b101 6
#823470000000
1!
1%
1-
12
#823480000000
0!
0%
b110 *
0-
02
b110 6
#823490000000
1!
1%
1-
12
#823500000000
0!
0%
b111 *
0-
02
b111 6
#823510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#823520000000
0!
0%
b0 *
0-
02
b0 6
#823530000000
1!
1%
1-
12
#823540000000
0!
0%
b1 *
0-
02
b1 6
#823550000000
1!
1%
1-
12
#823560000000
0!
0%
b10 *
0-
02
b10 6
#823570000000
1!
1%
1-
12
#823580000000
0!
0%
b11 *
0-
02
b11 6
#823590000000
1!
1%
1-
12
15
#823600000000
0!
0%
b100 *
0-
02
b100 6
#823610000000
1!
1%
1-
12
#823620000000
0!
0%
b101 *
0-
02
b101 6
#823630000000
1!
1%
1-
12
#823640000000
0!
0%
b110 *
0-
02
b110 6
#823650000000
1!
1%
1-
12
#823660000000
0!
0%
b111 *
0-
02
b111 6
#823670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#823680000000
0!
0%
b0 *
0-
02
b0 6
#823690000000
1!
1%
1-
12
#823700000000
0!
0%
b1 *
0-
02
b1 6
#823710000000
1!
1%
1-
12
#823720000000
0!
0%
b10 *
0-
02
b10 6
#823730000000
1!
1%
1-
12
#823740000000
0!
0%
b11 *
0-
02
b11 6
#823750000000
1!
1%
1-
12
15
#823760000000
0!
0%
b100 *
0-
02
b100 6
#823770000000
1!
1%
1-
12
#823780000000
0!
0%
b101 *
0-
02
b101 6
#823790000000
1!
1%
1-
12
#823800000000
0!
0%
b110 *
0-
02
b110 6
#823810000000
1!
1%
1-
12
#823820000000
0!
0%
b111 *
0-
02
b111 6
#823830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#823840000000
0!
0%
b0 *
0-
02
b0 6
#823850000000
1!
1%
1-
12
#823860000000
0!
0%
b1 *
0-
02
b1 6
#823870000000
1!
1%
1-
12
#823880000000
0!
0%
b10 *
0-
02
b10 6
#823890000000
1!
1%
1-
12
#823900000000
0!
0%
b11 *
0-
02
b11 6
#823910000000
1!
1%
1-
12
15
#823920000000
0!
0%
b100 *
0-
02
b100 6
#823930000000
1!
1%
1-
12
#823940000000
0!
0%
b101 *
0-
02
b101 6
#823950000000
1!
1%
1-
12
#823960000000
0!
0%
b110 *
0-
02
b110 6
#823970000000
1!
1%
1-
12
#823980000000
0!
0%
b111 *
0-
02
b111 6
#823990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#824000000000
0!
0%
b0 *
0-
02
b0 6
#824010000000
1!
1%
1-
12
#824020000000
0!
0%
b1 *
0-
02
b1 6
#824030000000
1!
1%
1-
12
#824040000000
0!
0%
b10 *
0-
02
b10 6
#824050000000
1!
1%
1-
12
#824060000000
0!
0%
b11 *
0-
02
b11 6
#824070000000
1!
1%
1-
12
15
#824080000000
0!
0%
b100 *
0-
02
b100 6
#824090000000
1!
1%
1-
12
#824100000000
0!
0%
b101 *
0-
02
b101 6
#824110000000
1!
1%
1-
12
#824120000000
0!
0%
b110 *
0-
02
b110 6
#824130000000
1!
1%
1-
12
#824140000000
0!
0%
b111 *
0-
02
b111 6
#824150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#824160000000
0!
0%
b0 *
0-
02
b0 6
#824170000000
1!
1%
1-
12
#824180000000
0!
0%
b1 *
0-
02
b1 6
#824190000000
1!
1%
1-
12
#824200000000
0!
0%
b10 *
0-
02
b10 6
#824210000000
1!
1%
1-
12
#824220000000
0!
0%
b11 *
0-
02
b11 6
#824230000000
1!
1%
1-
12
15
#824240000000
0!
0%
b100 *
0-
02
b100 6
#824250000000
1!
1%
1-
12
#824260000000
0!
0%
b101 *
0-
02
b101 6
#824270000000
1!
1%
1-
12
#824280000000
0!
0%
b110 *
0-
02
b110 6
#824290000000
1!
1%
1-
12
#824300000000
0!
0%
b111 *
0-
02
b111 6
#824310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#824320000000
0!
0%
b0 *
0-
02
b0 6
#824330000000
1!
1%
1-
12
#824340000000
0!
0%
b1 *
0-
02
b1 6
#824350000000
1!
1%
1-
12
#824360000000
0!
0%
b10 *
0-
02
b10 6
#824370000000
1!
1%
1-
12
#824380000000
0!
0%
b11 *
0-
02
b11 6
#824390000000
1!
1%
1-
12
15
#824400000000
0!
0%
b100 *
0-
02
b100 6
#824410000000
1!
1%
1-
12
#824420000000
0!
0%
b101 *
0-
02
b101 6
#824430000000
1!
1%
1-
12
#824440000000
0!
0%
b110 *
0-
02
b110 6
#824450000000
1!
1%
1-
12
#824460000000
0!
0%
b111 *
0-
02
b111 6
#824470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#824480000000
0!
0%
b0 *
0-
02
b0 6
#824490000000
1!
1%
1-
12
#824500000000
0!
0%
b1 *
0-
02
b1 6
#824510000000
1!
1%
1-
12
#824520000000
0!
0%
b10 *
0-
02
b10 6
#824530000000
1!
1%
1-
12
#824540000000
0!
0%
b11 *
0-
02
b11 6
#824550000000
1!
1%
1-
12
15
#824560000000
0!
0%
b100 *
0-
02
b100 6
#824570000000
1!
1%
1-
12
#824580000000
0!
0%
b101 *
0-
02
b101 6
#824590000000
1!
1%
1-
12
#824600000000
0!
0%
b110 *
0-
02
b110 6
#824610000000
1!
1%
1-
12
#824620000000
0!
0%
b111 *
0-
02
b111 6
#824630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#824640000000
0!
0%
b0 *
0-
02
b0 6
#824650000000
1!
1%
1-
12
#824660000000
0!
0%
b1 *
0-
02
b1 6
#824670000000
1!
1%
1-
12
#824680000000
0!
0%
b10 *
0-
02
b10 6
#824690000000
1!
1%
1-
12
#824700000000
0!
0%
b11 *
0-
02
b11 6
#824710000000
1!
1%
1-
12
15
#824720000000
0!
0%
b100 *
0-
02
b100 6
#824730000000
1!
1%
1-
12
#824740000000
0!
0%
b101 *
0-
02
b101 6
#824750000000
1!
1%
1-
12
#824760000000
0!
0%
b110 *
0-
02
b110 6
#824770000000
1!
1%
1-
12
#824780000000
0!
0%
b111 *
0-
02
b111 6
#824790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#824800000000
0!
0%
b0 *
0-
02
b0 6
#824810000000
1!
1%
1-
12
#824820000000
0!
0%
b1 *
0-
02
b1 6
#824830000000
1!
1%
1-
12
#824840000000
0!
0%
b10 *
0-
02
b10 6
#824850000000
1!
1%
1-
12
#824860000000
0!
0%
b11 *
0-
02
b11 6
#824870000000
1!
1%
1-
12
15
#824880000000
0!
0%
b100 *
0-
02
b100 6
#824890000000
1!
1%
1-
12
#824900000000
0!
0%
b101 *
0-
02
b101 6
#824910000000
1!
1%
1-
12
#824920000000
0!
0%
b110 *
0-
02
b110 6
#824930000000
1!
1%
1-
12
#824940000000
0!
0%
b111 *
0-
02
b111 6
#824950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#824960000000
0!
0%
b0 *
0-
02
b0 6
#824970000000
1!
1%
1-
12
#824980000000
0!
0%
b1 *
0-
02
b1 6
#824990000000
1!
1%
1-
12
#825000000000
0!
0%
b10 *
0-
02
b10 6
#825010000000
1!
1%
1-
12
#825020000000
0!
0%
b11 *
0-
02
b11 6
#825030000000
1!
1%
1-
12
15
#825040000000
0!
0%
b100 *
0-
02
b100 6
#825050000000
1!
1%
1-
12
#825060000000
0!
0%
b101 *
0-
02
b101 6
#825070000000
1!
1%
1-
12
#825080000000
0!
0%
b110 *
0-
02
b110 6
#825090000000
1!
1%
1-
12
#825100000000
0!
0%
b111 *
0-
02
b111 6
#825110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#825120000000
0!
0%
b0 *
0-
02
b0 6
#825130000000
1!
1%
1-
12
#825140000000
0!
0%
b1 *
0-
02
b1 6
#825150000000
1!
1%
1-
12
#825160000000
0!
0%
b10 *
0-
02
b10 6
#825170000000
1!
1%
1-
12
#825180000000
0!
0%
b11 *
0-
02
b11 6
#825190000000
1!
1%
1-
12
15
#825200000000
0!
0%
b100 *
0-
02
b100 6
#825210000000
1!
1%
1-
12
#825220000000
0!
0%
b101 *
0-
02
b101 6
#825230000000
1!
1%
1-
12
#825240000000
0!
0%
b110 *
0-
02
b110 6
#825250000000
1!
1%
1-
12
#825260000000
0!
0%
b111 *
0-
02
b111 6
#825270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#825280000000
0!
0%
b0 *
0-
02
b0 6
#825290000000
1!
1%
1-
12
#825300000000
0!
0%
b1 *
0-
02
b1 6
#825310000000
1!
1%
1-
12
#825320000000
0!
0%
b10 *
0-
02
b10 6
#825330000000
1!
1%
1-
12
#825340000000
0!
0%
b11 *
0-
02
b11 6
#825350000000
1!
1%
1-
12
15
#825360000000
0!
0%
b100 *
0-
02
b100 6
#825370000000
1!
1%
1-
12
#825380000000
0!
0%
b101 *
0-
02
b101 6
#825390000000
1!
1%
1-
12
#825400000000
0!
0%
b110 *
0-
02
b110 6
#825410000000
1!
1%
1-
12
#825420000000
0!
0%
b111 *
0-
02
b111 6
#825430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#825440000000
0!
0%
b0 *
0-
02
b0 6
#825450000000
1!
1%
1-
12
#825460000000
0!
0%
b1 *
0-
02
b1 6
#825470000000
1!
1%
1-
12
#825480000000
0!
0%
b10 *
0-
02
b10 6
#825490000000
1!
1%
1-
12
#825500000000
0!
0%
b11 *
0-
02
b11 6
#825510000000
1!
1%
1-
12
15
#825520000000
0!
0%
b100 *
0-
02
b100 6
#825530000000
1!
1%
1-
12
#825540000000
0!
0%
b101 *
0-
02
b101 6
#825550000000
1!
1%
1-
12
#825560000000
0!
0%
b110 *
0-
02
b110 6
#825570000000
1!
1%
1-
12
#825580000000
0!
0%
b111 *
0-
02
b111 6
#825590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#825600000000
0!
0%
b0 *
0-
02
b0 6
#825610000000
1!
1%
1-
12
#825620000000
0!
0%
b1 *
0-
02
b1 6
#825630000000
1!
1%
1-
12
#825640000000
0!
0%
b10 *
0-
02
b10 6
#825650000000
1!
1%
1-
12
#825660000000
0!
0%
b11 *
0-
02
b11 6
#825670000000
1!
1%
1-
12
15
#825680000000
0!
0%
b100 *
0-
02
b100 6
#825690000000
1!
1%
1-
12
#825700000000
0!
0%
b101 *
0-
02
b101 6
#825710000000
1!
1%
1-
12
#825720000000
0!
0%
b110 *
0-
02
b110 6
#825730000000
1!
1%
1-
12
#825740000000
0!
0%
b111 *
0-
02
b111 6
#825750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#825760000000
0!
0%
b0 *
0-
02
b0 6
#825770000000
1!
1%
1-
12
#825780000000
0!
0%
b1 *
0-
02
b1 6
#825790000000
1!
1%
1-
12
#825800000000
0!
0%
b10 *
0-
02
b10 6
#825810000000
1!
1%
1-
12
#825820000000
0!
0%
b11 *
0-
02
b11 6
#825830000000
1!
1%
1-
12
15
#825840000000
0!
0%
b100 *
0-
02
b100 6
#825850000000
1!
1%
1-
12
#825860000000
0!
0%
b101 *
0-
02
b101 6
#825870000000
1!
1%
1-
12
#825880000000
0!
0%
b110 *
0-
02
b110 6
#825890000000
1!
1%
1-
12
#825900000000
0!
0%
b111 *
0-
02
b111 6
#825910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#825920000000
0!
0%
b0 *
0-
02
b0 6
#825930000000
1!
1%
1-
12
#825940000000
0!
0%
b1 *
0-
02
b1 6
#825950000000
1!
1%
1-
12
#825960000000
0!
0%
b10 *
0-
02
b10 6
#825970000000
1!
1%
1-
12
#825980000000
0!
0%
b11 *
0-
02
b11 6
#825990000000
1!
1%
1-
12
15
#826000000000
0!
0%
b100 *
0-
02
b100 6
#826010000000
1!
1%
1-
12
#826020000000
0!
0%
b101 *
0-
02
b101 6
#826030000000
1!
1%
1-
12
#826040000000
0!
0%
b110 *
0-
02
b110 6
#826050000000
1!
1%
1-
12
#826060000000
0!
0%
b111 *
0-
02
b111 6
#826070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#826080000000
0!
0%
b0 *
0-
02
b0 6
#826090000000
1!
1%
1-
12
#826100000000
0!
0%
b1 *
0-
02
b1 6
#826110000000
1!
1%
1-
12
#826120000000
0!
0%
b10 *
0-
02
b10 6
#826130000000
1!
1%
1-
12
#826140000000
0!
0%
b11 *
0-
02
b11 6
#826150000000
1!
1%
1-
12
15
#826160000000
0!
0%
b100 *
0-
02
b100 6
#826170000000
1!
1%
1-
12
#826180000000
0!
0%
b101 *
0-
02
b101 6
#826190000000
1!
1%
1-
12
#826200000000
0!
0%
b110 *
0-
02
b110 6
#826210000000
1!
1%
1-
12
#826220000000
0!
0%
b111 *
0-
02
b111 6
#826230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#826240000000
0!
0%
b0 *
0-
02
b0 6
#826250000000
1!
1%
1-
12
#826260000000
0!
0%
b1 *
0-
02
b1 6
#826270000000
1!
1%
1-
12
#826280000000
0!
0%
b10 *
0-
02
b10 6
#826290000000
1!
1%
1-
12
#826300000000
0!
0%
b11 *
0-
02
b11 6
#826310000000
1!
1%
1-
12
15
#826320000000
0!
0%
b100 *
0-
02
b100 6
#826330000000
1!
1%
1-
12
#826340000000
0!
0%
b101 *
0-
02
b101 6
#826350000000
1!
1%
1-
12
#826360000000
0!
0%
b110 *
0-
02
b110 6
#826370000000
1!
1%
1-
12
#826380000000
0!
0%
b111 *
0-
02
b111 6
#826390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#826400000000
0!
0%
b0 *
0-
02
b0 6
#826410000000
1!
1%
1-
12
#826420000000
0!
0%
b1 *
0-
02
b1 6
#826430000000
1!
1%
1-
12
#826440000000
0!
0%
b10 *
0-
02
b10 6
#826450000000
1!
1%
1-
12
#826460000000
0!
0%
b11 *
0-
02
b11 6
#826470000000
1!
1%
1-
12
15
#826480000000
0!
0%
b100 *
0-
02
b100 6
#826490000000
1!
1%
1-
12
#826500000000
0!
0%
b101 *
0-
02
b101 6
#826510000000
1!
1%
1-
12
#826520000000
0!
0%
b110 *
0-
02
b110 6
#826530000000
1!
1%
1-
12
#826540000000
0!
0%
b111 *
0-
02
b111 6
#826550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#826560000000
0!
0%
b0 *
0-
02
b0 6
#826570000000
1!
1%
1-
12
#826580000000
0!
0%
b1 *
0-
02
b1 6
#826590000000
1!
1%
1-
12
#826600000000
0!
0%
b10 *
0-
02
b10 6
#826610000000
1!
1%
1-
12
#826620000000
0!
0%
b11 *
0-
02
b11 6
#826630000000
1!
1%
1-
12
15
#826640000000
0!
0%
b100 *
0-
02
b100 6
#826650000000
1!
1%
1-
12
#826660000000
0!
0%
b101 *
0-
02
b101 6
#826670000000
1!
1%
1-
12
#826680000000
0!
0%
b110 *
0-
02
b110 6
#826690000000
1!
1%
1-
12
#826700000000
0!
0%
b111 *
0-
02
b111 6
#826710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#826720000000
0!
0%
b0 *
0-
02
b0 6
#826730000000
1!
1%
1-
12
#826740000000
0!
0%
b1 *
0-
02
b1 6
#826750000000
1!
1%
1-
12
#826760000000
0!
0%
b10 *
0-
02
b10 6
#826770000000
1!
1%
1-
12
#826780000000
0!
0%
b11 *
0-
02
b11 6
#826790000000
1!
1%
1-
12
15
#826800000000
0!
0%
b100 *
0-
02
b100 6
#826810000000
1!
1%
1-
12
#826820000000
0!
0%
b101 *
0-
02
b101 6
#826830000000
1!
1%
1-
12
#826840000000
0!
0%
b110 *
0-
02
b110 6
#826850000000
1!
1%
1-
12
#826860000000
0!
0%
b111 *
0-
02
b111 6
#826870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#826880000000
0!
0%
b0 *
0-
02
b0 6
#826890000000
1!
1%
1-
12
#826900000000
0!
0%
b1 *
0-
02
b1 6
#826910000000
1!
1%
1-
12
#826920000000
0!
0%
b10 *
0-
02
b10 6
#826930000000
1!
1%
1-
12
#826940000000
0!
0%
b11 *
0-
02
b11 6
#826950000000
1!
1%
1-
12
15
#826960000000
0!
0%
b100 *
0-
02
b100 6
#826970000000
1!
1%
1-
12
#826980000000
0!
0%
b101 *
0-
02
b101 6
#826990000000
1!
1%
1-
12
#827000000000
0!
0%
b110 *
0-
02
b110 6
#827010000000
1!
1%
1-
12
#827020000000
0!
0%
b111 *
0-
02
b111 6
#827030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#827040000000
0!
0%
b0 *
0-
02
b0 6
#827050000000
1!
1%
1-
12
#827060000000
0!
0%
b1 *
0-
02
b1 6
#827070000000
1!
1%
1-
12
#827080000000
0!
0%
b10 *
0-
02
b10 6
#827090000000
1!
1%
1-
12
#827100000000
0!
0%
b11 *
0-
02
b11 6
#827110000000
1!
1%
1-
12
15
#827120000000
0!
0%
b100 *
0-
02
b100 6
#827130000000
1!
1%
1-
12
#827140000000
0!
0%
b101 *
0-
02
b101 6
#827150000000
1!
1%
1-
12
#827160000000
0!
0%
b110 *
0-
02
b110 6
#827170000000
1!
1%
1-
12
#827180000000
0!
0%
b111 *
0-
02
b111 6
#827190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#827200000000
0!
0%
b0 *
0-
02
b0 6
#827210000000
1!
1%
1-
12
#827220000000
0!
0%
b1 *
0-
02
b1 6
#827230000000
1!
1%
1-
12
#827240000000
0!
0%
b10 *
0-
02
b10 6
#827250000000
1!
1%
1-
12
#827260000000
0!
0%
b11 *
0-
02
b11 6
#827270000000
1!
1%
1-
12
15
#827280000000
0!
0%
b100 *
0-
02
b100 6
#827290000000
1!
1%
1-
12
#827300000000
0!
0%
b101 *
0-
02
b101 6
#827310000000
1!
1%
1-
12
#827320000000
0!
0%
b110 *
0-
02
b110 6
#827330000000
1!
1%
1-
12
#827340000000
0!
0%
b111 *
0-
02
b111 6
#827350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#827360000000
0!
0%
b0 *
0-
02
b0 6
#827370000000
1!
1%
1-
12
#827380000000
0!
0%
b1 *
0-
02
b1 6
#827390000000
1!
1%
1-
12
#827400000000
0!
0%
b10 *
0-
02
b10 6
#827410000000
1!
1%
1-
12
#827420000000
0!
0%
b11 *
0-
02
b11 6
#827430000000
1!
1%
1-
12
15
#827440000000
0!
0%
b100 *
0-
02
b100 6
#827450000000
1!
1%
1-
12
#827460000000
0!
0%
b101 *
0-
02
b101 6
#827470000000
1!
1%
1-
12
#827480000000
0!
0%
b110 *
0-
02
b110 6
#827490000000
1!
1%
1-
12
#827500000000
0!
0%
b111 *
0-
02
b111 6
#827510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#827520000000
0!
0%
b0 *
0-
02
b0 6
#827530000000
1!
1%
1-
12
#827540000000
0!
0%
b1 *
0-
02
b1 6
#827550000000
1!
1%
1-
12
#827560000000
0!
0%
b10 *
0-
02
b10 6
#827570000000
1!
1%
1-
12
#827580000000
0!
0%
b11 *
0-
02
b11 6
#827590000000
1!
1%
1-
12
15
#827600000000
0!
0%
b100 *
0-
02
b100 6
#827610000000
1!
1%
1-
12
#827620000000
0!
0%
b101 *
0-
02
b101 6
#827630000000
1!
1%
1-
12
#827640000000
0!
0%
b110 *
0-
02
b110 6
#827650000000
1!
1%
1-
12
#827660000000
0!
0%
b111 *
0-
02
b111 6
#827670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#827680000000
0!
0%
b0 *
0-
02
b0 6
#827690000000
1!
1%
1-
12
#827700000000
0!
0%
b1 *
0-
02
b1 6
#827710000000
1!
1%
1-
12
#827720000000
0!
0%
b10 *
0-
02
b10 6
#827730000000
1!
1%
1-
12
#827740000000
0!
0%
b11 *
0-
02
b11 6
#827750000000
1!
1%
1-
12
15
#827760000000
0!
0%
b100 *
0-
02
b100 6
#827770000000
1!
1%
1-
12
#827780000000
0!
0%
b101 *
0-
02
b101 6
#827790000000
1!
1%
1-
12
#827800000000
0!
0%
b110 *
0-
02
b110 6
#827810000000
1!
1%
1-
12
#827820000000
0!
0%
b111 *
0-
02
b111 6
#827830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#827840000000
0!
0%
b0 *
0-
02
b0 6
#827850000000
1!
1%
1-
12
#827860000000
0!
0%
b1 *
0-
02
b1 6
#827870000000
1!
1%
1-
12
#827880000000
0!
0%
b10 *
0-
02
b10 6
#827890000000
1!
1%
1-
12
#827900000000
0!
0%
b11 *
0-
02
b11 6
#827910000000
1!
1%
1-
12
15
#827920000000
0!
0%
b100 *
0-
02
b100 6
#827930000000
1!
1%
1-
12
#827940000000
0!
0%
b101 *
0-
02
b101 6
#827950000000
1!
1%
1-
12
#827960000000
0!
0%
b110 *
0-
02
b110 6
#827970000000
1!
1%
1-
12
#827980000000
0!
0%
b111 *
0-
02
b111 6
#827990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#828000000000
0!
0%
b0 *
0-
02
b0 6
#828010000000
1!
1%
1-
12
#828020000000
0!
0%
b1 *
0-
02
b1 6
#828030000000
1!
1%
1-
12
#828040000000
0!
0%
b10 *
0-
02
b10 6
#828050000000
1!
1%
1-
12
#828060000000
0!
0%
b11 *
0-
02
b11 6
#828070000000
1!
1%
1-
12
15
#828080000000
0!
0%
b100 *
0-
02
b100 6
#828090000000
1!
1%
1-
12
#828100000000
0!
0%
b101 *
0-
02
b101 6
#828110000000
1!
1%
1-
12
#828120000000
0!
0%
b110 *
0-
02
b110 6
#828130000000
1!
1%
1-
12
#828140000000
0!
0%
b111 *
0-
02
b111 6
#828150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#828160000000
0!
0%
b0 *
0-
02
b0 6
#828170000000
1!
1%
1-
12
#828180000000
0!
0%
b1 *
0-
02
b1 6
#828190000000
1!
1%
1-
12
#828200000000
0!
0%
b10 *
0-
02
b10 6
#828210000000
1!
1%
1-
12
#828220000000
0!
0%
b11 *
0-
02
b11 6
#828230000000
1!
1%
1-
12
15
#828240000000
0!
0%
b100 *
0-
02
b100 6
#828250000000
1!
1%
1-
12
#828260000000
0!
0%
b101 *
0-
02
b101 6
#828270000000
1!
1%
1-
12
#828280000000
0!
0%
b110 *
0-
02
b110 6
#828290000000
1!
1%
1-
12
#828300000000
0!
0%
b111 *
0-
02
b111 6
#828310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#828320000000
0!
0%
b0 *
0-
02
b0 6
#828330000000
1!
1%
1-
12
#828340000000
0!
0%
b1 *
0-
02
b1 6
#828350000000
1!
1%
1-
12
#828360000000
0!
0%
b10 *
0-
02
b10 6
#828370000000
1!
1%
1-
12
#828380000000
0!
0%
b11 *
0-
02
b11 6
#828390000000
1!
1%
1-
12
15
#828400000000
0!
0%
b100 *
0-
02
b100 6
#828410000000
1!
1%
1-
12
#828420000000
0!
0%
b101 *
0-
02
b101 6
#828430000000
1!
1%
1-
12
#828440000000
0!
0%
b110 *
0-
02
b110 6
#828450000000
1!
1%
1-
12
#828460000000
0!
0%
b111 *
0-
02
b111 6
#828470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#828480000000
0!
0%
b0 *
0-
02
b0 6
#828490000000
1!
1%
1-
12
#828500000000
0!
0%
b1 *
0-
02
b1 6
#828510000000
1!
1%
1-
12
#828520000000
0!
0%
b10 *
0-
02
b10 6
#828530000000
1!
1%
1-
12
#828540000000
0!
0%
b11 *
0-
02
b11 6
#828550000000
1!
1%
1-
12
15
#828560000000
0!
0%
b100 *
0-
02
b100 6
#828570000000
1!
1%
1-
12
#828580000000
0!
0%
b101 *
0-
02
b101 6
#828590000000
1!
1%
1-
12
#828600000000
0!
0%
b110 *
0-
02
b110 6
#828610000000
1!
1%
1-
12
#828620000000
0!
0%
b111 *
0-
02
b111 6
#828630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#828640000000
0!
0%
b0 *
0-
02
b0 6
#828650000000
1!
1%
1-
12
#828660000000
0!
0%
b1 *
0-
02
b1 6
#828670000000
1!
1%
1-
12
#828680000000
0!
0%
b10 *
0-
02
b10 6
#828690000000
1!
1%
1-
12
#828700000000
0!
0%
b11 *
0-
02
b11 6
#828710000000
1!
1%
1-
12
15
#828720000000
0!
0%
b100 *
0-
02
b100 6
#828730000000
1!
1%
1-
12
#828740000000
0!
0%
b101 *
0-
02
b101 6
#828750000000
1!
1%
1-
12
#828760000000
0!
0%
b110 *
0-
02
b110 6
#828770000000
1!
1%
1-
12
#828780000000
0!
0%
b111 *
0-
02
b111 6
#828790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#828800000000
0!
0%
b0 *
0-
02
b0 6
#828810000000
1!
1%
1-
12
#828820000000
0!
0%
b1 *
0-
02
b1 6
#828830000000
1!
1%
1-
12
#828840000000
0!
0%
b10 *
0-
02
b10 6
#828850000000
1!
1%
1-
12
#828860000000
0!
0%
b11 *
0-
02
b11 6
#828870000000
1!
1%
1-
12
15
#828880000000
0!
0%
b100 *
0-
02
b100 6
#828890000000
1!
1%
1-
12
#828900000000
0!
0%
b101 *
0-
02
b101 6
#828910000000
1!
1%
1-
12
#828920000000
0!
0%
b110 *
0-
02
b110 6
#828930000000
1!
1%
1-
12
#828940000000
0!
0%
b111 *
0-
02
b111 6
#828950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#828960000000
0!
0%
b0 *
0-
02
b0 6
#828970000000
1!
1%
1-
12
#828980000000
0!
0%
b1 *
0-
02
b1 6
#828990000000
1!
1%
1-
12
#829000000000
0!
0%
b10 *
0-
02
b10 6
#829010000000
1!
1%
1-
12
#829020000000
0!
0%
b11 *
0-
02
b11 6
#829030000000
1!
1%
1-
12
15
#829040000000
0!
0%
b100 *
0-
02
b100 6
#829050000000
1!
1%
1-
12
#829060000000
0!
0%
b101 *
0-
02
b101 6
#829070000000
1!
1%
1-
12
#829080000000
0!
0%
b110 *
0-
02
b110 6
#829090000000
1!
1%
1-
12
#829100000000
0!
0%
b111 *
0-
02
b111 6
#829110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#829120000000
0!
0%
b0 *
0-
02
b0 6
#829130000000
1!
1%
1-
12
#829140000000
0!
0%
b1 *
0-
02
b1 6
#829150000000
1!
1%
1-
12
#829160000000
0!
0%
b10 *
0-
02
b10 6
#829170000000
1!
1%
1-
12
#829180000000
0!
0%
b11 *
0-
02
b11 6
#829190000000
1!
1%
1-
12
15
#829200000000
0!
0%
b100 *
0-
02
b100 6
#829210000000
1!
1%
1-
12
#829220000000
0!
0%
b101 *
0-
02
b101 6
#829230000000
1!
1%
1-
12
#829240000000
0!
0%
b110 *
0-
02
b110 6
#829250000000
1!
1%
1-
12
#829260000000
0!
0%
b111 *
0-
02
b111 6
#829270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#829280000000
0!
0%
b0 *
0-
02
b0 6
#829290000000
1!
1%
1-
12
#829300000000
0!
0%
b1 *
0-
02
b1 6
#829310000000
1!
1%
1-
12
#829320000000
0!
0%
b10 *
0-
02
b10 6
#829330000000
1!
1%
1-
12
#829340000000
0!
0%
b11 *
0-
02
b11 6
#829350000000
1!
1%
1-
12
15
#829360000000
0!
0%
b100 *
0-
02
b100 6
#829370000000
1!
1%
1-
12
#829380000000
0!
0%
b101 *
0-
02
b101 6
#829390000000
1!
1%
1-
12
#829400000000
0!
0%
b110 *
0-
02
b110 6
#829410000000
1!
1%
1-
12
#829420000000
0!
0%
b111 *
0-
02
b111 6
#829430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#829440000000
0!
0%
b0 *
0-
02
b0 6
#829450000000
1!
1%
1-
12
#829460000000
0!
0%
b1 *
0-
02
b1 6
#829470000000
1!
1%
1-
12
#829480000000
0!
0%
b10 *
0-
02
b10 6
#829490000000
1!
1%
1-
12
#829500000000
0!
0%
b11 *
0-
02
b11 6
#829510000000
1!
1%
1-
12
15
#829520000000
0!
0%
b100 *
0-
02
b100 6
#829530000000
1!
1%
1-
12
#829540000000
0!
0%
b101 *
0-
02
b101 6
#829550000000
1!
1%
1-
12
#829560000000
0!
0%
b110 *
0-
02
b110 6
#829570000000
1!
1%
1-
12
#829580000000
0!
0%
b111 *
0-
02
b111 6
#829590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#829600000000
0!
0%
b0 *
0-
02
b0 6
#829610000000
1!
1%
1-
12
#829620000000
0!
0%
b1 *
0-
02
b1 6
#829630000000
1!
1%
1-
12
#829640000000
0!
0%
b10 *
0-
02
b10 6
#829650000000
1!
1%
1-
12
#829660000000
0!
0%
b11 *
0-
02
b11 6
#829670000000
1!
1%
1-
12
15
#829680000000
0!
0%
b100 *
0-
02
b100 6
#829690000000
1!
1%
1-
12
#829700000000
0!
0%
b101 *
0-
02
b101 6
#829710000000
1!
1%
1-
12
#829720000000
0!
0%
b110 *
0-
02
b110 6
#829730000000
1!
1%
1-
12
#829740000000
0!
0%
b111 *
0-
02
b111 6
#829750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#829760000000
0!
0%
b0 *
0-
02
b0 6
#829770000000
1!
1%
1-
12
#829780000000
0!
0%
b1 *
0-
02
b1 6
#829790000000
1!
1%
1-
12
#829800000000
0!
0%
b10 *
0-
02
b10 6
#829810000000
1!
1%
1-
12
#829820000000
0!
0%
b11 *
0-
02
b11 6
#829830000000
1!
1%
1-
12
15
#829840000000
0!
0%
b100 *
0-
02
b100 6
#829850000000
1!
1%
1-
12
#829860000000
0!
0%
b101 *
0-
02
b101 6
#829870000000
1!
1%
1-
12
#829880000000
0!
0%
b110 *
0-
02
b110 6
#829890000000
1!
1%
1-
12
#829900000000
0!
0%
b111 *
0-
02
b111 6
#829910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#829920000000
0!
0%
b0 *
0-
02
b0 6
#829930000000
1!
1%
1-
12
#829940000000
0!
0%
b1 *
0-
02
b1 6
#829950000000
1!
1%
1-
12
#829960000000
0!
0%
b10 *
0-
02
b10 6
#829970000000
1!
1%
1-
12
#829980000000
0!
0%
b11 *
0-
02
b11 6
#829990000000
1!
1%
1-
12
15
#830000000000
0!
0%
b100 *
0-
02
b100 6
#830010000000
1!
1%
1-
12
#830020000000
0!
0%
b101 *
0-
02
b101 6
#830030000000
1!
1%
1-
12
#830040000000
0!
0%
b110 *
0-
02
b110 6
#830050000000
1!
1%
1-
12
#830060000000
0!
0%
b111 *
0-
02
b111 6
#830070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#830080000000
0!
0%
b0 *
0-
02
b0 6
#830090000000
1!
1%
1-
12
#830100000000
0!
0%
b1 *
0-
02
b1 6
#830110000000
1!
1%
1-
12
#830120000000
0!
0%
b10 *
0-
02
b10 6
#830130000000
1!
1%
1-
12
#830140000000
0!
0%
b11 *
0-
02
b11 6
#830150000000
1!
1%
1-
12
15
#830160000000
0!
0%
b100 *
0-
02
b100 6
#830170000000
1!
1%
1-
12
#830180000000
0!
0%
b101 *
0-
02
b101 6
#830190000000
1!
1%
1-
12
#830200000000
0!
0%
b110 *
0-
02
b110 6
#830210000000
1!
1%
1-
12
#830220000000
0!
0%
b111 *
0-
02
b111 6
#830230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#830240000000
0!
0%
b0 *
0-
02
b0 6
#830250000000
1!
1%
1-
12
#830260000000
0!
0%
b1 *
0-
02
b1 6
#830270000000
1!
1%
1-
12
#830280000000
0!
0%
b10 *
0-
02
b10 6
#830290000000
1!
1%
1-
12
#830300000000
0!
0%
b11 *
0-
02
b11 6
#830310000000
1!
1%
1-
12
15
#830320000000
0!
0%
b100 *
0-
02
b100 6
#830330000000
1!
1%
1-
12
#830340000000
0!
0%
b101 *
0-
02
b101 6
#830350000000
1!
1%
1-
12
#830360000000
0!
0%
b110 *
0-
02
b110 6
#830370000000
1!
1%
1-
12
#830380000000
0!
0%
b111 *
0-
02
b111 6
#830390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#830400000000
0!
0%
b0 *
0-
02
b0 6
#830410000000
1!
1%
1-
12
#830420000000
0!
0%
b1 *
0-
02
b1 6
#830430000000
1!
1%
1-
12
#830440000000
0!
0%
b10 *
0-
02
b10 6
#830450000000
1!
1%
1-
12
#830460000000
0!
0%
b11 *
0-
02
b11 6
#830470000000
1!
1%
1-
12
15
#830480000000
0!
0%
b100 *
0-
02
b100 6
#830490000000
1!
1%
1-
12
#830500000000
0!
0%
b101 *
0-
02
b101 6
#830510000000
1!
1%
1-
12
#830520000000
0!
0%
b110 *
0-
02
b110 6
#830530000000
1!
1%
1-
12
#830540000000
0!
0%
b111 *
0-
02
b111 6
#830550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#830560000000
0!
0%
b0 *
0-
02
b0 6
#830570000000
1!
1%
1-
12
#830580000000
0!
0%
b1 *
0-
02
b1 6
#830590000000
1!
1%
1-
12
#830600000000
0!
0%
b10 *
0-
02
b10 6
#830610000000
1!
1%
1-
12
#830620000000
0!
0%
b11 *
0-
02
b11 6
#830630000000
1!
1%
1-
12
15
#830640000000
0!
0%
b100 *
0-
02
b100 6
#830650000000
1!
1%
1-
12
#830660000000
0!
0%
b101 *
0-
02
b101 6
#830670000000
1!
1%
1-
12
#830680000000
0!
0%
b110 *
0-
02
b110 6
#830690000000
1!
1%
1-
12
#830700000000
0!
0%
b111 *
0-
02
b111 6
#830710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#830720000000
0!
0%
b0 *
0-
02
b0 6
#830730000000
1!
1%
1-
12
#830740000000
0!
0%
b1 *
0-
02
b1 6
#830750000000
1!
1%
1-
12
#830760000000
0!
0%
b10 *
0-
02
b10 6
#830770000000
1!
1%
1-
12
#830780000000
0!
0%
b11 *
0-
02
b11 6
#830790000000
1!
1%
1-
12
15
#830800000000
0!
0%
b100 *
0-
02
b100 6
#830810000000
1!
1%
1-
12
#830820000000
0!
0%
b101 *
0-
02
b101 6
#830830000000
1!
1%
1-
12
#830840000000
0!
0%
b110 *
0-
02
b110 6
#830850000000
1!
1%
1-
12
#830860000000
0!
0%
b111 *
0-
02
b111 6
#830870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#830880000000
0!
0%
b0 *
0-
02
b0 6
#830890000000
1!
1%
1-
12
#830900000000
0!
0%
b1 *
0-
02
b1 6
#830910000000
1!
1%
1-
12
#830920000000
0!
0%
b10 *
0-
02
b10 6
#830930000000
1!
1%
1-
12
#830940000000
0!
0%
b11 *
0-
02
b11 6
#830950000000
1!
1%
1-
12
15
#830960000000
0!
0%
b100 *
0-
02
b100 6
#830970000000
1!
1%
1-
12
#830980000000
0!
0%
b101 *
0-
02
b101 6
#830990000000
1!
1%
1-
12
#831000000000
0!
0%
b110 *
0-
02
b110 6
#831010000000
1!
1%
1-
12
#831020000000
0!
0%
b111 *
0-
02
b111 6
#831030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#831040000000
0!
0%
b0 *
0-
02
b0 6
#831050000000
1!
1%
1-
12
#831060000000
0!
0%
b1 *
0-
02
b1 6
#831070000000
1!
1%
1-
12
#831080000000
0!
0%
b10 *
0-
02
b10 6
#831090000000
1!
1%
1-
12
#831100000000
0!
0%
b11 *
0-
02
b11 6
#831110000000
1!
1%
1-
12
15
#831120000000
0!
0%
b100 *
0-
02
b100 6
#831130000000
1!
1%
1-
12
#831140000000
0!
0%
b101 *
0-
02
b101 6
#831150000000
1!
1%
1-
12
#831160000000
0!
0%
b110 *
0-
02
b110 6
#831170000000
1!
1%
1-
12
#831180000000
0!
0%
b111 *
0-
02
b111 6
#831190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#831200000000
0!
0%
b0 *
0-
02
b0 6
#831210000000
1!
1%
1-
12
#831220000000
0!
0%
b1 *
0-
02
b1 6
#831230000000
1!
1%
1-
12
#831240000000
0!
0%
b10 *
0-
02
b10 6
#831250000000
1!
1%
1-
12
#831260000000
0!
0%
b11 *
0-
02
b11 6
#831270000000
1!
1%
1-
12
15
#831280000000
0!
0%
b100 *
0-
02
b100 6
#831290000000
1!
1%
1-
12
#831300000000
0!
0%
b101 *
0-
02
b101 6
#831310000000
1!
1%
1-
12
#831320000000
0!
0%
b110 *
0-
02
b110 6
#831330000000
1!
1%
1-
12
#831340000000
0!
0%
b111 *
0-
02
b111 6
#831350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#831360000000
0!
0%
b0 *
0-
02
b0 6
#831370000000
1!
1%
1-
12
#831380000000
0!
0%
b1 *
0-
02
b1 6
#831390000000
1!
1%
1-
12
#831400000000
0!
0%
b10 *
0-
02
b10 6
#831410000000
1!
1%
1-
12
#831420000000
0!
0%
b11 *
0-
02
b11 6
#831430000000
1!
1%
1-
12
15
#831440000000
0!
0%
b100 *
0-
02
b100 6
#831450000000
1!
1%
1-
12
#831460000000
0!
0%
b101 *
0-
02
b101 6
#831470000000
1!
1%
1-
12
#831480000000
0!
0%
b110 *
0-
02
b110 6
#831490000000
1!
1%
1-
12
#831500000000
0!
0%
b111 *
0-
02
b111 6
#831510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#831520000000
0!
0%
b0 *
0-
02
b0 6
#831530000000
1!
1%
1-
12
#831540000000
0!
0%
b1 *
0-
02
b1 6
#831550000000
1!
1%
1-
12
#831560000000
0!
0%
b10 *
0-
02
b10 6
#831570000000
1!
1%
1-
12
#831580000000
0!
0%
b11 *
0-
02
b11 6
#831590000000
1!
1%
1-
12
15
#831600000000
0!
0%
b100 *
0-
02
b100 6
#831610000000
1!
1%
1-
12
#831620000000
0!
0%
b101 *
0-
02
b101 6
#831630000000
1!
1%
1-
12
#831640000000
0!
0%
b110 *
0-
02
b110 6
#831650000000
1!
1%
1-
12
#831660000000
0!
0%
b111 *
0-
02
b111 6
#831670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#831680000000
0!
0%
b0 *
0-
02
b0 6
#831690000000
1!
1%
1-
12
#831700000000
0!
0%
b1 *
0-
02
b1 6
#831710000000
1!
1%
1-
12
#831720000000
0!
0%
b10 *
0-
02
b10 6
#831730000000
1!
1%
1-
12
#831740000000
0!
0%
b11 *
0-
02
b11 6
#831750000000
1!
1%
1-
12
15
#831760000000
0!
0%
b100 *
0-
02
b100 6
#831770000000
1!
1%
1-
12
#831780000000
0!
0%
b101 *
0-
02
b101 6
#831790000000
1!
1%
1-
12
#831800000000
0!
0%
b110 *
0-
02
b110 6
#831810000000
1!
1%
1-
12
#831820000000
0!
0%
b111 *
0-
02
b111 6
#831830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#831840000000
0!
0%
b0 *
0-
02
b0 6
#831850000000
1!
1%
1-
12
#831860000000
0!
0%
b1 *
0-
02
b1 6
#831870000000
1!
1%
1-
12
#831880000000
0!
0%
b10 *
0-
02
b10 6
#831890000000
1!
1%
1-
12
#831900000000
0!
0%
b11 *
0-
02
b11 6
#831910000000
1!
1%
1-
12
15
#831920000000
0!
0%
b100 *
0-
02
b100 6
#831930000000
1!
1%
1-
12
#831940000000
0!
0%
b101 *
0-
02
b101 6
#831950000000
1!
1%
1-
12
#831960000000
0!
0%
b110 *
0-
02
b110 6
#831970000000
1!
1%
1-
12
#831980000000
0!
0%
b111 *
0-
02
b111 6
#831990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#832000000000
0!
0%
b0 *
0-
02
b0 6
#832010000000
1!
1%
1-
12
#832020000000
0!
0%
b1 *
0-
02
b1 6
#832030000000
1!
1%
1-
12
#832040000000
0!
0%
b10 *
0-
02
b10 6
#832050000000
1!
1%
1-
12
#832060000000
0!
0%
b11 *
0-
02
b11 6
#832070000000
1!
1%
1-
12
15
#832080000000
0!
0%
b100 *
0-
02
b100 6
#832090000000
1!
1%
1-
12
#832100000000
0!
0%
b101 *
0-
02
b101 6
#832110000000
1!
1%
1-
12
#832120000000
0!
0%
b110 *
0-
02
b110 6
#832130000000
1!
1%
1-
12
#832140000000
0!
0%
b111 *
0-
02
b111 6
#832150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#832160000000
0!
0%
b0 *
0-
02
b0 6
#832170000000
1!
1%
1-
12
#832180000000
0!
0%
b1 *
0-
02
b1 6
#832190000000
1!
1%
1-
12
#832200000000
0!
0%
b10 *
0-
02
b10 6
#832210000000
1!
1%
1-
12
#832220000000
0!
0%
b11 *
0-
02
b11 6
#832230000000
1!
1%
1-
12
15
#832240000000
0!
0%
b100 *
0-
02
b100 6
#832250000000
1!
1%
1-
12
#832260000000
0!
0%
b101 *
0-
02
b101 6
#832270000000
1!
1%
1-
12
#832280000000
0!
0%
b110 *
0-
02
b110 6
#832290000000
1!
1%
1-
12
#832300000000
0!
0%
b111 *
0-
02
b111 6
#832310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#832320000000
0!
0%
b0 *
0-
02
b0 6
#832330000000
1!
1%
1-
12
#832340000000
0!
0%
b1 *
0-
02
b1 6
#832350000000
1!
1%
1-
12
#832360000000
0!
0%
b10 *
0-
02
b10 6
#832370000000
1!
1%
1-
12
#832380000000
0!
0%
b11 *
0-
02
b11 6
#832390000000
1!
1%
1-
12
15
#832400000000
0!
0%
b100 *
0-
02
b100 6
#832410000000
1!
1%
1-
12
#832420000000
0!
0%
b101 *
0-
02
b101 6
#832430000000
1!
1%
1-
12
#832440000000
0!
0%
b110 *
0-
02
b110 6
#832450000000
1!
1%
1-
12
#832460000000
0!
0%
b111 *
0-
02
b111 6
#832470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#832480000000
0!
0%
b0 *
0-
02
b0 6
#832490000000
1!
1%
1-
12
#832500000000
0!
0%
b1 *
0-
02
b1 6
#832510000000
1!
1%
1-
12
#832520000000
0!
0%
b10 *
0-
02
b10 6
#832530000000
1!
1%
1-
12
#832540000000
0!
0%
b11 *
0-
02
b11 6
#832550000000
1!
1%
1-
12
15
#832560000000
0!
0%
b100 *
0-
02
b100 6
#832570000000
1!
1%
1-
12
#832580000000
0!
0%
b101 *
0-
02
b101 6
#832590000000
1!
1%
1-
12
#832600000000
0!
0%
b110 *
0-
02
b110 6
#832610000000
1!
1%
1-
12
#832620000000
0!
0%
b111 *
0-
02
b111 6
#832630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#832640000000
0!
0%
b0 *
0-
02
b0 6
#832650000000
1!
1%
1-
12
#832660000000
0!
0%
b1 *
0-
02
b1 6
#832670000000
1!
1%
1-
12
#832680000000
0!
0%
b10 *
0-
02
b10 6
#832690000000
1!
1%
1-
12
#832700000000
0!
0%
b11 *
0-
02
b11 6
#832710000000
1!
1%
1-
12
15
#832720000000
0!
0%
b100 *
0-
02
b100 6
#832730000000
1!
1%
1-
12
#832740000000
0!
0%
b101 *
0-
02
b101 6
#832750000000
1!
1%
1-
12
#832760000000
0!
0%
b110 *
0-
02
b110 6
#832770000000
1!
1%
1-
12
#832780000000
0!
0%
b111 *
0-
02
b111 6
#832790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#832800000000
0!
0%
b0 *
0-
02
b0 6
#832810000000
1!
1%
1-
12
#832820000000
0!
0%
b1 *
0-
02
b1 6
#832830000000
1!
1%
1-
12
#832840000000
0!
0%
b10 *
0-
02
b10 6
#832850000000
1!
1%
1-
12
#832860000000
0!
0%
b11 *
0-
02
b11 6
#832870000000
1!
1%
1-
12
15
#832880000000
0!
0%
b100 *
0-
02
b100 6
#832890000000
1!
1%
1-
12
#832900000000
0!
0%
b101 *
0-
02
b101 6
#832910000000
1!
1%
1-
12
#832920000000
0!
0%
b110 *
0-
02
b110 6
#832930000000
1!
1%
1-
12
#832940000000
0!
0%
b111 *
0-
02
b111 6
#832950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#832960000000
0!
0%
b0 *
0-
02
b0 6
#832970000000
1!
1%
1-
12
#832980000000
0!
0%
b1 *
0-
02
b1 6
#832990000000
1!
1%
1-
12
#833000000000
0!
0%
b10 *
0-
02
b10 6
#833010000000
1!
1%
1-
12
#833020000000
0!
0%
b11 *
0-
02
b11 6
#833030000000
1!
1%
1-
12
15
#833040000000
0!
0%
b100 *
0-
02
b100 6
#833050000000
1!
1%
1-
12
#833060000000
0!
0%
b101 *
0-
02
b101 6
#833070000000
1!
1%
1-
12
#833080000000
0!
0%
b110 *
0-
02
b110 6
#833090000000
1!
1%
1-
12
#833100000000
0!
0%
b111 *
0-
02
b111 6
#833110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#833120000000
0!
0%
b0 *
0-
02
b0 6
#833130000000
1!
1%
1-
12
#833140000000
0!
0%
b1 *
0-
02
b1 6
#833150000000
1!
1%
1-
12
#833160000000
0!
0%
b10 *
0-
02
b10 6
#833170000000
1!
1%
1-
12
#833180000000
0!
0%
b11 *
0-
02
b11 6
#833190000000
1!
1%
1-
12
15
#833200000000
0!
0%
b100 *
0-
02
b100 6
#833210000000
1!
1%
1-
12
#833220000000
0!
0%
b101 *
0-
02
b101 6
#833230000000
1!
1%
1-
12
#833240000000
0!
0%
b110 *
0-
02
b110 6
#833250000000
1!
1%
1-
12
#833260000000
0!
0%
b111 *
0-
02
b111 6
#833270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#833280000000
0!
0%
b0 *
0-
02
b0 6
#833290000000
1!
1%
1-
12
#833300000000
0!
0%
b1 *
0-
02
b1 6
#833310000000
1!
1%
1-
12
#833320000000
0!
0%
b10 *
0-
02
b10 6
#833330000000
1!
1%
1-
12
#833340000000
0!
0%
b11 *
0-
02
b11 6
#833350000000
1!
1%
1-
12
15
#833360000000
0!
0%
b100 *
0-
02
b100 6
#833370000000
1!
1%
1-
12
#833380000000
0!
0%
b101 *
0-
02
b101 6
#833390000000
1!
1%
1-
12
#833400000000
0!
0%
b110 *
0-
02
b110 6
#833410000000
1!
1%
1-
12
#833420000000
0!
0%
b111 *
0-
02
b111 6
#833430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#833440000000
0!
0%
b0 *
0-
02
b0 6
#833450000000
1!
1%
1-
12
#833460000000
0!
0%
b1 *
0-
02
b1 6
#833470000000
1!
1%
1-
12
#833480000000
0!
0%
b10 *
0-
02
b10 6
#833490000000
1!
1%
1-
12
#833500000000
0!
0%
b11 *
0-
02
b11 6
#833510000000
1!
1%
1-
12
15
#833520000000
0!
0%
b100 *
0-
02
b100 6
#833530000000
1!
1%
1-
12
#833540000000
0!
0%
b101 *
0-
02
b101 6
#833550000000
1!
1%
1-
12
#833560000000
0!
0%
b110 *
0-
02
b110 6
#833570000000
1!
1%
1-
12
#833580000000
0!
0%
b111 *
0-
02
b111 6
#833590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#833600000000
0!
0%
b0 *
0-
02
b0 6
#833610000000
1!
1%
1-
12
#833620000000
0!
0%
b1 *
0-
02
b1 6
#833630000000
1!
1%
1-
12
#833640000000
0!
0%
b10 *
0-
02
b10 6
#833650000000
1!
1%
1-
12
#833660000000
0!
0%
b11 *
0-
02
b11 6
#833670000000
1!
1%
1-
12
15
#833680000000
0!
0%
b100 *
0-
02
b100 6
#833690000000
1!
1%
1-
12
#833700000000
0!
0%
b101 *
0-
02
b101 6
#833710000000
1!
1%
1-
12
#833720000000
0!
0%
b110 *
0-
02
b110 6
#833730000000
1!
1%
1-
12
#833740000000
0!
0%
b111 *
0-
02
b111 6
#833750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#833760000000
0!
0%
b0 *
0-
02
b0 6
#833770000000
1!
1%
1-
12
#833780000000
0!
0%
b1 *
0-
02
b1 6
#833790000000
1!
1%
1-
12
#833800000000
0!
0%
b10 *
0-
02
b10 6
#833810000000
1!
1%
1-
12
#833820000000
0!
0%
b11 *
0-
02
b11 6
#833830000000
1!
1%
1-
12
15
#833840000000
0!
0%
b100 *
0-
02
b100 6
#833850000000
1!
1%
1-
12
#833860000000
0!
0%
b101 *
0-
02
b101 6
#833870000000
1!
1%
1-
12
#833880000000
0!
0%
b110 *
0-
02
b110 6
#833890000000
1!
1%
1-
12
#833900000000
0!
0%
b111 *
0-
02
b111 6
#833910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#833920000000
0!
0%
b0 *
0-
02
b0 6
#833930000000
1!
1%
1-
12
#833940000000
0!
0%
b1 *
0-
02
b1 6
#833950000000
1!
1%
1-
12
#833960000000
0!
0%
b10 *
0-
02
b10 6
#833970000000
1!
1%
1-
12
#833980000000
0!
0%
b11 *
0-
02
b11 6
#833990000000
1!
1%
1-
12
15
#834000000000
0!
0%
b100 *
0-
02
b100 6
#834010000000
1!
1%
1-
12
#834020000000
0!
0%
b101 *
0-
02
b101 6
#834030000000
1!
1%
1-
12
#834040000000
0!
0%
b110 *
0-
02
b110 6
#834050000000
1!
1%
1-
12
#834060000000
0!
0%
b111 *
0-
02
b111 6
#834070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#834080000000
0!
0%
b0 *
0-
02
b0 6
#834090000000
1!
1%
1-
12
#834100000000
0!
0%
b1 *
0-
02
b1 6
#834110000000
1!
1%
1-
12
#834120000000
0!
0%
b10 *
0-
02
b10 6
#834130000000
1!
1%
1-
12
#834140000000
0!
0%
b11 *
0-
02
b11 6
#834150000000
1!
1%
1-
12
15
#834160000000
0!
0%
b100 *
0-
02
b100 6
#834170000000
1!
1%
1-
12
#834180000000
0!
0%
b101 *
0-
02
b101 6
#834190000000
1!
1%
1-
12
#834200000000
0!
0%
b110 *
0-
02
b110 6
#834210000000
1!
1%
1-
12
#834220000000
0!
0%
b111 *
0-
02
b111 6
#834230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#834240000000
0!
0%
b0 *
0-
02
b0 6
#834250000000
1!
1%
1-
12
#834260000000
0!
0%
b1 *
0-
02
b1 6
#834270000000
1!
1%
1-
12
#834280000000
0!
0%
b10 *
0-
02
b10 6
#834290000000
1!
1%
1-
12
#834300000000
0!
0%
b11 *
0-
02
b11 6
#834310000000
1!
1%
1-
12
15
#834320000000
0!
0%
b100 *
0-
02
b100 6
#834330000000
1!
1%
1-
12
#834340000000
0!
0%
b101 *
0-
02
b101 6
#834350000000
1!
1%
1-
12
#834360000000
0!
0%
b110 *
0-
02
b110 6
#834370000000
1!
1%
1-
12
#834380000000
0!
0%
b111 *
0-
02
b111 6
#834390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#834400000000
0!
0%
b0 *
0-
02
b0 6
#834410000000
1!
1%
1-
12
#834420000000
0!
0%
b1 *
0-
02
b1 6
#834430000000
1!
1%
1-
12
#834440000000
0!
0%
b10 *
0-
02
b10 6
#834450000000
1!
1%
1-
12
#834460000000
0!
0%
b11 *
0-
02
b11 6
#834470000000
1!
1%
1-
12
15
#834480000000
0!
0%
b100 *
0-
02
b100 6
#834490000000
1!
1%
1-
12
#834500000000
0!
0%
b101 *
0-
02
b101 6
#834510000000
1!
1%
1-
12
#834520000000
0!
0%
b110 *
0-
02
b110 6
#834530000000
1!
1%
1-
12
#834540000000
0!
0%
b111 *
0-
02
b111 6
#834550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#834560000000
0!
0%
b0 *
0-
02
b0 6
#834570000000
1!
1%
1-
12
#834580000000
0!
0%
b1 *
0-
02
b1 6
#834590000000
1!
1%
1-
12
#834600000000
0!
0%
b10 *
0-
02
b10 6
#834610000000
1!
1%
1-
12
#834620000000
0!
0%
b11 *
0-
02
b11 6
#834630000000
1!
1%
1-
12
15
#834640000000
0!
0%
b100 *
0-
02
b100 6
#834650000000
1!
1%
1-
12
#834660000000
0!
0%
b101 *
0-
02
b101 6
#834670000000
1!
1%
1-
12
#834680000000
0!
0%
b110 *
0-
02
b110 6
#834690000000
1!
1%
1-
12
#834700000000
0!
0%
b111 *
0-
02
b111 6
#834710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#834720000000
0!
0%
b0 *
0-
02
b0 6
#834730000000
1!
1%
1-
12
#834740000000
0!
0%
b1 *
0-
02
b1 6
#834750000000
1!
1%
1-
12
#834760000000
0!
0%
b10 *
0-
02
b10 6
#834770000000
1!
1%
1-
12
#834780000000
0!
0%
b11 *
0-
02
b11 6
#834790000000
1!
1%
1-
12
15
#834800000000
0!
0%
b100 *
0-
02
b100 6
#834810000000
1!
1%
1-
12
#834820000000
0!
0%
b101 *
0-
02
b101 6
#834830000000
1!
1%
1-
12
#834840000000
0!
0%
b110 *
0-
02
b110 6
#834850000000
1!
1%
1-
12
#834860000000
0!
0%
b111 *
0-
02
b111 6
#834870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#834880000000
0!
0%
b0 *
0-
02
b0 6
#834890000000
1!
1%
1-
12
#834900000000
0!
0%
b1 *
0-
02
b1 6
#834910000000
1!
1%
1-
12
#834920000000
0!
0%
b10 *
0-
02
b10 6
#834930000000
1!
1%
1-
12
#834940000000
0!
0%
b11 *
0-
02
b11 6
#834950000000
1!
1%
1-
12
15
#834960000000
0!
0%
b100 *
0-
02
b100 6
#834970000000
1!
1%
1-
12
#834980000000
0!
0%
b101 *
0-
02
b101 6
#834990000000
1!
1%
1-
12
#835000000000
0!
0%
b110 *
0-
02
b110 6
#835010000000
1!
1%
1-
12
#835020000000
0!
0%
b111 *
0-
02
b111 6
#835030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#835040000000
0!
0%
b0 *
0-
02
b0 6
#835050000000
1!
1%
1-
12
#835060000000
0!
0%
b1 *
0-
02
b1 6
#835070000000
1!
1%
1-
12
#835080000000
0!
0%
b10 *
0-
02
b10 6
#835090000000
1!
1%
1-
12
#835100000000
0!
0%
b11 *
0-
02
b11 6
#835110000000
1!
1%
1-
12
15
#835120000000
0!
0%
b100 *
0-
02
b100 6
#835130000000
1!
1%
1-
12
#835140000000
0!
0%
b101 *
0-
02
b101 6
#835150000000
1!
1%
1-
12
#835160000000
0!
0%
b110 *
0-
02
b110 6
#835170000000
1!
1%
1-
12
#835180000000
0!
0%
b111 *
0-
02
b111 6
#835190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#835200000000
0!
0%
b0 *
0-
02
b0 6
#835210000000
1!
1%
1-
12
#835220000000
0!
0%
b1 *
0-
02
b1 6
#835230000000
1!
1%
1-
12
#835240000000
0!
0%
b10 *
0-
02
b10 6
#835250000000
1!
1%
1-
12
#835260000000
0!
0%
b11 *
0-
02
b11 6
#835270000000
1!
1%
1-
12
15
#835280000000
0!
0%
b100 *
0-
02
b100 6
#835290000000
1!
1%
1-
12
#835300000000
0!
0%
b101 *
0-
02
b101 6
#835310000000
1!
1%
1-
12
#835320000000
0!
0%
b110 *
0-
02
b110 6
#835330000000
1!
1%
1-
12
#835340000000
0!
0%
b111 *
0-
02
b111 6
#835350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#835360000000
0!
0%
b0 *
0-
02
b0 6
#835370000000
1!
1%
1-
12
#835380000000
0!
0%
b1 *
0-
02
b1 6
#835390000000
1!
1%
1-
12
#835400000000
0!
0%
b10 *
0-
02
b10 6
#835410000000
1!
1%
1-
12
#835420000000
0!
0%
b11 *
0-
02
b11 6
#835430000000
1!
1%
1-
12
15
#835440000000
0!
0%
b100 *
0-
02
b100 6
#835450000000
1!
1%
1-
12
#835460000000
0!
0%
b101 *
0-
02
b101 6
#835470000000
1!
1%
1-
12
#835480000000
0!
0%
b110 *
0-
02
b110 6
#835490000000
1!
1%
1-
12
#835500000000
0!
0%
b111 *
0-
02
b111 6
#835510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#835520000000
0!
0%
b0 *
0-
02
b0 6
#835530000000
1!
1%
1-
12
#835540000000
0!
0%
b1 *
0-
02
b1 6
#835550000000
1!
1%
1-
12
#835560000000
0!
0%
b10 *
0-
02
b10 6
#835570000000
1!
1%
1-
12
#835580000000
0!
0%
b11 *
0-
02
b11 6
#835590000000
1!
1%
1-
12
15
#835600000000
0!
0%
b100 *
0-
02
b100 6
#835610000000
1!
1%
1-
12
#835620000000
0!
0%
b101 *
0-
02
b101 6
#835630000000
1!
1%
1-
12
#835640000000
0!
0%
b110 *
0-
02
b110 6
#835650000000
1!
1%
1-
12
#835660000000
0!
0%
b111 *
0-
02
b111 6
#835670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#835680000000
0!
0%
b0 *
0-
02
b0 6
#835690000000
1!
1%
1-
12
#835700000000
0!
0%
b1 *
0-
02
b1 6
#835710000000
1!
1%
1-
12
#835720000000
0!
0%
b10 *
0-
02
b10 6
#835730000000
1!
1%
1-
12
#835740000000
0!
0%
b11 *
0-
02
b11 6
#835750000000
1!
1%
1-
12
15
#835760000000
0!
0%
b100 *
0-
02
b100 6
#835770000000
1!
1%
1-
12
#835780000000
0!
0%
b101 *
0-
02
b101 6
#835790000000
1!
1%
1-
12
#835800000000
0!
0%
b110 *
0-
02
b110 6
#835810000000
1!
1%
1-
12
#835820000000
0!
0%
b111 *
0-
02
b111 6
#835830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#835840000000
0!
0%
b0 *
0-
02
b0 6
#835850000000
1!
1%
1-
12
#835860000000
0!
0%
b1 *
0-
02
b1 6
#835870000000
1!
1%
1-
12
#835880000000
0!
0%
b10 *
0-
02
b10 6
#835890000000
1!
1%
1-
12
#835900000000
0!
0%
b11 *
0-
02
b11 6
#835910000000
1!
1%
1-
12
15
#835920000000
0!
0%
b100 *
0-
02
b100 6
#835930000000
1!
1%
1-
12
#835940000000
0!
0%
b101 *
0-
02
b101 6
#835950000000
1!
1%
1-
12
#835960000000
0!
0%
b110 *
0-
02
b110 6
#835970000000
1!
1%
1-
12
#835980000000
0!
0%
b111 *
0-
02
b111 6
#835990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#836000000000
0!
0%
b0 *
0-
02
b0 6
#836010000000
1!
1%
1-
12
#836020000000
0!
0%
b1 *
0-
02
b1 6
#836030000000
1!
1%
1-
12
#836040000000
0!
0%
b10 *
0-
02
b10 6
#836050000000
1!
1%
1-
12
#836060000000
0!
0%
b11 *
0-
02
b11 6
#836070000000
1!
1%
1-
12
15
#836080000000
0!
0%
b100 *
0-
02
b100 6
#836090000000
1!
1%
1-
12
#836100000000
0!
0%
b101 *
0-
02
b101 6
#836110000000
1!
1%
1-
12
#836120000000
0!
0%
b110 *
0-
02
b110 6
#836130000000
1!
1%
1-
12
#836140000000
0!
0%
b111 *
0-
02
b111 6
#836150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#836160000000
0!
0%
b0 *
0-
02
b0 6
#836170000000
1!
1%
1-
12
#836180000000
0!
0%
b1 *
0-
02
b1 6
#836190000000
1!
1%
1-
12
#836200000000
0!
0%
b10 *
0-
02
b10 6
#836210000000
1!
1%
1-
12
#836220000000
0!
0%
b11 *
0-
02
b11 6
#836230000000
1!
1%
1-
12
15
#836240000000
0!
0%
b100 *
0-
02
b100 6
#836250000000
1!
1%
1-
12
#836260000000
0!
0%
b101 *
0-
02
b101 6
#836270000000
1!
1%
1-
12
#836280000000
0!
0%
b110 *
0-
02
b110 6
#836290000000
1!
1%
1-
12
#836300000000
0!
0%
b111 *
0-
02
b111 6
#836310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#836320000000
0!
0%
b0 *
0-
02
b0 6
#836330000000
1!
1%
1-
12
#836340000000
0!
0%
b1 *
0-
02
b1 6
#836350000000
1!
1%
1-
12
#836360000000
0!
0%
b10 *
0-
02
b10 6
#836370000000
1!
1%
1-
12
#836380000000
0!
0%
b11 *
0-
02
b11 6
#836390000000
1!
1%
1-
12
15
#836400000000
0!
0%
b100 *
0-
02
b100 6
#836410000000
1!
1%
1-
12
#836420000000
0!
0%
b101 *
0-
02
b101 6
#836430000000
1!
1%
1-
12
#836440000000
0!
0%
b110 *
0-
02
b110 6
#836450000000
1!
1%
1-
12
#836460000000
0!
0%
b111 *
0-
02
b111 6
#836470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#836480000000
0!
0%
b0 *
0-
02
b0 6
#836490000000
1!
1%
1-
12
#836500000000
0!
0%
b1 *
0-
02
b1 6
#836510000000
1!
1%
1-
12
#836520000000
0!
0%
b10 *
0-
02
b10 6
#836530000000
1!
1%
1-
12
#836540000000
0!
0%
b11 *
0-
02
b11 6
#836550000000
1!
1%
1-
12
15
#836560000000
0!
0%
b100 *
0-
02
b100 6
#836570000000
1!
1%
1-
12
#836580000000
0!
0%
b101 *
0-
02
b101 6
#836590000000
1!
1%
1-
12
#836600000000
0!
0%
b110 *
0-
02
b110 6
#836610000000
1!
1%
1-
12
#836620000000
0!
0%
b111 *
0-
02
b111 6
#836630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#836640000000
0!
0%
b0 *
0-
02
b0 6
#836650000000
1!
1%
1-
12
#836660000000
0!
0%
b1 *
0-
02
b1 6
#836670000000
1!
1%
1-
12
#836680000000
0!
0%
b10 *
0-
02
b10 6
#836690000000
1!
1%
1-
12
#836700000000
0!
0%
b11 *
0-
02
b11 6
#836710000000
1!
1%
1-
12
15
#836720000000
0!
0%
b100 *
0-
02
b100 6
#836730000000
1!
1%
1-
12
#836740000000
0!
0%
b101 *
0-
02
b101 6
#836750000000
1!
1%
1-
12
#836760000000
0!
0%
b110 *
0-
02
b110 6
#836770000000
1!
1%
1-
12
#836780000000
0!
0%
b111 *
0-
02
b111 6
#836790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#836800000000
0!
0%
b0 *
0-
02
b0 6
#836810000000
1!
1%
1-
12
#836820000000
0!
0%
b1 *
0-
02
b1 6
#836830000000
1!
1%
1-
12
#836840000000
0!
0%
b10 *
0-
02
b10 6
#836850000000
1!
1%
1-
12
#836860000000
0!
0%
b11 *
0-
02
b11 6
#836870000000
1!
1%
1-
12
15
#836880000000
0!
0%
b100 *
0-
02
b100 6
#836890000000
1!
1%
1-
12
#836900000000
0!
0%
b101 *
0-
02
b101 6
#836910000000
1!
1%
1-
12
#836920000000
0!
0%
b110 *
0-
02
b110 6
#836930000000
1!
1%
1-
12
#836940000000
0!
0%
b111 *
0-
02
b111 6
#836950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#836960000000
0!
0%
b0 *
0-
02
b0 6
#836970000000
1!
1%
1-
12
#836980000000
0!
0%
b1 *
0-
02
b1 6
#836990000000
1!
1%
1-
12
#837000000000
0!
0%
b10 *
0-
02
b10 6
#837010000000
1!
1%
1-
12
#837020000000
0!
0%
b11 *
0-
02
b11 6
#837030000000
1!
1%
1-
12
15
#837040000000
0!
0%
b100 *
0-
02
b100 6
#837050000000
1!
1%
1-
12
#837060000000
0!
0%
b101 *
0-
02
b101 6
#837070000000
1!
1%
1-
12
#837080000000
0!
0%
b110 *
0-
02
b110 6
#837090000000
1!
1%
1-
12
#837100000000
0!
0%
b111 *
0-
02
b111 6
#837110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#837120000000
0!
0%
b0 *
0-
02
b0 6
#837130000000
1!
1%
1-
12
#837140000000
0!
0%
b1 *
0-
02
b1 6
#837150000000
1!
1%
1-
12
#837160000000
0!
0%
b10 *
0-
02
b10 6
#837170000000
1!
1%
1-
12
#837180000000
0!
0%
b11 *
0-
02
b11 6
#837190000000
1!
1%
1-
12
15
#837200000000
0!
0%
b100 *
0-
02
b100 6
#837210000000
1!
1%
1-
12
#837220000000
0!
0%
b101 *
0-
02
b101 6
#837230000000
1!
1%
1-
12
#837240000000
0!
0%
b110 *
0-
02
b110 6
#837250000000
1!
1%
1-
12
#837260000000
0!
0%
b111 *
0-
02
b111 6
#837270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#837280000000
0!
0%
b0 *
0-
02
b0 6
#837290000000
1!
1%
1-
12
#837300000000
0!
0%
b1 *
0-
02
b1 6
#837310000000
1!
1%
1-
12
#837320000000
0!
0%
b10 *
0-
02
b10 6
#837330000000
1!
1%
1-
12
#837340000000
0!
0%
b11 *
0-
02
b11 6
#837350000000
1!
1%
1-
12
15
#837360000000
0!
0%
b100 *
0-
02
b100 6
#837370000000
1!
1%
1-
12
#837380000000
0!
0%
b101 *
0-
02
b101 6
#837390000000
1!
1%
1-
12
#837400000000
0!
0%
b110 *
0-
02
b110 6
#837410000000
1!
1%
1-
12
#837420000000
0!
0%
b111 *
0-
02
b111 6
#837430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#837440000000
0!
0%
b0 *
0-
02
b0 6
#837450000000
1!
1%
1-
12
#837460000000
0!
0%
b1 *
0-
02
b1 6
#837470000000
1!
1%
1-
12
#837480000000
0!
0%
b10 *
0-
02
b10 6
#837490000000
1!
1%
1-
12
#837500000000
0!
0%
b11 *
0-
02
b11 6
#837510000000
1!
1%
1-
12
15
#837520000000
0!
0%
b100 *
0-
02
b100 6
#837530000000
1!
1%
1-
12
#837540000000
0!
0%
b101 *
0-
02
b101 6
#837550000000
1!
1%
1-
12
#837560000000
0!
0%
b110 *
0-
02
b110 6
#837570000000
1!
1%
1-
12
#837580000000
0!
0%
b111 *
0-
02
b111 6
#837590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#837600000000
0!
0%
b0 *
0-
02
b0 6
#837610000000
1!
1%
1-
12
#837620000000
0!
0%
b1 *
0-
02
b1 6
#837630000000
1!
1%
1-
12
#837640000000
0!
0%
b10 *
0-
02
b10 6
#837650000000
1!
1%
1-
12
#837660000000
0!
0%
b11 *
0-
02
b11 6
#837670000000
1!
1%
1-
12
15
#837680000000
0!
0%
b100 *
0-
02
b100 6
#837690000000
1!
1%
1-
12
#837700000000
0!
0%
b101 *
0-
02
b101 6
#837710000000
1!
1%
1-
12
#837720000000
0!
0%
b110 *
0-
02
b110 6
#837730000000
1!
1%
1-
12
#837740000000
0!
0%
b111 *
0-
02
b111 6
#837750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#837760000000
0!
0%
b0 *
0-
02
b0 6
#837770000000
1!
1%
1-
12
#837780000000
0!
0%
b1 *
0-
02
b1 6
#837790000000
1!
1%
1-
12
#837800000000
0!
0%
b10 *
0-
02
b10 6
#837810000000
1!
1%
1-
12
#837820000000
0!
0%
b11 *
0-
02
b11 6
#837830000000
1!
1%
1-
12
15
#837840000000
0!
0%
b100 *
0-
02
b100 6
#837850000000
1!
1%
1-
12
#837860000000
0!
0%
b101 *
0-
02
b101 6
#837870000000
1!
1%
1-
12
#837880000000
0!
0%
b110 *
0-
02
b110 6
#837890000000
1!
1%
1-
12
#837900000000
0!
0%
b111 *
0-
02
b111 6
#837910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#837920000000
0!
0%
b0 *
0-
02
b0 6
#837930000000
1!
1%
1-
12
#837940000000
0!
0%
b1 *
0-
02
b1 6
#837950000000
1!
1%
1-
12
#837960000000
0!
0%
b10 *
0-
02
b10 6
#837970000000
1!
1%
1-
12
#837980000000
0!
0%
b11 *
0-
02
b11 6
#837990000000
1!
1%
1-
12
15
#838000000000
0!
0%
b100 *
0-
02
b100 6
#838010000000
1!
1%
1-
12
#838020000000
0!
0%
b101 *
0-
02
b101 6
#838030000000
1!
1%
1-
12
#838040000000
0!
0%
b110 *
0-
02
b110 6
#838050000000
1!
1%
1-
12
#838060000000
0!
0%
b111 *
0-
02
b111 6
#838070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#838080000000
0!
0%
b0 *
0-
02
b0 6
#838090000000
1!
1%
1-
12
#838100000000
0!
0%
b1 *
0-
02
b1 6
#838110000000
1!
1%
1-
12
#838120000000
0!
0%
b10 *
0-
02
b10 6
#838130000000
1!
1%
1-
12
#838140000000
0!
0%
b11 *
0-
02
b11 6
#838150000000
1!
1%
1-
12
15
#838160000000
0!
0%
b100 *
0-
02
b100 6
#838170000000
1!
1%
1-
12
#838180000000
0!
0%
b101 *
0-
02
b101 6
#838190000000
1!
1%
1-
12
#838200000000
0!
0%
b110 *
0-
02
b110 6
#838210000000
1!
1%
1-
12
#838220000000
0!
0%
b111 *
0-
02
b111 6
#838230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#838240000000
0!
0%
b0 *
0-
02
b0 6
#838250000000
1!
1%
1-
12
#838260000000
0!
0%
b1 *
0-
02
b1 6
#838270000000
1!
1%
1-
12
#838280000000
0!
0%
b10 *
0-
02
b10 6
#838290000000
1!
1%
1-
12
#838300000000
0!
0%
b11 *
0-
02
b11 6
#838310000000
1!
1%
1-
12
15
#838320000000
0!
0%
b100 *
0-
02
b100 6
#838330000000
1!
1%
1-
12
#838340000000
0!
0%
b101 *
0-
02
b101 6
#838350000000
1!
1%
1-
12
#838360000000
0!
0%
b110 *
0-
02
b110 6
#838370000000
1!
1%
1-
12
#838380000000
0!
0%
b111 *
0-
02
b111 6
#838390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#838400000000
0!
0%
b0 *
0-
02
b0 6
#838410000000
1!
1%
1-
12
#838420000000
0!
0%
b1 *
0-
02
b1 6
#838430000000
1!
1%
1-
12
#838440000000
0!
0%
b10 *
0-
02
b10 6
#838450000000
1!
1%
1-
12
#838460000000
0!
0%
b11 *
0-
02
b11 6
#838470000000
1!
1%
1-
12
15
#838480000000
0!
0%
b100 *
0-
02
b100 6
#838490000000
1!
1%
1-
12
#838500000000
0!
0%
b101 *
0-
02
b101 6
#838510000000
1!
1%
1-
12
#838520000000
0!
0%
b110 *
0-
02
b110 6
#838530000000
1!
1%
1-
12
#838540000000
0!
0%
b111 *
0-
02
b111 6
#838550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#838560000000
0!
0%
b0 *
0-
02
b0 6
#838570000000
1!
1%
1-
12
#838580000000
0!
0%
b1 *
0-
02
b1 6
#838590000000
1!
1%
1-
12
#838600000000
0!
0%
b10 *
0-
02
b10 6
#838610000000
1!
1%
1-
12
#838620000000
0!
0%
b11 *
0-
02
b11 6
#838630000000
1!
1%
1-
12
15
#838640000000
0!
0%
b100 *
0-
02
b100 6
#838650000000
1!
1%
1-
12
#838660000000
0!
0%
b101 *
0-
02
b101 6
#838670000000
1!
1%
1-
12
#838680000000
0!
0%
b110 *
0-
02
b110 6
#838690000000
1!
1%
1-
12
#838700000000
0!
0%
b111 *
0-
02
b111 6
#838710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#838720000000
0!
0%
b0 *
0-
02
b0 6
#838730000000
1!
1%
1-
12
#838740000000
0!
0%
b1 *
0-
02
b1 6
#838750000000
1!
1%
1-
12
#838760000000
0!
0%
b10 *
0-
02
b10 6
#838770000000
1!
1%
1-
12
#838780000000
0!
0%
b11 *
0-
02
b11 6
#838790000000
1!
1%
1-
12
15
#838800000000
0!
0%
b100 *
0-
02
b100 6
#838810000000
1!
1%
1-
12
#838820000000
0!
0%
b101 *
0-
02
b101 6
#838830000000
1!
1%
1-
12
#838840000000
0!
0%
b110 *
0-
02
b110 6
#838850000000
1!
1%
1-
12
#838860000000
0!
0%
b111 *
0-
02
b111 6
#838870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#838880000000
0!
0%
b0 *
0-
02
b0 6
#838890000000
1!
1%
1-
12
#838900000000
0!
0%
b1 *
0-
02
b1 6
#838910000000
1!
1%
1-
12
#838920000000
0!
0%
b10 *
0-
02
b10 6
#838930000000
1!
1%
1-
12
#838940000000
0!
0%
b11 *
0-
02
b11 6
#838950000000
1!
1%
1-
12
15
#838960000000
0!
0%
b100 *
0-
02
b100 6
#838970000000
1!
1%
1-
12
#838980000000
0!
0%
b101 *
0-
02
b101 6
#838990000000
1!
1%
1-
12
#839000000000
0!
0%
b110 *
0-
02
b110 6
#839010000000
1!
1%
1-
12
#839020000000
0!
0%
b111 *
0-
02
b111 6
#839030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#839040000000
0!
0%
b0 *
0-
02
b0 6
#839050000000
1!
1%
1-
12
#839060000000
0!
0%
b1 *
0-
02
b1 6
#839070000000
1!
1%
1-
12
#839080000000
0!
0%
b10 *
0-
02
b10 6
#839090000000
1!
1%
1-
12
#839100000000
0!
0%
b11 *
0-
02
b11 6
#839110000000
1!
1%
1-
12
15
#839120000000
0!
0%
b100 *
0-
02
b100 6
#839130000000
1!
1%
1-
12
#839140000000
0!
0%
b101 *
0-
02
b101 6
#839150000000
1!
1%
1-
12
#839160000000
0!
0%
b110 *
0-
02
b110 6
#839170000000
1!
1%
1-
12
#839180000000
0!
0%
b111 *
0-
02
b111 6
#839190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#839200000000
0!
0%
b0 *
0-
02
b0 6
#839210000000
1!
1%
1-
12
#839220000000
0!
0%
b1 *
0-
02
b1 6
#839230000000
1!
1%
1-
12
#839240000000
0!
0%
b10 *
0-
02
b10 6
#839250000000
1!
1%
1-
12
#839260000000
0!
0%
b11 *
0-
02
b11 6
#839270000000
1!
1%
1-
12
15
#839280000000
0!
0%
b100 *
0-
02
b100 6
#839290000000
1!
1%
1-
12
#839300000000
0!
0%
b101 *
0-
02
b101 6
#839310000000
1!
1%
1-
12
#839320000000
0!
0%
b110 *
0-
02
b110 6
#839330000000
1!
1%
1-
12
#839340000000
0!
0%
b111 *
0-
02
b111 6
#839350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#839360000000
0!
0%
b0 *
0-
02
b0 6
#839370000000
1!
1%
1-
12
#839380000000
0!
0%
b1 *
0-
02
b1 6
#839390000000
1!
1%
1-
12
#839400000000
0!
0%
b10 *
0-
02
b10 6
#839410000000
1!
1%
1-
12
#839420000000
0!
0%
b11 *
0-
02
b11 6
#839430000000
1!
1%
1-
12
15
#839440000000
0!
0%
b100 *
0-
02
b100 6
#839450000000
1!
1%
1-
12
#839460000000
0!
0%
b101 *
0-
02
b101 6
#839470000000
1!
1%
1-
12
#839480000000
0!
0%
b110 *
0-
02
b110 6
#839490000000
1!
1%
1-
12
#839500000000
0!
0%
b111 *
0-
02
b111 6
#839510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#839520000000
0!
0%
b0 *
0-
02
b0 6
#839530000000
1!
1%
1-
12
#839540000000
0!
0%
b1 *
0-
02
b1 6
#839550000000
1!
1%
1-
12
#839560000000
0!
0%
b10 *
0-
02
b10 6
#839570000000
1!
1%
1-
12
#839580000000
0!
0%
b11 *
0-
02
b11 6
#839590000000
1!
1%
1-
12
15
#839600000000
0!
0%
b100 *
0-
02
b100 6
#839610000000
1!
1%
1-
12
#839620000000
0!
0%
b101 *
0-
02
b101 6
#839630000000
1!
1%
1-
12
#839640000000
0!
0%
b110 *
0-
02
b110 6
#839650000000
1!
1%
1-
12
#839660000000
0!
0%
b111 *
0-
02
b111 6
#839670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#839680000000
0!
0%
b0 *
0-
02
b0 6
#839690000000
1!
1%
1-
12
#839700000000
0!
0%
b1 *
0-
02
b1 6
#839710000000
1!
1%
1-
12
#839720000000
0!
0%
b10 *
0-
02
b10 6
#839730000000
1!
1%
1-
12
#839740000000
0!
0%
b11 *
0-
02
b11 6
#839750000000
1!
1%
1-
12
15
#839760000000
0!
0%
b100 *
0-
02
b100 6
#839770000000
1!
1%
1-
12
#839780000000
0!
0%
b101 *
0-
02
b101 6
#839790000000
1!
1%
1-
12
#839800000000
0!
0%
b110 *
0-
02
b110 6
#839810000000
1!
1%
1-
12
#839820000000
0!
0%
b111 *
0-
02
b111 6
#839830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#839840000000
0!
0%
b0 *
0-
02
b0 6
#839850000000
1!
1%
1-
12
#839860000000
0!
0%
b1 *
0-
02
b1 6
#839870000000
1!
1%
1-
12
#839880000000
0!
0%
b10 *
0-
02
b10 6
#839890000000
1!
1%
1-
12
#839900000000
0!
0%
b11 *
0-
02
b11 6
#839910000000
1!
1%
1-
12
15
#839920000000
0!
0%
b100 *
0-
02
b100 6
#839930000000
1!
1%
1-
12
#839940000000
0!
0%
b101 *
0-
02
b101 6
#839950000000
1!
1%
1-
12
#839960000000
0!
0%
b110 *
0-
02
b110 6
#839970000000
1!
1%
1-
12
#839980000000
0!
0%
b111 *
0-
02
b111 6
#839990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#840000000000
0!
0%
b0 *
0-
02
b0 6
#840010000000
1!
1%
1-
12
#840020000000
0!
0%
b1 *
0-
02
b1 6
#840030000000
1!
1%
1-
12
#840040000000
0!
0%
b10 *
0-
02
b10 6
#840050000000
1!
1%
1-
12
#840060000000
0!
0%
b11 *
0-
02
b11 6
#840070000000
1!
1%
1-
12
15
#840080000000
0!
0%
b100 *
0-
02
b100 6
#840090000000
1!
1%
1-
12
#840100000000
0!
0%
b101 *
0-
02
b101 6
#840110000000
1!
1%
1-
12
#840120000000
0!
0%
b110 *
0-
02
b110 6
#840130000000
1!
1%
1-
12
#840140000000
0!
0%
b111 *
0-
02
b111 6
#840150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#840160000000
0!
0%
b0 *
0-
02
b0 6
#840170000000
1!
1%
1-
12
#840180000000
0!
0%
b1 *
0-
02
b1 6
#840190000000
1!
1%
1-
12
#840200000000
0!
0%
b10 *
0-
02
b10 6
#840210000000
1!
1%
1-
12
#840220000000
0!
0%
b11 *
0-
02
b11 6
#840230000000
1!
1%
1-
12
15
#840240000000
0!
0%
b100 *
0-
02
b100 6
#840250000000
1!
1%
1-
12
#840260000000
0!
0%
b101 *
0-
02
b101 6
#840270000000
1!
1%
1-
12
#840280000000
0!
0%
b110 *
0-
02
b110 6
#840290000000
1!
1%
1-
12
#840300000000
0!
0%
b111 *
0-
02
b111 6
#840310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#840320000000
0!
0%
b0 *
0-
02
b0 6
#840330000000
1!
1%
1-
12
#840340000000
0!
0%
b1 *
0-
02
b1 6
#840350000000
1!
1%
1-
12
#840360000000
0!
0%
b10 *
0-
02
b10 6
#840370000000
1!
1%
1-
12
#840380000000
0!
0%
b11 *
0-
02
b11 6
#840390000000
1!
1%
1-
12
15
#840400000000
0!
0%
b100 *
0-
02
b100 6
#840410000000
1!
1%
1-
12
#840420000000
0!
0%
b101 *
0-
02
b101 6
#840430000000
1!
1%
1-
12
#840440000000
0!
0%
b110 *
0-
02
b110 6
#840450000000
1!
1%
1-
12
#840460000000
0!
0%
b111 *
0-
02
b111 6
#840470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#840480000000
0!
0%
b0 *
0-
02
b0 6
#840490000000
1!
1%
1-
12
#840500000000
0!
0%
b1 *
0-
02
b1 6
#840510000000
1!
1%
1-
12
#840520000000
0!
0%
b10 *
0-
02
b10 6
#840530000000
1!
1%
1-
12
#840540000000
0!
0%
b11 *
0-
02
b11 6
#840550000000
1!
1%
1-
12
15
#840560000000
0!
0%
b100 *
0-
02
b100 6
#840570000000
1!
1%
1-
12
#840580000000
0!
0%
b101 *
0-
02
b101 6
#840590000000
1!
1%
1-
12
#840600000000
0!
0%
b110 *
0-
02
b110 6
#840610000000
1!
1%
1-
12
#840620000000
0!
0%
b111 *
0-
02
b111 6
#840630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#840640000000
0!
0%
b0 *
0-
02
b0 6
#840650000000
1!
1%
1-
12
#840660000000
0!
0%
b1 *
0-
02
b1 6
#840670000000
1!
1%
1-
12
#840680000000
0!
0%
b10 *
0-
02
b10 6
#840690000000
1!
1%
1-
12
#840700000000
0!
0%
b11 *
0-
02
b11 6
#840710000000
1!
1%
1-
12
15
#840720000000
0!
0%
b100 *
0-
02
b100 6
#840730000000
1!
1%
1-
12
#840740000000
0!
0%
b101 *
0-
02
b101 6
#840750000000
1!
1%
1-
12
#840760000000
0!
0%
b110 *
0-
02
b110 6
#840770000000
1!
1%
1-
12
#840780000000
0!
0%
b111 *
0-
02
b111 6
#840790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#840800000000
0!
0%
b0 *
0-
02
b0 6
#840810000000
1!
1%
1-
12
#840820000000
0!
0%
b1 *
0-
02
b1 6
#840830000000
1!
1%
1-
12
#840840000000
0!
0%
b10 *
0-
02
b10 6
#840850000000
1!
1%
1-
12
#840860000000
0!
0%
b11 *
0-
02
b11 6
#840870000000
1!
1%
1-
12
15
#840880000000
0!
0%
b100 *
0-
02
b100 6
#840890000000
1!
1%
1-
12
#840900000000
0!
0%
b101 *
0-
02
b101 6
#840910000000
1!
1%
1-
12
#840920000000
0!
0%
b110 *
0-
02
b110 6
#840930000000
1!
1%
1-
12
#840940000000
0!
0%
b111 *
0-
02
b111 6
#840950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#840960000000
0!
0%
b0 *
0-
02
b0 6
#840970000000
1!
1%
1-
12
#840980000000
0!
0%
b1 *
0-
02
b1 6
#840990000000
1!
1%
1-
12
#841000000000
0!
0%
b10 *
0-
02
b10 6
#841010000000
1!
1%
1-
12
#841020000000
0!
0%
b11 *
0-
02
b11 6
#841030000000
1!
1%
1-
12
15
#841040000000
0!
0%
b100 *
0-
02
b100 6
#841050000000
1!
1%
1-
12
#841060000000
0!
0%
b101 *
0-
02
b101 6
#841070000000
1!
1%
1-
12
#841080000000
0!
0%
b110 *
0-
02
b110 6
#841090000000
1!
1%
1-
12
#841100000000
0!
0%
b111 *
0-
02
b111 6
#841110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#841120000000
0!
0%
b0 *
0-
02
b0 6
#841130000000
1!
1%
1-
12
#841140000000
0!
0%
b1 *
0-
02
b1 6
#841150000000
1!
1%
1-
12
#841160000000
0!
0%
b10 *
0-
02
b10 6
#841170000000
1!
1%
1-
12
#841180000000
0!
0%
b11 *
0-
02
b11 6
#841190000000
1!
1%
1-
12
15
#841200000000
0!
0%
b100 *
0-
02
b100 6
#841210000000
1!
1%
1-
12
#841220000000
0!
0%
b101 *
0-
02
b101 6
#841230000000
1!
1%
1-
12
#841240000000
0!
0%
b110 *
0-
02
b110 6
#841250000000
1!
1%
1-
12
#841260000000
0!
0%
b111 *
0-
02
b111 6
#841270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#841280000000
0!
0%
b0 *
0-
02
b0 6
#841290000000
1!
1%
1-
12
#841300000000
0!
0%
b1 *
0-
02
b1 6
#841310000000
1!
1%
1-
12
#841320000000
0!
0%
b10 *
0-
02
b10 6
#841330000000
1!
1%
1-
12
#841340000000
0!
0%
b11 *
0-
02
b11 6
#841350000000
1!
1%
1-
12
15
#841360000000
0!
0%
b100 *
0-
02
b100 6
#841370000000
1!
1%
1-
12
#841380000000
0!
0%
b101 *
0-
02
b101 6
#841390000000
1!
1%
1-
12
#841400000000
0!
0%
b110 *
0-
02
b110 6
#841410000000
1!
1%
1-
12
#841420000000
0!
0%
b111 *
0-
02
b111 6
#841430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#841440000000
0!
0%
b0 *
0-
02
b0 6
#841450000000
1!
1%
1-
12
#841460000000
0!
0%
b1 *
0-
02
b1 6
#841470000000
1!
1%
1-
12
#841480000000
0!
0%
b10 *
0-
02
b10 6
#841490000000
1!
1%
1-
12
#841500000000
0!
0%
b11 *
0-
02
b11 6
#841510000000
1!
1%
1-
12
15
#841520000000
0!
0%
b100 *
0-
02
b100 6
#841530000000
1!
1%
1-
12
#841540000000
0!
0%
b101 *
0-
02
b101 6
#841550000000
1!
1%
1-
12
#841560000000
0!
0%
b110 *
0-
02
b110 6
#841570000000
1!
1%
1-
12
#841580000000
0!
0%
b111 *
0-
02
b111 6
#841590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#841600000000
0!
0%
b0 *
0-
02
b0 6
#841610000000
1!
1%
1-
12
#841620000000
0!
0%
b1 *
0-
02
b1 6
#841630000000
1!
1%
1-
12
#841640000000
0!
0%
b10 *
0-
02
b10 6
#841650000000
1!
1%
1-
12
#841660000000
0!
0%
b11 *
0-
02
b11 6
#841670000000
1!
1%
1-
12
15
#841680000000
0!
0%
b100 *
0-
02
b100 6
#841690000000
1!
1%
1-
12
#841700000000
0!
0%
b101 *
0-
02
b101 6
#841710000000
1!
1%
1-
12
#841720000000
0!
0%
b110 *
0-
02
b110 6
#841730000000
1!
1%
1-
12
#841740000000
0!
0%
b111 *
0-
02
b111 6
#841750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#841760000000
0!
0%
b0 *
0-
02
b0 6
#841770000000
1!
1%
1-
12
#841780000000
0!
0%
b1 *
0-
02
b1 6
#841790000000
1!
1%
1-
12
#841800000000
0!
0%
b10 *
0-
02
b10 6
#841810000000
1!
1%
1-
12
#841820000000
0!
0%
b11 *
0-
02
b11 6
#841830000000
1!
1%
1-
12
15
#841840000000
0!
0%
b100 *
0-
02
b100 6
#841850000000
1!
1%
1-
12
#841860000000
0!
0%
b101 *
0-
02
b101 6
#841870000000
1!
1%
1-
12
#841880000000
0!
0%
b110 *
0-
02
b110 6
#841890000000
1!
1%
1-
12
#841900000000
0!
0%
b111 *
0-
02
b111 6
#841910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#841920000000
0!
0%
b0 *
0-
02
b0 6
#841930000000
1!
1%
1-
12
#841940000000
0!
0%
b1 *
0-
02
b1 6
#841950000000
1!
1%
1-
12
#841960000000
0!
0%
b10 *
0-
02
b10 6
#841970000000
1!
1%
1-
12
#841980000000
0!
0%
b11 *
0-
02
b11 6
#841990000000
1!
1%
1-
12
15
#842000000000
0!
0%
b100 *
0-
02
b100 6
#842010000000
1!
1%
1-
12
#842020000000
0!
0%
b101 *
0-
02
b101 6
#842030000000
1!
1%
1-
12
#842040000000
0!
0%
b110 *
0-
02
b110 6
#842050000000
1!
1%
1-
12
#842060000000
0!
0%
b111 *
0-
02
b111 6
#842070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#842080000000
0!
0%
b0 *
0-
02
b0 6
#842090000000
1!
1%
1-
12
#842100000000
0!
0%
b1 *
0-
02
b1 6
#842110000000
1!
1%
1-
12
#842120000000
0!
0%
b10 *
0-
02
b10 6
#842130000000
1!
1%
1-
12
#842140000000
0!
0%
b11 *
0-
02
b11 6
#842150000000
1!
1%
1-
12
15
#842160000000
0!
0%
b100 *
0-
02
b100 6
#842170000000
1!
1%
1-
12
#842180000000
0!
0%
b101 *
0-
02
b101 6
#842190000000
1!
1%
1-
12
#842200000000
0!
0%
b110 *
0-
02
b110 6
#842210000000
1!
1%
1-
12
#842220000000
0!
0%
b111 *
0-
02
b111 6
#842230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#842240000000
0!
0%
b0 *
0-
02
b0 6
#842250000000
1!
1%
1-
12
#842260000000
0!
0%
b1 *
0-
02
b1 6
#842270000000
1!
1%
1-
12
#842280000000
0!
0%
b10 *
0-
02
b10 6
#842290000000
1!
1%
1-
12
#842300000000
0!
0%
b11 *
0-
02
b11 6
#842310000000
1!
1%
1-
12
15
#842320000000
0!
0%
b100 *
0-
02
b100 6
#842330000000
1!
1%
1-
12
#842340000000
0!
0%
b101 *
0-
02
b101 6
#842350000000
1!
1%
1-
12
#842360000000
0!
0%
b110 *
0-
02
b110 6
#842370000000
1!
1%
1-
12
#842380000000
0!
0%
b111 *
0-
02
b111 6
#842390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#842400000000
0!
0%
b0 *
0-
02
b0 6
#842410000000
1!
1%
1-
12
#842420000000
0!
0%
b1 *
0-
02
b1 6
#842430000000
1!
1%
1-
12
#842440000000
0!
0%
b10 *
0-
02
b10 6
#842450000000
1!
1%
1-
12
#842460000000
0!
0%
b11 *
0-
02
b11 6
#842470000000
1!
1%
1-
12
15
#842480000000
0!
0%
b100 *
0-
02
b100 6
#842490000000
1!
1%
1-
12
#842500000000
0!
0%
b101 *
0-
02
b101 6
#842510000000
1!
1%
1-
12
#842520000000
0!
0%
b110 *
0-
02
b110 6
#842530000000
1!
1%
1-
12
#842540000000
0!
0%
b111 *
0-
02
b111 6
#842550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#842560000000
0!
0%
b0 *
0-
02
b0 6
#842570000000
1!
1%
1-
12
#842580000000
0!
0%
b1 *
0-
02
b1 6
#842590000000
1!
1%
1-
12
#842600000000
0!
0%
b10 *
0-
02
b10 6
#842610000000
1!
1%
1-
12
#842620000000
0!
0%
b11 *
0-
02
b11 6
#842630000000
1!
1%
1-
12
15
#842640000000
0!
0%
b100 *
0-
02
b100 6
#842650000000
1!
1%
1-
12
#842660000000
0!
0%
b101 *
0-
02
b101 6
#842670000000
1!
1%
1-
12
#842680000000
0!
0%
b110 *
0-
02
b110 6
#842690000000
1!
1%
1-
12
#842700000000
0!
0%
b111 *
0-
02
b111 6
#842710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#842720000000
0!
0%
b0 *
0-
02
b0 6
#842730000000
1!
1%
1-
12
#842740000000
0!
0%
b1 *
0-
02
b1 6
#842750000000
1!
1%
1-
12
#842760000000
0!
0%
b10 *
0-
02
b10 6
#842770000000
1!
1%
1-
12
#842780000000
0!
0%
b11 *
0-
02
b11 6
#842790000000
1!
1%
1-
12
15
#842800000000
0!
0%
b100 *
0-
02
b100 6
#842810000000
1!
1%
1-
12
#842820000000
0!
0%
b101 *
0-
02
b101 6
#842830000000
1!
1%
1-
12
#842840000000
0!
0%
b110 *
0-
02
b110 6
#842850000000
1!
1%
1-
12
#842860000000
0!
0%
b111 *
0-
02
b111 6
#842870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#842880000000
0!
0%
b0 *
0-
02
b0 6
#842890000000
1!
1%
1-
12
#842900000000
0!
0%
b1 *
0-
02
b1 6
#842910000000
1!
1%
1-
12
#842920000000
0!
0%
b10 *
0-
02
b10 6
#842930000000
1!
1%
1-
12
#842940000000
0!
0%
b11 *
0-
02
b11 6
#842950000000
1!
1%
1-
12
15
#842960000000
0!
0%
b100 *
0-
02
b100 6
#842970000000
1!
1%
1-
12
#842980000000
0!
0%
b101 *
0-
02
b101 6
#842990000000
1!
1%
1-
12
#843000000000
0!
0%
b110 *
0-
02
b110 6
#843010000000
1!
1%
1-
12
#843020000000
0!
0%
b111 *
0-
02
b111 6
#843030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#843040000000
0!
0%
b0 *
0-
02
b0 6
#843050000000
1!
1%
1-
12
#843060000000
0!
0%
b1 *
0-
02
b1 6
#843070000000
1!
1%
1-
12
#843080000000
0!
0%
b10 *
0-
02
b10 6
#843090000000
1!
1%
1-
12
#843100000000
0!
0%
b11 *
0-
02
b11 6
#843110000000
1!
1%
1-
12
15
#843120000000
0!
0%
b100 *
0-
02
b100 6
#843130000000
1!
1%
1-
12
#843140000000
0!
0%
b101 *
0-
02
b101 6
#843150000000
1!
1%
1-
12
#843160000000
0!
0%
b110 *
0-
02
b110 6
#843170000000
1!
1%
1-
12
#843180000000
0!
0%
b111 *
0-
02
b111 6
#843190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#843200000000
0!
0%
b0 *
0-
02
b0 6
#843210000000
1!
1%
1-
12
#843220000000
0!
0%
b1 *
0-
02
b1 6
#843230000000
1!
1%
1-
12
#843240000000
0!
0%
b10 *
0-
02
b10 6
#843250000000
1!
1%
1-
12
#843260000000
0!
0%
b11 *
0-
02
b11 6
#843270000000
1!
1%
1-
12
15
#843280000000
0!
0%
b100 *
0-
02
b100 6
#843290000000
1!
1%
1-
12
#843300000000
0!
0%
b101 *
0-
02
b101 6
#843310000000
1!
1%
1-
12
#843320000000
0!
0%
b110 *
0-
02
b110 6
#843330000000
1!
1%
1-
12
#843340000000
0!
0%
b111 *
0-
02
b111 6
#843350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#843360000000
0!
0%
b0 *
0-
02
b0 6
#843370000000
1!
1%
1-
12
#843380000000
0!
0%
b1 *
0-
02
b1 6
#843390000000
1!
1%
1-
12
#843400000000
0!
0%
b10 *
0-
02
b10 6
#843410000000
1!
1%
1-
12
#843420000000
0!
0%
b11 *
0-
02
b11 6
#843430000000
1!
1%
1-
12
15
#843440000000
0!
0%
b100 *
0-
02
b100 6
#843450000000
1!
1%
1-
12
#843460000000
0!
0%
b101 *
0-
02
b101 6
#843470000000
1!
1%
1-
12
#843480000000
0!
0%
b110 *
0-
02
b110 6
#843490000000
1!
1%
1-
12
#843500000000
0!
0%
b111 *
0-
02
b111 6
#843510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#843520000000
0!
0%
b0 *
0-
02
b0 6
#843530000000
1!
1%
1-
12
#843540000000
0!
0%
b1 *
0-
02
b1 6
#843550000000
1!
1%
1-
12
#843560000000
0!
0%
b10 *
0-
02
b10 6
#843570000000
1!
1%
1-
12
#843580000000
0!
0%
b11 *
0-
02
b11 6
#843590000000
1!
1%
1-
12
15
#843600000000
0!
0%
b100 *
0-
02
b100 6
#843610000000
1!
1%
1-
12
#843620000000
0!
0%
b101 *
0-
02
b101 6
#843630000000
1!
1%
1-
12
#843640000000
0!
0%
b110 *
0-
02
b110 6
#843650000000
1!
1%
1-
12
#843660000000
0!
0%
b111 *
0-
02
b111 6
#843670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#843680000000
0!
0%
b0 *
0-
02
b0 6
#843690000000
1!
1%
1-
12
#843700000000
0!
0%
b1 *
0-
02
b1 6
#843710000000
1!
1%
1-
12
#843720000000
0!
0%
b10 *
0-
02
b10 6
#843730000000
1!
1%
1-
12
#843740000000
0!
0%
b11 *
0-
02
b11 6
#843750000000
1!
1%
1-
12
15
#843760000000
0!
0%
b100 *
0-
02
b100 6
#843770000000
1!
1%
1-
12
#843780000000
0!
0%
b101 *
0-
02
b101 6
#843790000000
1!
1%
1-
12
#843800000000
0!
0%
b110 *
0-
02
b110 6
#843810000000
1!
1%
1-
12
#843820000000
0!
0%
b111 *
0-
02
b111 6
#843830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#843840000000
0!
0%
b0 *
0-
02
b0 6
#843850000000
1!
1%
1-
12
#843860000000
0!
0%
b1 *
0-
02
b1 6
#843870000000
1!
1%
1-
12
#843880000000
0!
0%
b10 *
0-
02
b10 6
#843890000000
1!
1%
1-
12
#843900000000
0!
0%
b11 *
0-
02
b11 6
#843910000000
1!
1%
1-
12
15
#843920000000
0!
0%
b100 *
0-
02
b100 6
#843930000000
1!
1%
1-
12
#843940000000
0!
0%
b101 *
0-
02
b101 6
#843950000000
1!
1%
1-
12
#843960000000
0!
0%
b110 *
0-
02
b110 6
#843970000000
1!
1%
1-
12
#843980000000
0!
0%
b111 *
0-
02
b111 6
#843990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#844000000000
0!
0%
b0 *
0-
02
b0 6
#844010000000
1!
1%
1-
12
#844020000000
0!
0%
b1 *
0-
02
b1 6
#844030000000
1!
1%
1-
12
#844040000000
0!
0%
b10 *
0-
02
b10 6
#844050000000
1!
1%
1-
12
#844060000000
0!
0%
b11 *
0-
02
b11 6
#844070000000
1!
1%
1-
12
15
#844080000000
0!
0%
b100 *
0-
02
b100 6
#844090000000
1!
1%
1-
12
#844100000000
0!
0%
b101 *
0-
02
b101 6
#844110000000
1!
1%
1-
12
#844120000000
0!
0%
b110 *
0-
02
b110 6
#844130000000
1!
1%
1-
12
#844140000000
0!
0%
b111 *
0-
02
b111 6
#844150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#844160000000
0!
0%
b0 *
0-
02
b0 6
#844170000000
1!
1%
1-
12
#844180000000
0!
0%
b1 *
0-
02
b1 6
#844190000000
1!
1%
1-
12
#844200000000
0!
0%
b10 *
0-
02
b10 6
#844210000000
1!
1%
1-
12
#844220000000
0!
0%
b11 *
0-
02
b11 6
#844230000000
1!
1%
1-
12
15
#844240000000
0!
0%
b100 *
0-
02
b100 6
#844250000000
1!
1%
1-
12
#844260000000
0!
0%
b101 *
0-
02
b101 6
#844270000000
1!
1%
1-
12
#844280000000
0!
0%
b110 *
0-
02
b110 6
#844290000000
1!
1%
1-
12
#844300000000
0!
0%
b111 *
0-
02
b111 6
#844310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#844320000000
0!
0%
b0 *
0-
02
b0 6
#844330000000
1!
1%
1-
12
#844340000000
0!
0%
b1 *
0-
02
b1 6
#844350000000
1!
1%
1-
12
#844360000000
0!
0%
b10 *
0-
02
b10 6
#844370000000
1!
1%
1-
12
#844380000000
0!
0%
b11 *
0-
02
b11 6
#844390000000
1!
1%
1-
12
15
#844400000000
0!
0%
b100 *
0-
02
b100 6
#844410000000
1!
1%
1-
12
#844420000000
0!
0%
b101 *
0-
02
b101 6
#844430000000
1!
1%
1-
12
#844440000000
0!
0%
b110 *
0-
02
b110 6
#844450000000
1!
1%
1-
12
#844460000000
0!
0%
b111 *
0-
02
b111 6
#844470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#844480000000
0!
0%
b0 *
0-
02
b0 6
#844490000000
1!
1%
1-
12
#844500000000
0!
0%
b1 *
0-
02
b1 6
#844510000000
1!
1%
1-
12
#844520000000
0!
0%
b10 *
0-
02
b10 6
#844530000000
1!
1%
1-
12
#844540000000
0!
0%
b11 *
0-
02
b11 6
#844550000000
1!
1%
1-
12
15
#844560000000
0!
0%
b100 *
0-
02
b100 6
#844570000000
1!
1%
1-
12
#844580000000
0!
0%
b101 *
0-
02
b101 6
#844590000000
1!
1%
1-
12
#844600000000
0!
0%
b110 *
0-
02
b110 6
#844610000000
1!
1%
1-
12
#844620000000
0!
0%
b111 *
0-
02
b111 6
#844630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#844640000000
0!
0%
b0 *
0-
02
b0 6
#844650000000
1!
1%
1-
12
#844660000000
0!
0%
b1 *
0-
02
b1 6
#844670000000
1!
1%
1-
12
#844680000000
0!
0%
b10 *
0-
02
b10 6
#844690000000
1!
1%
1-
12
#844700000000
0!
0%
b11 *
0-
02
b11 6
#844710000000
1!
1%
1-
12
15
#844720000000
0!
0%
b100 *
0-
02
b100 6
#844730000000
1!
1%
1-
12
#844740000000
0!
0%
b101 *
0-
02
b101 6
#844750000000
1!
1%
1-
12
#844760000000
0!
0%
b110 *
0-
02
b110 6
#844770000000
1!
1%
1-
12
#844780000000
0!
0%
b111 *
0-
02
b111 6
#844790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#844800000000
0!
0%
b0 *
0-
02
b0 6
#844810000000
1!
1%
1-
12
#844820000000
0!
0%
b1 *
0-
02
b1 6
#844830000000
1!
1%
1-
12
#844840000000
0!
0%
b10 *
0-
02
b10 6
#844850000000
1!
1%
1-
12
#844860000000
0!
0%
b11 *
0-
02
b11 6
#844870000000
1!
1%
1-
12
15
#844880000000
0!
0%
b100 *
0-
02
b100 6
#844890000000
1!
1%
1-
12
#844900000000
0!
0%
b101 *
0-
02
b101 6
#844910000000
1!
1%
1-
12
#844920000000
0!
0%
b110 *
0-
02
b110 6
#844930000000
1!
1%
1-
12
#844940000000
0!
0%
b111 *
0-
02
b111 6
#844950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#844960000000
0!
0%
b0 *
0-
02
b0 6
#844970000000
1!
1%
1-
12
#844980000000
0!
0%
b1 *
0-
02
b1 6
#844990000000
1!
1%
1-
12
#845000000000
0!
0%
b10 *
0-
02
b10 6
#845010000000
1!
1%
1-
12
#845020000000
0!
0%
b11 *
0-
02
b11 6
#845030000000
1!
1%
1-
12
15
#845040000000
0!
0%
b100 *
0-
02
b100 6
#845050000000
1!
1%
1-
12
#845060000000
0!
0%
b101 *
0-
02
b101 6
#845070000000
1!
1%
1-
12
#845080000000
0!
0%
b110 *
0-
02
b110 6
#845090000000
1!
1%
1-
12
#845100000000
0!
0%
b111 *
0-
02
b111 6
#845110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#845120000000
0!
0%
b0 *
0-
02
b0 6
#845130000000
1!
1%
1-
12
#845140000000
0!
0%
b1 *
0-
02
b1 6
#845150000000
1!
1%
1-
12
#845160000000
0!
0%
b10 *
0-
02
b10 6
#845170000000
1!
1%
1-
12
#845180000000
0!
0%
b11 *
0-
02
b11 6
#845190000000
1!
1%
1-
12
15
#845200000000
0!
0%
b100 *
0-
02
b100 6
#845210000000
1!
1%
1-
12
#845220000000
0!
0%
b101 *
0-
02
b101 6
#845230000000
1!
1%
1-
12
#845240000000
0!
0%
b110 *
0-
02
b110 6
#845250000000
1!
1%
1-
12
#845260000000
0!
0%
b111 *
0-
02
b111 6
#845270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#845280000000
0!
0%
b0 *
0-
02
b0 6
#845290000000
1!
1%
1-
12
#845300000000
0!
0%
b1 *
0-
02
b1 6
#845310000000
1!
1%
1-
12
#845320000000
0!
0%
b10 *
0-
02
b10 6
#845330000000
1!
1%
1-
12
#845340000000
0!
0%
b11 *
0-
02
b11 6
#845350000000
1!
1%
1-
12
15
#845360000000
0!
0%
b100 *
0-
02
b100 6
#845370000000
1!
1%
1-
12
#845380000000
0!
0%
b101 *
0-
02
b101 6
#845390000000
1!
1%
1-
12
#845400000000
0!
0%
b110 *
0-
02
b110 6
#845410000000
1!
1%
1-
12
#845420000000
0!
0%
b111 *
0-
02
b111 6
#845430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#845440000000
0!
0%
b0 *
0-
02
b0 6
#845450000000
1!
1%
1-
12
#845460000000
0!
0%
b1 *
0-
02
b1 6
#845470000000
1!
1%
1-
12
#845480000000
0!
0%
b10 *
0-
02
b10 6
#845490000000
1!
1%
1-
12
#845500000000
0!
0%
b11 *
0-
02
b11 6
#845510000000
1!
1%
1-
12
15
#845520000000
0!
0%
b100 *
0-
02
b100 6
#845530000000
1!
1%
1-
12
#845540000000
0!
0%
b101 *
0-
02
b101 6
#845550000000
1!
1%
1-
12
#845560000000
0!
0%
b110 *
0-
02
b110 6
#845570000000
1!
1%
1-
12
#845580000000
0!
0%
b111 *
0-
02
b111 6
#845590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#845600000000
0!
0%
b0 *
0-
02
b0 6
#845610000000
1!
1%
1-
12
#845620000000
0!
0%
b1 *
0-
02
b1 6
#845630000000
1!
1%
1-
12
#845640000000
0!
0%
b10 *
0-
02
b10 6
#845650000000
1!
1%
1-
12
#845660000000
0!
0%
b11 *
0-
02
b11 6
#845670000000
1!
1%
1-
12
15
#845680000000
0!
0%
b100 *
0-
02
b100 6
#845690000000
1!
1%
1-
12
#845700000000
0!
0%
b101 *
0-
02
b101 6
#845710000000
1!
1%
1-
12
#845720000000
0!
0%
b110 *
0-
02
b110 6
#845730000000
1!
1%
1-
12
#845740000000
0!
0%
b111 *
0-
02
b111 6
#845750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#845760000000
0!
0%
b0 *
0-
02
b0 6
#845770000000
1!
1%
1-
12
#845780000000
0!
0%
b1 *
0-
02
b1 6
#845790000000
1!
1%
1-
12
#845800000000
0!
0%
b10 *
0-
02
b10 6
#845810000000
1!
1%
1-
12
#845820000000
0!
0%
b11 *
0-
02
b11 6
#845830000000
1!
1%
1-
12
15
#845840000000
0!
0%
b100 *
0-
02
b100 6
#845850000000
1!
1%
1-
12
#845860000000
0!
0%
b101 *
0-
02
b101 6
#845870000000
1!
1%
1-
12
#845880000000
0!
0%
b110 *
0-
02
b110 6
#845890000000
1!
1%
1-
12
#845900000000
0!
0%
b111 *
0-
02
b111 6
#845910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#845920000000
0!
0%
b0 *
0-
02
b0 6
#845930000000
1!
1%
1-
12
#845940000000
0!
0%
b1 *
0-
02
b1 6
#845950000000
1!
1%
1-
12
#845960000000
0!
0%
b10 *
0-
02
b10 6
#845970000000
1!
1%
1-
12
#845980000000
0!
0%
b11 *
0-
02
b11 6
#845990000000
1!
1%
1-
12
15
#846000000000
0!
0%
b100 *
0-
02
b100 6
#846010000000
1!
1%
1-
12
#846020000000
0!
0%
b101 *
0-
02
b101 6
#846030000000
1!
1%
1-
12
#846040000000
0!
0%
b110 *
0-
02
b110 6
#846050000000
1!
1%
1-
12
#846060000000
0!
0%
b111 *
0-
02
b111 6
#846070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#846080000000
0!
0%
b0 *
0-
02
b0 6
#846090000000
1!
1%
1-
12
#846100000000
0!
0%
b1 *
0-
02
b1 6
#846110000000
1!
1%
1-
12
#846120000000
0!
0%
b10 *
0-
02
b10 6
#846130000000
1!
1%
1-
12
#846140000000
0!
0%
b11 *
0-
02
b11 6
#846150000000
1!
1%
1-
12
15
#846160000000
0!
0%
b100 *
0-
02
b100 6
#846170000000
1!
1%
1-
12
#846180000000
0!
0%
b101 *
0-
02
b101 6
#846190000000
1!
1%
1-
12
#846200000000
0!
0%
b110 *
0-
02
b110 6
#846210000000
1!
1%
1-
12
#846220000000
0!
0%
b111 *
0-
02
b111 6
#846230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#846240000000
0!
0%
b0 *
0-
02
b0 6
#846250000000
1!
1%
1-
12
#846260000000
0!
0%
b1 *
0-
02
b1 6
#846270000000
1!
1%
1-
12
#846280000000
0!
0%
b10 *
0-
02
b10 6
#846290000000
1!
1%
1-
12
#846300000000
0!
0%
b11 *
0-
02
b11 6
#846310000000
1!
1%
1-
12
15
#846320000000
0!
0%
b100 *
0-
02
b100 6
#846330000000
1!
1%
1-
12
#846340000000
0!
0%
b101 *
0-
02
b101 6
#846350000000
1!
1%
1-
12
#846360000000
0!
0%
b110 *
0-
02
b110 6
#846370000000
1!
1%
1-
12
#846380000000
0!
0%
b111 *
0-
02
b111 6
#846390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#846400000000
0!
0%
b0 *
0-
02
b0 6
#846410000000
1!
1%
1-
12
#846420000000
0!
0%
b1 *
0-
02
b1 6
#846430000000
1!
1%
1-
12
#846440000000
0!
0%
b10 *
0-
02
b10 6
#846450000000
1!
1%
1-
12
#846460000000
0!
0%
b11 *
0-
02
b11 6
#846470000000
1!
1%
1-
12
15
#846480000000
0!
0%
b100 *
0-
02
b100 6
#846490000000
1!
1%
1-
12
#846500000000
0!
0%
b101 *
0-
02
b101 6
#846510000000
1!
1%
1-
12
#846520000000
0!
0%
b110 *
0-
02
b110 6
#846530000000
1!
1%
1-
12
#846540000000
0!
0%
b111 *
0-
02
b111 6
#846550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#846560000000
0!
0%
b0 *
0-
02
b0 6
#846570000000
1!
1%
1-
12
#846580000000
0!
0%
b1 *
0-
02
b1 6
#846590000000
1!
1%
1-
12
#846600000000
0!
0%
b10 *
0-
02
b10 6
#846610000000
1!
1%
1-
12
#846620000000
0!
0%
b11 *
0-
02
b11 6
#846630000000
1!
1%
1-
12
15
#846640000000
0!
0%
b100 *
0-
02
b100 6
#846650000000
1!
1%
1-
12
#846660000000
0!
0%
b101 *
0-
02
b101 6
#846670000000
1!
1%
1-
12
#846680000000
0!
0%
b110 *
0-
02
b110 6
#846690000000
1!
1%
1-
12
#846700000000
0!
0%
b111 *
0-
02
b111 6
#846710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#846720000000
0!
0%
b0 *
0-
02
b0 6
#846730000000
1!
1%
1-
12
#846740000000
0!
0%
b1 *
0-
02
b1 6
#846750000000
1!
1%
1-
12
#846760000000
0!
0%
b10 *
0-
02
b10 6
#846770000000
1!
1%
1-
12
#846780000000
0!
0%
b11 *
0-
02
b11 6
#846790000000
1!
1%
1-
12
15
#846800000000
0!
0%
b100 *
0-
02
b100 6
#846810000000
1!
1%
1-
12
#846820000000
0!
0%
b101 *
0-
02
b101 6
#846830000000
1!
1%
1-
12
#846840000000
0!
0%
b110 *
0-
02
b110 6
#846850000000
1!
1%
1-
12
#846860000000
0!
0%
b111 *
0-
02
b111 6
#846870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#846880000000
0!
0%
b0 *
0-
02
b0 6
#846890000000
1!
1%
1-
12
#846900000000
0!
0%
b1 *
0-
02
b1 6
#846910000000
1!
1%
1-
12
#846920000000
0!
0%
b10 *
0-
02
b10 6
#846930000000
1!
1%
1-
12
#846940000000
0!
0%
b11 *
0-
02
b11 6
#846950000000
1!
1%
1-
12
15
#846960000000
0!
0%
b100 *
0-
02
b100 6
#846970000000
1!
1%
1-
12
#846980000000
0!
0%
b101 *
0-
02
b101 6
#846990000000
1!
1%
1-
12
#847000000000
0!
0%
b110 *
0-
02
b110 6
#847010000000
1!
1%
1-
12
#847020000000
0!
0%
b111 *
0-
02
b111 6
#847030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#847040000000
0!
0%
b0 *
0-
02
b0 6
#847050000000
1!
1%
1-
12
#847060000000
0!
0%
b1 *
0-
02
b1 6
#847070000000
1!
1%
1-
12
#847080000000
0!
0%
b10 *
0-
02
b10 6
#847090000000
1!
1%
1-
12
#847100000000
0!
0%
b11 *
0-
02
b11 6
#847110000000
1!
1%
1-
12
15
#847120000000
0!
0%
b100 *
0-
02
b100 6
#847130000000
1!
1%
1-
12
#847140000000
0!
0%
b101 *
0-
02
b101 6
#847150000000
1!
1%
1-
12
#847160000000
0!
0%
b110 *
0-
02
b110 6
#847170000000
1!
1%
1-
12
#847180000000
0!
0%
b111 *
0-
02
b111 6
#847190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#847200000000
0!
0%
b0 *
0-
02
b0 6
#847210000000
1!
1%
1-
12
#847220000000
0!
0%
b1 *
0-
02
b1 6
#847230000000
1!
1%
1-
12
#847240000000
0!
0%
b10 *
0-
02
b10 6
#847250000000
1!
1%
1-
12
#847260000000
0!
0%
b11 *
0-
02
b11 6
#847270000000
1!
1%
1-
12
15
#847280000000
0!
0%
b100 *
0-
02
b100 6
#847290000000
1!
1%
1-
12
#847300000000
0!
0%
b101 *
0-
02
b101 6
#847310000000
1!
1%
1-
12
#847320000000
0!
0%
b110 *
0-
02
b110 6
#847330000000
1!
1%
1-
12
#847340000000
0!
0%
b111 *
0-
02
b111 6
#847350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#847360000000
0!
0%
b0 *
0-
02
b0 6
#847370000000
1!
1%
1-
12
#847380000000
0!
0%
b1 *
0-
02
b1 6
#847390000000
1!
1%
1-
12
#847400000000
0!
0%
b10 *
0-
02
b10 6
#847410000000
1!
1%
1-
12
#847420000000
0!
0%
b11 *
0-
02
b11 6
#847430000000
1!
1%
1-
12
15
#847440000000
0!
0%
b100 *
0-
02
b100 6
#847450000000
1!
1%
1-
12
#847460000000
0!
0%
b101 *
0-
02
b101 6
#847470000000
1!
1%
1-
12
#847480000000
0!
0%
b110 *
0-
02
b110 6
#847490000000
1!
1%
1-
12
#847500000000
0!
0%
b111 *
0-
02
b111 6
#847510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#847520000000
0!
0%
b0 *
0-
02
b0 6
#847530000000
1!
1%
1-
12
#847540000000
0!
0%
b1 *
0-
02
b1 6
#847550000000
1!
1%
1-
12
#847560000000
0!
0%
b10 *
0-
02
b10 6
#847570000000
1!
1%
1-
12
#847580000000
0!
0%
b11 *
0-
02
b11 6
#847590000000
1!
1%
1-
12
15
#847600000000
0!
0%
b100 *
0-
02
b100 6
#847610000000
1!
1%
1-
12
#847620000000
0!
0%
b101 *
0-
02
b101 6
#847630000000
1!
1%
1-
12
#847640000000
0!
0%
b110 *
0-
02
b110 6
#847650000000
1!
1%
1-
12
#847660000000
0!
0%
b111 *
0-
02
b111 6
#847670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#847680000000
0!
0%
b0 *
0-
02
b0 6
#847690000000
1!
1%
1-
12
#847700000000
0!
0%
b1 *
0-
02
b1 6
#847710000000
1!
1%
1-
12
#847720000000
0!
0%
b10 *
0-
02
b10 6
#847730000000
1!
1%
1-
12
#847740000000
0!
0%
b11 *
0-
02
b11 6
#847750000000
1!
1%
1-
12
15
#847760000000
0!
0%
b100 *
0-
02
b100 6
#847770000000
1!
1%
1-
12
#847780000000
0!
0%
b101 *
0-
02
b101 6
#847790000000
1!
1%
1-
12
#847800000000
0!
0%
b110 *
0-
02
b110 6
#847810000000
1!
1%
1-
12
#847820000000
0!
0%
b111 *
0-
02
b111 6
#847830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#847840000000
0!
0%
b0 *
0-
02
b0 6
#847850000000
1!
1%
1-
12
#847860000000
0!
0%
b1 *
0-
02
b1 6
#847870000000
1!
1%
1-
12
#847880000000
0!
0%
b10 *
0-
02
b10 6
#847890000000
1!
1%
1-
12
#847900000000
0!
0%
b11 *
0-
02
b11 6
#847910000000
1!
1%
1-
12
15
#847920000000
0!
0%
b100 *
0-
02
b100 6
#847930000000
1!
1%
1-
12
#847940000000
0!
0%
b101 *
0-
02
b101 6
#847950000000
1!
1%
1-
12
#847960000000
0!
0%
b110 *
0-
02
b110 6
#847970000000
1!
1%
1-
12
#847980000000
0!
0%
b111 *
0-
02
b111 6
#847990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#848000000000
0!
0%
b0 *
0-
02
b0 6
#848010000000
1!
1%
1-
12
#848020000000
0!
0%
b1 *
0-
02
b1 6
#848030000000
1!
1%
1-
12
#848040000000
0!
0%
b10 *
0-
02
b10 6
#848050000000
1!
1%
1-
12
#848060000000
0!
0%
b11 *
0-
02
b11 6
#848070000000
1!
1%
1-
12
15
#848080000000
0!
0%
b100 *
0-
02
b100 6
#848090000000
1!
1%
1-
12
#848100000000
0!
0%
b101 *
0-
02
b101 6
#848110000000
1!
1%
1-
12
#848120000000
0!
0%
b110 *
0-
02
b110 6
#848130000000
1!
1%
1-
12
#848140000000
0!
0%
b111 *
0-
02
b111 6
#848150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#848160000000
0!
0%
b0 *
0-
02
b0 6
#848170000000
1!
1%
1-
12
#848180000000
0!
0%
b1 *
0-
02
b1 6
#848190000000
1!
1%
1-
12
#848200000000
0!
0%
b10 *
0-
02
b10 6
#848210000000
1!
1%
1-
12
#848220000000
0!
0%
b11 *
0-
02
b11 6
#848230000000
1!
1%
1-
12
15
#848240000000
0!
0%
b100 *
0-
02
b100 6
#848250000000
1!
1%
1-
12
#848260000000
0!
0%
b101 *
0-
02
b101 6
#848270000000
1!
1%
1-
12
#848280000000
0!
0%
b110 *
0-
02
b110 6
#848290000000
1!
1%
1-
12
#848300000000
0!
0%
b111 *
0-
02
b111 6
#848310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#848320000000
0!
0%
b0 *
0-
02
b0 6
#848330000000
1!
1%
1-
12
#848340000000
0!
0%
b1 *
0-
02
b1 6
#848350000000
1!
1%
1-
12
#848360000000
0!
0%
b10 *
0-
02
b10 6
#848370000000
1!
1%
1-
12
#848380000000
0!
0%
b11 *
0-
02
b11 6
#848390000000
1!
1%
1-
12
15
#848400000000
0!
0%
b100 *
0-
02
b100 6
#848410000000
1!
1%
1-
12
#848420000000
0!
0%
b101 *
0-
02
b101 6
#848430000000
1!
1%
1-
12
#848440000000
0!
0%
b110 *
0-
02
b110 6
#848450000000
1!
1%
1-
12
#848460000000
0!
0%
b111 *
0-
02
b111 6
#848470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#848480000000
0!
0%
b0 *
0-
02
b0 6
#848490000000
1!
1%
1-
12
#848500000000
0!
0%
b1 *
0-
02
b1 6
#848510000000
1!
1%
1-
12
#848520000000
0!
0%
b10 *
0-
02
b10 6
#848530000000
1!
1%
1-
12
#848540000000
0!
0%
b11 *
0-
02
b11 6
#848550000000
1!
1%
1-
12
15
#848560000000
0!
0%
b100 *
0-
02
b100 6
#848570000000
1!
1%
1-
12
#848580000000
0!
0%
b101 *
0-
02
b101 6
#848590000000
1!
1%
1-
12
#848600000000
0!
0%
b110 *
0-
02
b110 6
#848610000000
1!
1%
1-
12
#848620000000
0!
0%
b111 *
0-
02
b111 6
#848630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#848640000000
0!
0%
b0 *
0-
02
b0 6
#848650000000
1!
1%
1-
12
#848660000000
0!
0%
b1 *
0-
02
b1 6
#848670000000
1!
1%
1-
12
#848680000000
0!
0%
b10 *
0-
02
b10 6
#848690000000
1!
1%
1-
12
#848700000000
0!
0%
b11 *
0-
02
b11 6
#848710000000
1!
1%
1-
12
15
#848720000000
0!
0%
b100 *
0-
02
b100 6
#848730000000
1!
1%
1-
12
#848740000000
0!
0%
b101 *
0-
02
b101 6
#848750000000
1!
1%
1-
12
#848760000000
0!
0%
b110 *
0-
02
b110 6
#848770000000
1!
1%
1-
12
#848780000000
0!
0%
b111 *
0-
02
b111 6
#848790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#848800000000
0!
0%
b0 *
0-
02
b0 6
#848810000000
1!
1%
1-
12
#848820000000
0!
0%
b1 *
0-
02
b1 6
#848830000000
1!
1%
1-
12
#848840000000
0!
0%
b10 *
0-
02
b10 6
#848850000000
1!
1%
1-
12
#848860000000
0!
0%
b11 *
0-
02
b11 6
#848870000000
1!
1%
1-
12
15
#848880000000
0!
0%
b100 *
0-
02
b100 6
#848890000000
1!
1%
1-
12
#848900000000
0!
0%
b101 *
0-
02
b101 6
#848910000000
1!
1%
1-
12
#848920000000
0!
0%
b110 *
0-
02
b110 6
#848930000000
1!
1%
1-
12
#848940000000
0!
0%
b111 *
0-
02
b111 6
#848950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#848960000000
0!
0%
b0 *
0-
02
b0 6
#848970000000
1!
1%
1-
12
#848980000000
0!
0%
b1 *
0-
02
b1 6
#848990000000
1!
1%
1-
12
#849000000000
0!
0%
b10 *
0-
02
b10 6
#849010000000
1!
1%
1-
12
#849020000000
0!
0%
b11 *
0-
02
b11 6
#849030000000
1!
1%
1-
12
15
#849040000000
0!
0%
b100 *
0-
02
b100 6
#849050000000
1!
1%
1-
12
#849060000000
0!
0%
b101 *
0-
02
b101 6
#849070000000
1!
1%
1-
12
#849080000000
0!
0%
b110 *
0-
02
b110 6
#849090000000
1!
1%
1-
12
#849100000000
0!
0%
b111 *
0-
02
b111 6
#849110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#849120000000
0!
0%
b0 *
0-
02
b0 6
#849130000000
1!
1%
1-
12
#849140000000
0!
0%
b1 *
0-
02
b1 6
#849150000000
1!
1%
1-
12
#849160000000
0!
0%
b10 *
0-
02
b10 6
#849170000000
1!
1%
1-
12
#849180000000
0!
0%
b11 *
0-
02
b11 6
#849190000000
1!
1%
1-
12
15
#849200000000
0!
0%
b100 *
0-
02
b100 6
#849210000000
1!
1%
1-
12
#849220000000
0!
0%
b101 *
0-
02
b101 6
#849230000000
1!
1%
1-
12
#849240000000
0!
0%
b110 *
0-
02
b110 6
#849250000000
1!
1%
1-
12
#849260000000
0!
0%
b111 *
0-
02
b111 6
#849270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#849280000000
0!
0%
b0 *
0-
02
b0 6
#849290000000
1!
1%
1-
12
#849300000000
0!
0%
b1 *
0-
02
b1 6
#849310000000
1!
1%
1-
12
#849320000000
0!
0%
b10 *
0-
02
b10 6
#849330000000
1!
1%
1-
12
#849340000000
0!
0%
b11 *
0-
02
b11 6
#849350000000
1!
1%
1-
12
15
#849360000000
0!
0%
b100 *
0-
02
b100 6
#849370000000
1!
1%
1-
12
#849380000000
0!
0%
b101 *
0-
02
b101 6
#849390000000
1!
1%
1-
12
#849400000000
0!
0%
b110 *
0-
02
b110 6
#849410000000
1!
1%
1-
12
#849420000000
0!
0%
b111 *
0-
02
b111 6
#849430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#849440000000
0!
0%
b0 *
0-
02
b0 6
#849450000000
1!
1%
1-
12
#849460000000
0!
0%
b1 *
0-
02
b1 6
#849470000000
1!
1%
1-
12
#849480000000
0!
0%
b10 *
0-
02
b10 6
#849490000000
1!
1%
1-
12
#849500000000
0!
0%
b11 *
0-
02
b11 6
#849510000000
1!
1%
1-
12
15
#849520000000
0!
0%
b100 *
0-
02
b100 6
#849530000000
1!
1%
1-
12
#849540000000
0!
0%
b101 *
0-
02
b101 6
#849550000000
1!
1%
1-
12
#849560000000
0!
0%
b110 *
0-
02
b110 6
#849570000000
1!
1%
1-
12
#849580000000
0!
0%
b111 *
0-
02
b111 6
#849590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#849600000000
0!
0%
b0 *
0-
02
b0 6
#849610000000
1!
1%
1-
12
#849620000000
0!
0%
b1 *
0-
02
b1 6
#849630000000
1!
1%
1-
12
#849640000000
0!
0%
b10 *
0-
02
b10 6
#849650000000
1!
1%
1-
12
#849660000000
0!
0%
b11 *
0-
02
b11 6
#849670000000
1!
1%
1-
12
15
#849680000000
0!
0%
b100 *
0-
02
b100 6
#849690000000
1!
1%
1-
12
#849700000000
0!
0%
b101 *
0-
02
b101 6
#849710000000
1!
1%
1-
12
#849720000000
0!
0%
b110 *
0-
02
b110 6
#849730000000
1!
1%
1-
12
#849740000000
0!
0%
b111 *
0-
02
b111 6
#849750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#849760000000
0!
0%
b0 *
0-
02
b0 6
#849770000000
1!
1%
1-
12
#849780000000
0!
0%
b1 *
0-
02
b1 6
#849790000000
1!
1%
1-
12
#849800000000
0!
0%
b10 *
0-
02
b10 6
#849810000000
1!
1%
1-
12
#849820000000
0!
0%
b11 *
0-
02
b11 6
#849830000000
1!
1%
1-
12
15
#849840000000
0!
0%
b100 *
0-
02
b100 6
#849850000000
1!
1%
1-
12
#849860000000
0!
0%
b101 *
0-
02
b101 6
#849870000000
1!
1%
1-
12
#849880000000
0!
0%
b110 *
0-
02
b110 6
#849890000000
1!
1%
1-
12
#849900000000
0!
0%
b111 *
0-
02
b111 6
#849910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#849920000000
0!
0%
b0 *
0-
02
b0 6
#849930000000
1!
1%
1-
12
#849940000000
0!
0%
b1 *
0-
02
b1 6
#849950000000
1!
1%
1-
12
#849960000000
0!
0%
b10 *
0-
02
b10 6
#849970000000
1!
1%
1-
12
#849980000000
0!
0%
b11 *
0-
02
b11 6
#849990000000
1!
1%
1-
12
15
#850000000000
0!
0%
b100 *
0-
02
b100 6
#850010000000
1!
1%
1-
12
#850020000000
0!
0%
b101 *
0-
02
b101 6
#850030000000
1!
1%
1-
12
#850040000000
0!
0%
b110 *
0-
02
b110 6
#850050000000
1!
1%
1-
12
#850060000000
0!
0%
b111 *
0-
02
b111 6
#850070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#850080000000
0!
0%
b0 *
0-
02
b0 6
#850090000000
1!
1%
1-
12
#850100000000
0!
0%
b1 *
0-
02
b1 6
#850110000000
1!
1%
1-
12
#850120000000
0!
0%
b10 *
0-
02
b10 6
#850130000000
1!
1%
1-
12
#850140000000
0!
0%
b11 *
0-
02
b11 6
#850150000000
1!
1%
1-
12
15
#850160000000
0!
0%
b100 *
0-
02
b100 6
#850170000000
1!
1%
1-
12
#850180000000
0!
0%
b101 *
0-
02
b101 6
#850190000000
1!
1%
1-
12
#850200000000
0!
0%
b110 *
0-
02
b110 6
#850210000000
1!
1%
1-
12
#850220000000
0!
0%
b111 *
0-
02
b111 6
#850230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#850240000000
0!
0%
b0 *
0-
02
b0 6
#850250000000
1!
1%
1-
12
#850260000000
0!
0%
b1 *
0-
02
b1 6
#850270000000
1!
1%
1-
12
#850280000000
0!
0%
b10 *
0-
02
b10 6
#850290000000
1!
1%
1-
12
#850300000000
0!
0%
b11 *
0-
02
b11 6
#850310000000
1!
1%
1-
12
15
#850320000000
0!
0%
b100 *
0-
02
b100 6
#850330000000
1!
1%
1-
12
#850340000000
0!
0%
b101 *
0-
02
b101 6
#850350000000
1!
1%
1-
12
#850360000000
0!
0%
b110 *
0-
02
b110 6
#850370000000
1!
1%
1-
12
#850380000000
0!
0%
b111 *
0-
02
b111 6
#850390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#850400000000
0!
0%
b0 *
0-
02
b0 6
#850410000000
1!
1%
1-
12
#850420000000
0!
0%
b1 *
0-
02
b1 6
#850430000000
1!
1%
1-
12
#850440000000
0!
0%
b10 *
0-
02
b10 6
#850450000000
1!
1%
1-
12
#850460000000
0!
0%
b11 *
0-
02
b11 6
#850470000000
1!
1%
1-
12
15
#850480000000
0!
0%
b100 *
0-
02
b100 6
#850490000000
1!
1%
1-
12
#850500000000
0!
0%
b101 *
0-
02
b101 6
#850510000000
1!
1%
1-
12
#850520000000
0!
0%
b110 *
0-
02
b110 6
#850530000000
1!
1%
1-
12
#850540000000
0!
0%
b111 *
0-
02
b111 6
#850550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#850560000000
0!
0%
b0 *
0-
02
b0 6
#850570000000
1!
1%
1-
12
#850580000000
0!
0%
b1 *
0-
02
b1 6
#850590000000
1!
1%
1-
12
#850600000000
0!
0%
b10 *
0-
02
b10 6
#850610000000
1!
1%
1-
12
#850620000000
0!
0%
b11 *
0-
02
b11 6
#850630000000
1!
1%
1-
12
15
#850640000000
0!
0%
b100 *
0-
02
b100 6
#850650000000
1!
1%
1-
12
#850660000000
0!
0%
b101 *
0-
02
b101 6
#850670000000
1!
1%
1-
12
#850680000000
0!
0%
b110 *
0-
02
b110 6
#850690000000
1!
1%
1-
12
#850700000000
0!
0%
b111 *
0-
02
b111 6
#850710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#850720000000
0!
0%
b0 *
0-
02
b0 6
#850730000000
1!
1%
1-
12
#850740000000
0!
0%
b1 *
0-
02
b1 6
#850750000000
1!
1%
1-
12
#850760000000
0!
0%
b10 *
0-
02
b10 6
#850770000000
1!
1%
1-
12
#850780000000
0!
0%
b11 *
0-
02
b11 6
#850790000000
1!
1%
1-
12
15
#850800000000
0!
0%
b100 *
0-
02
b100 6
#850810000000
1!
1%
1-
12
#850820000000
0!
0%
b101 *
0-
02
b101 6
#850830000000
1!
1%
1-
12
#850840000000
0!
0%
b110 *
0-
02
b110 6
#850850000000
1!
1%
1-
12
#850860000000
0!
0%
b111 *
0-
02
b111 6
#850870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#850880000000
0!
0%
b0 *
0-
02
b0 6
#850890000000
1!
1%
1-
12
#850900000000
0!
0%
b1 *
0-
02
b1 6
#850910000000
1!
1%
1-
12
#850920000000
0!
0%
b10 *
0-
02
b10 6
#850930000000
1!
1%
1-
12
#850940000000
0!
0%
b11 *
0-
02
b11 6
#850950000000
1!
1%
1-
12
15
#850960000000
0!
0%
b100 *
0-
02
b100 6
#850970000000
1!
1%
1-
12
#850980000000
0!
0%
b101 *
0-
02
b101 6
#850990000000
1!
1%
1-
12
#851000000000
0!
0%
b110 *
0-
02
b110 6
#851010000000
1!
1%
1-
12
#851020000000
0!
0%
b111 *
0-
02
b111 6
#851030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#851040000000
0!
0%
b0 *
0-
02
b0 6
#851050000000
1!
1%
1-
12
#851060000000
0!
0%
b1 *
0-
02
b1 6
#851070000000
1!
1%
1-
12
#851080000000
0!
0%
b10 *
0-
02
b10 6
#851090000000
1!
1%
1-
12
#851100000000
0!
0%
b11 *
0-
02
b11 6
#851110000000
1!
1%
1-
12
15
#851120000000
0!
0%
b100 *
0-
02
b100 6
#851130000000
1!
1%
1-
12
#851140000000
0!
0%
b101 *
0-
02
b101 6
#851150000000
1!
1%
1-
12
#851160000000
0!
0%
b110 *
0-
02
b110 6
#851170000000
1!
1%
1-
12
#851180000000
0!
0%
b111 *
0-
02
b111 6
#851190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#851200000000
0!
0%
b0 *
0-
02
b0 6
#851210000000
1!
1%
1-
12
#851220000000
0!
0%
b1 *
0-
02
b1 6
#851230000000
1!
1%
1-
12
#851240000000
0!
0%
b10 *
0-
02
b10 6
#851250000000
1!
1%
1-
12
#851260000000
0!
0%
b11 *
0-
02
b11 6
#851270000000
1!
1%
1-
12
15
#851280000000
0!
0%
b100 *
0-
02
b100 6
#851290000000
1!
1%
1-
12
#851300000000
0!
0%
b101 *
0-
02
b101 6
#851310000000
1!
1%
1-
12
#851320000000
0!
0%
b110 *
0-
02
b110 6
#851330000000
1!
1%
1-
12
#851340000000
0!
0%
b111 *
0-
02
b111 6
#851350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#851360000000
0!
0%
b0 *
0-
02
b0 6
#851370000000
1!
1%
1-
12
#851380000000
0!
0%
b1 *
0-
02
b1 6
#851390000000
1!
1%
1-
12
#851400000000
0!
0%
b10 *
0-
02
b10 6
#851410000000
1!
1%
1-
12
#851420000000
0!
0%
b11 *
0-
02
b11 6
#851430000000
1!
1%
1-
12
15
#851440000000
0!
0%
b100 *
0-
02
b100 6
#851450000000
1!
1%
1-
12
#851460000000
0!
0%
b101 *
0-
02
b101 6
#851470000000
1!
1%
1-
12
#851480000000
0!
0%
b110 *
0-
02
b110 6
#851490000000
1!
1%
1-
12
#851500000000
0!
0%
b111 *
0-
02
b111 6
#851510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#851520000000
0!
0%
b0 *
0-
02
b0 6
#851530000000
1!
1%
1-
12
#851540000000
0!
0%
b1 *
0-
02
b1 6
#851550000000
1!
1%
1-
12
#851560000000
0!
0%
b10 *
0-
02
b10 6
#851570000000
1!
1%
1-
12
#851580000000
0!
0%
b11 *
0-
02
b11 6
#851590000000
1!
1%
1-
12
15
#851600000000
0!
0%
b100 *
0-
02
b100 6
#851610000000
1!
1%
1-
12
#851620000000
0!
0%
b101 *
0-
02
b101 6
#851630000000
1!
1%
1-
12
#851640000000
0!
0%
b110 *
0-
02
b110 6
#851650000000
1!
1%
1-
12
#851660000000
0!
0%
b111 *
0-
02
b111 6
#851670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#851680000000
0!
0%
b0 *
0-
02
b0 6
#851690000000
1!
1%
1-
12
#851700000000
0!
0%
b1 *
0-
02
b1 6
#851710000000
1!
1%
1-
12
#851720000000
0!
0%
b10 *
0-
02
b10 6
#851730000000
1!
1%
1-
12
#851740000000
0!
0%
b11 *
0-
02
b11 6
#851750000000
1!
1%
1-
12
15
#851760000000
0!
0%
b100 *
0-
02
b100 6
#851770000000
1!
1%
1-
12
#851780000000
0!
0%
b101 *
0-
02
b101 6
#851790000000
1!
1%
1-
12
#851800000000
0!
0%
b110 *
0-
02
b110 6
#851810000000
1!
1%
1-
12
#851820000000
0!
0%
b111 *
0-
02
b111 6
#851830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#851840000000
0!
0%
b0 *
0-
02
b0 6
#851850000000
1!
1%
1-
12
#851860000000
0!
0%
b1 *
0-
02
b1 6
#851870000000
1!
1%
1-
12
#851880000000
0!
0%
b10 *
0-
02
b10 6
#851890000000
1!
1%
1-
12
#851900000000
0!
0%
b11 *
0-
02
b11 6
#851910000000
1!
1%
1-
12
15
#851920000000
0!
0%
b100 *
0-
02
b100 6
#851930000000
1!
1%
1-
12
#851940000000
0!
0%
b101 *
0-
02
b101 6
#851950000000
1!
1%
1-
12
#851960000000
0!
0%
b110 *
0-
02
b110 6
#851970000000
1!
1%
1-
12
#851980000000
0!
0%
b111 *
0-
02
b111 6
#851990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#852000000000
0!
0%
b0 *
0-
02
b0 6
#852010000000
1!
1%
1-
12
#852020000000
0!
0%
b1 *
0-
02
b1 6
#852030000000
1!
1%
1-
12
#852040000000
0!
0%
b10 *
0-
02
b10 6
#852050000000
1!
1%
1-
12
#852060000000
0!
0%
b11 *
0-
02
b11 6
#852070000000
1!
1%
1-
12
15
#852080000000
0!
0%
b100 *
0-
02
b100 6
#852090000000
1!
1%
1-
12
#852100000000
0!
0%
b101 *
0-
02
b101 6
#852110000000
1!
1%
1-
12
#852120000000
0!
0%
b110 *
0-
02
b110 6
#852130000000
1!
1%
1-
12
#852140000000
0!
0%
b111 *
0-
02
b111 6
#852150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#852160000000
0!
0%
b0 *
0-
02
b0 6
#852170000000
1!
1%
1-
12
#852180000000
0!
0%
b1 *
0-
02
b1 6
#852190000000
1!
1%
1-
12
#852200000000
0!
0%
b10 *
0-
02
b10 6
#852210000000
1!
1%
1-
12
#852220000000
0!
0%
b11 *
0-
02
b11 6
#852230000000
1!
1%
1-
12
15
#852240000000
0!
0%
b100 *
0-
02
b100 6
#852250000000
1!
1%
1-
12
#852260000000
0!
0%
b101 *
0-
02
b101 6
#852270000000
1!
1%
1-
12
#852280000000
0!
0%
b110 *
0-
02
b110 6
#852290000000
1!
1%
1-
12
#852300000000
0!
0%
b111 *
0-
02
b111 6
#852310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#852320000000
0!
0%
b0 *
0-
02
b0 6
#852330000000
1!
1%
1-
12
#852340000000
0!
0%
b1 *
0-
02
b1 6
#852350000000
1!
1%
1-
12
#852360000000
0!
0%
b10 *
0-
02
b10 6
#852370000000
1!
1%
1-
12
#852380000000
0!
0%
b11 *
0-
02
b11 6
#852390000000
1!
1%
1-
12
15
#852400000000
0!
0%
b100 *
0-
02
b100 6
#852410000000
1!
1%
1-
12
#852420000000
0!
0%
b101 *
0-
02
b101 6
#852430000000
1!
1%
1-
12
#852440000000
0!
0%
b110 *
0-
02
b110 6
#852450000000
1!
1%
1-
12
#852460000000
0!
0%
b111 *
0-
02
b111 6
#852470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#852480000000
0!
0%
b0 *
0-
02
b0 6
#852490000000
1!
1%
1-
12
#852500000000
0!
0%
b1 *
0-
02
b1 6
#852510000000
1!
1%
1-
12
#852520000000
0!
0%
b10 *
0-
02
b10 6
#852530000000
1!
1%
1-
12
#852540000000
0!
0%
b11 *
0-
02
b11 6
#852550000000
1!
1%
1-
12
15
#852560000000
0!
0%
b100 *
0-
02
b100 6
#852570000000
1!
1%
1-
12
#852580000000
0!
0%
b101 *
0-
02
b101 6
#852590000000
1!
1%
1-
12
#852600000000
0!
0%
b110 *
0-
02
b110 6
#852610000000
1!
1%
1-
12
#852620000000
0!
0%
b111 *
0-
02
b111 6
#852630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#852640000000
0!
0%
b0 *
0-
02
b0 6
#852650000000
1!
1%
1-
12
#852660000000
0!
0%
b1 *
0-
02
b1 6
#852670000000
1!
1%
1-
12
#852680000000
0!
0%
b10 *
0-
02
b10 6
#852690000000
1!
1%
1-
12
#852700000000
0!
0%
b11 *
0-
02
b11 6
#852710000000
1!
1%
1-
12
15
#852720000000
0!
0%
b100 *
0-
02
b100 6
#852730000000
1!
1%
1-
12
#852740000000
0!
0%
b101 *
0-
02
b101 6
#852750000000
1!
1%
1-
12
#852760000000
0!
0%
b110 *
0-
02
b110 6
#852770000000
1!
1%
1-
12
#852780000000
0!
0%
b111 *
0-
02
b111 6
#852790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#852800000000
0!
0%
b0 *
0-
02
b0 6
#852810000000
1!
1%
1-
12
#852820000000
0!
0%
b1 *
0-
02
b1 6
#852830000000
1!
1%
1-
12
#852840000000
0!
0%
b10 *
0-
02
b10 6
#852850000000
1!
1%
1-
12
#852860000000
0!
0%
b11 *
0-
02
b11 6
#852870000000
1!
1%
1-
12
15
#852880000000
0!
0%
b100 *
0-
02
b100 6
#852890000000
1!
1%
1-
12
#852900000000
0!
0%
b101 *
0-
02
b101 6
#852910000000
1!
1%
1-
12
#852920000000
0!
0%
b110 *
0-
02
b110 6
#852930000000
1!
1%
1-
12
#852940000000
0!
0%
b111 *
0-
02
b111 6
#852950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#852960000000
0!
0%
b0 *
0-
02
b0 6
#852970000000
1!
1%
1-
12
#852980000000
0!
0%
b1 *
0-
02
b1 6
#852990000000
1!
1%
1-
12
#853000000000
0!
0%
b10 *
0-
02
b10 6
#853010000000
1!
1%
1-
12
#853020000000
0!
0%
b11 *
0-
02
b11 6
#853030000000
1!
1%
1-
12
15
#853040000000
0!
0%
b100 *
0-
02
b100 6
#853050000000
1!
1%
1-
12
#853060000000
0!
0%
b101 *
0-
02
b101 6
#853070000000
1!
1%
1-
12
#853080000000
0!
0%
b110 *
0-
02
b110 6
#853090000000
1!
1%
1-
12
#853100000000
0!
0%
b111 *
0-
02
b111 6
#853110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#853120000000
0!
0%
b0 *
0-
02
b0 6
#853130000000
1!
1%
1-
12
#853140000000
0!
0%
b1 *
0-
02
b1 6
#853150000000
1!
1%
1-
12
#853160000000
0!
0%
b10 *
0-
02
b10 6
#853170000000
1!
1%
1-
12
#853180000000
0!
0%
b11 *
0-
02
b11 6
#853190000000
1!
1%
1-
12
15
#853200000000
0!
0%
b100 *
0-
02
b100 6
#853210000000
1!
1%
1-
12
#853220000000
0!
0%
b101 *
0-
02
b101 6
#853230000000
1!
1%
1-
12
#853240000000
0!
0%
b110 *
0-
02
b110 6
#853250000000
1!
1%
1-
12
#853260000000
0!
0%
b111 *
0-
02
b111 6
#853270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#853280000000
0!
0%
b0 *
0-
02
b0 6
#853290000000
1!
1%
1-
12
#853300000000
0!
0%
b1 *
0-
02
b1 6
#853310000000
1!
1%
1-
12
#853320000000
0!
0%
b10 *
0-
02
b10 6
#853330000000
1!
1%
1-
12
#853340000000
0!
0%
b11 *
0-
02
b11 6
#853350000000
1!
1%
1-
12
15
#853360000000
0!
0%
b100 *
0-
02
b100 6
#853370000000
1!
1%
1-
12
#853380000000
0!
0%
b101 *
0-
02
b101 6
#853390000000
1!
1%
1-
12
#853400000000
0!
0%
b110 *
0-
02
b110 6
#853410000000
1!
1%
1-
12
#853420000000
0!
0%
b111 *
0-
02
b111 6
#853430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#853440000000
0!
0%
b0 *
0-
02
b0 6
#853450000000
1!
1%
1-
12
#853460000000
0!
0%
b1 *
0-
02
b1 6
#853470000000
1!
1%
1-
12
#853480000000
0!
0%
b10 *
0-
02
b10 6
#853490000000
1!
1%
1-
12
#853500000000
0!
0%
b11 *
0-
02
b11 6
#853510000000
1!
1%
1-
12
15
#853520000000
0!
0%
b100 *
0-
02
b100 6
#853530000000
1!
1%
1-
12
#853540000000
0!
0%
b101 *
0-
02
b101 6
#853550000000
1!
1%
1-
12
#853560000000
0!
0%
b110 *
0-
02
b110 6
#853570000000
1!
1%
1-
12
#853580000000
0!
0%
b111 *
0-
02
b111 6
#853590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#853600000000
0!
0%
b0 *
0-
02
b0 6
#853610000000
1!
1%
1-
12
#853620000000
0!
0%
b1 *
0-
02
b1 6
#853630000000
1!
1%
1-
12
#853640000000
0!
0%
b10 *
0-
02
b10 6
#853650000000
1!
1%
1-
12
#853660000000
0!
0%
b11 *
0-
02
b11 6
#853670000000
1!
1%
1-
12
15
#853680000000
0!
0%
b100 *
0-
02
b100 6
#853690000000
1!
1%
1-
12
#853700000000
0!
0%
b101 *
0-
02
b101 6
#853710000000
1!
1%
1-
12
#853720000000
0!
0%
b110 *
0-
02
b110 6
#853730000000
1!
1%
1-
12
#853740000000
0!
0%
b111 *
0-
02
b111 6
#853750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#853760000000
0!
0%
b0 *
0-
02
b0 6
#853770000000
1!
1%
1-
12
#853780000000
0!
0%
b1 *
0-
02
b1 6
#853790000000
1!
1%
1-
12
#853800000000
0!
0%
b10 *
0-
02
b10 6
#853810000000
1!
1%
1-
12
#853820000000
0!
0%
b11 *
0-
02
b11 6
#853830000000
1!
1%
1-
12
15
#853840000000
0!
0%
b100 *
0-
02
b100 6
#853850000000
1!
1%
1-
12
#853860000000
0!
0%
b101 *
0-
02
b101 6
#853870000000
1!
1%
1-
12
#853880000000
0!
0%
b110 *
0-
02
b110 6
#853890000000
1!
1%
1-
12
#853900000000
0!
0%
b111 *
0-
02
b111 6
#853910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#853920000000
0!
0%
b0 *
0-
02
b0 6
#853930000000
1!
1%
1-
12
#853940000000
0!
0%
b1 *
0-
02
b1 6
#853950000000
1!
1%
1-
12
#853960000000
0!
0%
b10 *
0-
02
b10 6
#853970000000
1!
1%
1-
12
#853980000000
0!
0%
b11 *
0-
02
b11 6
#853990000000
1!
1%
1-
12
15
#854000000000
0!
0%
b100 *
0-
02
b100 6
#854010000000
1!
1%
1-
12
#854020000000
0!
0%
b101 *
0-
02
b101 6
#854030000000
1!
1%
1-
12
#854040000000
0!
0%
b110 *
0-
02
b110 6
#854050000000
1!
1%
1-
12
#854060000000
0!
0%
b111 *
0-
02
b111 6
#854070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#854080000000
0!
0%
b0 *
0-
02
b0 6
#854090000000
1!
1%
1-
12
#854100000000
0!
0%
b1 *
0-
02
b1 6
#854110000000
1!
1%
1-
12
#854120000000
0!
0%
b10 *
0-
02
b10 6
#854130000000
1!
1%
1-
12
#854140000000
0!
0%
b11 *
0-
02
b11 6
#854150000000
1!
1%
1-
12
15
#854160000000
0!
0%
b100 *
0-
02
b100 6
#854170000000
1!
1%
1-
12
#854180000000
0!
0%
b101 *
0-
02
b101 6
#854190000000
1!
1%
1-
12
#854200000000
0!
0%
b110 *
0-
02
b110 6
#854210000000
1!
1%
1-
12
#854220000000
0!
0%
b111 *
0-
02
b111 6
#854230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#854240000000
0!
0%
b0 *
0-
02
b0 6
#854250000000
1!
1%
1-
12
#854260000000
0!
0%
b1 *
0-
02
b1 6
#854270000000
1!
1%
1-
12
#854280000000
0!
0%
b10 *
0-
02
b10 6
#854290000000
1!
1%
1-
12
#854300000000
0!
0%
b11 *
0-
02
b11 6
#854310000000
1!
1%
1-
12
15
#854320000000
0!
0%
b100 *
0-
02
b100 6
#854330000000
1!
1%
1-
12
#854340000000
0!
0%
b101 *
0-
02
b101 6
#854350000000
1!
1%
1-
12
#854360000000
0!
0%
b110 *
0-
02
b110 6
#854370000000
1!
1%
1-
12
#854380000000
0!
0%
b111 *
0-
02
b111 6
#854390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#854400000000
0!
0%
b0 *
0-
02
b0 6
#854410000000
1!
1%
1-
12
#854420000000
0!
0%
b1 *
0-
02
b1 6
#854430000000
1!
1%
1-
12
#854440000000
0!
0%
b10 *
0-
02
b10 6
#854450000000
1!
1%
1-
12
#854460000000
0!
0%
b11 *
0-
02
b11 6
#854470000000
1!
1%
1-
12
15
#854480000000
0!
0%
b100 *
0-
02
b100 6
#854490000000
1!
1%
1-
12
#854500000000
0!
0%
b101 *
0-
02
b101 6
#854510000000
1!
1%
1-
12
#854520000000
0!
0%
b110 *
0-
02
b110 6
#854530000000
1!
1%
1-
12
#854540000000
0!
0%
b111 *
0-
02
b111 6
#854550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#854560000000
0!
0%
b0 *
0-
02
b0 6
#854570000000
1!
1%
1-
12
#854580000000
0!
0%
b1 *
0-
02
b1 6
#854590000000
1!
1%
1-
12
#854600000000
0!
0%
b10 *
0-
02
b10 6
#854610000000
1!
1%
1-
12
#854620000000
0!
0%
b11 *
0-
02
b11 6
#854630000000
1!
1%
1-
12
15
#854640000000
0!
0%
b100 *
0-
02
b100 6
#854650000000
1!
1%
1-
12
#854660000000
0!
0%
b101 *
0-
02
b101 6
#854670000000
1!
1%
1-
12
#854680000000
0!
0%
b110 *
0-
02
b110 6
#854690000000
1!
1%
1-
12
#854700000000
0!
0%
b111 *
0-
02
b111 6
#854710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#854720000000
0!
0%
b0 *
0-
02
b0 6
#854730000000
1!
1%
1-
12
#854740000000
0!
0%
b1 *
0-
02
b1 6
#854750000000
1!
1%
1-
12
#854760000000
0!
0%
b10 *
0-
02
b10 6
#854770000000
1!
1%
1-
12
#854780000000
0!
0%
b11 *
0-
02
b11 6
#854790000000
1!
1%
1-
12
15
#854800000000
0!
0%
b100 *
0-
02
b100 6
#854810000000
1!
1%
1-
12
#854820000000
0!
0%
b101 *
0-
02
b101 6
#854830000000
1!
1%
1-
12
#854840000000
0!
0%
b110 *
0-
02
b110 6
#854850000000
1!
1%
1-
12
#854860000000
0!
0%
b111 *
0-
02
b111 6
#854870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#854880000000
0!
0%
b0 *
0-
02
b0 6
#854890000000
1!
1%
1-
12
#854900000000
0!
0%
b1 *
0-
02
b1 6
#854910000000
1!
1%
1-
12
#854920000000
0!
0%
b10 *
0-
02
b10 6
#854930000000
1!
1%
1-
12
#854940000000
0!
0%
b11 *
0-
02
b11 6
#854950000000
1!
1%
1-
12
15
#854960000000
0!
0%
b100 *
0-
02
b100 6
#854970000000
1!
1%
1-
12
#854980000000
0!
0%
b101 *
0-
02
b101 6
#854990000000
1!
1%
1-
12
#855000000000
0!
0%
b110 *
0-
02
b110 6
#855010000000
1!
1%
1-
12
#855020000000
0!
0%
b111 *
0-
02
b111 6
#855030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#855040000000
0!
0%
b0 *
0-
02
b0 6
#855050000000
1!
1%
1-
12
#855060000000
0!
0%
b1 *
0-
02
b1 6
#855070000000
1!
1%
1-
12
#855080000000
0!
0%
b10 *
0-
02
b10 6
#855090000000
1!
1%
1-
12
#855100000000
0!
0%
b11 *
0-
02
b11 6
#855110000000
1!
1%
1-
12
15
#855120000000
0!
0%
b100 *
0-
02
b100 6
#855130000000
1!
1%
1-
12
#855140000000
0!
0%
b101 *
0-
02
b101 6
#855150000000
1!
1%
1-
12
#855160000000
0!
0%
b110 *
0-
02
b110 6
#855170000000
1!
1%
1-
12
#855180000000
0!
0%
b111 *
0-
02
b111 6
#855190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#855200000000
0!
0%
b0 *
0-
02
b0 6
#855210000000
1!
1%
1-
12
#855220000000
0!
0%
b1 *
0-
02
b1 6
#855230000000
1!
1%
1-
12
#855240000000
0!
0%
b10 *
0-
02
b10 6
#855250000000
1!
1%
1-
12
#855260000000
0!
0%
b11 *
0-
02
b11 6
#855270000000
1!
1%
1-
12
15
#855280000000
0!
0%
b100 *
0-
02
b100 6
#855290000000
1!
1%
1-
12
#855300000000
0!
0%
b101 *
0-
02
b101 6
#855310000000
1!
1%
1-
12
#855320000000
0!
0%
b110 *
0-
02
b110 6
#855330000000
1!
1%
1-
12
#855340000000
0!
0%
b111 *
0-
02
b111 6
#855350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#855360000000
0!
0%
b0 *
0-
02
b0 6
#855370000000
1!
1%
1-
12
#855380000000
0!
0%
b1 *
0-
02
b1 6
#855390000000
1!
1%
1-
12
#855400000000
0!
0%
b10 *
0-
02
b10 6
#855410000000
1!
1%
1-
12
#855420000000
0!
0%
b11 *
0-
02
b11 6
#855430000000
1!
1%
1-
12
15
#855440000000
0!
0%
b100 *
0-
02
b100 6
#855450000000
1!
1%
1-
12
#855460000000
0!
0%
b101 *
0-
02
b101 6
#855470000000
1!
1%
1-
12
#855480000000
0!
0%
b110 *
0-
02
b110 6
#855490000000
1!
1%
1-
12
#855500000000
0!
0%
b111 *
0-
02
b111 6
#855510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#855520000000
0!
0%
b0 *
0-
02
b0 6
#855530000000
1!
1%
1-
12
#855540000000
0!
0%
b1 *
0-
02
b1 6
#855550000000
1!
1%
1-
12
#855560000000
0!
0%
b10 *
0-
02
b10 6
#855570000000
1!
1%
1-
12
#855580000000
0!
0%
b11 *
0-
02
b11 6
#855590000000
1!
1%
1-
12
15
#855600000000
0!
0%
b100 *
0-
02
b100 6
#855610000000
1!
1%
1-
12
#855620000000
0!
0%
b101 *
0-
02
b101 6
#855630000000
1!
1%
1-
12
#855640000000
0!
0%
b110 *
0-
02
b110 6
#855650000000
1!
1%
1-
12
#855660000000
0!
0%
b111 *
0-
02
b111 6
#855670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#855680000000
0!
0%
b0 *
0-
02
b0 6
#855690000000
1!
1%
1-
12
#855700000000
0!
0%
b1 *
0-
02
b1 6
#855710000000
1!
1%
1-
12
#855720000000
0!
0%
b10 *
0-
02
b10 6
#855730000000
1!
1%
1-
12
#855740000000
0!
0%
b11 *
0-
02
b11 6
#855750000000
1!
1%
1-
12
15
#855760000000
0!
0%
b100 *
0-
02
b100 6
#855770000000
1!
1%
1-
12
#855780000000
0!
0%
b101 *
0-
02
b101 6
#855790000000
1!
1%
1-
12
#855800000000
0!
0%
b110 *
0-
02
b110 6
#855810000000
1!
1%
1-
12
#855820000000
0!
0%
b111 *
0-
02
b111 6
#855830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#855840000000
0!
0%
b0 *
0-
02
b0 6
#855850000000
1!
1%
1-
12
#855860000000
0!
0%
b1 *
0-
02
b1 6
#855870000000
1!
1%
1-
12
#855880000000
0!
0%
b10 *
0-
02
b10 6
#855890000000
1!
1%
1-
12
#855900000000
0!
0%
b11 *
0-
02
b11 6
#855910000000
1!
1%
1-
12
15
#855920000000
0!
0%
b100 *
0-
02
b100 6
#855930000000
1!
1%
1-
12
#855940000000
0!
0%
b101 *
0-
02
b101 6
#855950000000
1!
1%
1-
12
#855960000000
0!
0%
b110 *
0-
02
b110 6
#855970000000
1!
1%
1-
12
#855980000000
0!
0%
b111 *
0-
02
b111 6
#855990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#856000000000
0!
0%
b0 *
0-
02
b0 6
#856010000000
1!
1%
1-
12
#856020000000
0!
0%
b1 *
0-
02
b1 6
#856030000000
1!
1%
1-
12
#856040000000
0!
0%
b10 *
0-
02
b10 6
#856050000000
1!
1%
1-
12
#856060000000
0!
0%
b11 *
0-
02
b11 6
#856070000000
1!
1%
1-
12
15
#856080000000
0!
0%
b100 *
0-
02
b100 6
#856090000000
1!
1%
1-
12
#856100000000
0!
0%
b101 *
0-
02
b101 6
#856110000000
1!
1%
1-
12
#856120000000
0!
0%
b110 *
0-
02
b110 6
#856130000000
1!
1%
1-
12
#856140000000
0!
0%
b111 *
0-
02
b111 6
#856150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#856160000000
0!
0%
b0 *
0-
02
b0 6
#856170000000
1!
1%
1-
12
#856180000000
0!
0%
b1 *
0-
02
b1 6
#856190000000
1!
1%
1-
12
#856200000000
0!
0%
b10 *
0-
02
b10 6
#856210000000
1!
1%
1-
12
#856220000000
0!
0%
b11 *
0-
02
b11 6
#856230000000
1!
1%
1-
12
15
#856240000000
0!
0%
b100 *
0-
02
b100 6
#856250000000
1!
1%
1-
12
#856260000000
0!
0%
b101 *
0-
02
b101 6
#856270000000
1!
1%
1-
12
#856280000000
0!
0%
b110 *
0-
02
b110 6
#856290000000
1!
1%
1-
12
#856300000000
0!
0%
b111 *
0-
02
b111 6
#856310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#856320000000
0!
0%
b0 *
0-
02
b0 6
#856330000000
1!
1%
1-
12
#856340000000
0!
0%
b1 *
0-
02
b1 6
#856350000000
1!
1%
1-
12
#856360000000
0!
0%
b10 *
0-
02
b10 6
#856370000000
1!
1%
1-
12
#856380000000
0!
0%
b11 *
0-
02
b11 6
#856390000000
1!
1%
1-
12
15
#856400000000
0!
0%
b100 *
0-
02
b100 6
#856410000000
1!
1%
1-
12
#856420000000
0!
0%
b101 *
0-
02
b101 6
#856430000000
1!
1%
1-
12
#856440000000
0!
0%
b110 *
0-
02
b110 6
#856450000000
1!
1%
1-
12
#856460000000
0!
0%
b111 *
0-
02
b111 6
#856470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#856480000000
0!
0%
b0 *
0-
02
b0 6
#856490000000
1!
1%
1-
12
#856500000000
0!
0%
b1 *
0-
02
b1 6
#856510000000
1!
1%
1-
12
#856520000000
0!
0%
b10 *
0-
02
b10 6
#856530000000
1!
1%
1-
12
#856540000000
0!
0%
b11 *
0-
02
b11 6
#856550000000
1!
1%
1-
12
15
#856560000000
0!
0%
b100 *
0-
02
b100 6
#856570000000
1!
1%
1-
12
#856580000000
0!
0%
b101 *
0-
02
b101 6
#856590000000
1!
1%
1-
12
#856600000000
0!
0%
b110 *
0-
02
b110 6
#856610000000
1!
1%
1-
12
#856620000000
0!
0%
b111 *
0-
02
b111 6
#856630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#856640000000
0!
0%
b0 *
0-
02
b0 6
#856650000000
1!
1%
1-
12
#856660000000
0!
0%
b1 *
0-
02
b1 6
#856670000000
1!
1%
1-
12
#856680000000
0!
0%
b10 *
0-
02
b10 6
#856690000000
1!
1%
1-
12
#856700000000
0!
0%
b11 *
0-
02
b11 6
#856710000000
1!
1%
1-
12
15
#856720000000
0!
0%
b100 *
0-
02
b100 6
#856730000000
1!
1%
1-
12
#856740000000
0!
0%
b101 *
0-
02
b101 6
#856750000000
1!
1%
1-
12
#856760000000
0!
0%
b110 *
0-
02
b110 6
#856770000000
1!
1%
1-
12
#856780000000
0!
0%
b111 *
0-
02
b111 6
#856790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#856800000000
0!
0%
b0 *
0-
02
b0 6
#856810000000
1!
1%
1-
12
#856820000000
0!
0%
b1 *
0-
02
b1 6
#856830000000
1!
1%
1-
12
#856840000000
0!
0%
b10 *
0-
02
b10 6
#856850000000
1!
1%
1-
12
#856860000000
0!
0%
b11 *
0-
02
b11 6
#856870000000
1!
1%
1-
12
15
#856880000000
0!
0%
b100 *
0-
02
b100 6
#856890000000
1!
1%
1-
12
#856900000000
0!
0%
b101 *
0-
02
b101 6
#856910000000
1!
1%
1-
12
#856920000000
0!
0%
b110 *
0-
02
b110 6
#856930000000
1!
1%
1-
12
#856940000000
0!
0%
b111 *
0-
02
b111 6
#856950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#856960000000
0!
0%
b0 *
0-
02
b0 6
#856970000000
1!
1%
1-
12
#856980000000
0!
0%
b1 *
0-
02
b1 6
#856990000000
1!
1%
1-
12
#857000000000
0!
0%
b10 *
0-
02
b10 6
#857010000000
1!
1%
1-
12
#857020000000
0!
0%
b11 *
0-
02
b11 6
#857030000000
1!
1%
1-
12
15
#857040000000
0!
0%
b100 *
0-
02
b100 6
#857050000000
1!
1%
1-
12
#857060000000
0!
0%
b101 *
0-
02
b101 6
#857070000000
1!
1%
1-
12
#857080000000
0!
0%
b110 *
0-
02
b110 6
#857090000000
1!
1%
1-
12
#857100000000
0!
0%
b111 *
0-
02
b111 6
#857110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#857120000000
0!
0%
b0 *
0-
02
b0 6
#857130000000
1!
1%
1-
12
#857140000000
0!
0%
b1 *
0-
02
b1 6
#857150000000
1!
1%
1-
12
#857160000000
0!
0%
b10 *
0-
02
b10 6
#857170000000
1!
1%
1-
12
#857180000000
0!
0%
b11 *
0-
02
b11 6
#857190000000
1!
1%
1-
12
15
#857200000000
0!
0%
b100 *
0-
02
b100 6
#857210000000
1!
1%
1-
12
#857220000000
0!
0%
b101 *
0-
02
b101 6
#857230000000
1!
1%
1-
12
#857240000000
0!
0%
b110 *
0-
02
b110 6
#857250000000
1!
1%
1-
12
#857260000000
0!
0%
b111 *
0-
02
b111 6
#857270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#857280000000
0!
0%
b0 *
0-
02
b0 6
#857290000000
1!
1%
1-
12
#857300000000
0!
0%
b1 *
0-
02
b1 6
#857310000000
1!
1%
1-
12
#857320000000
0!
0%
b10 *
0-
02
b10 6
#857330000000
1!
1%
1-
12
#857340000000
0!
0%
b11 *
0-
02
b11 6
#857350000000
1!
1%
1-
12
15
#857360000000
0!
0%
b100 *
0-
02
b100 6
#857370000000
1!
1%
1-
12
#857380000000
0!
0%
b101 *
0-
02
b101 6
#857390000000
1!
1%
1-
12
#857400000000
0!
0%
b110 *
0-
02
b110 6
#857410000000
1!
1%
1-
12
#857420000000
0!
0%
b111 *
0-
02
b111 6
#857430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#857440000000
0!
0%
b0 *
0-
02
b0 6
#857450000000
1!
1%
1-
12
#857460000000
0!
0%
b1 *
0-
02
b1 6
#857470000000
1!
1%
1-
12
#857480000000
0!
0%
b10 *
0-
02
b10 6
#857490000000
1!
1%
1-
12
#857500000000
0!
0%
b11 *
0-
02
b11 6
#857510000000
1!
1%
1-
12
15
#857520000000
0!
0%
b100 *
0-
02
b100 6
#857530000000
1!
1%
1-
12
#857540000000
0!
0%
b101 *
0-
02
b101 6
#857550000000
1!
1%
1-
12
#857560000000
0!
0%
b110 *
0-
02
b110 6
#857570000000
1!
1%
1-
12
#857580000000
0!
0%
b111 *
0-
02
b111 6
#857590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#857600000000
0!
0%
b0 *
0-
02
b0 6
#857610000000
1!
1%
1-
12
#857620000000
0!
0%
b1 *
0-
02
b1 6
#857630000000
1!
1%
1-
12
#857640000000
0!
0%
b10 *
0-
02
b10 6
#857650000000
1!
1%
1-
12
#857660000000
0!
0%
b11 *
0-
02
b11 6
#857670000000
1!
1%
1-
12
15
#857680000000
0!
0%
b100 *
0-
02
b100 6
#857690000000
1!
1%
1-
12
#857700000000
0!
0%
b101 *
0-
02
b101 6
#857710000000
1!
1%
1-
12
#857720000000
0!
0%
b110 *
0-
02
b110 6
#857730000000
1!
1%
1-
12
#857740000000
0!
0%
b111 *
0-
02
b111 6
#857750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#857760000000
0!
0%
b0 *
0-
02
b0 6
#857770000000
1!
1%
1-
12
#857780000000
0!
0%
b1 *
0-
02
b1 6
#857790000000
1!
1%
1-
12
#857800000000
0!
0%
b10 *
0-
02
b10 6
#857810000000
1!
1%
1-
12
#857820000000
0!
0%
b11 *
0-
02
b11 6
#857830000000
1!
1%
1-
12
15
#857840000000
0!
0%
b100 *
0-
02
b100 6
#857850000000
1!
1%
1-
12
#857860000000
0!
0%
b101 *
0-
02
b101 6
#857870000000
1!
1%
1-
12
#857880000000
0!
0%
b110 *
0-
02
b110 6
#857890000000
1!
1%
1-
12
#857900000000
0!
0%
b111 *
0-
02
b111 6
#857910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#857920000000
0!
0%
b0 *
0-
02
b0 6
#857930000000
1!
1%
1-
12
#857940000000
0!
0%
b1 *
0-
02
b1 6
#857950000000
1!
1%
1-
12
#857960000000
0!
0%
b10 *
0-
02
b10 6
#857970000000
1!
1%
1-
12
#857980000000
0!
0%
b11 *
0-
02
b11 6
#857990000000
1!
1%
1-
12
15
#858000000000
0!
0%
b100 *
0-
02
b100 6
#858010000000
1!
1%
1-
12
#858020000000
0!
0%
b101 *
0-
02
b101 6
#858030000000
1!
1%
1-
12
#858040000000
0!
0%
b110 *
0-
02
b110 6
#858050000000
1!
1%
1-
12
#858060000000
0!
0%
b111 *
0-
02
b111 6
#858070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#858080000000
0!
0%
b0 *
0-
02
b0 6
#858090000000
1!
1%
1-
12
#858100000000
0!
0%
b1 *
0-
02
b1 6
#858110000000
1!
1%
1-
12
#858120000000
0!
0%
b10 *
0-
02
b10 6
#858130000000
1!
1%
1-
12
#858140000000
0!
0%
b11 *
0-
02
b11 6
#858150000000
1!
1%
1-
12
15
#858160000000
0!
0%
b100 *
0-
02
b100 6
#858170000000
1!
1%
1-
12
#858180000000
0!
0%
b101 *
0-
02
b101 6
#858190000000
1!
1%
1-
12
#858200000000
0!
0%
b110 *
0-
02
b110 6
#858210000000
1!
1%
1-
12
#858220000000
0!
0%
b111 *
0-
02
b111 6
#858230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#858240000000
0!
0%
b0 *
0-
02
b0 6
#858250000000
1!
1%
1-
12
#858260000000
0!
0%
b1 *
0-
02
b1 6
#858270000000
1!
1%
1-
12
#858280000000
0!
0%
b10 *
0-
02
b10 6
#858290000000
1!
1%
1-
12
#858300000000
0!
0%
b11 *
0-
02
b11 6
#858310000000
1!
1%
1-
12
15
#858320000000
0!
0%
b100 *
0-
02
b100 6
#858330000000
1!
1%
1-
12
#858340000000
0!
0%
b101 *
0-
02
b101 6
#858350000000
1!
1%
1-
12
#858360000000
0!
0%
b110 *
0-
02
b110 6
#858370000000
1!
1%
1-
12
#858380000000
0!
0%
b111 *
0-
02
b111 6
#858390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#858400000000
0!
0%
b0 *
0-
02
b0 6
#858410000000
1!
1%
1-
12
#858420000000
0!
0%
b1 *
0-
02
b1 6
#858430000000
1!
1%
1-
12
#858440000000
0!
0%
b10 *
0-
02
b10 6
#858450000000
1!
1%
1-
12
#858460000000
0!
0%
b11 *
0-
02
b11 6
#858470000000
1!
1%
1-
12
15
#858480000000
0!
0%
b100 *
0-
02
b100 6
#858490000000
1!
1%
1-
12
#858500000000
0!
0%
b101 *
0-
02
b101 6
#858510000000
1!
1%
1-
12
#858520000000
0!
0%
b110 *
0-
02
b110 6
#858530000000
1!
1%
1-
12
#858540000000
0!
0%
b111 *
0-
02
b111 6
#858550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#858560000000
0!
0%
b0 *
0-
02
b0 6
#858570000000
1!
1%
1-
12
#858580000000
0!
0%
b1 *
0-
02
b1 6
#858590000000
1!
1%
1-
12
#858600000000
0!
0%
b10 *
0-
02
b10 6
#858610000000
1!
1%
1-
12
#858620000000
0!
0%
b11 *
0-
02
b11 6
#858630000000
1!
1%
1-
12
15
#858640000000
0!
0%
b100 *
0-
02
b100 6
#858650000000
1!
1%
1-
12
#858660000000
0!
0%
b101 *
0-
02
b101 6
#858670000000
1!
1%
1-
12
#858680000000
0!
0%
b110 *
0-
02
b110 6
#858690000000
1!
1%
1-
12
#858700000000
0!
0%
b111 *
0-
02
b111 6
#858710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#858720000000
0!
0%
b0 *
0-
02
b0 6
#858730000000
1!
1%
1-
12
#858740000000
0!
0%
b1 *
0-
02
b1 6
#858750000000
1!
1%
1-
12
#858760000000
0!
0%
b10 *
0-
02
b10 6
#858770000000
1!
1%
1-
12
#858780000000
0!
0%
b11 *
0-
02
b11 6
#858790000000
1!
1%
1-
12
15
#858800000000
0!
0%
b100 *
0-
02
b100 6
#858810000000
1!
1%
1-
12
#858820000000
0!
0%
b101 *
0-
02
b101 6
#858830000000
1!
1%
1-
12
#858840000000
0!
0%
b110 *
0-
02
b110 6
#858850000000
1!
1%
1-
12
#858860000000
0!
0%
b111 *
0-
02
b111 6
#858870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#858880000000
0!
0%
b0 *
0-
02
b0 6
#858890000000
1!
1%
1-
12
#858900000000
0!
0%
b1 *
0-
02
b1 6
#858910000000
1!
1%
1-
12
#858920000000
0!
0%
b10 *
0-
02
b10 6
#858930000000
1!
1%
1-
12
#858940000000
0!
0%
b11 *
0-
02
b11 6
#858950000000
1!
1%
1-
12
15
#858960000000
0!
0%
b100 *
0-
02
b100 6
#858970000000
1!
1%
1-
12
#858980000000
0!
0%
b101 *
0-
02
b101 6
#858990000000
1!
1%
1-
12
#859000000000
0!
0%
b110 *
0-
02
b110 6
#859010000000
1!
1%
1-
12
#859020000000
0!
0%
b111 *
0-
02
b111 6
#859030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#859040000000
0!
0%
b0 *
0-
02
b0 6
#859050000000
1!
1%
1-
12
#859060000000
0!
0%
b1 *
0-
02
b1 6
#859070000000
1!
1%
1-
12
#859080000000
0!
0%
b10 *
0-
02
b10 6
#859090000000
1!
1%
1-
12
#859100000000
0!
0%
b11 *
0-
02
b11 6
#859110000000
1!
1%
1-
12
15
#859120000000
0!
0%
b100 *
0-
02
b100 6
#859130000000
1!
1%
1-
12
#859140000000
0!
0%
b101 *
0-
02
b101 6
#859150000000
1!
1%
1-
12
#859160000000
0!
0%
b110 *
0-
02
b110 6
#859170000000
1!
1%
1-
12
#859180000000
0!
0%
b111 *
0-
02
b111 6
#859190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#859200000000
0!
0%
b0 *
0-
02
b0 6
#859210000000
1!
1%
1-
12
#859220000000
0!
0%
b1 *
0-
02
b1 6
#859230000000
1!
1%
1-
12
#859240000000
0!
0%
b10 *
0-
02
b10 6
#859250000000
1!
1%
1-
12
#859260000000
0!
0%
b11 *
0-
02
b11 6
#859270000000
1!
1%
1-
12
15
#859280000000
0!
0%
b100 *
0-
02
b100 6
#859290000000
1!
1%
1-
12
#859300000000
0!
0%
b101 *
0-
02
b101 6
#859310000000
1!
1%
1-
12
#859320000000
0!
0%
b110 *
0-
02
b110 6
#859330000000
1!
1%
1-
12
#859340000000
0!
0%
b111 *
0-
02
b111 6
#859350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#859360000000
0!
0%
b0 *
0-
02
b0 6
#859370000000
1!
1%
1-
12
#859380000000
0!
0%
b1 *
0-
02
b1 6
#859390000000
1!
1%
1-
12
#859400000000
0!
0%
b10 *
0-
02
b10 6
#859410000000
1!
1%
1-
12
#859420000000
0!
0%
b11 *
0-
02
b11 6
#859430000000
1!
1%
1-
12
15
#859440000000
0!
0%
b100 *
0-
02
b100 6
#859450000000
1!
1%
1-
12
#859460000000
0!
0%
b101 *
0-
02
b101 6
#859470000000
1!
1%
1-
12
#859480000000
0!
0%
b110 *
0-
02
b110 6
#859490000000
1!
1%
1-
12
#859500000000
0!
0%
b111 *
0-
02
b111 6
#859510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#859520000000
0!
0%
b0 *
0-
02
b0 6
#859530000000
1!
1%
1-
12
#859540000000
0!
0%
b1 *
0-
02
b1 6
#859550000000
1!
1%
1-
12
#859560000000
0!
0%
b10 *
0-
02
b10 6
#859570000000
1!
1%
1-
12
#859580000000
0!
0%
b11 *
0-
02
b11 6
#859590000000
1!
1%
1-
12
15
#859600000000
0!
0%
b100 *
0-
02
b100 6
#859610000000
1!
1%
1-
12
#859620000000
0!
0%
b101 *
0-
02
b101 6
#859630000000
1!
1%
1-
12
#859640000000
0!
0%
b110 *
0-
02
b110 6
#859650000000
1!
1%
1-
12
#859660000000
0!
0%
b111 *
0-
02
b111 6
#859670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#859680000000
0!
0%
b0 *
0-
02
b0 6
#859690000000
1!
1%
1-
12
#859700000000
0!
0%
b1 *
0-
02
b1 6
#859710000000
1!
1%
1-
12
#859720000000
0!
0%
b10 *
0-
02
b10 6
#859730000000
1!
1%
1-
12
#859740000000
0!
0%
b11 *
0-
02
b11 6
#859750000000
1!
1%
1-
12
15
#859760000000
0!
0%
b100 *
0-
02
b100 6
#859770000000
1!
1%
1-
12
#859780000000
0!
0%
b101 *
0-
02
b101 6
#859790000000
1!
1%
1-
12
#859800000000
0!
0%
b110 *
0-
02
b110 6
#859810000000
1!
1%
1-
12
#859820000000
0!
0%
b111 *
0-
02
b111 6
#859830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#859840000000
0!
0%
b0 *
0-
02
b0 6
#859850000000
1!
1%
1-
12
#859860000000
0!
0%
b1 *
0-
02
b1 6
#859870000000
1!
1%
1-
12
#859880000000
0!
0%
b10 *
0-
02
b10 6
#859890000000
1!
1%
1-
12
#859900000000
0!
0%
b11 *
0-
02
b11 6
#859910000000
1!
1%
1-
12
15
#859920000000
0!
0%
b100 *
0-
02
b100 6
#859930000000
1!
1%
1-
12
#859940000000
0!
0%
b101 *
0-
02
b101 6
#859950000000
1!
1%
1-
12
#859960000000
0!
0%
b110 *
0-
02
b110 6
#859970000000
1!
1%
1-
12
#859980000000
0!
0%
b111 *
0-
02
b111 6
#859990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#860000000000
0!
0%
b0 *
0-
02
b0 6
#860010000000
1!
1%
1-
12
#860020000000
0!
0%
b1 *
0-
02
b1 6
#860030000000
1!
1%
1-
12
#860040000000
0!
0%
b10 *
0-
02
b10 6
#860050000000
1!
1%
1-
12
#860060000000
0!
0%
b11 *
0-
02
b11 6
#860070000000
1!
1%
1-
12
15
#860080000000
0!
0%
b100 *
0-
02
b100 6
#860090000000
1!
1%
1-
12
#860100000000
0!
0%
b101 *
0-
02
b101 6
#860110000000
1!
1%
1-
12
#860120000000
0!
0%
b110 *
0-
02
b110 6
#860130000000
1!
1%
1-
12
#860140000000
0!
0%
b111 *
0-
02
b111 6
#860150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#860160000000
0!
0%
b0 *
0-
02
b0 6
#860170000000
1!
1%
1-
12
#860180000000
0!
0%
b1 *
0-
02
b1 6
#860190000000
1!
1%
1-
12
#860200000000
0!
0%
b10 *
0-
02
b10 6
#860210000000
1!
1%
1-
12
#860220000000
0!
0%
b11 *
0-
02
b11 6
#860230000000
1!
1%
1-
12
15
#860240000000
0!
0%
b100 *
0-
02
b100 6
#860250000000
1!
1%
1-
12
#860260000000
0!
0%
b101 *
0-
02
b101 6
#860270000000
1!
1%
1-
12
#860280000000
0!
0%
b110 *
0-
02
b110 6
#860290000000
1!
1%
1-
12
#860300000000
0!
0%
b111 *
0-
02
b111 6
#860310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#860320000000
0!
0%
b0 *
0-
02
b0 6
#860330000000
1!
1%
1-
12
#860340000000
0!
0%
b1 *
0-
02
b1 6
#860350000000
1!
1%
1-
12
#860360000000
0!
0%
b10 *
0-
02
b10 6
#860370000000
1!
1%
1-
12
#860380000000
0!
0%
b11 *
0-
02
b11 6
#860390000000
1!
1%
1-
12
15
#860400000000
0!
0%
b100 *
0-
02
b100 6
#860410000000
1!
1%
1-
12
#860420000000
0!
0%
b101 *
0-
02
b101 6
#860430000000
1!
1%
1-
12
#860440000000
0!
0%
b110 *
0-
02
b110 6
#860450000000
1!
1%
1-
12
#860460000000
0!
0%
b111 *
0-
02
b111 6
#860470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#860480000000
0!
0%
b0 *
0-
02
b0 6
#860490000000
1!
1%
1-
12
#860500000000
0!
0%
b1 *
0-
02
b1 6
#860510000000
1!
1%
1-
12
#860520000000
0!
0%
b10 *
0-
02
b10 6
#860530000000
1!
1%
1-
12
#860540000000
0!
0%
b11 *
0-
02
b11 6
#860550000000
1!
1%
1-
12
15
#860560000000
0!
0%
b100 *
0-
02
b100 6
#860570000000
1!
1%
1-
12
#860580000000
0!
0%
b101 *
0-
02
b101 6
#860590000000
1!
1%
1-
12
#860600000000
0!
0%
b110 *
0-
02
b110 6
#860610000000
1!
1%
1-
12
#860620000000
0!
0%
b111 *
0-
02
b111 6
#860630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#860640000000
0!
0%
b0 *
0-
02
b0 6
#860650000000
1!
1%
1-
12
#860660000000
0!
0%
b1 *
0-
02
b1 6
#860670000000
1!
1%
1-
12
#860680000000
0!
0%
b10 *
0-
02
b10 6
#860690000000
1!
1%
1-
12
#860700000000
0!
0%
b11 *
0-
02
b11 6
#860710000000
1!
1%
1-
12
15
#860720000000
0!
0%
b100 *
0-
02
b100 6
#860730000000
1!
1%
1-
12
#860740000000
0!
0%
b101 *
0-
02
b101 6
#860750000000
1!
1%
1-
12
#860760000000
0!
0%
b110 *
0-
02
b110 6
#860770000000
1!
1%
1-
12
#860780000000
0!
0%
b111 *
0-
02
b111 6
#860790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#860800000000
0!
0%
b0 *
0-
02
b0 6
#860810000000
1!
1%
1-
12
#860820000000
0!
0%
b1 *
0-
02
b1 6
#860830000000
1!
1%
1-
12
#860840000000
0!
0%
b10 *
0-
02
b10 6
#860850000000
1!
1%
1-
12
#860860000000
0!
0%
b11 *
0-
02
b11 6
#860870000000
1!
1%
1-
12
15
#860880000000
0!
0%
b100 *
0-
02
b100 6
#860890000000
1!
1%
1-
12
#860900000000
0!
0%
b101 *
0-
02
b101 6
#860910000000
1!
1%
1-
12
#860920000000
0!
0%
b110 *
0-
02
b110 6
#860930000000
1!
1%
1-
12
#860940000000
0!
0%
b111 *
0-
02
b111 6
#860950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#860960000000
0!
0%
b0 *
0-
02
b0 6
#860970000000
1!
1%
1-
12
#860980000000
0!
0%
b1 *
0-
02
b1 6
#860990000000
1!
1%
1-
12
#861000000000
0!
0%
b10 *
0-
02
b10 6
#861010000000
1!
1%
1-
12
#861020000000
0!
0%
b11 *
0-
02
b11 6
#861030000000
1!
1%
1-
12
15
#861040000000
0!
0%
b100 *
0-
02
b100 6
#861050000000
1!
1%
1-
12
#861060000000
0!
0%
b101 *
0-
02
b101 6
#861070000000
1!
1%
1-
12
#861080000000
0!
0%
b110 *
0-
02
b110 6
#861090000000
1!
1%
1-
12
#861100000000
0!
0%
b111 *
0-
02
b111 6
#861110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#861120000000
0!
0%
b0 *
0-
02
b0 6
#861130000000
1!
1%
1-
12
#861140000000
0!
0%
b1 *
0-
02
b1 6
#861150000000
1!
1%
1-
12
#861160000000
0!
0%
b10 *
0-
02
b10 6
#861170000000
1!
1%
1-
12
#861180000000
0!
0%
b11 *
0-
02
b11 6
#861190000000
1!
1%
1-
12
15
#861200000000
0!
0%
b100 *
0-
02
b100 6
#861210000000
1!
1%
1-
12
#861220000000
0!
0%
b101 *
0-
02
b101 6
#861230000000
1!
1%
1-
12
#861240000000
0!
0%
b110 *
0-
02
b110 6
#861250000000
1!
1%
1-
12
#861260000000
0!
0%
b111 *
0-
02
b111 6
#861270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#861280000000
0!
0%
b0 *
0-
02
b0 6
#861290000000
1!
1%
1-
12
#861300000000
0!
0%
b1 *
0-
02
b1 6
#861310000000
1!
1%
1-
12
#861320000000
0!
0%
b10 *
0-
02
b10 6
#861330000000
1!
1%
1-
12
#861340000000
0!
0%
b11 *
0-
02
b11 6
#861350000000
1!
1%
1-
12
15
#861360000000
0!
0%
b100 *
0-
02
b100 6
#861370000000
1!
1%
1-
12
#861380000000
0!
0%
b101 *
0-
02
b101 6
#861390000000
1!
1%
1-
12
#861400000000
0!
0%
b110 *
0-
02
b110 6
#861410000000
1!
1%
1-
12
#861420000000
0!
0%
b111 *
0-
02
b111 6
#861430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#861440000000
0!
0%
b0 *
0-
02
b0 6
#861450000000
1!
1%
1-
12
#861460000000
0!
0%
b1 *
0-
02
b1 6
#861470000000
1!
1%
1-
12
#861480000000
0!
0%
b10 *
0-
02
b10 6
#861490000000
1!
1%
1-
12
#861500000000
0!
0%
b11 *
0-
02
b11 6
#861510000000
1!
1%
1-
12
15
#861520000000
0!
0%
b100 *
0-
02
b100 6
#861530000000
1!
1%
1-
12
#861540000000
0!
0%
b101 *
0-
02
b101 6
#861550000000
1!
1%
1-
12
#861560000000
0!
0%
b110 *
0-
02
b110 6
#861570000000
1!
1%
1-
12
#861580000000
0!
0%
b111 *
0-
02
b111 6
#861590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#861600000000
0!
0%
b0 *
0-
02
b0 6
#861610000000
1!
1%
1-
12
#861620000000
0!
0%
b1 *
0-
02
b1 6
#861630000000
1!
1%
1-
12
#861640000000
0!
0%
b10 *
0-
02
b10 6
#861650000000
1!
1%
1-
12
#861660000000
0!
0%
b11 *
0-
02
b11 6
#861670000000
1!
1%
1-
12
15
#861680000000
0!
0%
b100 *
0-
02
b100 6
#861690000000
1!
1%
1-
12
#861700000000
0!
0%
b101 *
0-
02
b101 6
#861710000000
1!
1%
1-
12
#861720000000
0!
0%
b110 *
0-
02
b110 6
#861730000000
1!
1%
1-
12
#861740000000
0!
0%
b111 *
0-
02
b111 6
#861750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#861760000000
0!
0%
b0 *
0-
02
b0 6
#861770000000
1!
1%
1-
12
#861780000000
0!
0%
b1 *
0-
02
b1 6
#861790000000
1!
1%
1-
12
#861800000000
0!
0%
b10 *
0-
02
b10 6
#861810000000
1!
1%
1-
12
#861820000000
0!
0%
b11 *
0-
02
b11 6
#861830000000
1!
1%
1-
12
15
#861840000000
0!
0%
b100 *
0-
02
b100 6
#861850000000
1!
1%
1-
12
#861860000000
0!
0%
b101 *
0-
02
b101 6
#861870000000
1!
1%
1-
12
#861880000000
0!
0%
b110 *
0-
02
b110 6
#861890000000
1!
1%
1-
12
#861900000000
0!
0%
b111 *
0-
02
b111 6
#861910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#861920000000
0!
0%
b0 *
0-
02
b0 6
#861930000000
1!
1%
1-
12
#861940000000
0!
0%
b1 *
0-
02
b1 6
#861950000000
1!
1%
1-
12
#861960000000
0!
0%
b10 *
0-
02
b10 6
#861970000000
1!
1%
1-
12
#861980000000
0!
0%
b11 *
0-
02
b11 6
#861990000000
1!
1%
1-
12
15
#862000000000
0!
0%
b100 *
0-
02
b100 6
#862010000000
1!
1%
1-
12
#862020000000
0!
0%
b101 *
0-
02
b101 6
#862030000000
1!
1%
1-
12
#862040000000
0!
0%
b110 *
0-
02
b110 6
#862050000000
1!
1%
1-
12
#862060000000
0!
0%
b111 *
0-
02
b111 6
#862070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#862080000000
0!
0%
b0 *
0-
02
b0 6
#862090000000
1!
1%
1-
12
#862100000000
0!
0%
b1 *
0-
02
b1 6
#862110000000
1!
1%
1-
12
#862120000000
0!
0%
b10 *
0-
02
b10 6
#862130000000
1!
1%
1-
12
#862140000000
0!
0%
b11 *
0-
02
b11 6
#862150000000
1!
1%
1-
12
15
#862160000000
0!
0%
b100 *
0-
02
b100 6
#862170000000
1!
1%
1-
12
#862180000000
0!
0%
b101 *
0-
02
b101 6
#862190000000
1!
1%
1-
12
#862200000000
0!
0%
b110 *
0-
02
b110 6
#862210000000
1!
1%
1-
12
#862220000000
0!
0%
b111 *
0-
02
b111 6
#862230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#862240000000
0!
0%
b0 *
0-
02
b0 6
#862250000000
1!
1%
1-
12
#862260000000
0!
0%
b1 *
0-
02
b1 6
#862270000000
1!
1%
1-
12
#862280000000
0!
0%
b10 *
0-
02
b10 6
#862290000000
1!
1%
1-
12
#862300000000
0!
0%
b11 *
0-
02
b11 6
#862310000000
1!
1%
1-
12
15
#862320000000
0!
0%
b100 *
0-
02
b100 6
#862330000000
1!
1%
1-
12
#862340000000
0!
0%
b101 *
0-
02
b101 6
#862350000000
1!
1%
1-
12
#862360000000
0!
0%
b110 *
0-
02
b110 6
#862370000000
1!
1%
1-
12
#862380000000
0!
0%
b111 *
0-
02
b111 6
#862390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#862400000000
0!
0%
b0 *
0-
02
b0 6
#862410000000
1!
1%
1-
12
#862420000000
0!
0%
b1 *
0-
02
b1 6
#862430000000
1!
1%
1-
12
#862440000000
0!
0%
b10 *
0-
02
b10 6
#862450000000
1!
1%
1-
12
#862460000000
0!
0%
b11 *
0-
02
b11 6
#862470000000
1!
1%
1-
12
15
#862480000000
0!
0%
b100 *
0-
02
b100 6
#862490000000
1!
1%
1-
12
#862500000000
0!
0%
b101 *
0-
02
b101 6
#862510000000
1!
1%
1-
12
#862520000000
0!
0%
b110 *
0-
02
b110 6
#862530000000
1!
1%
1-
12
#862540000000
0!
0%
b111 *
0-
02
b111 6
#862550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#862560000000
0!
0%
b0 *
0-
02
b0 6
#862570000000
1!
1%
1-
12
#862580000000
0!
0%
b1 *
0-
02
b1 6
#862590000000
1!
1%
1-
12
#862600000000
0!
0%
b10 *
0-
02
b10 6
#862610000000
1!
1%
1-
12
#862620000000
0!
0%
b11 *
0-
02
b11 6
#862630000000
1!
1%
1-
12
15
#862640000000
0!
0%
b100 *
0-
02
b100 6
#862650000000
1!
1%
1-
12
#862660000000
0!
0%
b101 *
0-
02
b101 6
#862670000000
1!
1%
1-
12
#862680000000
0!
0%
b110 *
0-
02
b110 6
#862690000000
1!
1%
1-
12
#862700000000
0!
0%
b111 *
0-
02
b111 6
#862710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#862720000000
0!
0%
b0 *
0-
02
b0 6
#862730000000
1!
1%
1-
12
#862740000000
0!
0%
b1 *
0-
02
b1 6
#862750000000
1!
1%
1-
12
#862760000000
0!
0%
b10 *
0-
02
b10 6
#862770000000
1!
1%
1-
12
#862780000000
0!
0%
b11 *
0-
02
b11 6
#862790000000
1!
1%
1-
12
15
#862800000000
0!
0%
b100 *
0-
02
b100 6
#862810000000
1!
1%
1-
12
#862820000000
0!
0%
b101 *
0-
02
b101 6
#862830000000
1!
1%
1-
12
#862840000000
0!
0%
b110 *
0-
02
b110 6
#862850000000
1!
1%
1-
12
#862860000000
0!
0%
b111 *
0-
02
b111 6
#862870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#862880000000
0!
0%
b0 *
0-
02
b0 6
#862890000000
1!
1%
1-
12
#862900000000
0!
0%
b1 *
0-
02
b1 6
#862910000000
1!
1%
1-
12
#862920000000
0!
0%
b10 *
0-
02
b10 6
#862930000000
1!
1%
1-
12
#862940000000
0!
0%
b11 *
0-
02
b11 6
#862950000000
1!
1%
1-
12
15
#862960000000
0!
0%
b100 *
0-
02
b100 6
#862970000000
1!
1%
1-
12
#862980000000
0!
0%
b101 *
0-
02
b101 6
#862990000000
1!
1%
1-
12
#863000000000
0!
0%
b110 *
0-
02
b110 6
#863010000000
1!
1%
1-
12
#863020000000
0!
0%
b111 *
0-
02
b111 6
#863030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#863040000000
0!
0%
b0 *
0-
02
b0 6
#863050000000
1!
1%
1-
12
#863060000000
0!
0%
b1 *
0-
02
b1 6
#863070000000
1!
1%
1-
12
#863080000000
0!
0%
b10 *
0-
02
b10 6
#863090000000
1!
1%
1-
12
#863100000000
0!
0%
b11 *
0-
02
b11 6
#863110000000
1!
1%
1-
12
15
#863120000000
0!
0%
b100 *
0-
02
b100 6
#863130000000
1!
1%
1-
12
#863140000000
0!
0%
b101 *
0-
02
b101 6
#863150000000
1!
1%
1-
12
#863160000000
0!
0%
b110 *
0-
02
b110 6
#863170000000
1!
1%
1-
12
#863180000000
0!
0%
b111 *
0-
02
b111 6
#863190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#863200000000
0!
0%
b0 *
0-
02
b0 6
#863210000000
1!
1%
1-
12
#863220000000
0!
0%
b1 *
0-
02
b1 6
#863230000000
1!
1%
1-
12
#863240000000
0!
0%
b10 *
0-
02
b10 6
#863250000000
1!
1%
1-
12
#863260000000
0!
0%
b11 *
0-
02
b11 6
#863270000000
1!
1%
1-
12
15
#863280000000
0!
0%
b100 *
0-
02
b100 6
#863290000000
1!
1%
1-
12
#863300000000
0!
0%
b101 *
0-
02
b101 6
#863310000000
1!
1%
1-
12
#863320000000
0!
0%
b110 *
0-
02
b110 6
#863330000000
1!
1%
1-
12
#863340000000
0!
0%
b111 *
0-
02
b111 6
#863350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#863360000000
0!
0%
b0 *
0-
02
b0 6
#863370000000
1!
1%
1-
12
#863380000000
0!
0%
b1 *
0-
02
b1 6
#863390000000
1!
1%
1-
12
#863400000000
0!
0%
b10 *
0-
02
b10 6
#863410000000
1!
1%
1-
12
#863420000000
0!
0%
b11 *
0-
02
b11 6
#863430000000
1!
1%
1-
12
15
#863440000000
0!
0%
b100 *
0-
02
b100 6
#863450000000
1!
1%
1-
12
#863460000000
0!
0%
b101 *
0-
02
b101 6
#863470000000
1!
1%
1-
12
#863480000000
0!
0%
b110 *
0-
02
b110 6
#863490000000
1!
1%
1-
12
#863500000000
0!
0%
b111 *
0-
02
b111 6
#863510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#863520000000
0!
0%
b0 *
0-
02
b0 6
#863530000000
1!
1%
1-
12
#863540000000
0!
0%
b1 *
0-
02
b1 6
#863550000000
1!
1%
1-
12
#863560000000
0!
0%
b10 *
0-
02
b10 6
#863570000000
1!
1%
1-
12
#863580000000
0!
0%
b11 *
0-
02
b11 6
#863590000000
1!
1%
1-
12
15
#863600000000
0!
0%
b100 *
0-
02
b100 6
#863610000000
1!
1%
1-
12
#863620000000
0!
0%
b101 *
0-
02
b101 6
#863630000000
1!
1%
1-
12
#863640000000
0!
0%
b110 *
0-
02
b110 6
#863650000000
1!
1%
1-
12
#863660000000
0!
0%
b111 *
0-
02
b111 6
#863670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#863680000000
0!
0%
b0 *
0-
02
b0 6
#863690000000
1!
1%
1-
12
#863700000000
0!
0%
b1 *
0-
02
b1 6
#863710000000
1!
1%
1-
12
#863720000000
0!
0%
b10 *
0-
02
b10 6
#863730000000
1!
1%
1-
12
#863740000000
0!
0%
b11 *
0-
02
b11 6
#863750000000
1!
1%
1-
12
15
#863760000000
0!
0%
b100 *
0-
02
b100 6
#863770000000
1!
1%
1-
12
#863780000000
0!
0%
b101 *
0-
02
b101 6
#863790000000
1!
1%
1-
12
#863800000000
0!
0%
b110 *
0-
02
b110 6
#863810000000
1!
1%
1-
12
#863820000000
0!
0%
b111 *
0-
02
b111 6
#863830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#863840000000
0!
0%
b0 *
0-
02
b0 6
#863850000000
1!
1%
1-
12
#863860000000
0!
0%
b1 *
0-
02
b1 6
#863870000000
1!
1%
1-
12
#863880000000
0!
0%
b10 *
0-
02
b10 6
#863890000000
1!
1%
1-
12
#863900000000
0!
0%
b11 *
0-
02
b11 6
#863910000000
1!
1%
1-
12
15
#863920000000
0!
0%
b100 *
0-
02
b100 6
#863930000000
1!
1%
1-
12
#863940000000
0!
0%
b101 *
0-
02
b101 6
#863950000000
1!
1%
1-
12
#863960000000
0!
0%
b110 *
0-
02
b110 6
#863970000000
1!
1%
1-
12
#863980000000
0!
0%
b111 *
0-
02
b111 6
#863990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#864000000000
0!
0%
b0 *
0-
02
b0 6
#864010000000
1!
1%
1-
12
#864020000000
0!
0%
b1 *
0-
02
b1 6
#864030000000
1!
1%
1-
12
#864040000000
0!
0%
b10 *
0-
02
b10 6
#864050000000
1!
1%
1-
12
#864060000000
0!
0%
b11 *
0-
02
b11 6
#864070000000
1!
1%
1-
12
15
#864080000000
0!
0%
b100 *
0-
02
b100 6
#864090000000
1!
1%
1-
12
#864100000000
0!
0%
b101 *
0-
02
b101 6
#864110000000
1!
1%
1-
12
#864120000000
0!
0%
b110 *
0-
02
b110 6
#864130000000
1!
1%
1-
12
#864140000000
0!
0%
b111 *
0-
02
b111 6
#864150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#864160000000
0!
0%
b0 *
0-
02
b0 6
#864170000000
1!
1%
1-
12
#864180000000
0!
0%
b1 *
0-
02
b1 6
#864190000000
1!
1%
1-
12
#864200000000
0!
0%
b10 *
0-
02
b10 6
#864210000000
1!
1%
1-
12
#864220000000
0!
0%
b11 *
0-
02
b11 6
#864230000000
1!
1%
1-
12
15
#864240000000
0!
0%
b100 *
0-
02
b100 6
#864250000000
1!
1%
1-
12
#864260000000
0!
0%
b101 *
0-
02
b101 6
#864270000000
1!
1%
1-
12
#864280000000
0!
0%
b110 *
0-
02
b110 6
#864290000000
1!
1%
1-
12
#864300000000
0!
0%
b111 *
0-
02
b111 6
#864310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#864320000000
0!
0%
b0 *
0-
02
b0 6
#864330000000
1!
1%
1-
12
#864340000000
0!
0%
b1 *
0-
02
b1 6
#864350000000
1!
1%
1-
12
#864360000000
0!
0%
b10 *
0-
02
b10 6
#864370000000
1!
1%
1-
12
#864380000000
0!
0%
b11 *
0-
02
b11 6
#864390000000
1!
1%
1-
12
15
#864400000000
0!
0%
b100 *
0-
02
b100 6
#864410000000
1!
1%
1-
12
#864420000000
0!
0%
b101 *
0-
02
b101 6
#864430000000
1!
1%
1-
12
#864440000000
0!
0%
b110 *
0-
02
b110 6
#864450000000
1!
1%
1-
12
#864460000000
0!
0%
b111 *
0-
02
b111 6
#864470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#864480000000
0!
0%
b0 *
0-
02
b0 6
#864490000000
1!
1%
1-
12
#864500000000
0!
0%
b1 *
0-
02
b1 6
#864510000000
1!
1%
1-
12
#864520000000
0!
0%
b10 *
0-
02
b10 6
#864530000000
1!
1%
1-
12
#864540000000
0!
0%
b11 *
0-
02
b11 6
#864550000000
1!
1%
1-
12
15
#864560000000
0!
0%
b100 *
0-
02
b100 6
#864570000000
1!
1%
1-
12
#864580000000
0!
0%
b101 *
0-
02
b101 6
#864590000000
1!
1%
1-
12
#864600000000
0!
0%
b110 *
0-
02
b110 6
#864610000000
1!
1%
1-
12
#864620000000
0!
0%
b111 *
0-
02
b111 6
#864630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#864640000000
0!
0%
b0 *
0-
02
b0 6
#864650000000
1!
1%
1-
12
#864660000000
0!
0%
b1 *
0-
02
b1 6
#864670000000
1!
1%
1-
12
#864680000000
0!
0%
b10 *
0-
02
b10 6
#864690000000
1!
1%
1-
12
#864700000000
0!
0%
b11 *
0-
02
b11 6
#864710000000
1!
1%
1-
12
15
#864720000000
0!
0%
b100 *
0-
02
b100 6
#864730000000
1!
1%
1-
12
#864740000000
0!
0%
b101 *
0-
02
b101 6
#864750000000
1!
1%
1-
12
#864760000000
0!
0%
b110 *
0-
02
b110 6
#864770000000
1!
1%
1-
12
#864780000000
0!
0%
b111 *
0-
02
b111 6
#864790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#864800000000
0!
0%
b0 *
0-
02
b0 6
#864810000000
1!
1%
1-
12
#864820000000
0!
0%
b1 *
0-
02
b1 6
#864830000000
1!
1%
1-
12
#864840000000
0!
0%
b10 *
0-
02
b10 6
#864850000000
1!
1%
1-
12
#864860000000
0!
0%
b11 *
0-
02
b11 6
#864870000000
1!
1%
1-
12
15
#864880000000
0!
0%
b100 *
0-
02
b100 6
#864890000000
1!
1%
1-
12
#864900000000
0!
0%
b101 *
0-
02
b101 6
#864910000000
1!
1%
1-
12
#864920000000
0!
0%
b110 *
0-
02
b110 6
#864930000000
1!
1%
1-
12
#864940000000
0!
0%
b111 *
0-
02
b111 6
#864950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#864960000000
0!
0%
b0 *
0-
02
b0 6
#864970000000
1!
1%
1-
12
#864980000000
0!
0%
b1 *
0-
02
b1 6
#864990000000
1!
1%
1-
12
#865000000000
0!
0%
b10 *
0-
02
b10 6
#865010000000
1!
1%
1-
12
#865020000000
0!
0%
b11 *
0-
02
b11 6
#865030000000
1!
1%
1-
12
15
#865040000000
0!
0%
b100 *
0-
02
b100 6
#865050000000
1!
1%
1-
12
#865060000000
0!
0%
b101 *
0-
02
b101 6
#865070000000
1!
1%
1-
12
#865080000000
0!
0%
b110 *
0-
02
b110 6
#865090000000
1!
1%
1-
12
#865100000000
0!
0%
b111 *
0-
02
b111 6
#865110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#865120000000
0!
0%
b0 *
0-
02
b0 6
#865130000000
1!
1%
1-
12
#865140000000
0!
0%
b1 *
0-
02
b1 6
#865150000000
1!
1%
1-
12
#865160000000
0!
0%
b10 *
0-
02
b10 6
#865170000000
1!
1%
1-
12
#865180000000
0!
0%
b11 *
0-
02
b11 6
#865190000000
1!
1%
1-
12
15
#865200000000
0!
0%
b100 *
0-
02
b100 6
#865210000000
1!
1%
1-
12
#865220000000
0!
0%
b101 *
0-
02
b101 6
#865230000000
1!
1%
1-
12
#865240000000
0!
0%
b110 *
0-
02
b110 6
#865250000000
1!
1%
1-
12
#865260000000
0!
0%
b111 *
0-
02
b111 6
#865270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#865280000000
0!
0%
b0 *
0-
02
b0 6
#865290000000
1!
1%
1-
12
#865300000000
0!
0%
b1 *
0-
02
b1 6
#865310000000
1!
1%
1-
12
#865320000000
0!
0%
b10 *
0-
02
b10 6
#865330000000
1!
1%
1-
12
#865340000000
0!
0%
b11 *
0-
02
b11 6
#865350000000
1!
1%
1-
12
15
#865360000000
0!
0%
b100 *
0-
02
b100 6
#865370000000
1!
1%
1-
12
#865380000000
0!
0%
b101 *
0-
02
b101 6
#865390000000
1!
1%
1-
12
#865400000000
0!
0%
b110 *
0-
02
b110 6
#865410000000
1!
1%
1-
12
#865420000000
0!
0%
b111 *
0-
02
b111 6
#865430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#865440000000
0!
0%
b0 *
0-
02
b0 6
#865450000000
1!
1%
1-
12
#865460000000
0!
0%
b1 *
0-
02
b1 6
#865470000000
1!
1%
1-
12
#865480000000
0!
0%
b10 *
0-
02
b10 6
#865490000000
1!
1%
1-
12
#865500000000
0!
0%
b11 *
0-
02
b11 6
#865510000000
1!
1%
1-
12
15
#865520000000
0!
0%
b100 *
0-
02
b100 6
#865530000000
1!
1%
1-
12
#865540000000
0!
0%
b101 *
0-
02
b101 6
#865550000000
1!
1%
1-
12
#865560000000
0!
0%
b110 *
0-
02
b110 6
#865570000000
1!
1%
1-
12
#865580000000
0!
0%
b111 *
0-
02
b111 6
#865590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#865600000000
0!
0%
b0 *
0-
02
b0 6
#865610000000
1!
1%
1-
12
#865620000000
0!
0%
b1 *
0-
02
b1 6
#865630000000
1!
1%
1-
12
#865640000000
0!
0%
b10 *
0-
02
b10 6
#865650000000
1!
1%
1-
12
#865660000000
0!
0%
b11 *
0-
02
b11 6
#865670000000
1!
1%
1-
12
15
#865680000000
0!
0%
b100 *
0-
02
b100 6
#865690000000
1!
1%
1-
12
#865700000000
0!
0%
b101 *
0-
02
b101 6
#865710000000
1!
1%
1-
12
#865720000000
0!
0%
b110 *
0-
02
b110 6
#865730000000
1!
1%
1-
12
#865740000000
0!
0%
b111 *
0-
02
b111 6
#865750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#865760000000
0!
0%
b0 *
0-
02
b0 6
#865770000000
1!
1%
1-
12
#865780000000
0!
0%
b1 *
0-
02
b1 6
#865790000000
1!
1%
1-
12
#865800000000
0!
0%
b10 *
0-
02
b10 6
#865810000000
1!
1%
1-
12
#865820000000
0!
0%
b11 *
0-
02
b11 6
#865830000000
1!
1%
1-
12
15
#865840000000
0!
0%
b100 *
0-
02
b100 6
#865850000000
1!
1%
1-
12
#865860000000
0!
0%
b101 *
0-
02
b101 6
#865870000000
1!
1%
1-
12
#865880000000
0!
0%
b110 *
0-
02
b110 6
#865890000000
1!
1%
1-
12
#865900000000
0!
0%
b111 *
0-
02
b111 6
#865910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#865920000000
0!
0%
b0 *
0-
02
b0 6
#865930000000
1!
1%
1-
12
#865940000000
0!
0%
b1 *
0-
02
b1 6
#865950000000
1!
1%
1-
12
#865960000000
0!
0%
b10 *
0-
02
b10 6
#865970000000
1!
1%
1-
12
#865980000000
0!
0%
b11 *
0-
02
b11 6
#865990000000
1!
1%
1-
12
15
#866000000000
0!
0%
b100 *
0-
02
b100 6
#866010000000
1!
1%
1-
12
#866020000000
0!
0%
b101 *
0-
02
b101 6
#866030000000
1!
1%
1-
12
#866040000000
0!
0%
b110 *
0-
02
b110 6
#866050000000
1!
1%
1-
12
#866060000000
0!
0%
b111 *
0-
02
b111 6
#866070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#866080000000
0!
0%
b0 *
0-
02
b0 6
#866090000000
1!
1%
1-
12
#866100000000
0!
0%
b1 *
0-
02
b1 6
#866110000000
1!
1%
1-
12
#866120000000
0!
0%
b10 *
0-
02
b10 6
#866130000000
1!
1%
1-
12
#866140000000
0!
0%
b11 *
0-
02
b11 6
#866150000000
1!
1%
1-
12
15
#866160000000
0!
0%
b100 *
0-
02
b100 6
#866170000000
1!
1%
1-
12
#866180000000
0!
0%
b101 *
0-
02
b101 6
#866190000000
1!
1%
1-
12
#866200000000
0!
0%
b110 *
0-
02
b110 6
#866210000000
1!
1%
1-
12
#866220000000
0!
0%
b111 *
0-
02
b111 6
#866230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#866240000000
0!
0%
b0 *
0-
02
b0 6
#866250000000
1!
1%
1-
12
#866260000000
0!
0%
b1 *
0-
02
b1 6
#866270000000
1!
1%
1-
12
#866280000000
0!
0%
b10 *
0-
02
b10 6
#866290000000
1!
1%
1-
12
#866300000000
0!
0%
b11 *
0-
02
b11 6
#866310000000
1!
1%
1-
12
15
#866320000000
0!
0%
b100 *
0-
02
b100 6
#866330000000
1!
1%
1-
12
#866340000000
0!
0%
b101 *
0-
02
b101 6
#866350000000
1!
1%
1-
12
#866360000000
0!
0%
b110 *
0-
02
b110 6
#866370000000
1!
1%
1-
12
#866380000000
0!
0%
b111 *
0-
02
b111 6
#866390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#866400000000
0!
0%
b0 *
0-
02
b0 6
#866410000000
1!
1%
1-
12
#866420000000
0!
0%
b1 *
0-
02
b1 6
#866430000000
1!
1%
1-
12
#866440000000
0!
0%
b10 *
0-
02
b10 6
#866450000000
1!
1%
1-
12
#866460000000
0!
0%
b11 *
0-
02
b11 6
#866470000000
1!
1%
1-
12
15
#866480000000
0!
0%
b100 *
0-
02
b100 6
#866490000000
1!
1%
1-
12
#866500000000
0!
0%
b101 *
0-
02
b101 6
#866510000000
1!
1%
1-
12
#866520000000
0!
0%
b110 *
0-
02
b110 6
#866530000000
1!
1%
1-
12
#866540000000
0!
0%
b111 *
0-
02
b111 6
#866550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#866560000000
0!
0%
b0 *
0-
02
b0 6
#866570000000
1!
1%
1-
12
#866580000000
0!
0%
b1 *
0-
02
b1 6
#866590000000
1!
1%
1-
12
#866600000000
0!
0%
b10 *
0-
02
b10 6
#866610000000
1!
1%
1-
12
#866620000000
0!
0%
b11 *
0-
02
b11 6
#866630000000
1!
1%
1-
12
15
#866640000000
0!
0%
b100 *
0-
02
b100 6
#866650000000
1!
1%
1-
12
#866660000000
0!
0%
b101 *
0-
02
b101 6
#866670000000
1!
1%
1-
12
#866680000000
0!
0%
b110 *
0-
02
b110 6
#866690000000
1!
1%
1-
12
#866700000000
0!
0%
b111 *
0-
02
b111 6
#866710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#866720000000
0!
0%
b0 *
0-
02
b0 6
#866730000000
1!
1%
1-
12
#866740000000
0!
0%
b1 *
0-
02
b1 6
#866750000000
1!
1%
1-
12
#866760000000
0!
0%
b10 *
0-
02
b10 6
#866770000000
1!
1%
1-
12
#866780000000
0!
0%
b11 *
0-
02
b11 6
#866790000000
1!
1%
1-
12
15
#866800000000
0!
0%
b100 *
0-
02
b100 6
#866810000000
1!
1%
1-
12
#866820000000
0!
0%
b101 *
0-
02
b101 6
#866830000000
1!
1%
1-
12
#866840000000
0!
0%
b110 *
0-
02
b110 6
#866850000000
1!
1%
1-
12
#866860000000
0!
0%
b111 *
0-
02
b111 6
#866870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#866880000000
0!
0%
b0 *
0-
02
b0 6
#866890000000
1!
1%
1-
12
#866900000000
0!
0%
b1 *
0-
02
b1 6
#866910000000
1!
1%
1-
12
#866920000000
0!
0%
b10 *
0-
02
b10 6
#866930000000
1!
1%
1-
12
#866940000000
0!
0%
b11 *
0-
02
b11 6
#866950000000
1!
1%
1-
12
15
#866960000000
0!
0%
b100 *
0-
02
b100 6
#866970000000
1!
1%
1-
12
#866980000000
0!
0%
b101 *
0-
02
b101 6
#866990000000
1!
1%
1-
12
#867000000000
0!
0%
b110 *
0-
02
b110 6
#867010000000
1!
1%
1-
12
#867020000000
0!
0%
b111 *
0-
02
b111 6
#867030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#867040000000
0!
0%
b0 *
0-
02
b0 6
#867050000000
1!
1%
1-
12
#867060000000
0!
0%
b1 *
0-
02
b1 6
#867070000000
1!
1%
1-
12
#867080000000
0!
0%
b10 *
0-
02
b10 6
#867090000000
1!
1%
1-
12
#867100000000
0!
0%
b11 *
0-
02
b11 6
#867110000000
1!
1%
1-
12
15
#867120000000
0!
0%
b100 *
0-
02
b100 6
#867130000000
1!
1%
1-
12
#867140000000
0!
0%
b101 *
0-
02
b101 6
#867150000000
1!
1%
1-
12
#867160000000
0!
0%
b110 *
0-
02
b110 6
#867170000000
1!
1%
1-
12
#867180000000
0!
0%
b111 *
0-
02
b111 6
#867190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#867200000000
0!
0%
b0 *
0-
02
b0 6
#867210000000
1!
1%
1-
12
#867220000000
0!
0%
b1 *
0-
02
b1 6
#867230000000
1!
1%
1-
12
#867240000000
0!
0%
b10 *
0-
02
b10 6
#867250000000
1!
1%
1-
12
#867260000000
0!
0%
b11 *
0-
02
b11 6
#867270000000
1!
1%
1-
12
15
#867280000000
0!
0%
b100 *
0-
02
b100 6
#867290000000
1!
1%
1-
12
#867300000000
0!
0%
b101 *
0-
02
b101 6
#867310000000
1!
1%
1-
12
#867320000000
0!
0%
b110 *
0-
02
b110 6
#867330000000
1!
1%
1-
12
#867340000000
0!
0%
b111 *
0-
02
b111 6
#867350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#867360000000
0!
0%
b0 *
0-
02
b0 6
#867370000000
1!
1%
1-
12
#867380000000
0!
0%
b1 *
0-
02
b1 6
#867390000000
1!
1%
1-
12
#867400000000
0!
0%
b10 *
0-
02
b10 6
#867410000000
1!
1%
1-
12
#867420000000
0!
0%
b11 *
0-
02
b11 6
#867430000000
1!
1%
1-
12
15
#867440000000
0!
0%
b100 *
0-
02
b100 6
#867450000000
1!
1%
1-
12
#867460000000
0!
0%
b101 *
0-
02
b101 6
#867470000000
1!
1%
1-
12
#867480000000
0!
0%
b110 *
0-
02
b110 6
#867490000000
1!
1%
1-
12
#867500000000
0!
0%
b111 *
0-
02
b111 6
#867510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#867520000000
0!
0%
b0 *
0-
02
b0 6
#867530000000
1!
1%
1-
12
#867540000000
0!
0%
b1 *
0-
02
b1 6
#867550000000
1!
1%
1-
12
#867560000000
0!
0%
b10 *
0-
02
b10 6
#867570000000
1!
1%
1-
12
#867580000000
0!
0%
b11 *
0-
02
b11 6
#867590000000
1!
1%
1-
12
15
#867600000000
0!
0%
b100 *
0-
02
b100 6
#867610000000
1!
1%
1-
12
#867620000000
0!
0%
b101 *
0-
02
b101 6
#867630000000
1!
1%
1-
12
#867640000000
0!
0%
b110 *
0-
02
b110 6
#867650000000
1!
1%
1-
12
#867660000000
0!
0%
b111 *
0-
02
b111 6
#867670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#867680000000
0!
0%
b0 *
0-
02
b0 6
#867690000000
1!
1%
1-
12
#867700000000
0!
0%
b1 *
0-
02
b1 6
#867710000000
1!
1%
1-
12
#867720000000
0!
0%
b10 *
0-
02
b10 6
#867730000000
1!
1%
1-
12
#867740000000
0!
0%
b11 *
0-
02
b11 6
#867750000000
1!
1%
1-
12
15
#867760000000
0!
0%
b100 *
0-
02
b100 6
#867770000000
1!
1%
1-
12
#867780000000
0!
0%
b101 *
0-
02
b101 6
#867790000000
1!
1%
1-
12
#867800000000
0!
0%
b110 *
0-
02
b110 6
#867810000000
1!
1%
1-
12
#867820000000
0!
0%
b111 *
0-
02
b111 6
#867830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#867840000000
0!
0%
b0 *
0-
02
b0 6
#867850000000
1!
1%
1-
12
#867860000000
0!
0%
b1 *
0-
02
b1 6
#867870000000
1!
1%
1-
12
#867880000000
0!
0%
b10 *
0-
02
b10 6
#867890000000
1!
1%
1-
12
#867900000000
0!
0%
b11 *
0-
02
b11 6
#867910000000
1!
1%
1-
12
15
#867920000000
0!
0%
b100 *
0-
02
b100 6
#867930000000
1!
1%
1-
12
#867940000000
0!
0%
b101 *
0-
02
b101 6
#867950000000
1!
1%
1-
12
#867960000000
0!
0%
b110 *
0-
02
b110 6
#867970000000
1!
1%
1-
12
#867980000000
0!
0%
b111 *
0-
02
b111 6
#867990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#868000000000
0!
0%
b0 *
0-
02
b0 6
#868010000000
1!
1%
1-
12
#868020000000
0!
0%
b1 *
0-
02
b1 6
#868030000000
1!
1%
1-
12
#868040000000
0!
0%
b10 *
0-
02
b10 6
#868050000000
1!
1%
1-
12
#868060000000
0!
0%
b11 *
0-
02
b11 6
#868070000000
1!
1%
1-
12
15
#868080000000
0!
0%
b100 *
0-
02
b100 6
#868090000000
1!
1%
1-
12
#868100000000
0!
0%
b101 *
0-
02
b101 6
#868110000000
1!
1%
1-
12
#868120000000
0!
0%
b110 *
0-
02
b110 6
#868130000000
1!
1%
1-
12
#868140000000
0!
0%
b111 *
0-
02
b111 6
#868150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#868160000000
0!
0%
b0 *
0-
02
b0 6
#868170000000
1!
1%
1-
12
#868180000000
0!
0%
b1 *
0-
02
b1 6
#868190000000
1!
1%
1-
12
#868200000000
0!
0%
b10 *
0-
02
b10 6
#868210000000
1!
1%
1-
12
#868220000000
0!
0%
b11 *
0-
02
b11 6
#868230000000
1!
1%
1-
12
15
#868240000000
0!
0%
b100 *
0-
02
b100 6
#868250000000
1!
1%
1-
12
#868260000000
0!
0%
b101 *
0-
02
b101 6
#868270000000
1!
1%
1-
12
#868280000000
0!
0%
b110 *
0-
02
b110 6
#868290000000
1!
1%
1-
12
#868300000000
0!
0%
b111 *
0-
02
b111 6
#868310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#868320000000
0!
0%
b0 *
0-
02
b0 6
#868330000000
1!
1%
1-
12
#868340000000
0!
0%
b1 *
0-
02
b1 6
#868350000000
1!
1%
1-
12
#868360000000
0!
0%
b10 *
0-
02
b10 6
#868370000000
1!
1%
1-
12
#868380000000
0!
0%
b11 *
0-
02
b11 6
#868390000000
1!
1%
1-
12
15
#868400000000
0!
0%
b100 *
0-
02
b100 6
#868410000000
1!
1%
1-
12
#868420000000
0!
0%
b101 *
0-
02
b101 6
#868430000000
1!
1%
1-
12
#868440000000
0!
0%
b110 *
0-
02
b110 6
#868450000000
1!
1%
1-
12
#868460000000
0!
0%
b111 *
0-
02
b111 6
#868470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#868480000000
0!
0%
b0 *
0-
02
b0 6
#868490000000
1!
1%
1-
12
#868500000000
0!
0%
b1 *
0-
02
b1 6
#868510000000
1!
1%
1-
12
#868520000000
0!
0%
b10 *
0-
02
b10 6
#868530000000
1!
1%
1-
12
#868540000000
0!
0%
b11 *
0-
02
b11 6
#868550000000
1!
1%
1-
12
15
#868560000000
0!
0%
b100 *
0-
02
b100 6
#868570000000
1!
1%
1-
12
#868580000000
0!
0%
b101 *
0-
02
b101 6
#868590000000
1!
1%
1-
12
#868600000000
0!
0%
b110 *
0-
02
b110 6
#868610000000
1!
1%
1-
12
#868620000000
0!
0%
b111 *
0-
02
b111 6
#868630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#868640000000
0!
0%
b0 *
0-
02
b0 6
#868650000000
1!
1%
1-
12
#868660000000
0!
0%
b1 *
0-
02
b1 6
#868670000000
1!
1%
1-
12
#868680000000
0!
0%
b10 *
0-
02
b10 6
#868690000000
1!
1%
1-
12
#868700000000
0!
0%
b11 *
0-
02
b11 6
#868710000000
1!
1%
1-
12
15
#868720000000
0!
0%
b100 *
0-
02
b100 6
#868730000000
1!
1%
1-
12
#868740000000
0!
0%
b101 *
0-
02
b101 6
#868750000000
1!
1%
1-
12
#868760000000
0!
0%
b110 *
0-
02
b110 6
#868770000000
1!
1%
1-
12
#868780000000
0!
0%
b111 *
0-
02
b111 6
#868790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#868800000000
0!
0%
b0 *
0-
02
b0 6
#868810000000
1!
1%
1-
12
#868820000000
0!
0%
b1 *
0-
02
b1 6
#868830000000
1!
1%
1-
12
#868840000000
0!
0%
b10 *
0-
02
b10 6
#868850000000
1!
1%
1-
12
#868860000000
0!
0%
b11 *
0-
02
b11 6
#868870000000
1!
1%
1-
12
15
#868880000000
0!
0%
b100 *
0-
02
b100 6
#868890000000
1!
1%
1-
12
#868900000000
0!
0%
b101 *
0-
02
b101 6
#868910000000
1!
1%
1-
12
#868920000000
0!
0%
b110 *
0-
02
b110 6
#868930000000
1!
1%
1-
12
#868940000000
0!
0%
b111 *
0-
02
b111 6
#868950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#868960000000
0!
0%
b0 *
0-
02
b0 6
#868970000000
1!
1%
1-
12
#868980000000
0!
0%
b1 *
0-
02
b1 6
#868990000000
1!
1%
1-
12
#869000000000
0!
0%
b10 *
0-
02
b10 6
#869010000000
1!
1%
1-
12
#869020000000
0!
0%
b11 *
0-
02
b11 6
#869030000000
1!
1%
1-
12
15
#869040000000
0!
0%
b100 *
0-
02
b100 6
#869050000000
1!
1%
1-
12
#869060000000
0!
0%
b101 *
0-
02
b101 6
#869070000000
1!
1%
1-
12
#869080000000
0!
0%
b110 *
0-
02
b110 6
#869090000000
1!
1%
1-
12
#869100000000
0!
0%
b111 *
0-
02
b111 6
#869110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#869120000000
0!
0%
b0 *
0-
02
b0 6
#869130000000
1!
1%
1-
12
#869140000000
0!
0%
b1 *
0-
02
b1 6
#869150000000
1!
1%
1-
12
#869160000000
0!
0%
b10 *
0-
02
b10 6
#869170000000
1!
1%
1-
12
#869180000000
0!
0%
b11 *
0-
02
b11 6
#869190000000
1!
1%
1-
12
15
#869200000000
0!
0%
b100 *
0-
02
b100 6
#869210000000
1!
1%
1-
12
#869220000000
0!
0%
b101 *
0-
02
b101 6
#869230000000
1!
1%
1-
12
#869240000000
0!
0%
b110 *
0-
02
b110 6
#869250000000
1!
1%
1-
12
#869260000000
0!
0%
b111 *
0-
02
b111 6
#869270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#869280000000
0!
0%
b0 *
0-
02
b0 6
#869290000000
1!
1%
1-
12
#869300000000
0!
0%
b1 *
0-
02
b1 6
#869310000000
1!
1%
1-
12
#869320000000
0!
0%
b10 *
0-
02
b10 6
#869330000000
1!
1%
1-
12
#869340000000
0!
0%
b11 *
0-
02
b11 6
#869350000000
1!
1%
1-
12
15
#869360000000
0!
0%
b100 *
0-
02
b100 6
#869370000000
1!
1%
1-
12
#869380000000
0!
0%
b101 *
0-
02
b101 6
#869390000000
1!
1%
1-
12
#869400000000
0!
0%
b110 *
0-
02
b110 6
#869410000000
1!
1%
1-
12
#869420000000
0!
0%
b111 *
0-
02
b111 6
#869430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#869440000000
0!
0%
b0 *
0-
02
b0 6
#869450000000
1!
1%
1-
12
#869460000000
0!
0%
b1 *
0-
02
b1 6
#869470000000
1!
1%
1-
12
#869480000000
0!
0%
b10 *
0-
02
b10 6
#869490000000
1!
1%
1-
12
#869500000000
0!
0%
b11 *
0-
02
b11 6
#869510000000
1!
1%
1-
12
15
#869520000000
0!
0%
b100 *
0-
02
b100 6
#869530000000
1!
1%
1-
12
#869540000000
0!
0%
b101 *
0-
02
b101 6
#869550000000
1!
1%
1-
12
#869560000000
0!
0%
b110 *
0-
02
b110 6
#869570000000
1!
1%
1-
12
#869580000000
0!
0%
b111 *
0-
02
b111 6
#869590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#869600000000
0!
0%
b0 *
0-
02
b0 6
#869610000000
1!
1%
1-
12
#869620000000
0!
0%
b1 *
0-
02
b1 6
#869630000000
1!
1%
1-
12
#869640000000
0!
0%
b10 *
0-
02
b10 6
#869650000000
1!
1%
1-
12
#869660000000
0!
0%
b11 *
0-
02
b11 6
#869670000000
1!
1%
1-
12
15
#869680000000
0!
0%
b100 *
0-
02
b100 6
#869690000000
1!
1%
1-
12
#869700000000
0!
0%
b101 *
0-
02
b101 6
#869710000000
1!
1%
1-
12
#869720000000
0!
0%
b110 *
0-
02
b110 6
#869730000000
1!
1%
1-
12
#869740000000
0!
0%
b111 *
0-
02
b111 6
#869750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#869760000000
0!
0%
b0 *
0-
02
b0 6
#869770000000
1!
1%
1-
12
#869780000000
0!
0%
b1 *
0-
02
b1 6
#869790000000
1!
1%
1-
12
#869800000000
0!
0%
b10 *
0-
02
b10 6
#869810000000
1!
1%
1-
12
#869820000000
0!
0%
b11 *
0-
02
b11 6
#869830000000
1!
1%
1-
12
15
#869840000000
0!
0%
b100 *
0-
02
b100 6
#869850000000
1!
1%
1-
12
#869860000000
0!
0%
b101 *
0-
02
b101 6
#869870000000
1!
1%
1-
12
#869880000000
0!
0%
b110 *
0-
02
b110 6
#869890000000
1!
1%
1-
12
#869900000000
0!
0%
b111 *
0-
02
b111 6
#869910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#869920000000
0!
0%
b0 *
0-
02
b0 6
#869930000000
1!
1%
1-
12
#869940000000
0!
0%
b1 *
0-
02
b1 6
#869950000000
1!
1%
1-
12
#869960000000
0!
0%
b10 *
0-
02
b10 6
#869970000000
1!
1%
1-
12
#869980000000
0!
0%
b11 *
0-
02
b11 6
#869990000000
1!
1%
1-
12
15
#870000000000
0!
0%
b100 *
0-
02
b100 6
#870010000000
1!
1%
1-
12
#870020000000
0!
0%
b101 *
0-
02
b101 6
#870030000000
1!
1%
1-
12
#870040000000
0!
0%
b110 *
0-
02
b110 6
#870050000000
1!
1%
1-
12
#870060000000
0!
0%
b111 *
0-
02
b111 6
#870070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#870080000000
0!
0%
b0 *
0-
02
b0 6
#870090000000
1!
1%
1-
12
#870100000000
0!
0%
b1 *
0-
02
b1 6
#870110000000
1!
1%
1-
12
#870120000000
0!
0%
b10 *
0-
02
b10 6
#870130000000
1!
1%
1-
12
#870140000000
0!
0%
b11 *
0-
02
b11 6
#870150000000
1!
1%
1-
12
15
#870160000000
0!
0%
b100 *
0-
02
b100 6
#870170000000
1!
1%
1-
12
#870180000000
0!
0%
b101 *
0-
02
b101 6
#870190000000
1!
1%
1-
12
#870200000000
0!
0%
b110 *
0-
02
b110 6
#870210000000
1!
1%
1-
12
#870220000000
0!
0%
b111 *
0-
02
b111 6
#870230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#870240000000
0!
0%
b0 *
0-
02
b0 6
#870250000000
1!
1%
1-
12
#870260000000
0!
0%
b1 *
0-
02
b1 6
#870270000000
1!
1%
1-
12
#870280000000
0!
0%
b10 *
0-
02
b10 6
#870290000000
1!
1%
1-
12
#870300000000
0!
0%
b11 *
0-
02
b11 6
#870310000000
1!
1%
1-
12
15
#870320000000
0!
0%
b100 *
0-
02
b100 6
#870330000000
1!
1%
1-
12
#870340000000
0!
0%
b101 *
0-
02
b101 6
#870350000000
1!
1%
1-
12
#870360000000
0!
0%
b110 *
0-
02
b110 6
#870370000000
1!
1%
1-
12
#870380000000
0!
0%
b111 *
0-
02
b111 6
#870390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#870400000000
0!
0%
b0 *
0-
02
b0 6
#870410000000
1!
1%
1-
12
#870420000000
0!
0%
b1 *
0-
02
b1 6
#870430000000
1!
1%
1-
12
#870440000000
0!
0%
b10 *
0-
02
b10 6
#870450000000
1!
1%
1-
12
#870460000000
0!
0%
b11 *
0-
02
b11 6
#870470000000
1!
1%
1-
12
15
#870480000000
0!
0%
b100 *
0-
02
b100 6
#870490000000
1!
1%
1-
12
#870500000000
0!
0%
b101 *
0-
02
b101 6
#870510000000
1!
1%
1-
12
#870520000000
0!
0%
b110 *
0-
02
b110 6
#870530000000
1!
1%
1-
12
#870540000000
0!
0%
b111 *
0-
02
b111 6
#870550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#870560000000
0!
0%
b0 *
0-
02
b0 6
#870570000000
1!
1%
1-
12
#870580000000
0!
0%
b1 *
0-
02
b1 6
#870590000000
1!
1%
1-
12
#870600000000
0!
0%
b10 *
0-
02
b10 6
#870610000000
1!
1%
1-
12
#870620000000
0!
0%
b11 *
0-
02
b11 6
#870630000000
1!
1%
1-
12
15
#870640000000
0!
0%
b100 *
0-
02
b100 6
#870650000000
1!
1%
1-
12
#870660000000
0!
0%
b101 *
0-
02
b101 6
#870670000000
1!
1%
1-
12
#870680000000
0!
0%
b110 *
0-
02
b110 6
#870690000000
1!
1%
1-
12
#870700000000
0!
0%
b111 *
0-
02
b111 6
#870710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#870720000000
0!
0%
b0 *
0-
02
b0 6
#870730000000
1!
1%
1-
12
#870740000000
0!
0%
b1 *
0-
02
b1 6
#870750000000
1!
1%
1-
12
#870760000000
0!
0%
b10 *
0-
02
b10 6
#870770000000
1!
1%
1-
12
#870780000000
0!
0%
b11 *
0-
02
b11 6
#870790000000
1!
1%
1-
12
15
#870800000000
0!
0%
b100 *
0-
02
b100 6
#870810000000
1!
1%
1-
12
#870820000000
0!
0%
b101 *
0-
02
b101 6
#870830000000
1!
1%
1-
12
#870840000000
0!
0%
b110 *
0-
02
b110 6
#870850000000
1!
1%
1-
12
#870860000000
0!
0%
b111 *
0-
02
b111 6
#870870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#870880000000
0!
0%
b0 *
0-
02
b0 6
#870890000000
1!
1%
1-
12
#870900000000
0!
0%
b1 *
0-
02
b1 6
#870910000000
1!
1%
1-
12
#870920000000
0!
0%
b10 *
0-
02
b10 6
#870930000000
1!
1%
1-
12
#870940000000
0!
0%
b11 *
0-
02
b11 6
#870950000000
1!
1%
1-
12
15
#870960000000
0!
0%
b100 *
0-
02
b100 6
#870970000000
1!
1%
1-
12
#870980000000
0!
0%
b101 *
0-
02
b101 6
#870990000000
1!
1%
1-
12
#871000000000
0!
0%
b110 *
0-
02
b110 6
#871010000000
1!
1%
1-
12
#871020000000
0!
0%
b111 *
0-
02
b111 6
#871030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#871040000000
0!
0%
b0 *
0-
02
b0 6
#871050000000
1!
1%
1-
12
#871060000000
0!
0%
b1 *
0-
02
b1 6
#871070000000
1!
1%
1-
12
#871080000000
0!
0%
b10 *
0-
02
b10 6
#871090000000
1!
1%
1-
12
#871100000000
0!
0%
b11 *
0-
02
b11 6
#871110000000
1!
1%
1-
12
15
#871120000000
0!
0%
b100 *
0-
02
b100 6
#871130000000
1!
1%
1-
12
#871140000000
0!
0%
b101 *
0-
02
b101 6
#871150000000
1!
1%
1-
12
#871160000000
0!
0%
b110 *
0-
02
b110 6
#871170000000
1!
1%
1-
12
#871180000000
0!
0%
b111 *
0-
02
b111 6
#871190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#871200000000
0!
0%
b0 *
0-
02
b0 6
#871210000000
1!
1%
1-
12
#871220000000
0!
0%
b1 *
0-
02
b1 6
#871230000000
1!
1%
1-
12
#871240000000
0!
0%
b10 *
0-
02
b10 6
#871250000000
1!
1%
1-
12
#871260000000
0!
0%
b11 *
0-
02
b11 6
#871270000000
1!
1%
1-
12
15
#871280000000
0!
0%
b100 *
0-
02
b100 6
#871290000000
1!
1%
1-
12
#871300000000
0!
0%
b101 *
0-
02
b101 6
#871310000000
1!
1%
1-
12
#871320000000
0!
0%
b110 *
0-
02
b110 6
#871330000000
1!
1%
1-
12
#871340000000
0!
0%
b111 *
0-
02
b111 6
#871350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#871360000000
0!
0%
b0 *
0-
02
b0 6
#871370000000
1!
1%
1-
12
#871380000000
0!
0%
b1 *
0-
02
b1 6
#871390000000
1!
1%
1-
12
#871400000000
0!
0%
b10 *
0-
02
b10 6
#871410000000
1!
1%
1-
12
#871420000000
0!
0%
b11 *
0-
02
b11 6
#871430000000
1!
1%
1-
12
15
#871440000000
0!
0%
b100 *
0-
02
b100 6
#871450000000
1!
1%
1-
12
#871460000000
0!
0%
b101 *
0-
02
b101 6
#871470000000
1!
1%
1-
12
#871480000000
0!
0%
b110 *
0-
02
b110 6
#871490000000
1!
1%
1-
12
#871500000000
0!
0%
b111 *
0-
02
b111 6
#871510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#871520000000
0!
0%
b0 *
0-
02
b0 6
#871530000000
1!
1%
1-
12
#871540000000
0!
0%
b1 *
0-
02
b1 6
#871550000000
1!
1%
1-
12
#871560000000
0!
0%
b10 *
0-
02
b10 6
#871570000000
1!
1%
1-
12
#871580000000
0!
0%
b11 *
0-
02
b11 6
#871590000000
1!
1%
1-
12
15
#871600000000
0!
0%
b100 *
0-
02
b100 6
#871610000000
1!
1%
1-
12
#871620000000
0!
0%
b101 *
0-
02
b101 6
#871630000000
1!
1%
1-
12
#871640000000
0!
0%
b110 *
0-
02
b110 6
#871650000000
1!
1%
1-
12
#871660000000
0!
0%
b111 *
0-
02
b111 6
#871670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#871680000000
0!
0%
b0 *
0-
02
b0 6
#871690000000
1!
1%
1-
12
#871700000000
0!
0%
b1 *
0-
02
b1 6
#871710000000
1!
1%
1-
12
#871720000000
0!
0%
b10 *
0-
02
b10 6
#871730000000
1!
1%
1-
12
#871740000000
0!
0%
b11 *
0-
02
b11 6
#871750000000
1!
1%
1-
12
15
#871760000000
0!
0%
b100 *
0-
02
b100 6
#871770000000
1!
1%
1-
12
#871780000000
0!
0%
b101 *
0-
02
b101 6
#871790000000
1!
1%
1-
12
#871800000000
0!
0%
b110 *
0-
02
b110 6
#871810000000
1!
1%
1-
12
#871820000000
0!
0%
b111 *
0-
02
b111 6
#871830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#871840000000
0!
0%
b0 *
0-
02
b0 6
#871850000000
1!
1%
1-
12
#871860000000
0!
0%
b1 *
0-
02
b1 6
#871870000000
1!
1%
1-
12
#871880000000
0!
0%
b10 *
0-
02
b10 6
#871890000000
1!
1%
1-
12
#871900000000
0!
0%
b11 *
0-
02
b11 6
#871910000000
1!
1%
1-
12
15
#871920000000
0!
0%
b100 *
0-
02
b100 6
#871930000000
1!
1%
1-
12
#871940000000
0!
0%
b101 *
0-
02
b101 6
#871950000000
1!
1%
1-
12
#871960000000
0!
0%
b110 *
0-
02
b110 6
#871970000000
1!
1%
1-
12
#871980000000
0!
0%
b111 *
0-
02
b111 6
#871990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#872000000000
0!
0%
b0 *
0-
02
b0 6
#872010000000
1!
1%
1-
12
#872020000000
0!
0%
b1 *
0-
02
b1 6
#872030000000
1!
1%
1-
12
#872040000000
0!
0%
b10 *
0-
02
b10 6
#872050000000
1!
1%
1-
12
#872060000000
0!
0%
b11 *
0-
02
b11 6
#872070000000
1!
1%
1-
12
15
#872080000000
0!
0%
b100 *
0-
02
b100 6
#872090000000
1!
1%
1-
12
#872100000000
0!
0%
b101 *
0-
02
b101 6
#872110000000
1!
1%
1-
12
#872120000000
0!
0%
b110 *
0-
02
b110 6
#872130000000
1!
1%
1-
12
#872140000000
0!
0%
b111 *
0-
02
b111 6
#872150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#872160000000
0!
0%
b0 *
0-
02
b0 6
#872170000000
1!
1%
1-
12
#872180000000
0!
0%
b1 *
0-
02
b1 6
#872190000000
1!
1%
1-
12
#872200000000
0!
0%
b10 *
0-
02
b10 6
#872210000000
1!
1%
1-
12
#872220000000
0!
0%
b11 *
0-
02
b11 6
#872230000000
1!
1%
1-
12
15
#872240000000
0!
0%
b100 *
0-
02
b100 6
#872250000000
1!
1%
1-
12
#872260000000
0!
0%
b101 *
0-
02
b101 6
#872270000000
1!
1%
1-
12
#872280000000
0!
0%
b110 *
0-
02
b110 6
#872290000000
1!
1%
1-
12
#872300000000
0!
0%
b111 *
0-
02
b111 6
#872310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#872320000000
0!
0%
b0 *
0-
02
b0 6
#872330000000
1!
1%
1-
12
#872340000000
0!
0%
b1 *
0-
02
b1 6
#872350000000
1!
1%
1-
12
#872360000000
0!
0%
b10 *
0-
02
b10 6
#872370000000
1!
1%
1-
12
#872380000000
0!
0%
b11 *
0-
02
b11 6
#872390000000
1!
1%
1-
12
15
#872400000000
0!
0%
b100 *
0-
02
b100 6
#872410000000
1!
1%
1-
12
#872420000000
0!
0%
b101 *
0-
02
b101 6
#872430000000
1!
1%
1-
12
#872440000000
0!
0%
b110 *
0-
02
b110 6
#872450000000
1!
1%
1-
12
#872460000000
0!
0%
b111 *
0-
02
b111 6
#872470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#872480000000
0!
0%
b0 *
0-
02
b0 6
#872490000000
1!
1%
1-
12
#872500000000
0!
0%
b1 *
0-
02
b1 6
#872510000000
1!
1%
1-
12
#872520000000
0!
0%
b10 *
0-
02
b10 6
#872530000000
1!
1%
1-
12
#872540000000
0!
0%
b11 *
0-
02
b11 6
#872550000000
1!
1%
1-
12
15
#872560000000
0!
0%
b100 *
0-
02
b100 6
#872570000000
1!
1%
1-
12
#872580000000
0!
0%
b101 *
0-
02
b101 6
#872590000000
1!
1%
1-
12
#872600000000
0!
0%
b110 *
0-
02
b110 6
#872610000000
1!
1%
1-
12
#872620000000
0!
0%
b111 *
0-
02
b111 6
#872630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#872640000000
0!
0%
b0 *
0-
02
b0 6
#872650000000
1!
1%
1-
12
#872660000000
0!
0%
b1 *
0-
02
b1 6
#872670000000
1!
1%
1-
12
#872680000000
0!
0%
b10 *
0-
02
b10 6
#872690000000
1!
1%
1-
12
#872700000000
0!
0%
b11 *
0-
02
b11 6
#872710000000
1!
1%
1-
12
15
#872720000000
0!
0%
b100 *
0-
02
b100 6
#872730000000
1!
1%
1-
12
#872740000000
0!
0%
b101 *
0-
02
b101 6
#872750000000
1!
1%
1-
12
#872760000000
0!
0%
b110 *
0-
02
b110 6
#872770000000
1!
1%
1-
12
#872780000000
0!
0%
b111 *
0-
02
b111 6
#872790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#872800000000
0!
0%
b0 *
0-
02
b0 6
#872810000000
1!
1%
1-
12
#872820000000
0!
0%
b1 *
0-
02
b1 6
#872830000000
1!
1%
1-
12
#872840000000
0!
0%
b10 *
0-
02
b10 6
#872850000000
1!
1%
1-
12
#872860000000
0!
0%
b11 *
0-
02
b11 6
#872870000000
1!
1%
1-
12
15
#872880000000
0!
0%
b100 *
0-
02
b100 6
#872890000000
1!
1%
1-
12
#872900000000
0!
0%
b101 *
0-
02
b101 6
#872910000000
1!
1%
1-
12
#872920000000
0!
0%
b110 *
0-
02
b110 6
#872930000000
1!
1%
1-
12
#872940000000
0!
0%
b111 *
0-
02
b111 6
#872950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#872960000000
0!
0%
b0 *
0-
02
b0 6
#872970000000
1!
1%
1-
12
#872980000000
0!
0%
b1 *
0-
02
b1 6
#872990000000
1!
1%
1-
12
#873000000000
0!
0%
b10 *
0-
02
b10 6
#873010000000
1!
1%
1-
12
#873020000000
0!
0%
b11 *
0-
02
b11 6
#873030000000
1!
1%
1-
12
15
#873040000000
0!
0%
b100 *
0-
02
b100 6
#873050000000
1!
1%
1-
12
#873060000000
0!
0%
b101 *
0-
02
b101 6
#873070000000
1!
1%
1-
12
#873080000000
0!
0%
b110 *
0-
02
b110 6
#873090000000
1!
1%
1-
12
#873100000000
0!
0%
b111 *
0-
02
b111 6
#873110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#873120000000
0!
0%
b0 *
0-
02
b0 6
#873130000000
1!
1%
1-
12
#873140000000
0!
0%
b1 *
0-
02
b1 6
#873150000000
1!
1%
1-
12
#873160000000
0!
0%
b10 *
0-
02
b10 6
#873170000000
1!
1%
1-
12
#873180000000
0!
0%
b11 *
0-
02
b11 6
#873190000000
1!
1%
1-
12
15
#873200000000
0!
0%
b100 *
0-
02
b100 6
#873210000000
1!
1%
1-
12
#873220000000
0!
0%
b101 *
0-
02
b101 6
#873230000000
1!
1%
1-
12
#873240000000
0!
0%
b110 *
0-
02
b110 6
#873250000000
1!
1%
1-
12
#873260000000
0!
0%
b111 *
0-
02
b111 6
#873270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#873280000000
0!
0%
b0 *
0-
02
b0 6
#873290000000
1!
1%
1-
12
#873300000000
0!
0%
b1 *
0-
02
b1 6
#873310000000
1!
1%
1-
12
#873320000000
0!
0%
b10 *
0-
02
b10 6
#873330000000
1!
1%
1-
12
#873340000000
0!
0%
b11 *
0-
02
b11 6
#873350000000
1!
1%
1-
12
15
#873360000000
0!
0%
b100 *
0-
02
b100 6
#873370000000
1!
1%
1-
12
#873380000000
0!
0%
b101 *
0-
02
b101 6
#873390000000
1!
1%
1-
12
#873400000000
0!
0%
b110 *
0-
02
b110 6
#873410000000
1!
1%
1-
12
#873420000000
0!
0%
b111 *
0-
02
b111 6
#873430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#873440000000
0!
0%
b0 *
0-
02
b0 6
#873450000000
1!
1%
1-
12
#873460000000
0!
0%
b1 *
0-
02
b1 6
#873470000000
1!
1%
1-
12
#873480000000
0!
0%
b10 *
0-
02
b10 6
#873490000000
1!
1%
1-
12
#873500000000
0!
0%
b11 *
0-
02
b11 6
#873510000000
1!
1%
1-
12
15
#873520000000
0!
0%
b100 *
0-
02
b100 6
#873530000000
1!
1%
1-
12
#873540000000
0!
0%
b101 *
0-
02
b101 6
#873550000000
1!
1%
1-
12
#873560000000
0!
0%
b110 *
0-
02
b110 6
#873570000000
1!
1%
1-
12
#873580000000
0!
0%
b111 *
0-
02
b111 6
#873590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#873600000000
0!
0%
b0 *
0-
02
b0 6
#873610000000
1!
1%
1-
12
#873620000000
0!
0%
b1 *
0-
02
b1 6
#873630000000
1!
1%
1-
12
#873640000000
0!
0%
b10 *
0-
02
b10 6
#873650000000
1!
1%
1-
12
#873660000000
0!
0%
b11 *
0-
02
b11 6
#873670000000
1!
1%
1-
12
15
#873680000000
0!
0%
b100 *
0-
02
b100 6
#873690000000
1!
1%
1-
12
#873700000000
0!
0%
b101 *
0-
02
b101 6
#873710000000
1!
1%
1-
12
#873720000000
0!
0%
b110 *
0-
02
b110 6
#873730000000
1!
1%
1-
12
#873740000000
0!
0%
b111 *
0-
02
b111 6
#873750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#873760000000
0!
0%
b0 *
0-
02
b0 6
#873770000000
1!
1%
1-
12
#873780000000
0!
0%
b1 *
0-
02
b1 6
#873790000000
1!
1%
1-
12
#873800000000
0!
0%
b10 *
0-
02
b10 6
#873810000000
1!
1%
1-
12
#873820000000
0!
0%
b11 *
0-
02
b11 6
#873830000000
1!
1%
1-
12
15
#873840000000
0!
0%
b100 *
0-
02
b100 6
#873850000000
1!
1%
1-
12
#873860000000
0!
0%
b101 *
0-
02
b101 6
#873870000000
1!
1%
1-
12
#873880000000
0!
0%
b110 *
0-
02
b110 6
#873890000000
1!
1%
1-
12
#873900000000
0!
0%
b111 *
0-
02
b111 6
#873910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#873920000000
0!
0%
b0 *
0-
02
b0 6
#873930000000
1!
1%
1-
12
#873940000000
0!
0%
b1 *
0-
02
b1 6
#873950000000
1!
1%
1-
12
#873960000000
0!
0%
b10 *
0-
02
b10 6
#873970000000
1!
1%
1-
12
#873980000000
0!
0%
b11 *
0-
02
b11 6
#873990000000
1!
1%
1-
12
15
#874000000000
0!
0%
b100 *
0-
02
b100 6
#874010000000
1!
1%
1-
12
#874020000000
0!
0%
b101 *
0-
02
b101 6
#874030000000
1!
1%
1-
12
#874040000000
0!
0%
b110 *
0-
02
b110 6
#874050000000
1!
1%
1-
12
#874060000000
0!
0%
b111 *
0-
02
b111 6
#874070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#874080000000
0!
0%
b0 *
0-
02
b0 6
#874090000000
1!
1%
1-
12
#874100000000
0!
0%
b1 *
0-
02
b1 6
#874110000000
1!
1%
1-
12
#874120000000
0!
0%
b10 *
0-
02
b10 6
#874130000000
1!
1%
1-
12
#874140000000
0!
0%
b11 *
0-
02
b11 6
#874150000000
1!
1%
1-
12
15
#874160000000
0!
0%
b100 *
0-
02
b100 6
#874170000000
1!
1%
1-
12
#874180000000
0!
0%
b101 *
0-
02
b101 6
#874190000000
1!
1%
1-
12
#874200000000
0!
0%
b110 *
0-
02
b110 6
#874210000000
1!
1%
1-
12
#874220000000
0!
0%
b111 *
0-
02
b111 6
#874230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#874240000000
0!
0%
b0 *
0-
02
b0 6
#874250000000
1!
1%
1-
12
#874260000000
0!
0%
b1 *
0-
02
b1 6
#874270000000
1!
1%
1-
12
#874280000000
0!
0%
b10 *
0-
02
b10 6
#874290000000
1!
1%
1-
12
#874300000000
0!
0%
b11 *
0-
02
b11 6
#874310000000
1!
1%
1-
12
15
#874320000000
0!
0%
b100 *
0-
02
b100 6
#874330000000
1!
1%
1-
12
#874340000000
0!
0%
b101 *
0-
02
b101 6
#874350000000
1!
1%
1-
12
#874360000000
0!
0%
b110 *
0-
02
b110 6
#874370000000
1!
1%
1-
12
#874380000000
0!
0%
b111 *
0-
02
b111 6
#874390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#874400000000
0!
0%
b0 *
0-
02
b0 6
#874410000000
1!
1%
1-
12
#874420000000
0!
0%
b1 *
0-
02
b1 6
#874430000000
1!
1%
1-
12
#874440000000
0!
0%
b10 *
0-
02
b10 6
#874450000000
1!
1%
1-
12
#874460000000
0!
0%
b11 *
0-
02
b11 6
#874470000000
1!
1%
1-
12
15
#874480000000
0!
0%
b100 *
0-
02
b100 6
#874490000000
1!
1%
1-
12
#874500000000
0!
0%
b101 *
0-
02
b101 6
#874510000000
1!
1%
1-
12
#874520000000
0!
0%
b110 *
0-
02
b110 6
#874530000000
1!
1%
1-
12
#874540000000
0!
0%
b111 *
0-
02
b111 6
#874550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#874560000000
0!
0%
b0 *
0-
02
b0 6
#874570000000
1!
1%
1-
12
#874580000000
0!
0%
b1 *
0-
02
b1 6
#874590000000
1!
1%
1-
12
#874600000000
0!
0%
b10 *
0-
02
b10 6
#874610000000
1!
1%
1-
12
#874620000000
0!
0%
b11 *
0-
02
b11 6
#874630000000
1!
1%
1-
12
15
#874640000000
0!
0%
b100 *
0-
02
b100 6
#874650000000
1!
1%
1-
12
#874660000000
0!
0%
b101 *
0-
02
b101 6
#874670000000
1!
1%
1-
12
#874680000000
0!
0%
b110 *
0-
02
b110 6
#874690000000
1!
1%
1-
12
#874700000000
0!
0%
b111 *
0-
02
b111 6
#874710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#874720000000
0!
0%
b0 *
0-
02
b0 6
#874730000000
1!
1%
1-
12
#874740000000
0!
0%
b1 *
0-
02
b1 6
#874750000000
1!
1%
1-
12
#874760000000
0!
0%
b10 *
0-
02
b10 6
#874770000000
1!
1%
1-
12
#874780000000
0!
0%
b11 *
0-
02
b11 6
#874790000000
1!
1%
1-
12
15
#874800000000
0!
0%
b100 *
0-
02
b100 6
#874810000000
1!
1%
1-
12
#874820000000
0!
0%
b101 *
0-
02
b101 6
#874830000000
1!
1%
1-
12
#874840000000
0!
0%
b110 *
0-
02
b110 6
#874850000000
1!
1%
1-
12
#874860000000
0!
0%
b111 *
0-
02
b111 6
#874870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#874880000000
0!
0%
b0 *
0-
02
b0 6
#874890000000
1!
1%
1-
12
#874900000000
0!
0%
b1 *
0-
02
b1 6
#874910000000
1!
1%
1-
12
#874920000000
0!
0%
b10 *
0-
02
b10 6
#874930000000
1!
1%
1-
12
#874940000000
0!
0%
b11 *
0-
02
b11 6
#874950000000
1!
1%
1-
12
15
#874960000000
0!
0%
b100 *
0-
02
b100 6
#874970000000
1!
1%
1-
12
#874980000000
0!
0%
b101 *
0-
02
b101 6
#874990000000
1!
1%
1-
12
#875000000000
0!
0%
b110 *
0-
02
b110 6
#875010000000
1!
1%
1-
12
#875020000000
0!
0%
b111 *
0-
02
b111 6
#875030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#875040000000
0!
0%
b0 *
0-
02
b0 6
#875050000000
1!
1%
1-
12
#875060000000
0!
0%
b1 *
0-
02
b1 6
#875070000000
1!
1%
1-
12
#875080000000
0!
0%
b10 *
0-
02
b10 6
#875090000000
1!
1%
1-
12
#875100000000
0!
0%
b11 *
0-
02
b11 6
#875110000000
1!
1%
1-
12
15
#875120000000
0!
0%
b100 *
0-
02
b100 6
#875130000000
1!
1%
1-
12
#875140000000
0!
0%
b101 *
0-
02
b101 6
#875150000000
1!
1%
1-
12
#875160000000
0!
0%
b110 *
0-
02
b110 6
#875170000000
1!
1%
1-
12
#875180000000
0!
0%
b111 *
0-
02
b111 6
#875190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#875200000000
0!
0%
b0 *
0-
02
b0 6
#875210000000
1!
1%
1-
12
#875220000000
0!
0%
b1 *
0-
02
b1 6
#875230000000
1!
1%
1-
12
#875240000000
0!
0%
b10 *
0-
02
b10 6
#875250000000
1!
1%
1-
12
#875260000000
0!
0%
b11 *
0-
02
b11 6
#875270000000
1!
1%
1-
12
15
#875280000000
0!
0%
b100 *
0-
02
b100 6
#875290000000
1!
1%
1-
12
#875300000000
0!
0%
b101 *
0-
02
b101 6
#875310000000
1!
1%
1-
12
#875320000000
0!
0%
b110 *
0-
02
b110 6
#875330000000
1!
1%
1-
12
#875340000000
0!
0%
b111 *
0-
02
b111 6
#875350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#875360000000
0!
0%
b0 *
0-
02
b0 6
#875370000000
1!
1%
1-
12
#875380000000
0!
0%
b1 *
0-
02
b1 6
#875390000000
1!
1%
1-
12
#875400000000
0!
0%
b10 *
0-
02
b10 6
#875410000000
1!
1%
1-
12
#875420000000
0!
0%
b11 *
0-
02
b11 6
#875430000000
1!
1%
1-
12
15
#875440000000
0!
0%
b100 *
0-
02
b100 6
#875450000000
1!
1%
1-
12
#875460000000
0!
0%
b101 *
0-
02
b101 6
#875470000000
1!
1%
1-
12
#875480000000
0!
0%
b110 *
0-
02
b110 6
#875490000000
1!
1%
1-
12
#875500000000
0!
0%
b111 *
0-
02
b111 6
#875510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#875520000000
0!
0%
b0 *
0-
02
b0 6
#875530000000
1!
1%
1-
12
#875540000000
0!
0%
b1 *
0-
02
b1 6
#875550000000
1!
1%
1-
12
#875560000000
0!
0%
b10 *
0-
02
b10 6
#875570000000
1!
1%
1-
12
#875580000000
0!
0%
b11 *
0-
02
b11 6
#875590000000
1!
1%
1-
12
15
#875600000000
0!
0%
b100 *
0-
02
b100 6
#875610000000
1!
1%
1-
12
#875620000000
0!
0%
b101 *
0-
02
b101 6
#875630000000
1!
1%
1-
12
#875640000000
0!
0%
b110 *
0-
02
b110 6
#875650000000
1!
1%
1-
12
#875660000000
0!
0%
b111 *
0-
02
b111 6
#875670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#875680000000
0!
0%
b0 *
0-
02
b0 6
#875690000000
1!
1%
1-
12
#875700000000
0!
0%
b1 *
0-
02
b1 6
#875710000000
1!
1%
1-
12
#875720000000
0!
0%
b10 *
0-
02
b10 6
#875730000000
1!
1%
1-
12
#875740000000
0!
0%
b11 *
0-
02
b11 6
#875750000000
1!
1%
1-
12
15
#875760000000
0!
0%
b100 *
0-
02
b100 6
#875770000000
1!
1%
1-
12
#875780000000
0!
0%
b101 *
0-
02
b101 6
#875790000000
1!
1%
1-
12
#875800000000
0!
0%
b110 *
0-
02
b110 6
#875810000000
1!
1%
1-
12
#875820000000
0!
0%
b111 *
0-
02
b111 6
#875830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#875840000000
0!
0%
b0 *
0-
02
b0 6
#875850000000
1!
1%
1-
12
#875860000000
0!
0%
b1 *
0-
02
b1 6
#875870000000
1!
1%
1-
12
#875880000000
0!
0%
b10 *
0-
02
b10 6
#875890000000
1!
1%
1-
12
#875900000000
0!
0%
b11 *
0-
02
b11 6
#875910000000
1!
1%
1-
12
15
#875920000000
0!
0%
b100 *
0-
02
b100 6
#875930000000
1!
1%
1-
12
#875940000000
0!
0%
b101 *
0-
02
b101 6
#875950000000
1!
1%
1-
12
#875960000000
0!
0%
b110 *
0-
02
b110 6
#875970000000
1!
1%
1-
12
#875980000000
0!
0%
b111 *
0-
02
b111 6
#875990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#876000000000
0!
0%
b0 *
0-
02
b0 6
#876010000000
1!
1%
1-
12
#876020000000
0!
0%
b1 *
0-
02
b1 6
#876030000000
1!
1%
1-
12
#876040000000
0!
0%
b10 *
0-
02
b10 6
#876050000000
1!
1%
1-
12
#876060000000
0!
0%
b11 *
0-
02
b11 6
#876070000000
1!
1%
1-
12
15
#876080000000
0!
0%
b100 *
0-
02
b100 6
#876090000000
1!
1%
1-
12
#876100000000
0!
0%
b101 *
0-
02
b101 6
#876110000000
1!
1%
1-
12
#876120000000
0!
0%
b110 *
0-
02
b110 6
#876130000000
1!
1%
1-
12
#876140000000
0!
0%
b111 *
0-
02
b111 6
#876150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#876160000000
0!
0%
b0 *
0-
02
b0 6
#876170000000
1!
1%
1-
12
#876180000000
0!
0%
b1 *
0-
02
b1 6
#876190000000
1!
1%
1-
12
#876200000000
0!
0%
b10 *
0-
02
b10 6
#876210000000
1!
1%
1-
12
#876220000000
0!
0%
b11 *
0-
02
b11 6
#876230000000
1!
1%
1-
12
15
#876240000000
0!
0%
b100 *
0-
02
b100 6
#876250000000
1!
1%
1-
12
#876260000000
0!
0%
b101 *
0-
02
b101 6
#876270000000
1!
1%
1-
12
#876280000000
0!
0%
b110 *
0-
02
b110 6
#876290000000
1!
1%
1-
12
#876300000000
0!
0%
b111 *
0-
02
b111 6
#876310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#876320000000
0!
0%
b0 *
0-
02
b0 6
#876330000000
1!
1%
1-
12
#876340000000
0!
0%
b1 *
0-
02
b1 6
#876350000000
1!
1%
1-
12
#876360000000
0!
0%
b10 *
0-
02
b10 6
#876370000000
1!
1%
1-
12
#876380000000
0!
0%
b11 *
0-
02
b11 6
#876390000000
1!
1%
1-
12
15
#876400000000
0!
0%
b100 *
0-
02
b100 6
#876410000000
1!
1%
1-
12
#876420000000
0!
0%
b101 *
0-
02
b101 6
#876430000000
1!
1%
1-
12
#876440000000
0!
0%
b110 *
0-
02
b110 6
#876450000000
1!
1%
1-
12
#876460000000
0!
0%
b111 *
0-
02
b111 6
#876470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#876480000000
0!
0%
b0 *
0-
02
b0 6
#876490000000
1!
1%
1-
12
#876500000000
0!
0%
b1 *
0-
02
b1 6
#876510000000
1!
1%
1-
12
#876520000000
0!
0%
b10 *
0-
02
b10 6
#876530000000
1!
1%
1-
12
#876540000000
0!
0%
b11 *
0-
02
b11 6
#876550000000
1!
1%
1-
12
15
#876560000000
0!
0%
b100 *
0-
02
b100 6
#876570000000
1!
1%
1-
12
#876580000000
0!
0%
b101 *
0-
02
b101 6
#876590000000
1!
1%
1-
12
#876600000000
0!
0%
b110 *
0-
02
b110 6
#876610000000
1!
1%
1-
12
#876620000000
0!
0%
b111 *
0-
02
b111 6
#876630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#876640000000
0!
0%
b0 *
0-
02
b0 6
#876650000000
1!
1%
1-
12
#876660000000
0!
0%
b1 *
0-
02
b1 6
#876670000000
1!
1%
1-
12
#876680000000
0!
0%
b10 *
0-
02
b10 6
#876690000000
1!
1%
1-
12
#876700000000
0!
0%
b11 *
0-
02
b11 6
#876710000000
1!
1%
1-
12
15
#876720000000
0!
0%
b100 *
0-
02
b100 6
#876730000000
1!
1%
1-
12
#876740000000
0!
0%
b101 *
0-
02
b101 6
#876750000000
1!
1%
1-
12
#876760000000
0!
0%
b110 *
0-
02
b110 6
#876770000000
1!
1%
1-
12
#876780000000
0!
0%
b111 *
0-
02
b111 6
#876790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#876800000000
0!
0%
b0 *
0-
02
b0 6
#876810000000
1!
1%
1-
12
#876820000000
0!
0%
b1 *
0-
02
b1 6
#876830000000
1!
1%
1-
12
#876840000000
0!
0%
b10 *
0-
02
b10 6
#876850000000
1!
1%
1-
12
#876860000000
0!
0%
b11 *
0-
02
b11 6
#876870000000
1!
1%
1-
12
15
#876880000000
0!
0%
b100 *
0-
02
b100 6
#876890000000
1!
1%
1-
12
#876900000000
0!
0%
b101 *
0-
02
b101 6
#876910000000
1!
1%
1-
12
#876920000000
0!
0%
b110 *
0-
02
b110 6
#876930000000
1!
1%
1-
12
#876940000000
0!
0%
b111 *
0-
02
b111 6
#876950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#876960000000
0!
0%
b0 *
0-
02
b0 6
#876970000000
1!
1%
1-
12
#876980000000
0!
0%
b1 *
0-
02
b1 6
#876990000000
1!
1%
1-
12
#877000000000
0!
0%
b10 *
0-
02
b10 6
#877010000000
1!
1%
1-
12
#877020000000
0!
0%
b11 *
0-
02
b11 6
#877030000000
1!
1%
1-
12
15
#877040000000
0!
0%
b100 *
0-
02
b100 6
#877050000000
1!
1%
1-
12
#877060000000
0!
0%
b101 *
0-
02
b101 6
#877070000000
1!
1%
1-
12
#877080000000
0!
0%
b110 *
0-
02
b110 6
#877090000000
1!
1%
1-
12
#877100000000
0!
0%
b111 *
0-
02
b111 6
#877110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#877120000000
0!
0%
b0 *
0-
02
b0 6
#877130000000
1!
1%
1-
12
#877140000000
0!
0%
b1 *
0-
02
b1 6
#877150000000
1!
1%
1-
12
#877160000000
0!
0%
b10 *
0-
02
b10 6
#877170000000
1!
1%
1-
12
#877180000000
0!
0%
b11 *
0-
02
b11 6
#877190000000
1!
1%
1-
12
15
#877200000000
0!
0%
b100 *
0-
02
b100 6
#877210000000
1!
1%
1-
12
#877220000000
0!
0%
b101 *
0-
02
b101 6
#877230000000
1!
1%
1-
12
#877240000000
0!
0%
b110 *
0-
02
b110 6
#877250000000
1!
1%
1-
12
#877260000000
0!
0%
b111 *
0-
02
b111 6
#877270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#877280000000
0!
0%
b0 *
0-
02
b0 6
#877290000000
1!
1%
1-
12
#877300000000
0!
0%
b1 *
0-
02
b1 6
#877310000000
1!
1%
1-
12
#877320000000
0!
0%
b10 *
0-
02
b10 6
#877330000000
1!
1%
1-
12
#877340000000
0!
0%
b11 *
0-
02
b11 6
#877350000000
1!
1%
1-
12
15
#877360000000
0!
0%
b100 *
0-
02
b100 6
#877370000000
1!
1%
1-
12
#877380000000
0!
0%
b101 *
0-
02
b101 6
#877390000000
1!
1%
1-
12
#877400000000
0!
0%
b110 *
0-
02
b110 6
#877410000000
1!
1%
1-
12
#877420000000
0!
0%
b111 *
0-
02
b111 6
#877430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#877440000000
0!
0%
b0 *
0-
02
b0 6
#877450000000
1!
1%
1-
12
#877460000000
0!
0%
b1 *
0-
02
b1 6
#877470000000
1!
1%
1-
12
#877480000000
0!
0%
b10 *
0-
02
b10 6
#877490000000
1!
1%
1-
12
#877500000000
0!
0%
b11 *
0-
02
b11 6
#877510000000
1!
1%
1-
12
15
#877520000000
0!
0%
b100 *
0-
02
b100 6
#877530000000
1!
1%
1-
12
#877540000000
0!
0%
b101 *
0-
02
b101 6
#877550000000
1!
1%
1-
12
#877560000000
0!
0%
b110 *
0-
02
b110 6
#877570000000
1!
1%
1-
12
#877580000000
0!
0%
b111 *
0-
02
b111 6
#877590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#877600000000
0!
0%
b0 *
0-
02
b0 6
#877610000000
1!
1%
1-
12
#877620000000
0!
0%
b1 *
0-
02
b1 6
#877630000000
1!
1%
1-
12
#877640000000
0!
0%
b10 *
0-
02
b10 6
#877650000000
1!
1%
1-
12
#877660000000
0!
0%
b11 *
0-
02
b11 6
#877670000000
1!
1%
1-
12
15
#877680000000
0!
0%
b100 *
0-
02
b100 6
#877690000000
1!
1%
1-
12
#877700000000
0!
0%
b101 *
0-
02
b101 6
#877710000000
1!
1%
1-
12
#877720000000
0!
0%
b110 *
0-
02
b110 6
#877730000000
1!
1%
1-
12
#877740000000
0!
0%
b111 *
0-
02
b111 6
#877750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#877760000000
0!
0%
b0 *
0-
02
b0 6
#877770000000
1!
1%
1-
12
#877780000000
0!
0%
b1 *
0-
02
b1 6
#877790000000
1!
1%
1-
12
#877800000000
0!
0%
b10 *
0-
02
b10 6
#877810000000
1!
1%
1-
12
#877820000000
0!
0%
b11 *
0-
02
b11 6
#877830000000
1!
1%
1-
12
15
#877840000000
0!
0%
b100 *
0-
02
b100 6
#877850000000
1!
1%
1-
12
#877860000000
0!
0%
b101 *
0-
02
b101 6
#877870000000
1!
1%
1-
12
#877880000000
0!
0%
b110 *
0-
02
b110 6
#877890000000
1!
1%
1-
12
#877900000000
0!
0%
b111 *
0-
02
b111 6
#877910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#877920000000
0!
0%
b0 *
0-
02
b0 6
#877930000000
1!
1%
1-
12
#877940000000
0!
0%
b1 *
0-
02
b1 6
#877950000000
1!
1%
1-
12
#877960000000
0!
0%
b10 *
0-
02
b10 6
#877970000000
1!
1%
1-
12
#877980000000
0!
0%
b11 *
0-
02
b11 6
#877990000000
1!
1%
1-
12
15
#878000000000
0!
0%
b100 *
0-
02
b100 6
#878010000000
1!
1%
1-
12
#878020000000
0!
0%
b101 *
0-
02
b101 6
#878030000000
1!
1%
1-
12
#878040000000
0!
0%
b110 *
0-
02
b110 6
#878050000000
1!
1%
1-
12
#878060000000
0!
0%
b111 *
0-
02
b111 6
#878070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#878080000000
0!
0%
b0 *
0-
02
b0 6
#878090000000
1!
1%
1-
12
#878100000000
0!
0%
b1 *
0-
02
b1 6
#878110000000
1!
1%
1-
12
#878120000000
0!
0%
b10 *
0-
02
b10 6
#878130000000
1!
1%
1-
12
#878140000000
0!
0%
b11 *
0-
02
b11 6
#878150000000
1!
1%
1-
12
15
#878160000000
0!
0%
b100 *
0-
02
b100 6
#878170000000
1!
1%
1-
12
#878180000000
0!
0%
b101 *
0-
02
b101 6
#878190000000
1!
1%
1-
12
#878200000000
0!
0%
b110 *
0-
02
b110 6
#878210000000
1!
1%
1-
12
#878220000000
0!
0%
b111 *
0-
02
b111 6
#878230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#878240000000
0!
0%
b0 *
0-
02
b0 6
#878250000000
1!
1%
1-
12
#878260000000
0!
0%
b1 *
0-
02
b1 6
#878270000000
1!
1%
1-
12
#878280000000
0!
0%
b10 *
0-
02
b10 6
#878290000000
1!
1%
1-
12
#878300000000
0!
0%
b11 *
0-
02
b11 6
#878310000000
1!
1%
1-
12
15
#878320000000
0!
0%
b100 *
0-
02
b100 6
#878330000000
1!
1%
1-
12
#878340000000
0!
0%
b101 *
0-
02
b101 6
#878350000000
1!
1%
1-
12
#878360000000
0!
0%
b110 *
0-
02
b110 6
#878370000000
1!
1%
1-
12
#878380000000
0!
0%
b111 *
0-
02
b111 6
#878390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#878400000000
0!
0%
b0 *
0-
02
b0 6
#878410000000
1!
1%
1-
12
#878420000000
0!
0%
b1 *
0-
02
b1 6
#878430000000
1!
1%
1-
12
#878440000000
0!
0%
b10 *
0-
02
b10 6
#878450000000
1!
1%
1-
12
#878460000000
0!
0%
b11 *
0-
02
b11 6
#878470000000
1!
1%
1-
12
15
#878480000000
0!
0%
b100 *
0-
02
b100 6
#878490000000
1!
1%
1-
12
#878500000000
0!
0%
b101 *
0-
02
b101 6
#878510000000
1!
1%
1-
12
#878520000000
0!
0%
b110 *
0-
02
b110 6
#878530000000
1!
1%
1-
12
#878540000000
0!
0%
b111 *
0-
02
b111 6
#878550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#878560000000
0!
0%
b0 *
0-
02
b0 6
#878570000000
1!
1%
1-
12
#878580000000
0!
0%
b1 *
0-
02
b1 6
#878590000000
1!
1%
1-
12
#878600000000
0!
0%
b10 *
0-
02
b10 6
#878610000000
1!
1%
1-
12
#878620000000
0!
0%
b11 *
0-
02
b11 6
#878630000000
1!
1%
1-
12
15
#878640000000
0!
0%
b100 *
0-
02
b100 6
#878650000000
1!
1%
1-
12
#878660000000
0!
0%
b101 *
0-
02
b101 6
#878670000000
1!
1%
1-
12
#878680000000
0!
0%
b110 *
0-
02
b110 6
#878690000000
1!
1%
1-
12
#878700000000
0!
0%
b111 *
0-
02
b111 6
#878710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#878720000000
0!
0%
b0 *
0-
02
b0 6
#878730000000
1!
1%
1-
12
#878740000000
0!
0%
b1 *
0-
02
b1 6
#878750000000
1!
1%
1-
12
#878760000000
0!
0%
b10 *
0-
02
b10 6
#878770000000
1!
1%
1-
12
#878780000000
0!
0%
b11 *
0-
02
b11 6
#878790000000
1!
1%
1-
12
15
#878800000000
0!
0%
b100 *
0-
02
b100 6
#878810000000
1!
1%
1-
12
#878820000000
0!
0%
b101 *
0-
02
b101 6
#878830000000
1!
1%
1-
12
#878840000000
0!
0%
b110 *
0-
02
b110 6
#878850000000
1!
1%
1-
12
#878860000000
0!
0%
b111 *
0-
02
b111 6
#878870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#878880000000
0!
0%
b0 *
0-
02
b0 6
#878890000000
1!
1%
1-
12
#878900000000
0!
0%
b1 *
0-
02
b1 6
#878910000000
1!
1%
1-
12
#878920000000
0!
0%
b10 *
0-
02
b10 6
#878930000000
1!
1%
1-
12
#878940000000
0!
0%
b11 *
0-
02
b11 6
#878950000000
1!
1%
1-
12
15
#878960000000
0!
0%
b100 *
0-
02
b100 6
#878970000000
1!
1%
1-
12
#878980000000
0!
0%
b101 *
0-
02
b101 6
#878990000000
1!
1%
1-
12
#879000000000
0!
0%
b110 *
0-
02
b110 6
#879010000000
1!
1%
1-
12
#879020000000
0!
0%
b111 *
0-
02
b111 6
#879030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#879040000000
0!
0%
b0 *
0-
02
b0 6
#879050000000
1!
1%
1-
12
#879060000000
0!
0%
b1 *
0-
02
b1 6
#879070000000
1!
1%
1-
12
#879080000000
0!
0%
b10 *
0-
02
b10 6
#879090000000
1!
1%
1-
12
#879100000000
0!
0%
b11 *
0-
02
b11 6
#879110000000
1!
1%
1-
12
15
#879120000000
0!
0%
b100 *
0-
02
b100 6
#879130000000
1!
1%
1-
12
#879140000000
0!
0%
b101 *
0-
02
b101 6
#879150000000
1!
1%
1-
12
#879160000000
0!
0%
b110 *
0-
02
b110 6
#879170000000
1!
1%
1-
12
#879180000000
0!
0%
b111 *
0-
02
b111 6
#879190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#879200000000
0!
0%
b0 *
0-
02
b0 6
#879210000000
1!
1%
1-
12
#879220000000
0!
0%
b1 *
0-
02
b1 6
#879230000000
1!
1%
1-
12
#879240000000
0!
0%
b10 *
0-
02
b10 6
#879250000000
1!
1%
1-
12
#879260000000
0!
0%
b11 *
0-
02
b11 6
#879270000000
1!
1%
1-
12
15
#879280000000
0!
0%
b100 *
0-
02
b100 6
#879290000000
1!
1%
1-
12
#879300000000
0!
0%
b101 *
0-
02
b101 6
#879310000000
1!
1%
1-
12
#879320000000
0!
0%
b110 *
0-
02
b110 6
#879330000000
1!
1%
1-
12
#879340000000
0!
0%
b111 *
0-
02
b111 6
#879350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#879360000000
0!
0%
b0 *
0-
02
b0 6
#879370000000
1!
1%
1-
12
#879380000000
0!
0%
b1 *
0-
02
b1 6
#879390000000
1!
1%
1-
12
#879400000000
0!
0%
b10 *
0-
02
b10 6
#879410000000
1!
1%
1-
12
#879420000000
0!
0%
b11 *
0-
02
b11 6
#879430000000
1!
1%
1-
12
15
#879440000000
0!
0%
b100 *
0-
02
b100 6
#879450000000
1!
1%
1-
12
#879460000000
0!
0%
b101 *
0-
02
b101 6
#879470000000
1!
1%
1-
12
#879480000000
0!
0%
b110 *
0-
02
b110 6
#879490000000
1!
1%
1-
12
#879500000000
0!
0%
b111 *
0-
02
b111 6
#879510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#879520000000
0!
0%
b0 *
0-
02
b0 6
#879530000000
1!
1%
1-
12
#879540000000
0!
0%
b1 *
0-
02
b1 6
#879550000000
1!
1%
1-
12
#879560000000
0!
0%
b10 *
0-
02
b10 6
#879570000000
1!
1%
1-
12
#879580000000
0!
0%
b11 *
0-
02
b11 6
#879590000000
1!
1%
1-
12
15
#879600000000
0!
0%
b100 *
0-
02
b100 6
#879610000000
1!
1%
1-
12
#879620000000
0!
0%
b101 *
0-
02
b101 6
#879630000000
1!
1%
1-
12
#879640000000
0!
0%
b110 *
0-
02
b110 6
#879650000000
1!
1%
1-
12
#879660000000
0!
0%
b111 *
0-
02
b111 6
#879670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#879680000000
0!
0%
b0 *
0-
02
b0 6
#879690000000
1!
1%
1-
12
#879700000000
0!
0%
b1 *
0-
02
b1 6
#879710000000
1!
1%
1-
12
#879720000000
0!
0%
b10 *
0-
02
b10 6
#879730000000
1!
1%
1-
12
#879740000000
0!
0%
b11 *
0-
02
b11 6
#879750000000
1!
1%
1-
12
15
#879760000000
0!
0%
b100 *
0-
02
b100 6
#879770000000
1!
1%
1-
12
#879780000000
0!
0%
b101 *
0-
02
b101 6
#879790000000
1!
1%
1-
12
#879800000000
0!
0%
b110 *
0-
02
b110 6
#879810000000
1!
1%
1-
12
#879820000000
0!
0%
b111 *
0-
02
b111 6
#879830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#879840000000
0!
0%
b0 *
0-
02
b0 6
#879850000000
1!
1%
1-
12
#879860000000
0!
0%
b1 *
0-
02
b1 6
#879870000000
1!
1%
1-
12
#879880000000
0!
0%
b10 *
0-
02
b10 6
#879890000000
1!
1%
1-
12
#879900000000
0!
0%
b11 *
0-
02
b11 6
#879910000000
1!
1%
1-
12
15
#879920000000
0!
0%
b100 *
0-
02
b100 6
#879930000000
1!
1%
1-
12
#879940000000
0!
0%
b101 *
0-
02
b101 6
#879950000000
1!
1%
1-
12
#879960000000
0!
0%
b110 *
0-
02
b110 6
#879970000000
1!
1%
1-
12
#879980000000
0!
0%
b111 *
0-
02
b111 6
#879990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#880000000000
0!
0%
b0 *
0-
02
b0 6
#880010000000
1!
1%
1-
12
#880020000000
0!
0%
b1 *
0-
02
b1 6
#880030000000
1!
1%
1-
12
#880040000000
0!
0%
b10 *
0-
02
b10 6
#880050000000
1!
1%
1-
12
#880060000000
0!
0%
b11 *
0-
02
b11 6
#880070000000
1!
1%
1-
12
15
#880080000000
0!
0%
b100 *
0-
02
b100 6
#880090000000
1!
1%
1-
12
#880100000000
0!
0%
b101 *
0-
02
b101 6
#880110000000
1!
1%
1-
12
#880120000000
0!
0%
b110 *
0-
02
b110 6
#880130000000
1!
1%
1-
12
#880140000000
0!
0%
b111 *
0-
02
b111 6
#880150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#880160000000
0!
0%
b0 *
0-
02
b0 6
#880170000000
1!
1%
1-
12
#880180000000
0!
0%
b1 *
0-
02
b1 6
#880190000000
1!
1%
1-
12
#880200000000
0!
0%
b10 *
0-
02
b10 6
#880210000000
1!
1%
1-
12
#880220000000
0!
0%
b11 *
0-
02
b11 6
#880230000000
1!
1%
1-
12
15
#880240000000
0!
0%
b100 *
0-
02
b100 6
#880250000000
1!
1%
1-
12
#880260000000
0!
0%
b101 *
0-
02
b101 6
#880270000000
1!
1%
1-
12
#880280000000
0!
0%
b110 *
0-
02
b110 6
#880290000000
1!
1%
1-
12
#880300000000
0!
0%
b111 *
0-
02
b111 6
#880310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#880320000000
0!
0%
b0 *
0-
02
b0 6
#880330000000
1!
1%
1-
12
#880340000000
0!
0%
b1 *
0-
02
b1 6
#880350000000
1!
1%
1-
12
#880360000000
0!
0%
b10 *
0-
02
b10 6
#880370000000
1!
1%
1-
12
#880380000000
0!
0%
b11 *
0-
02
b11 6
#880390000000
1!
1%
1-
12
15
#880400000000
0!
0%
b100 *
0-
02
b100 6
#880410000000
1!
1%
1-
12
#880420000000
0!
0%
b101 *
0-
02
b101 6
#880430000000
1!
1%
1-
12
#880440000000
0!
0%
b110 *
0-
02
b110 6
#880450000000
1!
1%
1-
12
#880460000000
0!
0%
b111 *
0-
02
b111 6
#880470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#880480000000
0!
0%
b0 *
0-
02
b0 6
#880490000000
1!
1%
1-
12
#880500000000
0!
0%
b1 *
0-
02
b1 6
#880510000000
1!
1%
1-
12
#880520000000
0!
0%
b10 *
0-
02
b10 6
#880530000000
1!
1%
1-
12
#880540000000
0!
0%
b11 *
0-
02
b11 6
#880550000000
1!
1%
1-
12
15
#880560000000
0!
0%
b100 *
0-
02
b100 6
#880570000000
1!
1%
1-
12
#880580000000
0!
0%
b101 *
0-
02
b101 6
#880590000000
1!
1%
1-
12
#880600000000
0!
0%
b110 *
0-
02
b110 6
#880610000000
1!
1%
1-
12
#880620000000
0!
0%
b111 *
0-
02
b111 6
#880630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#880640000000
0!
0%
b0 *
0-
02
b0 6
#880650000000
1!
1%
1-
12
#880660000000
0!
0%
b1 *
0-
02
b1 6
#880670000000
1!
1%
1-
12
#880680000000
0!
0%
b10 *
0-
02
b10 6
#880690000000
1!
1%
1-
12
#880700000000
0!
0%
b11 *
0-
02
b11 6
#880710000000
1!
1%
1-
12
15
#880720000000
0!
0%
b100 *
0-
02
b100 6
#880730000000
1!
1%
1-
12
#880740000000
0!
0%
b101 *
0-
02
b101 6
#880750000000
1!
1%
1-
12
#880760000000
0!
0%
b110 *
0-
02
b110 6
#880770000000
1!
1%
1-
12
#880780000000
0!
0%
b111 *
0-
02
b111 6
#880790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#880800000000
0!
0%
b0 *
0-
02
b0 6
#880810000000
1!
1%
1-
12
#880820000000
0!
0%
b1 *
0-
02
b1 6
#880830000000
1!
1%
1-
12
#880840000000
0!
0%
b10 *
0-
02
b10 6
#880850000000
1!
1%
1-
12
#880860000000
0!
0%
b11 *
0-
02
b11 6
#880870000000
1!
1%
1-
12
15
#880880000000
0!
0%
b100 *
0-
02
b100 6
#880890000000
1!
1%
1-
12
#880900000000
0!
0%
b101 *
0-
02
b101 6
#880910000000
1!
1%
1-
12
#880920000000
0!
0%
b110 *
0-
02
b110 6
#880930000000
1!
1%
1-
12
#880940000000
0!
0%
b111 *
0-
02
b111 6
#880950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#880960000000
0!
0%
b0 *
0-
02
b0 6
#880970000000
1!
1%
1-
12
#880980000000
0!
0%
b1 *
0-
02
b1 6
#880990000000
1!
1%
1-
12
#881000000000
0!
0%
b10 *
0-
02
b10 6
#881010000000
1!
1%
1-
12
#881020000000
0!
0%
b11 *
0-
02
b11 6
#881030000000
1!
1%
1-
12
15
#881040000000
0!
0%
b100 *
0-
02
b100 6
#881050000000
1!
1%
1-
12
#881060000000
0!
0%
b101 *
0-
02
b101 6
#881070000000
1!
1%
1-
12
#881080000000
0!
0%
b110 *
0-
02
b110 6
#881090000000
1!
1%
1-
12
#881100000000
0!
0%
b111 *
0-
02
b111 6
#881110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#881120000000
0!
0%
b0 *
0-
02
b0 6
#881130000000
1!
1%
1-
12
#881140000000
0!
0%
b1 *
0-
02
b1 6
#881150000000
1!
1%
1-
12
#881160000000
0!
0%
b10 *
0-
02
b10 6
#881170000000
1!
1%
1-
12
#881180000000
0!
0%
b11 *
0-
02
b11 6
#881190000000
1!
1%
1-
12
15
#881200000000
0!
0%
b100 *
0-
02
b100 6
#881210000000
1!
1%
1-
12
#881220000000
0!
0%
b101 *
0-
02
b101 6
#881230000000
1!
1%
1-
12
#881240000000
0!
0%
b110 *
0-
02
b110 6
#881250000000
1!
1%
1-
12
#881260000000
0!
0%
b111 *
0-
02
b111 6
#881270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#881280000000
0!
0%
b0 *
0-
02
b0 6
#881290000000
1!
1%
1-
12
#881300000000
0!
0%
b1 *
0-
02
b1 6
#881310000000
1!
1%
1-
12
#881320000000
0!
0%
b10 *
0-
02
b10 6
#881330000000
1!
1%
1-
12
#881340000000
0!
0%
b11 *
0-
02
b11 6
#881350000000
1!
1%
1-
12
15
#881360000000
0!
0%
b100 *
0-
02
b100 6
#881370000000
1!
1%
1-
12
#881380000000
0!
0%
b101 *
0-
02
b101 6
#881390000000
1!
1%
1-
12
#881400000000
0!
0%
b110 *
0-
02
b110 6
#881410000000
1!
1%
1-
12
#881420000000
0!
0%
b111 *
0-
02
b111 6
#881430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#881440000000
0!
0%
b0 *
0-
02
b0 6
#881450000000
1!
1%
1-
12
#881460000000
0!
0%
b1 *
0-
02
b1 6
#881470000000
1!
1%
1-
12
#881480000000
0!
0%
b10 *
0-
02
b10 6
#881490000000
1!
1%
1-
12
#881500000000
0!
0%
b11 *
0-
02
b11 6
#881510000000
1!
1%
1-
12
15
#881520000000
0!
0%
b100 *
0-
02
b100 6
#881530000000
1!
1%
1-
12
#881540000000
0!
0%
b101 *
0-
02
b101 6
#881550000000
1!
1%
1-
12
#881560000000
0!
0%
b110 *
0-
02
b110 6
#881570000000
1!
1%
1-
12
#881580000000
0!
0%
b111 *
0-
02
b111 6
#881590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#881600000000
0!
0%
b0 *
0-
02
b0 6
#881610000000
1!
1%
1-
12
#881620000000
0!
0%
b1 *
0-
02
b1 6
#881630000000
1!
1%
1-
12
#881640000000
0!
0%
b10 *
0-
02
b10 6
#881650000000
1!
1%
1-
12
#881660000000
0!
0%
b11 *
0-
02
b11 6
#881670000000
1!
1%
1-
12
15
#881680000000
0!
0%
b100 *
0-
02
b100 6
#881690000000
1!
1%
1-
12
#881700000000
0!
0%
b101 *
0-
02
b101 6
#881710000000
1!
1%
1-
12
#881720000000
0!
0%
b110 *
0-
02
b110 6
#881730000000
1!
1%
1-
12
#881740000000
0!
0%
b111 *
0-
02
b111 6
#881750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#881760000000
0!
0%
b0 *
0-
02
b0 6
#881770000000
1!
1%
1-
12
#881780000000
0!
0%
b1 *
0-
02
b1 6
#881790000000
1!
1%
1-
12
#881800000000
0!
0%
b10 *
0-
02
b10 6
#881810000000
1!
1%
1-
12
#881820000000
0!
0%
b11 *
0-
02
b11 6
#881830000000
1!
1%
1-
12
15
#881840000000
0!
0%
b100 *
0-
02
b100 6
#881850000000
1!
1%
1-
12
#881860000000
0!
0%
b101 *
0-
02
b101 6
#881870000000
1!
1%
1-
12
#881880000000
0!
0%
b110 *
0-
02
b110 6
#881890000000
1!
1%
1-
12
#881900000000
0!
0%
b111 *
0-
02
b111 6
#881910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#881920000000
0!
0%
b0 *
0-
02
b0 6
#881930000000
1!
1%
1-
12
#881940000000
0!
0%
b1 *
0-
02
b1 6
#881950000000
1!
1%
1-
12
#881960000000
0!
0%
b10 *
0-
02
b10 6
#881970000000
1!
1%
1-
12
#881980000000
0!
0%
b11 *
0-
02
b11 6
#881990000000
1!
1%
1-
12
15
#882000000000
0!
0%
b100 *
0-
02
b100 6
#882010000000
1!
1%
1-
12
#882020000000
0!
0%
b101 *
0-
02
b101 6
#882030000000
1!
1%
1-
12
#882040000000
0!
0%
b110 *
0-
02
b110 6
#882050000000
1!
1%
1-
12
#882060000000
0!
0%
b111 *
0-
02
b111 6
#882070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#882080000000
0!
0%
b0 *
0-
02
b0 6
#882090000000
1!
1%
1-
12
#882100000000
0!
0%
b1 *
0-
02
b1 6
#882110000000
1!
1%
1-
12
#882120000000
0!
0%
b10 *
0-
02
b10 6
#882130000000
1!
1%
1-
12
#882140000000
0!
0%
b11 *
0-
02
b11 6
#882150000000
1!
1%
1-
12
15
#882160000000
0!
0%
b100 *
0-
02
b100 6
#882170000000
1!
1%
1-
12
#882180000000
0!
0%
b101 *
0-
02
b101 6
#882190000000
1!
1%
1-
12
#882200000000
0!
0%
b110 *
0-
02
b110 6
#882210000000
1!
1%
1-
12
#882220000000
0!
0%
b111 *
0-
02
b111 6
#882230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#882240000000
0!
0%
b0 *
0-
02
b0 6
#882250000000
1!
1%
1-
12
#882260000000
0!
0%
b1 *
0-
02
b1 6
#882270000000
1!
1%
1-
12
#882280000000
0!
0%
b10 *
0-
02
b10 6
#882290000000
1!
1%
1-
12
#882300000000
0!
0%
b11 *
0-
02
b11 6
#882310000000
1!
1%
1-
12
15
#882320000000
0!
0%
b100 *
0-
02
b100 6
#882330000000
1!
1%
1-
12
#882340000000
0!
0%
b101 *
0-
02
b101 6
#882350000000
1!
1%
1-
12
#882360000000
0!
0%
b110 *
0-
02
b110 6
#882370000000
1!
1%
1-
12
#882380000000
0!
0%
b111 *
0-
02
b111 6
#882390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#882400000000
0!
0%
b0 *
0-
02
b0 6
#882410000000
1!
1%
1-
12
#882420000000
0!
0%
b1 *
0-
02
b1 6
#882430000000
1!
1%
1-
12
#882440000000
0!
0%
b10 *
0-
02
b10 6
#882450000000
1!
1%
1-
12
#882460000000
0!
0%
b11 *
0-
02
b11 6
#882470000000
1!
1%
1-
12
15
#882480000000
0!
0%
b100 *
0-
02
b100 6
#882490000000
1!
1%
1-
12
#882500000000
0!
0%
b101 *
0-
02
b101 6
#882510000000
1!
1%
1-
12
#882520000000
0!
0%
b110 *
0-
02
b110 6
#882530000000
1!
1%
1-
12
#882540000000
0!
0%
b111 *
0-
02
b111 6
#882550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#882560000000
0!
0%
b0 *
0-
02
b0 6
#882570000000
1!
1%
1-
12
#882580000000
0!
0%
b1 *
0-
02
b1 6
#882590000000
1!
1%
1-
12
#882600000000
0!
0%
b10 *
0-
02
b10 6
#882610000000
1!
1%
1-
12
#882620000000
0!
0%
b11 *
0-
02
b11 6
#882630000000
1!
1%
1-
12
15
#882640000000
0!
0%
b100 *
0-
02
b100 6
#882650000000
1!
1%
1-
12
#882660000000
0!
0%
b101 *
0-
02
b101 6
#882670000000
1!
1%
1-
12
#882680000000
0!
0%
b110 *
0-
02
b110 6
#882690000000
1!
1%
1-
12
#882700000000
0!
0%
b111 *
0-
02
b111 6
#882710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#882720000000
0!
0%
b0 *
0-
02
b0 6
#882730000000
1!
1%
1-
12
#882740000000
0!
0%
b1 *
0-
02
b1 6
#882750000000
1!
1%
1-
12
#882760000000
0!
0%
b10 *
0-
02
b10 6
#882770000000
1!
1%
1-
12
#882780000000
0!
0%
b11 *
0-
02
b11 6
#882790000000
1!
1%
1-
12
15
#882800000000
0!
0%
b100 *
0-
02
b100 6
#882810000000
1!
1%
1-
12
#882820000000
0!
0%
b101 *
0-
02
b101 6
#882830000000
1!
1%
1-
12
#882840000000
0!
0%
b110 *
0-
02
b110 6
#882850000000
1!
1%
1-
12
#882860000000
0!
0%
b111 *
0-
02
b111 6
#882870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#882880000000
0!
0%
b0 *
0-
02
b0 6
#882890000000
1!
1%
1-
12
#882900000000
0!
0%
b1 *
0-
02
b1 6
#882910000000
1!
1%
1-
12
#882920000000
0!
0%
b10 *
0-
02
b10 6
#882930000000
1!
1%
1-
12
#882940000000
0!
0%
b11 *
0-
02
b11 6
#882950000000
1!
1%
1-
12
15
#882960000000
0!
0%
b100 *
0-
02
b100 6
#882970000000
1!
1%
1-
12
#882980000000
0!
0%
b101 *
0-
02
b101 6
#882990000000
1!
1%
1-
12
#883000000000
0!
0%
b110 *
0-
02
b110 6
#883010000000
1!
1%
1-
12
#883020000000
0!
0%
b111 *
0-
02
b111 6
#883030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#883040000000
0!
0%
b0 *
0-
02
b0 6
#883050000000
1!
1%
1-
12
#883060000000
0!
0%
b1 *
0-
02
b1 6
#883070000000
1!
1%
1-
12
#883080000000
0!
0%
b10 *
0-
02
b10 6
#883090000000
1!
1%
1-
12
#883100000000
0!
0%
b11 *
0-
02
b11 6
#883110000000
1!
1%
1-
12
15
#883120000000
0!
0%
b100 *
0-
02
b100 6
#883130000000
1!
1%
1-
12
#883140000000
0!
0%
b101 *
0-
02
b101 6
#883150000000
1!
1%
1-
12
#883160000000
0!
0%
b110 *
0-
02
b110 6
#883170000000
1!
1%
1-
12
#883180000000
0!
0%
b111 *
0-
02
b111 6
#883190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#883200000000
0!
0%
b0 *
0-
02
b0 6
#883210000000
1!
1%
1-
12
#883220000000
0!
0%
b1 *
0-
02
b1 6
#883230000000
1!
1%
1-
12
#883240000000
0!
0%
b10 *
0-
02
b10 6
#883250000000
1!
1%
1-
12
#883260000000
0!
0%
b11 *
0-
02
b11 6
#883270000000
1!
1%
1-
12
15
#883280000000
0!
0%
b100 *
0-
02
b100 6
#883290000000
1!
1%
1-
12
#883300000000
0!
0%
b101 *
0-
02
b101 6
#883310000000
1!
1%
1-
12
#883320000000
0!
0%
b110 *
0-
02
b110 6
#883330000000
1!
1%
1-
12
#883340000000
0!
0%
b111 *
0-
02
b111 6
#883350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#883360000000
0!
0%
b0 *
0-
02
b0 6
#883370000000
1!
1%
1-
12
#883380000000
0!
0%
b1 *
0-
02
b1 6
#883390000000
1!
1%
1-
12
#883400000000
0!
0%
b10 *
0-
02
b10 6
#883410000000
1!
1%
1-
12
#883420000000
0!
0%
b11 *
0-
02
b11 6
#883430000000
1!
1%
1-
12
15
#883440000000
0!
0%
b100 *
0-
02
b100 6
#883450000000
1!
1%
1-
12
#883460000000
0!
0%
b101 *
0-
02
b101 6
#883470000000
1!
1%
1-
12
#883480000000
0!
0%
b110 *
0-
02
b110 6
#883490000000
1!
1%
1-
12
#883500000000
0!
0%
b111 *
0-
02
b111 6
#883510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#883520000000
0!
0%
b0 *
0-
02
b0 6
#883530000000
1!
1%
1-
12
#883540000000
0!
0%
b1 *
0-
02
b1 6
#883550000000
1!
1%
1-
12
#883560000000
0!
0%
b10 *
0-
02
b10 6
#883570000000
1!
1%
1-
12
#883580000000
0!
0%
b11 *
0-
02
b11 6
#883590000000
1!
1%
1-
12
15
#883600000000
0!
0%
b100 *
0-
02
b100 6
#883610000000
1!
1%
1-
12
#883620000000
0!
0%
b101 *
0-
02
b101 6
#883630000000
1!
1%
1-
12
#883640000000
0!
0%
b110 *
0-
02
b110 6
#883650000000
1!
1%
1-
12
#883660000000
0!
0%
b111 *
0-
02
b111 6
#883670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#883680000000
0!
0%
b0 *
0-
02
b0 6
#883690000000
1!
1%
1-
12
#883700000000
0!
0%
b1 *
0-
02
b1 6
#883710000000
1!
1%
1-
12
#883720000000
0!
0%
b10 *
0-
02
b10 6
#883730000000
1!
1%
1-
12
#883740000000
0!
0%
b11 *
0-
02
b11 6
#883750000000
1!
1%
1-
12
15
#883760000000
0!
0%
b100 *
0-
02
b100 6
#883770000000
1!
1%
1-
12
#883780000000
0!
0%
b101 *
0-
02
b101 6
#883790000000
1!
1%
1-
12
#883800000000
0!
0%
b110 *
0-
02
b110 6
#883810000000
1!
1%
1-
12
#883820000000
0!
0%
b111 *
0-
02
b111 6
#883830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#883840000000
0!
0%
b0 *
0-
02
b0 6
#883850000000
1!
1%
1-
12
#883860000000
0!
0%
b1 *
0-
02
b1 6
#883870000000
1!
1%
1-
12
#883880000000
0!
0%
b10 *
0-
02
b10 6
#883890000000
1!
1%
1-
12
#883900000000
0!
0%
b11 *
0-
02
b11 6
#883910000000
1!
1%
1-
12
15
#883920000000
0!
0%
b100 *
0-
02
b100 6
#883930000000
1!
1%
1-
12
#883940000000
0!
0%
b101 *
0-
02
b101 6
#883950000000
1!
1%
1-
12
#883960000000
0!
0%
b110 *
0-
02
b110 6
#883970000000
1!
1%
1-
12
#883980000000
0!
0%
b111 *
0-
02
b111 6
#883990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#884000000000
0!
0%
b0 *
0-
02
b0 6
#884010000000
1!
1%
1-
12
#884020000000
0!
0%
b1 *
0-
02
b1 6
#884030000000
1!
1%
1-
12
#884040000000
0!
0%
b10 *
0-
02
b10 6
#884050000000
1!
1%
1-
12
#884060000000
0!
0%
b11 *
0-
02
b11 6
#884070000000
1!
1%
1-
12
15
#884080000000
0!
0%
b100 *
0-
02
b100 6
#884090000000
1!
1%
1-
12
#884100000000
0!
0%
b101 *
0-
02
b101 6
#884110000000
1!
1%
1-
12
#884120000000
0!
0%
b110 *
0-
02
b110 6
#884130000000
1!
1%
1-
12
#884140000000
0!
0%
b111 *
0-
02
b111 6
#884150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#884160000000
0!
0%
b0 *
0-
02
b0 6
#884170000000
1!
1%
1-
12
#884180000000
0!
0%
b1 *
0-
02
b1 6
#884190000000
1!
1%
1-
12
#884200000000
0!
0%
b10 *
0-
02
b10 6
#884210000000
1!
1%
1-
12
#884220000000
0!
0%
b11 *
0-
02
b11 6
#884230000000
1!
1%
1-
12
15
#884240000000
0!
0%
b100 *
0-
02
b100 6
#884250000000
1!
1%
1-
12
#884260000000
0!
0%
b101 *
0-
02
b101 6
#884270000000
1!
1%
1-
12
#884280000000
0!
0%
b110 *
0-
02
b110 6
#884290000000
1!
1%
1-
12
#884300000000
0!
0%
b111 *
0-
02
b111 6
#884310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#884320000000
0!
0%
b0 *
0-
02
b0 6
#884330000000
1!
1%
1-
12
#884340000000
0!
0%
b1 *
0-
02
b1 6
#884350000000
1!
1%
1-
12
#884360000000
0!
0%
b10 *
0-
02
b10 6
#884370000000
1!
1%
1-
12
#884380000000
0!
0%
b11 *
0-
02
b11 6
#884390000000
1!
1%
1-
12
15
#884400000000
0!
0%
b100 *
0-
02
b100 6
#884410000000
1!
1%
1-
12
#884420000000
0!
0%
b101 *
0-
02
b101 6
#884430000000
1!
1%
1-
12
#884440000000
0!
0%
b110 *
0-
02
b110 6
#884450000000
1!
1%
1-
12
#884460000000
0!
0%
b111 *
0-
02
b111 6
#884470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#884480000000
0!
0%
b0 *
0-
02
b0 6
#884490000000
1!
1%
1-
12
#884500000000
0!
0%
b1 *
0-
02
b1 6
#884510000000
1!
1%
1-
12
#884520000000
0!
0%
b10 *
0-
02
b10 6
#884530000000
1!
1%
1-
12
#884540000000
0!
0%
b11 *
0-
02
b11 6
#884550000000
1!
1%
1-
12
15
#884560000000
0!
0%
b100 *
0-
02
b100 6
#884570000000
1!
1%
1-
12
#884580000000
0!
0%
b101 *
0-
02
b101 6
#884590000000
1!
1%
1-
12
#884600000000
0!
0%
b110 *
0-
02
b110 6
#884610000000
1!
1%
1-
12
#884620000000
0!
0%
b111 *
0-
02
b111 6
#884630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#884640000000
0!
0%
b0 *
0-
02
b0 6
#884650000000
1!
1%
1-
12
#884660000000
0!
0%
b1 *
0-
02
b1 6
#884670000000
1!
1%
1-
12
#884680000000
0!
0%
b10 *
0-
02
b10 6
#884690000000
1!
1%
1-
12
#884700000000
0!
0%
b11 *
0-
02
b11 6
#884710000000
1!
1%
1-
12
15
#884720000000
0!
0%
b100 *
0-
02
b100 6
#884730000000
1!
1%
1-
12
#884740000000
0!
0%
b101 *
0-
02
b101 6
#884750000000
1!
1%
1-
12
#884760000000
0!
0%
b110 *
0-
02
b110 6
#884770000000
1!
1%
1-
12
#884780000000
0!
0%
b111 *
0-
02
b111 6
#884790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#884800000000
0!
0%
b0 *
0-
02
b0 6
#884810000000
1!
1%
1-
12
#884820000000
0!
0%
b1 *
0-
02
b1 6
#884830000000
1!
1%
1-
12
#884840000000
0!
0%
b10 *
0-
02
b10 6
#884850000000
1!
1%
1-
12
#884860000000
0!
0%
b11 *
0-
02
b11 6
#884870000000
1!
1%
1-
12
15
#884880000000
0!
0%
b100 *
0-
02
b100 6
#884890000000
1!
1%
1-
12
#884900000000
0!
0%
b101 *
0-
02
b101 6
#884910000000
1!
1%
1-
12
#884920000000
0!
0%
b110 *
0-
02
b110 6
#884930000000
1!
1%
1-
12
#884940000000
0!
0%
b111 *
0-
02
b111 6
#884950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#884960000000
0!
0%
b0 *
0-
02
b0 6
#884970000000
1!
1%
1-
12
#884980000000
0!
0%
b1 *
0-
02
b1 6
#884990000000
1!
1%
1-
12
#885000000000
0!
0%
b10 *
0-
02
b10 6
#885010000000
1!
1%
1-
12
#885020000000
0!
0%
b11 *
0-
02
b11 6
#885030000000
1!
1%
1-
12
15
#885040000000
0!
0%
b100 *
0-
02
b100 6
#885050000000
1!
1%
1-
12
#885060000000
0!
0%
b101 *
0-
02
b101 6
#885070000000
1!
1%
1-
12
#885080000000
0!
0%
b110 *
0-
02
b110 6
#885090000000
1!
1%
1-
12
#885100000000
0!
0%
b111 *
0-
02
b111 6
#885110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#885120000000
0!
0%
b0 *
0-
02
b0 6
#885130000000
1!
1%
1-
12
#885140000000
0!
0%
b1 *
0-
02
b1 6
#885150000000
1!
1%
1-
12
#885160000000
0!
0%
b10 *
0-
02
b10 6
#885170000000
1!
1%
1-
12
#885180000000
0!
0%
b11 *
0-
02
b11 6
#885190000000
1!
1%
1-
12
15
#885200000000
0!
0%
b100 *
0-
02
b100 6
#885210000000
1!
1%
1-
12
#885220000000
0!
0%
b101 *
0-
02
b101 6
#885230000000
1!
1%
1-
12
#885240000000
0!
0%
b110 *
0-
02
b110 6
#885250000000
1!
1%
1-
12
#885260000000
0!
0%
b111 *
0-
02
b111 6
#885270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#885280000000
0!
0%
b0 *
0-
02
b0 6
#885290000000
1!
1%
1-
12
#885300000000
0!
0%
b1 *
0-
02
b1 6
#885310000000
1!
1%
1-
12
#885320000000
0!
0%
b10 *
0-
02
b10 6
#885330000000
1!
1%
1-
12
#885340000000
0!
0%
b11 *
0-
02
b11 6
#885350000000
1!
1%
1-
12
15
#885360000000
0!
0%
b100 *
0-
02
b100 6
#885370000000
1!
1%
1-
12
#885380000000
0!
0%
b101 *
0-
02
b101 6
#885390000000
1!
1%
1-
12
#885400000000
0!
0%
b110 *
0-
02
b110 6
#885410000000
1!
1%
1-
12
#885420000000
0!
0%
b111 *
0-
02
b111 6
#885430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#885440000000
0!
0%
b0 *
0-
02
b0 6
#885450000000
1!
1%
1-
12
#885460000000
0!
0%
b1 *
0-
02
b1 6
#885470000000
1!
1%
1-
12
#885480000000
0!
0%
b10 *
0-
02
b10 6
#885490000000
1!
1%
1-
12
#885500000000
0!
0%
b11 *
0-
02
b11 6
#885510000000
1!
1%
1-
12
15
#885520000000
0!
0%
b100 *
0-
02
b100 6
#885530000000
1!
1%
1-
12
#885540000000
0!
0%
b101 *
0-
02
b101 6
#885550000000
1!
1%
1-
12
#885560000000
0!
0%
b110 *
0-
02
b110 6
#885570000000
1!
1%
1-
12
#885580000000
0!
0%
b111 *
0-
02
b111 6
#885590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#885600000000
0!
0%
b0 *
0-
02
b0 6
#885610000000
1!
1%
1-
12
#885620000000
0!
0%
b1 *
0-
02
b1 6
#885630000000
1!
1%
1-
12
#885640000000
0!
0%
b10 *
0-
02
b10 6
#885650000000
1!
1%
1-
12
#885660000000
0!
0%
b11 *
0-
02
b11 6
#885670000000
1!
1%
1-
12
15
#885680000000
0!
0%
b100 *
0-
02
b100 6
#885690000000
1!
1%
1-
12
#885700000000
0!
0%
b101 *
0-
02
b101 6
#885710000000
1!
1%
1-
12
#885720000000
0!
0%
b110 *
0-
02
b110 6
#885730000000
1!
1%
1-
12
#885740000000
0!
0%
b111 *
0-
02
b111 6
#885750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#885760000000
0!
0%
b0 *
0-
02
b0 6
#885770000000
1!
1%
1-
12
#885780000000
0!
0%
b1 *
0-
02
b1 6
#885790000000
1!
1%
1-
12
#885800000000
0!
0%
b10 *
0-
02
b10 6
#885810000000
1!
1%
1-
12
#885820000000
0!
0%
b11 *
0-
02
b11 6
#885830000000
1!
1%
1-
12
15
#885840000000
0!
0%
b100 *
0-
02
b100 6
#885850000000
1!
1%
1-
12
#885860000000
0!
0%
b101 *
0-
02
b101 6
#885870000000
1!
1%
1-
12
#885880000000
0!
0%
b110 *
0-
02
b110 6
#885890000000
1!
1%
1-
12
#885900000000
0!
0%
b111 *
0-
02
b111 6
#885910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#885920000000
0!
0%
b0 *
0-
02
b0 6
#885930000000
1!
1%
1-
12
#885940000000
0!
0%
b1 *
0-
02
b1 6
#885950000000
1!
1%
1-
12
#885960000000
0!
0%
b10 *
0-
02
b10 6
#885970000000
1!
1%
1-
12
#885980000000
0!
0%
b11 *
0-
02
b11 6
#885990000000
1!
1%
1-
12
15
#886000000000
0!
0%
b100 *
0-
02
b100 6
#886010000000
1!
1%
1-
12
#886020000000
0!
0%
b101 *
0-
02
b101 6
#886030000000
1!
1%
1-
12
#886040000000
0!
0%
b110 *
0-
02
b110 6
#886050000000
1!
1%
1-
12
#886060000000
0!
0%
b111 *
0-
02
b111 6
#886070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#886080000000
0!
0%
b0 *
0-
02
b0 6
#886090000000
1!
1%
1-
12
#886100000000
0!
0%
b1 *
0-
02
b1 6
#886110000000
1!
1%
1-
12
#886120000000
0!
0%
b10 *
0-
02
b10 6
#886130000000
1!
1%
1-
12
#886140000000
0!
0%
b11 *
0-
02
b11 6
#886150000000
1!
1%
1-
12
15
#886160000000
0!
0%
b100 *
0-
02
b100 6
#886170000000
1!
1%
1-
12
#886180000000
0!
0%
b101 *
0-
02
b101 6
#886190000000
1!
1%
1-
12
#886200000000
0!
0%
b110 *
0-
02
b110 6
#886210000000
1!
1%
1-
12
#886220000000
0!
0%
b111 *
0-
02
b111 6
#886230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#886240000000
0!
0%
b0 *
0-
02
b0 6
#886250000000
1!
1%
1-
12
#886260000000
0!
0%
b1 *
0-
02
b1 6
#886270000000
1!
1%
1-
12
#886280000000
0!
0%
b10 *
0-
02
b10 6
#886290000000
1!
1%
1-
12
#886300000000
0!
0%
b11 *
0-
02
b11 6
#886310000000
1!
1%
1-
12
15
#886320000000
0!
0%
b100 *
0-
02
b100 6
#886330000000
1!
1%
1-
12
#886340000000
0!
0%
b101 *
0-
02
b101 6
#886350000000
1!
1%
1-
12
#886360000000
0!
0%
b110 *
0-
02
b110 6
#886370000000
1!
1%
1-
12
#886380000000
0!
0%
b111 *
0-
02
b111 6
#886390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#886400000000
0!
0%
b0 *
0-
02
b0 6
#886410000000
1!
1%
1-
12
#886420000000
0!
0%
b1 *
0-
02
b1 6
#886430000000
1!
1%
1-
12
#886440000000
0!
0%
b10 *
0-
02
b10 6
#886450000000
1!
1%
1-
12
#886460000000
0!
0%
b11 *
0-
02
b11 6
#886470000000
1!
1%
1-
12
15
#886480000000
0!
0%
b100 *
0-
02
b100 6
#886490000000
1!
1%
1-
12
#886500000000
0!
0%
b101 *
0-
02
b101 6
#886510000000
1!
1%
1-
12
#886520000000
0!
0%
b110 *
0-
02
b110 6
#886530000000
1!
1%
1-
12
#886540000000
0!
0%
b111 *
0-
02
b111 6
#886550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#886560000000
0!
0%
b0 *
0-
02
b0 6
#886570000000
1!
1%
1-
12
#886580000000
0!
0%
b1 *
0-
02
b1 6
#886590000000
1!
1%
1-
12
#886600000000
0!
0%
b10 *
0-
02
b10 6
#886610000000
1!
1%
1-
12
#886620000000
0!
0%
b11 *
0-
02
b11 6
#886630000000
1!
1%
1-
12
15
#886640000000
0!
0%
b100 *
0-
02
b100 6
#886650000000
1!
1%
1-
12
#886660000000
0!
0%
b101 *
0-
02
b101 6
#886670000000
1!
1%
1-
12
#886680000000
0!
0%
b110 *
0-
02
b110 6
#886690000000
1!
1%
1-
12
#886700000000
0!
0%
b111 *
0-
02
b111 6
#886710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#886720000000
0!
0%
b0 *
0-
02
b0 6
#886730000000
1!
1%
1-
12
#886740000000
0!
0%
b1 *
0-
02
b1 6
#886750000000
1!
1%
1-
12
#886760000000
0!
0%
b10 *
0-
02
b10 6
#886770000000
1!
1%
1-
12
#886780000000
0!
0%
b11 *
0-
02
b11 6
#886790000000
1!
1%
1-
12
15
#886800000000
0!
0%
b100 *
0-
02
b100 6
#886810000000
1!
1%
1-
12
#886820000000
0!
0%
b101 *
0-
02
b101 6
#886830000000
1!
1%
1-
12
#886840000000
0!
0%
b110 *
0-
02
b110 6
#886850000000
1!
1%
1-
12
#886860000000
0!
0%
b111 *
0-
02
b111 6
#886870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#886880000000
0!
0%
b0 *
0-
02
b0 6
#886890000000
1!
1%
1-
12
#886900000000
0!
0%
b1 *
0-
02
b1 6
#886910000000
1!
1%
1-
12
#886920000000
0!
0%
b10 *
0-
02
b10 6
#886930000000
1!
1%
1-
12
#886940000000
0!
0%
b11 *
0-
02
b11 6
#886950000000
1!
1%
1-
12
15
#886960000000
0!
0%
b100 *
0-
02
b100 6
#886970000000
1!
1%
1-
12
#886980000000
0!
0%
b101 *
0-
02
b101 6
#886990000000
1!
1%
1-
12
#887000000000
0!
0%
b110 *
0-
02
b110 6
#887010000000
1!
1%
1-
12
#887020000000
0!
0%
b111 *
0-
02
b111 6
#887030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#887040000000
0!
0%
b0 *
0-
02
b0 6
#887050000000
1!
1%
1-
12
#887060000000
0!
0%
b1 *
0-
02
b1 6
#887070000000
1!
1%
1-
12
#887080000000
0!
0%
b10 *
0-
02
b10 6
#887090000000
1!
1%
1-
12
#887100000000
0!
0%
b11 *
0-
02
b11 6
#887110000000
1!
1%
1-
12
15
#887120000000
0!
0%
b100 *
0-
02
b100 6
#887130000000
1!
1%
1-
12
#887140000000
0!
0%
b101 *
0-
02
b101 6
#887150000000
1!
1%
1-
12
#887160000000
0!
0%
b110 *
0-
02
b110 6
#887170000000
1!
1%
1-
12
#887180000000
0!
0%
b111 *
0-
02
b111 6
#887190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#887200000000
0!
0%
b0 *
0-
02
b0 6
#887210000000
1!
1%
1-
12
#887220000000
0!
0%
b1 *
0-
02
b1 6
#887230000000
1!
1%
1-
12
#887240000000
0!
0%
b10 *
0-
02
b10 6
#887250000000
1!
1%
1-
12
#887260000000
0!
0%
b11 *
0-
02
b11 6
#887270000000
1!
1%
1-
12
15
#887280000000
0!
0%
b100 *
0-
02
b100 6
#887290000000
1!
1%
1-
12
#887300000000
0!
0%
b101 *
0-
02
b101 6
#887310000000
1!
1%
1-
12
#887320000000
0!
0%
b110 *
0-
02
b110 6
#887330000000
1!
1%
1-
12
#887340000000
0!
0%
b111 *
0-
02
b111 6
#887350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#887360000000
0!
0%
b0 *
0-
02
b0 6
#887370000000
1!
1%
1-
12
#887380000000
0!
0%
b1 *
0-
02
b1 6
#887390000000
1!
1%
1-
12
#887400000000
0!
0%
b10 *
0-
02
b10 6
#887410000000
1!
1%
1-
12
#887420000000
0!
0%
b11 *
0-
02
b11 6
#887430000000
1!
1%
1-
12
15
#887440000000
0!
0%
b100 *
0-
02
b100 6
#887450000000
1!
1%
1-
12
#887460000000
0!
0%
b101 *
0-
02
b101 6
#887470000000
1!
1%
1-
12
#887480000000
0!
0%
b110 *
0-
02
b110 6
#887490000000
1!
1%
1-
12
#887500000000
0!
0%
b111 *
0-
02
b111 6
#887510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#887520000000
0!
0%
b0 *
0-
02
b0 6
#887530000000
1!
1%
1-
12
#887540000000
0!
0%
b1 *
0-
02
b1 6
#887550000000
1!
1%
1-
12
#887560000000
0!
0%
b10 *
0-
02
b10 6
#887570000000
1!
1%
1-
12
#887580000000
0!
0%
b11 *
0-
02
b11 6
#887590000000
1!
1%
1-
12
15
#887600000000
0!
0%
b100 *
0-
02
b100 6
#887610000000
1!
1%
1-
12
#887620000000
0!
0%
b101 *
0-
02
b101 6
#887630000000
1!
1%
1-
12
#887640000000
0!
0%
b110 *
0-
02
b110 6
#887650000000
1!
1%
1-
12
#887660000000
0!
0%
b111 *
0-
02
b111 6
#887670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#887680000000
0!
0%
b0 *
0-
02
b0 6
#887690000000
1!
1%
1-
12
#887700000000
0!
0%
b1 *
0-
02
b1 6
#887710000000
1!
1%
1-
12
#887720000000
0!
0%
b10 *
0-
02
b10 6
#887730000000
1!
1%
1-
12
#887740000000
0!
0%
b11 *
0-
02
b11 6
#887750000000
1!
1%
1-
12
15
#887760000000
0!
0%
b100 *
0-
02
b100 6
#887770000000
1!
1%
1-
12
#887780000000
0!
0%
b101 *
0-
02
b101 6
#887790000000
1!
1%
1-
12
#887800000000
0!
0%
b110 *
0-
02
b110 6
#887810000000
1!
1%
1-
12
#887820000000
0!
0%
b111 *
0-
02
b111 6
#887830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#887840000000
0!
0%
b0 *
0-
02
b0 6
#887850000000
1!
1%
1-
12
#887860000000
0!
0%
b1 *
0-
02
b1 6
#887870000000
1!
1%
1-
12
#887880000000
0!
0%
b10 *
0-
02
b10 6
#887890000000
1!
1%
1-
12
#887900000000
0!
0%
b11 *
0-
02
b11 6
#887910000000
1!
1%
1-
12
15
#887920000000
0!
0%
b100 *
0-
02
b100 6
#887930000000
1!
1%
1-
12
#887940000000
0!
0%
b101 *
0-
02
b101 6
#887950000000
1!
1%
1-
12
#887960000000
0!
0%
b110 *
0-
02
b110 6
#887970000000
1!
1%
1-
12
#887980000000
0!
0%
b111 *
0-
02
b111 6
#887990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#888000000000
0!
0%
b0 *
0-
02
b0 6
#888010000000
1!
1%
1-
12
#888020000000
0!
0%
b1 *
0-
02
b1 6
#888030000000
1!
1%
1-
12
#888040000000
0!
0%
b10 *
0-
02
b10 6
#888050000000
1!
1%
1-
12
#888060000000
0!
0%
b11 *
0-
02
b11 6
#888070000000
1!
1%
1-
12
15
#888080000000
0!
0%
b100 *
0-
02
b100 6
#888090000000
1!
1%
1-
12
#888100000000
0!
0%
b101 *
0-
02
b101 6
#888110000000
1!
1%
1-
12
#888120000000
0!
0%
b110 *
0-
02
b110 6
#888130000000
1!
1%
1-
12
#888140000000
0!
0%
b111 *
0-
02
b111 6
#888150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#888160000000
0!
0%
b0 *
0-
02
b0 6
#888170000000
1!
1%
1-
12
#888180000000
0!
0%
b1 *
0-
02
b1 6
#888190000000
1!
1%
1-
12
#888200000000
0!
0%
b10 *
0-
02
b10 6
#888210000000
1!
1%
1-
12
#888220000000
0!
0%
b11 *
0-
02
b11 6
#888230000000
1!
1%
1-
12
15
#888240000000
0!
0%
b100 *
0-
02
b100 6
#888250000000
1!
1%
1-
12
#888260000000
0!
0%
b101 *
0-
02
b101 6
#888270000000
1!
1%
1-
12
#888280000000
0!
0%
b110 *
0-
02
b110 6
#888290000000
1!
1%
1-
12
#888300000000
0!
0%
b111 *
0-
02
b111 6
#888310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#888320000000
0!
0%
b0 *
0-
02
b0 6
#888330000000
1!
1%
1-
12
#888340000000
0!
0%
b1 *
0-
02
b1 6
#888350000000
1!
1%
1-
12
#888360000000
0!
0%
b10 *
0-
02
b10 6
#888370000000
1!
1%
1-
12
#888380000000
0!
0%
b11 *
0-
02
b11 6
#888390000000
1!
1%
1-
12
15
#888400000000
0!
0%
b100 *
0-
02
b100 6
#888410000000
1!
1%
1-
12
#888420000000
0!
0%
b101 *
0-
02
b101 6
#888430000000
1!
1%
1-
12
#888440000000
0!
0%
b110 *
0-
02
b110 6
#888450000000
1!
1%
1-
12
#888460000000
0!
0%
b111 *
0-
02
b111 6
#888470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#888480000000
0!
0%
b0 *
0-
02
b0 6
#888490000000
1!
1%
1-
12
#888500000000
0!
0%
b1 *
0-
02
b1 6
#888510000000
1!
1%
1-
12
#888520000000
0!
0%
b10 *
0-
02
b10 6
#888530000000
1!
1%
1-
12
#888540000000
0!
0%
b11 *
0-
02
b11 6
#888550000000
1!
1%
1-
12
15
#888560000000
0!
0%
b100 *
0-
02
b100 6
#888570000000
1!
1%
1-
12
#888580000000
0!
0%
b101 *
0-
02
b101 6
#888590000000
1!
1%
1-
12
#888600000000
0!
0%
b110 *
0-
02
b110 6
#888610000000
1!
1%
1-
12
#888620000000
0!
0%
b111 *
0-
02
b111 6
#888630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#888640000000
0!
0%
b0 *
0-
02
b0 6
#888650000000
1!
1%
1-
12
#888660000000
0!
0%
b1 *
0-
02
b1 6
#888670000000
1!
1%
1-
12
#888680000000
0!
0%
b10 *
0-
02
b10 6
#888690000000
1!
1%
1-
12
#888700000000
0!
0%
b11 *
0-
02
b11 6
#888710000000
1!
1%
1-
12
15
#888720000000
0!
0%
b100 *
0-
02
b100 6
#888730000000
1!
1%
1-
12
#888740000000
0!
0%
b101 *
0-
02
b101 6
#888750000000
1!
1%
1-
12
#888760000000
0!
0%
b110 *
0-
02
b110 6
#888770000000
1!
1%
1-
12
#888780000000
0!
0%
b111 *
0-
02
b111 6
#888790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#888800000000
0!
0%
b0 *
0-
02
b0 6
#888810000000
1!
1%
1-
12
#888820000000
0!
0%
b1 *
0-
02
b1 6
#888830000000
1!
1%
1-
12
#888840000000
0!
0%
b10 *
0-
02
b10 6
#888850000000
1!
1%
1-
12
#888860000000
0!
0%
b11 *
0-
02
b11 6
#888870000000
1!
1%
1-
12
15
#888880000000
0!
0%
b100 *
0-
02
b100 6
#888890000000
1!
1%
1-
12
#888900000000
0!
0%
b101 *
0-
02
b101 6
#888910000000
1!
1%
1-
12
#888920000000
0!
0%
b110 *
0-
02
b110 6
#888930000000
1!
1%
1-
12
#888940000000
0!
0%
b111 *
0-
02
b111 6
#888950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#888960000000
0!
0%
b0 *
0-
02
b0 6
#888970000000
1!
1%
1-
12
#888980000000
0!
0%
b1 *
0-
02
b1 6
#888990000000
1!
1%
1-
12
#889000000000
0!
0%
b10 *
0-
02
b10 6
#889010000000
1!
1%
1-
12
#889020000000
0!
0%
b11 *
0-
02
b11 6
#889030000000
1!
1%
1-
12
15
#889040000000
0!
0%
b100 *
0-
02
b100 6
#889050000000
1!
1%
1-
12
#889060000000
0!
0%
b101 *
0-
02
b101 6
#889070000000
1!
1%
1-
12
#889080000000
0!
0%
b110 *
0-
02
b110 6
#889090000000
1!
1%
1-
12
#889100000000
0!
0%
b111 *
0-
02
b111 6
#889110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#889120000000
0!
0%
b0 *
0-
02
b0 6
#889130000000
1!
1%
1-
12
#889140000000
0!
0%
b1 *
0-
02
b1 6
#889150000000
1!
1%
1-
12
#889160000000
0!
0%
b10 *
0-
02
b10 6
#889170000000
1!
1%
1-
12
#889180000000
0!
0%
b11 *
0-
02
b11 6
#889190000000
1!
1%
1-
12
15
#889200000000
0!
0%
b100 *
0-
02
b100 6
#889210000000
1!
1%
1-
12
#889220000000
0!
0%
b101 *
0-
02
b101 6
#889230000000
1!
1%
1-
12
#889240000000
0!
0%
b110 *
0-
02
b110 6
#889250000000
1!
1%
1-
12
#889260000000
0!
0%
b111 *
0-
02
b111 6
#889270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#889280000000
0!
0%
b0 *
0-
02
b0 6
#889290000000
1!
1%
1-
12
#889300000000
0!
0%
b1 *
0-
02
b1 6
#889310000000
1!
1%
1-
12
#889320000000
0!
0%
b10 *
0-
02
b10 6
#889330000000
1!
1%
1-
12
#889340000000
0!
0%
b11 *
0-
02
b11 6
#889350000000
1!
1%
1-
12
15
#889360000000
0!
0%
b100 *
0-
02
b100 6
#889370000000
1!
1%
1-
12
#889380000000
0!
0%
b101 *
0-
02
b101 6
#889390000000
1!
1%
1-
12
#889400000000
0!
0%
b110 *
0-
02
b110 6
#889410000000
1!
1%
1-
12
#889420000000
0!
0%
b111 *
0-
02
b111 6
#889430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#889440000000
0!
0%
b0 *
0-
02
b0 6
#889450000000
1!
1%
1-
12
#889460000000
0!
0%
b1 *
0-
02
b1 6
#889470000000
1!
1%
1-
12
#889480000000
0!
0%
b10 *
0-
02
b10 6
#889490000000
1!
1%
1-
12
#889500000000
0!
0%
b11 *
0-
02
b11 6
#889510000000
1!
1%
1-
12
15
#889520000000
0!
0%
b100 *
0-
02
b100 6
#889530000000
1!
1%
1-
12
#889540000000
0!
0%
b101 *
0-
02
b101 6
#889550000000
1!
1%
1-
12
#889560000000
0!
0%
b110 *
0-
02
b110 6
#889570000000
1!
1%
1-
12
#889580000000
0!
0%
b111 *
0-
02
b111 6
#889590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#889600000000
0!
0%
b0 *
0-
02
b0 6
#889610000000
1!
1%
1-
12
#889620000000
0!
0%
b1 *
0-
02
b1 6
#889630000000
1!
1%
1-
12
#889640000000
0!
0%
b10 *
0-
02
b10 6
#889650000000
1!
1%
1-
12
#889660000000
0!
0%
b11 *
0-
02
b11 6
#889670000000
1!
1%
1-
12
15
#889680000000
0!
0%
b100 *
0-
02
b100 6
#889690000000
1!
1%
1-
12
#889700000000
0!
0%
b101 *
0-
02
b101 6
#889710000000
1!
1%
1-
12
#889720000000
0!
0%
b110 *
0-
02
b110 6
#889730000000
1!
1%
1-
12
#889740000000
0!
0%
b111 *
0-
02
b111 6
#889750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#889760000000
0!
0%
b0 *
0-
02
b0 6
#889770000000
1!
1%
1-
12
#889780000000
0!
0%
b1 *
0-
02
b1 6
#889790000000
1!
1%
1-
12
#889800000000
0!
0%
b10 *
0-
02
b10 6
#889810000000
1!
1%
1-
12
#889820000000
0!
0%
b11 *
0-
02
b11 6
#889830000000
1!
1%
1-
12
15
#889840000000
0!
0%
b100 *
0-
02
b100 6
#889850000000
1!
1%
1-
12
#889860000000
0!
0%
b101 *
0-
02
b101 6
#889870000000
1!
1%
1-
12
#889880000000
0!
0%
b110 *
0-
02
b110 6
#889890000000
1!
1%
1-
12
#889900000000
0!
0%
b111 *
0-
02
b111 6
#889910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#889920000000
0!
0%
b0 *
0-
02
b0 6
#889930000000
1!
1%
1-
12
#889940000000
0!
0%
b1 *
0-
02
b1 6
#889950000000
1!
1%
1-
12
#889960000000
0!
0%
b10 *
0-
02
b10 6
#889970000000
1!
1%
1-
12
#889980000000
0!
0%
b11 *
0-
02
b11 6
#889990000000
1!
1%
1-
12
15
#890000000000
0!
0%
b100 *
0-
02
b100 6
#890010000000
1!
1%
1-
12
#890020000000
0!
0%
b101 *
0-
02
b101 6
#890030000000
1!
1%
1-
12
#890040000000
0!
0%
b110 *
0-
02
b110 6
#890050000000
1!
1%
1-
12
#890060000000
0!
0%
b111 *
0-
02
b111 6
#890070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#890080000000
0!
0%
b0 *
0-
02
b0 6
#890090000000
1!
1%
1-
12
#890100000000
0!
0%
b1 *
0-
02
b1 6
#890110000000
1!
1%
1-
12
#890120000000
0!
0%
b10 *
0-
02
b10 6
#890130000000
1!
1%
1-
12
#890140000000
0!
0%
b11 *
0-
02
b11 6
#890150000000
1!
1%
1-
12
15
#890160000000
0!
0%
b100 *
0-
02
b100 6
#890170000000
1!
1%
1-
12
#890180000000
0!
0%
b101 *
0-
02
b101 6
#890190000000
1!
1%
1-
12
#890200000000
0!
0%
b110 *
0-
02
b110 6
#890210000000
1!
1%
1-
12
#890220000000
0!
0%
b111 *
0-
02
b111 6
#890230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#890240000000
0!
0%
b0 *
0-
02
b0 6
#890250000000
1!
1%
1-
12
#890260000000
0!
0%
b1 *
0-
02
b1 6
#890270000000
1!
1%
1-
12
#890280000000
0!
0%
b10 *
0-
02
b10 6
#890290000000
1!
1%
1-
12
#890300000000
0!
0%
b11 *
0-
02
b11 6
#890310000000
1!
1%
1-
12
15
#890320000000
0!
0%
b100 *
0-
02
b100 6
#890330000000
1!
1%
1-
12
#890340000000
0!
0%
b101 *
0-
02
b101 6
#890350000000
1!
1%
1-
12
#890360000000
0!
0%
b110 *
0-
02
b110 6
#890370000000
1!
1%
1-
12
#890380000000
0!
0%
b111 *
0-
02
b111 6
#890390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#890400000000
0!
0%
b0 *
0-
02
b0 6
#890410000000
1!
1%
1-
12
#890420000000
0!
0%
b1 *
0-
02
b1 6
#890430000000
1!
1%
1-
12
#890440000000
0!
0%
b10 *
0-
02
b10 6
#890450000000
1!
1%
1-
12
#890460000000
0!
0%
b11 *
0-
02
b11 6
#890470000000
1!
1%
1-
12
15
#890480000000
0!
0%
b100 *
0-
02
b100 6
#890490000000
1!
1%
1-
12
#890500000000
0!
0%
b101 *
0-
02
b101 6
#890510000000
1!
1%
1-
12
#890520000000
0!
0%
b110 *
0-
02
b110 6
#890530000000
1!
1%
1-
12
#890540000000
0!
0%
b111 *
0-
02
b111 6
#890550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#890560000000
0!
0%
b0 *
0-
02
b0 6
#890570000000
1!
1%
1-
12
#890580000000
0!
0%
b1 *
0-
02
b1 6
#890590000000
1!
1%
1-
12
#890600000000
0!
0%
b10 *
0-
02
b10 6
#890610000000
1!
1%
1-
12
#890620000000
0!
0%
b11 *
0-
02
b11 6
#890630000000
1!
1%
1-
12
15
#890640000000
0!
0%
b100 *
0-
02
b100 6
#890650000000
1!
1%
1-
12
#890660000000
0!
0%
b101 *
0-
02
b101 6
#890670000000
1!
1%
1-
12
#890680000000
0!
0%
b110 *
0-
02
b110 6
#890690000000
1!
1%
1-
12
#890700000000
0!
0%
b111 *
0-
02
b111 6
#890710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#890720000000
0!
0%
b0 *
0-
02
b0 6
#890730000000
1!
1%
1-
12
#890740000000
0!
0%
b1 *
0-
02
b1 6
#890750000000
1!
1%
1-
12
#890760000000
0!
0%
b10 *
0-
02
b10 6
#890770000000
1!
1%
1-
12
#890780000000
0!
0%
b11 *
0-
02
b11 6
#890790000000
1!
1%
1-
12
15
#890800000000
0!
0%
b100 *
0-
02
b100 6
#890810000000
1!
1%
1-
12
#890820000000
0!
0%
b101 *
0-
02
b101 6
#890830000000
1!
1%
1-
12
#890840000000
0!
0%
b110 *
0-
02
b110 6
#890850000000
1!
1%
1-
12
#890860000000
0!
0%
b111 *
0-
02
b111 6
#890870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#890880000000
0!
0%
b0 *
0-
02
b0 6
#890890000000
1!
1%
1-
12
#890900000000
0!
0%
b1 *
0-
02
b1 6
#890910000000
1!
1%
1-
12
#890920000000
0!
0%
b10 *
0-
02
b10 6
#890930000000
1!
1%
1-
12
#890940000000
0!
0%
b11 *
0-
02
b11 6
#890950000000
1!
1%
1-
12
15
#890960000000
0!
0%
b100 *
0-
02
b100 6
#890970000000
1!
1%
1-
12
#890980000000
0!
0%
b101 *
0-
02
b101 6
#890990000000
1!
1%
1-
12
#891000000000
0!
0%
b110 *
0-
02
b110 6
#891010000000
1!
1%
1-
12
#891020000000
0!
0%
b111 *
0-
02
b111 6
#891030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#891040000000
0!
0%
b0 *
0-
02
b0 6
#891050000000
1!
1%
1-
12
#891060000000
0!
0%
b1 *
0-
02
b1 6
#891070000000
1!
1%
1-
12
#891080000000
0!
0%
b10 *
0-
02
b10 6
#891090000000
1!
1%
1-
12
#891100000000
0!
0%
b11 *
0-
02
b11 6
#891110000000
1!
1%
1-
12
15
#891120000000
0!
0%
b100 *
0-
02
b100 6
#891130000000
1!
1%
1-
12
#891140000000
0!
0%
b101 *
0-
02
b101 6
#891150000000
1!
1%
1-
12
#891160000000
0!
0%
b110 *
0-
02
b110 6
#891170000000
1!
1%
1-
12
#891180000000
0!
0%
b111 *
0-
02
b111 6
#891190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#891200000000
0!
0%
b0 *
0-
02
b0 6
#891210000000
1!
1%
1-
12
#891220000000
0!
0%
b1 *
0-
02
b1 6
#891230000000
1!
1%
1-
12
#891240000000
0!
0%
b10 *
0-
02
b10 6
#891250000000
1!
1%
1-
12
#891260000000
0!
0%
b11 *
0-
02
b11 6
#891270000000
1!
1%
1-
12
15
#891280000000
0!
0%
b100 *
0-
02
b100 6
#891290000000
1!
1%
1-
12
#891300000000
0!
0%
b101 *
0-
02
b101 6
#891310000000
1!
1%
1-
12
#891320000000
0!
0%
b110 *
0-
02
b110 6
#891330000000
1!
1%
1-
12
#891340000000
0!
0%
b111 *
0-
02
b111 6
#891350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#891360000000
0!
0%
b0 *
0-
02
b0 6
#891370000000
1!
1%
1-
12
#891380000000
0!
0%
b1 *
0-
02
b1 6
#891390000000
1!
1%
1-
12
#891400000000
0!
0%
b10 *
0-
02
b10 6
#891410000000
1!
1%
1-
12
#891420000000
0!
0%
b11 *
0-
02
b11 6
#891430000000
1!
1%
1-
12
15
#891440000000
0!
0%
b100 *
0-
02
b100 6
#891450000000
1!
1%
1-
12
#891460000000
0!
0%
b101 *
0-
02
b101 6
#891470000000
1!
1%
1-
12
#891480000000
0!
0%
b110 *
0-
02
b110 6
#891490000000
1!
1%
1-
12
#891500000000
0!
0%
b111 *
0-
02
b111 6
#891510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#891520000000
0!
0%
b0 *
0-
02
b0 6
#891530000000
1!
1%
1-
12
#891540000000
0!
0%
b1 *
0-
02
b1 6
#891550000000
1!
1%
1-
12
#891560000000
0!
0%
b10 *
0-
02
b10 6
#891570000000
1!
1%
1-
12
#891580000000
0!
0%
b11 *
0-
02
b11 6
#891590000000
1!
1%
1-
12
15
#891600000000
0!
0%
b100 *
0-
02
b100 6
#891610000000
1!
1%
1-
12
#891620000000
0!
0%
b101 *
0-
02
b101 6
#891630000000
1!
1%
1-
12
#891640000000
0!
0%
b110 *
0-
02
b110 6
#891650000000
1!
1%
1-
12
#891660000000
0!
0%
b111 *
0-
02
b111 6
#891670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#891680000000
0!
0%
b0 *
0-
02
b0 6
#891690000000
1!
1%
1-
12
#891700000000
0!
0%
b1 *
0-
02
b1 6
#891710000000
1!
1%
1-
12
#891720000000
0!
0%
b10 *
0-
02
b10 6
#891730000000
1!
1%
1-
12
#891740000000
0!
0%
b11 *
0-
02
b11 6
#891750000000
1!
1%
1-
12
15
#891760000000
0!
0%
b100 *
0-
02
b100 6
#891770000000
1!
1%
1-
12
#891780000000
0!
0%
b101 *
0-
02
b101 6
#891790000000
1!
1%
1-
12
#891800000000
0!
0%
b110 *
0-
02
b110 6
#891810000000
1!
1%
1-
12
#891820000000
0!
0%
b111 *
0-
02
b111 6
#891830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#891840000000
0!
0%
b0 *
0-
02
b0 6
#891850000000
1!
1%
1-
12
#891860000000
0!
0%
b1 *
0-
02
b1 6
#891870000000
1!
1%
1-
12
#891880000000
0!
0%
b10 *
0-
02
b10 6
#891890000000
1!
1%
1-
12
#891900000000
0!
0%
b11 *
0-
02
b11 6
#891910000000
1!
1%
1-
12
15
#891920000000
0!
0%
b100 *
0-
02
b100 6
#891930000000
1!
1%
1-
12
#891940000000
0!
0%
b101 *
0-
02
b101 6
#891950000000
1!
1%
1-
12
#891960000000
0!
0%
b110 *
0-
02
b110 6
#891970000000
1!
1%
1-
12
#891980000000
0!
0%
b111 *
0-
02
b111 6
#891990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#892000000000
0!
0%
b0 *
0-
02
b0 6
#892010000000
1!
1%
1-
12
#892020000000
0!
0%
b1 *
0-
02
b1 6
#892030000000
1!
1%
1-
12
#892040000000
0!
0%
b10 *
0-
02
b10 6
#892050000000
1!
1%
1-
12
#892060000000
0!
0%
b11 *
0-
02
b11 6
#892070000000
1!
1%
1-
12
15
#892080000000
0!
0%
b100 *
0-
02
b100 6
#892090000000
1!
1%
1-
12
#892100000000
0!
0%
b101 *
0-
02
b101 6
#892110000000
1!
1%
1-
12
#892120000000
0!
0%
b110 *
0-
02
b110 6
#892130000000
1!
1%
1-
12
#892140000000
0!
0%
b111 *
0-
02
b111 6
#892150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#892160000000
0!
0%
b0 *
0-
02
b0 6
#892170000000
1!
1%
1-
12
#892180000000
0!
0%
b1 *
0-
02
b1 6
#892190000000
1!
1%
1-
12
#892200000000
0!
0%
b10 *
0-
02
b10 6
#892210000000
1!
1%
1-
12
#892220000000
0!
0%
b11 *
0-
02
b11 6
#892230000000
1!
1%
1-
12
15
#892240000000
0!
0%
b100 *
0-
02
b100 6
#892250000000
1!
1%
1-
12
#892260000000
0!
0%
b101 *
0-
02
b101 6
#892270000000
1!
1%
1-
12
#892280000000
0!
0%
b110 *
0-
02
b110 6
#892290000000
1!
1%
1-
12
#892300000000
0!
0%
b111 *
0-
02
b111 6
#892310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#892320000000
0!
0%
b0 *
0-
02
b0 6
#892330000000
1!
1%
1-
12
#892340000000
0!
0%
b1 *
0-
02
b1 6
#892350000000
1!
1%
1-
12
#892360000000
0!
0%
b10 *
0-
02
b10 6
#892370000000
1!
1%
1-
12
#892380000000
0!
0%
b11 *
0-
02
b11 6
#892390000000
1!
1%
1-
12
15
#892400000000
0!
0%
b100 *
0-
02
b100 6
#892410000000
1!
1%
1-
12
#892420000000
0!
0%
b101 *
0-
02
b101 6
#892430000000
1!
1%
1-
12
#892440000000
0!
0%
b110 *
0-
02
b110 6
#892450000000
1!
1%
1-
12
#892460000000
0!
0%
b111 *
0-
02
b111 6
#892470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#892480000000
0!
0%
b0 *
0-
02
b0 6
#892490000000
1!
1%
1-
12
#892500000000
0!
0%
b1 *
0-
02
b1 6
#892510000000
1!
1%
1-
12
#892520000000
0!
0%
b10 *
0-
02
b10 6
#892530000000
1!
1%
1-
12
#892540000000
0!
0%
b11 *
0-
02
b11 6
#892550000000
1!
1%
1-
12
15
#892560000000
0!
0%
b100 *
0-
02
b100 6
#892570000000
1!
1%
1-
12
#892580000000
0!
0%
b101 *
0-
02
b101 6
#892590000000
1!
1%
1-
12
#892600000000
0!
0%
b110 *
0-
02
b110 6
#892610000000
1!
1%
1-
12
#892620000000
0!
0%
b111 *
0-
02
b111 6
#892630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#892640000000
0!
0%
b0 *
0-
02
b0 6
#892650000000
1!
1%
1-
12
#892660000000
0!
0%
b1 *
0-
02
b1 6
#892670000000
1!
1%
1-
12
#892680000000
0!
0%
b10 *
0-
02
b10 6
#892690000000
1!
1%
1-
12
#892700000000
0!
0%
b11 *
0-
02
b11 6
#892710000000
1!
1%
1-
12
15
#892720000000
0!
0%
b100 *
0-
02
b100 6
#892730000000
1!
1%
1-
12
#892740000000
0!
0%
b101 *
0-
02
b101 6
#892750000000
1!
1%
1-
12
#892760000000
0!
0%
b110 *
0-
02
b110 6
#892770000000
1!
1%
1-
12
#892780000000
0!
0%
b111 *
0-
02
b111 6
#892790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#892800000000
0!
0%
b0 *
0-
02
b0 6
#892810000000
1!
1%
1-
12
#892820000000
0!
0%
b1 *
0-
02
b1 6
#892830000000
1!
1%
1-
12
#892840000000
0!
0%
b10 *
0-
02
b10 6
#892850000000
1!
1%
1-
12
#892860000000
0!
0%
b11 *
0-
02
b11 6
#892870000000
1!
1%
1-
12
15
#892880000000
0!
0%
b100 *
0-
02
b100 6
#892890000000
1!
1%
1-
12
#892900000000
0!
0%
b101 *
0-
02
b101 6
#892910000000
1!
1%
1-
12
#892920000000
0!
0%
b110 *
0-
02
b110 6
#892930000000
1!
1%
1-
12
#892940000000
0!
0%
b111 *
0-
02
b111 6
#892950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#892960000000
0!
0%
b0 *
0-
02
b0 6
#892970000000
1!
1%
1-
12
#892980000000
0!
0%
b1 *
0-
02
b1 6
#892990000000
1!
1%
1-
12
#893000000000
0!
0%
b10 *
0-
02
b10 6
#893010000000
1!
1%
1-
12
#893020000000
0!
0%
b11 *
0-
02
b11 6
#893030000000
1!
1%
1-
12
15
#893040000000
0!
0%
b100 *
0-
02
b100 6
#893050000000
1!
1%
1-
12
#893060000000
0!
0%
b101 *
0-
02
b101 6
#893070000000
1!
1%
1-
12
#893080000000
0!
0%
b110 *
0-
02
b110 6
#893090000000
1!
1%
1-
12
#893100000000
0!
0%
b111 *
0-
02
b111 6
#893110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#893120000000
0!
0%
b0 *
0-
02
b0 6
#893130000000
1!
1%
1-
12
#893140000000
0!
0%
b1 *
0-
02
b1 6
#893150000000
1!
1%
1-
12
#893160000000
0!
0%
b10 *
0-
02
b10 6
#893170000000
1!
1%
1-
12
#893180000000
0!
0%
b11 *
0-
02
b11 6
#893190000000
1!
1%
1-
12
15
#893200000000
0!
0%
b100 *
0-
02
b100 6
#893210000000
1!
1%
1-
12
#893220000000
0!
0%
b101 *
0-
02
b101 6
#893230000000
1!
1%
1-
12
#893240000000
0!
0%
b110 *
0-
02
b110 6
#893250000000
1!
1%
1-
12
#893260000000
0!
0%
b111 *
0-
02
b111 6
#893270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#893280000000
0!
0%
b0 *
0-
02
b0 6
#893290000000
1!
1%
1-
12
#893300000000
0!
0%
b1 *
0-
02
b1 6
#893310000000
1!
1%
1-
12
#893320000000
0!
0%
b10 *
0-
02
b10 6
#893330000000
1!
1%
1-
12
#893340000000
0!
0%
b11 *
0-
02
b11 6
#893350000000
1!
1%
1-
12
15
#893360000000
0!
0%
b100 *
0-
02
b100 6
#893370000000
1!
1%
1-
12
#893380000000
0!
0%
b101 *
0-
02
b101 6
#893390000000
1!
1%
1-
12
#893400000000
0!
0%
b110 *
0-
02
b110 6
#893410000000
1!
1%
1-
12
#893420000000
0!
0%
b111 *
0-
02
b111 6
#893430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#893440000000
0!
0%
b0 *
0-
02
b0 6
#893450000000
1!
1%
1-
12
#893460000000
0!
0%
b1 *
0-
02
b1 6
#893470000000
1!
1%
1-
12
#893480000000
0!
0%
b10 *
0-
02
b10 6
#893490000000
1!
1%
1-
12
#893500000000
0!
0%
b11 *
0-
02
b11 6
#893510000000
1!
1%
1-
12
15
#893520000000
0!
0%
b100 *
0-
02
b100 6
#893530000000
1!
1%
1-
12
#893540000000
0!
0%
b101 *
0-
02
b101 6
#893550000000
1!
1%
1-
12
#893560000000
0!
0%
b110 *
0-
02
b110 6
#893570000000
1!
1%
1-
12
#893580000000
0!
0%
b111 *
0-
02
b111 6
#893590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#893600000000
0!
0%
b0 *
0-
02
b0 6
#893610000000
1!
1%
1-
12
#893620000000
0!
0%
b1 *
0-
02
b1 6
#893630000000
1!
1%
1-
12
#893640000000
0!
0%
b10 *
0-
02
b10 6
#893650000000
1!
1%
1-
12
#893660000000
0!
0%
b11 *
0-
02
b11 6
#893670000000
1!
1%
1-
12
15
#893680000000
0!
0%
b100 *
0-
02
b100 6
#893690000000
1!
1%
1-
12
#893700000000
0!
0%
b101 *
0-
02
b101 6
#893710000000
1!
1%
1-
12
#893720000000
0!
0%
b110 *
0-
02
b110 6
#893730000000
1!
1%
1-
12
#893740000000
0!
0%
b111 *
0-
02
b111 6
#893750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#893760000000
0!
0%
b0 *
0-
02
b0 6
#893770000000
1!
1%
1-
12
#893780000000
0!
0%
b1 *
0-
02
b1 6
#893790000000
1!
1%
1-
12
#893800000000
0!
0%
b10 *
0-
02
b10 6
#893810000000
1!
1%
1-
12
#893820000000
0!
0%
b11 *
0-
02
b11 6
#893830000000
1!
1%
1-
12
15
#893840000000
0!
0%
b100 *
0-
02
b100 6
#893850000000
1!
1%
1-
12
#893860000000
0!
0%
b101 *
0-
02
b101 6
#893870000000
1!
1%
1-
12
#893880000000
0!
0%
b110 *
0-
02
b110 6
#893890000000
1!
1%
1-
12
#893900000000
0!
0%
b111 *
0-
02
b111 6
#893910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#893920000000
0!
0%
b0 *
0-
02
b0 6
#893930000000
1!
1%
1-
12
#893940000000
0!
0%
b1 *
0-
02
b1 6
#893950000000
1!
1%
1-
12
#893960000000
0!
0%
b10 *
0-
02
b10 6
#893970000000
1!
1%
1-
12
#893980000000
0!
0%
b11 *
0-
02
b11 6
#893990000000
1!
1%
1-
12
15
#894000000000
0!
0%
b100 *
0-
02
b100 6
#894010000000
1!
1%
1-
12
#894020000000
0!
0%
b101 *
0-
02
b101 6
#894030000000
1!
1%
1-
12
#894040000000
0!
0%
b110 *
0-
02
b110 6
#894050000000
1!
1%
1-
12
#894060000000
0!
0%
b111 *
0-
02
b111 6
#894070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#894080000000
0!
0%
b0 *
0-
02
b0 6
#894090000000
1!
1%
1-
12
#894100000000
0!
0%
b1 *
0-
02
b1 6
#894110000000
1!
1%
1-
12
#894120000000
0!
0%
b10 *
0-
02
b10 6
#894130000000
1!
1%
1-
12
#894140000000
0!
0%
b11 *
0-
02
b11 6
#894150000000
1!
1%
1-
12
15
#894160000000
0!
0%
b100 *
0-
02
b100 6
#894170000000
1!
1%
1-
12
#894180000000
0!
0%
b101 *
0-
02
b101 6
#894190000000
1!
1%
1-
12
#894200000000
0!
0%
b110 *
0-
02
b110 6
#894210000000
1!
1%
1-
12
#894220000000
0!
0%
b111 *
0-
02
b111 6
#894230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#894240000000
0!
0%
b0 *
0-
02
b0 6
#894250000000
1!
1%
1-
12
#894260000000
0!
0%
b1 *
0-
02
b1 6
#894270000000
1!
1%
1-
12
#894280000000
0!
0%
b10 *
0-
02
b10 6
#894290000000
1!
1%
1-
12
#894300000000
0!
0%
b11 *
0-
02
b11 6
#894310000000
1!
1%
1-
12
15
#894320000000
0!
0%
b100 *
0-
02
b100 6
#894330000000
1!
1%
1-
12
#894340000000
0!
0%
b101 *
0-
02
b101 6
#894350000000
1!
1%
1-
12
#894360000000
0!
0%
b110 *
0-
02
b110 6
#894370000000
1!
1%
1-
12
#894380000000
0!
0%
b111 *
0-
02
b111 6
#894390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#894400000000
0!
0%
b0 *
0-
02
b0 6
#894410000000
1!
1%
1-
12
#894420000000
0!
0%
b1 *
0-
02
b1 6
#894430000000
1!
1%
1-
12
#894440000000
0!
0%
b10 *
0-
02
b10 6
#894450000000
1!
1%
1-
12
#894460000000
0!
0%
b11 *
0-
02
b11 6
#894470000000
1!
1%
1-
12
15
#894480000000
0!
0%
b100 *
0-
02
b100 6
#894490000000
1!
1%
1-
12
#894500000000
0!
0%
b101 *
0-
02
b101 6
#894510000000
1!
1%
1-
12
#894520000000
0!
0%
b110 *
0-
02
b110 6
#894530000000
1!
1%
1-
12
#894540000000
0!
0%
b111 *
0-
02
b111 6
#894550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#894560000000
0!
0%
b0 *
0-
02
b0 6
#894570000000
1!
1%
1-
12
#894580000000
0!
0%
b1 *
0-
02
b1 6
#894590000000
1!
1%
1-
12
#894600000000
0!
0%
b10 *
0-
02
b10 6
#894610000000
1!
1%
1-
12
#894620000000
0!
0%
b11 *
0-
02
b11 6
#894630000000
1!
1%
1-
12
15
#894640000000
0!
0%
b100 *
0-
02
b100 6
#894650000000
1!
1%
1-
12
#894660000000
0!
0%
b101 *
0-
02
b101 6
#894670000000
1!
1%
1-
12
#894680000000
0!
0%
b110 *
0-
02
b110 6
#894690000000
1!
1%
1-
12
#894700000000
0!
0%
b111 *
0-
02
b111 6
#894710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#894720000000
0!
0%
b0 *
0-
02
b0 6
#894730000000
1!
1%
1-
12
#894740000000
0!
0%
b1 *
0-
02
b1 6
#894750000000
1!
1%
1-
12
#894760000000
0!
0%
b10 *
0-
02
b10 6
#894770000000
1!
1%
1-
12
#894780000000
0!
0%
b11 *
0-
02
b11 6
#894790000000
1!
1%
1-
12
15
#894800000000
0!
0%
b100 *
0-
02
b100 6
#894810000000
1!
1%
1-
12
#894820000000
0!
0%
b101 *
0-
02
b101 6
#894830000000
1!
1%
1-
12
#894840000000
0!
0%
b110 *
0-
02
b110 6
#894850000000
1!
1%
1-
12
#894860000000
0!
0%
b111 *
0-
02
b111 6
#894870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#894880000000
0!
0%
b0 *
0-
02
b0 6
#894890000000
1!
1%
1-
12
#894900000000
0!
0%
b1 *
0-
02
b1 6
#894910000000
1!
1%
1-
12
#894920000000
0!
0%
b10 *
0-
02
b10 6
#894930000000
1!
1%
1-
12
#894940000000
0!
0%
b11 *
0-
02
b11 6
#894950000000
1!
1%
1-
12
15
#894960000000
0!
0%
b100 *
0-
02
b100 6
#894970000000
1!
1%
1-
12
#894980000000
0!
0%
b101 *
0-
02
b101 6
#894990000000
1!
1%
1-
12
#895000000000
0!
0%
b110 *
0-
02
b110 6
#895010000000
1!
1%
1-
12
#895020000000
0!
0%
b111 *
0-
02
b111 6
#895030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#895040000000
0!
0%
b0 *
0-
02
b0 6
#895050000000
1!
1%
1-
12
#895060000000
0!
0%
b1 *
0-
02
b1 6
#895070000000
1!
1%
1-
12
#895080000000
0!
0%
b10 *
0-
02
b10 6
#895090000000
1!
1%
1-
12
#895100000000
0!
0%
b11 *
0-
02
b11 6
#895110000000
1!
1%
1-
12
15
#895120000000
0!
0%
b100 *
0-
02
b100 6
#895130000000
1!
1%
1-
12
#895140000000
0!
0%
b101 *
0-
02
b101 6
#895150000000
1!
1%
1-
12
#895160000000
0!
0%
b110 *
0-
02
b110 6
#895170000000
1!
1%
1-
12
#895180000000
0!
0%
b111 *
0-
02
b111 6
#895190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#895200000000
0!
0%
b0 *
0-
02
b0 6
#895210000000
1!
1%
1-
12
#895220000000
0!
0%
b1 *
0-
02
b1 6
#895230000000
1!
1%
1-
12
#895240000000
0!
0%
b10 *
0-
02
b10 6
#895250000000
1!
1%
1-
12
#895260000000
0!
0%
b11 *
0-
02
b11 6
#895270000000
1!
1%
1-
12
15
#895280000000
0!
0%
b100 *
0-
02
b100 6
#895290000000
1!
1%
1-
12
#895300000000
0!
0%
b101 *
0-
02
b101 6
#895310000000
1!
1%
1-
12
#895320000000
0!
0%
b110 *
0-
02
b110 6
#895330000000
1!
1%
1-
12
#895340000000
0!
0%
b111 *
0-
02
b111 6
#895350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#895360000000
0!
0%
b0 *
0-
02
b0 6
#895370000000
1!
1%
1-
12
#895380000000
0!
0%
b1 *
0-
02
b1 6
#895390000000
1!
1%
1-
12
#895400000000
0!
0%
b10 *
0-
02
b10 6
#895410000000
1!
1%
1-
12
#895420000000
0!
0%
b11 *
0-
02
b11 6
#895430000000
1!
1%
1-
12
15
#895440000000
0!
0%
b100 *
0-
02
b100 6
#895450000000
1!
1%
1-
12
#895460000000
0!
0%
b101 *
0-
02
b101 6
#895470000000
1!
1%
1-
12
#895480000000
0!
0%
b110 *
0-
02
b110 6
#895490000000
1!
1%
1-
12
#895500000000
0!
0%
b111 *
0-
02
b111 6
#895510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#895520000000
0!
0%
b0 *
0-
02
b0 6
#895530000000
1!
1%
1-
12
#895540000000
0!
0%
b1 *
0-
02
b1 6
#895550000000
1!
1%
1-
12
#895560000000
0!
0%
b10 *
0-
02
b10 6
#895570000000
1!
1%
1-
12
#895580000000
0!
0%
b11 *
0-
02
b11 6
#895590000000
1!
1%
1-
12
15
#895600000000
0!
0%
b100 *
0-
02
b100 6
#895610000000
1!
1%
1-
12
#895620000000
0!
0%
b101 *
0-
02
b101 6
#895630000000
1!
1%
1-
12
#895640000000
0!
0%
b110 *
0-
02
b110 6
#895650000000
1!
1%
1-
12
#895660000000
0!
0%
b111 *
0-
02
b111 6
#895670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#895680000000
0!
0%
b0 *
0-
02
b0 6
#895690000000
1!
1%
1-
12
#895700000000
0!
0%
b1 *
0-
02
b1 6
#895710000000
1!
1%
1-
12
#895720000000
0!
0%
b10 *
0-
02
b10 6
#895730000000
1!
1%
1-
12
#895740000000
0!
0%
b11 *
0-
02
b11 6
#895750000000
1!
1%
1-
12
15
#895760000000
0!
0%
b100 *
0-
02
b100 6
#895770000000
1!
1%
1-
12
#895780000000
0!
0%
b101 *
0-
02
b101 6
#895790000000
1!
1%
1-
12
#895800000000
0!
0%
b110 *
0-
02
b110 6
#895810000000
1!
1%
1-
12
#895820000000
0!
0%
b111 *
0-
02
b111 6
#895830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#895840000000
0!
0%
b0 *
0-
02
b0 6
#895850000000
1!
1%
1-
12
#895860000000
0!
0%
b1 *
0-
02
b1 6
#895870000000
1!
1%
1-
12
#895880000000
0!
0%
b10 *
0-
02
b10 6
#895890000000
1!
1%
1-
12
#895900000000
0!
0%
b11 *
0-
02
b11 6
#895910000000
1!
1%
1-
12
15
#895920000000
0!
0%
b100 *
0-
02
b100 6
#895930000000
1!
1%
1-
12
#895940000000
0!
0%
b101 *
0-
02
b101 6
#895950000000
1!
1%
1-
12
#895960000000
0!
0%
b110 *
0-
02
b110 6
#895970000000
1!
1%
1-
12
#895980000000
0!
0%
b111 *
0-
02
b111 6
#895990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#896000000000
0!
0%
b0 *
0-
02
b0 6
#896010000000
1!
1%
1-
12
#896020000000
0!
0%
b1 *
0-
02
b1 6
#896030000000
1!
1%
1-
12
#896040000000
0!
0%
b10 *
0-
02
b10 6
#896050000000
1!
1%
1-
12
#896060000000
0!
0%
b11 *
0-
02
b11 6
#896070000000
1!
1%
1-
12
15
#896080000000
0!
0%
b100 *
0-
02
b100 6
#896090000000
1!
1%
1-
12
#896100000000
0!
0%
b101 *
0-
02
b101 6
#896110000000
1!
1%
1-
12
#896120000000
0!
0%
b110 *
0-
02
b110 6
#896130000000
1!
1%
1-
12
#896140000000
0!
0%
b111 *
0-
02
b111 6
#896150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#896160000000
0!
0%
b0 *
0-
02
b0 6
#896170000000
1!
1%
1-
12
#896180000000
0!
0%
b1 *
0-
02
b1 6
#896190000000
1!
1%
1-
12
#896200000000
0!
0%
b10 *
0-
02
b10 6
#896210000000
1!
1%
1-
12
#896220000000
0!
0%
b11 *
0-
02
b11 6
#896230000000
1!
1%
1-
12
15
#896240000000
0!
0%
b100 *
0-
02
b100 6
#896250000000
1!
1%
1-
12
#896260000000
0!
0%
b101 *
0-
02
b101 6
#896270000000
1!
1%
1-
12
#896280000000
0!
0%
b110 *
0-
02
b110 6
#896290000000
1!
1%
1-
12
#896300000000
0!
0%
b111 *
0-
02
b111 6
#896310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#896320000000
0!
0%
b0 *
0-
02
b0 6
#896330000000
1!
1%
1-
12
#896340000000
0!
0%
b1 *
0-
02
b1 6
#896350000000
1!
1%
1-
12
#896360000000
0!
0%
b10 *
0-
02
b10 6
#896370000000
1!
1%
1-
12
#896380000000
0!
0%
b11 *
0-
02
b11 6
#896390000000
1!
1%
1-
12
15
#896400000000
0!
0%
b100 *
0-
02
b100 6
#896410000000
1!
1%
1-
12
#896420000000
0!
0%
b101 *
0-
02
b101 6
#896430000000
1!
1%
1-
12
#896440000000
0!
0%
b110 *
0-
02
b110 6
#896450000000
1!
1%
1-
12
#896460000000
0!
0%
b111 *
0-
02
b111 6
#896470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#896480000000
0!
0%
b0 *
0-
02
b0 6
#896490000000
1!
1%
1-
12
#896500000000
0!
0%
b1 *
0-
02
b1 6
#896510000000
1!
1%
1-
12
#896520000000
0!
0%
b10 *
0-
02
b10 6
#896530000000
1!
1%
1-
12
#896540000000
0!
0%
b11 *
0-
02
b11 6
#896550000000
1!
1%
1-
12
15
#896560000000
0!
0%
b100 *
0-
02
b100 6
#896570000000
1!
1%
1-
12
#896580000000
0!
0%
b101 *
0-
02
b101 6
#896590000000
1!
1%
1-
12
#896600000000
0!
0%
b110 *
0-
02
b110 6
#896610000000
1!
1%
1-
12
#896620000000
0!
0%
b111 *
0-
02
b111 6
#896630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#896640000000
0!
0%
b0 *
0-
02
b0 6
#896650000000
1!
1%
1-
12
#896660000000
0!
0%
b1 *
0-
02
b1 6
#896670000000
1!
1%
1-
12
#896680000000
0!
0%
b10 *
0-
02
b10 6
#896690000000
1!
1%
1-
12
#896700000000
0!
0%
b11 *
0-
02
b11 6
#896710000000
1!
1%
1-
12
15
#896720000000
0!
0%
b100 *
0-
02
b100 6
#896730000000
1!
1%
1-
12
#896740000000
0!
0%
b101 *
0-
02
b101 6
#896750000000
1!
1%
1-
12
#896760000000
0!
0%
b110 *
0-
02
b110 6
#896770000000
1!
1%
1-
12
#896780000000
0!
0%
b111 *
0-
02
b111 6
#896790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#896800000000
0!
0%
b0 *
0-
02
b0 6
#896810000000
1!
1%
1-
12
#896820000000
0!
0%
b1 *
0-
02
b1 6
#896830000000
1!
1%
1-
12
#896840000000
0!
0%
b10 *
0-
02
b10 6
#896850000000
1!
1%
1-
12
#896860000000
0!
0%
b11 *
0-
02
b11 6
#896870000000
1!
1%
1-
12
15
#896880000000
0!
0%
b100 *
0-
02
b100 6
#896890000000
1!
1%
1-
12
#896900000000
0!
0%
b101 *
0-
02
b101 6
#896910000000
1!
1%
1-
12
#896920000000
0!
0%
b110 *
0-
02
b110 6
#896930000000
1!
1%
1-
12
#896940000000
0!
0%
b111 *
0-
02
b111 6
#896950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#896960000000
0!
0%
b0 *
0-
02
b0 6
#896970000000
1!
1%
1-
12
#896980000000
0!
0%
b1 *
0-
02
b1 6
#896990000000
1!
1%
1-
12
#897000000000
0!
0%
b10 *
0-
02
b10 6
#897010000000
1!
1%
1-
12
#897020000000
0!
0%
b11 *
0-
02
b11 6
#897030000000
1!
1%
1-
12
15
#897040000000
0!
0%
b100 *
0-
02
b100 6
#897050000000
1!
1%
1-
12
#897060000000
0!
0%
b101 *
0-
02
b101 6
#897070000000
1!
1%
1-
12
#897080000000
0!
0%
b110 *
0-
02
b110 6
#897090000000
1!
1%
1-
12
#897100000000
0!
0%
b111 *
0-
02
b111 6
#897110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#897120000000
0!
0%
b0 *
0-
02
b0 6
#897130000000
1!
1%
1-
12
#897140000000
0!
0%
b1 *
0-
02
b1 6
#897150000000
1!
1%
1-
12
#897160000000
0!
0%
b10 *
0-
02
b10 6
#897170000000
1!
1%
1-
12
#897180000000
0!
0%
b11 *
0-
02
b11 6
#897190000000
1!
1%
1-
12
15
#897200000000
0!
0%
b100 *
0-
02
b100 6
#897210000000
1!
1%
1-
12
#897220000000
0!
0%
b101 *
0-
02
b101 6
#897230000000
1!
1%
1-
12
#897240000000
0!
0%
b110 *
0-
02
b110 6
#897250000000
1!
1%
1-
12
#897260000000
0!
0%
b111 *
0-
02
b111 6
#897270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#897280000000
0!
0%
b0 *
0-
02
b0 6
#897290000000
1!
1%
1-
12
#897300000000
0!
0%
b1 *
0-
02
b1 6
#897310000000
1!
1%
1-
12
#897320000000
0!
0%
b10 *
0-
02
b10 6
#897330000000
1!
1%
1-
12
#897340000000
0!
0%
b11 *
0-
02
b11 6
#897350000000
1!
1%
1-
12
15
#897360000000
0!
0%
b100 *
0-
02
b100 6
#897370000000
1!
1%
1-
12
#897380000000
0!
0%
b101 *
0-
02
b101 6
#897390000000
1!
1%
1-
12
#897400000000
0!
0%
b110 *
0-
02
b110 6
#897410000000
1!
1%
1-
12
#897420000000
0!
0%
b111 *
0-
02
b111 6
#897430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#897440000000
0!
0%
b0 *
0-
02
b0 6
#897450000000
1!
1%
1-
12
#897460000000
0!
0%
b1 *
0-
02
b1 6
#897470000000
1!
1%
1-
12
#897480000000
0!
0%
b10 *
0-
02
b10 6
#897490000000
1!
1%
1-
12
#897500000000
0!
0%
b11 *
0-
02
b11 6
#897510000000
1!
1%
1-
12
15
#897520000000
0!
0%
b100 *
0-
02
b100 6
#897530000000
1!
1%
1-
12
#897540000000
0!
0%
b101 *
0-
02
b101 6
#897550000000
1!
1%
1-
12
#897560000000
0!
0%
b110 *
0-
02
b110 6
#897570000000
1!
1%
1-
12
#897580000000
0!
0%
b111 *
0-
02
b111 6
#897590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#897600000000
0!
0%
b0 *
0-
02
b0 6
#897610000000
1!
1%
1-
12
#897620000000
0!
0%
b1 *
0-
02
b1 6
#897630000000
1!
1%
1-
12
#897640000000
0!
0%
b10 *
0-
02
b10 6
#897650000000
1!
1%
1-
12
#897660000000
0!
0%
b11 *
0-
02
b11 6
#897670000000
1!
1%
1-
12
15
#897680000000
0!
0%
b100 *
0-
02
b100 6
#897690000000
1!
1%
1-
12
#897700000000
0!
0%
b101 *
0-
02
b101 6
#897710000000
1!
1%
1-
12
#897720000000
0!
0%
b110 *
0-
02
b110 6
#897730000000
1!
1%
1-
12
#897740000000
0!
0%
b111 *
0-
02
b111 6
#897750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#897760000000
0!
0%
b0 *
0-
02
b0 6
#897770000000
1!
1%
1-
12
#897780000000
0!
0%
b1 *
0-
02
b1 6
#897790000000
1!
1%
1-
12
#897800000000
0!
0%
b10 *
0-
02
b10 6
#897810000000
1!
1%
1-
12
#897820000000
0!
0%
b11 *
0-
02
b11 6
#897830000000
1!
1%
1-
12
15
#897840000000
0!
0%
b100 *
0-
02
b100 6
#897850000000
1!
1%
1-
12
#897860000000
0!
0%
b101 *
0-
02
b101 6
#897870000000
1!
1%
1-
12
#897880000000
0!
0%
b110 *
0-
02
b110 6
#897890000000
1!
1%
1-
12
#897900000000
0!
0%
b111 *
0-
02
b111 6
#897910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#897920000000
0!
0%
b0 *
0-
02
b0 6
#897930000000
1!
1%
1-
12
#897940000000
0!
0%
b1 *
0-
02
b1 6
#897950000000
1!
1%
1-
12
#897960000000
0!
0%
b10 *
0-
02
b10 6
#897970000000
1!
1%
1-
12
#897980000000
0!
0%
b11 *
0-
02
b11 6
#897990000000
1!
1%
1-
12
15
#898000000000
0!
0%
b100 *
0-
02
b100 6
#898010000000
1!
1%
1-
12
#898020000000
0!
0%
b101 *
0-
02
b101 6
#898030000000
1!
1%
1-
12
#898040000000
0!
0%
b110 *
0-
02
b110 6
#898050000000
1!
1%
1-
12
#898060000000
0!
0%
b111 *
0-
02
b111 6
#898070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#898080000000
0!
0%
b0 *
0-
02
b0 6
#898090000000
1!
1%
1-
12
#898100000000
0!
0%
b1 *
0-
02
b1 6
#898110000000
1!
1%
1-
12
#898120000000
0!
0%
b10 *
0-
02
b10 6
#898130000000
1!
1%
1-
12
#898140000000
0!
0%
b11 *
0-
02
b11 6
#898150000000
1!
1%
1-
12
15
#898160000000
0!
0%
b100 *
0-
02
b100 6
#898170000000
1!
1%
1-
12
#898180000000
0!
0%
b101 *
0-
02
b101 6
#898190000000
1!
1%
1-
12
#898200000000
0!
0%
b110 *
0-
02
b110 6
#898210000000
1!
1%
1-
12
#898220000000
0!
0%
b111 *
0-
02
b111 6
#898230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#898240000000
0!
0%
b0 *
0-
02
b0 6
#898250000000
1!
1%
1-
12
#898260000000
0!
0%
b1 *
0-
02
b1 6
#898270000000
1!
1%
1-
12
#898280000000
0!
0%
b10 *
0-
02
b10 6
#898290000000
1!
1%
1-
12
#898300000000
0!
0%
b11 *
0-
02
b11 6
#898310000000
1!
1%
1-
12
15
#898320000000
0!
0%
b100 *
0-
02
b100 6
#898330000000
1!
1%
1-
12
#898340000000
0!
0%
b101 *
0-
02
b101 6
#898350000000
1!
1%
1-
12
#898360000000
0!
0%
b110 *
0-
02
b110 6
#898370000000
1!
1%
1-
12
#898380000000
0!
0%
b111 *
0-
02
b111 6
#898390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#898400000000
0!
0%
b0 *
0-
02
b0 6
#898410000000
1!
1%
1-
12
#898420000000
0!
0%
b1 *
0-
02
b1 6
#898430000000
1!
1%
1-
12
#898440000000
0!
0%
b10 *
0-
02
b10 6
#898450000000
1!
1%
1-
12
#898460000000
0!
0%
b11 *
0-
02
b11 6
#898470000000
1!
1%
1-
12
15
#898480000000
0!
0%
b100 *
0-
02
b100 6
#898490000000
1!
1%
1-
12
#898500000000
0!
0%
b101 *
0-
02
b101 6
#898510000000
1!
1%
1-
12
#898520000000
0!
0%
b110 *
0-
02
b110 6
#898530000000
1!
1%
1-
12
#898540000000
0!
0%
b111 *
0-
02
b111 6
#898550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#898560000000
0!
0%
b0 *
0-
02
b0 6
#898570000000
1!
1%
1-
12
#898580000000
0!
0%
b1 *
0-
02
b1 6
#898590000000
1!
1%
1-
12
#898600000000
0!
0%
b10 *
0-
02
b10 6
#898610000000
1!
1%
1-
12
#898620000000
0!
0%
b11 *
0-
02
b11 6
#898630000000
1!
1%
1-
12
15
#898640000000
0!
0%
b100 *
0-
02
b100 6
#898650000000
1!
1%
1-
12
#898660000000
0!
0%
b101 *
0-
02
b101 6
#898670000000
1!
1%
1-
12
#898680000000
0!
0%
b110 *
0-
02
b110 6
#898690000000
1!
1%
1-
12
#898700000000
0!
0%
b111 *
0-
02
b111 6
#898710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#898720000000
0!
0%
b0 *
0-
02
b0 6
#898730000000
1!
1%
1-
12
#898740000000
0!
0%
b1 *
0-
02
b1 6
#898750000000
1!
1%
1-
12
#898760000000
0!
0%
b10 *
0-
02
b10 6
#898770000000
1!
1%
1-
12
#898780000000
0!
0%
b11 *
0-
02
b11 6
#898790000000
1!
1%
1-
12
15
#898800000000
0!
0%
b100 *
0-
02
b100 6
#898810000000
1!
1%
1-
12
#898820000000
0!
0%
b101 *
0-
02
b101 6
#898830000000
1!
1%
1-
12
#898840000000
0!
0%
b110 *
0-
02
b110 6
#898850000000
1!
1%
1-
12
#898860000000
0!
0%
b111 *
0-
02
b111 6
#898870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#898880000000
0!
0%
b0 *
0-
02
b0 6
#898890000000
1!
1%
1-
12
#898900000000
0!
0%
b1 *
0-
02
b1 6
#898910000000
1!
1%
1-
12
#898920000000
0!
0%
b10 *
0-
02
b10 6
#898930000000
1!
1%
1-
12
#898940000000
0!
0%
b11 *
0-
02
b11 6
#898950000000
1!
1%
1-
12
15
#898960000000
0!
0%
b100 *
0-
02
b100 6
#898970000000
1!
1%
1-
12
#898980000000
0!
0%
b101 *
0-
02
b101 6
#898990000000
1!
1%
1-
12
#899000000000
0!
0%
b110 *
0-
02
b110 6
#899010000000
1!
1%
1-
12
#899020000000
0!
0%
b111 *
0-
02
b111 6
#899030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#899040000000
0!
0%
b0 *
0-
02
b0 6
#899050000000
1!
1%
1-
12
#899060000000
0!
0%
b1 *
0-
02
b1 6
#899070000000
1!
1%
1-
12
#899080000000
0!
0%
b10 *
0-
02
b10 6
#899090000000
1!
1%
1-
12
#899100000000
0!
0%
b11 *
0-
02
b11 6
#899110000000
1!
1%
1-
12
15
#899120000000
0!
0%
b100 *
0-
02
b100 6
#899130000000
1!
1%
1-
12
#899140000000
0!
0%
b101 *
0-
02
b101 6
#899150000000
1!
1%
1-
12
#899160000000
0!
0%
b110 *
0-
02
b110 6
#899170000000
1!
1%
1-
12
#899180000000
0!
0%
b111 *
0-
02
b111 6
#899190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#899200000000
0!
0%
b0 *
0-
02
b0 6
#899210000000
1!
1%
1-
12
#899220000000
0!
0%
b1 *
0-
02
b1 6
#899230000000
1!
1%
1-
12
#899240000000
0!
0%
b10 *
0-
02
b10 6
#899250000000
1!
1%
1-
12
#899260000000
0!
0%
b11 *
0-
02
b11 6
#899270000000
1!
1%
1-
12
15
#899280000000
0!
0%
b100 *
0-
02
b100 6
#899290000000
1!
1%
1-
12
#899300000000
0!
0%
b101 *
0-
02
b101 6
#899310000000
1!
1%
1-
12
#899320000000
0!
0%
b110 *
0-
02
b110 6
#899330000000
1!
1%
1-
12
#899340000000
0!
0%
b111 *
0-
02
b111 6
#899350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#899360000000
0!
0%
b0 *
0-
02
b0 6
#899370000000
1!
1%
1-
12
#899380000000
0!
0%
b1 *
0-
02
b1 6
#899390000000
1!
1%
1-
12
#899400000000
0!
0%
b10 *
0-
02
b10 6
#899410000000
1!
1%
1-
12
#899420000000
0!
0%
b11 *
0-
02
b11 6
#899430000000
1!
1%
1-
12
15
#899440000000
0!
0%
b100 *
0-
02
b100 6
#899450000000
1!
1%
1-
12
#899460000000
0!
0%
b101 *
0-
02
b101 6
#899470000000
1!
1%
1-
12
#899480000000
0!
0%
b110 *
0-
02
b110 6
#899490000000
1!
1%
1-
12
#899500000000
0!
0%
b111 *
0-
02
b111 6
#899510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#899520000000
0!
0%
b0 *
0-
02
b0 6
#899530000000
1!
1%
1-
12
#899540000000
0!
0%
b1 *
0-
02
b1 6
#899550000000
1!
1%
1-
12
#899560000000
0!
0%
b10 *
0-
02
b10 6
#899570000000
1!
1%
1-
12
#899580000000
0!
0%
b11 *
0-
02
b11 6
#899590000000
1!
1%
1-
12
15
#899600000000
0!
0%
b100 *
0-
02
b100 6
#899610000000
1!
1%
1-
12
#899620000000
0!
0%
b101 *
0-
02
b101 6
#899630000000
1!
1%
1-
12
#899640000000
0!
0%
b110 *
0-
02
b110 6
#899650000000
1!
1%
1-
12
#899660000000
0!
0%
b111 *
0-
02
b111 6
#899670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#899680000000
0!
0%
b0 *
0-
02
b0 6
#899690000000
1!
1%
1-
12
#899700000000
0!
0%
b1 *
0-
02
b1 6
#899710000000
1!
1%
1-
12
#899720000000
0!
0%
b10 *
0-
02
b10 6
#899730000000
1!
1%
1-
12
#899740000000
0!
0%
b11 *
0-
02
b11 6
#899750000000
1!
1%
1-
12
15
#899760000000
0!
0%
b100 *
0-
02
b100 6
#899770000000
1!
1%
1-
12
#899780000000
0!
0%
b101 *
0-
02
b101 6
#899790000000
1!
1%
1-
12
#899800000000
0!
0%
b110 *
0-
02
b110 6
#899810000000
1!
1%
1-
12
#899820000000
0!
0%
b111 *
0-
02
b111 6
#899830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#899840000000
0!
0%
b0 *
0-
02
b0 6
#899850000000
1!
1%
1-
12
#899860000000
0!
0%
b1 *
0-
02
b1 6
#899870000000
1!
1%
1-
12
#899880000000
0!
0%
b10 *
0-
02
b10 6
#899890000000
1!
1%
1-
12
#899900000000
0!
0%
b11 *
0-
02
b11 6
#899910000000
1!
1%
1-
12
15
#899920000000
0!
0%
b100 *
0-
02
b100 6
#899930000000
1!
1%
1-
12
#899940000000
0!
0%
b101 *
0-
02
b101 6
#899950000000
1!
1%
1-
12
#899960000000
0!
0%
b110 *
0-
02
b110 6
#899970000000
1!
1%
1-
12
#899980000000
0!
0%
b111 *
0-
02
b111 6
#899990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#900000000000
0!
0%
b0 *
0-
02
b0 6
#900010000000
1!
1%
1-
12
#900020000000
0!
0%
b1 *
0-
02
b1 6
#900030000000
1!
1%
1-
12
#900040000000
0!
0%
b10 *
0-
02
b10 6
#900050000000
1!
1%
1-
12
#900060000000
0!
0%
b11 *
0-
02
b11 6
#900070000000
1!
1%
1-
12
15
#900080000000
0!
0%
b100 *
0-
02
b100 6
#900090000000
1!
1%
1-
12
#900100000000
0!
0%
b101 *
0-
02
b101 6
#900110000000
1!
1%
1-
12
#900120000000
0!
0%
b110 *
0-
02
b110 6
#900130000000
1!
1%
1-
12
#900140000000
0!
0%
b111 *
0-
02
b111 6
#900150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#900160000000
0!
0%
b0 *
0-
02
b0 6
#900170000000
1!
1%
1-
12
#900180000000
0!
0%
b1 *
0-
02
b1 6
#900190000000
1!
1%
1-
12
#900200000000
0!
0%
b10 *
0-
02
b10 6
#900210000000
1!
1%
1-
12
#900220000000
0!
0%
b11 *
0-
02
b11 6
#900230000000
1!
1%
1-
12
15
#900240000000
0!
0%
b100 *
0-
02
b100 6
#900250000000
1!
1%
1-
12
#900260000000
0!
0%
b101 *
0-
02
b101 6
#900270000000
1!
1%
1-
12
#900280000000
0!
0%
b110 *
0-
02
b110 6
#900290000000
1!
1%
1-
12
#900300000000
0!
0%
b111 *
0-
02
b111 6
#900310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#900320000000
0!
0%
b0 *
0-
02
b0 6
#900330000000
1!
1%
1-
12
#900340000000
0!
0%
b1 *
0-
02
b1 6
#900350000000
1!
1%
1-
12
#900360000000
0!
0%
b10 *
0-
02
b10 6
#900370000000
1!
1%
1-
12
#900380000000
0!
0%
b11 *
0-
02
b11 6
#900390000000
1!
1%
1-
12
15
#900400000000
0!
0%
b100 *
0-
02
b100 6
#900410000000
1!
1%
1-
12
#900420000000
0!
0%
b101 *
0-
02
b101 6
#900430000000
1!
1%
1-
12
#900440000000
0!
0%
b110 *
0-
02
b110 6
#900450000000
1!
1%
1-
12
#900460000000
0!
0%
b111 *
0-
02
b111 6
#900470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#900480000000
0!
0%
b0 *
0-
02
b0 6
#900490000000
1!
1%
1-
12
#900500000000
0!
0%
b1 *
0-
02
b1 6
#900510000000
1!
1%
1-
12
#900520000000
0!
0%
b10 *
0-
02
b10 6
#900530000000
1!
1%
1-
12
#900540000000
0!
0%
b11 *
0-
02
b11 6
#900550000000
1!
1%
1-
12
15
#900560000000
0!
0%
b100 *
0-
02
b100 6
#900570000000
1!
1%
1-
12
#900580000000
0!
0%
b101 *
0-
02
b101 6
#900590000000
1!
1%
1-
12
#900600000000
0!
0%
b110 *
0-
02
b110 6
#900610000000
1!
1%
1-
12
#900620000000
0!
0%
b111 *
0-
02
b111 6
#900630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#900640000000
0!
0%
b0 *
0-
02
b0 6
#900650000000
1!
1%
1-
12
#900660000000
0!
0%
b1 *
0-
02
b1 6
#900670000000
1!
1%
1-
12
#900680000000
0!
0%
b10 *
0-
02
b10 6
#900690000000
1!
1%
1-
12
#900700000000
0!
0%
b11 *
0-
02
b11 6
#900710000000
1!
1%
1-
12
15
#900720000000
0!
0%
b100 *
0-
02
b100 6
#900730000000
1!
1%
1-
12
#900740000000
0!
0%
b101 *
0-
02
b101 6
#900750000000
1!
1%
1-
12
#900760000000
0!
0%
b110 *
0-
02
b110 6
#900770000000
1!
1%
1-
12
#900780000000
0!
0%
b111 *
0-
02
b111 6
#900790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#900800000000
0!
0%
b0 *
0-
02
b0 6
#900810000000
1!
1%
1-
12
#900820000000
0!
0%
b1 *
0-
02
b1 6
#900830000000
1!
1%
1-
12
#900840000000
0!
0%
b10 *
0-
02
b10 6
#900850000000
1!
1%
1-
12
#900860000000
0!
0%
b11 *
0-
02
b11 6
#900870000000
1!
1%
1-
12
15
#900880000000
0!
0%
b100 *
0-
02
b100 6
#900890000000
1!
1%
1-
12
#900900000000
0!
0%
b101 *
0-
02
b101 6
#900910000000
1!
1%
1-
12
#900920000000
0!
0%
b110 *
0-
02
b110 6
#900930000000
1!
1%
1-
12
#900940000000
0!
0%
b111 *
0-
02
b111 6
#900950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#900960000000
0!
0%
b0 *
0-
02
b0 6
#900970000000
1!
1%
1-
12
#900980000000
0!
0%
b1 *
0-
02
b1 6
#900990000000
1!
1%
1-
12
#901000000000
0!
0%
b10 *
0-
02
b10 6
#901010000000
1!
1%
1-
12
#901020000000
0!
0%
b11 *
0-
02
b11 6
#901030000000
1!
1%
1-
12
15
#901040000000
0!
0%
b100 *
0-
02
b100 6
#901050000000
1!
1%
1-
12
#901060000000
0!
0%
b101 *
0-
02
b101 6
#901070000000
1!
1%
1-
12
#901080000000
0!
0%
b110 *
0-
02
b110 6
#901090000000
1!
1%
1-
12
#901100000000
0!
0%
b111 *
0-
02
b111 6
#901110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#901120000000
0!
0%
b0 *
0-
02
b0 6
#901130000000
1!
1%
1-
12
#901140000000
0!
0%
b1 *
0-
02
b1 6
#901150000000
1!
1%
1-
12
#901160000000
0!
0%
b10 *
0-
02
b10 6
#901170000000
1!
1%
1-
12
#901180000000
0!
0%
b11 *
0-
02
b11 6
#901190000000
1!
1%
1-
12
15
#901200000000
0!
0%
b100 *
0-
02
b100 6
#901210000000
1!
1%
1-
12
#901220000000
0!
0%
b101 *
0-
02
b101 6
#901230000000
1!
1%
1-
12
#901240000000
0!
0%
b110 *
0-
02
b110 6
#901250000000
1!
1%
1-
12
#901260000000
0!
0%
b111 *
0-
02
b111 6
#901270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#901280000000
0!
0%
b0 *
0-
02
b0 6
#901290000000
1!
1%
1-
12
#901300000000
0!
0%
b1 *
0-
02
b1 6
#901310000000
1!
1%
1-
12
#901320000000
0!
0%
b10 *
0-
02
b10 6
#901330000000
1!
1%
1-
12
#901340000000
0!
0%
b11 *
0-
02
b11 6
#901350000000
1!
1%
1-
12
15
#901360000000
0!
0%
b100 *
0-
02
b100 6
#901370000000
1!
1%
1-
12
#901380000000
0!
0%
b101 *
0-
02
b101 6
#901390000000
1!
1%
1-
12
#901400000000
0!
0%
b110 *
0-
02
b110 6
#901410000000
1!
1%
1-
12
#901420000000
0!
0%
b111 *
0-
02
b111 6
#901430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#901440000000
0!
0%
b0 *
0-
02
b0 6
#901450000000
1!
1%
1-
12
#901460000000
0!
0%
b1 *
0-
02
b1 6
#901470000000
1!
1%
1-
12
#901480000000
0!
0%
b10 *
0-
02
b10 6
#901490000000
1!
1%
1-
12
#901500000000
0!
0%
b11 *
0-
02
b11 6
#901510000000
1!
1%
1-
12
15
#901520000000
0!
0%
b100 *
0-
02
b100 6
#901530000000
1!
1%
1-
12
#901540000000
0!
0%
b101 *
0-
02
b101 6
#901550000000
1!
1%
1-
12
#901560000000
0!
0%
b110 *
0-
02
b110 6
#901570000000
1!
1%
1-
12
#901580000000
0!
0%
b111 *
0-
02
b111 6
#901590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#901600000000
0!
0%
b0 *
0-
02
b0 6
#901610000000
1!
1%
1-
12
#901620000000
0!
0%
b1 *
0-
02
b1 6
#901630000000
1!
1%
1-
12
#901640000000
0!
0%
b10 *
0-
02
b10 6
#901650000000
1!
1%
1-
12
#901660000000
0!
0%
b11 *
0-
02
b11 6
#901670000000
1!
1%
1-
12
15
#901680000000
0!
0%
b100 *
0-
02
b100 6
#901690000000
1!
1%
1-
12
#901700000000
0!
0%
b101 *
0-
02
b101 6
#901710000000
1!
1%
1-
12
#901720000000
0!
0%
b110 *
0-
02
b110 6
#901730000000
1!
1%
1-
12
#901740000000
0!
0%
b111 *
0-
02
b111 6
#901750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#901760000000
0!
0%
b0 *
0-
02
b0 6
#901770000000
1!
1%
1-
12
#901780000000
0!
0%
b1 *
0-
02
b1 6
#901790000000
1!
1%
1-
12
#901800000000
0!
0%
b10 *
0-
02
b10 6
#901810000000
1!
1%
1-
12
#901820000000
0!
0%
b11 *
0-
02
b11 6
#901830000000
1!
1%
1-
12
15
#901840000000
0!
0%
b100 *
0-
02
b100 6
#901850000000
1!
1%
1-
12
#901860000000
0!
0%
b101 *
0-
02
b101 6
#901870000000
1!
1%
1-
12
#901880000000
0!
0%
b110 *
0-
02
b110 6
#901890000000
1!
1%
1-
12
#901900000000
0!
0%
b111 *
0-
02
b111 6
#901910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#901920000000
0!
0%
b0 *
0-
02
b0 6
#901930000000
1!
1%
1-
12
#901940000000
0!
0%
b1 *
0-
02
b1 6
#901950000000
1!
1%
1-
12
#901960000000
0!
0%
b10 *
0-
02
b10 6
#901970000000
1!
1%
1-
12
#901980000000
0!
0%
b11 *
0-
02
b11 6
#901990000000
1!
1%
1-
12
15
#902000000000
0!
0%
b100 *
0-
02
b100 6
#902010000000
1!
1%
1-
12
#902020000000
0!
0%
b101 *
0-
02
b101 6
#902030000000
1!
1%
1-
12
#902040000000
0!
0%
b110 *
0-
02
b110 6
#902050000000
1!
1%
1-
12
#902060000000
0!
0%
b111 *
0-
02
b111 6
#902070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#902080000000
0!
0%
b0 *
0-
02
b0 6
#902090000000
1!
1%
1-
12
#902100000000
0!
0%
b1 *
0-
02
b1 6
#902110000000
1!
1%
1-
12
#902120000000
0!
0%
b10 *
0-
02
b10 6
#902130000000
1!
1%
1-
12
#902140000000
0!
0%
b11 *
0-
02
b11 6
#902150000000
1!
1%
1-
12
15
#902160000000
0!
0%
b100 *
0-
02
b100 6
#902170000000
1!
1%
1-
12
#902180000000
0!
0%
b101 *
0-
02
b101 6
#902190000000
1!
1%
1-
12
#902200000000
0!
0%
b110 *
0-
02
b110 6
#902210000000
1!
1%
1-
12
#902220000000
0!
0%
b111 *
0-
02
b111 6
#902230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#902240000000
0!
0%
b0 *
0-
02
b0 6
#902250000000
1!
1%
1-
12
#902260000000
0!
0%
b1 *
0-
02
b1 6
#902270000000
1!
1%
1-
12
#902280000000
0!
0%
b10 *
0-
02
b10 6
#902290000000
1!
1%
1-
12
#902300000000
0!
0%
b11 *
0-
02
b11 6
#902310000000
1!
1%
1-
12
15
#902320000000
0!
0%
b100 *
0-
02
b100 6
#902330000000
1!
1%
1-
12
#902340000000
0!
0%
b101 *
0-
02
b101 6
#902350000000
1!
1%
1-
12
#902360000000
0!
0%
b110 *
0-
02
b110 6
#902370000000
1!
1%
1-
12
#902380000000
0!
0%
b111 *
0-
02
b111 6
#902390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#902400000000
0!
0%
b0 *
0-
02
b0 6
#902410000000
1!
1%
1-
12
#902420000000
0!
0%
b1 *
0-
02
b1 6
#902430000000
1!
1%
1-
12
#902440000000
0!
0%
b10 *
0-
02
b10 6
#902450000000
1!
1%
1-
12
#902460000000
0!
0%
b11 *
0-
02
b11 6
#902470000000
1!
1%
1-
12
15
#902480000000
0!
0%
b100 *
0-
02
b100 6
#902490000000
1!
1%
1-
12
#902500000000
0!
0%
b101 *
0-
02
b101 6
#902510000000
1!
1%
1-
12
#902520000000
0!
0%
b110 *
0-
02
b110 6
#902530000000
1!
1%
1-
12
#902540000000
0!
0%
b111 *
0-
02
b111 6
#902550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#902560000000
0!
0%
b0 *
0-
02
b0 6
#902570000000
1!
1%
1-
12
#902580000000
0!
0%
b1 *
0-
02
b1 6
#902590000000
1!
1%
1-
12
#902600000000
0!
0%
b10 *
0-
02
b10 6
#902610000000
1!
1%
1-
12
#902620000000
0!
0%
b11 *
0-
02
b11 6
#902630000000
1!
1%
1-
12
15
#902640000000
0!
0%
b100 *
0-
02
b100 6
#902650000000
1!
1%
1-
12
#902660000000
0!
0%
b101 *
0-
02
b101 6
#902670000000
1!
1%
1-
12
#902680000000
0!
0%
b110 *
0-
02
b110 6
#902690000000
1!
1%
1-
12
#902700000000
0!
0%
b111 *
0-
02
b111 6
#902710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#902720000000
0!
0%
b0 *
0-
02
b0 6
#902730000000
1!
1%
1-
12
#902740000000
0!
0%
b1 *
0-
02
b1 6
#902750000000
1!
1%
1-
12
#902760000000
0!
0%
b10 *
0-
02
b10 6
#902770000000
1!
1%
1-
12
#902780000000
0!
0%
b11 *
0-
02
b11 6
#902790000000
1!
1%
1-
12
15
#902800000000
0!
0%
b100 *
0-
02
b100 6
#902810000000
1!
1%
1-
12
#902820000000
0!
0%
b101 *
0-
02
b101 6
#902830000000
1!
1%
1-
12
#902840000000
0!
0%
b110 *
0-
02
b110 6
#902850000000
1!
1%
1-
12
#902860000000
0!
0%
b111 *
0-
02
b111 6
#902870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#902880000000
0!
0%
b0 *
0-
02
b0 6
#902890000000
1!
1%
1-
12
#902900000000
0!
0%
b1 *
0-
02
b1 6
#902910000000
1!
1%
1-
12
#902920000000
0!
0%
b10 *
0-
02
b10 6
#902930000000
1!
1%
1-
12
#902940000000
0!
0%
b11 *
0-
02
b11 6
#902950000000
1!
1%
1-
12
15
#902960000000
0!
0%
b100 *
0-
02
b100 6
#902970000000
1!
1%
1-
12
#902980000000
0!
0%
b101 *
0-
02
b101 6
#902990000000
1!
1%
1-
12
#903000000000
0!
0%
b110 *
0-
02
b110 6
#903010000000
1!
1%
1-
12
#903020000000
0!
0%
b111 *
0-
02
b111 6
#903030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#903040000000
0!
0%
b0 *
0-
02
b0 6
#903050000000
1!
1%
1-
12
#903060000000
0!
0%
b1 *
0-
02
b1 6
#903070000000
1!
1%
1-
12
#903080000000
0!
0%
b10 *
0-
02
b10 6
#903090000000
1!
1%
1-
12
#903100000000
0!
0%
b11 *
0-
02
b11 6
#903110000000
1!
1%
1-
12
15
#903120000000
0!
0%
b100 *
0-
02
b100 6
#903130000000
1!
1%
1-
12
#903140000000
0!
0%
b101 *
0-
02
b101 6
#903150000000
1!
1%
1-
12
#903160000000
0!
0%
b110 *
0-
02
b110 6
#903170000000
1!
1%
1-
12
#903180000000
0!
0%
b111 *
0-
02
b111 6
#903190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#903200000000
0!
0%
b0 *
0-
02
b0 6
#903210000000
1!
1%
1-
12
#903220000000
0!
0%
b1 *
0-
02
b1 6
#903230000000
1!
1%
1-
12
#903240000000
0!
0%
b10 *
0-
02
b10 6
#903250000000
1!
1%
1-
12
#903260000000
0!
0%
b11 *
0-
02
b11 6
#903270000000
1!
1%
1-
12
15
#903280000000
0!
0%
b100 *
0-
02
b100 6
#903290000000
1!
1%
1-
12
#903300000000
0!
0%
b101 *
0-
02
b101 6
#903310000000
1!
1%
1-
12
#903320000000
0!
0%
b110 *
0-
02
b110 6
#903330000000
1!
1%
1-
12
#903340000000
0!
0%
b111 *
0-
02
b111 6
#903350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#903360000000
0!
0%
b0 *
0-
02
b0 6
#903370000000
1!
1%
1-
12
#903380000000
0!
0%
b1 *
0-
02
b1 6
#903390000000
1!
1%
1-
12
#903400000000
0!
0%
b10 *
0-
02
b10 6
#903410000000
1!
1%
1-
12
#903420000000
0!
0%
b11 *
0-
02
b11 6
#903430000000
1!
1%
1-
12
15
#903440000000
0!
0%
b100 *
0-
02
b100 6
#903450000000
1!
1%
1-
12
#903460000000
0!
0%
b101 *
0-
02
b101 6
#903470000000
1!
1%
1-
12
#903480000000
0!
0%
b110 *
0-
02
b110 6
#903490000000
1!
1%
1-
12
#903500000000
0!
0%
b111 *
0-
02
b111 6
#903510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#903520000000
0!
0%
b0 *
0-
02
b0 6
#903530000000
1!
1%
1-
12
#903540000000
0!
0%
b1 *
0-
02
b1 6
#903550000000
1!
1%
1-
12
#903560000000
0!
0%
b10 *
0-
02
b10 6
#903570000000
1!
1%
1-
12
#903580000000
0!
0%
b11 *
0-
02
b11 6
#903590000000
1!
1%
1-
12
15
#903600000000
0!
0%
b100 *
0-
02
b100 6
#903610000000
1!
1%
1-
12
#903620000000
0!
0%
b101 *
0-
02
b101 6
#903630000000
1!
1%
1-
12
#903640000000
0!
0%
b110 *
0-
02
b110 6
#903650000000
1!
1%
1-
12
#903660000000
0!
0%
b111 *
0-
02
b111 6
#903670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#903680000000
0!
0%
b0 *
0-
02
b0 6
#903690000000
1!
1%
1-
12
#903700000000
0!
0%
b1 *
0-
02
b1 6
#903710000000
1!
1%
1-
12
#903720000000
0!
0%
b10 *
0-
02
b10 6
#903730000000
1!
1%
1-
12
#903740000000
0!
0%
b11 *
0-
02
b11 6
#903750000000
1!
1%
1-
12
15
#903760000000
0!
0%
b100 *
0-
02
b100 6
#903770000000
1!
1%
1-
12
#903780000000
0!
0%
b101 *
0-
02
b101 6
#903790000000
1!
1%
1-
12
#903800000000
0!
0%
b110 *
0-
02
b110 6
#903810000000
1!
1%
1-
12
#903820000000
0!
0%
b111 *
0-
02
b111 6
#903830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#903840000000
0!
0%
b0 *
0-
02
b0 6
#903850000000
1!
1%
1-
12
#903860000000
0!
0%
b1 *
0-
02
b1 6
#903870000000
1!
1%
1-
12
#903880000000
0!
0%
b10 *
0-
02
b10 6
#903890000000
1!
1%
1-
12
#903900000000
0!
0%
b11 *
0-
02
b11 6
#903910000000
1!
1%
1-
12
15
#903920000000
0!
0%
b100 *
0-
02
b100 6
#903930000000
1!
1%
1-
12
#903940000000
0!
0%
b101 *
0-
02
b101 6
#903950000000
1!
1%
1-
12
#903960000000
0!
0%
b110 *
0-
02
b110 6
#903970000000
1!
1%
1-
12
#903980000000
0!
0%
b111 *
0-
02
b111 6
#903990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#904000000000
0!
0%
b0 *
0-
02
b0 6
#904010000000
1!
1%
1-
12
#904020000000
0!
0%
b1 *
0-
02
b1 6
#904030000000
1!
1%
1-
12
#904040000000
0!
0%
b10 *
0-
02
b10 6
#904050000000
1!
1%
1-
12
#904060000000
0!
0%
b11 *
0-
02
b11 6
#904070000000
1!
1%
1-
12
15
#904080000000
0!
0%
b100 *
0-
02
b100 6
#904090000000
1!
1%
1-
12
#904100000000
0!
0%
b101 *
0-
02
b101 6
#904110000000
1!
1%
1-
12
#904120000000
0!
0%
b110 *
0-
02
b110 6
#904130000000
1!
1%
1-
12
#904140000000
0!
0%
b111 *
0-
02
b111 6
#904150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#904160000000
0!
0%
b0 *
0-
02
b0 6
#904170000000
1!
1%
1-
12
#904180000000
0!
0%
b1 *
0-
02
b1 6
#904190000000
1!
1%
1-
12
#904200000000
0!
0%
b10 *
0-
02
b10 6
#904210000000
1!
1%
1-
12
#904220000000
0!
0%
b11 *
0-
02
b11 6
#904230000000
1!
1%
1-
12
15
#904240000000
0!
0%
b100 *
0-
02
b100 6
#904250000000
1!
1%
1-
12
#904260000000
0!
0%
b101 *
0-
02
b101 6
#904270000000
1!
1%
1-
12
#904280000000
0!
0%
b110 *
0-
02
b110 6
#904290000000
1!
1%
1-
12
#904300000000
0!
0%
b111 *
0-
02
b111 6
#904310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#904320000000
0!
0%
b0 *
0-
02
b0 6
#904330000000
1!
1%
1-
12
#904340000000
0!
0%
b1 *
0-
02
b1 6
#904350000000
1!
1%
1-
12
#904360000000
0!
0%
b10 *
0-
02
b10 6
#904370000000
1!
1%
1-
12
#904380000000
0!
0%
b11 *
0-
02
b11 6
#904390000000
1!
1%
1-
12
15
#904400000000
0!
0%
b100 *
0-
02
b100 6
#904410000000
1!
1%
1-
12
#904420000000
0!
0%
b101 *
0-
02
b101 6
#904430000000
1!
1%
1-
12
#904440000000
0!
0%
b110 *
0-
02
b110 6
#904450000000
1!
1%
1-
12
#904460000000
0!
0%
b111 *
0-
02
b111 6
#904470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#904480000000
0!
0%
b0 *
0-
02
b0 6
#904490000000
1!
1%
1-
12
#904500000000
0!
0%
b1 *
0-
02
b1 6
#904510000000
1!
1%
1-
12
#904520000000
0!
0%
b10 *
0-
02
b10 6
#904530000000
1!
1%
1-
12
#904540000000
0!
0%
b11 *
0-
02
b11 6
#904550000000
1!
1%
1-
12
15
#904560000000
0!
0%
b100 *
0-
02
b100 6
#904570000000
1!
1%
1-
12
#904580000000
0!
0%
b101 *
0-
02
b101 6
#904590000000
1!
1%
1-
12
#904600000000
0!
0%
b110 *
0-
02
b110 6
#904610000000
1!
1%
1-
12
#904620000000
0!
0%
b111 *
0-
02
b111 6
#904630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#904640000000
0!
0%
b0 *
0-
02
b0 6
#904650000000
1!
1%
1-
12
#904660000000
0!
0%
b1 *
0-
02
b1 6
#904670000000
1!
1%
1-
12
#904680000000
0!
0%
b10 *
0-
02
b10 6
#904690000000
1!
1%
1-
12
#904700000000
0!
0%
b11 *
0-
02
b11 6
#904710000000
1!
1%
1-
12
15
#904720000000
0!
0%
b100 *
0-
02
b100 6
#904730000000
1!
1%
1-
12
#904740000000
0!
0%
b101 *
0-
02
b101 6
#904750000000
1!
1%
1-
12
#904760000000
0!
0%
b110 *
0-
02
b110 6
#904770000000
1!
1%
1-
12
#904780000000
0!
0%
b111 *
0-
02
b111 6
#904790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#904800000000
0!
0%
b0 *
0-
02
b0 6
#904810000000
1!
1%
1-
12
#904820000000
0!
0%
b1 *
0-
02
b1 6
#904830000000
1!
1%
1-
12
#904840000000
0!
0%
b10 *
0-
02
b10 6
#904850000000
1!
1%
1-
12
#904860000000
0!
0%
b11 *
0-
02
b11 6
#904870000000
1!
1%
1-
12
15
#904880000000
0!
0%
b100 *
0-
02
b100 6
#904890000000
1!
1%
1-
12
#904900000000
0!
0%
b101 *
0-
02
b101 6
#904910000000
1!
1%
1-
12
#904920000000
0!
0%
b110 *
0-
02
b110 6
#904930000000
1!
1%
1-
12
#904940000000
0!
0%
b111 *
0-
02
b111 6
#904950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#904960000000
0!
0%
b0 *
0-
02
b0 6
#904970000000
1!
1%
1-
12
#904980000000
0!
0%
b1 *
0-
02
b1 6
#904990000000
1!
1%
1-
12
#905000000000
0!
0%
b10 *
0-
02
b10 6
#905010000000
1!
1%
1-
12
#905020000000
0!
0%
b11 *
0-
02
b11 6
#905030000000
1!
1%
1-
12
15
#905040000000
0!
0%
b100 *
0-
02
b100 6
#905050000000
1!
1%
1-
12
#905060000000
0!
0%
b101 *
0-
02
b101 6
#905070000000
1!
1%
1-
12
#905080000000
0!
0%
b110 *
0-
02
b110 6
#905090000000
1!
1%
1-
12
#905100000000
0!
0%
b111 *
0-
02
b111 6
#905110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#905120000000
0!
0%
b0 *
0-
02
b0 6
#905130000000
1!
1%
1-
12
#905140000000
0!
0%
b1 *
0-
02
b1 6
#905150000000
1!
1%
1-
12
#905160000000
0!
0%
b10 *
0-
02
b10 6
#905170000000
1!
1%
1-
12
#905180000000
0!
0%
b11 *
0-
02
b11 6
#905190000000
1!
1%
1-
12
15
#905200000000
0!
0%
b100 *
0-
02
b100 6
#905210000000
1!
1%
1-
12
#905220000000
0!
0%
b101 *
0-
02
b101 6
#905230000000
1!
1%
1-
12
#905240000000
0!
0%
b110 *
0-
02
b110 6
#905250000000
1!
1%
1-
12
#905260000000
0!
0%
b111 *
0-
02
b111 6
#905270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#905280000000
0!
0%
b0 *
0-
02
b0 6
#905290000000
1!
1%
1-
12
#905300000000
0!
0%
b1 *
0-
02
b1 6
#905310000000
1!
1%
1-
12
#905320000000
0!
0%
b10 *
0-
02
b10 6
#905330000000
1!
1%
1-
12
#905340000000
0!
0%
b11 *
0-
02
b11 6
#905350000000
1!
1%
1-
12
15
#905360000000
0!
0%
b100 *
0-
02
b100 6
#905370000000
1!
1%
1-
12
#905380000000
0!
0%
b101 *
0-
02
b101 6
#905390000000
1!
1%
1-
12
#905400000000
0!
0%
b110 *
0-
02
b110 6
#905410000000
1!
1%
1-
12
#905420000000
0!
0%
b111 *
0-
02
b111 6
#905430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#905440000000
0!
0%
b0 *
0-
02
b0 6
#905450000000
1!
1%
1-
12
#905460000000
0!
0%
b1 *
0-
02
b1 6
#905470000000
1!
1%
1-
12
#905480000000
0!
0%
b10 *
0-
02
b10 6
#905490000000
1!
1%
1-
12
#905500000000
0!
0%
b11 *
0-
02
b11 6
#905510000000
1!
1%
1-
12
15
#905520000000
0!
0%
b100 *
0-
02
b100 6
#905530000000
1!
1%
1-
12
#905540000000
0!
0%
b101 *
0-
02
b101 6
#905550000000
1!
1%
1-
12
#905560000000
0!
0%
b110 *
0-
02
b110 6
#905570000000
1!
1%
1-
12
#905580000000
0!
0%
b111 *
0-
02
b111 6
#905590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#905600000000
0!
0%
b0 *
0-
02
b0 6
#905610000000
1!
1%
1-
12
#905620000000
0!
0%
b1 *
0-
02
b1 6
#905630000000
1!
1%
1-
12
#905640000000
0!
0%
b10 *
0-
02
b10 6
#905650000000
1!
1%
1-
12
#905660000000
0!
0%
b11 *
0-
02
b11 6
#905670000000
1!
1%
1-
12
15
#905680000000
0!
0%
b100 *
0-
02
b100 6
#905690000000
1!
1%
1-
12
#905700000000
0!
0%
b101 *
0-
02
b101 6
#905710000000
1!
1%
1-
12
#905720000000
0!
0%
b110 *
0-
02
b110 6
#905730000000
1!
1%
1-
12
#905740000000
0!
0%
b111 *
0-
02
b111 6
#905750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#905760000000
0!
0%
b0 *
0-
02
b0 6
#905770000000
1!
1%
1-
12
#905780000000
0!
0%
b1 *
0-
02
b1 6
#905790000000
1!
1%
1-
12
#905800000000
0!
0%
b10 *
0-
02
b10 6
#905810000000
1!
1%
1-
12
#905820000000
0!
0%
b11 *
0-
02
b11 6
#905830000000
1!
1%
1-
12
15
#905840000000
0!
0%
b100 *
0-
02
b100 6
#905850000000
1!
1%
1-
12
#905860000000
0!
0%
b101 *
0-
02
b101 6
#905870000000
1!
1%
1-
12
#905880000000
0!
0%
b110 *
0-
02
b110 6
#905890000000
1!
1%
1-
12
#905900000000
0!
0%
b111 *
0-
02
b111 6
#905910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#905920000000
0!
0%
b0 *
0-
02
b0 6
#905930000000
1!
1%
1-
12
#905940000000
0!
0%
b1 *
0-
02
b1 6
#905950000000
1!
1%
1-
12
#905960000000
0!
0%
b10 *
0-
02
b10 6
#905970000000
1!
1%
1-
12
#905980000000
0!
0%
b11 *
0-
02
b11 6
#905990000000
1!
1%
1-
12
15
#906000000000
0!
0%
b100 *
0-
02
b100 6
#906010000000
1!
1%
1-
12
#906020000000
0!
0%
b101 *
0-
02
b101 6
#906030000000
1!
1%
1-
12
#906040000000
0!
0%
b110 *
0-
02
b110 6
#906050000000
1!
1%
1-
12
#906060000000
0!
0%
b111 *
0-
02
b111 6
#906070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#906080000000
0!
0%
b0 *
0-
02
b0 6
#906090000000
1!
1%
1-
12
#906100000000
0!
0%
b1 *
0-
02
b1 6
#906110000000
1!
1%
1-
12
#906120000000
0!
0%
b10 *
0-
02
b10 6
#906130000000
1!
1%
1-
12
#906140000000
0!
0%
b11 *
0-
02
b11 6
#906150000000
1!
1%
1-
12
15
#906160000000
0!
0%
b100 *
0-
02
b100 6
#906170000000
1!
1%
1-
12
#906180000000
0!
0%
b101 *
0-
02
b101 6
#906190000000
1!
1%
1-
12
#906200000000
0!
0%
b110 *
0-
02
b110 6
#906210000000
1!
1%
1-
12
#906220000000
0!
0%
b111 *
0-
02
b111 6
#906230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#906240000000
0!
0%
b0 *
0-
02
b0 6
#906250000000
1!
1%
1-
12
#906260000000
0!
0%
b1 *
0-
02
b1 6
#906270000000
1!
1%
1-
12
#906280000000
0!
0%
b10 *
0-
02
b10 6
#906290000000
1!
1%
1-
12
#906300000000
0!
0%
b11 *
0-
02
b11 6
#906310000000
1!
1%
1-
12
15
#906320000000
0!
0%
b100 *
0-
02
b100 6
#906330000000
1!
1%
1-
12
#906340000000
0!
0%
b101 *
0-
02
b101 6
#906350000000
1!
1%
1-
12
#906360000000
0!
0%
b110 *
0-
02
b110 6
#906370000000
1!
1%
1-
12
#906380000000
0!
0%
b111 *
0-
02
b111 6
#906390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#906400000000
0!
0%
b0 *
0-
02
b0 6
#906410000000
1!
1%
1-
12
#906420000000
0!
0%
b1 *
0-
02
b1 6
#906430000000
1!
1%
1-
12
#906440000000
0!
0%
b10 *
0-
02
b10 6
#906450000000
1!
1%
1-
12
#906460000000
0!
0%
b11 *
0-
02
b11 6
#906470000000
1!
1%
1-
12
15
#906480000000
0!
0%
b100 *
0-
02
b100 6
#906490000000
1!
1%
1-
12
#906500000000
0!
0%
b101 *
0-
02
b101 6
#906510000000
1!
1%
1-
12
#906520000000
0!
0%
b110 *
0-
02
b110 6
#906530000000
1!
1%
1-
12
#906540000000
0!
0%
b111 *
0-
02
b111 6
#906550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#906560000000
0!
0%
b0 *
0-
02
b0 6
#906570000000
1!
1%
1-
12
#906580000000
0!
0%
b1 *
0-
02
b1 6
#906590000000
1!
1%
1-
12
#906600000000
0!
0%
b10 *
0-
02
b10 6
#906610000000
1!
1%
1-
12
#906620000000
0!
0%
b11 *
0-
02
b11 6
#906630000000
1!
1%
1-
12
15
#906640000000
0!
0%
b100 *
0-
02
b100 6
#906650000000
1!
1%
1-
12
#906660000000
0!
0%
b101 *
0-
02
b101 6
#906670000000
1!
1%
1-
12
#906680000000
0!
0%
b110 *
0-
02
b110 6
#906690000000
1!
1%
1-
12
#906700000000
0!
0%
b111 *
0-
02
b111 6
#906710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#906720000000
0!
0%
b0 *
0-
02
b0 6
#906730000000
1!
1%
1-
12
#906740000000
0!
0%
b1 *
0-
02
b1 6
#906750000000
1!
1%
1-
12
#906760000000
0!
0%
b10 *
0-
02
b10 6
#906770000000
1!
1%
1-
12
#906780000000
0!
0%
b11 *
0-
02
b11 6
#906790000000
1!
1%
1-
12
15
#906800000000
0!
0%
b100 *
0-
02
b100 6
#906810000000
1!
1%
1-
12
#906820000000
0!
0%
b101 *
0-
02
b101 6
#906830000000
1!
1%
1-
12
#906840000000
0!
0%
b110 *
0-
02
b110 6
#906850000000
1!
1%
1-
12
#906860000000
0!
0%
b111 *
0-
02
b111 6
#906870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#906880000000
0!
0%
b0 *
0-
02
b0 6
#906890000000
1!
1%
1-
12
#906900000000
0!
0%
b1 *
0-
02
b1 6
#906910000000
1!
1%
1-
12
#906920000000
0!
0%
b10 *
0-
02
b10 6
#906930000000
1!
1%
1-
12
#906940000000
0!
0%
b11 *
0-
02
b11 6
#906950000000
1!
1%
1-
12
15
#906960000000
0!
0%
b100 *
0-
02
b100 6
#906970000000
1!
1%
1-
12
#906980000000
0!
0%
b101 *
0-
02
b101 6
#906990000000
1!
1%
1-
12
#907000000000
0!
0%
b110 *
0-
02
b110 6
#907010000000
1!
1%
1-
12
#907020000000
0!
0%
b111 *
0-
02
b111 6
#907030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#907040000000
0!
0%
b0 *
0-
02
b0 6
#907050000000
1!
1%
1-
12
#907060000000
0!
0%
b1 *
0-
02
b1 6
#907070000000
1!
1%
1-
12
#907080000000
0!
0%
b10 *
0-
02
b10 6
#907090000000
1!
1%
1-
12
#907100000000
0!
0%
b11 *
0-
02
b11 6
#907110000000
1!
1%
1-
12
15
#907120000000
0!
0%
b100 *
0-
02
b100 6
#907130000000
1!
1%
1-
12
#907140000000
0!
0%
b101 *
0-
02
b101 6
#907150000000
1!
1%
1-
12
#907160000000
0!
0%
b110 *
0-
02
b110 6
#907170000000
1!
1%
1-
12
#907180000000
0!
0%
b111 *
0-
02
b111 6
#907190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#907200000000
0!
0%
b0 *
0-
02
b0 6
#907210000000
1!
1%
1-
12
#907220000000
0!
0%
b1 *
0-
02
b1 6
#907230000000
1!
1%
1-
12
#907240000000
0!
0%
b10 *
0-
02
b10 6
#907250000000
1!
1%
1-
12
#907260000000
0!
0%
b11 *
0-
02
b11 6
#907270000000
1!
1%
1-
12
15
#907280000000
0!
0%
b100 *
0-
02
b100 6
#907290000000
1!
1%
1-
12
#907300000000
0!
0%
b101 *
0-
02
b101 6
#907310000000
1!
1%
1-
12
#907320000000
0!
0%
b110 *
0-
02
b110 6
#907330000000
1!
1%
1-
12
#907340000000
0!
0%
b111 *
0-
02
b111 6
#907350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#907360000000
0!
0%
b0 *
0-
02
b0 6
#907370000000
1!
1%
1-
12
#907380000000
0!
0%
b1 *
0-
02
b1 6
#907390000000
1!
1%
1-
12
#907400000000
0!
0%
b10 *
0-
02
b10 6
#907410000000
1!
1%
1-
12
#907420000000
0!
0%
b11 *
0-
02
b11 6
#907430000000
1!
1%
1-
12
15
#907440000000
0!
0%
b100 *
0-
02
b100 6
#907450000000
1!
1%
1-
12
#907460000000
0!
0%
b101 *
0-
02
b101 6
#907470000000
1!
1%
1-
12
#907480000000
0!
0%
b110 *
0-
02
b110 6
#907490000000
1!
1%
1-
12
#907500000000
0!
0%
b111 *
0-
02
b111 6
#907510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#907520000000
0!
0%
b0 *
0-
02
b0 6
#907530000000
1!
1%
1-
12
#907540000000
0!
0%
b1 *
0-
02
b1 6
#907550000000
1!
1%
1-
12
#907560000000
0!
0%
b10 *
0-
02
b10 6
#907570000000
1!
1%
1-
12
#907580000000
0!
0%
b11 *
0-
02
b11 6
#907590000000
1!
1%
1-
12
15
#907600000000
0!
0%
b100 *
0-
02
b100 6
#907610000000
1!
1%
1-
12
#907620000000
0!
0%
b101 *
0-
02
b101 6
#907630000000
1!
1%
1-
12
#907640000000
0!
0%
b110 *
0-
02
b110 6
#907650000000
1!
1%
1-
12
#907660000000
0!
0%
b111 *
0-
02
b111 6
#907670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#907680000000
0!
0%
b0 *
0-
02
b0 6
#907690000000
1!
1%
1-
12
#907700000000
0!
0%
b1 *
0-
02
b1 6
#907710000000
1!
1%
1-
12
#907720000000
0!
0%
b10 *
0-
02
b10 6
#907730000000
1!
1%
1-
12
#907740000000
0!
0%
b11 *
0-
02
b11 6
#907750000000
1!
1%
1-
12
15
#907760000000
0!
0%
b100 *
0-
02
b100 6
#907770000000
1!
1%
1-
12
#907780000000
0!
0%
b101 *
0-
02
b101 6
#907790000000
1!
1%
1-
12
#907800000000
0!
0%
b110 *
0-
02
b110 6
#907810000000
1!
1%
1-
12
#907820000000
0!
0%
b111 *
0-
02
b111 6
#907830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#907840000000
0!
0%
b0 *
0-
02
b0 6
#907850000000
1!
1%
1-
12
#907860000000
0!
0%
b1 *
0-
02
b1 6
#907870000000
1!
1%
1-
12
#907880000000
0!
0%
b10 *
0-
02
b10 6
#907890000000
1!
1%
1-
12
#907900000000
0!
0%
b11 *
0-
02
b11 6
#907910000000
1!
1%
1-
12
15
#907920000000
0!
0%
b100 *
0-
02
b100 6
#907930000000
1!
1%
1-
12
#907940000000
0!
0%
b101 *
0-
02
b101 6
#907950000000
1!
1%
1-
12
#907960000000
0!
0%
b110 *
0-
02
b110 6
#907970000000
1!
1%
1-
12
#907980000000
0!
0%
b111 *
0-
02
b111 6
#907990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#908000000000
0!
0%
b0 *
0-
02
b0 6
#908010000000
1!
1%
1-
12
#908020000000
0!
0%
b1 *
0-
02
b1 6
#908030000000
1!
1%
1-
12
#908040000000
0!
0%
b10 *
0-
02
b10 6
#908050000000
1!
1%
1-
12
#908060000000
0!
0%
b11 *
0-
02
b11 6
#908070000000
1!
1%
1-
12
15
#908080000000
0!
0%
b100 *
0-
02
b100 6
#908090000000
1!
1%
1-
12
#908100000000
0!
0%
b101 *
0-
02
b101 6
#908110000000
1!
1%
1-
12
#908120000000
0!
0%
b110 *
0-
02
b110 6
#908130000000
1!
1%
1-
12
#908140000000
0!
0%
b111 *
0-
02
b111 6
#908150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#908160000000
0!
0%
b0 *
0-
02
b0 6
#908170000000
1!
1%
1-
12
#908180000000
0!
0%
b1 *
0-
02
b1 6
#908190000000
1!
1%
1-
12
#908200000000
0!
0%
b10 *
0-
02
b10 6
#908210000000
1!
1%
1-
12
#908220000000
0!
0%
b11 *
0-
02
b11 6
#908230000000
1!
1%
1-
12
15
#908240000000
0!
0%
b100 *
0-
02
b100 6
#908250000000
1!
1%
1-
12
#908260000000
0!
0%
b101 *
0-
02
b101 6
#908270000000
1!
1%
1-
12
#908280000000
0!
0%
b110 *
0-
02
b110 6
#908290000000
1!
1%
1-
12
#908300000000
0!
0%
b111 *
0-
02
b111 6
#908310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#908320000000
0!
0%
b0 *
0-
02
b0 6
#908330000000
1!
1%
1-
12
#908340000000
0!
0%
b1 *
0-
02
b1 6
#908350000000
1!
1%
1-
12
#908360000000
0!
0%
b10 *
0-
02
b10 6
#908370000000
1!
1%
1-
12
#908380000000
0!
0%
b11 *
0-
02
b11 6
#908390000000
1!
1%
1-
12
15
#908400000000
0!
0%
b100 *
0-
02
b100 6
#908410000000
1!
1%
1-
12
#908420000000
0!
0%
b101 *
0-
02
b101 6
#908430000000
1!
1%
1-
12
#908440000000
0!
0%
b110 *
0-
02
b110 6
#908450000000
1!
1%
1-
12
#908460000000
0!
0%
b111 *
0-
02
b111 6
#908470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#908480000000
0!
0%
b0 *
0-
02
b0 6
#908490000000
1!
1%
1-
12
#908500000000
0!
0%
b1 *
0-
02
b1 6
#908510000000
1!
1%
1-
12
#908520000000
0!
0%
b10 *
0-
02
b10 6
#908530000000
1!
1%
1-
12
#908540000000
0!
0%
b11 *
0-
02
b11 6
#908550000000
1!
1%
1-
12
15
#908560000000
0!
0%
b100 *
0-
02
b100 6
#908570000000
1!
1%
1-
12
#908580000000
0!
0%
b101 *
0-
02
b101 6
#908590000000
1!
1%
1-
12
#908600000000
0!
0%
b110 *
0-
02
b110 6
#908610000000
1!
1%
1-
12
#908620000000
0!
0%
b111 *
0-
02
b111 6
#908630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#908640000000
0!
0%
b0 *
0-
02
b0 6
#908650000000
1!
1%
1-
12
#908660000000
0!
0%
b1 *
0-
02
b1 6
#908670000000
1!
1%
1-
12
#908680000000
0!
0%
b10 *
0-
02
b10 6
#908690000000
1!
1%
1-
12
#908700000000
0!
0%
b11 *
0-
02
b11 6
#908710000000
1!
1%
1-
12
15
#908720000000
0!
0%
b100 *
0-
02
b100 6
#908730000000
1!
1%
1-
12
#908740000000
0!
0%
b101 *
0-
02
b101 6
#908750000000
1!
1%
1-
12
#908760000000
0!
0%
b110 *
0-
02
b110 6
#908770000000
1!
1%
1-
12
#908780000000
0!
0%
b111 *
0-
02
b111 6
#908790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#908800000000
0!
0%
b0 *
0-
02
b0 6
#908810000000
1!
1%
1-
12
#908820000000
0!
0%
b1 *
0-
02
b1 6
#908830000000
1!
1%
1-
12
#908840000000
0!
0%
b10 *
0-
02
b10 6
#908850000000
1!
1%
1-
12
#908860000000
0!
0%
b11 *
0-
02
b11 6
#908870000000
1!
1%
1-
12
15
#908880000000
0!
0%
b100 *
0-
02
b100 6
#908890000000
1!
1%
1-
12
#908900000000
0!
0%
b101 *
0-
02
b101 6
#908910000000
1!
1%
1-
12
#908920000000
0!
0%
b110 *
0-
02
b110 6
#908930000000
1!
1%
1-
12
#908940000000
0!
0%
b111 *
0-
02
b111 6
#908950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#908960000000
0!
0%
b0 *
0-
02
b0 6
#908970000000
1!
1%
1-
12
#908980000000
0!
0%
b1 *
0-
02
b1 6
#908990000000
1!
1%
1-
12
#909000000000
0!
0%
b10 *
0-
02
b10 6
#909010000000
1!
1%
1-
12
#909020000000
0!
0%
b11 *
0-
02
b11 6
#909030000000
1!
1%
1-
12
15
#909040000000
0!
0%
b100 *
0-
02
b100 6
#909050000000
1!
1%
1-
12
#909060000000
0!
0%
b101 *
0-
02
b101 6
#909070000000
1!
1%
1-
12
#909080000000
0!
0%
b110 *
0-
02
b110 6
#909090000000
1!
1%
1-
12
#909100000000
0!
0%
b111 *
0-
02
b111 6
#909110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#909120000000
0!
0%
b0 *
0-
02
b0 6
#909130000000
1!
1%
1-
12
#909140000000
0!
0%
b1 *
0-
02
b1 6
#909150000000
1!
1%
1-
12
#909160000000
0!
0%
b10 *
0-
02
b10 6
#909170000000
1!
1%
1-
12
#909180000000
0!
0%
b11 *
0-
02
b11 6
#909190000000
1!
1%
1-
12
15
#909200000000
0!
0%
b100 *
0-
02
b100 6
#909210000000
1!
1%
1-
12
#909220000000
0!
0%
b101 *
0-
02
b101 6
#909230000000
1!
1%
1-
12
#909240000000
0!
0%
b110 *
0-
02
b110 6
#909250000000
1!
1%
1-
12
#909260000000
0!
0%
b111 *
0-
02
b111 6
#909270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#909280000000
0!
0%
b0 *
0-
02
b0 6
#909290000000
1!
1%
1-
12
#909300000000
0!
0%
b1 *
0-
02
b1 6
#909310000000
1!
1%
1-
12
#909320000000
0!
0%
b10 *
0-
02
b10 6
#909330000000
1!
1%
1-
12
#909340000000
0!
0%
b11 *
0-
02
b11 6
#909350000000
1!
1%
1-
12
15
#909360000000
0!
0%
b100 *
0-
02
b100 6
#909370000000
1!
1%
1-
12
#909380000000
0!
0%
b101 *
0-
02
b101 6
#909390000000
1!
1%
1-
12
#909400000000
0!
0%
b110 *
0-
02
b110 6
#909410000000
1!
1%
1-
12
#909420000000
0!
0%
b111 *
0-
02
b111 6
#909430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#909440000000
0!
0%
b0 *
0-
02
b0 6
#909450000000
1!
1%
1-
12
#909460000000
0!
0%
b1 *
0-
02
b1 6
#909470000000
1!
1%
1-
12
#909480000000
0!
0%
b10 *
0-
02
b10 6
#909490000000
1!
1%
1-
12
#909500000000
0!
0%
b11 *
0-
02
b11 6
#909510000000
1!
1%
1-
12
15
#909520000000
0!
0%
b100 *
0-
02
b100 6
#909530000000
1!
1%
1-
12
#909540000000
0!
0%
b101 *
0-
02
b101 6
#909550000000
1!
1%
1-
12
#909560000000
0!
0%
b110 *
0-
02
b110 6
#909570000000
1!
1%
1-
12
#909580000000
0!
0%
b111 *
0-
02
b111 6
#909590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#909600000000
0!
0%
b0 *
0-
02
b0 6
#909610000000
1!
1%
1-
12
#909620000000
0!
0%
b1 *
0-
02
b1 6
#909630000000
1!
1%
1-
12
#909640000000
0!
0%
b10 *
0-
02
b10 6
#909650000000
1!
1%
1-
12
#909660000000
0!
0%
b11 *
0-
02
b11 6
#909670000000
1!
1%
1-
12
15
#909680000000
0!
0%
b100 *
0-
02
b100 6
#909690000000
1!
1%
1-
12
#909700000000
0!
0%
b101 *
0-
02
b101 6
#909710000000
1!
1%
1-
12
#909720000000
0!
0%
b110 *
0-
02
b110 6
#909730000000
1!
1%
1-
12
#909740000000
0!
0%
b111 *
0-
02
b111 6
#909750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#909760000000
0!
0%
b0 *
0-
02
b0 6
#909770000000
1!
1%
1-
12
#909780000000
0!
0%
b1 *
0-
02
b1 6
#909790000000
1!
1%
1-
12
#909800000000
0!
0%
b10 *
0-
02
b10 6
#909810000000
1!
1%
1-
12
#909820000000
0!
0%
b11 *
0-
02
b11 6
#909830000000
1!
1%
1-
12
15
#909840000000
0!
0%
b100 *
0-
02
b100 6
#909850000000
1!
1%
1-
12
#909860000000
0!
0%
b101 *
0-
02
b101 6
#909870000000
1!
1%
1-
12
#909880000000
0!
0%
b110 *
0-
02
b110 6
#909890000000
1!
1%
1-
12
#909900000000
0!
0%
b111 *
0-
02
b111 6
#909910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#909920000000
0!
0%
b0 *
0-
02
b0 6
#909930000000
1!
1%
1-
12
#909940000000
0!
0%
b1 *
0-
02
b1 6
#909950000000
1!
1%
1-
12
#909960000000
0!
0%
b10 *
0-
02
b10 6
#909970000000
1!
1%
1-
12
#909980000000
0!
0%
b11 *
0-
02
b11 6
#909990000000
1!
1%
1-
12
15
#910000000000
0!
0%
b100 *
0-
02
b100 6
#910010000000
1!
1%
1-
12
#910020000000
0!
0%
b101 *
0-
02
b101 6
#910030000000
1!
1%
1-
12
#910040000000
0!
0%
b110 *
0-
02
b110 6
#910050000000
1!
1%
1-
12
#910060000000
0!
0%
b111 *
0-
02
b111 6
#910070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#910080000000
0!
0%
b0 *
0-
02
b0 6
#910090000000
1!
1%
1-
12
#910100000000
0!
0%
b1 *
0-
02
b1 6
#910110000000
1!
1%
1-
12
#910120000000
0!
0%
b10 *
0-
02
b10 6
#910130000000
1!
1%
1-
12
#910140000000
0!
0%
b11 *
0-
02
b11 6
#910150000000
1!
1%
1-
12
15
#910160000000
0!
0%
b100 *
0-
02
b100 6
#910170000000
1!
1%
1-
12
#910180000000
0!
0%
b101 *
0-
02
b101 6
#910190000000
1!
1%
1-
12
#910200000000
0!
0%
b110 *
0-
02
b110 6
#910210000000
1!
1%
1-
12
#910220000000
0!
0%
b111 *
0-
02
b111 6
#910230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#910240000000
0!
0%
b0 *
0-
02
b0 6
#910250000000
1!
1%
1-
12
#910260000000
0!
0%
b1 *
0-
02
b1 6
#910270000000
1!
1%
1-
12
#910280000000
0!
0%
b10 *
0-
02
b10 6
#910290000000
1!
1%
1-
12
#910300000000
0!
0%
b11 *
0-
02
b11 6
#910310000000
1!
1%
1-
12
15
#910320000000
0!
0%
b100 *
0-
02
b100 6
#910330000000
1!
1%
1-
12
#910340000000
0!
0%
b101 *
0-
02
b101 6
#910350000000
1!
1%
1-
12
#910360000000
0!
0%
b110 *
0-
02
b110 6
#910370000000
1!
1%
1-
12
#910380000000
0!
0%
b111 *
0-
02
b111 6
#910390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#910400000000
0!
0%
b0 *
0-
02
b0 6
#910410000000
1!
1%
1-
12
#910420000000
0!
0%
b1 *
0-
02
b1 6
#910430000000
1!
1%
1-
12
#910440000000
0!
0%
b10 *
0-
02
b10 6
#910450000000
1!
1%
1-
12
#910460000000
0!
0%
b11 *
0-
02
b11 6
#910470000000
1!
1%
1-
12
15
#910480000000
0!
0%
b100 *
0-
02
b100 6
#910490000000
1!
1%
1-
12
#910500000000
0!
0%
b101 *
0-
02
b101 6
#910510000000
1!
1%
1-
12
#910520000000
0!
0%
b110 *
0-
02
b110 6
#910530000000
1!
1%
1-
12
#910540000000
0!
0%
b111 *
0-
02
b111 6
#910550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#910560000000
0!
0%
b0 *
0-
02
b0 6
#910570000000
1!
1%
1-
12
#910580000000
0!
0%
b1 *
0-
02
b1 6
#910590000000
1!
1%
1-
12
#910600000000
0!
0%
b10 *
0-
02
b10 6
#910610000000
1!
1%
1-
12
#910620000000
0!
0%
b11 *
0-
02
b11 6
#910630000000
1!
1%
1-
12
15
#910640000000
0!
0%
b100 *
0-
02
b100 6
#910650000000
1!
1%
1-
12
#910660000000
0!
0%
b101 *
0-
02
b101 6
#910670000000
1!
1%
1-
12
#910680000000
0!
0%
b110 *
0-
02
b110 6
#910690000000
1!
1%
1-
12
#910700000000
0!
0%
b111 *
0-
02
b111 6
#910710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#910720000000
0!
0%
b0 *
0-
02
b0 6
#910730000000
1!
1%
1-
12
#910740000000
0!
0%
b1 *
0-
02
b1 6
#910750000000
1!
1%
1-
12
#910760000000
0!
0%
b10 *
0-
02
b10 6
#910770000000
1!
1%
1-
12
#910780000000
0!
0%
b11 *
0-
02
b11 6
#910790000000
1!
1%
1-
12
15
#910800000000
0!
0%
b100 *
0-
02
b100 6
#910810000000
1!
1%
1-
12
#910820000000
0!
0%
b101 *
0-
02
b101 6
#910830000000
1!
1%
1-
12
#910840000000
0!
0%
b110 *
0-
02
b110 6
#910850000000
1!
1%
1-
12
#910860000000
0!
0%
b111 *
0-
02
b111 6
#910870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#910880000000
0!
0%
b0 *
0-
02
b0 6
#910890000000
1!
1%
1-
12
#910900000000
0!
0%
b1 *
0-
02
b1 6
#910910000000
1!
1%
1-
12
#910920000000
0!
0%
b10 *
0-
02
b10 6
#910930000000
1!
1%
1-
12
#910940000000
0!
0%
b11 *
0-
02
b11 6
#910950000000
1!
1%
1-
12
15
#910960000000
0!
0%
b100 *
0-
02
b100 6
#910970000000
1!
1%
1-
12
#910980000000
0!
0%
b101 *
0-
02
b101 6
#910990000000
1!
1%
1-
12
#911000000000
0!
0%
b110 *
0-
02
b110 6
#911010000000
1!
1%
1-
12
#911020000000
0!
0%
b111 *
0-
02
b111 6
#911030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#911040000000
0!
0%
b0 *
0-
02
b0 6
#911050000000
1!
1%
1-
12
#911060000000
0!
0%
b1 *
0-
02
b1 6
#911070000000
1!
1%
1-
12
#911080000000
0!
0%
b10 *
0-
02
b10 6
#911090000000
1!
1%
1-
12
#911100000000
0!
0%
b11 *
0-
02
b11 6
#911110000000
1!
1%
1-
12
15
#911120000000
0!
0%
b100 *
0-
02
b100 6
#911130000000
1!
1%
1-
12
#911140000000
0!
0%
b101 *
0-
02
b101 6
#911150000000
1!
1%
1-
12
#911160000000
0!
0%
b110 *
0-
02
b110 6
#911170000000
1!
1%
1-
12
#911180000000
0!
0%
b111 *
0-
02
b111 6
#911190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#911200000000
0!
0%
b0 *
0-
02
b0 6
#911210000000
1!
1%
1-
12
#911220000000
0!
0%
b1 *
0-
02
b1 6
#911230000000
1!
1%
1-
12
#911240000000
0!
0%
b10 *
0-
02
b10 6
#911250000000
1!
1%
1-
12
#911260000000
0!
0%
b11 *
0-
02
b11 6
#911270000000
1!
1%
1-
12
15
#911280000000
0!
0%
b100 *
0-
02
b100 6
#911290000000
1!
1%
1-
12
#911300000000
0!
0%
b101 *
0-
02
b101 6
#911310000000
1!
1%
1-
12
#911320000000
0!
0%
b110 *
0-
02
b110 6
#911330000000
1!
1%
1-
12
#911340000000
0!
0%
b111 *
0-
02
b111 6
#911350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#911360000000
0!
0%
b0 *
0-
02
b0 6
#911370000000
1!
1%
1-
12
#911380000000
0!
0%
b1 *
0-
02
b1 6
#911390000000
1!
1%
1-
12
#911400000000
0!
0%
b10 *
0-
02
b10 6
#911410000000
1!
1%
1-
12
#911420000000
0!
0%
b11 *
0-
02
b11 6
#911430000000
1!
1%
1-
12
15
#911440000000
0!
0%
b100 *
0-
02
b100 6
#911450000000
1!
1%
1-
12
#911460000000
0!
0%
b101 *
0-
02
b101 6
#911470000000
1!
1%
1-
12
#911480000000
0!
0%
b110 *
0-
02
b110 6
#911490000000
1!
1%
1-
12
#911500000000
0!
0%
b111 *
0-
02
b111 6
#911510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#911520000000
0!
0%
b0 *
0-
02
b0 6
#911530000000
1!
1%
1-
12
#911540000000
0!
0%
b1 *
0-
02
b1 6
#911550000000
1!
1%
1-
12
#911560000000
0!
0%
b10 *
0-
02
b10 6
#911570000000
1!
1%
1-
12
#911580000000
0!
0%
b11 *
0-
02
b11 6
#911590000000
1!
1%
1-
12
15
#911600000000
0!
0%
b100 *
0-
02
b100 6
#911610000000
1!
1%
1-
12
#911620000000
0!
0%
b101 *
0-
02
b101 6
#911630000000
1!
1%
1-
12
#911640000000
0!
0%
b110 *
0-
02
b110 6
#911650000000
1!
1%
1-
12
#911660000000
0!
0%
b111 *
0-
02
b111 6
#911670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#911680000000
0!
0%
b0 *
0-
02
b0 6
#911690000000
1!
1%
1-
12
#911700000000
0!
0%
b1 *
0-
02
b1 6
#911710000000
1!
1%
1-
12
#911720000000
0!
0%
b10 *
0-
02
b10 6
#911730000000
1!
1%
1-
12
#911740000000
0!
0%
b11 *
0-
02
b11 6
#911750000000
1!
1%
1-
12
15
#911760000000
0!
0%
b100 *
0-
02
b100 6
#911770000000
1!
1%
1-
12
#911780000000
0!
0%
b101 *
0-
02
b101 6
#911790000000
1!
1%
1-
12
#911800000000
0!
0%
b110 *
0-
02
b110 6
#911810000000
1!
1%
1-
12
#911820000000
0!
0%
b111 *
0-
02
b111 6
#911830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#911840000000
0!
0%
b0 *
0-
02
b0 6
#911850000000
1!
1%
1-
12
#911860000000
0!
0%
b1 *
0-
02
b1 6
#911870000000
1!
1%
1-
12
#911880000000
0!
0%
b10 *
0-
02
b10 6
#911890000000
1!
1%
1-
12
#911900000000
0!
0%
b11 *
0-
02
b11 6
#911910000000
1!
1%
1-
12
15
#911920000000
0!
0%
b100 *
0-
02
b100 6
#911930000000
1!
1%
1-
12
#911940000000
0!
0%
b101 *
0-
02
b101 6
#911950000000
1!
1%
1-
12
#911960000000
0!
0%
b110 *
0-
02
b110 6
#911970000000
1!
1%
1-
12
#911980000000
0!
0%
b111 *
0-
02
b111 6
#911990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#912000000000
0!
0%
b0 *
0-
02
b0 6
#912010000000
1!
1%
1-
12
#912020000000
0!
0%
b1 *
0-
02
b1 6
#912030000000
1!
1%
1-
12
#912040000000
0!
0%
b10 *
0-
02
b10 6
#912050000000
1!
1%
1-
12
#912060000000
0!
0%
b11 *
0-
02
b11 6
#912070000000
1!
1%
1-
12
15
#912080000000
0!
0%
b100 *
0-
02
b100 6
#912090000000
1!
1%
1-
12
#912100000000
0!
0%
b101 *
0-
02
b101 6
#912110000000
1!
1%
1-
12
#912120000000
0!
0%
b110 *
0-
02
b110 6
#912130000000
1!
1%
1-
12
#912140000000
0!
0%
b111 *
0-
02
b111 6
#912150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#912160000000
0!
0%
b0 *
0-
02
b0 6
#912170000000
1!
1%
1-
12
#912180000000
0!
0%
b1 *
0-
02
b1 6
#912190000000
1!
1%
1-
12
#912200000000
0!
0%
b10 *
0-
02
b10 6
#912210000000
1!
1%
1-
12
#912220000000
0!
0%
b11 *
0-
02
b11 6
#912230000000
1!
1%
1-
12
15
#912240000000
0!
0%
b100 *
0-
02
b100 6
#912250000000
1!
1%
1-
12
#912260000000
0!
0%
b101 *
0-
02
b101 6
#912270000000
1!
1%
1-
12
#912280000000
0!
0%
b110 *
0-
02
b110 6
#912290000000
1!
1%
1-
12
#912300000000
0!
0%
b111 *
0-
02
b111 6
#912310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#912320000000
0!
0%
b0 *
0-
02
b0 6
#912330000000
1!
1%
1-
12
#912340000000
0!
0%
b1 *
0-
02
b1 6
#912350000000
1!
1%
1-
12
#912360000000
0!
0%
b10 *
0-
02
b10 6
#912370000000
1!
1%
1-
12
#912380000000
0!
0%
b11 *
0-
02
b11 6
#912390000000
1!
1%
1-
12
15
#912400000000
0!
0%
b100 *
0-
02
b100 6
#912410000000
1!
1%
1-
12
#912420000000
0!
0%
b101 *
0-
02
b101 6
#912430000000
1!
1%
1-
12
#912440000000
0!
0%
b110 *
0-
02
b110 6
#912450000000
1!
1%
1-
12
#912460000000
0!
0%
b111 *
0-
02
b111 6
#912470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#912480000000
0!
0%
b0 *
0-
02
b0 6
#912490000000
1!
1%
1-
12
#912500000000
0!
0%
b1 *
0-
02
b1 6
#912510000000
1!
1%
1-
12
#912520000000
0!
0%
b10 *
0-
02
b10 6
#912530000000
1!
1%
1-
12
#912540000000
0!
0%
b11 *
0-
02
b11 6
#912550000000
1!
1%
1-
12
15
#912560000000
0!
0%
b100 *
0-
02
b100 6
#912570000000
1!
1%
1-
12
#912580000000
0!
0%
b101 *
0-
02
b101 6
#912590000000
1!
1%
1-
12
#912600000000
0!
0%
b110 *
0-
02
b110 6
#912610000000
1!
1%
1-
12
#912620000000
0!
0%
b111 *
0-
02
b111 6
#912630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#912640000000
0!
0%
b0 *
0-
02
b0 6
#912650000000
1!
1%
1-
12
#912660000000
0!
0%
b1 *
0-
02
b1 6
#912670000000
1!
1%
1-
12
#912680000000
0!
0%
b10 *
0-
02
b10 6
#912690000000
1!
1%
1-
12
#912700000000
0!
0%
b11 *
0-
02
b11 6
#912710000000
1!
1%
1-
12
15
#912720000000
0!
0%
b100 *
0-
02
b100 6
#912730000000
1!
1%
1-
12
#912740000000
0!
0%
b101 *
0-
02
b101 6
#912750000000
1!
1%
1-
12
#912760000000
0!
0%
b110 *
0-
02
b110 6
#912770000000
1!
1%
1-
12
#912780000000
0!
0%
b111 *
0-
02
b111 6
#912790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#912800000000
0!
0%
b0 *
0-
02
b0 6
#912810000000
1!
1%
1-
12
#912820000000
0!
0%
b1 *
0-
02
b1 6
#912830000000
1!
1%
1-
12
#912840000000
0!
0%
b10 *
0-
02
b10 6
#912850000000
1!
1%
1-
12
#912860000000
0!
0%
b11 *
0-
02
b11 6
#912870000000
1!
1%
1-
12
15
#912880000000
0!
0%
b100 *
0-
02
b100 6
#912890000000
1!
1%
1-
12
#912900000000
0!
0%
b101 *
0-
02
b101 6
#912910000000
1!
1%
1-
12
#912920000000
0!
0%
b110 *
0-
02
b110 6
#912930000000
1!
1%
1-
12
#912940000000
0!
0%
b111 *
0-
02
b111 6
#912950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#912960000000
0!
0%
b0 *
0-
02
b0 6
#912970000000
1!
1%
1-
12
#912980000000
0!
0%
b1 *
0-
02
b1 6
#912990000000
1!
1%
1-
12
#913000000000
0!
0%
b10 *
0-
02
b10 6
#913010000000
1!
1%
1-
12
#913020000000
0!
0%
b11 *
0-
02
b11 6
#913030000000
1!
1%
1-
12
15
#913040000000
0!
0%
b100 *
0-
02
b100 6
#913050000000
1!
1%
1-
12
#913060000000
0!
0%
b101 *
0-
02
b101 6
#913070000000
1!
1%
1-
12
#913080000000
0!
0%
b110 *
0-
02
b110 6
#913090000000
1!
1%
1-
12
#913100000000
0!
0%
b111 *
0-
02
b111 6
#913110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#913120000000
0!
0%
b0 *
0-
02
b0 6
#913130000000
1!
1%
1-
12
#913140000000
0!
0%
b1 *
0-
02
b1 6
#913150000000
1!
1%
1-
12
#913160000000
0!
0%
b10 *
0-
02
b10 6
#913170000000
1!
1%
1-
12
#913180000000
0!
0%
b11 *
0-
02
b11 6
#913190000000
1!
1%
1-
12
15
#913200000000
0!
0%
b100 *
0-
02
b100 6
#913210000000
1!
1%
1-
12
#913220000000
0!
0%
b101 *
0-
02
b101 6
#913230000000
1!
1%
1-
12
#913240000000
0!
0%
b110 *
0-
02
b110 6
#913250000000
1!
1%
1-
12
#913260000000
0!
0%
b111 *
0-
02
b111 6
#913270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#913280000000
0!
0%
b0 *
0-
02
b0 6
#913290000000
1!
1%
1-
12
#913300000000
0!
0%
b1 *
0-
02
b1 6
#913310000000
1!
1%
1-
12
#913320000000
0!
0%
b10 *
0-
02
b10 6
#913330000000
1!
1%
1-
12
#913340000000
0!
0%
b11 *
0-
02
b11 6
#913350000000
1!
1%
1-
12
15
#913360000000
0!
0%
b100 *
0-
02
b100 6
#913370000000
1!
1%
1-
12
#913380000000
0!
0%
b101 *
0-
02
b101 6
#913390000000
1!
1%
1-
12
#913400000000
0!
0%
b110 *
0-
02
b110 6
#913410000000
1!
1%
1-
12
#913420000000
0!
0%
b111 *
0-
02
b111 6
#913430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#913440000000
0!
0%
b0 *
0-
02
b0 6
#913450000000
1!
1%
1-
12
#913460000000
0!
0%
b1 *
0-
02
b1 6
#913470000000
1!
1%
1-
12
#913480000000
0!
0%
b10 *
0-
02
b10 6
#913490000000
1!
1%
1-
12
#913500000000
0!
0%
b11 *
0-
02
b11 6
#913510000000
1!
1%
1-
12
15
#913520000000
0!
0%
b100 *
0-
02
b100 6
#913530000000
1!
1%
1-
12
#913540000000
0!
0%
b101 *
0-
02
b101 6
#913550000000
1!
1%
1-
12
#913560000000
0!
0%
b110 *
0-
02
b110 6
#913570000000
1!
1%
1-
12
#913580000000
0!
0%
b111 *
0-
02
b111 6
#913590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#913600000000
0!
0%
b0 *
0-
02
b0 6
#913610000000
1!
1%
1-
12
#913620000000
0!
0%
b1 *
0-
02
b1 6
#913630000000
1!
1%
1-
12
#913640000000
0!
0%
b10 *
0-
02
b10 6
#913650000000
1!
1%
1-
12
#913660000000
0!
0%
b11 *
0-
02
b11 6
#913670000000
1!
1%
1-
12
15
#913680000000
0!
0%
b100 *
0-
02
b100 6
#913690000000
1!
1%
1-
12
#913700000000
0!
0%
b101 *
0-
02
b101 6
#913710000000
1!
1%
1-
12
#913720000000
0!
0%
b110 *
0-
02
b110 6
#913730000000
1!
1%
1-
12
#913740000000
0!
0%
b111 *
0-
02
b111 6
#913750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#913760000000
0!
0%
b0 *
0-
02
b0 6
#913770000000
1!
1%
1-
12
#913780000000
0!
0%
b1 *
0-
02
b1 6
#913790000000
1!
1%
1-
12
#913800000000
0!
0%
b10 *
0-
02
b10 6
#913810000000
1!
1%
1-
12
#913820000000
0!
0%
b11 *
0-
02
b11 6
#913830000000
1!
1%
1-
12
15
#913840000000
0!
0%
b100 *
0-
02
b100 6
#913850000000
1!
1%
1-
12
#913860000000
0!
0%
b101 *
0-
02
b101 6
#913870000000
1!
1%
1-
12
#913880000000
0!
0%
b110 *
0-
02
b110 6
#913890000000
1!
1%
1-
12
#913900000000
0!
0%
b111 *
0-
02
b111 6
#913910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#913920000000
0!
0%
b0 *
0-
02
b0 6
#913930000000
1!
1%
1-
12
#913940000000
0!
0%
b1 *
0-
02
b1 6
#913950000000
1!
1%
1-
12
#913960000000
0!
0%
b10 *
0-
02
b10 6
#913970000000
1!
1%
1-
12
#913980000000
0!
0%
b11 *
0-
02
b11 6
#913990000000
1!
1%
1-
12
15
#914000000000
0!
0%
b100 *
0-
02
b100 6
#914010000000
1!
1%
1-
12
#914020000000
0!
0%
b101 *
0-
02
b101 6
#914030000000
1!
1%
1-
12
#914040000000
0!
0%
b110 *
0-
02
b110 6
#914050000000
1!
1%
1-
12
#914060000000
0!
0%
b111 *
0-
02
b111 6
#914070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#914080000000
0!
0%
b0 *
0-
02
b0 6
#914090000000
1!
1%
1-
12
#914100000000
0!
0%
b1 *
0-
02
b1 6
#914110000000
1!
1%
1-
12
#914120000000
0!
0%
b10 *
0-
02
b10 6
#914130000000
1!
1%
1-
12
#914140000000
0!
0%
b11 *
0-
02
b11 6
#914150000000
1!
1%
1-
12
15
#914160000000
0!
0%
b100 *
0-
02
b100 6
#914170000000
1!
1%
1-
12
#914180000000
0!
0%
b101 *
0-
02
b101 6
#914190000000
1!
1%
1-
12
#914200000000
0!
0%
b110 *
0-
02
b110 6
#914210000000
1!
1%
1-
12
#914220000000
0!
0%
b111 *
0-
02
b111 6
#914230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#914240000000
0!
0%
b0 *
0-
02
b0 6
#914250000000
1!
1%
1-
12
#914260000000
0!
0%
b1 *
0-
02
b1 6
#914270000000
1!
1%
1-
12
#914280000000
0!
0%
b10 *
0-
02
b10 6
#914290000000
1!
1%
1-
12
#914300000000
0!
0%
b11 *
0-
02
b11 6
#914310000000
1!
1%
1-
12
15
#914320000000
0!
0%
b100 *
0-
02
b100 6
#914330000000
1!
1%
1-
12
#914340000000
0!
0%
b101 *
0-
02
b101 6
#914350000000
1!
1%
1-
12
#914360000000
0!
0%
b110 *
0-
02
b110 6
#914370000000
1!
1%
1-
12
#914380000000
0!
0%
b111 *
0-
02
b111 6
#914390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#914400000000
0!
0%
b0 *
0-
02
b0 6
#914410000000
1!
1%
1-
12
#914420000000
0!
0%
b1 *
0-
02
b1 6
#914430000000
1!
1%
1-
12
#914440000000
0!
0%
b10 *
0-
02
b10 6
#914450000000
1!
1%
1-
12
#914460000000
0!
0%
b11 *
0-
02
b11 6
#914470000000
1!
1%
1-
12
15
#914480000000
0!
0%
b100 *
0-
02
b100 6
#914490000000
1!
1%
1-
12
#914500000000
0!
0%
b101 *
0-
02
b101 6
#914510000000
1!
1%
1-
12
#914520000000
0!
0%
b110 *
0-
02
b110 6
#914530000000
1!
1%
1-
12
#914540000000
0!
0%
b111 *
0-
02
b111 6
#914550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#914560000000
0!
0%
b0 *
0-
02
b0 6
#914570000000
1!
1%
1-
12
#914580000000
0!
0%
b1 *
0-
02
b1 6
#914590000000
1!
1%
1-
12
#914600000000
0!
0%
b10 *
0-
02
b10 6
#914610000000
1!
1%
1-
12
#914620000000
0!
0%
b11 *
0-
02
b11 6
#914630000000
1!
1%
1-
12
15
#914640000000
0!
0%
b100 *
0-
02
b100 6
#914650000000
1!
1%
1-
12
#914660000000
0!
0%
b101 *
0-
02
b101 6
#914670000000
1!
1%
1-
12
#914680000000
0!
0%
b110 *
0-
02
b110 6
#914690000000
1!
1%
1-
12
#914700000000
0!
0%
b111 *
0-
02
b111 6
#914710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#914720000000
0!
0%
b0 *
0-
02
b0 6
#914730000000
1!
1%
1-
12
#914740000000
0!
0%
b1 *
0-
02
b1 6
#914750000000
1!
1%
1-
12
#914760000000
0!
0%
b10 *
0-
02
b10 6
#914770000000
1!
1%
1-
12
#914780000000
0!
0%
b11 *
0-
02
b11 6
#914790000000
1!
1%
1-
12
15
#914800000000
0!
0%
b100 *
0-
02
b100 6
#914810000000
1!
1%
1-
12
#914820000000
0!
0%
b101 *
0-
02
b101 6
#914830000000
1!
1%
1-
12
#914840000000
0!
0%
b110 *
0-
02
b110 6
#914850000000
1!
1%
1-
12
#914860000000
0!
0%
b111 *
0-
02
b111 6
#914870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#914880000000
0!
0%
b0 *
0-
02
b0 6
#914890000000
1!
1%
1-
12
#914900000000
0!
0%
b1 *
0-
02
b1 6
#914910000000
1!
1%
1-
12
#914920000000
0!
0%
b10 *
0-
02
b10 6
#914930000000
1!
1%
1-
12
#914940000000
0!
0%
b11 *
0-
02
b11 6
#914950000000
1!
1%
1-
12
15
#914960000000
0!
0%
b100 *
0-
02
b100 6
#914970000000
1!
1%
1-
12
#914980000000
0!
0%
b101 *
0-
02
b101 6
#914990000000
1!
1%
1-
12
#915000000000
0!
0%
b110 *
0-
02
b110 6
#915010000000
1!
1%
1-
12
#915020000000
0!
0%
b111 *
0-
02
b111 6
#915030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#915040000000
0!
0%
b0 *
0-
02
b0 6
#915050000000
1!
1%
1-
12
#915060000000
0!
0%
b1 *
0-
02
b1 6
#915070000000
1!
1%
1-
12
#915080000000
0!
0%
b10 *
0-
02
b10 6
#915090000000
1!
1%
1-
12
#915100000000
0!
0%
b11 *
0-
02
b11 6
#915110000000
1!
1%
1-
12
15
#915120000000
0!
0%
b100 *
0-
02
b100 6
#915130000000
1!
1%
1-
12
#915140000000
0!
0%
b101 *
0-
02
b101 6
#915150000000
1!
1%
1-
12
#915160000000
0!
0%
b110 *
0-
02
b110 6
#915170000000
1!
1%
1-
12
#915180000000
0!
0%
b111 *
0-
02
b111 6
#915190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#915200000000
0!
0%
b0 *
0-
02
b0 6
#915210000000
1!
1%
1-
12
#915220000000
0!
0%
b1 *
0-
02
b1 6
#915230000000
1!
1%
1-
12
#915240000000
0!
0%
b10 *
0-
02
b10 6
#915250000000
1!
1%
1-
12
#915260000000
0!
0%
b11 *
0-
02
b11 6
#915270000000
1!
1%
1-
12
15
#915280000000
0!
0%
b100 *
0-
02
b100 6
#915290000000
1!
1%
1-
12
#915300000000
0!
0%
b101 *
0-
02
b101 6
#915310000000
1!
1%
1-
12
#915320000000
0!
0%
b110 *
0-
02
b110 6
#915330000000
1!
1%
1-
12
#915340000000
0!
0%
b111 *
0-
02
b111 6
#915350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#915360000000
0!
0%
b0 *
0-
02
b0 6
#915370000000
1!
1%
1-
12
#915380000000
0!
0%
b1 *
0-
02
b1 6
#915390000000
1!
1%
1-
12
#915400000000
0!
0%
b10 *
0-
02
b10 6
#915410000000
1!
1%
1-
12
#915420000000
0!
0%
b11 *
0-
02
b11 6
#915430000000
1!
1%
1-
12
15
#915440000000
0!
0%
b100 *
0-
02
b100 6
#915450000000
1!
1%
1-
12
#915460000000
0!
0%
b101 *
0-
02
b101 6
#915470000000
1!
1%
1-
12
#915480000000
0!
0%
b110 *
0-
02
b110 6
#915490000000
1!
1%
1-
12
#915500000000
0!
0%
b111 *
0-
02
b111 6
#915510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#915520000000
0!
0%
b0 *
0-
02
b0 6
#915530000000
1!
1%
1-
12
#915540000000
0!
0%
b1 *
0-
02
b1 6
#915550000000
1!
1%
1-
12
#915560000000
0!
0%
b10 *
0-
02
b10 6
#915570000000
1!
1%
1-
12
#915580000000
0!
0%
b11 *
0-
02
b11 6
#915590000000
1!
1%
1-
12
15
#915600000000
0!
0%
b100 *
0-
02
b100 6
#915610000000
1!
1%
1-
12
#915620000000
0!
0%
b101 *
0-
02
b101 6
#915630000000
1!
1%
1-
12
#915640000000
0!
0%
b110 *
0-
02
b110 6
#915650000000
1!
1%
1-
12
#915660000000
0!
0%
b111 *
0-
02
b111 6
#915670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#915680000000
0!
0%
b0 *
0-
02
b0 6
#915690000000
1!
1%
1-
12
#915700000000
0!
0%
b1 *
0-
02
b1 6
#915710000000
1!
1%
1-
12
#915720000000
0!
0%
b10 *
0-
02
b10 6
#915730000000
1!
1%
1-
12
#915740000000
0!
0%
b11 *
0-
02
b11 6
#915750000000
1!
1%
1-
12
15
#915760000000
0!
0%
b100 *
0-
02
b100 6
#915770000000
1!
1%
1-
12
#915780000000
0!
0%
b101 *
0-
02
b101 6
#915790000000
1!
1%
1-
12
#915800000000
0!
0%
b110 *
0-
02
b110 6
#915810000000
1!
1%
1-
12
#915820000000
0!
0%
b111 *
0-
02
b111 6
#915830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#915840000000
0!
0%
b0 *
0-
02
b0 6
#915850000000
1!
1%
1-
12
#915860000000
0!
0%
b1 *
0-
02
b1 6
#915870000000
1!
1%
1-
12
#915880000000
0!
0%
b10 *
0-
02
b10 6
#915890000000
1!
1%
1-
12
#915900000000
0!
0%
b11 *
0-
02
b11 6
#915910000000
1!
1%
1-
12
15
#915920000000
0!
0%
b100 *
0-
02
b100 6
#915930000000
1!
1%
1-
12
#915940000000
0!
0%
b101 *
0-
02
b101 6
#915950000000
1!
1%
1-
12
#915960000000
0!
0%
b110 *
0-
02
b110 6
#915970000000
1!
1%
1-
12
#915980000000
0!
0%
b111 *
0-
02
b111 6
#915990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#916000000000
0!
0%
b0 *
0-
02
b0 6
#916010000000
1!
1%
1-
12
#916020000000
0!
0%
b1 *
0-
02
b1 6
#916030000000
1!
1%
1-
12
#916040000000
0!
0%
b10 *
0-
02
b10 6
#916050000000
1!
1%
1-
12
#916060000000
0!
0%
b11 *
0-
02
b11 6
#916070000000
1!
1%
1-
12
15
#916080000000
0!
0%
b100 *
0-
02
b100 6
#916090000000
1!
1%
1-
12
#916100000000
0!
0%
b101 *
0-
02
b101 6
#916110000000
1!
1%
1-
12
#916120000000
0!
0%
b110 *
0-
02
b110 6
#916130000000
1!
1%
1-
12
#916140000000
0!
0%
b111 *
0-
02
b111 6
#916150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#916160000000
0!
0%
b0 *
0-
02
b0 6
#916170000000
1!
1%
1-
12
#916180000000
0!
0%
b1 *
0-
02
b1 6
#916190000000
1!
1%
1-
12
#916200000000
0!
0%
b10 *
0-
02
b10 6
#916210000000
1!
1%
1-
12
#916220000000
0!
0%
b11 *
0-
02
b11 6
#916230000000
1!
1%
1-
12
15
#916240000000
0!
0%
b100 *
0-
02
b100 6
#916250000000
1!
1%
1-
12
#916260000000
0!
0%
b101 *
0-
02
b101 6
#916270000000
1!
1%
1-
12
#916280000000
0!
0%
b110 *
0-
02
b110 6
#916290000000
1!
1%
1-
12
#916300000000
0!
0%
b111 *
0-
02
b111 6
#916310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#916320000000
0!
0%
b0 *
0-
02
b0 6
#916330000000
1!
1%
1-
12
#916340000000
0!
0%
b1 *
0-
02
b1 6
#916350000000
1!
1%
1-
12
#916360000000
0!
0%
b10 *
0-
02
b10 6
#916370000000
1!
1%
1-
12
#916380000000
0!
0%
b11 *
0-
02
b11 6
#916390000000
1!
1%
1-
12
15
#916400000000
0!
0%
b100 *
0-
02
b100 6
#916410000000
1!
1%
1-
12
#916420000000
0!
0%
b101 *
0-
02
b101 6
#916430000000
1!
1%
1-
12
#916440000000
0!
0%
b110 *
0-
02
b110 6
#916450000000
1!
1%
1-
12
#916460000000
0!
0%
b111 *
0-
02
b111 6
#916470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#916480000000
0!
0%
b0 *
0-
02
b0 6
#916490000000
1!
1%
1-
12
#916500000000
0!
0%
b1 *
0-
02
b1 6
#916510000000
1!
1%
1-
12
#916520000000
0!
0%
b10 *
0-
02
b10 6
#916530000000
1!
1%
1-
12
#916540000000
0!
0%
b11 *
0-
02
b11 6
#916550000000
1!
1%
1-
12
15
#916560000000
0!
0%
b100 *
0-
02
b100 6
#916570000000
1!
1%
1-
12
#916580000000
0!
0%
b101 *
0-
02
b101 6
#916590000000
1!
1%
1-
12
#916600000000
0!
0%
b110 *
0-
02
b110 6
#916610000000
1!
1%
1-
12
#916620000000
0!
0%
b111 *
0-
02
b111 6
#916630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#916640000000
0!
0%
b0 *
0-
02
b0 6
#916650000000
1!
1%
1-
12
#916660000000
0!
0%
b1 *
0-
02
b1 6
#916670000000
1!
1%
1-
12
#916680000000
0!
0%
b10 *
0-
02
b10 6
#916690000000
1!
1%
1-
12
#916700000000
0!
0%
b11 *
0-
02
b11 6
#916710000000
1!
1%
1-
12
15
#916720000000
0!
0%
b100 *
0-
02
b100 6
#916730000000
1!
1%
1-
12
#916740000000
0!
0%
b101 *
0-
02
b101 6
#916750000000
1!
1%
1-
12
#916760000000
0!
0%
b110 *
0-
02
b110 6
#916770000000
1!
1%
1-
12
#916780000000
0!
0%
b111 *
0-
02
b111 6
#916790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#916800000000
0!
0%
b0 *
0-
02
b0 6
#916810000000
1!
1%
1-
12
#916820000000
0!
0%
b1 *
0-
02
b1 6
#916830000000
1!
1%
1-
12
#916840000000
0!
0%
b10 *
0-
02
b10 6
#916850000000
1!
1%
1-
12
#916860000000
0!
0%
b11 *
0-
02
b11 6
#916870000000
1!
1%
1-
12
15
#916880000000
0!
0%
b100 *
0-
02
b100 6
#916890000000
1!
1%
1-
12
#916900000000
0!
0%
b101 *
0-
02
b101 6
#916910000000
1!
1%
1-
12
#916920000000
0!
0%
b110 *
0-
02
b110 6
#916930000000
1!
1%
1-
12
#916940000000
0!
0%
b111 *
0-
02
b111 6
#916950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#916960000000
0!
0%
b0 *
0-
02
b0 6
#916970000000
1!
1%
1-
12
#916980000000
0!
0%
b1 *
0-
02
b1 6
#916990000000
1!
1%
1-
12
#917000000000
0!
0%
b10 *
0-
02
b10 6
#917010000000
1!
1%
1-
12
#917020000000
0!
0%
b11 *
0-
02
b11 6
#917030000000
1!
1%
1-
12
15
#917040000000
0!
0%
b100 *
0-
02
b100 6
#917050000000
1!
1%
1-
12
#917060000000
0!
0%
b101 *
0-
02
b101 6
#917070000000
1!
1%
1-
12
#917080000000
0!
0%
b110 *
0-
02
b110 6
#917090000000
1!
1%
1-
12
#917100000000
0!
0%
b111 *
0-
02
b111 6
#917110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#917120000000
0!
0%
b0 *
0-
02
b0 6
#917130000000
1!
1%
1-
12
#917140000000
0!
0%
b1 *
0-
02
b1 6
#917150000000
1!
1%
1-
12
#917160000000
0!
0%
b10 *
0-
02
b10 6
#917170000000
1!
1%
1-
12
#917180000000
0!
0%
b11 *
0-
02
b11 6
#917190000000
1!
1%
1-
12
15
#917200000000
0!
0%
b100 *
0-
02
b100 6
#917210000000
1!
1%
1-
12
#917220000000
0!
0%
b101 *
0-
02
b101 6
#917230000000
1!
1%
1-
12
#917240000000
0!
0%
b110 *
0-
02
b110 6
#917250000000
1!
1%
1-
12
#917260000000
0!
0%
b111 *
0-
02
b111 6
#917270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#917280000000
0!
0%
b0 *
0-
02
b0 6
#917290000000
1!
1%
1-
12
#917300000000
0!
0%
b1 *
0-
02
b1 6
#917310000000
1!
1%
1-
12
#917320000000
0!
0%
b10 *
0-
02
b10 6
#917330000000
1!
1%
1-
12
#917340000000
0!
0%
b11 *
0-
02
b11 6
#917350000000
1!
1%
1-
12
15
#917360000000
0!
0%
b100 *
0-
02
b100 6
#917370000000
1!
1%
1-
12
#917380000000
0!
0%
b101 *
0-
02
b101 6
#917390000000
1!
1%
1-
12
#917400000000
0!
0%
b110 *
0-
02
b110 6
#917410000000
1!
1%
1-
12
#917420000000
0!
0%
b111 *
0-
02
b111 6
#917430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#917440000000
0!
0%
b0 *
0-
02
b0 6
#917450000000
1!
1%
1-
12
#917460000000
0!
0%
b1 *
0-
02
b1 6
#917470000000
1!
1%
1-
12
#917480000000
0!
0%
b10 *
0-
02
b10 6
#917490000000
1!
1%
1-
12
#917500000000
0!
0%
b11 *
0-
02
b11 6
#917510000000
1!
1%
1-
12
15
#917520000000
0!
0%
b100 *
0-
02
b100 6
#917530000000
1!
1%
1-
12
#917540000000
0!
0%
b101 *
0-
02
b101 6
#917550000000
1!
1%
1-
12
#917560000000
0!
0%
b110 *
0-
02
b110 6
#917570000000
1!
1%
1-
12
#917580000000
0!
0%
b111 *
0-
02
b111 6
#917590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#917600000000
0!
0%
b0 *
0-
02
b0 6
#917610000000
1!
1%
1-
12
#917620000000
0!
0%
b1 *
0-
02
b1 6
#917630000000
1!
1%
1-
12
#917640000000
0!
0%
b10 *
0-
02
b10 6
#917650000000
1!
1%
1-
12
#917660000000
0!
0%
b11 *
0-
02
b11 6
#917670000000
1!
1%
1-
12
15
#917680000000
0!
0%
b100 *
0-
02
b100 6
#917690000000
1!
1%
1-
12
#917700000000
0!
0%
b101 *
0-
02
b101 6
#917710000000
1!
1%
1-
12
#917720000000
0!
0%
b110 *
0-
02
b110 6
#917730000000
1!
1%
1-
12
#917740000000
0!
0%
b111 *
0-
02
b111 6
#917750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#917760000000
0!
0%
b0 *
0-
02
b0 6
#917770000000
1!
1%
1-
12
#917780000000
0!
0%
b1 *
0-
02
b1 6
#917790000000
1!
1%
1-
12
#917800000000
0!
0%
b10 *
0-
02
b10 6
#917810000000
1!
1%
1-
12
#917820000000
0!
0%
b11 *
0-
02
b11 6
#917830000000
1!
1%
1-
12
15
#917840000000
0!
0%
b100 *
0-
02
b100 6
#917850000000
1!
1%
1-
12
#917860000000
0!
0%
b101 *
0-
02
b101 6
#917870000000
1!
1%
1-
12
#917880000000
0!
0%
b110 *
0-
02
b110 6
#917890000000
1!
1%
1-
12
#917900000000
0!
0%
b111 *
0-
02
b111 6
#917910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#917920000000
0!
0%
b0 *
0-
02
b0 6
#917930000000
1!
1%
1-
12
#917940000000
0!
0%
b1 *
0-
02
b1 6
#917950000000
1!
1%
1-
12
#917960000000
0!
0%
b10 *
0-
02
b10 6
#917970000000
1!
1%
1-
12
#917980000000
0!
0%
b11 *
0-
02
b11 6
#917990000000
1!
1%
1-
12
15
#918000000000
0!
0%
b100 *
0-
02
b100 6
#918010000000
1!
1%
1-
12
#918020000000
0!
0%
b101 *
0-
02
b101 6
#918030000000
1!
1%
1-
12
#918040000000
0!
0%
b110 *
0-
02
b110 6
#918050000000
1!
1%
1-
12
#918060000000
0!
0%
b111 *
0-
02
b111 6
#918070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#918080000000
0!
0%
b0 *
0-
02
b0 6
#918090000000
1!
1%
1-
12
#918100000000
0!
0%
b1 *
0-
02
b1 6
#918110000000
1!
1%
1-
12
#918120000000
0!
0%
b10 *
0-
02
b10 6
#918130000000
1!
1%
1-
12
#918140000000
0!
0%
b11 *
0-
02
b11 6
#918150000000
1!
1%
1-
12
15
#918160000000
0!
0%
b100 *
0-
02
b100 6
#918170000000
1!
1%
1-
12
#918180000000
0!
0%
b101 *
0-
02
b101 6
#918190000000
1!
1%
1-
12
#918200000000
0!
0%
b110 *
0-
02
b110 6
#918210000000
1!
1%
1-
12
#918220000000
0!
0%
b111 *
0-
02
b111 6
#918230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#918240000000
0!
0%
b0 *
0-
02
b0 6
#918250000000
1!
1%
1-
12
#918260000000
0!
0%
b1 *
0-
02
b1 6
#918270000000
1!
1%
1-
12
#918280000000
0!
0%
b10 *
0-
02
b10 6
#918290000000
1!
1%
1-
12
#918300000000
0!
0%
b11 *
0-
02
b11 6
#918310000000
1!
1%
1-
12
15
#918320000000
0!
0%
b100 *
0-
02
b100 6
#918330000000
1!
1%
1-
12
#918340000000
0!
0%
b101 *
0-
02
b101 6
#918350000000
1!
1%
1-
12
#918360000000
0!
0%
b110 *
0-
02
b110 6
#918370000000
1!
1%
1-
12
#918380000000
0!
0%
b111 *
0-
02
b111 6
#918390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#918400000000
0!
0%
b0 *
0-
02
b0 6
#918410000000
1!
1%
1-
12
#918420000000
0!
0%
b1 *
0-
02
b1 6
#918430000000
1!
1%
1-
12
#918440000000
0!
0%
b10 *
0-
02
b10 6
#918450000000
1!
1%
1-
12
#918460000000
0!
0%
b11 *
0-
02
b11 6
#918470000000
1!
1%
1-
12
15
#918480000000
0!
0%
b100 *
0-
02
b100 6
#918490000000
1!
1%
1-
12
#918500000000
0!
0%
b101 *
0-
02
b101 6
#918510000000
1!
1%
1-
12
#918520000000
0!
0%
b110 *
0-
02
b110 6
#918530000000
1!
1%
1-
12
#918540000000
0!
0%
b111 *
0-
02
b111 6
#918550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#918560000000
0!
0%
b0 *
0-
02
b0 6
#918570000000
1!
1%
1-
12
#918580000000
0!
0%
b1 *
0-
02
b1 6
#918590000000
1!
1%
1-
12
#918600000000
0!
0%
b10 *
0-
02
b10 6
#918610000000
1!
1%
1-
12
#918620000000
0!
0%
b11 *
0-
02
b11 6
#918630000000
1!
1%
1-
12
15
#918640000000
0!
0%
b100 *
0-
02
b100 6
#918650000000
1!
1%
1-
12
#918660000000
0!
0%
b101 *
0-
02
b101 6
#918670000000
1!
1%
1-
12
#918680000000
0!
0%
b110 *
0-
02
b110 6
#918690000000
1!
1%
1-
12
#918700000000
0!
0%
b111 *
0-
02
b111 6
#918710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#918720000000
0!
0%
b0 *
0-
02
b0 6
#918730000000
1!
1%
1-
12
#918740000000
0!
0%
b1 *
0-
02
b1 6
#918750000000
1!
1%
1-
12
#918760000000
0!
0%
b10 *
0-
02
b10 6
#918770000000
1!
1%
1-
12
#918780000000
0!
0%
b11 *
0-
02
b11 6
#918790000000
1!
1%
1-
12
15
#918800000000
0!
0%
b100 *
0-
02
b100 6
#918810000000
1!
1%
1-
12
#918820000000
0!
0%
b101 *
0-
02
b101 6
#918830000000
1!
1%
1-
12
#918840000000
0!
0%
b110 *
0-
02
b110 6
#918850000000
1!
1%
1-
12
#918860000000
0!
0%
b111 *
0-
02
b111 6
#918870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#918880000000
0!
0%
b0 *
0-
02
b0 6
#918890000000
1!
1%
1-
12
#918900000000
0!
0%
b1 *
0-
02
b1 6
#918910000000
1!
1%
1-
12
#918920000000
0!
0%
b10 *
0-
02
b10 6
#918930000000
1!
1%
1-
12
#918940000000
0!
0%
b11 *
0-
02
b11 6
#918950000000
1!
1%
1-
12
15
#918960000000
0!
0%
b100 *
0-
02
b100 6
#918970000000
1!
1%
1-
12
#918980000000
0!
0%
b101 *
0-
02
b101 6
#918990000000
1!
1%
1-
12
#919000000000
0!
0%
b110 *
0-
02
b110 6
#919010000000
1!
1%
1-
12
#919020000000
0!
0%
b111 *
0-
02
b111 6
#919030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#919040000000
0!
0%
b0 *
0-
02
b0 6
#919050000000
1!
1%
1-
12
#919060000000
0!
0%
b1 *
0-
02
b1 6
#919070000000
1!
1%
1-
12
#919080000000
0!
0%
b10 *
0-
02
b10 6
#919090000000
1!
1%
1-
12
#919100000000
0!
0%
b11 *
0-
02
b11 6
#919110000000
1!
1%
1-
12
15
#919120000000
0!
0%
b100 *
0-
02
b100 6
#919130000000
1!
1%
1-
12
#919140000000
0!
0%
b101 *
0-
02
b101 6
#919150000000
1!
1%
1-
12
#919160000000
0!
0%
b110 *
0-
02
b110 6
#919170000000
1!
1%
1-
12
#919180000000
0!
0%
b111 *
0-
02
b111 6
#919190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#919200000000
0!
0%
b0 *
0-
02
b0 6
#919210000000
1!
1%
1-
12
#919220000000
0!
0%
b1 *
0-
02
b1 6
#919230000000
1!
1%
1-
12
#919240000000
0!
0%
b10 *
0-
02
b10 6
#919250000000
1!
1%
1-
12
#919260000000
0!
0%
b11 *
0-
02
b11 6
#919270000000
1!
1%
1-
12
15
#919280000000
0!
0%
b100 *
0-
02
b100 6
#919290000000
1!
1%
1-
12
#919300000000
0!
0%
b101 *
0-
02
b101 6
#919310000000
1!
1%
1-
12
#919320000000
0!
0%
b110 *
0-
02
b110 6
#919330000000
1!
1%
1-
12
#919340000000
0!
0%
b111 *
0-
02
b111 6
#919350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#919360000000
0!
0%
b0 *
0-
02
b0 6
#919370000000
1!
1%
1-
12
#919380000000
0!
0%
b1 *
0-
02
b1 6
#919390000000
1!
1%
1-
12
#919400000000
0!
0%
b10 *
0-
02
b10 6
#919410000000
1!
1%
1-
12
#919420000000
0!
0%
b11 *
0-
02
b11 6
#919430000000
1!
1%
1-
12
15
#919440000000
0!
0%
b100 *
0-
02
b100 6
#919450000000
1!
1%
1-
12
#919460000000
0!
0%
b101 *
0-
02
b101 6
#919470000000
1!
1%
1-
12
#919480000000
0!
0%
b110 *
0-
02
b110 6
#919490000000
1!
1%
1-
12
#919500000000
0!
0%
b111 *
0-
02
b111 6
#919510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#919520000000
0!
0%
b0 *
0-
02
b0 6
#919530000000
1!
1%
1-
12
#919540000000
0!
0%
b1 *
0-
02
b1 6
#919550000000
1!
1%
1-
12
#919560000000
0!
0%
b10 *
0-
02
b10 6
#919570000000
1!
1%
1-
12
#919580000000
0!
0%
b11 *
0-
02
b11 6
#919590000000
1!
1%
1-
12
15
#919600000000
0!
0%
b100 *
0-
02
b100 6
#919610000000
1!
1%
1-
12
#919620000000
0!
0%
b101 *
0-
02
b101 6
#919630000000
1!
1%
1-
12
#919640000000
0!
0%
b110 *
0-
02
b110 6
#919650000000
1!
1%
1-
12
#919660000000
0!
0%
b111 *
0-
02
b111 6
#919670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#919680000000
0!
0%
b0 *
0-
02
b0 6
#919690000000
1!
1%
1-
12
#919700000000
0!
0%
b1 *
0-
02
b1 6
#919710000000
1!
1%
1-
12
#919720000000
0!
0%
b10 *
0-
02
b10 6
#919730000000
1!
1%
1-
12
#919740000000
0!
0%
b11 *
0-
02
b11 6
#919750000000
1!
1%
1-
12
15
#919760000000
0!
0%
b100 *
0-
02
b100 6
#919770000000
1!
1%
1-
12
#919780000000
0!
0%
b101 *
0-
02
b101 6
#919790000000
1!
1%
1-
12
#919800000000
0!
0%
b110 *
0-
02
b110 6
#919810000000
1!
1%
1-
12
#919820000000
0!
0%
b111 *
0-
02
b111 6
#919830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#919840000000
0!
0%
b0 *
0-
02
b0 6
#919850000000
1!
1%
1-
12
#919860000000
0!
0%
b1 *
0-
02
b1 6
#919870000000
1!
1%
1-
12
#919880000000
0!
0%
b10 *
0-
02
b10 6
#919890000000
1!
1%
1-
12
#919900000000
0!
0%
b11 *
0-
02
b11 6
#919910000000
1!
1%
1-
12
15
#919920000000
0!
0%
b100 *
0-
02
b100 6
#919930000000
1!
1%
1-
12
#919940000000
0!
0%
b101 *
0-
02
b101 6
#919950000000
1!
1%
1-
12
#919960000000
0!
0%
b110 *
0-
02
b110 6
#919970000000
1!
1%
1-
12
#919980000000
0!
0%
b111 *
0-
02
b111 6
#919990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#920000000000
0!
0%
b0 *
0-
02
b0 6
#920010000000
1!
1%
1-
12
#920020000000
0!
0%
b1 *
0-
02
b1 6
#920030000000
1!
1%
1-
12
#920040000000
0!
0%
b10 *
0-
02
b10 6
#920050000000
1!
1%
1-
12
#920060000000
0!
0%
b11 *
0-
02
b11 6
#920070000000
1!
1%
1-
12
15
#920080000000
0!
0%
b100 *
0-
02
b100 6
#920090000000
1!
1%
1-
12
#920100000000
0!
0%
b101 *
0-
02
b101 6
#920110000000
1!
1%
1-
12
#920120000000
0!
0%
b110 *
0-
02
b110 6
#920130000000
1!
1%
1-
12
#920140000000
0!
0%
b111 *
0-
02
b111 6
#920150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#920160000000
0!
0%
b0 *
0-
02
b0 6
#920170000000
1!
1%
1-
12
#920180000000
0!
0%
b1 *
0-
02
b1 6
#920190000000
1!
1%
1-
12
#920200000000
0!
0%
b10 *
0-
02
b10 6
#920210000000
1!
1%
1-
12
#920220000000
0!
0%
b11 *
0-
02
b11 6
#920230000000
1!
1%
1-
12
15
#920240000000
0!
0%
b100 *
0-
02
b100 6
#920250000000
1!
1%
1-
12
#920260000000
0!
0%
b101 *
0-
02
b101 6
#920270000000
1!
1%
1-
12
#920280000000
0!
0%
b110 *
0-
02
b110 6
#920290000000
1!
1%
1-
12
#920300000000
0!
0%
b111 *
0-
02
b111 6
#920310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#920320000000
0!
0%
b0 *
0-
02
b0 6
#920330000000
1!
1%
1-
12
#920340000000
0!
0%
b1 *
0-
02
b1 6
#920350000000
1!
1%
1-
12
#920360000000
0!
0%
b10 *
0-
02
b10 6
#920370000000
1!
1%
1-
12
#920380000000
0!
0%
b11 *
0-
02
b11 6
#920390000000
1!
1%
1-
12
15
#920400000000
0!
0%
b100 *
0-
02
b100 6
#920410000000
1!
1%
1-
12
#920420000000
0!
0%
b101 *
0-
02
b101 6
#920430000000
1!
1%
1-
12
#920440000000
0!
0%
b110 *
0-
02
b110 6
#920450000000
1!
1%
1-
12
#920460000000
0!
0%
b111 *
0-
02
b111 6
#920470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#920480000000
0!
0%
b0 *
0-
02
b0 6
#920490000000
1!
1%
1-
12
#920500000000
0!
0%
b1 *
0-
02
b1 6
#920510000000
1!
1%
1-
12
#920520000000
0!
0%
b10 *
0-
02
b10 6
#920530000000
1!
1%
1-
12
#920540000000
0!
0%
b11 *
0-
02
b11 6
#920550000000
1!
1%
1-
12
15
#920560000000
0!
0%
b100 *
0-
02
b100 6
#920570000000
1!
1%
1-
12
#920580000000
0!
0%
b101 *
0-
02
b101 6
#920590000000
1!
1%
1-
12
#920600000000
0!
0%
b110 *
0-
02
b110 6
#920610000000
1!
1%
1-
12
#920620000000
0!
0%
b111 *
0-
02
b111 6
#920630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#920640000000
0!
0%
b0 *
0-
02
b0 6
#920650000000
1!
1%
1-
12
#920660000000
0!
0%
b1 *
0-
02
b1 6
#920670000000
1!
1%
1-
12
#920680000000
0!
0%
b10 *
0-
02
b10 6
#920690000000
1!
1%
1-
12
#920700000000
0!
0%
b11 *
0-
02
b11 6
#920710000000
1!
1%
1-
12
15
#920720000000
0!
0%
b100 *
0-
02
b100 6
#920730000000
1!
1%
1-
12
#920740000000
0!
0%
b101 *
0-
02
b101 6
#920750000000
1!
1%
1-
12
#920760000000
0!
0%
b110 *
0-
02
b110 6
#920770000000
1!
1%
1-
12
#920780000000
0!
0%
b111 *
0-
02
b111 6
#920790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#920800000000
0!
0%
b0 *
0-
02
b0 6
#920810000000
1!
1%
1-
12
#920820000000
0!
0%
b1 *
0-
02
b1 6
#920830000000
1!
1%
1-
12
#920840000000
0!
0%
b10 *
0-
02
b10 6
#920850000000
1!
1%
1-
12
#920860000000
0!
0%
b11 *
0-
02
b11 6
#920870000000
1!
1%
1-
12
15
#920880000000
0!
0%
b100 *
0-
02
b100 6
#920890000000
1!
1%
1-
12
#920900000000
0!
0%
b101 *
0-
02
b101 6
#920910000000
1!
1%
1-
12
#920920000000
0!
0%
b110 *
0-
02
b110 6
#920930000000
1!
1%
1-
12
#920940000000
0!
0%
b111 *
0-
02
b111 6
#920950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#920960000000
0!
0%
b0 *
0-
02
b0 6
#920970000000
1!
1%
1-
12
#920980000000
0!
0%
b1 *
0-
02
b1 6
#920990000000
1!
1%
1-
12
#921000000000
0!
0%
b10 *
0-
02
b10 6
#921010000000
1!
1%
1-
12
#921020000000
0!
0%
b11 *
0-
02
b11 6
#921030000000
1!
1%
1-
12
15
#921040000000
0!
0%
b100 *
0-
02
b100 6
#921050000000
1!
1%
1-
12
#921060000000
0!
0%
b101 *
0-
02
b101 6
#921070000000
1!
1%
1-
12
#921080000000
0!
0%
b110 *
0-
02
b110 6
#921090000000
1!
1%
1-
12
#921100000000
0!
0%
b111 *
0-
02
b111 6
#921110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#921120000000
0!
0%
b0 *
0-
02
b0 6
#921130000000
1!
1%
1-
12
#921140000000
0!
0%
b1 *
0-
02
b1 6
#921150000000
1!
1%
1-
12
#921160000000
0!
0%
b10 *
0-
02
b10 6
#921170000000
1!
1%
1-
12
#921180000000
0!
0%
b11 *
0-
02
b11 6
#921190000000
1!
1%
1-
12
15
#921200000000
0!
0%
b100 *
0-
02
b100 6
#921210000000
1!
1%
1-
12
#921220000000
0!
0%
b101 *
0-
02
b101 6
#921230000000
1!
1%
1-
12
#921240000000
0!
0%
b110 *
0-
02
b110 6
#921250000000
1!
1%
1-
12
#921260000000
0!
0%
b111 *
0-
02
b111 6
#921270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#921280000000
0!
0%
b0 *
0-
02
b0 6
#921290000000
1!
1%
1-
12
#921300000000
0!
0%
b1 *
0-
02
b1 6
#921310000000
1!
1%
1-
12
#921320000000
0!
0%
b10 *
0-
02
b10 6
#921330000000
1!
1%
1-
12
#921340000000
0!
0%
b11 *
0-
02
b11 6
#921350000000
1!
1%
1-
12
15
#921360000000
0!
0%
b100 *
0-
02
b100 6
#921370000000
1!
1%
1-
12
#921380000000
0!
0%
b101 *
0-
02
b101 6
#921390000000
1!
1%
1-
12
#921400000000
0!
0%
b110 *
0-
02
b110 6
#921410000000
1!
1%
1-
12
#921420000000
0!
0%
b111 *
0-
02
b111 6
#921430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#921440000000
0!
0%
b0 *
0-
02
b0 6
#921450000000
1!
1%
1-
12
#921460000000
0!
0%
b1 *
0-
02
b1 6
#921470000000
1!
1%
1-
12
#921480000000
0!
0%
b10 *
0-
02
b10 6
#921490000000
1!
1%
1-
12
#921500000000
0!
0%
b11 *
0-
02
b11 6
#921510000000
1!
1%
1-
12
15
#921520000000
0!
0%
b100 *
0-
02
b100 6
#921530000000
1!
1%
1-
12
#921540000000
0!
0%
b101 *
0-
02
b101 6
#921550000000
1!
1%
1-
12
#921560000000
0!
0%
b110 *
0-
02
b110 6
#921570000000
1!
1%
1-
12
#921580000000
0!
0%
b111 *
0-
02
b111 6
#921590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#921600000000
0!
0%
b0 *
0-
02
b0 6
#921610000000
1!
1%
1-
12
#921620000000
0!
0%
b1 *
0-
02
b1 6
#921630000000
1!
1%
1-
12
#921640000000
0!
0%
b10 *
0-
02
b10 6
#921650000000
1!
1%
1-
12
#921660000000
0!
0%
b11 *
0-
02
b11 6
#921670000000
1!
1%
1-
12
15
#921680000000
0!
0%
b100 *
0-
02
b100 6
#921690000000
1!
1%
1-
12
#921700000000
0!
0%
b101 *
0-
02
b101 6
#921710000000
1!
1%
1-
12
#921720000000
0!
0%
b110 *
0-
02
b110 6
#921730000000
1!
1%
1-
12
#921740000000
0!
0%
b111 *
0-
02
b111 6
#921750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#921760000000
0!
0%
b0 *
0-
02
b0 6
#921770000000
1!
1%
1-
12
#921780000000
0!
0%
b1 *
0-
02
b1 6
#921790000000
1!
1%
1-
12
#921800000000
0!
0%
b10 *
0-
02
b10 6
#921810000000
1!
1%
1-
12
#921820000000
0!
0%
b11 *
0-
02
b11 6
#921830000000
1!
1%
1-
12
15
#921840000000
0!
0%
b100 *
0-
02
b100 6
#921850000000
1!
1%
1-
12
#921860000000
0!
0%
b101 *
0-
02
b101 6
#921870000000
1!
1%
1-
12
#921880000000
0!
0%
b110 *
0-
02
b110 6
#921890000000
1!
1%
1-
12
#921900000000
0!
0%
b111 *
0-
02
b111 6
#921910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#921920000000
0!
0%
b0 *
0-
02
b0 6
#921930000000
1!
1%
1-
12
#921940000000
0!
0%
b1 *
0-
02
b1 6
#921950000000
1!
1%
1-
12
#921960000000
0!
0%
b10 *
0-
02
b10 6
#921970000000
1!
1%
1-
12
#921980000000
0!
0%
b11 *
0-
02
b11 6
#921990000000
1!
1%
1-
12
15
#922000000000
0!
0%
b100 *
0-
02
b100 6
#922010000000
1!
1%
1-
12
#922020000000
0!
0%
b101 *
0-
02
b101 6
#922030000000
1!
1%
1-
12
#922040000000
0!
0%
b110 *
0-
02
b110 6
#922050000000
1!
1%
1-
12
#922060000000
0!
0%
b111 *
0-
02
b111 6
#922070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#922080000000
0!
0%
b0 *
0-
02
b0 6
#922090000000
1!
1%
1-
12
#922100000000
0!
0%
b1 *
0-
02
b1 6
#922110000000
1!
1%
1-
12
#922120000000
0!
0%
b10 *
0-
02
b10 6
#922130000000
1!
1%
1-
12
#922140000000
0!
0%
b11 *
0-
02
b11 6
#922150000000
1!
1%
1-
12
15
#922160000000
0!
0%
b100 *
0-
02
b100 6
#922170000000
1!
1%
1-
12
#922180000000
0!
0%
b101 *
0-
02
b101 6
#922190000000
1!
1%
1-
12
#922200000000
0!
0%
b110 *
0-
02
b110 6
#922210000000
1!
1%
1-
12
#922220000000
0!
0%
b111 *
0-
02
b111 6
#922230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#922240000000
0!
0%
b0 *
0-
02
b0 6
#922250000000
1!
1%
1-
12
#922260000000
0!
0%
b1 *
0-
02
b1 6
#922270000000
1!
1%
1-
12
#922280000000
0!
0%
b10 *
0-
02
b10 6
#922290000000
1!
1%
1-
12
#922300000000
0!
0%
b11 *
0-
02
b11 6
#922310000000
1!
1%
1-
12
15
#922320000000
0!
0%
b100 *
0-
02
b100 6
#922330000000
1!
1%
1-
12
#922340000000
0!
0%
b101 *
0-
02
b101 6
#922350000000
1!
1%
1-
12
#922360000000
0!
0%
b110 *
0-
02
b110 6
#922370000000
1!
1%
1-
12
#922380000000
0!
0%
b111 *
0-
02
b111 6
#922390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#922400000000
0!
0%
b0 *
0-
02
b0 6
#922410000000
1!
1%
1-
12
#922420000000
0!
0%
b1 *
0-
02
b1 6
#922430000000
1!
1%
1-
12
#922440000000
0!
0%
b10 *
0-
02
b10 6
#922450000000
1!
1%
1-
12
#922460000000
0!
0%
b11 *
0-
02
b11 6
#922470000000
1!
1%
1-
12
15
#922480000000
0!
0%
b100 *
0-
02
b100 6
#922490000000
1!
1%
1-
12
#922500000000
0!
0%
b101 *
0-
02
b101 6
#922510000000
1!
1%
1-
12
#922520000000
0!
0%
b110 *
0-
02
b110 6
#922530000000
1!
1%
1-
12
#922540000000
0!
0%
b111 *
0-
02
b111 6
#922550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#922560000000
0!
0%
b0 *
0-
02
b0 6
#922570000000
1!
1%
1-
12
#922580000000
0!
0%
b1 *
0-
02
b1 6
#922590000000
1!
1%
1-
12
#922600000000
0!
0%
b10 *
0-
02
b10 6
#922610000000
1!
1%
1-
12
#922620000000
0!
0%
b11 *
0-
02
b11 6
#922630000000
1!
1%
1-
12
15
#922640000000
0!
0%
b100 *
0-
02
b100 6
#922650000000
1!
1%
1-
12
#922660000000
0!
0%
b101 *
0-
02
b101 6
#922670000000
1!
1%
1-
12
#922680000000
0!
0%
b110 *
0-
02
b110 6
#922690000000
1!
1%
1-
12
#922700000000
0!
0%
b111 *
0-
02
b111 6
#922710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#922720000000
0!
0%
b0 *
0-
02
b0 6
#922730000000
1!
1%
1-
12
#922740000000
0!
0%
b1 *
0-
02
b1 6
#922750000000
1!
1%
1-
12
#922760000000
0!
0%
b10 *
0-
02
b10 6
#922770000000
1!
1%
1-
12
#922780000000
0!
0%
b11 *
0-
02
b11 6
#922790000000
1!
1%
1-
12
15
#922800000000
0!
0%
b100 *
0-
02
b100 6
#922810000000
1!
1%
1-
12
#922820000000
0!
0%
b101 *
0-
02
b101 6
#922830000000
1!
1%
1-
12
#922840000000
0!
0%
b110 *
0-
02
b110 6
#922850000000
1!
1%
1-
12
#922860000000
0!
0%
b111 *
0-
02
b111 6
#922870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#922880000000
0!
0%
b0 *
0-
02
b0 6
#922890000000
1!
1%
1-
12
#922900000000
0!
0%
b1 *
0-
02
b1 6
#922910000000
1!
1%
1-
12
#922920000000
0!
0%
b10 *
0-
02
b10 6
#922930000000
1!
1%
1-
12
#922940000000
0!
0%
b11 *
0-
02
b11 6
#922950000000
1!
1%
1-
12
15
#922960000000
0!
0%
b100 *
0-
02
b100 6
#922970000000
1!
1%
1-
12
#922980000000
0!
0%
b101 *
0-
02
b101 6
#922990000000
1!
1%
1-
12
#923000000000
0!
0%
b110 *
0-
02
b110 6
#923010000000
1!
1%
1-
12
#923020000000
0!
0%
b111 *
0-
02
b111 6
#923030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#923040000000
0!
0%
b0 *
0-
02
b0 6
#923050000000
1!
1%
1-
12
#923060000000
0!
0%
b1 *
0-
02
b1 6
#923070000000
1!
1%
1-
12
#923080000000
0!
0%
b10 *
0-
02
b10 6
#923090000000
1!
1%
1-
12
#923100000000
0!
0%
b11 *
0-
02
b11 6
#923110000000
1!
1%
1-
12
15
#923120000000
0!
0%
b100 *
0-
02
b100 6
#923130000000
1!
1%
1-
12
#923140000000
0!
0%
b101 *
0-
02
b101 6
#923150000000
1!
1%
1-
12
#923160000000
0!
0%
b110 *
0-
02
b110 6
#923170000000
1!
1%
1-
12
#923180000000
0!
0%
b111 *
0-
02
b111 6
#923190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#923200000000
0!
0%
b0 *
0-
02
b0 6
#923210000000
1!
1%
1-
12
#923220000000
0!
0%
b1 *
0-
02
b1 6
#923230000000
1!
1%
1-
12
#923240000000
0!
0%
b10 *
0-
02
b10 6
#923250000000
1!
1%
1-
12
#923260000000
0!
0%
b11 *
0-
02
b11 6
#923270000000
1!
1%
1-
12
15
#923280000000
0!
0%
b100 *
0-
02
b100 6
#923290000000
1!
1%
1-
12
#923300000000
0!
0%
b101 *
0-
02
b101 6
#923310000000
1!
1%
1-
12
#923320000000
0!
0%
b110 *
0-
02
b110 6
#923330000000
1!
1%
1-
12
#923340000000
0!
0%
b111 *
0-
02
b111 6
#923350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#923360000000
0!
0%
b0 *
0-
02
b0 6
#923370000000
1!
1%
1-
12
#923380000000
0!
0%
b1 *
0-
02
b1 6
#923390000000
1!
1%
1-
12
#923400000000
0!
0%
b10 *
0-
02
b10 6
#923410000000
1!
1%
1-
12
#923420000000
0!
0%
b11 *
0-
02
b11 6
#923430000000
1!
1%
1-
12
15
#923440000000
0!
0%
b100 *
0-
02
b100 6
#923450000000
1!
1%
1-
12
#923460000000
0!
0%
b101 *
0-
02
b101 6
#923470000000
1!
1%
1-
12
#923480000000
0!
0%
b110 *
0-
02
b110 6
#923490000000
1!
1%
1-
12
#923500000000
0!
0%
b111 *
0-
02
b111 6
#923510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#923520000000
0!
0%
b0 *
0-
02
b0 6
#923530000000
1!
1%
1-
12
#923540000000
0!
0%
b1 *
0-
02
b1 6
#923550000000
1!
1%
1-
12
#923560000000
0!
0%
b10 *
0-
02
b10 6
#923570000000
1!
1%
1-
12
#923580000000
0!
0%
b11 *
0-
02
b11 6
#923590000000
1!
1%
1-
12
15
#923600000000
0!
0%
b100 *
0-
02
b100 6
#923610000000
1!
1%
1-
12
#923620000000
0!
0%
b101 *
0-
02
b101 6
#923630000000
1!
1%
1-
12
#923640000000
0!
0%
b110 *
0-
02
b110 6
#923650000000
1!
1%
1-
12
#923660000000
0!
0%
b111 *
0-
02
b111 6
#923670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#923680000000
0!
0%
b0 *
0-
02
b0 6
#923690000000
1!
1%
1-
12
#923700000000
0!
0%
b1 *
0-
02
b1 6
#923710000000
1!
1%
1-
12
#923720000000
0!
0%
b10 *
0-
02
b10 6
#923730000000
1!
1%
1-
12
#923740000000
0!
0%
b11 *
0-
02
b11 6
#923750000000
1!
1%
1-
12
15
#923760000000
0!
0%
b100 *
0-
02
b100 6
#923770000000
1!
1%
1-
12
#923780000000
0!
0%
b101 *
0-
02
b101 6
#923790000000
1!
1%
1-
12
#923800000000
0!
0%
b110 *
0-
02
b110 6
#923810000000
1!
1%
1-
12
#923820000000
0!
0%
b111 *
0-
02
b111 6
#923830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#923840000000
0!
0%
b0 *
0-
02
b0 6
#923850000000
1!
1%
1-
12
#923860000000
0!
0%
b1 *
0-
02
b1 6
#923870000000
1!
1%
1-
12
#923880000000
0!
0%
b10 *
0-
02
b10 6
#923890000000
1!
1%
1-
12
#923900000000
0!
0%
b11 *
0-
02
b11 6
#923910000000
1!
1%
1-
12
15
#923920000000
0!
0%
b100 *
0-
02
b100 6
#923930000000
1!
1%
1-
12
#923940000000
0!
0%
b101 *
0-
02
b101 6
#923950000000
1!
1%
1-
12
#923960000000
0!
0%
b110 *
0-
02
b110 6
#923970000000
1!
1%
1-
12
#923980000000
0!
0%
b111 *
0-
02
b111 6
#923990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#924000000000
0!
0%
b0 *
0-
02
b0 6
#924010000000
1!
1%
1-
12
#924020000000
0!
0%
b1 *
0-
02
b1 6
#924030000000
1!
1%
1-
12
#924040000000
0!
0%
b10 *
0-
02
b10 6
#924050000000
1!
1%
1-
12
#924060000000
0!
0%
b11 *
0-
02
b11 6
#924070000000
1!
1%
1-
12
15
#924080000000
0!
0%
b100 *
0-
02
b100 6
#924090000000
1!
1%
1-
12
#924100000000
0!
0%
b101 *
0-
02
b101 6
#924110000000
1!
1%
1-
12
#924120000000
0!
0%
b110 *
0-
02
b110 6
#924130000000
1!
1%
1-
12
#924140000000
0!
0%
b111 *
0-
02
b111 6
#924150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#924160000000
0!
0%
b0 *
0-
02
b0 6
#924170000000
1!
1%
1-
12
#924180000000
0!
0%
b1 *
0-
02
b1 6
#924190000000
1!
1%
1-
12
#924200000000
0!
0%
b10 *
0-
02
b10 6
#924210000000
1!
1%
1-
12
#924220000000
0!
0%
b11 *
0-
02
b11 6
#924230000000
1!
1%
1-
12
15
#924240000000
0!
0%
b100 *
0-
02
b100 6
#924250000000
1!
1%
1-
12
#924260000000
0!
0%
b101 *
0-
02
b101 6
#924270000000
1!
1%
1-
12
#924280000000
0!
0%
b110 *
0-
02
b110 6
#924290000000
1!
1%
1-
12
#924300000000
0!
0%
b111 *
0-
02
b111 6
#924310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#924320000000
0!
0%
b0 *
0-
02
b0 6
#924330000000
1!
1%
1-
12
#924340000000
0!
0%
b1 *
0-
02
b1 6
#924350000000
1!
1%
1-
12
#924360000000
0!
0%
b10 *
0-
02
b10 6
#924370000000
1!
1%
1-
12
#924380000000
0!
0%
b11 *
0-
02
b11 6
#924390000000
1!
1%
1-
12
15
#924400000000
0!
0%
b100 *
0-
02
b100 6
#924410000000
1!
1%
1-
12
#924420000000
0!
0%
b101 *
0-
02
b101 6
#924430000000
1!
1%
1-
12
#924440000000
0!
0%
b110 *
0-
02
b110 6
#924450000000
1!
1%
1-
12
#924460000000
0!
0%
b111 *
0-
02
b111 6
#924470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#924480000000
0!
0%
b0 *
0-
02
b0 6
#924490000000
1!
1%
1-
12
#924500000000
0!
0%
b1 *
0-
02
b1 6
#924510000000
1!
1%
1-
12
#924520000000
0!
0%
b10 *
0-
02
b10 6
#924530000000
1!
1%
1-
12
#924540000000
0!
0%
b11 *
0-
02
b11 6
#924550000000
1!
1%
1-
12
15
#924560000000
0!
0%
b100 *
0-
02
b100 6
#924570000000
1!
1%
1-
12
#924580000000
0!
0%
b101 *
0-
02
b101 6
#924590000000
1!
1%
1-
12
#924600000000
0!
0%
b110 *
0-
02
b110 6
#924610000000
1!
1%
1-
12
#924620000000
0!
0%
b111 *
0-
02
b111 6
#924630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#924640000000
0!
0%
b0 *
0-
02
b0 6
#924650000000
1!
1%
1-
12
#924660000000
0!
0%
b1 *
0-
02
b1 6
#924670000000
1!
1%
1-
12
#924680000000
0!
0%
b10 *
0-
02
b10 6
#924690000000
1!
1%
1-
12
#924700000000
0!
0%
b11 *
0-
02
b11 6
#924710000000
1!
1%
1-
12
15
#924720000000
0!
0%
b100 *
0-
02
b100 6
#924730000000
1!
1%
1-
12
#924740000000
0!
0%
b101 *
0-
02
b101 6
#924750000000
1!
1%
1-
12
#924760000000
0!
0%
b110 *
0-
02
b110 6
#924770000000
1!
1%
1-
12
#924780000000
0!
0%
b111 *
0-
02
b111 6
#924790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#924800000000
0!
0%
b0 *
0-
02
b0 6
#924810000000
1!
1%
1-
12
#924820000000
0!
0%
b1 *
0-
02
b1 6
#924830000000
1!
1%
1-
12
#924840000000
0!
0%
b10 *
0-
02
b10 6
#924850000000
1!
1%
1-
12
#924860000000
0!
0%
b11 *
0-
02
b11 6
#924870000000
1!
1%
1-
12
15
#924880000000
0!
0%
b100 *
0-
02
b100 6
#924890000000
1!
1%
1-
12
#924900000000
0!
0%
b101 *
0-
02
b101 6
#924910000000
1!
1%
1-
12
#924920000000
0!
0%
b110 *
0-
02
b110 6
#924930000000
1!
1%
1-
12
#924940000000
0!
0%
b111 *
0-
02
b111 6
#924950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#924960000000
0!
0%
b0 *
0-
02
b0 6
#924970000000
1!
1%
1-
12
#924980000000
0!
0%
b1 *
0-
02
b1 6
#924990000000
1!
1%
1-
12
#925000000000
0!
0%
b10 *
0-
02
b10 6
#925010000000
1!
1%
1-
12
#925020000000
0!
0%
b11 *
0-
02
b11 6
#925030000000
1!
1%
1-
12
15
#925040000000
0!
0%
b100 *
0-
02
b100 6
#925050000000
1!
1%
1-
12
#925060000000
0!
0%
b101 *
0-
02
b101 6
#925070000000
1!
1%
1-
12
#925080000000
0!
0%
b110 *
0-
02
b110 6
#925090000000
1!
1%
1-
12
#925100000000
0!
0%
b111 *
0-
02
b111 6
#925110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#925120000000
0!
0%
b0 *
0-
02
b0 6
#925130000000
1!
1%
1-
12
#925140000000
0!
0%
b1 *
0-
02
b1 6
#925150000000
1!
1%
1-
12
#925160000000
0!
0%
b10 *
0-
02
b10 6
#925170000000
1!
1%
1-
12
#925180000000
0!
0%
b11 *
0-
02
b11 6
#925190000000
1!
1%
1-
12
15
#925200000000
0!
0%
b100 *
0-
02
b100 6
#925210000000
1!
1%
1-
12
#925220000000
0!
0%
b101 *
0-
02
b101 6
#925230000000
1!
1%
1-
12
#925240000000
0!
0%
b110 *
0-
02
b110 6
#925250000000
1!
1%
1-
12
#925260000000
0!
0%
b111 *
0-
02
b111 6
#925270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#925280000000
0!
0%
b0 *
0-
02
b0 6
#925290000000
1!
1%
1-
12
#925300000000
0!
0%
b1 *
0-
02
b1 6
#925310000000
1!
1%
1-
12
#925320000000
0!
0%
b10 *
0-
02
b10 6
#925330000000
1!
1%
1-
12
#925340000000
0!
0%
b11 *
0-
02
b11 6
#925350000000
1!
1%
1-
12
15
#925360000000
0!
0%
b100 *
0-
02
b100 6
#925370000000
1!
1%
1-
12
#925380000000
0!
0%
b101 *
0-
02
b101 6
#925390000000
1!
1%
1-
12
#925400000000
0!
0%
b110 *
0-
02
b110 6
#925410000000
1!
1%
1-
12
#925420000000
0!
0%
b111 *
0-
02
b111 6
#925430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#925440000000
0!
0%
b0 *
0-
02
b0 6
#925450000000
1!
1%
1-
12
#925460000000
0!
0%
b1 *
0-
02
b1 6
#925470000000
1!
1%
1-
12
#925480000000
0!
0%
b10 *
0-
02
b10 6
#925490000000
1!
1%
1-
12
#925500000000
0!
0%
b11 *
0-
02
b11 6
#925510000000
1!
1%
1-
12
15
#925520000000
0!
0%
b100 *
0-
02
b100 6
#925530000000
1!
1%
1-
12
#925540000000
0!
0%
b101 *
0-
02
b101 6
#925550000000
1!
1%
1-
12
#925560000000
0!
0%
b110 *
0-
02
b110 6
#925570000000
1!
1%
1-
12
#925580000000
0!
0%
b111 *
0-
02
b111 6
#925590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#925600000000
0!
0%
b0 *
0-
02
b0 6
#925610000000
1!
1%
1-
12
#925620000000
0!
0%
b1 *
0-
02
b1 6
#925630000000
1!
1%
1-
12
#925640000000
0!
0%
b10 *
0-
02
b10 6
#925650000000
1!
1%
1-
12
#925660000000
0!
0%
b11 *
0-
02
b11 6
#925670000000
1!
1%
1-
12
15
#925680000000
0!
0%
b100 *
0-
02
b100 6
#925690000000
1!
1%
1-
12
#925700000000
0!
0%
b101 *
0-
02
b101 6
#925710000000
1!
1%
1-
12
#925720000000
0!
0%
b110 *
0-
02
b110 6
#925730000000
1!
1%
1-
12
#925740000000
0!
0%
b111 *
0-
02
b111 6
#925750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#925760000000
0!
0%
b0 *
0-
02
b0 6
#925770000000
1!
1%
1-
12
#925780000000
0!
0%
b1 *
0-
02
b1 6
#925790000000
1!
1%
1-
12
#925800000000
0!
0%
b10 *
0-
02
b10 6
#925810000000
1!
1%
1-
12
#925820000000
0!
0%
b11 *
0-
02
b11 6
#925830000000
1!
1%
1-
12
15
#925840000000
0!
0%
b100 *
0-
02
b100 6
#925850000000
1!
1%
1-
12
#925860000000
0!
0%
b101 *
0-
02
b101 6
#925870000000
1!
1%
1-
12
#925880000000
0!
0%
b110 *
0-
02
b110 6
#925890000000
1!
1%
1-
12
#925900000000
0!
0%
b111 *
0-
02
b111 6
#925910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#925920000000
0!
0%
b0 *
0-
02
b0 6
#925930000000
1!
1%
1-
12
#925940000000
0!
0%
b1 *
0-
02
b1 6
#925950000000
1!
1%
1-
12
#925960000000
0!
0%
b10 *
0-
02
b10 6
#925970000000
1!
1%
1-
12
#925980000000
0!
0%
b11 *
0-
02
b11 6
#925990000000
1!
1%
1-
12
15
#926000000000
0!
0%
b100 *
0-
02
b100 6
#926010000000
1!
1%
1-
12
#926020000000
0!
0%
b101 *
0-
02
b101 6
#926030000000
1!
1%
1-
12
#926040000000
0!
0%
b110 *
0-
02
b110 6
#926050000000
1!
1%
1-
12
#926060000000
0!
0%
b111 *
0-
02
b111 6
#926070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#926080000000
0!
0%
b0 *
0-
02
b0 6
#926090000000
1!
1%
1-
12
#926100000000
0!
0%
b1 *
0-
02
b1 6
#926110000000
1!
1%
1-
12
#926120000000
0!
0%
b10 *
0-
02
b10 6
#926130000000
1!
1%
1-
12
#926140000000
0!
0%
b11 *
0-
02
b11 6
#926150000000
1!
1%
1-
12
15
#926160000000
0!
0%
b100 *
0-
02
b100 6
#926170000000
1!
1%
1-
12
#926180000000
0!
0%
b101 *
0-
02
b101 6
#926190000000
1!
1%
1-
12
#926200000000
0!
0%
b110 *
0-
02
b110 6
#926210000000
1!
1%
1-
12
#926220000000
0!
0%
b111 *
0-
02
b111 6
#926230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#926240000000
0!
0%
b0 *
0-
02
b0 6
#926250000000
1!
1%
1-
12
#926260000000
0!
0%
b1 *
0-
02
b1 6
#926270000000
1!
1%
1-
12
#926280000000
0!
0%
b10 *
0-
02
b10 6
#926290000000
1!
1%
1-
12
#926300000000
0!
0%
b11 *
0-
02
b11 6
#926310000000
1!
1%
1-
12
15
#926320000000
0!
0%
b100 *
0-
02
b100 6
#926330000000
1!
1%
1-
12
#926340000000
0!
0%
b101 *
0-
02
b101 6
#926350000000
1!
1%
1-
12
#926360000000
0!
0%
b110 *
0-
02
b110 6
#926370000000
1!
1%
1-
12
#926380000000
0!
0%
b111 *
0-
02
b111 6
#926390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#926400000000
0!
0%
b0 *
0-
02
b0 6
#926410000000
1!
1%
1-
12
#926420000000
0!
0%
b1 *
0-
02
b1 6
#926430000000
1!
1%
1-
12
#926440000000
0!
0%
b10 *
0-
02
b10 6
#926450000000
1!
1%
1-
12
#926460000000
0!
0%
b11 *
0-
02
b11 6
#926470000000
1!
1%
1-
12
15
#926480000000
0!
0%
b100 *
0-
02
b100 6
#926490000000
1!
1%
1-
12
#926500000000
0!
0%
b101 *
0-
02
b101 6
#926510000000
1!
1%
1-
12
#926520000000
0!
0%
b110 *
0-
02
b110 6
#926530000000
1!
1%
1-
12
#926540000000
0!
0%
b111 *
0-
02
b111 6
#926550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#926560000000
0!
0%
b0 *
0-
02
b0 6
#926570000000
1!
1%
1-
12
#926580000000
0!
0%
b1 *
0-
02
b1 6
#926590000000
1!
1%
1-
12
#926600000000
0!
0%
b10 *
0-
02
b10 6
#926610000000
1!
1%
1-
12
#926620000000
0!
0%
b11 *
0-
02
b11 6
#926630000000
1!
1%
1-
12
15
#926640000000
0!
0%
b100 *
0-
02
b100 6
#926650000000
1!
1%
1-
12
#926660000000
0!
0%
b101 *
0-
02
b101 6
#926670000000
1!
1%
1-
12
#926680000000
0!
0%
b110 *
0-
02
b110 6
#926690000000
1!
1%
1-
12
#926700000000
0!
0%
b111 *
0-
02
b111 6
#926710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#926720000000
0!
0%
b0 *
0-
02
b0 6
#926730000000
1!
1%
1-
12
#926740000000
0!
0%
b1 *
0-
02
b1 6
#926750000000
1!
1%
1-
12
#926760000000
0!
0%
b10 *
0-
02
b10 6
#926770000000
1!
1%
1-
12
#926780000000
0!
0%
b11 *
0-
02
b11 6
#926790000000
1!
1%
1-
12
15
#926800000000
0!
0%
b100 *
0-
02
b100 6
#926810000000
1!
1%
1-
12
#926820000000
0!
0%
b101 *
0-
02
b101 6
#926830000000
1!
1%
1-
12
#926840000000
0!
0%
b110 *
0-
02
b110 6
#926850000000
1!
1%
1-
12
#926860000000
0!
0%
b111 *
0-
02
b111 6
#926870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#926880000000
0!
0%
b0 *
0-
02
b0 6
#926890000000
1!
1%
1-
12
#926900000000
0!
0%
b1 *
0-
02
b1 6
#926910000000
1!
1%
1-
12
#926920000000
0!
0%
b10 *
0-
02
b10 6
#926930000000
1!
1%
1-
12
#926940000000
0!
0%
b11 *
0-
02
b11 6
#926950000000
1!
1%
1-
12
15
#926960000000
0!
0%
b100 *
0-
02
b100 6
#926970000000
1!
1%
1-
12
#926980000000
0!
0%
b101 *
0-
02
b101 6
#926990000000
1!
1%
1-
12
#927000000000
0!
0%
b110 *
0-
02
b110 6
#927010000000
1!
1%
1-
12
#927020000000
0!
0%
b111 *
0-
02
b111 6
#927030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#927040000000
0!
0%
b0 *
0-
02
b0 6
#927050000000
1!
1%
1-
12
#927060000000
0!
0%
b1 *
0-
02
b1 6
#927070000000
1!
1%
1-
12
#927080000000
0!
0%
b10 *
0-
02
b10 6
#927090000000
1!
1%
1-
12
#927100000000
0!
0%
b11 *
0-
02
b11 6
#927110000000
1!
1%
1-
12
15
#927120000000
0!
0%
b100 *
0-
02
b100 6
#927130000000
1!
1%
1-
12
#927140000000
0!
0%
b101 *
0-
02
b101 6
#927150000000
1!
1%
1-
12
#927160000000
0!
0%
b110 *
0-
02
b110 6
#927170000000
1!
1%
1-
12
#927180000000
0!
0%
b111 *
0-
02
b111 6
#927190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#927200000000
0!
0%
b0 *
0-
02
b0 6
#927210000000
1!
1%
1-
12
#927220000000
0!
0%
b1 *
0-
02
b1 6
#927230000000
1!
1%
1-
12
#927240000000
0!
0%
b10 *
0-
02
b10 6
#927250000000
1!
1%
1-
12
#927260000000
0!
0%
b11 *
0-
02
b11 6
#927270000000
1!
1%
1-
12
15
#927280000000
0!
0%
b100 *
0-
02
b100 6
#927290000000
1!
1%
1-
12
#927300000000
0!
0%
b101 *
0-
02
b101 6
#927310000000
1!
1%
1-
12
#927320000000
0!
0%
b110 *
0-
02
b110 6
#927330000000
1!
1%
1-
12
#927340000000
0!
0%
b111 *
0-
02
b111 6
#927350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#927360000000
0!
0%
b0 *
0-
02
b0 6
#927370000000
1!
1%
1-
12
#927380000000
0!
0%
b1 *
0-
02
b1 6
#927390000000
1!
1%
1-
12
#927400000000
0!
0%
b10 *
0-
02
b10 6
#927410000000
1!
1%
1-
12
#927420000000
0!
0%
b11 *
0-
02
b11 6
#927430000000
1!
1%
1-
12
15
#927440000000
0!
0%
b100 *
0-
02
b100 6
#927450000000
1!
1%
1-
12
#927460000000
0!
0%
b101 *
0-
02
b101 6
#927470000000
1!
1%
1-
12
#927480000000
0!
0%
b110 *
0-
02
b110 6
#927490000000
1!
1%
1-
12
#927500000000
0!
0%
b111 *
0-
02
b111 6
#927510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#927520000000
0!
0%
b0 *
0-
02
b0 6
#927530000000
1!
1%
1-
12
#927540000000
0!
0%
b1 *
0-
02
b1 6
#927550000000
1!
1%
1-
12
#927560000000
0!
0%
b10 *
0-
02
b10 6
#927570000000
1!
1%
1-
12
#927580000000
0!
0%
b11 *
0-
02
b11 6
#927590000000
1!
1%
1-
12
15
#927600000000
0!
0%
b100 *
0-
02
b100 6
#927610000000
1!
1%
1-
12
#927620000000
0!
0%
b101 *
0-
02
b101 6
#927630000000
1!
1%
1-
12
#927640000000
0!
0%
b110 *
0-
02
b110 6
#927650000000
1!
1%
1-
12
#927660000000
0!
0%
b111 *
0-
02
b111 6
#927670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#927680000000
0!
0%
b0 *
0-
02
b0 6
#927690000000
1!
1%
1-
12
#927700000000
0!
0%
b1 *
0-
02
b1 6
#927710000000
1!
1%
1-
12
#927720000000
0!
0%
b10 *
0-
02
b10 6
#927730000000
1!
1%
1-
12
#927740000000
0!
0%
b11 *
0-
02
b11 6
#927750000000
1!
1%
1-
12
15
#927760000000
0!
0%
b100 *
0-
02
b100 6
#927770000000
1!
1%
1-
12
#927780000000
0!
0%
b101 *
0-
02
b101 6
#927790000000
1!
1%
1-
12
#927800000000
0!
0%
b110 *
0-
02
b110 6
#927810000000
1!
1%
1-
12
#927820000000
0!
0%
b111 *
0-
02
b111 6
#927830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#927840000000
0!
0%
b0 *
0-
02
b0 6
#927850000000
1!
1%
1-
12
#927860000000
0!
0%
b1 *
0-
02
b1 6
#927870000000
1!
1%
1-
12
#927880000000
0!
0%
b10 *
0-
02
b10 6
#927890000000
1!
1%
1-
12
#927900000000
0!
0%
b11 *
0-
02
b11 6
#927910000000
1!
1%
1-
12
15
#927920000000
0!
0%
b100 *
0-
02
b100 6
#927930000000
1!
1%
1-
12
#927940000000
0!
0%
b101 *
0-
02
b101 6
#927950000000
1!
1%
1-
12
#927960000000
0!
0%
b110 *
0-
02
b110 6
#927970000000
1!
1%
1-
12
#927980000000
0!
0%
b111 *
0-
02
b111 6
#927990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#928000000000
0!
0%
b0 *
0-
02
b0 6
#928010000000
1!
1%
1-
12
#928020000000
0!
0%
b1 *
0-
02
b1 6
#928030000000
1!
1%
1-
12
#928040000000
0!
0%
b10 *
0-
02
b10 6
#928050000000
1!
1%
1-
12
#928060000000
0!
0%
b11 *
0-
02
b11 6
#928070000000
1!
1%
1-
12
15
#928080000000
0!
0%
b100 *
0-
02
b100 6
#928090000000
1!
1%
1-
12
#928100000000
0!
0%
b101 *
0-
02
b101 6
#928110000000
1!
1%
1-
12
#928120000000
0!
0%
b110 *
0-
02
b110 6
#928130000000
1!
1%
1-
12
#928140000000
0!
0%
b111 *
0-
02
b111 6
#928150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#928160000000
0!
0%
b0 *
0-
02
b0 6
#928170000000
1!
1%
1-
12
#928180000000
0!
0%
b1 *
0-
02
b1 6
#928190000000
1!
1%
1-
12
#928200000000
0!
0%
b10 *
0-
02
b10 6
#928210000000
1!
1%
1-
12
#928220000000
0!
0%
b11 *
0-
02
b11 6
#928230000000
1!
1%
1-
12
15
#928240000000
0!
0%
b100 *
0-
02
b100 6
#928250000000
1!
1%
1-
12
#928260000000
0!
0%
b101 *
0-
02
b101 6
#928270000000
1!
1%
1-
12
#928280000000
0!
0%
b110 *
0-
02
b110 6
#928290000000
1!
1%
1-
12
#928300000000
0!
0%
b111 *
0-
02
b111 6
#928310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#928320000000
0!
0%
b0 *
0-
02
b0 6
#928330000000
1!
1%
1-
12
#928340000000
0!
0%
b1 *
0-
02
b1 6
#928350000000
1!
1%
1-
12
#928360000000
0!
0%
b10 *
0-
02
b10 6
#928370000000
1!
1%
1-
12
#928380000000
0!
0%
b11 *
0-
02
b11 6
#928390000000
1!
1%
1-
12
15
#928400000000
0!
0%
b100 *
0-
02
b100 6
#928410000000
1!
1%
1-
12
#928420000000
0!
0%
b101 *
0-
02
b101 6
#928430000000
1!
1%
1-
12
#928440000000
0!
0%
b110 *
0-
02
b110 6
#928450000000
1!
1%
1-
12
#928460000000
0!
0%
b111 *
0-
02
b111 6
#928470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#928480000000
0!
0%
b0 *
0-
02
b0 6
#928490000000
1!
1%
1-
12
#928500000000
0!
0%
b1 *
0-
02
b1 6
#928510000000
1!
1%
1-
12
#928520000000
0!
0%
b10 *
0-
02
b10 6
#928530000000
1!
1%
1-
12
#928540000000
0!
0%
b11 *
0-
02
b11 6
#928550000000
1!
1%
1-
12
15
#928560000000
0!
0%
b100 *
0-
02
b100 6
#928570000000
1!
1%
1-
12
#928580000000
0!
0%
b101 *
0-
02
b101 6
#928590000000
1!
1%
1-
12
#928600000000
0!
0%
b110 *
0-
02
b110 6
#928610000000
1!
1%
1-
12
#928620000000
0!
0%
b111 *
0-
02
b111 6
#928630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#928640000000
0!
0%
b0 *
0-
02
b0 6
#928650000000
1!
1%
1-
12
#928660000000
0!
0%
b1 *
0-
02
b1 6
#928670000000
1!
1%
1-
12
#928680000000
0!
0%
b10 *
0-
02
b10 6
#928690000000
1!
1%
1-
12
#928700000000
0!
0%
b11 *
0-
02
b11 6
#928710000000
1!
1%
1-
12
15
#928720000000
0!
0%
b100 *
0-
02
b100 6
#928730000000
1!
1%
1-
12
#928740000000
0!
0%
b101 *
0-
02
b101 6
#928750000000
1!
1%
1-
12
#928760000000
0!
0%
b110 *
0-
02
b110 6
#928770000000
1!
1%
1-
12
#928780000000
0!
0%
b111 *
0-
02
b111 6
#928790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#928800000000
0!
0%
b0 *
0-
02
b0 6
#928810000000
1!
1%
1-
12
#928820000000
0!
0%
b1 *
0-
02
b1 6
#928830000000
1!
1%
1-
12
#928840000000
0!
0%
b10 *
0-
02
b10 6
#928850000000
1!
1%
1-
12
#928860000000
0!
0%
b11 *
0-
02
b11 6
#928870000000
1!
1%
1-
12
15
#928880000000
0!
0%
b100 *
0-
02
b100 6
#928890000000
1!
1%
1-
12
#928900000000
0!
0%
b101 *
0-
02
b101 6
#928910000000
1!
1%
1-
12
#928920000000
0!
0%
b110 *
0-
02
b110 6
#928930000000
1!
1%
1-
12
#928940000000
0!
0%
b111 *
0-
02
b111 6
#928950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#928960000000
0!
0%
b0 *
0-
02
b0 6
#928970000000
1!
1%
1-
12
#928980000000
0!
0%
b1 *
0-
02
b1 6
#928990000000
1!
1%
1-
12
#929000000000
0!
0%
b10 *
0-
02
b10 6
#929010000000
1!
1%
1-
12
#929020000000
0!
0%
b11 *
0-
02
b11 6
#929030000000
1!
1%
1-
12
15
#929040000000
0!
0%
b100 *
0-
02
b100 6
#929050000000
1!
1%
1-
12
#929060000000
0!
0%
b101 *
0-
02
b101 6
#929070000000
1!
1%
1-
12
#929080000000
0!
0%
b110 *
0-
02
b110 6
#929090000000
1!
1%
1-
12
#929100000000
0!
0%
b111 *
0-
02
b111 6
#929110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#929120000000
0!
0%
b0 *
0-
02
b0 6
#929130000000
1!
1%
1-
12
#929140000000
0!
0%
b1 *
0-
02
b1 6
#929150000000
1!
1%
1-
12
#929160000000
0!
0%
b10 *
0-
02
b10 6
#929170000000
1!
1%
1-
12
#929180000000
0!
0%
b11 *
0-
02
b11 6
#929190000000
1!
1%
1-
12
15
#929200000000
0!
0%
b100 *
0-
02
b100 6
#929210000000
1!
1%
1-
12
#929220000000
0!
0%
b101 *
0-
02
b101 6
#929230000000
1!
1%
1-
12
#929240000000
0!
0%
b110 *
0-
02
b110 6
#929250000000
1!
1%
1-
12
#929260000000
0!
0%
b111 *
0-
02
b111 6
#929270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#929280000000
0!
0%
b0 *
0-
02
b0 6
#929290000000
1!
1%
1-
12
#929300000000
0!
0%
b1 *
0-
02
b1 6
#929310000000
1!
1%
1-
12
#929320000000
0!
0%
b10 *
0-
02
b10 6
#929330000000
1!
1%
1-
12
#929340000000
0!
0%
b11 *
0-
02
b11 6
#929350000000
1!
1%
1-
12
15
#929360000000
0!
0%
b100 *
0-
02
b100 6
#929370000000
1!
1%
1-
12
#929380000000
0!
0%
b101 *
0-
02
b101 6
#929390000000
1!
1%
1-
12
#929400000000
0!
0%
b110 *
0-
02
b110 6
#929410000000
1!
1%
1-
12
#929420000000
0!
0%
b111 *
0-
02
b111 6
#929430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#929440000000
0!
0%
b0 *
0-
02
b0 6
#929450000000
1!
1%
1-
12
#929460000000
0!
0%
b1 *
0-
02
b1 6
#929470000000
1!
1%
1-
12
#929480000000
0!
0%
b10 *
0-
02
b10 6
#929490000000
1!
1%
1-
12
#929500000000
0!
0%
b11 *
0-
02
b11 6
#929510000000
1!
1%
1-
12
15
#929520000000
0!
0%
b100 *
0-
02
b100 6
#929530000000
1!
1%
1-
12
#929540000000
0!
0%
b101 *
0-
02
b101 6
#929550000000
1!
1%
1-
12
#929560000000
0!
0%
b110 *
0-
02
b110 6
#929570000000
1!
1%
1-
12
#929580000000
0!
0%
b111 *
0-
02
b111 6
#929590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#929600000000
0!
0%
b0 *
0-
02
b0 6
#929610000000
1!
1%
1-
12
#929620000000
0!
0%
b1 *
0-
02
b1 6
#929630000000
1!
1%
1-
12
#929640000000
0!
0%
b10 *
0-
02
b10 6
#929650000000
1!
1%
1-
12
#929660000000
0!
0%
b11 *
0-
02
b11 6
#929670000000
1!
1%
1-
12
15
#929680000000
0!
0%
b100 *
0-
02
b100 6
#929690000000
1!
1%
1-
12
#929700000000
0!
0%
b101 *
0-
02
b101 6
#929710000000
1!
1%
1-
12
#929720000000
0!
0%
b110 *
0-
02
b110 6
#929730000000
1!
1%
1-
12
#929740000000
0!
0%
b111 *
0-
02
b111 6
#929750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#929760000000
0!
0%
b0 *
0-
02
b0 6
#929770000000
1!
1%
1-
12
#929780000000
0!
0%
b1 *
0-
02
b1 6
#929790000000
1!
1%
1-
12
#929800000000
0!
0%
b10 *
0-
02
b10 6
#929810000000
1!
1%
1-
12
#929820000000
0!
0%
b11 *
0-
02
b11 6
#929830000000
1!
1%
1-
12
15
#929840000000
0!
0%
b100 *
0-
02
b100 6
#929850000000
1!
1%
1-
12
#929860000000
0!
0%
b101 *
0-
02
b101 6
#929870000000
1!
1%
1-
12
#929880000000
0!
0%
b110 *
0-
02
b110 6
#929890000000
1!
1%
1-
12
#929900000000
0!
0%
b111 *
0-
02
b111 6
#929910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#929920000000
0!
0%
b0 *
0-
02
b0 6
#929930000000
1!
1%
1-
12
#929940000000
0!
0%
b1 *
0-
02
b1 6
#929950000000
1!
1%
1-
12
#929960000000
0!
0%
b10 *
0-
02
b10 6
#929970000000
1!
1%
1-
12
#929980000000
0!
0%
b11 *
0-
02
b11 6
#929990000000
1!
1%
1-
12
15
#930000000000
0!
0%
b100 *
0-
02
b100 6
#930010000000
1!
1%
1-
12
#930020000000
0!
0%
b101 *
0-
02
b101 6
#930030000000
1!
1%
1-
12
#930040000000
0!
0%
b110 *
0-
02
b110 6
#930050000000
1!
1%
1-
12
#930060000000
0!
0%
b111 *
0-
02
b111 6
#930070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#930080000000
0!
0%
b0 *
0-
02
b0 6
#930090000000
1!
1%
1-
12
#930100000000
0!
0%
b1 *
0-
02
b1 6
#930110000000
1!
1%
1-
12
#930120000000
0!
0%
b10 *
0-
02
b10 6
#930130000000
1!
1%
1-
12
#930140000000
0!
0%
b11 *
0-
02
b11 6
#930150000000
1!
1%
1-
12
15
#930160000000
0!
0%
b100 *
0-
02
b100 6
#930170000000
1!
1%
1-
12
#930180000000
0!
0%
b101 *
0-
02
b101 6
#930190000000
1!
1%
1-
12
#930200000000
0!
0%
b110 *
0-
02
b110 6
#930210000000
1!
1%
1-
12
#930220000000
0!
0%
b111 *
0-
02
b111 6
#930230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#930240000000
0!
0%
b0 *
0-
02
b0 6
#930250000000
1!
1%
1-
12
#930260000000
0!
0%
b1 *
0-
02
b1 6
#930270000000
1!
1%
1-
12
#930280000000
0!
0%
b10 *
0-
02
b10 6
#930290000000
1!
1%
1-
12
#930300000000
0!
0%
b11 *
0-
02
b11 6
#930310000000
1!
1%
1-
12
15
#930320000000
0!
0%
b100 *
0-
02
b100 6
#930330000000
1!
1%
1-
12
#930340000000
0!
0%
b101 *
0-
02
b101 6
#930350000000
1!
1%
1-
12
#930360000000
0!
0%
b110 *
0-
02
b110 6
#930370000000
1!
1%
1-
12
#930380000000
0!
0%
b111 *
0-
02
b111 6
#930390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#930400000000
0!
0%
b0 *
0-
02
b0 6
#930410000000
1!
1%
1-
12
#930420000000
0!
0%
b1 *
0-
02
b1 6
#930430000000
1!
1%
1-
12
#930440000000
0!
0%
b10 *
0-
02
b10 6
#930450000000
1!
1%
1-
12
#930460000000
0!
0%
b11 *
0-
02
b11 6
#930470000000
1!
1%
1-
12
15
#930480000000
0!
0%
b100 *
0-
02
b100 6
#930490000000
1!
1%
1-
12
#930500000000
0!
0%
b101 *
0-
02
b101 6
#930510000000
1!
1%
1-
12
#930520000000
0!
0%
b110 *
0-
02
b110 6
#930530000000
1!
1%
1-
12
#930540000000
0!
0%
b111 *
0-
02
b111 6
#930550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#930560000000
0!
0%
b0 *
0-
02
b0 6
#930570000000
1!
1%
1-
12
#930580000000
0!
0%
b1 *
0-
02
b1 6
#930590000000
1!
1%
1-
12
#930600000000
0!
0%
b10 *
0-
02
b10 6
#930610000000
1!
1%
1-
12
#930620000000
0!
0%
b11 *
0-
02
b11 6
#930630000000
1!
1%
1-
12
15
#930640000000
0!
0%
b100 *
0-
02
b100 6
#930650000000
1!
1%
1-
12
#930660000000
0!
0%
b101 *
0-
02
b101 6
#930670000000
1!
1%
1-
12
#930680000000
0!
0%
b110 *
0-
02
b110 6
#930690000000
1!
1%
1-
12
#930700000000
0!
0%
b111 *
0-
02
b111 6
#930710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#930720000000
0!
0%
b0 *
0-
02
b0 6
#930730000000
1!
1%
1-
12
#930740000000
0!
0%
b1 *
0-
02
b1 6
#930750000000
1!
1%
1-
12
#930760000000
0!
0%
b10 *
0-
02
b10 6
#930770000000
1!
1%
1-
12
#930780000000
0!
0%
b11 *
0-
02
b11 6
#930790000000
1!
1%
1-
12
15
#930800000000
0!
0%
b100 *
0-
02
b100 6
#930810000000
1!
1%
1-
12
#930820000000
0!
0%
b101 *
0-
02
b101 6
#930830000000
1!
1%
1-
12
#930840000000
0!
0%
b110 *
0-
02
b110 6
#930850000000
1!
1%
1-
12
#930860000000
0!
0%
b111 *
0-
02
b111 6
#930870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#930880000000
0!
0%
b0 *
0-
02
b0 6
#930890000000
1!
1%
1-
12
#930900000000
0!
0%
b1 *
0-
02
b1 6
#930910000000
1!
1%
1-
12
#930920000000
0!
0%
b10 *
0-
02
b10 6
#930930000000
1!
1%
1-
12
#930940000000
0!
0%
b11 *
0-
02
b11 6
#930950000000
1!
1%
1-
12
15
#930960000000
0!
0%
b100 *
0-
02
b100 6
#930970000000
1!
1%
1-
12
#930980000000
0!
0%
b101 *
0-
02
b101 6
#930990000000
1!
1%
1-
12
#931000000000
0!
0%
b110 *
0-
02
b110 6
#931010000000
1!
1%
1-
12
#931020000000
0!
0%
b111 *
0-
02
b111 6
#931030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#931040000000
0!
0%
b0 *
0-
02
b0 6
#931050000000
1!
1%
1-
12
#931060000000
0!
0%
b1 *
0-
02
b1 6
#931070000000
1!
1%
1-
12
#931080000000
0!
0%
b10 *
0-
02
b10 6
#931090000000
1!
1%
1-
12
#931100000000
0!
0%
b11 *
0-
02
b11 6
#931110000000
1!
1%
1-
12
15
#931120000000
0!
0%
b100 *
0-
02
b100 6
#931130000000
1!
1%
1-
12
#931140000000
0!
0%
b101 *
0-
02
b101 6
#931150000000
1!
1%
1-
12
#931160000000
0!
0%
b110 *
0-
02
b110 6
#931170000000
1!
1%
1-
12
#931180000000
0!
0%
b111 *
0-
02
b111 6
#931190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#931200000000
0!
0%
b0 *
0-
02
b0 6
#931210000000
1!
1%
1-
12
#931220000000
0!
0%
b1 *
0-
02
b1 6
#931230000000
1!
1%
1-
12
#931240000000
0!
0%
b10 *
0-
02
b10 6
#931250000000
1!
1%
1-
12
#931260000000
0!
0%
b11 *
0-
02
b11 6
#931270000000
1!
1%
1-
12
15
#931280000000
0!
0%
b100 *
0-
02
b100 6
#931290000000
1!
1%
1-
12
#931300000000
0!
0%
b101 *
0-
02
b101 6
#931310000000
1!
1%
1-
12
#931320000000
0!
0%
b110 *
0-
02
b110 6
#931330000000
1!
1%
1-
12
#931340000000
0!
0%
b111 *
0-
02
b111 6
#931350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#931360000000
0!
0%
b0 *
0-
02
b0 6
#931370000000
1!
1%
1-
12
#931380000000
0!
0%
b1 *
0-
02
b1 6
#931390000000
1!
1%
1-
12
#931400000000
0!
0%
b10 *
0-
02
b10 6
#931410000000
1!
1%
1-
12
#931420000000
0!
0%
b11 *
0-
02
b11 6
#931430000000
1!
1%
1-
12
15
#931440000000
0!
0%
b100 *
0-
02
b100 6
#931450000000
1!
1%
1-
12
#931460000000
0!
0%
b101 *
0-
02
b101 6
#931470000000
1!
1%
1-
12
#931480000000
0!
0%
b110 *
0-
02
b110 6
#931490000000
1!
1%
1-
12
#931500000000
0!
0%
b111 *
0-
02
b111 6
#931510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#931520000000
0!
0%
b0 *
0-
02
b0 6
#931530000000
1!
1%
1-
12
#931540000000
0!
0%
b1 *
0-
02
b1 6
#931550000000
1!
1%
1-
12
#931560000000
0!
0%
b10 *
0-
02
b10 6
#931570000000
1!
1%
1-
12
#931580000000
0!
0%
b11 *
0-
02
b11 6
#931590000000
1!
1%
1-
12
15
#931600000000
0!
0%
b100 *
0-
02
b100 6
#931610000000
1!
1%
1-
12
#931620000000
0!
0%
b101 *
0-
02
b101 6
#931630000000
1!
1%
1-
12
#931640000000
0!
0%
b110 *
0-
02
b110 6
#931650000000
1!
1%
1-
12
#931660000000
0!
0%
b111 *
0-
02
b111 6
#931670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#931680000000
0!
0%
b0 *
0-
02
b0 6
#931690000000
1!
1%
1-
12
#931700000000
0!
0%
b1 *
0-
02
b1 6
#931710000000
1!
1%
1-
12
#931720000000
0!
0%
b10 *
0-
02
b10 6
#931730000000
1!
1%
1-
12
#931740000000
0!
0%
b11 *
0-
02
b11 6
#931750000000
1!
1%
1-
12
15
#931760000000
0!
0%
b100 *
0-
02
b100 6
#931770000000
1!
1%
1-
12
#931780000000
0!
0%
b101 *
0-
02
b101 6
#931790000000
1!
1%
1-
12
#931800000000
0!
0%
b110 *
0-
02
b110 6
#931810000000
1!
1%
1-
12
#931820000000
0!
0%
b111 *
0-
02
b111 6
#931830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#931840000000
0!
0%
b0 *
0-
02
b0 6
#931850000000
1!
1%
1-
12
#931860000000
0!
0%
b1 *
0-
02
b1 6
#931870000000
1!
1%
1-
12
#931880000000
0!
0%
b10 *
0-
02
b10 6
#931890000000
1!
1%
1-
12
#931900000000
0!
0%
b11 *
0-
02
b11 6
#931910000000
1!
1%
1-
12
15
#931920000000
0!
0%
b100 *
0-
02
b100 6
#931930000000
1!
1%
1-
12
#931940000000
0!
0%
b101 *
0-
02
b101 6
#931950000000
1!
1%
1-
12
#931960000000
0!
0%
b110 *
0-
02
b110 6
#931970000000
1!
1%
1-
12
#931980000000
0!
0%
b111 *
0-
02
b111 6
#931990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#932000000000
0!
0%
b0 *
0-
02
b0 6
#932010000000
1!
1%
1-
12
#932020000000
0!
0%
b1 *
0-
02
b1 6
#932030000000
1!
1%
1-
12
#932040000000
0!
0%
b10 *
0-
02
b10 6
#932050000000
1!
1%
1-
12
#932060000000
0!
0%
b11 *
0-
02
b11 6
#932070000000
1!
1%
1-
12
15
#932080000000
0!
0%
b100 *
0-
02
b100 6
#932090000000
1!
1%
1-
12
#932100000000
0!
0%
b101 *
0-
02
b101 6
#932110000000
1!
1%
1-
12
#932120000000
0!
0%
b110 *
0-
02
b110 6
#932130000000
1!
1%
1-
12
#932140000000
0!
0%
b111 *
0-
02
b111 6
#932150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#932160000000
0!
0%
b0 *
0-
02
b0 6
#932170000000
1!
1%
1-
12
#932180000000
0!
0%
b1 *
0-
02
b1 6
#932190000000
1!
1%
1-
12
#932200000000
0!
0%
b10 *
0-
02
b10 6
#932210000000
1!
1%
1-
12
#932220000000
0!
0%
b11 *
0-
02
b11 6
#932230000000
1!
1%
1-
12
15
#932240000000
0!
0%
b100 *
0-
02
b100 6
#932250000000
1!
1%
1-
12
#932260000000
0!
0%
b101 *
0-
02
b101 6
#932270000000
1!
1%
1-
12
#932280000000
0!
0%
b110 *
0-
02
b110 6
#932290000000
1!
1%
1-
12
#932300000000
0!
0%
b111 *
0-
02
b111 6
#932310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#932320000000
0!
0%
b0 *
0-
02
b0 6
#932330000000
1!
1%
1-
12
#932340000000
0!
0%
b1 *
0-
02
b1 6
#932350000000
1!
1%
1-
12
#932360000000
0!
0%
b10 *
0-
02
b10 6
#932370000000
1!
1%
1-
12
#932380000000
0!
0%
b11 *
0-
02
b11 6
#932390000000
1!
1%
1-
12
15
#932400000000
0!
0%
b100 *
0-
02
b100 6
#932410000000
1!
1%
1-
12
#932420000000
0!
0%
b101 *
0-
02
b101 6
#932430000000
1!
1%
1-
12
#932440000000
0!
0%
b110 *
0-
02
b110 6
#932450000000
1!
1%
1-
12
#932460000000
0!
0%
b111 *
0-
02
b111 6
#932470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#932480000000
0!
0%
b0 *
0-
02
b0 6
#932490000000
1!
1%
1-
12
#932500000000
0!
0%
b1 *
0-
02
b1 6
#932510000000
1!
1%
1-
12
#932520000000
0!
0%
b10 *
0-
02
b10 6
#932530000000
1!
1%
1-
12
#932540000000
0!
0%
b11 *
0-
02
b11 6
#932550000000
1!
1%
1-
12
15
#932560000000
0!
0%
b100 *
0-
02
b100 6
#932570000000
1!
1%
1-
12
#932580000000
0!
0%
b101 *
0-
02
b101 6
#932590000000
1!
1%
1-
12
#932600000000
0!
0%
b110 *
0-
02
b110 6
#932610000000
1!
1%
1-
12
#932620000000
0!
0%
b111 *
0-
02
b111 6
#932630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#932640000000
0!
0%
b0 *
0-
02
b0 6
#932650000000
1!
1%
1-
12
#932660000000
0!
0%
b1 *
0-
02
b1 6
#932670000000
1!
1%
1-
12
#932680000000
0!
0%
b10 *
0-
02
b10 6
#932690000000
1!
1%
1-
12
#932700000000
0!
0%
b11 *
0-
02
b11 6
#932710000000
1!
1%
1-
12
15
#932720000000
0!
0%
b100 *
0-
02
b100 6
#932730000000
1!
1%
1-
12
#932740000000
0!
0%
b101 *
0-
02
b101 6
#932750000000
1!
1%
1-
12
#932760000000
0!
0%
b110 *
0-
02
b110 6
#932770000000
1!
1%
1-
12
#932780000000
0!
0%
b111 *
0-
02
b111 6
#932790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#932800000000
0!
0%
b0 *
0-
02
b0 6
#932810000000
1!
1%
1-
12
#932820000000
0!
0%
b1 *
0-
02
b1 6
#932830000000
1!
1%
1-
12
#932840000000
0!
0%
b10 *
0-
02
b10 6
#932850000000
1!
1%
1-
12
#932860000000
0!
0%
b11 *
0-
02
b11 6
#932870000000
1!
1%
1-
12
15
#932880000000
0!
0%
b100 *
0-
02
b100 6
#932890000000
1!
1%
1-
12
#932900000000
0!
0%
b101 *
0-
02
b101 6
#932910000000
1!
1%
1-
12
#932920000000
0!
0%
b110 *
0-
02
b110 6
#932930000000
1!
1%
1-
12
#932940000000
0!
0%
b111 *
0-
02
b111 6
#932950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#932960000000
0!
0%
b0 *
0-
02
b0 6
#932970000000
1!
1%
1-
12
#932980000000
0!
0%
b1 *
0-
02
b1 6
#932990000000
1!
1%
1-
12
#933000000000
0!
0%
b10 *
0-
02
b10 6
#933010000000
1!
1%
1-
12
#933020000000
0!
0%
b11 *
0-
02
b11 6
#933030000000
1!
1%
1-
12
15
#933040000000
0!
0%
b100 *
0-
02
b100 6
#933050000000
1!
1%
1-
12
#933060000000
0!
0%
b101 *
0-
02
b101 6
#933070000000
1!
1%
1-
12
#933080000000
0!
0%
b110 *
0-
02
b110 6
#933090000000
1!
1%
1-
12
#933100000000
0!
0%
b111 *
0-
02
b111 6
#933110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#933120000000
0!
0%
b0 *
0-
02
b0 6
#933130000000
1!
1%
1-
12
#933140000000
0!
0%
b1 *
0-
02
b1 6
#933150000000
1!
1%
1-
12
#933160000000
0!
0%
b10 *
0-
02
b10 6
#933170000000
1!
1%
1-
12
#933180000000
0!
0%
b11 *
0-
02
b11 6
#933190000000
1!
1%
1-
12
15
#933200000000
0!
0%
b100 *
0-
02
b100 6
#933210000000
1!
1%
1-
12
#933220000000
0!
0%
b101 *
0-
02
b101 6
#933230000000
1!
1%
1-
12
#933240000000
0!
0%
b110 *
0-
02
b110 6
#933250000000
1!
1%
1-
12
#933260000000
0!
0%
b111 *
0-
02
b111 6
#933270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#933280000000
0!
0%
b0 *
0-
02
b0 6
#933290000000
1!
1%
1-
12
#933300000000
0!
0%
b1 *
0-
02
b1 6
#933310000000
1!
1%
1-
12
#933320000000
0!
0%
b10 *
0-
02
b10 6
#933330000000
1!
1%
1-
12
#933340000000
0!
0%
b11 *
0-
02
b11 6
#933350000000
1!
1%
1-
12
15
#933360000000
0!
0%
b100 *
0-
02
b100 6
#933370000000
1!
1%
1-
12
#933380000000
0!
0%
b101 *
0-
02
b101 6
#933390000000
1!
1%
1-
12
#933400000000
0!
0%
b110 *
0-
02
b110 6
#933410000000
1!
1%
1-
12
#933420000000
0!
0%
b111 *
0-
02
b111 6
#933430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#933440000000
0!
0%
b0 *
0-
02
b0 6
#933450000000
1!
1%
1-
12
#933460000000
0!
0%
b1 *
0-
02
b1 6
#933470000000
1!
1%
1-
12
#933480000000
0!
0%
b10 *
0-
02
b10 6
#933490000000
1!
1%
1-
12
#933500000000
0!
0%
b11 *
0-
02
b11 6
#933510000000
1!
1%
1-
12
15
#933520000000
0!
0%
b100 *
0-
02
b100 6
#933530000000
1!
1%
1-
12
#933540000000
0!
0%
b101 *
0-
02
b101 6
#933550000000
1!
1%
1-
12
#933560000000
0!
0%
b110 *
0-
02
b110 6
#933570000000
1!
1%
1-
12
#933580000000
0!
0%
b111 *
0-
02
b111 6
#933590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#933600000000
0!
0%
b0 *
0-
02
b0 6
#933610000000
1!
1%
1-
12
#933620000000
0!
0%
b1 *
0-
02
b1 6
#933630000000
1!
1%
1-
12
#933640000000
0!
0%
b10 *
0-
02
b10 6
#933650000000
1!
1%
1-
12
#933660000000
0!
0%
b11 *
0-
02
b11 6
#933670000000
1!
1%
1-
12
15
#933680000000
0!
0%
b100 *
0-
02
b100 6
#933690000000
1!
1%
1-
12
#933700000000
0!
0%
b101 *
0-
02
b101 6
#933710000000
1!
1%
1-
12
#933720000000
0!
0%
b110 *
0-
02
b110 6
#933730000000
1!
1%
1-
12
#933740000000
0!
0%
b111 *
0-
02
b111 6
#933750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#933760000000
0!
0%
b0 *
0-
02
b0 6
#933770000000
1!
1%
1-
12
#933780000000
0!
0%
b1 *
0-
02
b1 6
#933790000000
1!
1%
1-
12
#933800000000
0!
0%
b10 *
0-
02
b10 6
#933810000000
1!
1%
1-
12
#933820000000
0!
0%
b11 *
0-
02
b11 6
#933830000000
1!
1%
1-
12
15
#933840000000
0!
0%
b100 *
0-
02
b100 6
#933850000000
1!
1%
1-
12
#933860000000
0!
0%
b101 *
0-
02
b101 6
#933870000000
1!
1%
1-
12
#933880000000
0!
0%
b110 *
0-
02
b110 6
#933890000000
1!
1%
1-
12
#933900000000
0!
0%
b111 *
0-
02
b111 6
#933910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#933920000000
0!
0%
b0 *
0-
02
b0 6
#933930000000
1!
1%
1-
12
#933940000000
0!
0%
b1 *
0-
02
b1 6
#933950000000
1!
1%
1-
12
#933960000000
0!
0%
b10 *
0-
02
b10 6
#933970000000
1!
1%
1-
12
#933980000000
0!
0%
b11 *
0-
02
b11 6
#933990000000
1!
1%
1-
12
15
#934000000000
0!
0%
b100 *
0-
02
b100 6
#934010000000
1!
1%
1-
12
#934020000000
0!
0%
b101 *
0-
02
b101 6
#934030000000
1!
1%
1-
12
#934040000000
0!
0%
b110 *
0-
02
b110 6
#934050000000
1!
1%
1-
12
#934060000000
0!
0%
b111 *
0-
02
b111 6
#934070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#934080000000
0!
0%
b0 *
0-
02
b0 6
#934090000000
1!
1%
1-
12
#934100000000
0!
0%
b1 *
0-
02
b1 6
#934110000000
1!
1%
1-
12
#934120000000
0!
0%
b10 *
0-
02
b10 6
#934130000000
1!
1%
1-
12
#934140000000
0!
0%
b11 *
0-
02
b11 6
#934150000000
1!
1%
1-
12
15
#934160000000
0!
0%
b100 *
0-
02
b100 6
#934170000000
1!
1%
1-
12
#934180000000
0!
0%
b101 *
0-
02
b101 6
#934190000000
1!
1%
1-
12
#934200000000
0!
0%
b110 *
0-
02
b110 6
#934210000000
1!
1%
1-
12
#934220000000
0!
0%
b111 *
0-
02
b111 6
#934230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#934240000000
0!
0%
b0 *
0-
02
b0 6
#934250000000
1!
1%
1-
12
#934260000000
0!
0%
b1 *
0-
02
b1 6
#934270000000
1!
1%
1-
12
#934280000000
0!
0%
b10 *
0-
02
b10 6
#934290000000
1!
1%
1-
12
#934300000000
0!
0%
b11 *
0-
02
b11 6
#934310000000
1!
1%
1-
12
15
#934320000000
0!
0%
b100 *
0-
02
b100 6
#934330000000
1!
1%
1-
12
#934340000000
0!
0%
b101 *
0-
02
b101 6
#934350000000
1!
1%
1-
12
#934360000000
0!
0%
b110 *
0-
02
b110 6
#934370000000
1!
1%
1-
12
#934380000000
0!
0%
b111 *
0-
02
b111 6
#934390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#934400000000
0!
0%
b0 *
0-
02
b0 6
#934410000000
1!
1%
1-
12
#934420000000
0!
0%
b1 *
0-
02
b1 6
#934430000000
1!
1%
1-
12
#934440000000
0!
0%
b10 *
0-
02
b10 6
#934450000000
1!
1%
1-
12
#934460000000
0!
0%
b11 *
0-
02
b11 6
#934470000000
1!
1%
1-
12
15
#934480000000
0!
0%
b100 *
0-
02
b100 6
#934490000000
1!
1%
1-
12
#934500000000
0!
0%
b101 *
0-
02
b101 6
#934510000000
1!
1%
1-
12
#934520000000
0!
0%
b110 *
0-
02
b110 6
#934530000000
1!
1%
1-
12
#934540000000
0!
0%
b111 *
0-
02
b111 6
#934550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#934560000000
0!
0%
b0 *
0-
02
b0 6
#934570000000
1!
1%
1-
12
#934580000000
0!
0%
b1 *
0-
02
b1 6
#934590000000
1!
1%
1-
12
#934600000000
0!
0%
b10 *
0-
02
b10 6
#934610000000
1!
1%
1-
12
#934620000000
0!
0%
b11 *
0-
02
b11 6
#934630000000
1!
1%
1-
12
15
#934640000000
0!
0%
b100 *
0-
02
b100 6
#934650000000
1!
1%
1-
12
#934660000000
0!
0%
b101 *
0-
02
b101 6
#934670000000
1!
1%
1-
12
#934680000000
0!
0%
b110 *
0-
02
b110 6
#934690000000
1!
1%
1-
12
#934700000000
0!
0%
b111 *
0-
02
b111 6
#934710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#934720000000
0!
0%
b0 *
0-
02
b0 6
#934730000000
1!
1%
1-
12
#934740000000
0!
0%
b1 *
0-
02
b1 6
#934750000000
1!
1%
1-
12
#934760000000
0!
0%
b10 *
0-
02
b10 6
#934770000000
1!
1%
1-
12
#934780000000
0!
0%
b11 *
0-
02
b11 6
#934790000000
1!
1%
1-
12
15
#934800000000
0!
0%
b100 *
0-
02
b100 6
#934810000000
1!
1%
1-
12
#934820000000
0!
0%
b101 *
0-
02
b101 6
#934830000000
1!
1%
1-
12
#934840000000
0!
0%
b110 *
0-
02
b110 6
#934850000000
1!
1%
1-
12
#934860000000
0!
0%
b111 *
0-
02
b111 6
#934870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#934880000000
0!
0%
b0 *
0-
02
b0 6
#934890000000
1!
1%
1-
12
#934900000000
0!
0%
b1 *
0-
02
b1 6
#934910000000
1!
1%
1-
12
#934920000000
0!
0%
b10 *
0-
02
b10 6
#934930000000
1!
1%
1-
12
#934940000000
0!
0%
b11 *
0-
02
b11 6
#934950000000
1!
1%
1-
12
15
#934960000000
0!
0%
b100 *
0-
02
b100 6
#934970000000
1!
1%
1-
12
#934980000000
0!
0%
b101 *
0-
02
b101 6
#934990000000
1!
1%
1-
12
#935000000000
0!
0%
b110 *
0-
02
b110 6
#935010000000
1!
1%
1-
12
#935020000000
0!
0%
b111 *
0-
02
b111 6
#935030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#935040000000
0!
0%
b0 *
0-
02
b0 6
#935050000000
1!
1%
1-
12
#935060000000
0!
0%
b1 *
0-
02
b1 6
#935070000000
1!
1%
1-
12
#935080000000
0!
0%
b10 *
0-
02
b10 6
#935090000000
1!
1%
1-
12
#935100000000
0!
0%
b11 *
0-
02
b11 6
#935110000000
1!
1%
1-
12
15
#935120000000
0!
0%
b100 *
0-
02
b100 6
#935130000000
1!
1%
1-
12
#935140000000
0!
0%
b101 *
0-
02
b101 6
#935150000000
1!
1%
1-
12
#935160000000
0!
0%
b110 *
0-
02
b110 6
#935170000000
1!
1%
1-
12
#935180000000
0!
0%
b111 *
0-
02
b111 6
#935190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#935200000000
0!
0%
b0 *
0-
02
b0 6
#935210000000
1!
1%
1-
12
#935220000000
0!
0%
b1 *
0-
02
b1 6
#935230000000
1!
1%
1-
12
#935240000000
0!
0%
b10 *
0-
02
b10 6
#935250000000
1!
1%
1-
12
#935260000000
0!
0%
b11 *
0-
02
b11 6
#935270000000
1!
1%
1-
12
15
#935280000000
0!
0%
b100 *
0-
02
b100 6
#935290000000
1!
1%
1-
12
#935300000000
0!
0%
b101 *
0-
02
b101 6
#935310000000
1!
1%
1-
12
#935320000000
0!
0%
b110 *
0-
02
b110 6
#935330000000
1!
1%
1-
12
#935340000000
0!
0%
b111 *
0-
02
b111 6
#935350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#935360000000
0!
0%
b0 *
0-
02
b0 6
#935370000000
1!
1%
1-
12
#935380000000
0!
0%
b1 *
0-
02
b1 6
#935390000000
1!
1%
1-
12
#935400000000
0!
0%
b10 *
0-
02
b10 6
#935410000000
1!
1%
1-
12
#935420000000
0!
0%
b11 *
0-
02
b11 6
#935430000000
1!
1%
1-
12
15
#935440000000
0!
0%
b100 *
0-
02
b100 6
#935450000000
1!
1%
1-
12
#935460000000
0!
0%
b101 *
0-
02
b101 6
#935470000000
1!
1%
1-
12
#935480000000
0!
0%
b110 *
0-
02
b110 6
#935490000000
1!
1%
1-
12
#935500000000
0!
0%
b111 *
0-
02
b111 6
#935510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#935520000000
0!
0%
b0 *
0-
02
b0 6
#935530000000
1!
1%
1-
12
#935540000000
0!
0%
b1 *
0-
02
b1 6
#935550000000
1!
1%
1-
12
#935560000000
0!
0%
b10 *
0-
02
b10 6
#935570000000
1!
1%
1-
12
#935580000000
0!
0%
b11 *
0-
02
b11 6
#935590000000
1!
1%
1-
12
15
#935600000000
0!
0%
b100 *
0-
02
b100 6
#935610000000
1!
1%
1-
12
#935620000000
0!
0%
b101 *
0-
02
b101 6
#935630000000
1!
1%
1-
12
#935640000000
0!
0%
b110 *
0-
02
b110 6
#935650000000
1!
1%
1-
12
#935660000000
0!
0%
b111 *
0-
02
b111 6
#935670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#935680000000
0!
0%
b0 *
0-
02
b0 6
#935690000000
1!
1%
1-
12
#935700000000
0!
0%
b1 *
0-
02
b1 6
#935710000000
1!
1%
1-
12
#935720000000
0!
0%
b10 *
0-
02
b10 6
#935730000000
1!
1%
1-
12
#935740000000
0!
0%
b11 *
0-
02
b11 6
#935750000000
1!
1%
1-
12
15
#935760000000
0!
0%
b100 *
0-
02
b100 6
#935770000000
1!
1%
1-
12
#935780000000
0!
0%
b101 *
0-
02
b101 6
#935790000000
1!
1%
1-
12
#935800000000
0!
0%
b110 *
0-
02
b110 6
#935810000000
1!
1%
1-
12
#935820000000
0!
0%
b111 *
0-
02
b111 6
#935830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#935840000000
0!
0%
b0 *
0-
02
b0 6
#935850000000
1!
1%
1-
12
#935860000000
0!
0%
b1 *
0-
02
b1 6
#935870000000
1!
1%
1-
12
#935880000000
0!
0%
b10 *
0-
02
b10 6
#935890000000
1!
1%
1-
12
#935900000000
0!
0%
b11 *
0-
02
b11 6
#935910000000
1!
1%
1-
12
15
#935920000000
0!
0%
b100 *
0-
02
b100 6
#935930000000
1!
1%
1-
12
#935940000000
0!
0%
b101 *
0-
02
b101 6
#935950000000
1!
1%
1-
12
#935960000000
0!
0%
b110 *
0-
02
b110 6
#935970000000
1!
1%
1-
12
#935980000000
0!
0%
b111 *
0-
02
b111 6
#935990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#936000000000
0!
0%
b0 *
0-
02
b0 6
#936010000000
1!
1%
1-
12
#936020000000
0!
0%
b1 *
0-
02
b1 6
#936030000000
1!
1%
1-
12
#936040000000
0!
0%
b10 *
0-
02
b10 6
#936050000000
1!
1%
1-
12
#936060000000
0!
0%
b11 *
0-
02
b11 6
#936070000000
1!
1%
1-
12
15
#936080000000
0!
0%
b100 *
0-
02
b100 6
#936090000000
1!
1%
1-
12
#936100000000
0!
0%
b101 *
0-
02
b101 6
#936110000000
1!
1%
1-
12
#936120000000
0!
0%
b110 *
0-
02
b110 6
#936130000000
1!
1%
1-
12
#936140000000
0!
0%
b111 *
0-
02
b111 6
#936150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#936160000000
0!
0%
b0 *
0-
02
b0 6
#936170000000
1!
1%
1-
12
#936180000000
0!
0%
b1 *
0-
02
b1 6
#936190000000
1!
1%
1-
12
#936200000000
0!
0%
b10 *
0-
02
b10 6
#936210000000
1!
1%
1-
12
#936220000000
0!
0%
b11 *
0-
02
b11 6
#936230000000
1!
1%
1-
12
15
#936240000000
0!
0%
b100 *
0-
02
b100 6
#936250000000
1!
1%
1-
12
#936260000000
0!
0%
b101 *
0-
02
b101 6
#936270000000
1!
1%
1-
12
#936280000000
0!
0%
b110 *
0-
02
b110 6
#936290000000
1!
1%
1-
12
#936300000000
0!
0%
b111 *
0-
02
b111 6
#936310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#936320000000
0!
0%
b0 *
0-
02
b0 6
#936330000000
1!
1%
1-
12
#936340000000
0!
0%
b1 *
0-
02
b1 6
#936350000000
1!
1%
1-
12
#936360000000
0!
0%
b10 *
0-
02
b10 6
#936370000000
1!
1%
1-
12
#936380000000
0!
0%
b11 *
0-
02
b11 6
#936390000000
1!
1%
1-
12
15
#936400000000
0!
0%
b100 *
0-
02
b100 6
#936410000000
1!
1%
1-
12
#936420000000
0!
0%
b101 *
0-
02
b101 6
#936430000000
1!
1%
1-
12
#936440000000
0!
0%
b110 *
0-
02
b110 6
#936450000000
1!
1%
1-
12
#936460000000
0!
0%
b111 *
0-
02
b111 6
#936470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#936480000000
0!
0%
b0 *
0-
02
b0 6
#936490000000
1!
1%
1-
12
#936500000000
0!
0%
b1 *
0-
02
b1 6
#936510000000
1!
1%
1-
12
#936520000000
0!
0%
b10 *
0-
02
b10 6
#936530000000
1!
1%
1-
12
#936540000000
0!
0%
b11 *
0-
02
b11 6
#936550000000
1!
1%
1-
12
15
#936560000000
0!
0%
b100 *
0-
02
b100 6
#936570000000
1!
1%
1-
12
#936580000000
0!
0%
b101 *
0-
02
b101 6
#936590000000
1!
1%
1-
12
#936600000000
0!
0%
b110 *
0-
02
b110 6
#936610000000
1!
1%
1-
12
#936620000000
0!
0%
b111 *
0-
02
b111 6
#936630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#936640000000
0!
0%
b0 *
0-
02
b0 6
#936650000000
1!
1%
1-
12
#936660000000
0!
0%
b1 *
0-
02
b1 6
#936670000000
1!
1%
1-
12
#936680000000
0!
0%
b10 *
0-
02
b10 6
#936690000000
1!
1%
1-
12
#936700000000
0!
0%
b11 *
0-
02
b11 6
#936710000000
1!
1%
1-
12
15
#936720000000
0!
0%
b100 *
0-
02
b100 6
#936730000000
1!
1%
1-
12
#936740000000
0!
0%
b101 *
0-
02
b101 6
#936750000000
1!
1%
1-
12
#936760000000
0!
0%
b110 *
0-
02
b110 6
#936770000000
1!
1%
1-
12
#936780000000
0!
0%
b111 *
0-
02
b111 6
#936790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#936800000000
0!
0%
b0 *
0-
02
b0 6
#936810000000
1!
1%
1-
12
#936820000000
0!
0%
b1 *
0-
02
b1 6
#936830000000
1!
1%
1-
12
#936840000000
0!
0%
b10 *
0-
02
b10 6
#936850000000
1!
1%
1-
12
#936860000000
0!
0%
b11 *
0-
02
b11 6
#936870000000
1!
1%
1-
12
15
#936880000000
0!
0%
b100 *
0-
02
b100 6
#936890000000
1!
1%
1-
12
#936900000000
0!
0%
b101 *
0-
02
b101 6
#936910000000
1!
1%
1-
12
#936920000000
0!
0%
b110 *
0-
02
b110 6
#936930000000
1!
1%
1-
12
#936940000000
0!
0%
b111 *
0-
02
b111 6
#936950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#936960000000
0!
0%
b0 *
0-
02
b0 6
#936970000000
1!
1%
1-
12
#936980000000
0!
0%
b1 *
0-
02
b1 6
#936990000000
1!
1%
1-
12
#937000000000
0!
0%
b10 *
0-
02
b10 6
#937010000000
1!
1%
1-
12
#937020000000
0!
0%
b11 *
0-
02
b11 6
#937030000000
1!
1%
1-
12
15
#937040000000
0!
0%
b100 *
0-
02
b100 6
#937050000000
1!
1%
1-
12
#937060000000
0!
0%
b101 *
0-
02
b101 6
#937070000000
1!
1%
1-
12
#937080000000
0!
0%
b110 *
0-
02
b110 6
#937090000000
1!
1%
1-
12
#937100000000
0!
0%
b111 *
0-
02
b111 6
#937110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#937120000000
0!
0%
b0 *
0-
02
b0 6
#937130000000
1!
1%
1-
12
#937140000000
0!
0%
b1 *
0-
02
b1 6
#937150000000
1!
1%
1-
12
#937160000000
0!
0%
b10 *
0-
02
b10 6
#937170000000
1!
1%
1-
12
#937180000000
0!
0%
b11 *
0-
02
b11 6
#937190000000
1!
1%
1-
12
15
#937200000000
0!
0%
b100 *
0-
02
b100 6
#937210000000
1!
1%
1-
12
#937220000000
0!
0%
b101 *
0-
02
b101 6
#937230000000
1!
1%
1-
12
#937240000000
0!
0%
b110 *
0-
02
b110 6
#937250000000
1!
1%
1-
12
#937260000000
0!
0%
b111 *
0-
02
b111 6
#937270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#937280000000
0!
0%
b0 *
0-
02
b0 6
#937290000000
1!
1%
1-
12
#937300000000
0!
0%
b1 *
0-
02
b1 6
#937310000000
1!
1%
1-
12
#937320000000
0!
0%
b10 *
0-
02
b10 6
#937330000000
1!
1%
1-
12
#937340000000
0!
0%
b11 *
0-
02
b11 6
#937350000000
1!
1%
1-
12
15
#937360000000
0!
0%
b100 *
0-
02
b100 6
#937370000000
1!
1%
1-
12
#937380000000
0!
0%
b101 *
0-
02
b101 6
#937390000000
1!
1%
1-
12
#937400000000
0!
0%
b110 *
0-
02
b110 6
#937410000000
1!
1%
1-
12
#937420000000
0!
0%
b111 *
0-
02
b111 6
#937430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#937440000000
0!
0%
b0 *
0-
02
b0 6
#937450000000
1!
1%
1-
12
#937460000000
0!
0%
b1 *
0-
02
b1 6
#937470000000
1!
1%
1-
12
#937480000000
0!
0%
b10 *
0-
02
b10 6
#937490000000
1!
1%
1-
12
#937500000000
0!
0%
b11 *
0-
02
b11 6
#937510000000
1!
1%
1-
12
15
#937520000000
0!
0%
b100 *
0-
02
b100 6
#937530000000
1!
1%
1-
12
#937540000000
0!
0%
b101 *
0-
02
b101 6
#937550000000
1!
1%
1-
12
#937560000000
0!
0%
b110 *
0-
02
b110 6
#937570000000
1!
1%
1-
12
#937580000000
0!
0%
b111 *
0-
02
b111 6
#937590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#937600000000
0!
0%
b0 *
0-
02
b0 6
#937610000000
1!
1%
1-
12
#937620000000
0!
0%
b1 *
0-
02
b1 6
#937630000000
1!
1%
1-
12
#937640000000
0!
0%
b10 *
0-
02
b10 6
#937650000000
1!
1%
1-
12
#937660000000
0!
0%
b11 *
0-
02
b11 6
#937670000000
1!
1%
1-
12
15
#937680000000
0!
0%
b100 *
0-
02
b100 6
#937690000000
1!
1%
1-
12
#937700000000
0!
0%
b101 *
0-
02
b101 6
#937710000000
1!
1%
1-
12
#937720000000
0!
0%
b110 *
0-
02
b110 6
#937730000000
1!
1%
1-
12
#937740000000
0!
0%
b111 *
0-
02
b111 6
#937750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#937760000000
0!
0%
b0 *
0-
02
b0 6
#937770000000
1!
1%
1-
12
#937780000000
0!
0%
b1 *
0-
02
b1 6
#937790000000
1!
1%
1-
12
#937800000000
0!
0%
b10 *
0-
02
b10 6
#937810000000
1!
1%
1-
12
#937820000000
0!
0%
b11 *
0-
02
b11 6
#937830000000
1!
1%
1-
12
15
#937840000000
0!
0%
b100 *
0-
02
b100 6
#937850000000
1!
1%
1-
12
#937860000000
0!
0%
b101 *
0-
02
b101 6
#937870000000
1!
1%
1-
12
#937880000000
0!
0%
b110 *
0-
02
b110 6
#937890000000
1!
1%
1-
12
#937900000000
0!
0%
b111 *
0-
02
b111 6
#937910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#937920000000
0!
0%
b0 *
0-
02
b0 6
#937930000000
1!
1%
1-
12
#937940000000
0!
0%
b1 *
0-
02
b1 6
#937950000000
1!
1%
1-
12
#937960000000
0!
0%
b10 *
0-
02
b10 6
#937970000000
1!
1%
1-
12
#937980000000
0!
0%
b11 *
0-
02
b11 6
#937990000000
1!
1%
1-
12
15
#938000000000
0!
0%
b100 *
0-
02
b100 6
#938010000000
1!
1%
1-
12
#938020000000
0!
0%
b101 *
0-
02
b101 6
#938030000000
1!
1%
1-
12
#938040000000
0!
0%
b110 *
0-
02
b110 6
#938050000000
1!
1%
1-
12
#938060000000
0!
0%
b111 *
0-
02
b111 6
#938070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#938080000000
0!
0%
b0 *
0-
02
b0 6
#938090000000
1!
1%
1-
12
#938100000000
0!
0%
b1 *
0-
02
b1 6
#938110000000
1!
1%
1-
12
#938120000000
0!
0%
b10 *
0-
02
b10 6
#938130000000
1!
1%
1-
12
#938140000000
0!
0%
b11 *
0-
02
b11 6
#938150000000
1!
1%
1-
12
15
#938160000000
0!
0%
b100 *
0-
02
b100 6
#938170000000
1!
1%
1-
12
#938180000000
0!
0%
b101 *
0-
02
b101 6
#938190000000
1!
1%
1-
12
#938200000000
0!
0%
b110 *
0-
02
b110 6
#938210000000
1!
1%
1-
12
#938220000000
0!
0%
b111 *
0-
02
b111 6
#938230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#938240000000
0!
0%
b0 *
0-
02
b0 6
#938250000000
1!
1%
1-
12
#938260000000
0!
0%
b1 *
0-
02
b1 6
#938270000000
1!
1%
1-
12
#938280000000
0!
0%
b10 *
0-
02
b10 6
#938290000000
1!
1%
1-
12
#938300000000
0!
0%
b11 *
0-
02
b11 6
#938310000000
1!
1%
1-
12
15
#938320000000
0!
0%
b100 *
0-
02
b100 6
#938330000000
1!
1%
1-
12
#938340000000
0!
0%
b101 *
0-
02
b101 6
#938350000000
1!
1%
1-
12
#938360000000
0!
0%
b110 *
0-
02
b110 6
#938370000000
1!
1%
1-
12
#938380000000
0!
0%
b111 *
0-
02
b111 6
#938390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#938400000000
0!
0%
b0 *
0-
02
b0 6
#938410000000
1!
1%
1-
12
#938420000000
0!
0%
b1 *
0-
02
b1 6
#938430000000
1!
1%
1-
12
#938440000000
0!
0%
b10 *
0-
02
b10 6
#938450000000
1!
1%
1-
12
#938460000000
0!
0%
b11 *
0-
02
b11 6
#938470000000
1!
1%
1-
12
15
#938480000000
0!
0%
b100 *
0-
02
b100 6
#938490000000
1!
1%
1-
12
#938500000000
0!
0%
b101 *
0-
02
b101 6
#938510000000
1!
1%
1-
12
#938520000000
0!
0%
b110 *
0-
02
b110 6
#938530000000
1!
1%
1-
12
#938540000000
0!
0%
b111 *
0-
02
b111 6
#938550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#938560000000
0!
0%
b0 *
0-
02
b0 6
#938570000000
1!
1%
1-
12
#938580000000
0!
0%
b1 *
0-
02
b1 6
#938590000000
1!
1%
1-
12
#938600000000
0!
0%
b10 *
0-
02
b10 6
#938610000000
1!
1%
1-
12
#938620000000
0!
0%
b11 *
0-
02
b11 6
#938630000000
1!
1%
1-
12
15
#938640000000
0!
0%
b100 *
0-
02
b100 6
#938650000000
1!
1%
1-
12
#938660000000
0!
0%
b101 *
0-
02
b101 6
#938670000000
1!
1%
1-
12
#938680000000
0!
0%
b110 *
0-
02
b110 6
#938690000000
1!
1%
1-
12
#938700000000
0!
0%
b111 *
0-
02
b111 6
#938710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#938720000000
0!
0%
b0 *
0-
02
b0 6
#938730000000
1!
1%
1-
12
#938740000000
0!
0%
b1 *
0-
02
b1 6
#938750000000
1!
1%
1-
12
#938760000000
0!
0%
b10 *
0-
02
b10 6
#938770000000
1!
1%
1-
12
#938780000000
0!
0%
b11 *
0-
02
b11 6
#938790000000
1!
1%
1-
12
15
#938800000000
0!
0%
b100 *
0-
02
b100 6
#938810000000
1!
1%
1-
12
#938820000000
0!
0%
b101 *
0-
02
b101 6
#938830000000
1!
1%
1-
12
#938840000000
0!
0%
b110 *
0-
02
b110 6
#938850000000
1!
1%
1-
12
#938860000000
0!
0%
b111 *
0-
02
b111 6
#938870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#938880000000
0!
0%
b0 *
0-
02
b0 6
#938890000000
1!
1%
1-
12
#938900000000
0!
0%
b1 *
0-
02
b1 6
#938910000000
1!
1%
1-
12
#938920000000
0!
0%
b10 *
0-
02
b10 6
#938930000000
1!
1%
1-
12
#938940000000
0!
0%
b11 *
0-
02
b11 6
#938950000000
1!
1%
1-
12
15
#938960000000
0!
0%
b100 *
0-
02
b100 6
#938970000000
1!
1%
1-
12
#938980000000
0!
0%
b101 *
0-
02
b101 6
#938990000000
1!
1%
1-
12
#939000000000
0!
0%
b110 *
0-
02
b110 6
#939010000000
1!
1%
1-
12
#939020000000
0!
0%
b111 *
0-
02
b111 6
#939030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#939040000000
0!
0%
b0 *
0-
02
b0 6
#939050000000
1!
1%
1-
12
#939060000000
0!
0%
b1 *
0-
02
b1 6
#939070000000
1!
1%
1-
12
#939080000000
0!
0%
b10 *
0-
02
b10 6
#939090000000
1!
1%
1-
12
#939100000000
0!
0%
b11 *
0-
02
b11 6
#939110000000
1!
1%
1-
12
15
#939120000000
0!
0%
b100 *
0-
02
b100 6
#939130000000
1!
1%
1-
12
#939140000000
0!
0%
b101 *
0-
02
b101 6
#939150000000
1!
1%
1-
12
#939160000000
0!
0%
b110 *
0-
02
b110 6
#939170000000
1!
1%
1-
12
#939180000000
0!
0%
b111 *
0-
02
b111 6
#939190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#939200000000
0!
0%
b0 *
0-
02
b0 6
#939210000000
1!
1%
1-
12
#939220000000
0!
0%
b1 *
0-
02
b1 6
#939230000000
1!
1%
1-
12
#939240000000
0!
0%
b10 *
0-
02
b10 6
#939250000000
1!
1%
1-
12
#939260000000
0!
0%
b11 *
0-
02
b11 6
#939270000000
1!
1%
1-
12
15
#939280000000
0!
0%
b100 *
0-
02
b100 6
#939290000000
1!
1%
1-
12
#939300000000
0!
0%
b101 *
0-
02
b101 6
#939310000000
1!
1%
1-
12
#939320000000
0!
0%
b110 *
0-
02
b110 6
#939330000000
1!
1%
1-
12
#939340000000
0!
0%
b111 *
0-
02
b111 6
#939350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#939360000000
0!
0%
b0 *
0-
02
b0 6
#939370000000
1!
1%
1-
12
#939380000000
0!
0%
b1 *
0-
02
b1 6
#939390000000
1!
1%
1-
12
#939400000000
0!
0%
b10 *
0-
02
b10 6
#939410000000
1!
1%
1-
12
#939420000000
0!
0%
b11 *
0-
02
b11 6
#939430000000
1!
1%
1-
12
15
#939440000000
0!
0%
b100 *
0-
02
b100 6
#939450000000
1!
1%
1-
12
#939460000000
0!
0%
b101 *
0-
02
b101 6
#939470000000
1!
1%
1-
12
#939480000000
0!
0%
b110 *
0-
02
b110 6
#939490000000
1!
1%
1-
12
#939500000000
0!
0%
b111 *
0-
02
b111 6
#939510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#939520000000
0!
0%
b0 *
0-
02
b0 6
#939530000000
1!
1%
1-
12
#939540000000
0!
0%
b1 *
0-
02
b1 6
#939550000000
1!
1%
1-
12
#939560000000
0!
0%
b10 *
0-
02
b10 6
#939570000000
1!
1%
1-
12
#939580000000
0!
0%
b11 *
0-
02
b11 6
#939590000000
1!
1%
1-
12
15
#939600000000
0!
0%
b100 *
0-
02
b100 6
#939610000000
1!
1%
1-
12
#939620000000
0!
0%
b101 *
0-
02
b101 6
#939630000000
1!
1%
1-
12
#939640000000
0!
0%
b110 *
0-
02
b110 6
#939650000000
1!
1%
1-
12
#939660000000
0!
0%
b111 *
0-
02
b111 6
#939670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#939680000000
0!
0%
b0 *
0-
02
b0 6
#939690000000
1!
1%
1-
12
#939700000000
0!
0%
b1 *
0-
02
b1 6
#939710000000
1!
1%
1-
12
#939720000000
0!
0%
b10 *
0-
02
b10 6
#939730000000
1!
1%
1-
12
#939740000000
0!
0%
b11 *
0-
02
b11 6
#939750000000
1!
1%
1-
12
15
#939760000000
0!
0%
b100 *
0-
02
b100 6
#939770000000
1!
1%
1-
12
#939780000000
0!
0%
b101 *
0-
02
b101 6
#939790000000
1!
1%
1-
12
#939800000000
0!
0%
b110 *
0-
02
b110 6
#939810000000
1!
1%
1-
12
#939820000000
0!
0%
b111 *
0-
02
b111 6
#939830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#939840000000
0!
0%
b0 *
0-
02
b0 6
#939850000000
1!
1%
1-
12
#939860000000
0!
0%
b1 *
0-
02
b1 6
#939870000000
1!
1%
1-
12
#939880000000
0!
0%
b10 *
0-
02
b10 6
#939890000000
1!
1%
1-
12
#939900000000
0!
0%
b11 *
0-
02
b11 6
#939910000000
1!
1%
1-
12
15
#939920000000
0!
0%
b100 *
0-
02
b100 6
#939930000000
1!
1%
1-
12
#939940000000
0!
0%
b101 *
0-
02
b101 6
#939950000000
1!
1%
1-
12
#939960000000
0!
0%
b110 *
0-
02
b110 6
#939970000000
1!
1%
1-
12
#939980000000
0!
0%
b111 *
0-
02
b111 6
#939990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#940000000000
0!
0%
b0 *
0-
02
b0 6
#940010000000
1!
1%
1-
12
#940020000000
0!
0%
b1 *
0-
02
b1 6
#940030000000
1!
1%
1-
12
#940040000000
0!
0%
b10 *
0-
02
b10 6
#940050000000
1!
1%
1-
12
#940060000000
0!
0%
b11 *
0-
02
b11 6
#940070000000
1!
1%
1-
12
15
#940080000000
0!
0%
b100 *
0-
02
b100 6
#940090000000
1!
1%
1-
12
#940100000000
0!
0%
b101 *
0-
02
b101 6
#940110000000
1!
1%
1-
12
#940120000000
0!
0%
b110 *
0-
02
b110 6
#940130000000
1!
1%
1-
12
#940140000000
0!
0%
b111 *
0-
02
b111 6
#940150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#940160000000
0!
0%
b0 *
0-
02
b0 6
#940170000000
1!
1%
1-
12
#940180000000
0!
0%
b1 *
0-
02
b1 6
#940190000000
1!
1%
1-
12
#940200000000
0!
0%
b10 *
0-
02
b10 6
#940210000000
1!
1%
1-
12
#940220000000
0!
0%
b11 *
0-
02
b11 6
#940230000000
1!
1%
1-
12
15
#940240000000
0!
0%
b100 *
0-
02
b100 6
#940250000000
1!
1%
1-
12
#940260000000
0!
0%
b101 *
0-
02
b101 6
#940270000000
1!
1%
1-
12
#940280000000
0!
0%
b110 *
0-
02
b110 6
#940290000000
1!
1%
1-
12
#940300000000
0!
0%
b111 *
0-
02
b111 6
#940310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#940320000000
0!
0%
b0 *
0-
02
b0 6
#940330000000
1!
1%
1-
12
#940340000000
0!
0%
b1 *
0-
02
b1 6
#940350000000
1!
1%
1-
12
#940360000000
0!
0%
b10 *
0-
02
b10 6
#940370000000
1!
1%
1-
12
#940380000000
0!
0%
b11 *
0-
02
b11 6
#940390000000
1!
1%
1-
12
15
#940400000000
0!
0%
b100 *
0-
02
b100 6
#940410000000
1!
1%
1-
12
#940420000000
0!
0%
b101 *
0-
02
b101 6
#940430000000
1!
1%
1-
12
#940440000000
0!
0%
b110 *
0-
02
b110 6
#940450000000
1!
1%
1-
12
#940460000000
0!
0%
b111 *
0-
02
b111 6
#940470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#940480000000
0!
0%
b0 *
0-
02
b0 6
#940490000000
1!
1%
1-
12
#940500000000
0!
0%
b1 *
0-
02
b1 6
#940510000000
1!
1%
1-
12
#940520000000
0!
0%
b10 *
0-
02
b10 6
#940530000000
1!
1%
1-
12
#940540000000
0!
0%
b11 *
0-
02
b11 6
#940550000000
1!
1%
1-
12
15
#940560000000
0!
0%
b100 *
0-
02
b100 6
#940570000000
1!
1%
1-
12
#940580000000
0!
0%
b101 *
0-
02
b101 6
#940590000000
1!
1%
1-
12
#940600000000
0!
0%
b110 *
0-
02
b110 6
#940610000000
1!
1%
1-
12
#940620000000
0!
0%
b111 *
0-
02
b111 6
#940630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#940640000000
0!
0%
b0 *
0-
02
b0 6
#940650000000
1!
1%
1-
12
#940660000000
0!
0%
b1 *
0-
02
b1 6
#940670000000
1!
1%
1-
12
#940680000000
0!
0%
b10 *
0-
02
b10 6
#940690000000
1!
1%
1-
12
#940700000000
0!
0%
b11 *
0-
02
b11 6
#940710000000
1!
1%
1-
12
15
#940720000000
0!
0%
b100 *
0-
02
b100 6
#940730000000
1!
1%
1-
12
#940740000000
0!
0%
b101 *
0-
02
b101 6
#940750000000
1!
1%
1-
12
#940760000000
0!
0%
b110 *
0-
02
b110 6
#940770000000
1!
1%
1-
12
#940780000000
0!
0%
b111 *
0-
02
b111 6
#940790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#940800000000
0!
0%
b0 *
0-
02
b0 6
#940810000000
1!
1%
1-
12
#940820000000
0!
0%
b1 *
0-
02
b1 6
#940830000000
1!
1%
1-
12
#940840000000
0!
0%
b10 *
0-
02
b10 6
#940850000000
1!
1%
1-
12
#940860000000
0!
0%
b11 *
0-
02
b11 6
#940870000000
1!
1%
1-
12
15
#940880000000
0!
0%
b100 *
0-
02
b100 6
#940890000000
1!
1%
1-
12
#940900000000
0!
0%
b101 *
0-
02
b101 6
#940910000000
1!
1%
1-
12
#940920000000
0!
0%
b110 *
0-
02
b110 6
#940930000000
1!
1%
1-
12
#940940000000
0!
0%
b111 *
0-
02
b111 6
#940950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#940960000000
0!
0%
b0 *
0-
02
b0 6
#940970000000
1!
1%
1-
12
#940980000000
0!
0%
b1 *
0-
02
b1 6
#940990000000
1!
1%
1-
12
#941000000000
0!
0%
b10 *
0-
02
b10 6
#941010000000
1!
1%
1-
12
#941020000000
0!
0%
b11 *
0-
02
b11 6
#941030000000
1!
1%
1-
12
15
#941040000000
0!
0%
b100 *
0-
02
b100 6
#941050000000
1!
1%
1-
12
#941060000000
0!
0%
b101 *
0-
02
b101 6
#941070000000
1!
1%
1-
12
#941080000000
0!
0%
b110 *
0-
02
b110 6
#941090000000
1!
1%
1-
12
#941100000000
0!
0%
b111 *
0-
02
b111 6
#941110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#941120000000
0!
0%
b0 *
0-
02
b0 6
#941130000000
1!
1%
1-
12
#941140000000
0!
0%
b1 *
0-
02
b1 6
#941150000000
1!
1%
1-
12
#941160000000
0!
0%
b10 *
0-
02
b10 6
#941170000000
1!
1%
1-
12
#941180000000
0!
0%
b11 *
0-
02
b11 6
#941190000000
1!
1%
1-
12
15
#941200000000
0!
0%
b100 *
0-
02
b100 6
#941210000000
1!
1%
1-
12
#941220000000
0!
0%
b101 *
0-
02
b101 6
#941230000000
1!
1%
1-
12
#941240000000
0!
0%
b110 *
0-
02
b110 6
#941250000000
1!
1%
1-
12
#941260000000
0!
0%
b111 *
0-
02
b111 6
#941270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#941280000000
0!
0%
b0 *
0-
02
b0 6
#941290000000
1!
1%
1-
12
#941300000000
0!
0%
b1 *
0-
02
b1 6
#941310000000
1!
1%
1-
12
#941320000000
0!
0%
b10 *
0-
02
b10 6
#941330000000
1!
1%
1-
12
#941340000000
0!
0%
b11 *
0-
02
b11 6
#941350000000
1!
1%
1-
12
15
#941360000000
0!
0%
b100 *
0-
02
b100 6
#941370000000
1!
1%
1-
12
#941380000000
0!
0%
b101 *
0-
02
b101 6
#941390000000
1!
1%
1-
12
#941400000000
0!
0%
b110 *
0-
02
b110 6
#941410000000
1!
1%
1-
12
#941420000000
0!
0%
b111 *
0-
02
b111 6
#941430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#941440000000
0!
0%
b0 *
0-
02
b0 6
#941450000000
1!
1%
1-
12
#941460000000
0!
0%
b1 *
0-
02
b1 6
#941470000000
1!
1%
1-
12
#941480000000
0!
0%
b10 *
0-
02
b10 6
#941490000000
1!
1%
1-
12
#941500000000
0!
0%
b11 *
0-
02
b11 6
#941510000000
1!
1%
1-
12
15
#941520000000
0!
0%
b100 *
0-
02
b100 6
#941530000000
1!
1%
1-
12
#941540000000
0!
0%
b101 *
0-
02
b101 6
#941550000000
1!
1%
1-
12
#941560000000
0!
0%
b110 *
0-
02
b110 6
#941570000000
1!
1%
1-
12
#941580000000
0!
0%
b111 *
0-
02
b111 6
#941590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#941600000000
0!
0%
b0 *
0-
02
b0 6
#941610000000
1!
1%
1-
12
#941620000000
0!
0%
b1 *
0-
02
b1 6
#941630000000
1!
1%
1-
12
#941640000000
0!
0%
b10 *
0-
02
b10 6
#941650000000
1!
1%
1-
12
#941660000000
0!
0%
b11 *
0-
02
b11 6
#941670000000
1!
1%
1-
12
15
#941680000000
0!
0%
b100 *
0-
02
b100 6
#941690000000
1!
1%
1-
12
#941700000000
0!
0%
b101 *
0-
02
b101 6
#941710000000
1!
1%
1-
12
#941720000000
0!
0%
b110 *
0-
02
b110 6
#941730000000
1!
1%
1-
12
#941740000000
0!
0%
b111 *
0-
02
b111 6
#941750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#941760000000
0!
0%
b0 *
0-
02
b0 6
#941770000000
1!
1%
1-
12
#941780000000
0!
0%
b1 *
0-
02
b1 6
#941790000000
1!
1%
1-
12
#941800000000
0!
0%
b10 *
0-
02
b10 6
#941810000000
1!
1%
1-
12
#941820000000
0!
0%
b11 *
0-
02
b11 6
#941830000000
1!
1%
1-
12
15
#941840000000
0!
0%
b100 *
0-
02
b100 6
#941850000000
1!
1%
1-
12
#941860000000
0!
0%
b101 *
0-
02
b101 6
#941870000000
1!
1%
1-
12
#941880000000
0!
0%
b110 *
0-
02
b110 6
#941890000000
1!
1%
1-
12
#941900000000
0!
0%
b111 *
0-
02
b111 6
#941910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#941920000000
0!
0%
b0 *
0-
02
b0 6
#941930000000
1!
1%
1-
12
#941940000000
0!
0%
b1 *
0-
02
b1 6
#941950000000
1!
1%
1-
12
#941960000000
0!
0%
b10 *
0-
02
b10 6
#941970000000
1!
1%
1-
12
#941980000000
0!
0%
b11 *
0-
02
b11 6
#941990000000
1!
1%
1-
12
15
#942000000000
0!
0%
b100 *
0-
02
b100 6
#942010000000
1!
1%
1-
12
#942020000000
0!
0%
b101 *
0-
02
b101 6
#942030000000
1!
1%
1-
12
#942040000000
0!
0%
b110 *
0-
02
b110 6
#942050000000
1!
1%
1-
12
#942060000000
0!
0%
b111 *
0-
02
b111 6
#942070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#942080000000
0!
0%
b0 *
0-
02
b0 6
#942090000000
1!
1%
1-
12
#942100000000
0!
0%
b1 *
0-
02
b1 6
#942110000000
1!
1%
1-
12
#942120000000
0!
0%
b10 *
0-
02
b10 6
#942130000000
1!
1%
1-
12
#942140000000
0!
0%
b11 *
0-
02
b11 6
#942150000000
1!
1%
1-
12
15
#942160000000
0!
0%
b100 *
0-
02
b100 6
#942170000000
1!
1%
1-
12
#942180000000
0!
0%
b101 *
0-
02
b101 6
#942190000000
1!
1%
1-
12
#942200000000
0!
0%
b110 *
0-
02
b110 6
#942210000000
1!
1%
1-
12
#942220000000
0!
0%
b111 *
0-
02
b111 6
#942230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#942240000000
0!
0%
b0 *
0-
02
b0 6
#942250000000
1!
1%
1-
12
#942260000000
0!
0%
b1 *
0-
02
b1 6
#942270000000
1!
1%
1-
12
#942280000000
0!
0%
b10 *
0-
02
b10 6
#942290000000
1!
1%
1-
12
#942300000000
0!
0%
b11 *
0-
02
b11 6
#942310000000
1!
1%
1-
12
15
#942320000000
0!
0%
b100 *
0-
02
b100 6
#942330000000
1!
1%
1-
12
#942340000000
0!
0%
b101 *
0-
02
b101 6
#942350000000
1!
1%
1-
12
#942360000000
0!
0%
b110 *
0-
02
b110 6
#942370000000
1!
1%
1-
12
#942380000000
0!
0%
b111 *
0-
02
b111 6
#942390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#942400000000
0!
0%
b0 *
0-
02
b0 6
#942410000000
1!
1%
1-
12
#942420000000
0!
0%
b1 *
0-
02
b1 6
#942430000000
1!
1%
1-
12
#942440000000
0!
0%
b10 *
0-
02
b10 6
#942450000000
1!
1%
1-
12
#942460000000
0!
0%
b11 *
0-
02
b11 6
#942470000000
1!
1%
1-
12
15
#942480000000
0!
0%
b100 *
0-
02
b100 6
#942490000000
1!
1%
1-
12
#942500000000
0!
0%
b101 *
0-
02
b101 6
#942510000000
1!
1%
1-
12
#942520000000
0!
0%
b110 *
0-
02
b110 6
#942530000000
1!
1%
1-
12
#942540000000
0!
0%
b111 *
0-
02
b111 6
#942550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#942560000000
0!
0%
b0 *
0-
02
b0 6
#942570000000
1!
1%
1-
12
#942580000000
0!
0%
b1 *
0-
02
b1 6
#942590000000
1!
1%
1-
12
#942600000000
0!
0%
b10 *
0-
02
b10 6
#942610000000
1!
1%
1-
12
#942620000000
0!
0%
b11 *
0-
02
b11 6
#942630000000
1!
1%
1-
12
15
#942640000000
0!
0%
b100 *
0-
02
b100 6
#942650000000
1!
1%
1-
12
#942660000000
0!
0%
b101 *
0-
02
b101 6
#942670000000
1!
1%
1-
12
#942680000000
0!
0%
b110 *
0-
02
b110 6
#942690000000
1!
1%
1-
12
#942700000000
0!
0%
b111 *
0-
02
b111 6
#942710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#942720000000
0!
0%
b0 *
0-
02
b0 6
#942730000000
1!
1%
1-
12
#942740000000
0!
0%
b1 *
0-
02
b1 6
#942750000000
1!
1%
1-
12
#942760000000
0!
0%
b10 *
0-
02
b10 6
#942770000000
1!
1%
1-
12
#942780000000
0!
0%
b11 *
0-
02
b11 6
#942790000000
1!
1%
1-
12
15
#942800000000
0!
0%
b100 *
0-
02
b100 6
#942810000000
1!
1%
1-
12
#942820000000
0!
0%
b101 *
0-
02
b101 6
#942830000000
1!
1%
1-
12
#942840000000
0!
0%
b110 *
0-
02
b110 6
#942850000000
1!
1%
1-
12
#942860000000
0!
0%
b111 *
0-
02
b111 6
#942870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#942880000000
0!
0%
b0 *
0-
02
b0 6
#942890000000
1!
1%
1-
12
#942900000000
0!
0%
b1 *
0-
02
b1 6
#942910000000
1!
1%
1-
12
#942920000000
0!
0%
b10 *
0-
02
b10 6
#942930000000
1!
1%
1-
12
#942940000000
0!
0%
b11 *
0-
02
b11 6
#942950000000
1!
1%
1-
12
15
#942960000000
0!
0%
b100 *
0-
02
b100 6
#942970000000
1!
1%
1-
12
#942980000000
0!
0%
b101 *
0-
02
b101 6
#942990000000
1!
1%
1-
12
#943000000000
0!
0%
b110 *
0-
02
b110 6
#943010000000
1!
1%
1-
12
#943020000000
0!
0%
b111 *
0-
02
b111 6
#943030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#943040000000
0!
0%
b0 *
0-
02
b0 6
#943050000000
1!
1%
1-
12
#943060000000
0!
0%
b1 *
0-
02
b1 6
#943070000000
1!
1%
1-
12
#943080000000
0!
0%
b10 *
0-
02
b10 6
#943090000000
1!
1%
1-
12
#943100000000
0!
0%
b11 *
0-
02
b11 6
#943110000000
1!
1%
1-
12
15
#943120000000
0!
0%
b100 *
0-
02
b100 6
#943130000000
1!
1%
1-
12
#943140000000
0!
0%
b101 *
0-
02
b101 6
#943150000000
1!
1%
1-
12
#943160000000
0!
0%
b110 *
0-
02
b110 6
#943170000000
1!
1%
1-
12
#943180000000
0!
0%
b111 *
0-
02
b111 6
#943190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#943200000000
0!
0%
b0 *
0-
02
b0 6
#943210000000
1!
1%
1-
12
#943220000000
0!
0%
b1 *
0-
02
b1 6
#943230000000
1!
1%
1-
12
#943240000000
0!
0%
b10 *
0-
02
b10 6
#943250000000
1!
1%
1-
12
#943260000000
0!
0%
b11 *
0-
02
b11 6
#943270000000
1!
1%
1-
12
15
#943280000000
0!
0%
b100 *
0-
02
b100 6
#943290000000
1!
1%
1-
12
#943300000000
0!
0%
b101 *
0-
02
b101 6
#943310000000
1!
1%
1-
12
#943320000000
0!
0%
b110 *
0-
02
b110 6
#943330000000
1!
1%
1-
12
#943340000000
0!
0%
b111 *
0-
02
b111 6
#943350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#943360000000
0!
0%
b0 *
0-
02
b0 6
#943370000000
1!
1%
1-
12
#943380000000
0!
0%
b1 *
0-
02
b1 6
#943390000000
1!
1%
1-
12
#943400000000
0!
0%
b10 *
0-
02
b10 6
#943410000000
1!
1%
1-
12
#943420000000
0!
0%
b11 *
0-
02
b11 6
#943430000000
1!
1%
1-
12
15
#943440000000
0!
0%
b100 *
0-
02
b100 6
#943450000000
1!
1%
1-
12
#943460000000
0!
0%
b101 *
0-
02
b101 6
#943470000000
1!
1%
1-
12
#943480000000
0!
0%
b110 *
0-
02
b110 6
#943490000000
1!
1%
1-
12
#943500000000
0!
0%
b111 *
0-
02
b111 6
#943510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#943520000000
0!
0%
b0 *
0-
02
b0 6
#943530000000
1!
1%
1-
12
#943540000000
0!
0%
b1 *
0-
02
b1 6
#943550000000
1!
1%
1-
12
#943560000000
0!
0%
b10 *
0-
02
b10 6
#943570000000
1!
1%
1-
12
#943580000000
0!
0%
b11 *
0-
02
b11 6
#943590000000
1!
1%
1-
12
15
#943600000000
0!
0%
b100 *
0-
02
b100 6
#943610000000
1!
1%
1-
12
#943620000000
0!
0%
b101 *
0-
02
b101 6
#943630000000
1!
1%
1-
12
#943640000000
0!
0%
b110 *
0-
02
b110 6
#943650000000
1!
1%
1-
12
#943660000000
0!
0%
b111 *
0-
02
b111 6
#943670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#943680000000
0!
0%
b0 *
0-
02
b0 6
#943690000000
1!
1%
1-
12
#943700000000
0!
0%
b1 *
0-
02
b1 6
#943710000000
1!
1%
1-
12
#943720000000
0!
0%
b10 *
0-
02
b10 6
#943730000000
1!
1%
1-
12
#943740000000
0!
0%
b11 *
0-
02
b11 6
#943750000000
1!
1%
1-
12
15
#943760000000
0!
0%
b100 *
0-
02
b100 6
#943770000000
1!
1%
1-
12
#943780000000
0!
0%
b101 *
0-
02
b101 6
#943790000000
1!
1%
1-
12
#943800000000
0!
0%
b110 *
0-
02
b110 6
#943810000000
1!
1%
1-
12
#943820000000
0!
0%
b111 *
0-
02
b111 6
#943830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#943840000000
0!
0%
b0 *
0-
02
b0 6
#943850000000
1!
1%
1-
12
#943860000000
0!
0%
b1 *
0-
02
b1 6
#943870000000
1!
1%
1-
12
#943880000000
0!
0%
b10 *
0-
02
b10 6
#943890000000
1!
1%
1-
12
#943900000000
0!
0%
b11 *
0-
02
b11 6
#943910000000
1!
1%
1-
12
15
#943920000000
0!
0%
b100 *
0-
02
b100 6
#943930000000
1!
1%
1-
12
#943940000000
0!
0%
b101 *
0-
02
b101 6
#943950000000
1!
1%
1-
12
#943960000000
0!
0%
b110 *
0-
02
b110 6
#943970000000
1!
1%
1-
12
#943980000000
0!
0%
b111 *
0-
02
b111 6
#943990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#944000000000
0!
0%
b0 *
0-
02
b0 6
#944010000000
1!
1%
1-
12
#944020000000
0!
0%
b1 *
0-
02
b1 6
#944030000000
1!
1%
1-
12
#944040000000
0!
0%
b10 *
0-
02
b10 6
#944050000000
1!
1%
1-
12
#944060000000
0!
0%
b11 *
0-
02
b11 6
#944070000000
1!
1%
1-
12
15
#944080000000
0!
0%
b100 *
0-
02
b100 6
#944090000000
1!
1%
1-
12
#944100000000
0!
0%
b101 *
0-
02
b101 6
#944110000000
1!
1%
1-
12
#944120000000
0!
0%
b110 *
0-
02
b110 6
#944130000000
1!
1%
1-
12
#944140000000
0!
0%
b111 *
0-
02
b111 6
#944150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#944160000000
0!
0%
b0 *
0-
02
b0 6
#944170000000
1!
1%
1-
12
#944180000000
0!
0%
b1 *
0-
02
b1 6
#944190000000
1!
1%
1-
12
#944200000000
0!
0%
b10 *
0-
02
b10 6
#944210000000
1!
1%
1-
12
#944220000000
0!
0%
b11 *
0-
02
b11 6
#944230000000
1!
1%
1-
12
15
#944240000000
0!
0%
b100 *
0-
02
b100 6
#944250000000
1!
1%
1-
12
#944260000000
0!
0%
b101 *
0-
02
b101 6
#944270000000
1!
1%
1-
12
#944280000000
0!
0%
b110 *
0-
02
b110 6
#944290000000
1!
1%
1-
12
#944300000000
0!
0%
b111 *
0-
02
b111 6
#944310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#944320000000
0!
0%
b0 *
0-
02
b0 6
#944330000000
1!
1%
1-
12
#944340000000
0!
0%
b1 *
0-
02
b1 6
#944350000000
1!
1%
1-
12
#944360000000
0!
0%
b10 *
0-
02
b10 6
#944370000000
1!
1%
1-
12
#944380000000
0!
0%
b11 *
0-
02
b11 6
#944390000000
1!
1%
1-
12
15
#944400000000
0!
0%
b100 *
0-
02
b100 6
#944410000000
1!
1%
1-
12
#944420000000
0!
0%
b101 *
0-
02
b101 6
#944430000000
1!
1%
1-
12
#944440000000
0!
0%
b110 *
0-
02
b110 6
#944450000000
1!
1%
1-
12
#944460000000
0!
0%
b111 *
0-
02
b111 6
#944470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#944480000000
0!
0%
b0 *
0-
02
b0 6
#944490000000
1!
1%
1-
12
#944500000000
0!
0%
b1 *
0-
02
b1 6
#944510000000
1!
1%
1-
12
#944520000000
0!
0%
b10 *
0-
02
b10 6
#944530000000
1!
1%
1-
12
#944540000000
0!
0%
b11 *
0-
02
b11 6
#944550000000
1!
1%
1-
12
15
#944560000000
0!
0%
b100 *
0-
02
b100 6
#944570000000
1!
1%
1-
12
#944580000000
0!
0%
b101 *
0-
02
b101 6
#944590000000
1!
1%
1-
12
#944600000000
0!
0%
b110 *
0-
02
b110 6
#944610000000
1!
1%
1-
12
#944620000000
0!
0%
b111 *
0-
02
b111 6
#944630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#944640000000
0!
0%
b0 *
0-
02
b0 6
#944650000000
1!
1%
1-
12
#944660000000
0!
0%
b1 *
0-
02
b1 6
#944670000000
1!
1%
1-
12
#944680000000
0!
0%
b10 *
0-
02
b10 6
#944690000000
1!
1%
1-
12
#944700000000
0!
0%
b11 *
0-
02
b11 6
#944710000000
1!
1%
1-
12
15
#944720000000
0!
0%
b100 *
0-
02
b100 6
#944730000000
1!
1%
1-
12
#944740000000
0!
0%
b101 *
0-
02
b101 6
#944750000000
1!
1%
1-
12
#944760000000
0!
0%
b110 *
0-
02
b110 6
#944770000000
1!
1%
1-
12
#944780000000
0!
0%
b111 *
0-
02
b111 6
#944790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#944800000000
0!
0%
b0 *
0-
02
b0 6
#944810000000
1!
1%
1-
12
#944820000000
0!
0%
b1 *
0-
02
b1 6
#944830000000
1!
1%
1-
12
#944840000000
0!
0%
b10 *
0-
02
b10 6
#944850000000
1!
1%
1-
12
#944860000000
0!
0%
b11 *
0-
02
b11 6
#944870000000
1!
1%
1-
12
15
#944880000000
0!
0%
b100 *
0-
02
b100 6
#944890000000
1!
1%
1-
12
#944900000000
0!
0%
b101 *
0-
02
b101 6
#944910000000
1!
1%
1-
12
#944920000000
0!
0%
b110 *
0-
02
b110 6
#944930000000
1!
1%
1-
12
#944940000000
0!
0%
b111 *
0-
02
b111 6
#944950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#944960000000
0!
0%
b0 *
0-
02
b0 6
#944970000000
1!
1%
1-
12
#944980000000
0!
0%
b1 *
0-
02
b1 6
#944990000000
1!
1%
1-
12
#945000000000
0!
0%
b10 *
0-
02
b10 6
#945010000000
1!
1%
1-
12
#945020000000
0!
0%
b11 *
0-
02
b11 6
#945030000000
1!
1%
1-
12
15
#945040000000
0!
0%
b100 *
0-
02
b100 6
#945050000000
1!
1%
1-
12
#945060000000
0!
0%
b101 *
0-
02
b101 6
#945070000000
1!
1%
1-
12
#945080000000
0!
0%
b110 *
0-
02
b110 6
#945090000000
1!
1%
1-
12
#945100000000
0!
0%
b111 *
0-
02
b111 6
#945110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#945120000000
0!
0%
b0 *
0-
02
b0 6
#945130000000
1!
1%
1-
12
#945140000000
0!
0%
b1 *
0-
02
b1 6
#945150000000
1!
1%
1-
12
#945160000000
0!
0%
b10 *
0-
02
b10 6
#945170000000
1!
1%
1-
12
#945180000000
0!
0%
b11 *
0-
02
b11 6
#945190000000
1!
1%
1-
12
15
#945200000000
0!
0%
b100 *
0-
02
b100 6
#945210000000
1!
1%
1-
12
#945220000000
0!
0%
b101 *
0-
02
b101 6
#945230000000
1!
1%
1-
12
#945240000000
0!
0%
b110 *
0-
02
b110 6
#945250000000
1!
1%
1-
12
#945260000000
0!
0%
b111 *
0-
02
b111 6
#945270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#945280000000
0!
0%
b0 *
0-
02
b0 6
#945290000000
1!
1%
1-
12
#945300000000
0!
0%
b1 *
0-
02
b1 6
#945310000000
1!
1%
1-
12
#945320000000
0!
0%
b10 *
0-
02
b10 6
#945330000000
1!
1%
1-
12
#945340000000
0!
0%
b11 *
0-
02
b11 6
#945350000000
1!
1%
1-
12
15
#945360000000
0!
0%
b100 *
0-
02
b100 6
#945370000000
1!
1%
1-
12
#945380000000
0!
0%
b101 *
0-
02
b101 6
#945390000000
1!
1%
1-
12
#945400000000
0!
0%
b110 *
0-
02
b110 6
#945410000000
1!
1%
1-
12
#945420000000
0!
0%
b111 *
0-
02
b111 6
#945430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#945440000000
0!
0%
b0 *
0-
02
b0 6
#945450000000
1!
1%
1-
12
#945460000000
0!
0%
b1 *
0-
02
b1 6
#945470000000
1!
1%
1-
12
#945480000000
0!
0%
b10 *
0-
02
b10 6
#945490000000
1!
1%
1-
12
#945500000000
0!
0%
b11 *
0-
02
b11 6
#945510000000
1!
1%
1-
12
15
#945520000000
0!
0%
b100 *
0-
02
b100 6
#945530000000
1!
1%
1-
12
#945540000000
0!
0%
b101 *
0-
02
b101 6
#945550000000
1!
1%
1-
12
#945560000000
0!
0%
b110 *
0-
02
b110 6
#945570000000
1!
1%
1-
12
#945580000000
0!
0%
b111 *
0-
02
b111 6
#945590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#945600000000
0!
0%
b0 *
0-
02
b0 6
#945610000000
1!
1%
1-
12
#945620000000
0!
0%
b1 *
0-
02
b1 6
#945630000000
1!
1%
1-
12
#945640000000
0!
0%
b10 *
0-
02
b10 6
#945650000000
1!
1%
1-
12
#945660000000
0!
0%
b11 *
0-
02
b11 6
#945670000000
1!
1%
1-
12
15
#945680000000
0!
0%
b100 *
0-
02
b100 6
#945690000000
1!
1%
1-
12
#945700000000
0!
0%
b101 *
0-
02
b101 6
#945710000000
1!
1%
1-
12
#945720000000
0!
0%
b110 *
0-
02
b110 6
#945730000000
1!
1%
1-
12
#945740000000
0!
0%
b111 *
0-
02
b111 6
#945750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#945760000000
0!
0%
b0 *
0-
02
b0 6
#945770000000
1!
1%
1-
12
#945780000000
0!
0%
b1 *
0-
02
b1 6
#945790000000
1!
1%
1-
12
#945800000000
0!
0%
b10 *
0-
02
b10 6
#945810000000
1!
1%
1-
12
#945820000000
0!
0%
b11 *
0-
02
b11 6
#945830000000
1!
1%
1-
12
15
#945840000000
0!
0%
b100 *
0-
02
b100 6
#945850000000
1!
1%
1-
12
#945860000000
0!
0%
b101 *
0-
02
b101 6
#945870000000
1!
1%
1-
12
#945880000000
0!
0%
b110 *
0-
02
b110 6
#945890000000
1!
1%
1-
12
#945900000000
0!
0%
b111 *
0-
02
b111 6
#945910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#945920000000
0!
0%
b0 *
0-
02
b0 6
#945930000000
1!
1%
1-
12
#945940000000
0!
0%
b1 *
0-
02
b1 6
#945950000000
1!
1%
1-
12
#945960000000
0!
0%
b10 *
0-
02
b10 6
#945970000000
1!
1%
1-
12
#945980000000
0!
0%
b11 *
0-
02
b11 6
#945990000000
1!
1%
1-
12
15
#946000000000
0!
0%
b100 *
0-
02
b100 6
#946010000000
1!
1%
1-
12
#946020000000
0!
0%
b101 *
0-
02
b101 6
#946030000000
1!
1%
1-
12
#946040000000
0!
0%
b110 *
0-
02
b110 6
#946050000000
1!
1%
1-
12
#946060000000
0!
0%
b111 *
0-
02
b111 6
#946070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#946080000000
0!
0%
b0 *
0-
02
b0 6
#946090000000
1!
1%
1-
12
#946100000000
0!
0%
b1 *
0-
02
b1 6
#946110000000
1!
1%
1-
12
#946120000000
0!
0%
b10 *
0-
02
b10 6
#946130000000
1!
1%
1-
12
#946140000000
0!
0%
b11 *
0-
02
b11 6
#946150000000
1!
1%
1-
12
15
#946160000000
0!
0%
b100 *
0-
02
b100 6
#946170000000
1!
1%
1-
12
#946180000000
0!
0%
b101 *
0-
02
b101 6
#946190000000
1!
1%
1-
12
#946200000000
0!
0%
b110 *
0-
02
b110 6
#946210000000
1!
1%
1-
12
#946220000000
0!
0%
b111 *
0-
02
b111 6
#946230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#946240000000
0!
0%
b0 *
0-
02
b0 6
#946250000000
1!
1%
1-
12
#946260000000
0!
0%
b1 *
0-
02
b1 6
#946270000000
1!
1%
1-
12
#946280000000
0!
0%
b10 *
0-
02
b10 6
#946290000000
1!
1%
1-
12
#946300000000
0!
0%
b11 *
0-
02
b11 6
#946310000000
1!
1%
1-
12
15
#946320000000
0!
0%
b100 *
0-
02
b100 6
#946330000000
1!
1%
1-
12
#946340000000
0!
0%
b101 *
0-
02
b101 6
#946350000000
1!
1%
1-
12
#946360000000
0!
0%
b110 *
0-
02
b110 6
#946370000000
1!
1%
1-
12
#946380000000
0!
0%
b111 *
0-
02
b111 6
#946390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#946400000000
0!
0%
b0 *
0-
02
b0 6
#946410000000
1!
1%
1-
12
#946420000000
0!
0%
b1 *
0-
02
b1 6
#946430000000
1!
1%
1-
12
#946440000000
0!
0%
b10 *
0-
02
b10 6
#946450000000
1!
1%
1-
12
#946460000000
0!
0%
b11 *
0-
02
b11 6
#946470000000
1!
1%
1-
12
15
#946480000000
0!
0%
b100 *
0-
02
b100 6
#946490000000
1!
1%
1-
12
#946500000000
0!
0%
b101 *
0-
02
b101 6
#946510000000
1!
1%
1-
12
#946520000000
0!
0%
b110 *
0-
02
b110 6
#946530000000
1!
1%
1-
12
#946540000000
0!
0%
b111 *
0-
02
b111 6
#946550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#946560000000
0!
0%
b0 *
0-
02
b0 6
#946570000000
1!
1%
1-
12
#946580000000
0!
0%
b1 *
0-
02
b1 6
#946590000000
1!
1%
1-
12
#946600000000
0!
0%
b10 *
0-
02
b10 6
#946610000000
1!
1%
1-
12
#946620000000
0!
0%
b11 *
0-
02
b11 6
#946630000000
1!
1%
1-
12
15
#946640000000
0!
0%
b100 *
0-
02
b100 6
#946650000000
1!
1%
1-
12
#946660000000
0!
0%
b101 *
0-
02
b101 6
#946670000000
1!
1%
1-
12
#946680000000
0!
0%
b110 *
0-
02
b110 6
#946690000000
1!
1%
1-
12
#946700000000
0!
0%
b111 *
0-
02
b111 6
#946710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#946720000000
0!
0%
b0 *
0-
02
b0 6
#946730000000
1!
1%
1-
12
#946740000000
0!
0%
b1 *
0-
02
b1 6
#946750000000
1!
1%
1-
12
#946760000000
0!
0%
b10 *
0-
02
b10 6
#946770000000
1!
1%
1-
12
#946780000000
0!
0%
b11 *
0-
02
b11 6
#946790000000
1!
1%
1-
12
15
#946800000000
0!
0%
b100 *
0-
02
b100 6
#946810000000
1!
1%
1-
12
#946820000000
0!
0%
b101 *
0-
02
b101 6
#946830000000
1!
1%
1-
12
#946840000000
0!
0%
b110 *
0-
02
b110 6
#946850000000
1!
1%
1-
12
#946860000000
0!
0%
b111 *
0-
02
b111 6
#946870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#946880000000
0!
0%
b0 *
0-
02
b0 6
#946890000000
1!
1%
1-
12
#946900000000
0!
0%
b1 *
0-
02
b1 6
#946910000000
1!
1%
1-
12
#946920000000
0!
0%
b10 *
0-
02
b10 6
#946930000000
1!
1%
1-
12
#946940000000
0!
0%
b11 *
0-
02
b11 6
#946950000000
1!
1%
1-
12
15
#946960000000
0!
0%
b100 *
0-
02
b100 6
#946970000000
1!
1%
1-
12
#946980000000
0!
0%
b101 *
0-
02
b101 6
#946990000000
1!
1%
1-
12
#947000000000
0!
0%
b110 *
0-
02
b110 6
#947010000000
1!
1%
1-
12
#947020000000
0!
0%
b111 *
0-
02
b111 6
#947030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#947040000000
0!
0%
b0 *
0-
02
b0 6
#947050000000
1!
1%
1-
12
#947060000000
0!
0%
b1 *
0-
02
b1 6
#947070000000
1!
1%
1-
12
#947080000000
0!
0%
b10 *
0-
02
b10 6
#947090000000
1!
1%
1-
12
#947100000000
0!
0%
b11 *
0-
02
b11 6
#947110000000
1!
1%
1-
12
15
#947120000000
0!
0%
b100 *
0-
02
b100 6
#947130000000
1!
1%
1-
12
#947140000000
0!
0%
b101 *
0-
02
b101 6
#947150000000
1!
1%
1-
12
#947160000000
0!
0%
b110 *
0-
02
b110 6
#947170000000
1!
1%
1-
12
#947180000000
0!
0%
b111 *
0-
02
b111 6
#947190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#947200000000
0!
0%
b0 *
0-
02
b0 6
#947210000000
1!
1%
1-
12
#947220000000
0!
0%
b1 *
0-
02
b1 6
#947230000000
1!
1%
1-
12
#947240000000
0!
0%
b10 *
0-
02
b10 6
#947250000000
1!
1%
1-
12
#947260000000
0!
0%
b11 *
0-
02
b11 6
#947270000000
1!
1%
1-
12
15
#947280000000
0!
0%
b100 *
0-
02
b100 6
#947290000000
1!
1%
1-
12
#947300000000
0!
0%
b101 *
0-
02
b101 6
#947310000000
1!
1%
1-
12
#947320000000
0!
0%
b110 *
0-
02
b110 6
#947330000000
1!
1%
1-
12
#947340000000
0!
0%
b111 *
0-
02
b111 6
#947350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#947360000000
0!
0%
b0 *
0-
02
b0 6
#947370000000
1!
1%
1-
12
#947380000000
0!
0%
b1 *
0-
02
b1 6
#947390000000
1!
1%
1-
12
#947400000000
0!
0%
b10 *
0-
02
b10 6
#947410000000
1!
1%
1-
12
#947420000000
0!
0%
b11 *
0-
02
b11 6
#947430000000
1!
1%
1-
12
15
#947440000000
0!
0%
b100 *
0-
02
b100 6
#947450000000
1!
1%
1-
12
#947460000000
0!
0%
b101 *
0-
02
b101 6
#947470000000
1!
1%
1-
12
#947480000000
0!
0%
b110 *
0-
02
b110 6
#947490000000
1!
1%
1-
12
#947500000000
0!
0%
b111 *
0-
02
b111 6
#947510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#947520000000
0!
0%
b0 *
0-
02
b0 6
#947530000000
1!
1%
1-
12
#947540000000
0!
0%
b1 *
0-
02
b1 6
#947550000000
1!
1%
1-
12
#947560000000
0!
0%
b10 *
0-
02
b10 6
#947570000000
1!
1%
1-
12
#947580000000
0!
0%
b11 *
0-
02
b11 6
#947590000000
1!
1%
1-
12
15
#947600000000
0!
0%
b100 *
0-
02
b100 6
#947610000000
1!
1%
1-
12
#947620000000
0!
0%
b101 *
0-
02
b101 6
#947630000000
1!
1%
1-
12
#947640000000
0!
0%
b110 *
0-
02
b110 6
#947650000000
1!
1%
1-
12
#947660000000
0!
0%
b111 *
0-
02
b111 6
#947670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#947680000000
0!
0%
b0 *
0-
02
b0 6
#947690000000
1!
1%
1-
12
#947700000000
0!
0%
b1 *
0-
02
b1 6
#947710000000
1!
1%
1-
12
#947720000000
0!
0%
b10 *
0-
02
b10 6
#947730000000
1!
1%
1-
12
#947740000000
0!
0%
b11 *
0-
02
b11 6
#947750000000
1!
1%
1-
12
15
#947760000000
0!
0%
b100 *
0-
02
b100 6
#947770000000
1!
1%
1-
12
#947780000000
0!
0%
b101 *
0-
02
b101 6
#947790000000
1!
1%
1-
12
#947800000000
0!
0%
b110 *
0-
02
b110 6
#947810000000
1!
1%
1-
12
#947820000000
0!
0%
b111 *
0-
02
b111 6
#947830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#947840000000
0!
0%
b0 *
0-
02
b0 6
#947850000000
1!
1%
1-
12
#947860000000
0!
0%
b1 *
0-
02
b1 6
#947870000000
1!
1%
1-
12
#947880000000
0!
0%
b10 *
0-
02
b10 6
#947890000000
1!
1%
1-
12
#947900000000
0!
0%
b11 *
0-
02
b11 6
#947910000000
1!
1%
1-
12
15
#947920000000
0!
0%
b100 *
0-
02
b100 6
#947930000000
1!
1%
1-
12
#947940000000
0!
0%
b101 *
0-
02
b101 6
#947950000000
1!
1%
1-
12
#947960000000
0!
0%
b110 *
0-
02
b110 6
#947970000000
1!
1%
1-
12
#947980000000
0!
0%
b111 *
0-
02
b111 6
#947990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#948000000000
0!
0%
b0 *
0-
02
b0 6
#948010000000
1!
1%
1-
12
#948020000000
0!
0%
b1 *
0-
02
b1 6
#948030000000
1!
1%
1-
12
#948040000000
0!
0%
b10 *
0-
02
b10 6
#948050000000
1!
1%
1-
12
#948060000000
0!
0%
b11 *
0-
02
b11 6
#948070000000
1!
1%
1-
12
15
#948080000000
0!
0%
b100 *
0-
02
b100 6
#948090000000
1!
1%
1-
12
#948100000000
0!
0%
b101 *
0-
02
b101 6
#948110000000
1!
1%
1-
12
#948120000000
0!
0%
b110 *
0-
02
b110 6
#948130000000
1!
1%
1-
12
#948140000000
0!
0%
b111 *
0-
02
b111 6
#948150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#948160000000
0!
0%
b0 *
0-
02
b0 6
#948170000000
1!
1%
1-
12
#948180000000
0!
0%
b1 *
0-
02
b1 6
#948190000000
1!
1%
1-
12
#948200000000
0!
0%
b10 *
0-
02
b10 6
#948210000000
1!
1%
1-
12
#948220000000
0!
0%
b11 *
0-
02
b11 6
#948230000000
1!
1%
1-
12
15
#948240000000
0!
0%
b100 *
0-
02
b100 6
#948250000000
1!
1%
1-
12
#948260000000
0!
0%
b101 *
0-
02
b101 6
#948270000000
1!
1%
1-
12
#948280000000
0!
0%
b110 *
0-
02
b110 6
#948290000000
1!
1%
1-
12
#948300000000
0!
0%
b111 *
0-
02
b111 6
#948310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#948320000000
0!
0%
b0 *
0-
02
b0 6
#948330000000
1!
1%
1-
12
#948340000000
0!
0%
b1 *
0-
02
b1 6
#948350000000
1!
1%
1-
12
#948360000000
0!
0%
b10 *
0-
02
b10 6
#948370000000
1!
1%
1-
12
#948380000000
0!
0%
b11 *
0-
02
b11 6
#948390000000
1!
1%
1-
12
15
#948400000000
0!
0%
b100 *
0-
02
b100 6
#948410000000
1!
1%
1-
12
#948420000000
0!
0%
b101 *
0-
02
b101 6
#948430000000
1!
1%
1-
12
#948440000000
0!
0%
b110 *
0-
02
b110 6
#948450000000
1!
1%
1-
12
#948460000000
0!
0%
b111 *
0-
02
b111 6
#948470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#948480000000
0!
0%
b0 *
0-
02
b0 6
#948490000000
1!
1%
1-
12
#948500000000
0!
0%
b1 *
0-
02
b1 6
#948510000000
1!
1%
1-
12
#948520000000
0!
0%
b10 *
0-
02
b10 6
#948530000000
1!
1%
1-
12
#948540000000
0!
0%
b11 *
0-
02
b11 6
#948550000000
1!
1%
1-
12
15
#948560000000
0!
0%
b100 *
0-
02
b100 6
#948570000000
1!
1%
1-
12
#948580000000
0!
0%
b101 *
0-
02
b101 6
#948590000000
1!
1%
1-
12
#948600000000
0!
0%
b110 *
0-
02
b110 6
#948610000000
1!
1%
1-
12
#948620000000
0!
0%
b111 *
0-
02
b111 6
#948630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#948640000000
0!
0%
b0 *
0-
02
b0 6
#948650000000
1!
1%
1-
12
#948660000000
0!
0%
b1 *
0-
02
b1 6
#948670000000
1!
1%
1-
12
#948680000000
0!
0%
b10 *
0-
02
b10 6
#948690000000
1!
1%
1-
12
#948700000000
0!
0%
b11 *
0-
02
b11 6
#948710000000
1!
1%
1-
12
15
#948720000000
0!
0%
b100 *
0-
02
b100 6
#948730000000
1!
1%
1-
12
#948740000000
0!
0%
b101 *
0-
02
b101 6
#948750000000
1!
1%
1-
12
#948760000000
0!
0%
b110 *
0-
02
b110 6
#948770000000
1!
1%
1-
12
#948780000000
0!
0%
b111 *
0-
02
b111 6
#948790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#948800000000
0!
0%
b0 *
0-
02
b0 6
#948810000000
1!
1%
1-
12
#948820000000
0!
0%
b1 *
0-
02
b1 6
#948830000000
1!
1%
1-
12
#948840000000
0!
0%
b10 *
0-
02
b10 6
#948850000000
1!
1%
1-
12
#948860000000
0!
0%
b11 *
0-
02
b11 6
#948870000000
1!
1%
1-
12
15
#948880000000
0!
0%
b100 *
0-
02
b100 6
#948890000000
1!
1%
1-
12
#948900000000
0!
0%
b101 *
0-
02
b101 6
#948910000000
1!
1%
1-
12
#948920000000
0!
0%
b110 *
0-
02
b110 6
#948930000000
1!
1%
1-
12
#948940000000
0!
0%
b111 *
0-
02
b111 6
#948950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#948960000000
0!
0%
b0 *
0-
02
b0 6
#948970000000
1!
1%
1-
12
#948980000000
0!
0%
b1 *
0-
02
b1 6
#948990000000
1!
1%
1-
12
#949000000000
0!
0%
b10 *
0-
02
b10 6
#949010000000
1!
1%
1-
12
#949020000000
0!
0%
b11 *
0-
02
b11 6
#949030000000
1!
1%
1-
12
15
#949040000000
0!
0%
b100 *
0-
02
b100 6
#949050000000
1!
1%
1-
12
#949060000000
0!
0%
b101 *
0-
02
b101 6
#949070000000
1!
1%
1-
12
#949080000000
0!
0%
b110 *
0-
02
b110 6
#949090000000
1!
1%
1-
12
#949100000000
0!
0%
b111 *
0-
02
b111 6
#949110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#949120000000
0!
0%
b0 *
0-
02
b0 6
#949130000000
1!
1%
1-
12
#949140000000
0!
0%
b1 *
0-
02
b1 6
#949150000000
1!
1%
1-
12
#949160000000
0!
0%
b10 *
0-
02
b10 6
#949170000000
1!
1%
1-
12
#949180000000
0!
0%
b11 *
0-
02
b11 6
#949190000000
1!
1%
1-
12
15
#949200000000
0!
0%
b100 *
0-
02
b100 6
#949210000000
1!
1%
1-
12
#949220000000
0!
0%
b101 *
0-
02
b101 6
#949230000000
1!
1%
1-
12
#949240000000
0!
0%
b110 *
0-
02
b110 6
#949250000000
1!
1%
1-
12
#949260000000
0!
0%
b111 *
0-
02
b111 6
#949270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#949280000000
0!
0%
b0 *
0-
02
b0 6
#949290000000
1!
1%
1-
12
#949300000000
0!
0%
b1 *
0-
02
b1 6
#949310000000
1!
1%
1-
12
#949320000000
0!
0%
b10 *
0-
02
b10 6
#949330000000
1!
1%
1-
12
#949340000000
0!
0%
b11 *
0-
02
b11 6
#949350000000
1!
1%
1-
12
15
#949360000000
0!
0%
b100 *
0-
02
b100 6
#949370000000
1!
1%
1-
12
#949380000000
0!
0%
b101 *
0-
02
b101 6
#949390000000
1!
1%
1-
12
#949400000000
0!
0%
b110 *
0-
02
b110 6
#949410000000
1!
1%
1-
12
#949420000000
0!
0%
b111 *
0-
02
b111 6
#949430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#949440000000
0!
0%
b0 *
0-
02
b0 6
#949450000000
1!
1%
1-
12
#949460000000
0!
0%
b1 *
0-
02
b1 6
#949470000000
1!
1%
1-
12
#949480000000
0!
0%
b10 *
0-
02
b10 6
#949490000000
1!
1%
1-
12
#949500000000
0!
0%
b11 *
0-
02
b11 6
#949510000000
1!
1%
1-
12
15
#949520000000
0!
0%
b100 *
0-
02
b100 6
#949530000000
1!
1%
1-
12
#949540000000
0!
0%
b101 *
0-
02
b101 6
#949550000000
1!
1%
1-
12
#949560000000
0!
0%
b110 *
0-
02
b110 6
#949570000000
1!
1%
1-
12
#949580000000
0!
0%
b111 *
0-
02
b111 6
#949590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#949600000000
0!
0%
b0 *
0-
02
b0 6
#949610000000
1!
1%
1-
12
#949620000000
0!
0%
b1 *
0-
02
b1 6
#949630000000
1!
1%
1-
12
#949640000000
0!
0%
b10 *
0-
02
b10 6
#949650000000
1!
1%
1-
12
#949660000000
0!
0%
b11 *
0-
02
b11 6
#949670000000
1!
1%
1-
12
15
#949680000000
0!
0%
b100 *
0-
02
b100 6
#949690000000
1!
1%
1-
12
#949700000000
0!
0%
b101 *
0-
02
b101 6
#949710000000
1!
1%
1-
12
#949720000000
0!
0%
b110 *
0-
02
b110 6
#949730000000
1!
1%
1-
12
#949740000000
0!
0%
b111 *
0-
02
b111 6
#949750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#949760000000
0!
0%
b0 *
0-
02
b0 6
#949770000000
1!
1%
1-
12
#949780000000
0!
0%
b1 *
0-
02
b1 6
#949790000000
1!
1%
1-
12
#949800000000
0!
0%
b10 *
0-
02
b10 6
#949810000000
1!
1%
1-
12
#949820000000
0!
0%
b11 *
0-
02
b11 6
#949830000000
1!
1%
1-
12
15
#949840000000
0!
0%
b100 *
0-
02
b100 6
#949850000000
1!
1%
1-
12
#949860000000
0!
0%
b101 *
0-
02
b101 6
#949870000000
1!
1%
1-
12
#949880000000
0!
0%
b110 *
0-
02
b110 6
#949890000000
1!
1%
1-
12
#949900000000
0!
0%
b111 *
0-
02
b111 6
#949910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#949920000000
0!
0%
b0 *
0-
02
b0 6
#949930000000
1!
1%
1-
12
#949940000000
0!
0%
b1 *
0-
02
b1 6
#949950000000
1!
1%
1-
12
#949960000000
0!
0%
b10 *
0-
02
b10 6
#949970000000
1!
1%
1-
12
#949980000000
0!
0%
b11 *
0-
02
b11 6
#949990000000
1!
1%
1-
12
15
#950000000000
0!
0%
b100 *
0-
02
b100 6
#950010000000
1!
1%
1-
12
#950020000000
0!
0%
b101 *
0-
02
b101 6
#950030000000
1!
1%
1-
12
#950040000000
0!
0%
b110 *
0-
02
b110 6
#950050000000
1!
1%
1-
12
#950060000000
0!
0%
b111 *
0-
02
b111 6
#950070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#950080000000
0!
0%
b0 *
0-
02
b0 6
#950090000000
1!
1%
1-
12
#950100000000
0!
0%
b1 *
0-
02
b1 6
#950110000000
1!
1%
1-
12
#950120000000
0!
0%
b10 *
0-
02
b10 6
#950130000000
1!
1%
1-
12
#950140000000
0!
0%
b11 *
0-
02
b11 6
#950150000000
1!
1%
1-
12
15
#950160000000
0!
0%
b100 *
0-
02
b100 6
#950170000000
1!
1%
1-
12
#950180000000
0!
0%
b101 *
0-
02
b101 6
#950190000000
1!
1%
1-
12
#950200000000
0!
0%
b110 *
0-
02
b110 6
#950210000000
1!
1%
1-
12
#950220000000
0!
0%
b111 *
0-
02
b111 6
#950230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#950240000000
0!
0%
b0 *
0-
02
b0 6
#950250000000
1!
1%
1-
12
#950260000000
0!
0%
b1 *
0-
02
b1 6
#950270000000
1!
1%
1-
12
#950280000000
0!
0%
b10 *
0-
02
b10 6
#950290000000
1!
1%
1-
12
#950300000000
0!
0%
b11 *
0-
02
b11 6
#950310000000
1!
1%
1-
12
15
#950320000000
0!
0%
b100 *
0-
02
b100 6
#950330000000
1!
1%
1-
12
#950340000000
0!
0%
b101 *
0-
02
b101 6
#950350000000
1!
1%
1-
12
#950360000000
0!
0%
b110 *
0-
02
b110 6
#950370000000
1!
1%
1-
12
#950380000000
0!
0%
b111 *
0-
02
b111 6
#950390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#950400000000
0!
0%
b0 *
0-
02
b0 6
#950410000000
1!
1%
1-
12
#950420000000
0!
0%
b1 *
0-
02
b1 6
#950430000000
1!
1%
1-
12
#950440000000
0!
0%
b10 *
0-
02
b10 6
#950450000000
1!
1%
1-
12
#950460000000
0!
0%
b11 *
0-
02
b11 6
#950470000000
1!
1%
1-
12
15
#950480000000
0!
0%
b100 *
0-
02
b100 6
#950490000000
1!
1%
1-
12
#950500000000
0!
0%
b101 *
0-
02
b101 6
#950510000000
1!
1%
1-
12
#950520000000
0!
0%
b110 *
0-
02
b110 6
#950530000000
1!
1%
1-
12
#950540000000
0!
0%
b111 *
0-
02
b111 6
#950550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#950560000000
0!
0%
b0 *
0-
02
b0 6
#950570000000
1!
1%
1-
12
#950580000000
0!
0%
b1 *
0-
02
b1 6
#950590000000
1!
1%
1-
12
#950600000000
0!
0%
b10 *
0-
02
b10 6
#950610000000
1!
1%
1-
12
#950620000000
0!
0%
b11 *
0-
02
b11 6
#950630000000
1!
1%
1-
12
15
#950640000000
0!
0%
b100 *
0-
02
b100 6
#950650000000
1!
1%
1-
12
#950660000000
0!
0%
b101 *
0-
02
b101 6
#950670000000
1!
1%
1-
12
#950680000000
0!
0%
b110 *
0-
02
b110 6
#950690000000
1!
1%
1-
12
#950700000000
0!
0%
b111 *
0-
02
b111 6
#950710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#950720000000
0!
0%
b0 *
0-
02
b0 6
#950730000000
1!
1%
1-
12
#950740000000
0!
0%
b1 *
0-
02
b1 6
#950750000000
1!
1%
1-
12
#950760000000
0!
0%
b10 *
0-
02
b10 6
#950770000000
1!
1%
1-
12
#950780000000
0!
0%
b11 *
0-
02
b11 6
#950790000000
1!
1%
1-
12
15
#950800000000
0!
0%
b100 *
0-
02
b100 6
#950810000000
1!
1%
1-
12
#950820000000
0!
0%
b101 *
0-
02
b101 6
#950830000000
1!
1%
1-
12
#950840000000
0!
0%
b110 *
0-
02
b110 6
#950850000000
1!
1%
1-
12
#950860000000
0!
0%
b111 *
0-
02
b111 6
#950870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#950880000000
0!
0%
b0 *
0-
02
b0 6
#950890000000
1!
1%
1-
12
#950900000000
0!
0%
b1 *
0-
02
b1 6
#950910000000
1!
1%
1-
12
#950920000000
0!
0%
b10 *
0-
02
b10 6
#950930000000
1!
1%
1-
12
#950940000000
0!
0%
b11 *
0-
02
b11 6
#950950000000
1!
1%
1-
12
15
#950960000000
0!
0%
b100 *
0-
02
b100 6
#950970000000
1!
1%
1-
12
#950980000000
0!
0%
b101 *
0-
02
b101 6
#950990000000
1!
1%
1-
12
#951000000000
0!
0%
b110 *
0-
02
b110 6
#951010000000
1!
1%
1-
12
#951020000000
0!
0%
b111 *
0-
02
b111 6
#951030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#951040000000
0!
0%
b0 *
0-
02
b0 6
#951050000000
1!
1%
1-
12
#951060000000
0!
0%
b1 *
0-
02
b1 6
#951070000000
1!
1%
1-
12
#951080000000
0!
0%
b10 *
0-
02
b10 6
#951090000000
1!
1%
1-
12
#951100000000
0!
0%
b11 *
0-
02
b11 6
#951110000000
1!
1%
1-
12
15
#951120000000
0!
0%
b100 *
0-
02
b100 6
#951130000000
1!
1%
1-
12
#951140000000
0!
0%
b101 *
0-
02
b101 6
#951150000000
1!
1%
1-
12
#951160000000
0!
0%
b110 *
0-
02
b110 6
#951170000000
1!
1%
1-
12
#951180000000
0!
0%
b111 *
0-
02
b111 6
#951190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#951200000000
0!
0%
b0 *
0-
02
b0 6
#951210000000
1!
1%
1-
12
#951220000000
0!
0%
b1 *
0-
02
b1 6
#951230000000
1!
1%
1-
12
#951240000000
0!
0%
b10 *
0-
02
b10 6
#951250000000
1!
1%
1-
12
#951260000000
0!
0%
b11 *
0-
02
b11 6
#951270000000
1!
1%
1-
12
15
#951280000000
0!
0%
b100 *
0-
02
b100 6
#951290000000
1!
1%
1-
12
#951300000000
0!
0%
b101 *
0-
02
b101 6
#951310000000
1!
1%
1-
12
#951320000000
0!
0%
b110 *
0-
02
b110 6
#951330000000
1!
1%
1-
12
#951340000000
0!
0%
b111 *
0-
02
b111 6
#951350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#951360000000
0!
0%
b0 *
0-
02
b0 6
#951370000000
1!
1%
1-
12
#951380000000
0!
0%
b1 *
0-
02
b1 6
#951390000000
1!
1%
1-
12
#951400000000
0!
0%
b10 *
0-
02
b10 6
#951410000000
1!
1%
1-
12
#951420000000
0!
0%
b11 *
0-
02
b11 6
#951430000000
1!
1%
1-
12
15
#951440000000
0!
0%
b100 *
0-
02
b100 6
#951450000000
1!
1%
1-
12
#951460000000
0!
0%
b101 *
0-
02
b101 6
#951470000000
1!
1%
1-
12
#951480000000
0!
0%
b110 *
0-
02
b110 6
#951490000000
1!
1%
1-
12
#951500000000
0!
0%
b111 *
0-
02
b111 6
#951510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#951520000000
0!
0%
b0 *
0-
02
b0 6
#951530000000
1!
1%
1-
12
#951540000000
0!
0%
b1 *
0-
02
b1 6
#951550000000
1!
1%
1-
12
#951560000000
0!
0%
b10 *
0-
02
b10 6
#951570000000
1!
1%
1-
12
#951580000000
0!
0%
b11 *
0-
02
b11 6
#951590000000
1!
1%
1-
12
15
#951600000000
0!
0%
b100 *
0-
02
b100 6
#951610000000
1!
1%
1-
12
#951620000000
0!
0%
b101 *
0-
02
b101 6
#951630000000
1!
1%
1-
12
#951640000000
0!
0%
b110 *
0-
02
b110 6
#951650000000
1!
1%
1-
12
#951660000000
0!
0%
b111 *
0-
02
b111 6
#951670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#951680000000
0!
0%
b0 *
0-
02
b0 6
#951690000000
1!
1%
1-
12
#951700000000
0!
0%
b1 *
0-
02
b1 6
#951710000000
1!
1%
1-
12
#951720000000
0!
0%
b10 *
0-
02
b10 6
#951730000000
1!
1%
1-
12
#951740000000
0!
0%
b11 *
0-
02
b11 6
#951750000000
1!
1%
1-
12
15
#951760000000
0!
0%
b100 *
0-
02
b100 6
#951770000000
1!
1%
1-
12
#951780000000
0!
0%
b101 *
0-
02
b101 6
#951790000000
1!
1%
1-
12
#951800000000
0!
0%
b110 *
0-
02
b110 6
#951810000000
1!
1%
1-
12
#951820000000
0!
0%
b111 *
0-
02
b111 6
#951830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#951840000000
0!
0%
b0 *
0-
02
b0 6
#951850000000
1!
1%
1-
12
#951860000000
0!
0%
b1 *
0-
02
b1 6
#951870000000
1!
1%
1-
12
#951880000000
0!
0%
b10 *
0-
02
b10 6
#951890000000
1!
1%
1-
12
#951900000000
0!
0%
b11 *
0-
02
b11 6
#951910000000
1!
1%
1-
12
15
#951920000000
0!
0%
b100 *
0-
02
b100 6
#951930000000
1!
1%
1-
12
#951940000000
0!
0%
b101 *
0-
02
b101 6
#951950000000
1!
1%
1-
12
#951960000000
0!
0%
b110 *
0-
02
b110 6
#951970000000
1!
1%
1-
12
#951980000000
0!
0%
b111 *
0-
02
b111 6
#951990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#952000000000
0!
0%
b0 *
0-
02
b0 6
#952010000000
1!
1%
1-
12
#952020000000
0!
0%
b1 *
0-
02
b1 6
#952030000000
1!
1%
1-
12
#952040000000
0!
0%
b10 *
0-
02
b10 6
#952050000000
1!
1%
1-
12
#952060000000
0!
0%
b11 *
0-
02
b11 6
#952070000000
1!
1%
1-
12
15
#952080000000
0!
0%
b100 *
0-
02
b100 6
#952090000000
1!
1%
1-
12
#952100000000
0!
0%
b101 *
0-
02
b101 6
#952110000000
1!
1%
1-
12
#952120000000
0!
0%
b110 *
0-
02
b110 6
#952130000000
1!
1%
1-
12
#952140000000
0!
0%
b111 *
0-
02
b111 6
#952150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#952160000000
0!
0%
b0 *
0-
02
b0 6
#952170000000
1!
1%
1-
12
#952180000000
0!
0%
b1 *
0-
02
b1 6
#952190000000
1!
1%
1-
12
#952200000000
0!
0%
b10 *
0-
02
b10 6
#952210000000
1!
1%
1-
12
#952220000000
0!
0%
b11 *
0-
02
b11 6
#952230000000
1!
1%
1-
12
15
#952240000000
0!
0%
b100 *
0-
02
b100 6
#952250000000
1!
1%
1-
12
#952260000000
0!
0%
b101 *
0-
02
b101 6
#952270000000
1!
1%
1-
12
#952280000000
0!
0%
b110 *
0-
02
b110 6
#952290000000
1!
1%
1-
12
#952300000000
0!
0%
b111 *
0-
02
b111 6
#952310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#952320000000
0!
0%
b0 *
0-
02
b0 6
#952330000000
1!
1%
1-
12
#952340000000
0!
0%
b1 *
0-
02
b1 6
#952350000000
1!
1%
1-
12
#952360000000
0!
0%
b10 *
0-
02
b10 6
#952370000000
1!
1%
1-
12
#952380000000
0!
0%
b11 *
0-
02
b11 6
#952390000000
1!
1%
1-
12
15
#952400000000
0!
0%
b100 *
0-
02
b100 6
#952410000000
1!
1%
1-
12
#952420000000
0!
0%
b101 *
0-
02
b101 6
#952430000000
1!
1%
1-
12
#952440000000
0!
0%
b110 *
0-
02
b110 6
#952450000000
1!
1%
1-
12
#952460000000
0!
0%
b111 *
0-
02
b111 6
#952470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#952480000000
0!
0%
b0 *
0-
02
b0 6
#952490000000
1!
1%
1-
12
#952500000000
0!
0%
b1 *
0-
02
b1 6
#952510000000
1!
1%
1-
12
#952520000000
0!
0%
b10 *
0-
02
b10 6
#952530000000
1!
1%
1-
12
#952540000000
0!
0%
b11 *
0-
02
b11 6
#952550000000
1!
1%
1-
12
15
#952560000000
0!
0%
b100 *
0-
02
b100 6
#952570000000
1!
1%
1-
12
#952580000000
0!
0%
b101 *
0-
02
b101 6
#952590000000
1!
1%
1-
12
#952600000000
0!
0%
b110 *
0-
02
b110 6
#952610000000
1!
1%
1-
12
#952620000000
0!
0%
b111 *
0-
02
b111 6
#952630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#952640000000
0!
0%
b0 *
0-
02
b0 6
#952650000000
1!
1%
1-
12
#952660000000
0!
0%
b1 *
0-
02
b1 6
#952670000000
1!
1%
1-
12
#952680000000
0!
0%
b10 *
0-
02
b10 6
#952690000000
1!
1%
1-
12
#952700000000
0!
0%
b11 *
0-
02
b11 6
#952710000000
1!
1%
1-
12
15
#952720000000
0!
0%
b100 *
0-
02
b100 6
#952730000000
1!
1%
1-
12
#952740000000
0!
0%
b101 *
0-
02
b101 6
#952750000000
1!
1%
1-
12
#952760000000
0!
0%
b110 *
0-
02
b110 6
#952770000000
1!
1%
1-
12
#952780000000
0!
0%
b111 *
0-
02
b111 6
#952790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#952800000000
0!
0%
b0 *
0-
02
b0 6
#952810000000
1!
1%
1-
12
#952820000000
0!
0%
b1 *
0-
02
b1 6
#952830000000
1!
1%
1-
12
#952840000000
0!
0%
b10 *
0-
02
b10 6
#952850000000
1!
1%
1-
12
#952860000000
0!
0%
b11 *
0-
02
b11 6
#952870000000
1!
1%
1-
12
15
#952880000000
0!
0%
b100 *
0-
02
b100 6
#952890000000
1!
1%
1-
12
#952900000000
0!
0%
b101 *
0-
02
b101 6
#952910000000
1!
1%
1-
12
#952920000000
0!
0%
b110 *
0-
02
b110 6
#952930000000
1!
1%
1-
12
#952940000000
0!
0%
b111 *
0-
02
b111 6
#952950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#952960000000
0!
0%
b0 *
0-
02
b0 6
#952970000000
1!
1%
1-
12
#952980000000
0!
0%
b1 *
0-
02
b1 6
#952990000000
1!
1%
1-
12
#953000000000
0!
0%
b10 *
0-
02
b10 6
#953010000000
1!
1%
1-
12
#953020000000
0!
0%
b11 *
0-
02
b11 6
#953030000000
1!
1%
1-
12
15
#953040000000
0!
0%
b100 *
0-
02
b100 6
#953050000000
1!
1%
1-
12
#953060000000
0!
0%
b101 *
0-
02
b101 6
#953070000000
1!
1%
1-
12
#953080000000
0!
0%
b110 *
0-
02
b110 6
#953090000000
1!
1%
1-
12
#953100000000
0!
0%
b111 *
0-
02
b111 6
#953110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#953120000000
0!
0%
b0 *
0-
02
b0 6
#953130000000
1!
1%
1-
12
#953140000000
0!
0%
b1 *
0-
02
b1 6
#953150000000
1!
1%
1-
12
#953160000000
0!
0%
b10 *
0-
02
b10 6
#953170000000
1!
1%
1-
12
#953180000000
0!
0%
b11 *
0-
02
b11 6
#953190000000
1!
1%
1-
12
15
#953200000000
0!
0%
b100 *
0-
02
b100 6
#953210000000
1!
1%
1-
12
#953220000000
0!
0%
b101 *
0-
02
b101 6
#953230000000
1!
1%
1-
12
#953240000000
0!
0%
b110 *
0-
02
b110 6
#953250000000
1!
1%
1-
12
#953260000000
0!
0%
b111 *
0-
02
b111 6
#953270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#953280000000
0!
0%
b0 *
0-
02
b0 6
#953290000000
1!
1%
1-
12
#953300000000
0!
0%
b1 *
0-
02
b1 6
#953310000000
1!
1%
1-
12
#953320000000
0!
0%
b10 *
0-
02
b10 6
#953330000000
1!
1%
1-
12
#953340000000
0!
0%
b11 *
0-
02
b11 6
#953350000000
1!
1%
1-
12
15
#953360000000
0!
0%
b100 *
0-
02
b100 6
#953370000000
1!
1%
1-
12
#953380000000
0!
0%
b101 *
0-
02
b101 6
#953390000000
1!
1%
1-
12
#953400000000
0!
0%
b110 *
0-
02
b110 6
#953410000000
1!
1%
1-
12
#953420000000
0!
0%
b111 *
0-
02
b111 6
#953430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#953440000000
0!
0%
b0 *
0-
02
b0 6
#953450000000
1!
1%
1-
12
#953460000000
0!
0%
b1 *
0-
02
b1 6
#953470000000
1!
1%
1-
12
#953480000000
0!
0%
b10 *
0-
02
b10 6
#953490000000
1!
1%
1-
12
#953500000000
0!
0%
b11 *
0-
02
b11 6
#953510000000
1!
1%
1-
12
15
#953520000000
0!
0%
b100 *
0-
02
b100 6
#953530000000
1!
1%
1-
12
#953540000000
0!
0%
b101 *
0-
02
b101 6
#953550000000
1!
1%
1-
12
#953560000000
0!
0%
b110 *
0-
02
b110 6
#953570000000
1!
1%
1-
12
#953580000000
0!
0%
b111 *
0-
02
b111 6
#953590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#953600000000
0!
0%
b0 *
0-
02
b0 6
#953610000000
1!
1%
1-
12
#953620000000
0!
0%
b1 *
0-
02
b1 6
#953630000000
1!
1%
1-
12
#953640000000
0!
0%
b10 *
0-
02
b10 6
#953650000000
1!
1%
1-
12
#953660000000
0!
0%
b11 *
0-
02
b11 6
#953670000000
1!
1%
1-
12
15
#953680000000
0!
0%
b100 *
0-
02
b100 6
#953690000000
1!
1%
1-
12
#953700000000
0!
0%
b101 *
0-
02
b101 6
#953710000000
1!
1%
1-
12
#953720000000
0!
0%
b110 *
0-
02
b110 6
#953730000000
1!
1%
1-
12
#953740000000
0!
0%
b111 *
0-
02
b111 6
#953750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#953760000000
0!
0%
b0 *
0-
02
b0 6
#953770000000
1!
1%
1-
12
#953780000000
0!
0%
b1 *
0-
02
b1 6
#953790000000
1!
1%
1-
12
#953800000000
0!
0%
b10 *
0-
02
b10 6
#953810000000
1!
1%
1-
12
#953820000000
0!
0%
b11 *
0-
02
b11 6
#953830000000
1!
1%
1-
12
15
#953840000000
0!
0%
b100 *
0-
02
b100 6
#953850000000
1!
1%
1-
12
#953860000000
0!
0%
b101 *
0-
02
b101 6
#953870000000
1!
1%
1-
12
#953880000000
0!
0%
b110 *
0-
02
b110 6
#953890000000
1!
1%
1-
12
#953900000000
0!
0%
b111 *
0-
02
b111 6
#953910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#953920000000
0!
0%
b0 *
0-
02
b0 6
#953930000000
1!
1%
1-
12
#953940000000
0!
0%
b1 *
0-
02
b1 6
#953950000000
1!
1%
1-
12
#953960000000
0!
0%
b10 *
0-
02
b10 6
#953970000000
1!
1%
1-
12
#953980000000
0!
0%
b11 *
0-
02
b11 6
#953990000000
1!
1%
1-
12
15
#954000000000
0!
0%
b100 *
0-
02
b100 6
#954010000000
1!
1%
1-
12
#954020000000
0!
0%
b101 *
0-
02
b101 6
#954030000000
1!
1%
1-
12
#954040000000
0!
0%
b110 *
0-
02
b110 6
#954050000000
1!
1%
1-
12
#954060000000
0!
0%
b111 *
0-
02
b111 6
#954070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#954080000000
0!
0%
b0 *
0-
02
b0 6
#954090000000
1!
1%
1-
12
#954100000000
0!
0%
b1 *
0-
02
b1 6
#954110000000
1!
1%
1-
12
#954120000000
0!
0%
b10 *
0-
02
b10 6
#954130000000
1!
1%
1-
12
#954140000000
0!
0%
b11 *
0-
02
b11 6
#954150000000
1!
1%
1-
12
15
#954160000000
0!
0%
b100 *
0-
02
b100 6
#954170000000
1!
1%
1-
12
#954180000000
0!
0%
b101 *
0-
02
b101 6
#954190000000
1!
1%
1-
12
#954200000000
0!
0%
b110 *
0-
02
b110 6
#954210000000
1!
1%
1-
12
#954220000000
0!
0%
b111 *
0-
02
b111 6
#954230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#954240000000
0!
0%
b0 *
0-
02
b0 6
#954250000000
1!
1%
1-
12
#954260000000
0!
0%
b1 *
0-
02
b1 6
#954270000000
1!
1%
1-
12
#954280000000
0!
0%
b10 *
0-
02
b10 6
#954290000000
1!
1%
1-
12
#954300000000
0!
0%
b11 *
0-
02
b11 6
#954310000000
1!
1%
1-
12
15
#954320000000
0!
0%
b100 *
0-
02
b100 6
#954330000000
1!
1%
1-
12
#954340000000
0!
0%
b101 *
0-
02
b101 6
#954350000000
1!
1%
1-
12
#954360000000
0!
0%
b110 *
0-
02
b110 6
#954370000000
1!
1%
1-
12
#954380000000
0!
0%
b111 *
0-
02
b111 6
#954390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#954400000000
0!
0%
b0 *
0-
02
b0 6
#954410000000
1!
1%
1-
12
#954420000000
0!
0%
b1 *
0-
02
b1 6
#954430000000
1!
1%
1-
12
#954440000000
0!
0%
b10 *
0-
02
b10 6
#954450000000
1!
1%
1-
12
#954460000000
0!
0%
b11 *
0-
02
b11 6
#954470000000
1!
1%
1-
12
15
#954480000000
0!
0%
b100 *
0-
02
b100 6
#954490000000
1!
1%
1-
12
#954500000000
0!
0%
b101 *
0-
02
b101 6
#954510000000
1!
1%
1-
12
#954520000000
0!
0%
b110 *
0-
02
b110 6
#954530000000
1!
1%
1-
12
#954540000000
0!
0%
b111 *
0-
02
b111 6
#954550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#954560000000
0!
0%
b0 *
0-
02
b0 6
#954570000000
1!
1%
1-
12
#954580000000
0!
0%
b1 *
0-
02
b1 6
#954590000000
1!
1%
1-
12
#954600000000
0!
0%
b10 *
0-
02
b10 6
#954610000000
1!
1%
1-
12
#954620000000
0!
0%
b11 *
0-
02
b11 6
#954630000000
1!
1%
1-
12
15
#954640000000
0!
0%
b100 *
0-
02
b100 6
#954650000000
1!
1%
1-
12
#954660000000
0!
0%
b101 *
0-
02
b101 6
#954670000000
1!
1%
1-
12
#954680000000
0!
0%
b110 *
0-
02
b110 6
#954690000000
1!
1%
1-
12
#954700000000
0!
0%
b111 *
0-
02
b111 6
#954710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#954720000000
0!
0%
b0 *
0-
02
b0 6
#954730000000
1!
1%
1-
12
#954740000000
0!
0%
b1 *
0-
02
b1 6
#954750000000
1!
1%
1-
12
#954760000000
0!
0%
b10 *
0-
02
b10 6
#954770000000
1!
1%
1-
12
#954780000000
0!
0%
b11 *
0-
02
b11 6
#954790000000
1!
1%
1-
12
15
#954800000000
0!
0%
b100 *
0-
02
b100 6
#954810000000
1!
1%
1-
12
#954820000000
0!
0%
b101 *
0-
02
b101 6
#954830000000
1!
1%
1-
12
#954840000000
0!
0%
b110 *
0-
02
b110 6
#954850000000
1!
1%
1-
12
#954860000000
0!
0%
b111 *
0-
02
b111 6
#954870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#954880000000
0!
0%
b0 *
0-
02
b0 6
#954890000000
1!
1%
1-
12
#954900000000
0!
0%
b1 *
0-
02
b1 6
#954910000000
1!
1%
1-
12
#954920000000
0!
0%
b10 *
0-
02
b10 6
#954930000000
1!
1%
1-
12
#954940000000
0!
0%
b11 *
0-
02
b11 6
#954950000000
1!
1%
1-
12
15
#954960000000
0!
0%
b100 *
0-
02
b100 6
#954970000000
1!
1%
1-
12
#954980000000
0!
0%
b101 *
0-
02
b101 6
#954990000000
1!
1%
1-
12
#955000000000
0!
0%
b110 *
0-
02
b110 6
#955010000000
1!
1%
1-
12
#955020000000
0!
0%
b111 *
0-
02
b111 6
#955030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#955040000000
0!
0%
b0 *
0-
02
b0 6
#955050000000
1!
1%
1-
12
#955060000000
0!
0%
b1 *
0-
02
b1 6
#955070000000
1!
1%
1-
12
#955080000000
0!
0%
b10 *
0-
02
b10 6
#955090000000
1!
1%
1-
12
#955100000000
0!
0%
b11 *
0-
02
b11 6
#955110000000
1!
1%
1-
12
15
#955120000000
0!
0%
b100 *
0-
02
b100 6
#955130000000
1!
1%
1-
12
#955140000000
0!
0%
b101 *
0-
02
b101 6
#955150000000
1!
1%
1-
12
#955160000000
0!
0%
b110 *
0-
02
b110 6
#955170000000
1!
1%
1-
12
#955180000000
0!
0%
b111 *
0-
02
b111 6
#955190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#955200000000
0!
0%
b0 *
0-
02
b0 6
#955210000000
1!
1%
1-
12
#955220000000
0!
0%
b1 *
0-
02
b1 6
#955230000000
1!
1%
1-
12
#955240000000
0!
0%
b10 *
0-
02
b10 6
#955250000000
1!
1%
1-
12
#955260000000
0!
0%
b11 *
0-
02
b11 6
#955270000000
1!
1%
1-
12
15
#955280000000
0!
0%
b100 *
0-
02
b100 6
#955290000000
1!
1%
1-
12
#955300000000
0!
0%
b101 *
0-
02
b101 6
#955310000000
1!
1%
1-
12
#955320000000
0!
0%
b110 *
0-
02
b110 6
#955330000000
1!
1%
1-
12
#955340000000
0!
0%
b111 *
0-
02
b111 6
#955350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#955360000000
0!
0%
b0 *
0-
02
b0 6
#955370000000
1!
1%
1-
12
#955380000000
0!
0%
b1 *
0-
02
b1 6
#955390000000
1!
1%
1-
12
#955400000000
0!
0%
b10 *
0-
02
b10 6
#955410000000
1!
1%
1-
12
#955420000000
0!
0%
b11 *
0-
02
b11 6
#955430000000
1!
1%
1-
12
15
#955440000000
0!
0%
b100 *
0-
02
b100 6
#955450000000
1!
1%
1-
12
#955460000000
0!
0%
b101 *
0-
02
b101 6
#955470000000
1!
1%
1-
12
#955480000000
0!
0%
b110 *
0-
02
b110 6
#955490000000
1!
1%
1-
12
#955500000000
0!
0%
b111 *
0-
02
b111 6
#955510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#955520000000
0!
0%
b0 *
0-
02
b0 6
#955530000000
1!
1%
1-
12
#955540000000
0!
0%
b1 *
0-
02
b1 6
#955550000000
1!
1%
1-
12
#955560000000
0!
0%
b10 *
0-
02
b10 6
#955570000000
1!
1%
1-
12
#955580000000
0!
0%
b11 *
0-
02
b11 6
#955590000000
1!
1%
1-
12
15
#955600000000
0!
0%
b100 *
0-
02
b100 6
#955610000000
1!
1%
1-
12
#955620000000
0!
0%
b101 *
0-
02
b101 6
#955630000000
1!
1%
1-
12
#955640000000
0!
0%
b110 *
0-
02
b110 6
#955650000000
1!
1%
1-
12
#955660000000
0!
0%
b111 *
0-
02
b111 6
#955670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#955680000000
0!
0%
b0 *
0-
02
b0 6
#955690000000
1!
1%
1-
12
#955700000000
0!
0%
b1 *
0-
02
b1 6
#955710000000
1!
1%
1-
12
#955720000000
0!
0%
b10 *
0-
02
b10 6
#955730000000
1!
1%
1-
12
#955740000000
0!
0%
b11 *
0-
02
b11 6
#955750000000
1!
1%
1-
12
15
#955760000000
0!
0%
b100 *
0-
02
b100 6
#955770000000
1!
1%
1-
12
#955780000000
0!
0%
b101 *
0-
02
b101 6
#955790000000
1!
1%
1-
12
#955800000000
0!
0%
b110 *
0-
02
b110 6
#955810000000
1!
1%
1-
12
#955820000000
0!
0%
b111 *
0-
02
b111 6
#955830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#955840000000
0!
0%
b0 *
0-
02
b0 6
#955850000000
1!
1%
1-
12
#955860000000
0!
0%
b1 *
0-
02
b1 6
#955870000000
1!
1%
1-
12
#955880000000
0!
0%
b10 *
0-
02
b10 6
#955890000000
1!
1%
1-
12
#955900000000
0!
0%
b11 *
0-
02
b11 6
#955910000000
1!
1%
1-
12
15
#955920000000
0!
0%
b100 *
0-
02
b100 6
#955930000000
1!
1%
1-
12
#955940000000
0!
0%
b101 *
0-
02
b101 6
#955950000000
1!
1%
1-
12
#955960000000
0!
0%
b110 *
0-
02
b110 6
#955970000000
1!
1%
1-
12
#955980000000
0!
0%
b111 *
0-
02
b111 6
#955990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#956000000000
0!
0%
b0 *
0-
02
b0 6
#956010000000
1!
1%
1-
12
#956020000000
0!
0%
b1 *
0-
02
b1 6
#956030000000
1!
1%
1-
12
#956040000000
0!
0%
b10 *
0-
02
b10 6
#956050000000
1!
1%
1-
12
#956060000000
0!
0%
b11 *
0-
02
b11 6
#956070000000
1!
1%
1-
12
15
#956080000000
0!
0%
b100 *
0-
02
b100 6
#956090000000
1!
1%
1-
12
#956100000000
0!
0%
b101 *
0-
02
b101 6
#956110000000
1!
1%
1-
12
#956120000000
0!
0%
b110 *
0-
02
b110 6
#956130000000
1!
1%
1-
12
#956140000000
0!
0%
b111 *
0-
02
b111 6
#956150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#956160000000
0!
0%
b0 *
0-
02
b0 6
#956170000000
1!
1%
1-
12
#956180000000
0!
0%
b1 *
0-
02
b1 6
#956190000000
1!
1%
1-
12
#956200000000
0!
0%
b10 *
0-
02
b10 6
#956210000000
1!
1%
1-
12
#956220000000
0!
0%
b11 *
0-
02
b11 6
#956230000000
1!
1%
1-
12
15
#956240000000
0!
0%
b100 *
0-
02
b100 6
#956250000000
1!
1%
1-
12
#956260000000
0!
0%
b101 *
0-
02
b101 6
#956270000000
1!
1%
1-
12
#956280000000
0!
0%
b110 *
0-
02
b110 6
#956290000000
1!
1%
1-
12
#956300000000
0!
0%
b111 *
0-
02
b111 6
#956310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#956320000000
0!
0%
b0 *
0-
02
b0 6
#956330000000
1!
1%
1-
12
#956340000000
0!
0%
b1 *
0-
02
b1 6
#956350000000
1!
1%
1-
12
#956360000000
0!
0%
b10 *
0-
02
b10 6
#956370000000
1!
1%
1-
12
#956380000000
0!
0%
b11 *
0-
02
b11 6
#956390000000
1!
1%
1-
12
15
#956400000000
0!
0%
b100 *
0-
02
b100 6
#956410000000
1!
1%
1-
12
#956420000000
0!
0%
b101 *
0-
02
b101 6
#956430000000
1!
1%
1-
12
#956440000000
0!
0%
b110 *
0-
02
b110 6
#956450000000
1!
1%
1-
12
#956460000000
0!
0%
b111 *
0-
02
b111 6
#956470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#956480000000
0!
0%
b0 *
0-
02
b0 6
#956490000000
1!
1%
1-
12
#956500000000
0!
0%
b1 *
0-
02
b1 6
#956510000000
1!
1%
1-
12
#956520000000
0!
0%
b10 *
0-
02
b10 6
#956530000000
1!
1%
1-
12
#956540000000
0!
0%
b11 *
0-
02
b11 6
#956550000000
1!
1%
1-
12
15
#956560000000
0!
0%
b100 *
0-
02
b100 6
#956570000000
1!
1%
1-
12
#956580000000
0!
0%
b101 *
0-
02
b101 6
#956590000000
1!
1%
1-
12
#956600000000
0!
0%
b110 *
0-
02
b110 6
#956610000000
1!
1%
1-
12
#956620000000
0!
0%
b111 *
0-
02
b111 6
#956630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#956640000000
0!
0%
b0 *
0-
02
b0 6
#956650000000
1!
1%
1-
12
#956660000000
0!
0%
b1 *
0-
02
b1 6
#956670000000
1!
1%
1-
12
#956680000000
0!
0%
b10 *
0-
02
b10 6
#956690000000
1!
1%
1-
12
#956700000000
0!
0%
b11 *
0-
02
b11 6
#956710000000
1!
1%
1-
12
15
#956720000000
0!
0%
b100 *
0-
02
b100 6
#956730000000
1!
1%
1-
12
#956740000000
0!
0%
b101 *
0-
02
b101 6
#956750000000
1!
1%
1-
12
#956760000000
0!
0%
b110 *
0-
02
b110 6
#956770000000
1!
1%
1-
12
#956780000000
0!
0%
b111 *
0-
02
b111 6
#956790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#956800000000
0!
0%
b0 *
0-
02
b0 6
#956810000000
1!
1%
1-
12
#956820000000
0!
0%
b1 *
0-
02
b1 6
#956830000000
1!
1%
1-
12
#956840000000
0!
0%
b10 *
0-
02
b10 6
#956850000000
1!
1%
1-
12
#956860000000
0!
0%
b11 *
0-
02
b11 6
#956870000000
1!
1%
1-
12
15
#956880000000
0!
0%
b100 *
0-
02
b100 6
#956890000000
1!
1%
1-
12
#956900000000
0!
0%
b101 *
0-
02
b101 6
#956910000000
1!
1%
1-
12
#956920000000
0!
0%
b110 *
0-
02
b110 6
#956930000000
1!
1%
1-
12
#956940000000
0!
0%
b111 *
0-
02
b111 6
#956950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#956960000000
0!
0%
b0 *
0-
02
b0 6
#956970000000
1!
1%
1-
12
#956980000000
0!
0%
b1 *
0-
02
b1 6
#956990000000
1!
1%
1-
12
#957000000000
0!
0%
b10 *
0-
02
b10 6
#957010000000
1!
1%
1-
12
#957020000000
0!
0%
b11 *
0-
02
b11 6
#957030000000
1!
1%
1-
12
15
#957040000000
0!
0%
b100 *
0-
02
b100 6
#957050000000
1!
1%
1-
12
#957060000000
0!
0%
b101 *
0-
02
b101 6
#957070000000
1!
1%
1-
12
#957080000000
0!
0%
b110 *
0-
02
b110 6
#957090000000
1!
1%
1-
12
#957100000000
0!
0%
b111 *
0-
02
b111 6
#957110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#957120000000
0!
0%
b0 *
0-
02
b0 6
#957130000000
1!
1%
1-
12
#957140000000
0!
0%
b1 *
0-
02
b1 6
#957150000000
1!
1%
1-
12
#957160000000
0!
0%
b10 *
0-
02
b10 6
#957170000000
1!
1%
1-
12
#957180000000
0!
0%
b11 *
0-
02
b11 6
#957190000000
1!
1%
1-
12
15
#957200000000
0!
0%
b100 *
0-
02
b100 6
#957210000000
1!
1%
1-
12
#957220000000
0!
0%
b101 *
0-
02
b101 6
#957230000000
1!
1%
1-
12
#957240000000
0!
0%
b110 *
0-
02
b110 6
#957250000000
1!
1%
1-
12
#957260000000
0!
0%
b111 *
0-
02
b111 6
#957270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#957280000000
0!
0%
b0 *
0-
02
b0 6
#957290000000
1!
1%
1-
12
#957300000000
0!
0%
b1 *
0-
02
b1 6
#957310000000
1!
1%
1-
12
#957320000000
0!
0%
b10 *
0-
02
b10 6
#957330000000
1!
1%
1-
12
#957340000000
0!
0%
b11 *
0-
02
b11 6
#957350000000
1!
1%
1-
12
15
#957360000000
0!
0%
b100 *
0-
02
b100 6
#957370000000
1!
1%
1-
12
#957380000000
0!
0%
b101 *
0-
02
b101 6
#957390000000
1!
1%
1-
12
#957400000000
0!
0%
b110 *
0-
02
b110 6
#957410000000
1!
1%
1-
12
#957420000000
0!
0%
b111 *
0-
02
b111 6
#957430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#957440000000
0!
0%
b0 *
0-
02
b0 6
#957450000000
1!
1%
1-
12
#957460000000
0!
0%
b1 *
0-
02
b1 6
#957470000000
1!
1%
1-
12
#957480000000
0!
0%
b10 *
0-
02
b10 6
#957490000000
1!
1%
1-
12
#957500000000
0!
0%
b11 *
0-
02
b11 6
#957510000000
1!
1%
1-
12
15
#957520000000
0!
0%
b100 *
0-
02
b100 6
#957530000000
1!
1%
1-
12
#957540000000
0!
0%
b101 *
0-
02
b101 6
#957550000000
1!
1%
1-
12
#957560000000
0!
0%
b110 *
0-
02
b110 6
#957570000000
1!
1%
1-
12
#957580000000
0!
0%
b111 *
0-
02
b111 6
#957590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#957600000000
0!
0%
b0 *
0-
02
b0 6
#957610000000
1!
1%
1-
12
#957620000000
0!
0%
b1 *
0-
02
b1 6
#957630000000
1!
1%
1-
12
#957640000000
0!
0%
b10 *
0-
02
b10 6
#957650000000
1!
1%
1-
12
#957660000000
0!
0%
b11 *
0-
02
b11 6
#957670000000
1!
1%
1-
12
15
#957680000000
0!
0%
b100 *
0-
02
b100 6
#957690000000
1!
1%
1-
12
#957700000000
0!
0%
b101 *
0-
02
b101 6
#957710000000
1!
1%
1-
12
#957720000000
0!
0%
b110 *
0-
02
b110 6
#957730000000
1!
1%
1-
12
#957740000000
0!
0%
b111 *
0-
02
b111 6
#957750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#957760000000
0!
0%
b0 *
0-
02
b0 6
#957770000000
1!
1%
1-
12
#957780000000
0!
0%
b1 *
0-
02
b1 6
#957790000000
1!
1%
1-
12
#957800000000
0!
0%
b10 *
0-
02
b10 6
#957810000000
1!
1%
1-
12
#957820000000
0!
0%
b11 *
0-
02
b11 6
#957830000000
1!
1%
1-
12
15
#957840000000
0!
0%
b100 *
0-
02
b100 6
#957850000000
1!
1%
1-
12
#957860000000
0!
0%
b101 *
0-
02
b101 6
#957870000000
1!
1%
1-
12
#957880000000
0!
0%
b110 *
0-
02
b110 6
#957890000000
1!
1%
1-
12
#957900000000
0!
0%
b111 *
0-
02
b111 6
#957910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#957920000000
0!
0%
b0 *
0-
02
b0 6
#957930000000
1!
1%
1-
12
#957940000000
0!
0%
b1 *
0-
02
b1 6
#957950000000
1!
1%
1-
12
#957960000000
0!
0%
b10 *
0-
02
b10 6
#957970000000
1!
1%
1-
12
#957980000000
0!
0%
b11 *
0-
02
b11 6
#957990000000
1!
1%
1-
12
15
#958000000000
0!
0%
b100 *
0-
02
b100 6
#958010000000
1!
1%
1-
12
#958020000000
0!
0%
b101 *
0-
02
b101 6
#958030000000
1!
1%
1-
12
#958040000000
0!
0%
b110 *
0-
02
b110 6
#958050000000
1!
1%
1-
12
#958060000000
0!
0%
b111 *
0-
02
b111 6
#958070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#958080000000
0!
0%
b0 *
0-
02
b0 6
#958090000000
1!
1%
1-
12
#958100000000
0!
0%
b1 *
0-
02
b1 6
#958110000000
1!
1%
1-
12
#958120000000
0!
0%
b10 *
0-
02
b10 6
#958130000000
1!
1%
1-
12
#958140000000
0!
0%
b11 *
0-
02
b11 6
#958150000000
1!
1%
1-
12
15
#958160000000
0!
0%
b100 *
0-
02
b100 6
#958170000000
1!
1%
1-
12
#958180000000
0!
0%
b101 *
0-
02
b101 6
#958190000000
1!
1%
1-
12
#958200000000
0!
0%
b110 *
0-
02
b110 6
#958210000000
1!
1%
1-
12
#958220000000
0!
0%
b111 *
0-
02
b111 6
#958230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#958240000000
0!
0%
b0 *
0-
02
b0 6
#958250000000
1!
1%
1-
12
#958260000000
0!
0%
b1 *
0-
02
b1 6
#958270000000
1!
1%
1-
12
#958280000000
0!
0%
b10 *
0-
02
b10 6
#958290000000
1!
1%
1-
12
#958300000000
0!
0%
b11 *
0-
02
b11 6
#958310000000
1!
1%
1-
12
15
#958320000000
0!
0%
b100 *
0-
02
b100 6
#958330000000
1!
1%
1-
12
#958340000000
0!
0%
b101 *
0-
02
b101 6
#958350000000
1!
1%
1-
12
#958360000000
0!
0%
b110 *
0-
02
b110 6
#958370000000
1!
1%
1-
12
#958380000000
0!
0%
b111 *
0-
02
b111 6
#958390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#958400000000
0!
0%
b0 *
0-
02
b0 6
#958410000000
1!
1%
1-
12
#958420000000
0!
0%
b1 *
0-
02
b1 6
#958430000000
1!
1%
1-
12
#958440000000
0!
0%
b10 *
0-
02
b10 6
#958450000000
1!
1%
1-
12
#958460000000
0!
0%
b11 *
0-
02
b11 6
#958470000000
1!
1%
1-
12
15
#958480000000
0!
0%
b100 *
0-
02
b100 6
#958490000000
1!
1%
1-
12
#958500000000
0!
0%
b101 *
0-
02
b101 6
#958510000000
1!
1%
1-
12
#958520000000
0!
0%
b110 *
0-
02
b110 6
#958530000000
1!
1%
1-
12
#958540000000
0!
0%
b111 *
0-
02
b111 6
#958550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#958560000000
0!
0%
b0 *
0-
02
b0 6
#958570000000
1!
1%
1-
12
#958580000000
0!
0%
b1 *
0-
02
b1 6
#958590000000
1!
1%
1-
12
#958600000000
0!
0%
b10 *
0-
02
b10 6
#958610000000
1!
1%
1-
12
#958620000000
0!
0%
b11 *
0-
02
b11 6
#958630000000
1!
1%
1-
12
15
#958640000000
0!
0%
b100 *
0-
02
b100 6
#958650000000
1!
1%
1-
12
#958660000000
0!
0%
b101 *
0-
02
b101 6
#958670000000
1!
1%
1-
12
#958680000000
0!
0%
b110 *
0-
02
b110 6
#958690000000
1!
1%
1-
12
#958700000000
0!
0%
b111 *
0-
02
b111 6
#958710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#958720000000
0!
0%
b0 *
0-
02
b0 6
#958730000000
1!
1%
1-
12
#958740000000
0!
0%
b1 *
0-
02
b1 6
#958750000000
1!
1%
1-
12
#958760000000
0!
0%
b10 *
0-
02
b10 6
#958770000000
1!
1%
1-
12
#958780000000
0!
0%
b11 *
0-
02
b11 6
#958790000000
1!
1%
1-
12
15
#958800000000
0!
0%
b100 *
0-
02
b100 6
#958810000000
1!
1%
1-
12
#958820000000
0!
0%
b101 *
0-
02
b101 6
#958830000000
1!
1%
1-
12
#958840000000
0!
0%
b110 *
0-
02
b110 6
#958850000000
1!
1%
1-
12
#958860000000
0!
0%
b111 *
0-
02
b111 6
#958870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#958880000000
0!
0%
b0 *
0-
02
b0 6
#958890000000
1!
1%
1-
12
#958900000000
0!
0%
b1 *
0-
02
b1 6
#958910000000
1!
1%
1-
12
#958920000000
0!
0%
b10 *
0-
02
b10 6
#958930000000
1!
1%
1-
12
#958940000000
0!
0%
b11 *
0-
02
b11 6
#958950000000
1!
1%
1-
12
15
#958960000000
0!
0%
b100 *
0-
02
b100 6
#958970000000
1!
1%
1-
12
#958980000000
0!
0%
b101 *
0-
02
b101 6
#958990000000
1!
1%
1-
12
#959000000000
0!
0%
b110 *
0-
02
b110 6
#959010000000
1!
1%
1-
12
#959020000000
0!
0%
b111 *
0-
02
b111 6
#959030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#959040000000
0!
0%
b0 *
0-
02
b0 6
#959050000000
1!
1%
1-
12
#959060000000
0!
0%
b1 *
0-
02
b1 6
#959070000000
1!
1%
1-
12
#959080000000
0!
0%
b10 *
0-
02
b10 6
#959090000000
1!
1%
1-
12
#959100000000
0!
0%
b11 *
0-
02
b11 6
#959110000000
1!
1%
1-
12
15
#959120000000
0!
0%
b100 *
0-
02
b100 6
#959130000000
1!
1%
1-
12
#959140000000
0!
0%
b101 *
0-
02
b101 6
#959150000000
1!
1%
1-
12
#959160000000
0!
0%
b110 *
0-
02
b110 6
#959170000000
1!
1%
1-
12
#959180000000
0!
0%
b111 *
0-
02
b111 6
#959190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#959200000000
0!
0%
b0 *
0-
02
b0 6
#959210000000
1!
1%
1-
12
#959220000000
0!
0%
b1 *
0-
02
b1 6
#959230000000
1!
1%
1-
12
#959240000000
0!
0%
b10 *
0-
02
b10 6
#959250000000
1!
1%
1-
12
#959260000000
0!
0%
b11 *
0-
02
b11 6
#959270000000
1!
1%
1-
12
15
#959280000000
0!
0%
b100 *
0-
02
b100 6
#959290000000
1!
1%
1-
12
#959300000000
0!
0%
b101 *
0-
02
b101 6
#959310000000
1!
1%
1-
12
#959320000000
0!
0%
b110 *
0-
02
b110 6
#959330000000
1!
1%
1-
12
#959340000000
0!
0%
b111 *
0-
02
b111 6
#959350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#959360000000
0!
0%
b0 *
0-
02
b0 6
#959370000000
1!
1%
1-
12
#959380000000
0!
0%
b1 *
0-
02
b1 6
#959390000000
1!
1%
1-
12
#959400000000
0!
0%
b10 *
0-
02
b10 6
#959410000000
1!
1%
1-
12
#959420000000
0!
0%
b11 *
0-
02
b11 6
#959430000000
1!
1%
1-
12
15
#959440000000
0!
0%
b100 *
0-
02
b100 6
#959450000000
1!
1%
1-
12
#959460000000
0!
0%
b101 *
0-
02
b101 6
#959470000000
1!
1%
1-
12
#959480000000
0!
0%
b110 *
0-
02
b110 6
#959490000000
1!
1%
1-
12
#959500000000
0!
0%
b111 *
0-
02
b111 6
#959510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#959520000000
0!
0%
b0 *
0-
02
b0 6
#959530000000
1!
1%
1-
12
#959540000000
0!
0%
b1 *
0-
02
b1 6
#959550000000
1!
1%
1-
12
#959560000000
0!
0%
b10 *
0-
02
b10 6
#959570000000
1!
1%
1-
12
#959580000000
0!
0%
b11 *
0-
02
b11 6
#959590000000
1!
1%
1-
12
15
#959600000000
0!
0%
b100 *
0-
02
b100 6
#959610000000
1!
1%
1-
12
#959620000000
0!
0%
b101 *
0-
02
b101 6
#959630000000
1!
1%
1-
12
#959640000000
0!
0%
b110 *
0-
02
b110 6
#959650000000
1!
1%
1-
12
#959660000000
0!
0%
b111 *
0-
02
b111 6
#959670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#959680000000
0!
0%
b0 *
0-
02
b0 6
#959690000000
1!
1%
1-
12
#959700000000
0!
0%
b1 *
0-
02
b1 6
#959710000000
1!
1%
1-
12
#959720000000
0!
0%
b10 *
0-
02
b10 6
#959730000000
1!
1%
1-
12
#959740000000
0!
0%
b11 *
0-
02
b11 6
#959750000000
1!
1%
1-
12
15
#959760000000
0!
0%
b100 *
0-
02
b100 6
#959770000000
1!
1%
1-
12
#959780000000
0!
0%
b101 *
0-
02
b101 6
#959790000000
1!
1%
1-
12
#959800000000
0!
0%
b110 *
0-
02
b110 6
#959810000000
1!
1%
1-
12
#959820000000
0!
0%
b111 *
0-
02
b111 6
#959830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#959840000000
0!
0%
b0 *
0-
02
b0 6
#959850000000
1!
1%
1-
12
#959860000000
0!
0%
b1 *
0-
02
b1 6
#959870000000
1!
1%
1-
12
#959880000000
0!
0%
b10 *
0-
02
b10 6
#959890000000
1!
1%
1-
12
#959900000000
0!
0%
b11 *
0-
02
b11 6
#959910000000
1!
1%
1-
12
15
#959920000000
0!
0%
b100 *
0-
02
b100 6
#959930000000
1!
1%
1-
12
#959940000000
0!
0%
b101 *
0-
02
b101 6
#959950000000
1!
1%
1-
12
#959960000000
0!
0%
b110 *
0-
02
b110 6
#959970000000
1!
1%
1-
12
#959980000000
0!
0%
b111 *
0-
02
b111 6
#959990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#960000000000
0!
0%
b0 *
0-
02
b0 6
#960010000000
1!
1%
1-
12
#960020000000
0!
0%
b1 *
0-
02
b1 6
#960030000000
1!
1%
1-
12
#960040000000
0!
0%
b10 *
0-
02
b10 6
#960050000000
1!
1%
1-
12
#960060000000
0!
0%
b11 *
0-
02
b11 6
#960070000000
1!
1%
1-
12
15
#960080000000
0!
0%
b100 *
0-
02
b100 6
#960090000000
1!
1%
1-
12
#960100000000
0!
0%
b101 *
0-
02
b101 6
#960110000000
1!
1%
1-
12
#960120000000
0!
0%
b110 *
0-
02
b110 6
#960130000000
1!
1%
1-
12
#960140000000
0!
0%
b111 *
0-
02
b111 6
#960150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#960160000000
0!
0%
b0 *
0-
02
b0 6
#960170000000
1!
1%
1-
12
#960180000000
0!
0%
b1 *
0-
02
b1 6
#960190000000
1!
1%
1-
12
#960200000000
0!
0%
b10 *
0-
02
b10 6
#960210000000
1!
1%
1-
12
#960220000000
0!
0%
b11 *
0-
02
b11 6
#960230000000
1!
1%
1-
12
15
#960240000000
0!
0%
b100 *
0-
02
b100 6
#960250000000
1!
1%
1-
12
#960260000000
0!
0%
b101 *
0-
02
b101 6
#960270000000
1!
1%
1-
12
#960280000000
0!
0%
b110 *
0-
02
b110 6
#960290000000
1!
1%
1-
12
#960300000000
0!
0%
b111 *
0-
02
b111 6
#960310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#960320000000
0!
0%
b0 *
0-
02
b0 6
#960330000000
1!
1%
1-
12
#960340000000
0!
0%
b1 *
0-
02
b1 6
#960350000000
1!
1%
1-
12
#960360000000
0!
0%
b10 *
0-
02
b10 6
#960370000000
1!
1%
1-
12
#960380000000
0!
0%
b11 *
0-
02
b11 6
#960390000000
1!
1%
1-
12
15
#960400000000
0!
0%
b100 *
0-
02
b100 6
#960410000000
1!
1%
1-
12
#960420000000
0!
0%
b101 *
0-
02
b101 6
#960430000000
1!
1%
1-
12
#960440000000
0!
0%
b110 *
0-
02
b110 6
#960450000000
1!
1%
1-
12
#960460000000
0!
0%
b111 *
0-
02
b111 6
#960470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#960480000000
0!
0%
b0 *
0-
02
b0 6
#960490000000
1!
1%
1-
12
#960500000000
0!
0%
b1 *
0-
02
b1 6
#960510000000
1!
1%
1-
12
#960520000000
0!
0%
b10 *
0-
02
b10 6
#960530000000
1!
1%
1-
12
#960540000000
0!
0%
b11 *
0-
02
b11 6
#960550000000
1!
1%
1-
12
15
#960560000000
0!
0%
b100 *
0-
02
b100 6
#960570000000
1!
1%
1-
12
#960580000000
0!
0%
b101 *
0-
02
b101 6
#960590000000
1!
1%
1-
12
#960600000000
0!
0%
b110 *
0-
02
b110 6
#960610000000
1!
1%
1-
12
#960620000000
0!
0%
b111 *
0-
02
b111 6
#960630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#960640000000
0!
0%
b0 *
0-
02
b0 6
#960650000000
1!
1%
1-
12
#960660000000
0!
0%
b1 *
0-
02
b1 6
#960670000000
1!
1%
1-
12
#960680000000
0!
0%
b10 *
0-
02
b10 6
#960690000000
1!
1%
1-
12
#960700000000
0!
0%
b11 *
0-
02
b11 6
#960710000000
1!
1%
1-
12
15
#960720000000
0!
0%
b100 *
0-
02
b100 6
#960730000000
1!
1%
1-
12
#960740000000
0!
0%
b101 *
0-
02
b101 6
#960750000000
1!
1%
1-
12
#960760000000
0!
0%
b110 *
0-
02
b110 6
#960770000000
1!
1%
1-
12
#960780000000
0!
0%
b111 *
0-
02
b111 6
#960790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#960800000000
0!
0%
b0 *
0-
02
b0 6
#960810000000
1!
1%
1-
12
#960820000000
0!
0%
b1 *
0-
02
b1 6
#960830000000
1!
1%
1-
12
#960840000000
0!
0%
b10 *
0-
02
b10 6
#960850000000
1!
1%
1-
12
#960860000000
0!
0%
b11 *
0-
02
b11 6
#960870000000
1!
1%
1-
12
15
#960880000000
0!
0%
b100 *
0-
02
b100 6
#960890000000
1!
1%
1-
12
#960900000000
0!
0%
b101 *
0-
02
b101 6
#960910000000
1!
1%
1-
12
#960920000000
0!
0%
b110 *
0-
02
b110 6
#960930000000
1!
1%
1-
12
#960940000000
0!
0%
b111 *
0-
02
b111 6
#960950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#960960000000
0!
0%
b0 *
0-
02
b0 6
#960970000000
1!
1%
1-
12
#960980000000
0!
0%
b1 *
0-
02
b1 6
#960990000000
1!
1%
1-
12
#961000000000
0!
0%
b10 *
0-
02
b10 6
#961010000000
1!
1%
1-
12
#961020000000
0!
0%
b11 *
0-
02
b11 6
#961030000000
1!
1%
1-
12
15
#961040000000
0!
0%
b100 *
0-
02
b100 6
#961050000000
1!
1%
1-
12
#961060000000
0!
0%
b101 *
0-
02
b101 6
#961070000000
1!
1%
1-
12
#961080000000
0!
0%
b110 *
0-
02
b110 6
#961090000000
1!
1%
1-
12
#961100000000
0!
0%
b111 *
0-
02
b111 6
#961110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#961120000000
0!
0%
b0 *
0-
02
b0 6
#961130000000
1!
1%
1-
12
#961140000000
0!
0%
b1 *
0-
02
b1 6
#961150000000
1!
1%
1-
12
#961160000000
0!
0%
b10 *
0-
02
b10 6
#961170000000
1!
1%
1-
12
#961180000000
0!
0%
b11 *
0-
02
b11 6
#961190000000
1!
1%
1-
12
15
#961200000000
0!
0%
b100 *
0-
02
b100 6
#961210000000
1!
1%
1-
12
#961220000000
0!
0%
b101 *
0-
02
b101 6
#961230000000
1!
1%
1-
12
#961240000000
0!
0%
b110 *
0-
02
b110 6
#961250000000
1!
1%
1-
12
#961260000000
0!
0%
b111 *
0-
02
b111 6
#961270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#961280000000
0!
0%
b0 *
0-
02
b0 6
#961290000000
1!
1%
1-
12
#961300000000
0!
0%
b1 *
0-
02
b1 6
#961310000000
1!
1%
1-
12
#961320000000
0!
0%
b10 *
0-
02
b10 6
#961330000000
1!
1%
1-
12
#961340000000
0!
0%
b11 *
0-
02
b11 6
#961350000000
1!
1%
1-
12
15
#961360000000
0!
0%
b100 *
0-
02
b100 6
#961370000000
1!
1%
1-
12
#961380000000
0!
0%
b101 *
0-
02
b101 6
#961390000000
1!
1%
1-
12
#961400000000
0!
0%
b110 *
0-
02
b110 6
#961410000000
1!
1%
1-
12
#961420000000
0!
0%
b111 *
0-
02
b111 6
#961430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#961440000000
0!
0%
b0 *
0-
02
b0 6
#961450000000
1!
1%
1-
12
#961460000000
0!
0%
b1 *
0-
02
b1 6
#961470000000
1!
1%
1-
12
#961480000000
0!
0%
b10 *
0-
02
b10 6
#961490000000
1!
1%
1-
12
#961500000000
0!
0%
b11 *
0-
02
b11 6
#961510000000
1!
1%
1-
12
15
#961520000000
0!
0%
b100 *
0-
02
b100 6
#961530000000
1!
1%
1-
12
#961540000000
0!
0%
b101 *
0-
02
b101 6
#961550000000
1!
1%
1-
12
#961560000000
0!
0%
b110 *
0-
02
b110 6
#961570000000
1!
1%
1-
12
#961580000000
0!
0%
b111 *
0-
02
b111 6
#961590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#961600000000
0!
0%
b0 *
0-
02
b0 6
#961610000000
1!
1%
1-
12
#961620000000
0!
0%
b1 *
0-
02
b1 6
#961630000000
1!
1%
1-
12
#961640000000
0!
0%
b10 *
0-
02
b10 6
#961650000000
1!
1%
1-
12
#961660000000
0!
0%
b11 *
0-
02
b11 6
#961670000000
1!
1%
1-
12
15
#961680000000
0!
0%
b100 *
0-
02
b100 6
#961690000000
1!
1%
1-
12
#961700000000
0!
0%
b101 *
0-
02
b101 6
#961710000000
1!
1%
1-
12
#961720000000
0!
0%
b110 *
0-
02
b110 6
#961730000000
1!
1%
1-
12
#961740000000
0!
0%
b111 *
0-
02
b111 6
#961750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#961760000000
0!
0%
b0 *
0-
02
b0 6
#961770000000
1!
1%
1-
12
#961780000000
0!
0%
b1 *
0-
02
b1 6
#961790000000
1!
1%
1-
12
#961800000000
0!
0%
b10 *
0-
02
b10 6
#961810000000
1!
1%
1-
12
#961820000000
0!
0%
b11 *
0-
02
b11 6
#961830000000
1!
1%
1-
12
15
#961840000000
0!
0%
b100 *
0-
02
b100 6
#961850000000
1!
1%
1-
12
#961860000000
0!
0%
b101 *
0-
02
b101 6
#961870000000
1!
1%
1-
12
#961880000000
0!
0%
b110 *
0-
02
b110 6
#961890000000
1!
1%
1-
12
#961900000000
0!
0%
b111 *
0-
02
b111 6
#961910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#961920000000
0!
0%
b0 *
0-
02
b0 6
#961930000000
1!
1%
1-
12
#961940000000
0!
0%
b1 *
0-
02
b1 6
#961950000000
1!
1%
1-
12
#961960000000
0!
0%
b10 *
0-
02
b10 6
#961970000000
1!
1%
1-
12
#961980000000
0!
0%
b11 *
0-
02
b11 6
#961990000000
1!
1%
1-
12
15
#962000000000
0!
0%
b100 *
0-
02
b100 6
#962010000000
1!
1%
1-
12
#962020000000
0!
0%
b101 *
0-
02
b101 6
#962030000000
1!
1%
1-
12
#962040000000
0!
0%
b110 *
0-
02
b110 6
#962050000000
1!
1%
1-
12
#962060000000
0!
0%
b111 *
0-
02
b111 6
#962070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#962080000000
0!
0%
b0 *
0-
02
b0 6
#962090000000
1!
1%
1-
12
#962100000000
0!
0%
b1 *
0-
02
b1 6
#962110000000
1!
1%
1-
12
#962120000000
0!
0%
b10 *
0-
02
b10 6
#962130000000
1!
1%
1-
12
#962140000000
0!
0%
b11 *
0-
02
b11 6
#962150000000
1!
1%
1-
12
15
#962160000000
0!
0%
b100 *
0-
02
b100 6
#962170000000
1!
1%
1-
12
#962180000000
0!
0%
b101 *
0-
02
b101 6
#962190000000
1!
1%
1-
12
#962200000000
0!
0%
b110 *
0-
02
b110 6
#962210000000
1!
1%
1-
12
#962220000000
0!
0%
b111 *
0-
02
b111 6
#962230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#962240000000
0!
0%
b0 *
0-
02
b0 6
#962250000000
1!
1%
1-
12
#962260000000
0!
0%
b1 *
0-
02
b1 6
#962270000000
1!
1%
1-
12
#962280000000
0!
0%
b10 *
0-
02
b10 6
#962290000000
1!
1%
1-
12
#962300000000
0!
0%
b11 *
0-
02
b11 6
#962310000000
1!
1%
1-
12
15
#962320000000
0!
0%
b100 *
0-
02
b100 6
#962330000000
1!
1%
1-
12
#962340000000
0!
0%
b101 *
0-
02
b101 6
#962350000000
1!
1%
1-
12
#962360000000
0!
0%
b110 *
0-
02
b110 6
#962370000000
1!
1%
1-
12
#962380000000
0!
0%
b111 *
0-
02
b111 6
#962390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#962400000000
0!
0%
b0 *
0-
02
b0 6
#962410000000
1!
1%
1-
12
#962420000000
0!
0%
b1 *
0-
02
b1 6
#962430000000
1!
1%
1-
12
#962440000000
0!
0%
b10 *
0-
02
b10 6
#962450000000
1!
1%
1-
12
#962460000000
0!
0%
b11 *
0-
02
b11 6
#962470000000
1!
1%
1-
12
15
#962480000000
0!
0%
b100 *
0-
02
b100 6
#962490000000
1!
1%
1-
12
#962500000000
0!
0%
b101 *
0-
02
b101 6
#962510000000
1!
1%
1-
12
#962520000000
0!
0%
b110 *
0-
02
b110 6
#962530000000
1!
1%
1-
12
#962540000000
0!
0%
b111 *
0-
02
b111 6
#962550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#962560000000
0!
0%
b0 *
0-
02
b0 6
#962570000000
1!
1%
1-
12
#962580000000
0!
0%
b1 *
0-
02
b1 6
#962590000000
1!
1%
1-
12
#962600000000
0!
0%
b10 *
0-
02
b10 6
#962610000000
1!
1%
1-
12
#962620000000
0!
0%
b11 *
0-
02
b11 6
#962630000000
1!
1%
1-
12
15
#962640000000
0!
0%
b100 *
0-
02
b100 6
#962650000000
1!
1%
1-
12
#962660000000
0!
0%
b101 *
0-
02
b101 6
#962670000000
1!
1%
1-
12
#962680000000
0!
0%
b110 *
0-
02
b110 6
#962690000000
1!
1%
1-
12
#962700000000
0!
0%
b111 *
0-
02
b111 6
#962710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#962720000000
0!
0%
b0 *
0-
02
b0 6
#962730000000
1!
1%
1-
12
#962740000000
0!
0%
b1 *
0-
02
b1 6
#962750000000
1!
1%
1-
12
#962760000000
0!
0%
b10 *
0-
02
b10 6
#962770000000
1!
1%
1-
12
#962780000000
0!
0%
b11 *
0-
02
b11 6
#962790000000
1!
1%
1-
12
15
#962800000000
0!
0%
b100 *
0-
02
b100 6
#962810000000
1!
1%
1-
12
#962820000000
0!
0%
b101 *
0-
02
b101 6
#962830000000
1!
1%
1-
12
#962840000000
0!
0%
b110 *
0-
02
b110 6
#962850000000
1!
1%
1-
12
#962860000000
0!
0%
b111 *
0-
02
b111 6
#962870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#962880000000
0!
0%
b0 *
0-
02
b0 6
#962890000000
1!
1%
1-
12
#962900000000
0!
0%
b1 *
0-
02
b1 6
#962910000000
1!
1%
1-
12
#962920000000
0!
0%
b10 *
0-
02
b10 6
#962930000000
1!
1%
1-
12
#962940000000
0!
0%
b11 *
0-
02
b11 6
#962950000000
1!
1%
1-
12
15
#962960000000
0!
0%
b100 *
0-
02
b100 6
#962970000000
1!
1%
1-
12
#962980000000
0!
0%
b101 *
0-
02
b101 6
#962990000000
1!
1%
1-
12
#963000000000
0!
0%
b110 *
0-
02
b110 6
#963010000000
1!
1%
1-
12
#963020000000
0!
0%
b111 *
0-
02
b111 6
#963030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#963040000000
0!
0%
b0 *
0-
02
b0 6
#963050000000
1!
1%
1-
12
#963060000000
0!
0%
b1 *
0-
02
b1 6
#963070000000
1!
1%
1-
12
#963080000000
0!
0%
b10 *
0-
02
b10 6
#963090000000
1!
1%
1-
12
#963100000000
0!
0%
b11 *
0-
02
b11 6
#963110000000
1!
1%
1-
12
15
#963120000000
0!
0%
b100 *
0-
02
b100 6
#963130000000
1!
1%
1-
12
#963140000000
0!
0%
b101 *
0-
02
b101 6
#963150000000
1!
1%
1-
12
#963160000000
0!
0%
b110 *
0-
02
b110 6
#963170000000
1!
1%
1-
12
#963180000000
0!
0%
b111 *
0-
02
b111 6
#963190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#963200000000
0!
0%
b0 *
0-
02
b0 6
#963210000000
1!
1%
1-
12
#963220000000
0!
0%
b1 *
0-
02
b1 6
#963230000000
1!
1%
1-
12
#963240000000
0!
0%
b10 *
0-
02
b10 6
#963250000000
1!
1%
1-
12
#963260000000
0!
0%
b11 *
0-
02
b11 6
#963270000000
1!
1%
1-
12
15
#963280000000
0!
0%
b100 *
0-
02
b100 6
#963290000000
1!
1%
1-
12
#963300000000
0!
0%
b101 *
0-
02
b101 6
#963310000000
1!
1%
1-
12
#963320000000
0!
0%
b110 *
0-
02
b110 6
#963330000000
1!
1%
1-
12
#963340000000
0!
0%
b111 *
0-
02
b111 6
#963350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#963360000000
0!
0%
b0 *
0-
02
b0 6
#963370000000
1!
1%
1-
12
#963380000000
0!
0%
b1 *
0-
02
b1 6
#963390000000
1!
1%
1-
12
#963400000000
0!
0%
b10 *
0-
02
b10 6
#963410000000
1!
1%
1-
12
#963420000000
0!
0%
b11 *
0-
02
b11 6
#963430000000
1!
1%
1-
12
15
#963440000000
0!
0%
b100 *
0-
02
b100 6
#963450000000
1!
1%
1-
12
#963460000000
0!
0%
b101 *
0-
02
b101 6
#963470000000
1!
1%
1-
12
#963480000000
0!
0%
b110 *
0-
02
b110 6
#963490000000
1!
1%
1-
12
#963500000000
0!
0%
b111 *
0-
02
b111 6
#963510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#963520000000
0!
0%
b0 *
0-
02
b0 6
#963530000000
1!
1%
1-
12
#963540000000
0!
0%
b1 *
0-
02
b1 6
#963550000000
1!
1%
1-
12
#963560000000
0!
0%
b10 *
0-
02
b10 6
#963570000000
1!
1%
1-
12
#963580000000
0!
0%
b11 *
0-
02
b11 6
#963590000000
1!
1%
1-
12
15
#963600000000
0!
0%
b100 *
0-
02
b100 6
#963610000000
1!
1%
1-
12
#963620000000
0!
0%
b101 *
0-
02
b101 6
#963630000000
1!
1%
1-
12
#963640000000
0!
0%
b110 *
0-
02
b110 6
#963650000000
1!
1%
1-
12
#963660000000
0!
0%
b111 *
0-
02
b111 6
#963670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#963680000000
0!
0%
b0 *
0-
02
b0 6
#963690000000
1!
1%
1-
12
#963700000000
0!
0%
b1 *
0-
02
b1 6
#963710000000
1!
1%
1-
12
#963720000000
0!
0%
b10 *
0-
02
b10 6
#963730000000
1!
1%
1-
12
#963740000000
0!
0%
b11 *
0-
02
b11 6
#963750000000
1!
1%
1-
12
15
#963760000000
0!
0%
b100 *
0-
02
b100 6
#963770000000
1!
1%
1-
12
#963780000000
0!
0%
b101 *
0-
02
b101 6
#963790000000
1!
1%
1-
12
#963800000000
0!
0%
b110 *
0-
02
b110 6
#963810000000
1!
1%
1-
12
#963820000000
0!
0%
b111 *
0-
02
b111 6
#963830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#963840000000
0!
0%
b0 *
0-
02
b0 6
#963850000000
1!
1%
1-
12
#963860000000
0!
0%
b1 *
0-
02
b1 6
#963870000000
1!
1%
1-
12
#963880000000
0!
0%
b10 *
0-
02
b10 6
#963890000000
1!
1%
1-
12
#963900000000
0!
0%
b11 *
0-
02
b11 6
#963910000000
1!
1%
1-
12
15
#963920000000
0!
0%
b100 *
0-
02
b100 6
#963930000000
1!
1%
1-
12
#963940000000
0!
0%
b101 *
0-
02
b101 6
#963950000000
1!
1%
1-
12
#963960000000
0!
0%
b110 *
0-
02
b110 6
#963970000000
1!
1%
1-
12
#963980000000
0!
0%
b111 *
0-
02
b111 6
#963990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#964000000000
0!
0%
b0 *
0-
02
b0 6
#964010000000
1!
1%
1-
12
#964020000000
0!
0%
b1 *
0-
02
b1 6
#964030000000
1!
1%
1-
12
#964040000000
0!
0%
b10 *
0-
02
b10 6
#964050000000
1!
1%
1-
12
#964060000000
0!
0%
b11 *
0-
02
b11 6
#964070000000
1!
1%
1-
12
15
#964080000000
0!
0%
b100 *
0-
02
b100 6
#964090000000
1!
1%
1-
12
#964100000000
0!
0%
b101 *
0-
02
b101 6
#964110000000
1!
1%
1-
12
#964120000000
0!
0%
b110 *
0-
02
b110 6
#964130000000
1!
1%
1-
12
#964140000000
0!
0%
b111 *
0-
02
b111 6
#964150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#964160000000
0!
0%
b0 *
0-
02
b0 6
#964170000000
1!
1%
1-
12
#964180000000
0!
0%
b1 *
0-
02
b1 6
#964190000000
1!
1%
1-
12
#964200000000
0!
0%
b10 *
0-
02
b10 6
#964210000000
1!
1%
1-
12
#964220000000
0!
0%
b11 *
0-
02
b11 6
#964230000000
1!
1%
1-
12
15
#964240000000
0!
0%
b100 *
0-
02
b100 6
#964250000000
1!
1%
1-
12
#964260000000
0!
0%
b101 *
0-
02
b101 6
#964270000000
1!
1%
1-
12
#964280000000
0!
0%
b110 *
0-
02
b110 6
#964290000000
1!
1%
1-
12
#964300000000
0!
0%
b111 *
0-
02
b111 6
#964310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#964320000000
0!
0%
b0 *
0-
02
b0 6
#964330000000
1!
1%
1-
12
#964340000000
0!
0%
b1 *
0-
02
b1 6
#964350000000
1!
1%
1-
12
#964360000000
0!
0%
b10 *
0-
02
b10 6
#964370000000
1!
1%
1-
12
#964380000000
0!
0%
b11 *
0-
02
b11 6
#964390000000
1!
1%
1-
12
15
#964400000000
0!
0%
b100 *
0-
02
b100 6
#964410000000
1!
1%
1-
12
#964420000000
0!
0%
b101 *
0-
02
b101 6
#964430000000
1!
1%
1-
12
#964440000000
0!
0%
b110 *
0-
02
b110 6
#964450000000
1!
1%
1-
12
#964460000000
0!
0%
b111 *
0-
02
b111 6
#964470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#964480000000
0!
0%
b0 *
0-
02
b0 6
#964490000000
1!
1%
1-
12
#964500000000
0!
0%
b1 *
0-
02
b1 6
#964510000000
1!
1%
1-
12
#964520000000
0!
0%
b10 *
0-
02
b10 6
#964530000000
1!
1%
1-
12
#964540000000
0!
0%
b11 *
0-
02
b11 6
#964550000000
1!
1%
1-
12
15
#964560000000
0!
0%
b100 *
0-
02
b100 6
#964570000000
1!
1%
1-
12
#964580000000
0!
0%
b101 *
0-
02
b101 6
#964590000000
1!
1%
1-
12
#964600000000
0!
0%
b110 *
0-
02
b110 6
#964610000000
1!
1%
1-
12
#964620000000
0!
0%
b111 *
0-
02
b111 6
#964630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#964640000000
0!
0%
b0 *
0-
02
b0 6
#964650000000
1!
1%
1-
12
#964660000000
0!
0%
b1 *
0-
02
b1 6
#964670000000
1!
1%
1-
12
#964680000000
0!
0%
b10 *
0-
02
b10 6
#964690000000
1!
1%
1-
12
#964700000000
0!
0%
b11 *
0-
02
b11 6
#964710000000
1!
1%
1-
12
15
#964720000000
0!
0%
b100 *
0-
02
b100 6
#964730000000
1!
1%
1-
12
#964740000000
0!
0%
b101 *
0-
02
b101 6
#964750000000
1!
1%
1-
12
#964760000000
0!
0%
b110 *
0-
02
b110 6
#964770000000
1!
1%
1-
12
#964780000000
0!
0%
b111 *
0-
02
b111 6
#964790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#964800000000
0!
0%
b0 *
0-
02
b0 6
#964810000000
1!
1%
1-
12
#964820000000
0!
0%
b1 *
0-
02
b1 6
#964830000000
1!
1%
1-
12
#964840000000
0!
0%
b10 *
0-
02
b10 6
#964850000000
1!
1%
1-
12
#964860000000
0!
0%
b11 *
0-
02
b11 6
#964870000000
1!
1%
1-
12
15
#964880000000
0!
0%
b100 *
0-
02
b100 6
#964890000000
1!
1%
1-
12
#964900000000
0!
0%
b101 *
0-
02
b101 6
#964910000000
1!
1%
1-
12
#964920000000
0!
0%
b110 *
0-
02
b110 6
#964930000000
1!
1%
1-
12
#964940000000
0!
0%
b111 *
0-
02
b111 6
#964950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#964960000000
0!
0%
b0 *
0-
02
b0 6
#964970000000
1!
1%
1-
12
#964980000000
0!
0%
b1 *
0-
02
b1 6
#964990000000
1!
1%
1-
12
#965000000000
0!
0%
b10 *
0-
02
b10 6
#965010000000
1!
1%
1-
12
#965020000000
0!
0%
b11 *
0-
02
b11 6
#965030000000
1!
1%
1-
12
15
#965040000000
0!
0%
b100 *
0-
02
b100 6
#965050000000
1!
1%
1-
12
#965060000000
0!
0%
b101 *
0-
02
b101 6
#965070000000
1!
1%
1-
12
#965080000000
0!
0%
b110 *
0-
02
b110 6
#965090000000
1!
1%
1-
12
#965100000000
0!
0%
b111 *
0-
02
b111 6
#965110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#965120000000
0!
0%
b0 *
0-
02
b0 6
#965130000000
1!
1%
1-
12
#965140000000
0!
0%
b1 *
0-
02
b1 6
#965150000000
1!
1%
1-
12
#965160000000
0!
0%
b10 *
0-
02
b10 6
#965170000000
1!
1%
1-
12
#965180000000
0!
0%
b11 *
0-
02
b11 6
#965190000000
1!
1%
1-
12
15
#965200000000
0!
0%
b100 *
0-
02
b100 6
#965210000000
1!
1%
1-
12
#965220000000
0!
0%
b101 *
0-
02
b101 6
#965230000000
1!
1%
1-
12
#965240000000
0!
0%
b110 *
0-
02
b110 6
#965250000000
1!
1%
1-
12
#965260000000
0!
0%
b111 *
0-
02
b111 6
#965270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#965280000000
0!
0%
b0 *
0-
02
b0 6
#965290000000
1!
1%
1-
12
#965300000000
0!
0%
b1 *
0-
02
b1 6
#965310000000
1!
1%
1-
12
#965320000000
0!
0%
b10 *
0-
02
b10 6
#965330000000
1!
1%
1-
12
#965340000000
0!
0%
b11 *
0-
02
b11 6
#965350000000
1!
1%
1-
12
15
#965360000000
0!
0%
b100 *
0-
02
b100 6
#965370000000
1!
1%
1-
12
#965380000000
0!
0%
b101 *
0-
02
b101 6
#965390000000
1!
1%
1-
12
#965400000000
0!
0%
b110 *
0-
02
b110 6
#965410000000
1!
1%
1-
12
#965420000000
0!
0%
b111 *
0-
02
b111 6
#965430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#965440000000
0!
0%
b0 *
0-
02
b0 6
#965450000000
1!
1%
1-
12
#965460000000
0!
0%
b1 *
0-
02
b1 6
#965470000000
1!
1%
1-
12
#965480000000
0!
0%
b10 *
0-
02
b10 6
#965490000000
1!
1%
1-
12
#965500000000
0!
0%
b11 *
0-
02
b11 6
#965510000000
1!
1%
1-
12
15
#965520000000
0!
0%
b100 *
0-
02
b100 6
#965530000000
1!
1%
1-
12
#965540000000
0!
0%
b101 *
0-
02
b101 6
#965550000000
1!
1%
1-
12
#965560000000
0!
0%
b110 *
0-
02
b110 6
#965570000000
1!
1%
1-
12
#965580000000
0!
0%
b111 *
0-
02
b111 6
#965590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#965600000000
0!
0%
b0 *
0-
02
b0 6
#965610000000
1!
1%
1-
12
#965620000000
0!
0%
b1 *
0-
02
b1 6
#965630000000
1!
1%
1-
12
#965640000000
0!
0%
b10 *
0-
02
b10 6
#965650000000
1!
1%
1-
12
#965660000000
0!
0%
b11 *
0-
02
b11 6
#965670000000
1!
1%
1-
12
15
#965680000000
0!
0%
b100 *
0-
02
b100 6
#965690000000
1!
1%
1-
12
#965700000000
0!
0%
b101 *
0-
02
b101 6
#965710000000
1!
1%
1-
12
#965720000000
0!
0%
b110 *
0-
02
b110 6
#965730000000
1!
1%
1-
12
#965740000000
0!
0%
b111 *
0-
02
b111 6
#965750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#965760000000
0!
0%
b0 *
0-
02
b0 6
#965770000000
1!
1%
1-
12
#965780000000
0!
0%
b1 *
0-
02
b1 6
#965790000000
1!
1%
1-
12
#965800000000
0!
0%
b10 *
0-
02
b10 6
#965810000000
1!
1%
1-
12
#965820000000
0!
0%
b11 *
0-
02
b11 6
#965830000000
1!
1%
1-
12
15
#965840000000
0!
0%
b100 *
0-
02
b100 6
#965850000000
1!
1%
1-
12
#965860000000
0!
0%
b101 *
0-
02
b101 6
#965870000000
1!
1%
1-
12
#965880000000
0!
0%
b110 *
0-
02
b110 6
#965890000000
1!
1%
1-
12
#965900000000
0!
0%
b111 *
0-
02
b111 6
#965910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#965920000000
0!
0%
b0 *
0-
02
b0 6
#965930000000
1!
1%
1-
12
#965940000000
0!
0%
b1 *
0-
02
b1 6
#965950000000
1!
1%
1-
12
#965960000000
0!
0%
b10 *
0-
02
b10 6
#965970000000
1!
1%
1-
12
#965980000000
0!
0%
b11 *
0-
02
b11 6
#965990000000
1!
1%
1-
12
15
#966000000000
0!
0%
b100 *
0-
02
b100 6
#966010000000
1!
1%
1-
12
#966020000000
0!
0%
b101 *
0-
02
b101 6
#966030000000
1!
1%
1-
12
#966040000000
0!
0%
b110 *
0-
02
b110 6
#966050000000
1!
1%
1-
12
#966060000000
0!
0%
b111 *
0-
02
b111 6
#966070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#966080000000
0!
0%
b0 *
0-
02
b0 6
#966090000000
1!
1%
1-
12
#966100000000
0!
0%
b1 *
0-
02
b1 6
#966110000000
1!
1%
1-
12
#966120000000
0!
0%
b10 *
0-
02
b10 6
#966130000000
1!
1%
1-
12
#966140000000
0!
0%
b11 *
0-
02
b11 6
#966150000000
1!
1%
1-
12
15
#966160000000
0!
0%
b100 *
0-
02
b100 6
#966170000000
1!
1%
1-
12
#966180000000
0!
0%
b101 *
0-
02
b101 6
#966190000000
1!
1%
1-
12
#966200000000
0!
0%
b110 *
0-
02
b110 6
#966210000000
1!
1%
1-
12
#966220000000
0!
0%
b111 *
0-
02
b111 6
#966230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#966240000000
0!
0%
b0 *
0-
02
b0 6
#966250000000
1!
1%
1-
12
#966260000000
0!
0%
b1 *
0-
02
b1 6
#966270000000
1!
1%
1-
12
#966280000000
0!
0%
b10 *
0-
02
b10 6
#966290000000
1!
1%
1-
12
#966300000000
0!
0%
b11 *
0-
02
b11 6
#966310000000
1!
1%
1-
12
15
#966320000000
0!
0%
b100 *
0-
02
b100 6
#966330000000
1!
1%
1-
12
#966340000000
0!
0%
b101 *
0-
02
b101 6
#966350000000
1!
1%
1-
12
#966360000000
0!
0%
b110 *
0-
02
b110 6
#966370000000
1!
1%
1-
12
#966380000000
0!
0%
b111 *
0-
02
b111 6
#966390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#966400000000
0!
0%
b0 *
0-
02
b0 6
#966410000000
1!
1%
1-
12
#966420000000
0!
0%
b1 *
0-
02
b1 6
#966430000000
1!
1%
1-
12
#966440000000
0!
0%
b10 *
0-
02
b10 6
#966450000000
1!
1%
1-
12
#966460000000
0!
0%
b11 *
0-
02
b11 6
#966470000000
1!
1%
1-
12
15
#966480000000
0!
0%
b100 *
0-
02
b100 6
#966490000000
1!
1%
1-
12
#966500000000
0!
0%
b101 *
0-
02
b101 6
#966510000000
1!
1%
1-
12
#966520000000
0!
0%
b110 *
0-
02
b110 6
#966530000000
1!
1%
1-
12
#966540000000
0!
0%
b111 *
0-
02
b111 6
#966550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#966560000000
0!
0%
b0 *
0-
02
b0 6
#966570000000
1!
1%
1-
12
#966580000000
0!
0%
b1 *
0-
02
b1 6
#966590000000
1!
1%
1-
12
#966600000000
0!
0%
b10 *
0-
02
b10 6
#966610000000
1!
1%
1-
12
#966620000000
0!
0%
b11 *
0-
02
b11 6
#966630000000
1!
1%
1-
12
15
#966640000000
0!
0%
b100 *
0-
02
b100 6
#966650000000
1!
1%
1-
12
#966660000000
0!
0%
b101 *
0-
02
b101 6
#966670000000
1!
1%
1-
12
#966680000000
0!
0%
b110 *
0-
02
b110 6
#966690000000
1!
1%
1-
12
#966700000000
0!
0%
b111 *
0-
02
b111 6
#966710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#966720000000
0!
0%
b0 *
0-
02
b0 6
#966730000000
1!
1%
1-
12
#966740000000
0!
0%
b1 *
0-
02
b1 6
#966750000000
1!
1%
1-
12
#966760000000
0!
0%
b10 *
0-
02
b10 6
#966770000000
1!
1%
1-
12
#966780000000
0!
0%
b11 *
0-
02
b11 6
#966790000000
1!
1%
1-
12
15
#966800000000
0!
0%
b100 *
0-
02
b100 6
#966810000000
1!
1%
1-
12
#966820000000
0!
0%
b101 *
0-
02
b101 6
#966830000000
1!
1%
1-
12
#966840000000
0!
0%
b110 *
0-
02
b110 6
#966850000000
1!
1%
1-
12
#966860000000
0!
0%
b111 *
0-
02
b111 6
#966870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#966880000000
0!
0%
b0 *
0-
02
b0 6
#966890000000
1!
1%
1-
12
#966900000000
0!
0%
b1 *
0-
02
b1 6
#966910000000
1!
1%
1-
12
#966920000000
0!
0%
b10 *
0-
02
b10 6
#966930000000
1!
1%
1-
12
#966940000000
0!
0%
b11 *
0-
02
b11 6
#966950000000
1!
1%
1-
12
15
#966960000000
0!
0%
b100 *
0-
02
b100 6
#966970000000
1!
1%
1-
12
#966980000000
0!
0%
b101 *
0-
02
b101 6
#966990000000
1!
1%
1-
12
#967000000000
0!
0%
b110 *
0-
02
b110 6
#967010000000
1!
1%
1-
12
#967020000000
0!
0%
b111 *
0-
02
b111 6
#967030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#967040000000
0!
0%
b0 *
0-
02
b0 6
#967050000000
1!
1%
1-
12
#967060000000
0!
0%
b1 *
0-
02
b1 6
#967070000000
1!
1%
1-
12
#967080000000
0!
0%
b10 *
0-
02
b10 6
#967090000000
1!
1%
1-
12
#967100000000
0!
0%
b11 *
0-
02
b11 6
#967110000000
1!
1%
1-
12
15
#967120000000
0!
0%
b100 *
0-
02
b100 6
#967130000000
1!
1%
1-
12
#967140000000
0!
0%
b101 *
0-
02
b101 6
#967150000000
1!
1%
1-
12
#967160000000
0!
0%
b110 *
0-
02
b110 6
#967170000000
1!
1%
1-
12
#967180000000
0!
0%
b111 *
0-
02
b111 6
#967190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#967200000000
0!
0%
b0 *
0-
02
b0 6
#967210000000
1!
1%
1-
12
#967220000000
0!
0%
b1 *
0-
02
b1 6
#967230000000
1!
1%
1-
12
#967240000000
0!
0%
b10 *
0-
02
b10 6
#967250000000
1!
1%
1-
12
#967260000000
0!
0%
b11 *
0-
02
b11 6
#967270000000
1!
1%
1-
12
15
#967280000000
0!
0%
b100 *
0-
02
b100 6
#967290000000
1!
1%
1-
12
#967300000000
0!
0%
b101 *
0-
02
b101 6
#967310000000
1!
1%
1-
12
#967320000000
0!
0%
b110 *
0-
02
b110 6
#967330000000
1!
1%
1-
12
#967340000000
0!
0%
b111 *
0-
02
b111 6
#967350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#967360000000
0!
0%
b0 *
0-
02
b0 6
#967370000000
1!
1%
1-
12
#967380000000
0!
0%
b1 *
0-
02
b1 6
#967390000000
1!
1%
1-
12
#967400000000
0!
0%
b10 *
0-
02
b10 6
#967410000000
1!
1%
1-
12
#967420000000
0!
0%
b11 *
0-
02
b11 6
#967430000000
1!
1%
1-
12
15
#967440000000
0!
0%
b100 *
0-
02
b100 6
#967450000000
1!
1%
1-
12
#967460000000
0!
0%
b101 *
0-
02
b101 6
#967470000000
1!
1%
1-
12
#967480000000
0!
0%
b110 *
0-
02
b110 6
#967490000000
1!
1%
1-
12
#967500000000
0!
0%
b111 *
0-
02
b111 6
#967510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#967520000000
0!
0%
b0 *
0-
02
b0 6
#967530000000
1!
1%
1-
12
#967540000000
0!
0%
b1 *
0-
02
b1 6
#967550000000
1!
1%
1-
12
#967560000000
0!
0%
b10 *
0-
02
b10 6
#967570000000
1!
1%
1-
12
#967580000000
0!
0%
b11 *
0-
02
b11 6
#967590000000
1!
1%
1-
12
15
#967600000000
0!
0%
b100 *
0-
02
b100 6
#967610000000
1!
1%
1-
12
#967620000000
0!
0%
b101 *
0-
02
b101 6
#967630000000
1!
1%
1-
12
#967640000000
0!
0%
b110 *
0-
02
b110 6
#967650000000
1!
1%
1-
12
#967660000000
0!
0%
b111 *
0-
02
b111 6
#967670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#967680000000
0!
0%
b0 *
0-
02
b0 6
#967690000000
1!
1%
1-
12
#967700000000
0!
0%
b1 *
0-
02
b1 6
#967710000000
1!
1%
1-
12
#967720000000
0!
0%
b10 *
0-
02
b10 6
#967730000000
1!
1%
1-
12
#967740000000
0!
0%
b11 *
0-
02
b11 6
#967750000000
1!
1%
1-
12
15
#967760000000
0!
0%
b100 *
0-
02
b100 6
#967770000000
1!
1%
1-
12
#967780000000
0!
0%
b101 *
0-
02
b101 6
#967790000000
1!
1%
1-
12
#967800000000
0!
0%
b110 *
0-
02
b110 6
#967810000000
1!
1%
1-
12
#967820000000
0!
0%
b111 *
0-
02
b111 6
#967830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#967840000000
0!
0%
b0 *
0-
02
b0 6
#967850000000
1!
1%
1-
12
#967860000000
0!
0%
b1 *
0-
02
b1 6
#967870000000
1!
1%
1-
12
#967880000000
0!
0%
b10 *
0-
02
b10 6
#967890000000
1!
1%
1-
12
#967900000000
0!
0%
b11 *
0-
02
b11 6
#967910000000
1!
1%
1-
12
15
#967920000000
0!
0%
b100 *
0-
02
b100 6
#967930000000
1!
1%
1-
12
#967940000000
0!
0%
b101 *
0-
02
b101 6
#967950000000
1!
1%
1-
12
#967960000000
0!
0%
b110 *
0-
02
b110 6
#967970000000
1!
1%
1-
12
#967980000000
0!
0%
b111 *
0-
02
b111 6
#967990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#968000000000
0!
0%
b0 *
0-
02
b0 6
#968010000000
1!
1%
1-
12
#968020000000
0!
0%
b1 *
0-
02
b1 6
#968030000000
1!
1%
1-
12
#968040000000
0!
0%
b10 *
0-
02
b10 6
#968050000000
1!
1%
1-
12
#968060000000
0!
0%
b11 *
0-
02
b11 6
#968070000000
1!
1%
1-
12
15
#968080000000
0!
0%
b100 *
0-
02
b100 6
#968090000000
1!
1%
1-
12
#968100000000
0!
0%
b101 *
0-
02
b101 6
#968110000000
1!
1%
1-
12
#968120000000
0!
0%
b110 *
0-
02
b110 6
#968130000000
1!
1%
1-
12
#968140000000
0!
0%
b111 *
0-
02
b111 6
#968150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#968160000000
0!
0%
b0 *
0-
02
b0 6
#968170000000
1!
1%
1-
12
#968180000000
0!
0%
b1 *
0-
02
b1 6
#968190000000
1!
1%
1-
12
#968200000000
0!
0%
b10 *
0-
02
b10 6
#968210000000
1!
1%
1-
12
#968220000000
0!
0%
b11 *
0-
02
b11 6
#968230000000
1!
1%
1-
12
15
#968240000000
0!
0%
b100 *
0-
02
b100 6
#968250000000
1!
1%
1-
12
#968260000000
0!
0%
b101 *
0-
02
b101 6
#968270000000
1!
1%
1-
12
#968280000000
0!
0%
b110 *
0-
02
b110 6
#968290000000
1!
1%
1-
12
#968300000000
0!
0%
b111 *
0-
02
b111 6
#968310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#968320000000
0!
0%
b0 *
0-
02
b0 6
#968330000000
1!
1%
1-
12
#968340000000
0!
0%
b1 *
0-
02
b1 6
#968350000000
1!
1%
1-
12
#968360000000
0!
0%
b10 *
0-
02
b10 6
#968370000000
1!
1%
1-
12
#968380000000
0!
0%
b11 *
0-
02
b11 6
#968390000000
1!
1%
1-
12
15
#968400000000
0!
0%
b100 *
0-
02
b100 6
#968410000000
1!
1%
1-
12
#968420000000
0!
0%
b101 *
0-
02
b101 6
#968430000000
1!
1%
1-
12
#968440000000
0!
0%
b110 *
0-
02
b110 6
#968450000000
1!
1%
1-
12
#968460000000
0!
0%
b111 *
0-
02
b111 6
#968470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#968480000000
0!
0%
b0 *
0-
02
b0 6
#968490000000
1!
1%
1-
12
#968500000000
0!
0%
b1 *
0-
02
b1 6
#968510000000
1!
1%
1-
12
#968520000000
0!
0%
b10 *
0-
02
b10 6
#968530000000
1!
1%
1-
12
#968540000000
0!
0%
b11 *
0-
02
b11 6
#968550000000
1!
1%
1-
12
15
#968560000000
0!
0%
b100 *
0-
02
b100 6
#968570000000
1!
1%
1-
12
#968580000000
0!
0%
b101 *
0-
02
b101 6
#968590000000
1!
1%
1-
12
#968600000000
0!
0%
b110 *
0-
02
b110 6
#968610000000
1!
1%
1-
12
#968620000000
0!
0%
b111 *
0-
02
b111 6
#968630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#968640000000
0!
0%
b0 *
0-
02
b0 6
#968650000000
1!
1%
1-
12
#968660000000
0!
0%
b1 *
0-
02
b1 6
#968670000000
1!
1%
1-
12
#968680000000
0!
0%
b10 *
0-
02
b10 6
#968690000000
1!
1%
1-
12
#968700000000
0!
0%
b11 *
0-
02
b11 6
#968710000000
1!
1%
1-
12
15
#968720000000
0!
0%
b100 *
0-
02
b100 6
#968730000000
1!
1%
1-
12
#968740000000
0!
0%
b101 *
0-
02
b101 6
#968750000000
1!
1%
1-
12
#968760000000
0!
0%
b110 *
0-
02
b110 6
#968770000000
1!
1%
1-
12
#968780000000
0!
0%
b111 *
0-
02
b111 6
#968790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#968800000000
0!
0%
b0 *
0-
02
b0 6
#968810000000
1!
1%
1-
12
#968820000000
0!
0%
b1 *
0-
02
b1 6
#968830000000
1!
1%
1-
12
#968840000000
0!
0%
b10 *
0-
02
b10 6
#968850000000
1!
1%
1-
12
#968860000000
0!
0%
b11 *
0-
02
b11 6
#968870000000
1!
1%
1-
12
15
#968880000000
0!
0%
b100 *
0-
02
b100 6
#968890000000
1!
1%
1-
12
#968900000000
0!
0%
b101 *
0-
02
b101 6
#968910000000
1!
1%
1-
12
#968920000000
0!
0%
b110 *
0-
02
b110 6
#968930000000
1!
1%
1-
12
#968940000000
0!
0%
b111 *
0-
02
b111 6
#968950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#968960000000
0!
0%
b0 *
0-
02
b0 6
#968970000000
1!
1%
1-
12
#968980000000
0!
0%
b1 *
0-
02
b1 6
#968990000000
1!
1%
1-
12
#969000000000
0!
0%
b10 *
0-
02
b10 6
#969010000000
1!
1%
1-
12
#969020000000
0!
0%
b11 *
0-
02
b11 6
#969030000000
1!
1%
1-
12
15
#969040000000
0!
0%
b100 *
0-
02
b100 6
#969050000000
1!
1%
1-
12
#969060000000
0!
0%
b101 *
0-
02
b101 6
#969070000000
1!
1%
1-
12
#969080000000
0!
0%
b110 *
0-
02
b110 6
#969090000000
1!
1%
1-
12
#969100000000
0!
0%
b111 *
0-
02
b111 6
#969110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#969120000000
0!
0%
b0 *
0-
02
b0 6
#969130000000
1!
1%
1-
12
#969140000000
0!
0%
b1 *
0-
02
b1 6
#969150000000
1!
1%
1-
12
#969160000000
0!
0%
b10 *
0-
02
b10 6
#969170000000
1!
1%
1-
12
#969180000000
0!
0%
b11 *
0-
02
b11 6
#969190000000
1!
1%
1-
12
15
#969200000000
0!
0%
b100 *
0-
02
b100 6
#969210000000
1!
1%
1-
12
#969220000000
0!
0%
b101 *
0-
02
b101 6
#969230000000
1!
1%
1-
12
#969240000000
0!
0%
b110 *
0-
02
b110 6
#969250000000
1!
1%
1-
12
#969260000000
0!
0%
b111 *
0-
02
b111 6
#969270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#969280000000
0!
0%
b0 *
0-
02
b0 6
#969290000000
1!
1%
1-
12
#969300000000
0!
0%
b1 *
0-
02
b1 6
#969310000000
1!
1%
1-
12
#969320000000
0!
0%
b10 *
0-
02
b10 6
#969330000000
1!
1%
1-
12
#969340000000
0!
0%
b11 *
0-
02
b11 6
#969350000000
1!
1%
1-
12
15
#969360000000
0!
0%
b100 *
0-
02
b100 6
#969370000000
1!
1%
1-
12
#969380000000
0!
0%
b101 *
0-
02
b101 6
#969390000000
1!
1%
1-
12
#969400000000
0!
0%
b110 *
0-
02
b110 6
#969410000000
1!
1%
1-
12
#969420000000
0!
0%
b111 *
0-
02
b111 6
#969430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#969440000000
0!
0%
b0 *
0-
02
b0 6
#969450000000
1!
1%
1-
12
#969460000000
0!
0%
b1 *
0-
02
b1 6
#969470000000
1!
1%
1-
12
#969480000000
0!
0%
b10 *
0-
02
b10 6
#969490000000
1!
1%
1-
12
#969500000000
0!
0%
b11 *
0-
02
b11 6
#969510000000
1!
1%
1-
12
15
#969520000000
0!
0%
b100 *
0-
02
b100 6
#969530000000
1!
1%
1-
12
#969540000000
0!
0%
b101 *
0-
02
b101 6
#969550000000
1!
1%
1-
12
#969560000000
0!
0%
b110 *
0-
02
b110 6
#969570000000
1!
1%
1-
12
#969580000000
0!
0%
b111 *
0-
02
b111 6
#969590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#969600000000
0!
0%
b0 *
0-
02
b0 6
#969610000000
1!
1%
1-
12
#969620000000
0!
0%
b1 *
0-
02
b1 6
#969630000000
1!
1%
1-
12
#969640000000
0!
0%
b10 *
0-
02
b10 6
#969650000000
1!
1%
1-
12
#969660000000
0!
0%
b11 *
0-
02
b11 6
#969670000000
1!
1%
1-
12
15
#969680000000
0!
0%
b100 *
0-
02
b100 6
#969690000000
1!
1%
1-
12
#969700000000
0!
0%
b101 *
0-
02
b101 6
#969710000000
1!
1%
1-
12
#969720000000
0!
0%
b110 *
0-
02
b110 6
#969730000000
1!
1%
1-
12
#969740000000
0!
0%
b111 *
0-
02
b111 6
#969750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#969760000000
0!
0%
b0 *
0-
02
b0 6
#969770000000
1!
1%
1-
12
#969780000000
0!
0%
b1 *
0-
02
b1 6
#969790000000
1!
1%
1-
12
#969800000000
0!
0%
b10 *
0-
02
b10 6
#969810000000
1!
1%
1-
12
#969820000000
0!
0%
b11 *
0-
02
b11 6
#969830000000
1!
1%
1-
12
15
#969840000000
0!
0%
b100 *
0-
02
b100 6
#969850000000
1!
1%
1-
12
#969860000000
0!
0%
b101 *
0-
02
b101 6
#969870000000
1!
1%
1-
12
#969880000000
0!
0%
b110 *
0-
02
b110 6
#969890000000
1!
1%
1-
12
#969900000000
0!
0%
b111 *
0-
02
b111 6
#969910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#969920000000
0!
0%
b0 *
0-
02
b0 6
#969930000000
1!
1%
1-
12
#969940000000
0!
0%
b1 *
0-
02
b1 6
#969950000000
1!
1%
1-
12
#969960000000
0!
0%
b10 *
0-
02
b10 6
#969970000000
1!
1%
1-
12
#969980000000
0!
0%
b11 *
0-
02
b11 6
#969990000000
1!
1%
1-
12
15
#970000000000
0!
0%
b100 *
0-
02
b100 6
#970010000000
1!
1%
1-
12
#970020000000
0!
0%
b101 *
0-
02
b101 6
#970030000000
1!
1%
1-
12
#970040000000
0!
0%
b110 *
0-
02
b110 6
#970050000000
1!
1%
1-
12
#970060000000
0!
0%
b111 *
0-
02
b111 6
#970070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#970080000000
0!
0%
b0 *
0-
02
b0 6
#970090000000
1!
1%
1-
12
#970100000000
0!
0%
b1 *
0-
02
b1 6
#970110000000
1!
1%
1-
12
#970120000000
0!
0%
b10 *
0-
02
b10 6
#970130000000
1!
1%
1-
12
#970140000000
0!
0%
b11 *
0-
02
b11 6
#970150000000
1!
1%
1-
12
15
#970160000000
0!
0%
b100 *
0-
02
b100 6
#970170000000
1!
1%
1-
12
#970180000000
0!
0%
b101 *
0-
02
b101 6
#970190000000
1!
1%
1-
12
#970200000000
0!
0%
b110 *
0-
02
b110 6
#970210000000
1!
1%
1-
12
#970220000000
0!
0%
b111 *
0-
02
b111 6
#970230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#970240000000
0!
0%
b0 *
0-
02
b0 6
#970250000000
1!
1%
1-
12
#970260000000
0!
0%
b1 *
0-
02
b1 6
#970270000000
1!
1%
1-
12
#970280000000
0!
0%
b10 *
0-
02
b10 6
#970290000000
1!
1%
1-
12
#970300000000
0!
0%
b11 *
0-
02
b11 6
#970310000000
1!
1%
1-
12
15
#970320000000
0!
0%
b100 *
0-
02
b100 6
#970330000000
1!
1%
1-
12
#970340000000
0!
0%
b101 *
0-
02
b101 6
#970350000000
1!
1%
1-
12
#970360000000
0!
0%
b110 *
0-
02
b110 6
#970370000000
1!
1%
1-
12
#970380000000
0!
0%
b111 *
0-
02
b111 6
#970390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#970400000000
0!
0%
b0 *
0-
02
b0 6
#970410000000
1!
1%
1-
12
#970420000000
0!
0%
b1 *
0-
02
b1 6
#970430000000
1!
1%
1-
12
#970440000000
0!
0%
b10 *
0-
02
b10 6
#970450000000
1!
1%
1-
12
#970460000000
0!
0%
b11 *
0-
02
b11 6
#970470000000
1!
1%
1-
12
15
#970480000000
0!
0%
b100 *
0-
02
b100 6
#970490000000
1!
1%
1-
12
#970500000000
0!
0%
b101 *
0-
02
b101 6
#970510000000
1!
1%
1-
12
#970520000000
0!
0%
b110 *
0-
02
b110 6
#970530000000
1!
1%
1-
12
#970540000000
0!
0%
b111 *
0-
02
b111 6
#970550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#970560000000
0!
0%
b0 *
0-
02
b0 6
#970570000000
1!
1%
1-
12
#970580000000
0!
0%
b1 *
0-
02
b1 6
#970590000000
1!
1%
1-
12
#970600000000
0!
0%
b10 *
0-
02
b10 6
#970610000000
1!
1%
1-
12
#970620000000
0!
0%
b11 *
0-
02
b11 6
#970630000000
1!
1%
1-
12
15
#970640000000
0!
0%
b100 *
0-
02
b100 6
#970650000000
1!
1%
1-
12
#970660000000
0!
0%
b101 *
0-
02
b101 6
#970670000000
1!
1%
1-
12
#970680000000
0!
0%
b110 *
0-
02
b110 6
#970690000000
1!
1%
1-
12
#970700000000
0!
0%
b111 *
0-
02
b111 6
#970710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#970720000000
0!
0%
b0 *
0-
02
b0 6
#970730000000
1!
1%
1-
12
#970740000000
0!
0%
b1 *
0-
02
b1 6
#970750000000
1!
1%
1-
12
#970760000000
0!
0%
b10 *
0-
02
b10 6
#970770000000
1!
1%
1-
12
#970780000000
0!
0%
b11 *
0-
02
b11 6
#970790000000
1!
1%
1-
12
15
#970800000000
0!
0%
b100 *
0-
02
b100 6
#970810000000
1!
1%
1-
12
#970820000000
0!
0%
b101 *
0-
02
b101 6
#970830000000
1!
1%
1-
12
#970840000000
0!
0%
b110 *
0-
02
b110 6
#970850000000
1!
1%
1-
12
#970860000000
0!
0%
b111 *
0-
02
b111 6
#970870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#970880000000
0!
0%
b0 *
0-
02
b0 6
#970890000000
1!
1%
1-
12
#970900000000
0!
0%
b1 *
0-
02
b1 6
#970910000000
1!
1%
1-
12
#970920000000
0!
0%
b10 *
0-
02
b10 6
#970930000000
1!
1%
1-
12
#970940000000
0!
0%
b11 *
0-
02
b11 6
#970950000000
1!
1%
1-
12
15
#970960000000
0!
0%
b100 *
0-
02
b100 6
#970970000000
1!
1%
1-
12
#970980000000
0!
0%
b101 *
0-
02
b101 6
#970990000000
1!
1%
1-
12
#971000000000
0!
0%
b110 *
0-
02
b110 6
#971010000000
1!
1%
1-
12
#971020000000
0!
0%
b111 *
0-
02
b111 6
#971030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#971040000000
0!
0%
b0 *
0-
02
b0 6
#971050000000
1!
1%
1-
12
#971060000000
0!
0%
b1 *
0-
02
b1 6
#971070000000
1!
1%
1-
12
#971080000000
0!
0%
b10 *
0-
02
b10 6
#971090000000
1!
1%
1-
12
#971100000000
0!
0%
b11 *
0-
02
b11 6
#971110000000
1!
1%
1-
12
15
#971120000000
0!
0%
b100 *
0-
02
b100 6
#971130000000
1!
1%
1-
12
#971140000000
0!
0%
b101 *
0-
02
b101 6
#971150000000
1!
1%
1-
12
#971160000000
0!
0%
b110 *
0-
02
b110 6
#971170000000
1!
1%
1-
12
#971180000000
0!
0%
b111 *
0-
02
b111 6
#971190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#971200000000
0!
0%
b0 *
0-
02
b0 6
#971210000000
1!
1%
1-
12
#971220000000
0!
0%
b1 *
0-
02
b1 6
#971230000000
1!
1%
1-
12
#971240000000
0!
0%
b10 *
0-
02
b10 6
#971250000000
1!
1%
1-
12
#971260000000
0!
0%
b11 *
0-
02
b11 6
#971270000000
1!
1%
1-
12
15
#971280000000
0!
0%
b100 *
0-
02
b100 6
#971290000000
1!
1%
1-
12
#971300000000
0!
0%
b101 *
0-
02
b101 6
#971310000000
1!
1%
1-
12
#971320000000
0!
0%
b110 *
0-
02
b110 6
#971330000000
1!
1%
1-
12
#971340000000
0!
0%
b111 *
0-
02
b111 6
#971350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#971360000000
0!
0%
b0 *
0-
02
b0 6
#971370000000
1!
1%
1-
12
#971380000000
0!
0%
b1 *
0-
02
b1 6
#971390000000
1!
1%
1-
12
#971400000000
0!
0%
b10 *
0-
02
b10 6
#971410000000
1!
1%
1-
12
#971420000000
0!
0%
b11 *
0-
02
b11 6
#971430000000
1!
1%
1-
12
15
#971440000000
0!
0%
b100 *
0-
02
b100 6
#971450000000
1!
1%
1-
12
#971460000000
0!
0%
b101 *
0-
02
b101 6
#971470000000
1!
1%
1-
12
#971480000000
0!
0%
b110 *
0-
02
b110 6
#971490000000
1!
1%
1-
12
#971500000000
0!
0%
b111 *
0-
02
b111 6
#971510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#971520000000
0!
0%
b0 *
0-
02
b0 6
#971530000000
1!
1%
1-
12
#971540000000
0!
0%
b1 *
0-
02
b1 6
#971550000000
1!
1%
1-
12
#971560000000
0!
0%
b10 *
0-
02
b10 6
#971570000000
1!
1%
1-
12
#971580000000
0!
0%
b11 *
0-
02
b11 6
#971590000000
1!
1%
1-
12
15
#971600000000
0!
0%
b100 *
0-
02
b100 6
#971610000000
1!
1%
1-
12
#971620000000
0!
0%
b101 *
0-
02
b101 6
#971630000000
1!
1%
1-
12
#971640000000
0!
0%
b110 *
0-
02
b110 6
#971650000000
1!
1%
1-
12
#971660000000
0!
0%
b111 *
0-
02
b111 6
#971670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#971680000000
0!
0%
b0 *
0-
02
b0 6
#971690000000
1!
1%
1-
12
#971700000000
0!
0%
b1 *
0-
02
b1 6
#971710000000
1!
1%
1-
12
#971720000000
0!
0%
b10 *
0-
02
b10 6
#971730000000
1!
1%
1-
12
#971740000000
0!
0%
b11 *
0-
02
b11 6
#971750000000
1!
1%
1-
12
15
#971760000000
0!
0%
b100 *
0-
02
b100 6
#971770000000
1!
1%
1-
12
#971780000000
0!
0%
b101 *
0-
02
b101 6
#971790000000
1!
1%
1-
12
#971800000000
0!
0%
b110 *
0-
02
b110 6
#971810000000
1!
1%
1-
12
#971820000000
0!
0%
b111 *
0-
02
b111 6
#971830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#971840000000
0!
0%
b0 *
0-
02
b0 6
#971850000000
1!
1%
1-
12
#971860000000
0!
0%
b1 *
0-
02
b1 6
#971870000000
1!
1%
1-
12
#971880000000
0!
0%
b10 *
0-
02
b10 6
#971890000000
1!
1%
1-
12
#971900000000
0!
0%
b11 *
0-
02
b11 6
#971910000000
1!
1%
1-
12
15
#971920000000
0!
0%
b100 *
0-
02
b100 6
#971930000000
1!
1%
1-
12
#971940000000
0!
0%
b101 *
0-
02
b101 6
#971950000000
1!
1%
1-
12
#971960000000
0!
0%
b110 *
0-
02
b110 6
#971970000000
1!
1%
1-
12
#971980000000
0!
0%
b111 *
0-
02
b111 6
#971990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#972000000000
0!
0%
b0 *
0-
02
b0 6
#972010000000
1!
1%
1-
12
#972020000000
0!
0%
b1 *
0-
02
b1 6
#972030000000
1!
1%
1-
12
#972040000000
0!
0%
b10 *
0-
02
b10 6
#972050000000
1!
1%
1-
12
#972060000000
0!
0%
b11 *
0-
02
b11 6
#972070000000
1!
1%
1-
12
15
#972080000000
0!
0%
b100 *
0-
02
b100 6
#972090000000
1!
1%
1-
12
#972100000000
0!
0%
b101 *
0-
02
b101 6
#972110000000
1!
1%
1-
12
#972120000000
0!
0%
b110 *
0-
02
b110 6
#972130000000
1!
1%
1-
12
#972140000000
0!
0%
b111 *
0-
02
b111 6
#972150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#972160000000
0!
0%
b0 *
0-
02
b0 6
#972170000000
1!
1%
1-
12
#972180000000
0!
0%
b1 *
0-
02
b1 6
#972190000000
1!
1%
1-
12
#972200000000
0!
0%
b10 *
0-
02
b10 6
#972210000000
1!
1%
1-
12
#972220000000
0!
0%
b11 *
0-
02
b11 6
#972230000000
1!
1%
1-
12
15
#972240000000
0!
0%
b100 *
0-
02
b100 6
#972250000000
1!
1%
1-
12
#972260000000
0!
0%
b101 *
0-
02
b101 6
#972270000000
1!
1%
1-
12
#972280000000
0!
0%
b110 *
0-
02
b110 6
#972290000000
1!
1%
1-
12
#972300000000
0!
0%
b111 *
0-
02
b111 6
#972310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#972320000000
0!
0%
b0 *
0-
02
b0 6
#972330000000
1!
1%
1-
12
#972340000000
0!
0%
b1 *
0-
02
b1 6
#972350000000
1!
1%
1-
12
#972360000000
0!
0%
b10 *
0-
02
b10 6
#972370000000
1!
1%
1-
12
#972380000000
0!
0%
b11 *
0-
02
b11 6
#972390000000
1!
1%
1-
12
15
#972400000000
0!
0%
b100 *
0-
02
b100 6
#972410000000
1!
1%
1-
12
#972420000000
0!
0%
b101 *
0-
02
b101 6
#972430000000
1!
1%
1-
12
#972440000000
0!
0%
b110 *
0-
02
b110 6
#972450000000
1!
1%
1-
12
#972460000000
0!
0%
b111 *
0-
02
b111 6
#972470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#972480000000
0!
0%
b0 *
0-
02
b0 6
#972490000000
1!
1%
1-
12
#972500000000
0!
0%
b1 *
0-
02
b1 6
#972510000000
1!
1%
1-
12
#972520000000
0!
0%
b10 *
0-
02
b10 6
#972530000000
1!
1%
1-
12
#972540000000
0!
0%
b11 *
0-
02
b11 6
#972550000000
1!
1%
1-
12
15
#972560000000
0!
0%
b100 *
0-
02
b100 6
#972570000000
1!
1%
1-
12
#972580000000
0!
0%
b101 *
0-
02
b101 6
#972590000000
1!
1%
1-
12
#972600000000
0!
0%
b110 *
0-
02
b110 6
#972610000000
1!
1%
1-
12
#972620000000
0!
0%
b111 *
0-
02
b111 6
#972630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#972640000000
0!
0%
b0 *
0-
02
b0 6
#972650000000
1!
1%
1-
12
#972660000000
0!
0%
b1 *
0-
02
b1 6
#972670000000
1!
1%
1-
12
#972680000000
0!
0%
b10 *
0-
02
b10 6
#972690000000
1!
1%
1-
12
#972700000000
0!
0%
b11 *
0-
02
b11 6
#972710000000
1!
1%
1-
12
15
#972720000000
0!
0%
b100 *
0-
02
b100 6
#972730000000
1!
1%
1-
12
#972740000000
0!
0%
b101 *
0-
02
b101 6
#972750000000
1!
1%
1-
12
#972760000000
0!
0%
b110 *
0-
02
b110 6
#972770000000
1!
1%
1-
12
#972780000000
0!
0%
b111 *
0-
02
b111 6
#972790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#972800000000
0!
0%
b0 *
0-
02
b0 6
#972810000000
1!
1%
1-
12
#972820000000
0!
0%
b1 *
0-
02
b1 6
#972830000000
1!
1%
1-
12
#972840000000
0!
0%
b10 *
0-
02
b10 6
#972850000000
1!
1%
1-
12
#972860000000
0!
0%
b11 *
0-
02
b11 6
#972870000000
1!
1%
1-
12
15
#972880000000
0!
0%
b100 *
0-
02
b100 6
#972890000000
1!
1%
1-
12
#972900000000
0!
0%
b101 *
0-
02
b101 6
#972910000000
1!
1%
1-
12
#972920000000
0!
0%
b110 *
0-
02
b110 6
#972930000000
1!
1%
1-
12
#972940000000
0!
0%
b111 *
0-
02
b111 6
#972950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#972960000000
0!
0%
b0 *
0-
02
b0 6
#972970000000
1!
1%
1-
12
#972980000000
0!
0%
b1 *
0-
02
b1 6
#972990000000
1!
1%
1-
12
#973000000000
0!
0%
b10 *
0-
02
b10 6
#973010000000
1!
1%
1-
12
#973020000000
0!
0%
b11 *
0-
02
b11 6
#973030000000
1!
1%
1-
12
15
#973040000000
0!
0%
b100 *
0-
02
b100 6
#973050000000
1!
1%
1-
12
#973060000000
0!
0%
b101 *
0-
02
b101 6
#973070000000
1!
1%
1-
12
#973080000000
0!
0%
b110 *
0-
02
b110 6
#973090000000
1!
1%
1-
12
#973100000000
0!
0%
b111 *
0-
02
b111 6
#973110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#973120000000
0!
0%
b0 *
0-
02
b0 6
#973130000000
1!
1%
1-
12
#973140000000
0!
0%
b1 *
0-
02
b1 6
#973150000000
1!
1%
1-
12
#973160000000
0!
0%
b10 *
0-
02
b10 6
#973170000000
1!
1%
1-
12
#973180000000
0!
0%
b11 *
0-
02
b11 6
#973190000000
1!
1%
1-
12
15
#973200000000
0!
0%
b100 *
0-
02
b100 6
#973210000000
1!
1%
1-
12
#973220000000
0!
0%
b101 *
0-
02
b101 6
#973230000000
1!
1%
1-
12
#973240000000
0!
0%
b110 *
0-
02
b110 6
#973250000000
1!
1%
1-
12
#973260000000
0!
0%
b111 *
0-
02
b111 6
#973270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#973280000000
0!
0%
b0 *
0-
02
b0 6
#973290000000
1!
1%
1-
12
#973300000000
0!
0%
b1 *
0-
02
b1 6
#973310000000
1!
1%
1-
12
#973320000000
0!
0%
b10 *
0-
02
b10 6
#973330000000
1!
1%
1-
12
#973340000000
0!
0%
b11 *
0-
02
b11 6
#973350000000
1!
1%
1-
12
15
#973360000000
0!
0%
b100 *
0-
02
b100 6
#973370000000
1!
1%
1-
12
#973380000000
0!
0%
b101 *
0-
02
b101 6
#973390000000
1!
1%
1-
12
#973400000000
0!
0%
b110 *
0-
02
b110 6
#973410000000
1!
1%
1-
12
#973420000000
0!
0%
b111 *
0-
02
b111 6
#973430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#973440000000
0!
0%
b0 *
0-
02
b0 6
#973450000000
1!
1%
1-
12
#973460000000
0!
0%
b1 *
0-
02
b1 6
#973470000000
1!
1%
1-
12
#973480000000
0!
0%
b10 *
0-
02
b10 6
#973490000000
1!
1%
1-
12
#973500000000
0!
0%
b11 *
0-
02
b11 6
#973510000000
1!
1%
1-
12
15
#973520000000
0!
0%
b100 *
0-
02
b100 6
#973530000000
1!
1%
1-
12
#973540000000
0!
0%
b101 *
0-
02
b101 6
#973550000000
1!
1%
1-
12
#973560000000
0!
0%
b110 *
0-
02
b110 6
#973570000000
1!
1%
1-
12
#973580000000
0!
0%
b111 *
0-
02
b111 6
#973590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#973600000000
0!
0%
b0 *
0-
02
b0 6
#973610000000
1!
1%
1-
12
#973620000000
0!
0%
b1 *
0-
02
b1 6
#973630000000
1!
1%
1-
12
#973640000000
0!
0%
b10 *
0-
02
b10 6
#973650000000
1!
1%
1-
12
#973660000000
0!
0%
b11 *
0-
02
b11 6
#973670000000
1!
1%
1-
12
15
#973680000000
0!
0%
b100 *
0-
02
b100 6
#973690000000
1!
1%
1-
12
#973700000000
0!
0%
b101 *
0-
02
b101 6
#973710000000
1!
1%
1-
12
#973720000000
0!
0%
b110 *
0-
02
b110 6
#973730000000
1!
1%
1-
12
#973740000000
0!
0%
b111 *
0-
02
b111 6
#973750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#973760000000
0!
0%
b0 *
0-
02
b0 6
#973770000000
1!
1%
1-
12
#973780000000
0!
0%
b1 *
0-
02
b1 6
#973790000000
1!
1%
1-
12
#973800000000
0!
0%
b10 *
0-
02
b10 6
#973810000000
1!
1%
1-
12
#973820000000
0!
0%
b11 *
0-
02
b11 6
#973830000000
1!
1%
1-
12
15
#973840000000
0!
0%
b100 *
0-
02
b100 6
#973850000000
1!
1%
1-
12
#973860000000
0!
0%
b101 *
0-
02
b101 6
#973870000000
1!
1%
1-
12
#973880000000
0!
0%
b110 *
0-
02
b110 6
#973890000000
1!
1%
1-
12
#973900000000
0!
0%
b111 *
0-
02
b111 6
#973910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#973920000000
0!
0%
b0 *
0-
02
b0 6
#973930000000
1!
1%
1-
12
#973940000000
0!
0%
b1 *
0-
02
b1 6
#973950000000
1!
1%
1-
12
#973960000000
0!
0%
b10 *
0-
02
b10 6
#973970000000
1!
1%
1-
12
#973980000000
0!
0%
b11 *
0-
02
b11 6
#973990000000
1!
1%
1-
12
15
#974000000000
0!
0%
b100 *
0-
02
b100 6
#974010000000
1!
1%
1-
12
#974020000000
0!
0%
b101 *
0-
02
b101 6
#974030000000
1!
1%
1-
12
#974040000000
0!
0%
b110 *
0-
02
b110 6
#974050000000
1!
1%
1-
12
#974060000000
0!
0%
b111 *
0-
02
b111 6
#974070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#974080000000
0!
0%
b0 *
0-
02
b0 6
#974090000000
1!
1%
1-
12
#974100000000
0!
0%
b1 *
0-
02
b1 6
#974110000000
1!
1%
1-
12
#974120000000
0!
0%
b10 *
0-
02
b10 6
#974130000000
1!
1%
1-
12
#974140000000
0!
0%
b11 *
0-
02
b11 6
#974150000000
1!
1%
1-
12
15
#974160000000
0!
0%
b100 *
0-
02
b100 6
#974170000000
1!
1%
1-
12
#974180000000
0!
0%
b101 *
0-
02
b101 6
#974190000000
1!
1%
1-
12
#974200000000
0!
0%
b110 *
0-
02
b110 6
#974210000000
1!
1%
1-
12
#974220000000
0!
0%
b111 *
0-
02
b111 6
#974230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#974240000000
0!
0%
b0 *
0-
02
b0 6
#974250000000
1!
1%
1-
12
#974260000000
0!
0%
b1 *
0-
02
b1 6
#974270000000
1!
1%
1-
12
#974280000000
0!
0%
b10 *
0-
02
b10 6
#974290000000
1!
1%
1-
12
#974300000000
0!
0%
b11 *
0-
02
b11 6
#974310000000
1!
1%
1-
12
15
#974320000000
0!
0%
b100 *
0-
02
b100 6
#974330000000
1!
1%
1-
12
#974340000000
0!
0%
b101 *
0-
02
b101 6
#974350000000
1!
1%
1-
12
#974360000000
0!
0%
b110 *
0-
02
b110 6
#974370000000
1!
1%
1-
12
#974380000000
0!
0%
b111 *
0-
02
b111 6
#974390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#974400000000
0!
0%
b0 *
0-
02
b0 6
#974410000000
1!
1%
1-
12
#974420000000
0!
0%
b1 *
0-
02
b1 6
#974430000000
1!
1%
1-
12
#974440000000
0!
0%
b10 *
0-
02
b10 6
#974450000000
1!
1%
1-
12
#974460000000
0!
0%
b11 *
0-
02
b11 6
#974470000000
1!
1%
1-
12
15
#974480000000
0!
0%
b100 *
0-
02
b100 6
#974490000000
1!
1%
1-
12
#974500000000
0!
0%
b101 *
0-
02
b101 6
#974510000000
1!
1%
1-
12
#974520000000
0!
0%
b110 *
0-
02
b110 6
#974530000000
1!
1%
1-
12
#974540000000
0!
0%
b111 *
0-
02
b111 6
#974550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#974560000000
0!
0%
b0 *
0-
02
b0 6
#974570000000
1!
1%
1-
12
#974580000000
0!
0%
b1 *
0-
02
b1 6
#974590000000
1!
1%
1-
12
#974600000000
0!
0%
b10 *
0-
02
b10 6
#974610000000
1!
1%
1-
12
#974620000000
0!
0%
b11 *
0-
02
b11 6
#974630000000
1!
1%
1-
12
15
#974640000000
0!
0%
b100 *
0-
02
b100 6
#974650000000
1!
1%
1-
12
#974660000000
0!
0%
b101 *
0-
02
b101 6
#974670000000
1!
1%
1-
12
#974680000000
0!
0%
b110 *
0-
02
b110 6
#974690000000
1!
1%
1-
12
#974700000000
0!
0%
b111 *
0-
02
b111 6
#974710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#974720000000
0!
0%
b0 *
0-
02
b0 6
#974730000000
1!
1%
1-
12
#974740000000
0!
0%
b1 *
0-
02
b1 6
#974750000000
1!
1%
1-
12
#974760000000
0!
0%
b10 *
0-
02
b10 6
#974770000000
1!
1%
1-
12
#974780000000
0!
0%
b11 *
0-
02
b11 6
#974790000000
1!
1%
1-
12
15
#974800000000
0!
0%
b100 *
0-
02
b100 6
#974810000000
1!
1%
1-
12
#974820000000
0!
0%
b101 *
0-
02
b101 6
#974830000000
1!
1%
1-
12
#974840000000
0!
0%
b110 *
0-
02
b110 6
#974850000000
1!
1%
1-
12
#974860000000
0!
0%
b111 *
0-
02
b111 6
#974870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#974880000000
0!
0%
b0 *
0-
02
b0 6
#974890000000
1!
1%
1-
12
#974900000000
0!
0%
b1 *
0-
02
b1 6
#974910000000
1!
1%
1-
12
#974920000000
0!
0%
b10 *
0-
02
b10 6
#974930000000
1!
1%
1-
12
#974940000000
0!
0%
b11 *
0-
02
b11 6
#974950000000
1!
1%
1-
12
15
#974960000000
0!
0%
b100 *
0-
02
b100 6
#974970000000
1!
1%
1-
12
#974980000000
0!
0%
b101 *
0-
02
b101 6
#974990000000
1!
1%
1-
12
#975000000000
0!
0%
b110 *
0-
02
b110 6
#975010000000
1!
1%
1-
12
#975020000000
0!
0%
b111 *
0-
02
b111 6
#975030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#975040000000
0!
0%
b0 *
0-
02
b0 6
#975050000000
1!
1%
1-
12
#975060000000
0!
0%
b1 *
0-
02
b1 6
#975070000000
1!
1%
1-
12
#975080000000
0!
0%
b10 *
0-
02
b10 6
#975090000000
1!
1%
1-
12
#975100000000
0!
0%
b11 *
0-
02
b11 6
#975110000000
1!
1%
1-
12
15
#975120000000
0!
0%
b100 *
0-
02
b100 6
#975130000000
1!
1%
1-
12
#975140000000
0!
0%
b101 *
0-
02
b101 6
#975150000000
1!
1%
1-
12
#975160000000
0!
0%
b110 *
0-
02
b110 6
#975170000000
1!
1%
1-
12
#975180000000
0!
0%
b111 *
0-
02
b111 6
#975190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#975200000000
0!
0%
b0 *
0-
02
b0 6
#975210000000
1!
1%
1-
12
#975220000000
0!
0%
b1 *
0-
02
b1 6
#975230000000
1!
1%
1-
12
#975240000000
0!
0%
b10 *
0-
02
b10 6
#975250000000
1!
1%
1-
12
#975260000000
0!
0%
b11 *
0-
02
b11 6
#975270000000
1!
1%
1-
12
15
#975280000000
0!
0%
b100 *
0-
02
b100 6
#975290000000
1!
1%
1-
12
#975300000000
0!
0%
b101 *
0-
02
b101 6
#975310000000
1!
1%
1-
12
#975320000000
0!
0%
b110 *
0-
02
b110 6
#975330000000
1!
1%
1-
12
#975340000000
0!
0%
b111 *
0-
02
b111 6
#975350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#975360000000
0!
0%
b0 *
0-
02
b0 6
#975370000000
1!
1%
1-
12
#975380000000
0!
0%
b1 *
0-
02
b1 6
#975390000000
1!
1%
1-
12
#975400000000
0!
0%
b10 *
0-
02
b10 6
#975410000000
1!
1%
1-
12
#975420000000
0!
0%
b11 *
0-
02
b11 6
#975430000000
1!
1%
1-
12
15
#975440000000
0!
0%
b100 *
0-
02
b100 6
#975450000000
1!
1%
1-
12
#975460000000
0!
0%
b101 *
0-
02
b101 6
#975470000000
1!
1%
1-
12
#975480000000
0!
0%
b110 *
0-
02
b110 6
#975490000000
1!
1%
1-
12
#975500000000
0!
0%
b111 *
0-
02
b111 6
#975510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#975520000000
0!
0%
b0 *
0-
02
b0 6
#975530000000
1!
1%
1-
12
#975540000000
0!
0%
b1 *
0-
02
b1 6
#975550000000
1!
1%
1-
12
#975560000000
0!
0%
b10 *
0-
02
b10 6
#975570000000
1!
1%
1-
12
#975580000000
0!
0%
b11 *
0-
02
b11 6
#975590000000
1!
1%
1-
12
15
#975600000000
0!
0%
b100 *
0-
02
b100 6
#975610000000
1!
1%
1-
12
#975620000000
0!
0%
b101 *
0-
02
b101 6
#975630000000
1!
1%
1-
12
#975640000000
0!
0%
b110 *
0-
02
b110 6
#975650000000
1!
1%
1-
12
#975660000000
0!
0%
b111 *
0-
02
b111 6
#975670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#975680000000
0!
0%
b0 *
0-
02
b0 6
#975690000000
1!
1%
1-
12
#975700000000
0!
0%
b1 *
0-
02
b1 6
#975710000000
1!
1%
1-
12
#975720000000
0!
0%
b10 *
0-
02
b10 6
#975730000000
1!
1%
1-
12
#975740000000
0!
0%
b11 *
0-
02
b11 6
#975750000000
1!
1%
1-
12
15
#975760000000
0!
0%
b100 *
0-
02
b100 6
#975770000000
1!
1%
1-
12
#975780000000
0!
0%
b101 *
0-
02
b101 6
#975790000000
1!
1%
1-
12
#975800000000
0!
0%
b110 *
0-
02
b110 6
#975810000000
1!
1%
1-
12
#975820000000
0!
0%
b111 *
0-
02
b111 6
#975830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#975840000000
0!
0%
b0 *
0-
02
b0 6
#975850000000
1!
1%
1-
12
#975860000000
0!
0%
b1 *
0-
02
b1 6
#975870000000
1!
1%
1-
12
#975880000000
0!
0%
b10 *
0-
02
b10 6
#975890000000
1!
1%
1-
12
#975900000000
0!
0%
b11 *
0-
02
b11 6
#975910000000
1!
1%
1-
12
15
#975920000000
0!
0%
b100 *
0-
02
b100 6
#975930000000
1!
1%
1-
12
#975940000000
0!
0%
b101 *
0-
02
b101 6
#975950000000
1!
1%
1-
12
#975960000000
0!
0%
b110 *
0-
02
b110 6
#975970000000
1!
1%
1-
12
#975980000000
0!
0%
b111 *
0-
02
b111 6
#975990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#976000000000
0!
0%
b0 *
0-
02
b0 6
#976010000000
1!
1%
1-
12
#976020000000
0!
0%
b1 *
0-
02
b1 6
#976030000000
1!
1%
1-
12
#976040000000
0!
0%
b10 *
0-
02
b10 6
#976050000000
1!
1%
1-
12
#976060000000
0!
0%
b11 *
0-
02
b11 6
#976070000000
1!
1%
1-
12
15
#976080000000
0!
0%
b100 *
0-
02
b100 6
#976090000000
1!
1%
1-
12
#976100000000
0!
0%
b101 *
0-
02
b101 6
#976110000000
1!
1%
1-
12
#976120000000
0!
0%
b110 *
0-
02
b110 6
#976130000000
1!
1%
1-
12
#976140000000
0!
0%
b111 *
0-
02
b111 6
#976150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#976160000000
0!
0%
b0 *
0-
02
b0 6
#976170000000
1!
1%
1-
12
#976180000000
0!
0%
b1 *
0-
02
b1 6
#976190000000
1!
1%
1-
12
#976200000000
0!
0%
b10 *
0-
02
b10 6
#976210000000
1!
1%
1-
12
#976220000000
0!
0%
b11 *
0-
02
b11 6
#976230000000
1!
1%
1-
12
15
#976240000000
0!
0%
b100 *
0-
02
b100 6
#976250000000
1!
1%
1-
12
#976260000000
0!
0%
b101 *
0-
02
b101 6
#976270000000
1!
1%
1-
12
#976280000000
0!
0%
b110 *
0-
02
b110 6
#976290000000
1!
1%
1-
12
#976300000000
0!
0%
b111 *
0-
02
b111 6
#976310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#976320000000
0!
0%
b0 *
0-
02
b0 6
#976330000000
1!
1%
1-
12
#976340000000
0!
0%
b1 *
0-
02
b1 6
#976350000000
1!
1%
1-
12
#976360000000
0!
0%
b10 *
0-
02
b10 6
#976370000000
1!
1%
1-
12
#976380000000
0!
0%
b11 *
0-
02
b11 6
#976390000000
1!
1%
1-
12
15
#976400000000
0!
0%
b100 *
0-
02
b100 6
#976410000000
1!
1%
1-
12
#976420000000
0!
0%
b101 *
0-
02
b101 6
#976430000000
1!
1%
1-
12
#976440000000
0!
0%
b110 *
0-
02
b110 6
#976450000000
1!
1%
1-
12
#976460000000
0!
0%
b111 *
0-
02
b111 6
#976470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#976480000000
0!
0%
b0 *
0-
02
b0 6
#976490000000
1!
1%
1-
12
#976500000000
0!
0%
b1 *
0-
02
b1 6
#976510000000
1!
1%
1-
12
#976520000000
0!
0%
b10 *
0-
02
b10 6
#976530000000
1!
1%
1-
12
#976540000000
0!
0%
b11 *
0-
02
b11 6
#976550000000
1!
1%
1-
12
15
#976560000000
0!
0%
b100 *
0-
02
b100 6
#976570000000
1!
1%
1-
12
#976580000000
0!
0%
b101 *
0-
02
b101 6
#976590000000
1!
1%
1-
12
#976600000000
0!
0%
b110 *
0-
02
b110 6
#976610000000
1!
1%
1-
12
#976620000000
0!
0%
b111 *
0-
02
b111 6
#976630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#976640000000
0!
0%
b0 *
0-
02
b0 6
#976650000000
1!
1%
1-
12
#976660000000
0!
0%
b1 *
0-
02
b1 6
#976670000000
1!
1%
1-
12
#976680000000
0!
0%
b10 *
0-
02
b10 6
#976690000000
1!
1%
1-
12
#976700000000
0!
0%
b11 *
0-
02
b11 6
#976710000000
1!
1%
1-
12
15
#976720000000
0!
0%
b100 *
0-
02
b100 6
#976730000000
1!
1%
1-
12
#976740000000
0!
0%
b101 *
0-
02
b101 6
#976750000000
1!
1%
1-
12
#976760000000
0!
0%
b110 *
0-
02
b110 6
#976770000000
1!
1%
1-
12
#976780000000
0!
0%
b111 *
0-
02
b111 6
#976790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#976800000000
0!
0%
b0 *
0-
02
b0 6
#976810000000
1!
1%
1-
12
#976820000000
0!
0%
b1 *
0-
02
b1 6
#976830000000
1!
1%
1-
12
#976840000000
0!
0%
b10 *
0-
02
b10 6
#976850000000
1!
1%
1-
12
#976860000000
0!
0%
b11 *
0-
02
b11 6
#976870000000
1!
1%
1-
12
15
#976880000000
0!
0%
b100 *
0-
02
b100 6
#976890000000
1!
1%
1-
12
#976900000000
0!
0%
b101 *
0-
02
b101 6
#976910000000
1!
1%
1-
12
#976920000000
0!
0%
b110 *
0-
02
b110 6
#976930000000
1!
1%
1-
12
#976940000000
0!
0%
b111 *
0-
02
b111 6
#976950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#976960000000
0!
0%
b0 *
0-
02
b0 6
#976970000000
1!
1%
1-
12
#976980000000
0!
0%
b1 *
0-
02
b1 6
#976990000000
1!
1%
1-
12
#977000000000
0!
0%
b10 *
0-
02
b10 6
#977010000000
1!
1%
1-
12
#977020000000
0!
0%
b11 *
0-
02
b11 6
#977030000000
1!
1%
1-
12
15
#977040000000
0!
0%
b100 *
0-
02
b100 6
#977050000000
1!
1%
1-
12
#977060000000
0!
0%
b101 *
0-
02
b101 6
#977070000000
1!
1%
1-
12
#977080000000
0!
0%
b110 *
0-
02
b110 6
#977090000000
1!
1%
1-
12
#977100000000
0!
0%
b111 *
0-
02
b111 6
#977110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#977120000000
0!
0%
b0 *
0-
02
b0 6
#977130000000
1!
1%
1-
12
#977140000000
0!
0%
b1 *
0-
02
b1 6
#977150000000
1!
1%
1-
12
#977160000000
0!
0%
b10 *
0-
02
b10 6
#977170000000
1!
1%
1-
12
#977180000000
0!
0%
b11 *
0-
02
b11 6
#977190000000
1!
1%
1-
12
15
#977200000000
0!
0%
b100 *
0-
02
b100 6
#977210000000
1!
1%
1-
12
#977220000000
0!
0%
b101 *
0-
02
b101 6
#977230000000
1!
1%
1-
12
#977240000000
0!
0%
b110 *
0-
02
b110 6
#977250000000
1!
1%
1-
12
#977260000000
0!
0%
b111 *
0-
02
b111 6
#977270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#977280000000
0!
0%
b0 *
0-
02
b0 6
#977290000000
1!
1%
1-
12
#977300000000
0!
0%
b1 *
0-
02
b1 6
#977310000000
1!
1%
1-
12
#977320000000
0!
0%
b10 *
0-
02
b10 6
#977330000000
1!
1%
1-
12
#977340000000
0!
0%
b11 *
0-
02
b11 6
#977350000000
1!
1%
1-
12
15
#977360000000
0!
0%
b100 *
0-
02
b100 6
#977370000000
1!
1%
1-
12
#977380000000
0!
0%
b101 *
0-
02
b101 6
#977390000000
1!
1%
1-
12
#977400000000
0!
0%
b110 *
0-
02
b110 6
#977410000000
1!
1%
1-
12
#977420000000
0!
0%
b111 *
0-
02
b111 6
#977430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#977440000000
0!
0%
b0 *
0-
02
b0 6
#977450000000
1!
1%
1-
12
#977460000000
0!
0%
b1 *
0-
02
b1 6
#977470000000
1!
1%
1-
12
#977480000000
0!
0%
b10 *
0-
02
b10 6
#977490000000
1!
1%
1-
12
#977500000000
0!
0%
b11 *
0-
02
b11 6
#977510000000
1!
1%
1-
12
15
#977520000000
0!
0%
b100 *
0-
02
b100 6
#977530000000
1!
1%
1-
12
#977540000000
0!
0%
b101 *
0-
02
b101 6
#977550000000
1!
1%
1-
12
#977560000000
0!
0%
b110 *
0-
02
b110 6
#977570000000
1!
1%
1-
12
#977580000000
0!
0%
b111 *
0-
02
b111 6
#977590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#977600000000
0!
0%
b0 *
0-
02
b0 6
#977610000000
1!
1%
1-
12
#977620000000
0!
0%
b1 *
0-
02
b1 6
#977630000000
1!
1%
1-
12
#977640000000
0!
0%
b10 *
0-
02
b10 6
#977650000000
1!
1%
1-
12
#977660000000
0!
0%
b11 *
0-
02
b11 6
#977670000000
1!
1%
1-
12
15
#977680000000
0!
0%
b100 *
0-
02
b100 6
#977690000000
1!
1%
1-
12
#977700000000
0!
0%
b101 *
0-
02
b101 6
#977710000000
1!
1%
1-
12
#977720000000
0!
0%
b110 *
0-
02
b110 6
#977730000000
1!
1%
1-
12
#977740000000
0!
0%
b111 *
0-
02
b111 6
#977750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#977760000000
0!
0%
b0 *
0-
02
b0 6
#977770000000
1!
1%
1-
12
#977780000000
0!
0%
b1 *
0-
02
b1 6
#977790000000
1!
1%
1-
12
#977800000000
0!
0%
b10 *
0-
02
b10 6
#977810000000
1!
1%
1-
12
#977820000000
0!
0%
b11 *
0-
02
b11 6
#977830000000
1!
1%
1-
12
15
#977840000000
0!
0%
b100 *
0-
02
b100 6
#977850000000
1!
1%
1-
12
#977860000000
0!
0%
b101 *
0-
02
b101 6
#977870000000
1!
1%
1-
12
#977880000000
0!
0%
b110 *
0-
02
b110 6
#977890000000
1!
1%
1-
12
#977900000000
0!
0%
b111 *
0-
02
b111 6
#977910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#977920000000
0!
0%
b0 *
0-
02
b0 6
#977930000000
1!
1%
1-
12
#977940000000
0!
0%
b1 *
0-
02
b1 6
#977950000000
1!
1%
1-
12
#977960000000
0!
0%
b10 *
0-
02
b10 6
#977970000000
1!
1%
1-
12
#977980000000
0!
0%
b11 *
0-
02
b11 6
#977990000000
1!
1%
1-
12
15
#978000000000
0!
0%
b100 *
0-
02
b100 6
#978010000000
1!
1%
1-
12
#978020000000
0!
0%
b101 *
0-
02
b101 6
#978030000000
1!
1%
1-
12
#978040000000
0!
0%
b110 *
0-
02
b110 6
#978050000000
1!
1%
1-
12
#978060000000
0!
0%
b111 *
0-
02
b111 6
#978070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#978080000000
0!
0%
b0 *
0-
02
b0 6
#978090000000
1!
1%
1-
12
#978100000000
0!
0%
b1 *
0-
02
b1 6
#978110000000
1!
1%
1-
12
#978120000000
0!
0%
b10 *
0-
02
b10 6
#978130000000
1!
1%
1-
12
#978140000000
0!
0%
b11 *
0-
02
b11 6
#978150000000
1!
1%
1-
12
15
#978160000000
0!
0%
b100 *
0-
02
b100 6
#978170000000
1!
1%
1-
12
#978180000000
0!
0%
b101 *
0-
02
b101 6
#978190000000
1!
1%
1-
12
#978200000000
0!
0%
b110 *
0-
02
b110 6
#978210000000
1!
1%
1-
12
#978220000000
0!
0%
b111 *
0-
02
b111 6
#978230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#978240000000
0!
0%
b0 *
0-
02
b0 6
#978250000000
1!
1%
1-
12
#978260000000
0!
0%
b1 *
0-
02
b1 6
#978270000000
1!
1%
1-
12
#978280000000
0!
0%
b10 *
0-
02
b10 6
#978290000000
1!
1%
1-
12
#978300000000
0!
0%
b11 *
0-
02
b11 6
#978310000000
1!
1%
1-
12
15
#978320000000
0!
0%
b100 *
0-
02
b100 6
#978330000000
1!
1%
1-
12
#978340000000
0!
0%
b101 *
0-
02
b101 6
#978350000000
1!
1%
1-
12
#978360000000
0!
0%
b110 *
0-
02
b110 6
#978370000000
1!
1%
1-
12
#978380000000
0!
0%
b111 *
0-
02
b111 6
#978390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#978400000000
0!
0%
b0 *
0-
02
b0 6
#978410000000
1!
1%
1-
12
#978420000000
0!
0%
b1 *
0-
02
b1 6
#978430000000
1!
1%
1-
12
#978440000000
0!
0%
b10 *
0-
02
b10 6
#978450000000
1!
1%
1-
12
#978460000000
0!
0%
b11 *
0-
02
b11 6
#978470000000
1!
1%
1-
12
15
#978480000000
0!
0%
b100 *
0-
02
b100 6
#978490000000
1!
1%
1-
12
#978500000000
0!
0%
b101 *
0-
02
b101 6
#978510000000
1!
1%
1-
12
#978520000000
0!
0%
b110 *
0-
02
b110 6
#978530000000
1!
1%
1-
12
#978540000000
0!
0%
b111 *
0-
02
b111 6
#978550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#978560000000
0!
0%
b0 *
0-
02
b0 6
#978570000000
1!
1%
1-
12
#978580000000
0!
0%
b1 *
0-
02
b1 6
#978590000000
1!
1%
1-
12
#978600000000
0!
0%
b10 *
0-
02
b10 6
#978610000000
1!
1%
1-
12
#978620000000
0!
0%
b11 *
0-
02
b11 6
#978630000000
1!
1%
1-
12
15
#978640000000
0!
0%
b100 *
0-
02
b100 6
#978650000000
1!
1%
1-
12
#978660000000
0!
0%
b101 *
0-
02
b101 6
#978670000000
1!
1%
1-
12
#978680000000
0!
0%
b110 *
0-
02
b110 6
#978690000000
1!
1%
1-
12
#978700000000
0!
0%
b111 *
0-
02
b111 6
#978710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#978720000000
0!
0%
b0 *
0-
02
b0 6
#978730000000
1!
1%
1-
12
#978740000000
0!
0%
b1 *
0-
02
b1 6
#978750000000
1!
1%
1-
12
#978760000000
0!
0%
b10 *
0-
02
b10 6
#978770000000
1!
1%
1-
12
#978780000000
0!
0%
b11 *
0-
02
b11 6
#978790000000
1!
1%
1-
12
15
#978800000000
0!
0%
b100 *
0-
02
b100 6
#978810000000
1!
1%
1-
12
#978820000000
0!
0%
b101 *
0-
02
b101 6
#978830000000
1!
1%
1-
12
#978840000000
0!
0%
b110 *
0-
02
b110 6
#978850000000
1!
1%
1-
12
#978860000000
0!
0%
b111 *
0-
02
b111 6
#978870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#978880000000
0!
0%
b0 *
0-
02
b0 6
#978890000000
1!
1%
1-
12
#978900000000
0!
0%
b1 *
0-
02
b1 6
#978910000000
1!
1%
1-
12
#978920000000
0!
0%
b10 *
0-
02
b10 6
#978930000000
1!
1%
1-
12
#978940000000
0!
0%
b11 *
0-
02
b11 6
#978950000000
1!
1%
1-
12
15
#978960000000
0!
0%
b100 *
0-
02
b100 6
#978970000000
1!
1%
1-
12
#978980000000
0!
0%
b101 *
0-
02
b101 6
#978990000000
1!
1%
1-
12
#979000000000
0!
0%
b110 *
0-
02
b110 6
#979010000000
1!
1%
1-
12
#979020000000
0!
0%
b111 *
0-
02
b111 6
#979030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#979040000000
0!
0%
b0 *
0-
02
b0 6
#979050000000
1!
1%
1-
12
#979060000000
0!
0%
b1 *
0-
02
b1 6
#979070000000
1!
1%
1-
12
#979080000000
0!
0%
b10 *
0-
02
b10 6
#979090000000
1!
1%
1-
12
#979100000000
0!
0%
b11 *
0-
02
b11 6
#979110000000
1!
1%
1-
12
15
#979120000000
0!
0%
b100 *
0-
02
b100 6
#979130000000
1!
1%
1-
12
#979140000000
0!
0%
b101 *
0-
02
b101 6
#979150000000
1!
1%
1-
12
#979160000000
0!
0%
b110 *
0-
02
b110 6
#979170000000
1!
1%
1-
12
#979180000000
0!
0%
b111 *
0-
02
b111 6
#979190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#979200000000
0!
0%
b0 *
0-
02
b0 6
#979210000000
1!
1%
1-
12
#979220000000
0!
0%
b1 *
0-
02
b1 6
#979230000000
1!
1%
1-
12
#979240000000
0!
0%
b10 *
0-
02
b10 6
#979250000000
1!
1%
1-
12
#979260000000
0!
0%
b11 *
0-
02
b11 6
#979270000000
1!
1%
1-
12
15
#979280000000
0!
0%
b100 *
0-
02
b100 6
#979290000000
1!
1%
1-
12
#979300000000
0!
0%
b101 *
0-
02
b101 6
#979310000000
1!
1%
1-
12
#979320000000
0!
0%
b110 *
0-
02
b110 6
#979330000000
1!
1%
1-
12
#979340000000
0!
0%
b111 *
0-
02
b111 6
#979350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#979360000000
0!
0%
b0 *
0-
02
b0 6
#979370000000
1!
1%
1-
12
#979380000000
0!
0%
b1 *
0-
02
b1 6
#979390000000
1!
1%
1-
12
#979400000000
0!
0%
b10 *
0-
02
b10 6
#979410000000
1!
1%
1-
12
#979420000000
0!
0%
b11 *
0-
02
b11 6
#979430000000
1!
1%
1-
12
15
#979440000000
0!
0%
b100 *
0-
02
b100 6
#979450000000
1!
1%
1-
12
#979460000000
0!
0%
b101 *
0-
02
b101 6
#979470000000
1!
1%
1-
12
#979480000000
0!
0%
b110 *
0-
02
b110 6
#979490000000
1!
1%
1-
12
#979500000000
0!
0%
b111 *
0-
02
b111 6
#979510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#979520000000
0!
0%
b0 *
0-
02
b0 6
#979530000000
1!
1%
1-
12
#979540000000
0!
0%
b1 *
0-
02
b1 6
#979550000000
1!
1%
1-
12
#979560000000
0!
0%
b10 *
0-
02
b10 6
#979570000000
1!
1%
1-
12
#979580000000
0!
0%
b11 *
0-
02
b11 6
#979590000000
1!
1%
1-
12
15
#979600000000
0!
0%
b100 *
0-
02
b100 6
#979610000000
1!
1%
1-
12
#979620000000
0!
0%
b101 *
0-
02
b101 6
#979630000000
1!
1%
1-
12
#979640000000
0!
0%
b110 *
0-
02
b110 6
#979650000000
1!
1%
1-
12
#979660000000
0!
0%
b111 *
0-
02
b111 6
#979670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#979680000000
0!
0%
b0 *
0-
02
b0 6
#979690000000
1!
1%
1-
12
#979700000000
0!
0%
b1 *
0-
02
b1 6
#979710000000
1!
1%
1-
12
#979720000000
0!
0%
b10 *
0-
02
b10 6
#979730000000
1!
1%
1-
12
#979740000000
0!
0%
b11 *
0-
02
b11 6
#979750000000
1!
1%
1-
12
15
#979760000000
0!
0%
b100 *
0-
02
b100 6
#979770000000
1!
1%
1-
12
#979780000000
0!
0%
b101 *
0-
02
b101 6
#979790000000
1!
1%
1-
12
#979800000000
0!
0%
b110 *
0-
02
b110 6
#979810000000
1!
1%
1-
12
#979820000000
0!
0%
b111 *
0-
02
b111 6
#979830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#979840000000
0!
0%
b0 *
0-
02
b0 6
#979850000000
1!
1%
1-
12
#979860000000
0!
0%
b1 *
0-
02
b1 6
#979870000000
1!
1%
1-
12
#979880000000
0!
0%
b10 *
0-
02
b10 6
#979890000000
1!
1%
1-
12
#979900000000
0!
0%
b11 *
0-
02
b11 6
#979910000000
1!
1%
1-
12
15
#979920000000
0!
0%
b100 *
0-
02
b100 6
#979930000000
1!
1%
1-
12
#979940000000
0!
0%
b101 *
0-
02
b101 6
#979950000000
1!
1%
1-
12
#979960000000
0!
0%
b110 *
0-
02
b110 6
#979970000000
1!
1%
1-
12
#979980000000
0!
0%
b111 *
0-
02
b111 6
#979990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#980000000000
0!
0%
b0 *
0-
02
b0 6
#980010000000
1!
1%
1-
12
#980020000000
0!
0%
b1 *
0-
02
b1 6
#980030000000
1!
1%
1-
12
#980040000000
0!
0%
b10 *
0-
02
b10 6
#980050000000
1!
1%
1-
12
#980060000000
0!
0%
b11 *
0-
02
b11 6
#980070000000
1!
1%
1-
12
15
#980080000000
0!
0%
b100 *
0-
02
b100 6
#980090000000
1!
1%
1-
12
#980100000000
0!
0%
b101 *
0-
02
b101 6
#980110000000
1!
1%
1-
12
#980120000000
0!
0%
b110 *
0-
02
b110 6
#980130000000
1!
1%
1-
12
#980140000000
0!
0%
b111 *
0-
02
b111 6
#980150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#980160000000
0!
0%
b0 *
0-
02
b0 6
#980170000000
1!
1%
1-
12
#980180000000
0!
0%
b1 *
0-
02
b1 6
#980190000000
1!
1%
1-
12
#980200000000
0!
0%
b10 *
0-
02
b10 6
#980210000000
1!
1%
1-
12
#980220000000
0!
0%
b11 *
0-
02
b11 6
#980230000000
1!
1%
1-
12
15
#980240000000
0!
0%
b100 *
0-
02
b100 6
#980250000000
1!
1%
1-
12
#980260000000
0!
0%
b101 *
0-
02
b101 6
#980270000000
1!
1%
1-
12
#980280000000
0!
0%
b110 *
0-
02
b110 6
#980290000000
1!
1%
1-
12
#980300000000
0!
0%
b111 *
0-
02
b111 6
#980310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#980320000000
0!
0%
b0 *
0-
02
b0 6
#980330000000
1!
1%
1-
12
#980340000000
0!
0%
b1 *
0-
02
b1 6
#980350000000
1!
1%
1-
12
#980360000000
0!
0%
b10 *
0-
02
b10 6
#980370000000
1!
1%
1-
12
#980380000000
0!
0%
b11 *
0-
02
b11 6
#980390000000
1!
1%
1-
12
15
#980400000000
0!
0%
b100 *
0-
02
b100 6
#980410000000
1!
1%
1-
12
#980420000000
0!
0%
b101 *
0-
02
b101 6
#980430000000
1!
1%
1-
12
#980440000000
0!
0%
b110 *
0-
02
b110 6
#980450000000
1!
1%
1-
12
#980460000000
0!
0%
b111 *
0-
02
b111 6
#980470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#980480000000
0!
0%
b0 *
0-
02
b0 6
#980490000000
1!
1%
1-
12
#980500000000
0!
0%
b1 *
0-
02
b1 6
#980510000000
1!
1%
1-
12
#980520000000
0!
0%
b10 *
0-
02
b10 6
#980530000000
1!
1%
1-
12
#980540000000
0!
0%
b11 *
0-
02
b11 6
#980550000000
1!
1%
1-
12
15
#980560000000
0!
0%
b100 *
0-
02
b100 6
#980570000000
1!
1%
1-
12
#980580000000
0!
0%
b101 *
0-
02
b101 6
#980590000000
1!
1%
1-
12
#980600000000
0!
0%
b110 *
0-
02
b110 6
#980610000000
1!
1%
1-
12
#980620000000
0!
0%
b111 *
0-
02
b111 6
#980630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#980640000000
0!
0%
b0 *
0-
02
b0 6
#980650000000
1!
1%
1-
12
#980660000000
0!
0%
b1 *
0-
02
b1 6
#980670000000
1!
1%
1-
12
#980680000000
0!
0%
b10 *
0-
02
b10 6
#980690000000
1!
1%
1-
12
#980700000000
0!
0%
b11 *
0-
02
b11 6
#980710000000
1!
1%
1-
12
15
#980720000000
0!
0%
b100 *
0-
02
b100 6
#980730000000
1!
1%
1-
12
#980740000000
0!
0%
b101 *
0-
02
b101 6
#980750000000
1!
1%
1-
12
#980760000000
0!
0%
b110 *
0-
02
b110 6
#980770000000
1!
1%
1-
12
#980780000000
0!
0%
b111 *
0-
02
b111 6
#980790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#980800000000
0!
0%
b0 *
0-
02
b0 6
#980810000000
1!
1%
1-
12
#980820000000
0!
0%
b1 *
0-
02
b1 6
#980830000000
1!
1%
1-
12
#980840000000
0!
0%
b10 *
0-
02
b10 6
#980850000000
1!
1%
1-
12
#980860000000
0!
0%
b11 *
0-
02
b11 6
#980870000000
1!
1%
1-
12
15
#980880000000
0!
0%
b100 *
0-
02
b100 6
#980890000000
1!
1%
1-
12
#980900000000
0!
0%
b101 *
0-
02
b101 6
#980910000000
1!
1%
1-
12
#980920000000
0!
0%
b110 *
0-
02
b110 6
#980930000000
1!
1%
1-
12
#980940000000
0!
0%
b111 *
0-
02
b111 6
#980950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#980960000000
0!
0%
b0 *
0-
02
b0 6
#980970000000
1!
1%
1-
12
#980980000000
0!
0%
b1 *
0-
02
b1 6
#980990000000
1!
1%
1-
12
#981000000000
0!
0%
b10 *
0-
02
b10 6
#981010000000
1!
1%
1-
12
#981020000000
0!
0%
b11 *
0-
02
b11 6
#981030000000
1!
1%
1-
12
15
#981040000000
0!
0%
b100 *
0-
02
b100 6
#981050000000
1!
1%
1-
12
#981060000000
0!
0%
b101 *
0-
02
b101 6
#981070000000
1!
1%
1-
12
#981080000000
0!
0%
b110 *
0-
02
b110 6
#981090000000
1!
1%
1-
12
#981100000000
0!
0%
b111 *
0-
02
b111 6
#981110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#981120000000
0!
0%
b0 *
0-
02
b0 6
#981130000000
1!
1%
1-
12
#981140000000
0!
0%
b1 *
0-
02
b1 6
#981150000000
1!
1%
1-
12
#981160000000
0!
0%
b10 *
0-
02
b10 6
#981170000000
1!
1%
1-
12
#981180000000
0!
0%
b11 *
0-
02
b11 6
#981190000000
1!
1%
1-
12
15
#981200000000
0!
0%
b100 *
0-
02
b100 6
#981210000000
1!
1%
1-
12
#981220000000
0!
0%
b101 *
0-
02
b101 6
#981230000000
1!
1%
1-
12
#981240000000
0!
0%
b110 *
0-
02
b110 6
#981250000000
1!
1%
1-
12
#981260000000
0!
0%
b111 *
0-
02
b111 6
#981270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#981280000000
0!
0%
b0 *
0-
02
b0 6
#981290000000
1!
1%
1-
12
#981300000000
0!
0%
b1 *
0-
02
b1 6
#981310000000
1!
1%
1-
12
#981320000000
0!
0%
b10 *
0-
02
b10 6
#981330000000
1!
1%
1-
12
#981340000000
0!
0%
b11 *
0-
02
b11 6
#981350000000
1!
1%
1-
12
15
#981360000000
0!
0%
b100 *
0-
02
b100 6
#981370000000
1!
1%
1-
12
#981380000000
0!
0%
b101 *
0-
02
b101 6
#981390000000
1!
1%
1-
12
#981400000000
0!
0%
b110 *
0-
02
b110 6
#981410000000
1!
1%
1-
12
#981420000000
0!
0%
b111 *
0-
02
b111 6
#981430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#981440000000
0!
0%
b0 *
0-
02
b0 6
#981450000000
1!
1%
1-
12
#981460000000
0!
0%
b1 *
0-
02
b1 6
#981470000000
1!
1%
1-
12
#981480000000
0!
0%
b10 *
0-
02
b10 6
#981490000000
1!
1%
1-
12
#981500000000
0!
0%
b11 *
0-
02
b11 6
#981510000000
1!
1%
1-
12
15
#981520000000
0!
0%
b100 *
0-
02
b100 6
#981530000000
1!
1%
1-
12
#981540000000
0!
0%
b101 *
0-
02
b101 6
#981550000000
1!
1%
1-
12
#981560000000
0!
0%
b110 *
0-
02
b110 6
#981570000000
1!
1%
1-
12
#981580000000
0!
0%
b111 *
0-
02
b111 6
#981590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#981600000000
0!
0%
b0 *
0-
02
b0 6
#981610000000
1!
1%
1-
12
#981620000000
0!
0%
b1 *
0-
02
b1 6
#981630000000
1!
1%
1-
12
#981640000000
0!
0%
b10 *
0-
02
b10 6
#981650000000
1!
1%
1-
12
#981660000000
0!
0%
b11 *
0-
02
b11 6
#981670000000
1!
1%
1-
12
15
#981680000000
0!
0%
b100 *
0-
02
b100 6
#981690000000
1!
1%
1-
12
#981700000000
0!
0%
b101 *
0-
02
b101 6
#981710000000
1!
1%
1-
12
#981720000000
0!
0%
b110 *
0-
02
b110 6
#981730000000
1!
1%
1-
12
#981740000000
0!
0%
b111 *
0-
02
b111 6
#981750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#981760000000
0!
0%
b0 *
0-
02
b0 6
#981770000000
1!
1%
1-
12
#981780000000
0!
0%
b1 *
0-
02
b1 6
#981790000000
1!
1%
1-
12
#981800000000
0!
0%
b10 *
0-
02
b10 6
#981810000000
1!
1%
1-
12
#981820000000
0!
0%
b11 *
0-
02
b11 6
#981830000000
1!
1%
1-
12
15
#981840000000
0!
0%
b100 *
0-
02
b100 6
#981850000000
1!
1%
1-
12
#981860000000
0!
0%
b101 *
0-
02
b101 6
#981870000000
1!
1%
1-
12
#981880000000
0!
0%
b110 *
0-
02
b110 6
#981890000000
1!
1%
1-
12
#981900000000
0!
0%
b111 *
0-
02
b111 6
#981910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#981920000000
0!
0%
b0 *
0-
02
b0 6
#981930000000
1!
1%
1-
12
#981940000000
0!
0%
b1 *
0-
02
b1 6
#981950000000
1!
1%
1-
12
#981960000000
0!
0%
b10 *
0-
02
b10 6
#981970000000
1!
1%
1-
12
#981980000000
0!
0%
b11 *
0-
02
b11 6
#981990000000
1!
1%
1-
12
15
#982000000000
0!
0%
b100 *
0-
02
b100 6
#982010000000
1!
1%
1-
12
#982020000000
0!
0%
b101 *
0-
02
b101 6
#982030000000
1!
1%
1-
12
#982040000000
0!
0%
b110 *
0-
02
b110 6
#982050000000
1!
1%
1-
12
#982060000000
0!
0%
b111 *
0-
02
b111 6
#982070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#982080000000
0!
0%
b0 *
0-
02
b0 6
#982090000000
1!
1%
1-
12
#982100000000
0!
0%
b1 *
0-
02
b1 6
#982110000000
1!
1%
1-
12
#982120000000
0!
0%
b10 *
0-
02
b10 6
#982130000000
1!
1%
1-
12
#982140000000
0!
0%
b11 *
0-
02
b11 6
#982150000000
1!
1%
1-
12
15
#982160000000
0!
0%
b100 *
0-
02
b100 6
#982170000000
1!
1%
1-
12
#982180000000
0!
0%
b101 *
0-
02
b101 6
#982190000000
1!
1%
1-
12
#982200000000
0!
0%
b110 *
0-
02
b110 6
#982210000000
1!
1%
1-
12
#982220000000
0!
0%
b111 *
0-
02
b111 6
#982230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#982240000000
0!
0%
b0 *
0-
02
b0 6
#982250000000
1!
1%
1-
12
#982260000000
0!
0%
b1 *
0-
02
b1 6
#982270000000
1!
1%
1-
12
#982280000000
0!
0%
b10 *
0-
02
b10 6
#982290000000
1!
1%
1-
12
#982300000000
0!
0%
b11 *
0-
02
b11 6
#982310000000
1!
1%
1-
12
15
#982320000000
0!
0%
b100 *
0-
02
b100 6
#982330000000
1!
1%
1-
12
#982340000000
0!
0%
b101 *
0-
02
b101 6
#982350000000
1!
1%
1-
12
#982360000000
0!
0%
b110 *
0-
02
b110 6
#982370000000
1!
1%
1-
12
#982380000000
0!
0%
b111 *
0-
02
b111 6
#982390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#982400000000
0!
0%
b0 *
0-
02
b0 6
#982410000000
1!
1%
1-
12
#982420000000
0!
0%
b1 *
0-
02
b1 6
#982430000000
1!
1%
1-
12
#982440000000
0!
0%
b10 *
0-
02
b10 6
#982450000000
1!
1%
1-
12
#982460000000
0!
0%
b11 *
0-
02
b11 6
#982470000000
1!
1%
1-
12
15
#982480000000
0!
0%
b100 *
0-
02
b100 6
#982490000000
1!
1%
1-
12
#982500000000
0!
0%
b101 *
0-
02
b101 6
#982510000000
1!
1%
1-
12
#982520000000
0!
0%
b110 *
0-
02
b110 6
#982530000000
1!
1%
1-
12
#982540000000
0!
0%
b111 *
0-
02
b111 6
#982550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#982560000000
0!
0%
b0 *
0-
02
b0 6
#982570000000
1!
1%
1-
12
#982580000000
0!
0%
b1 *
0-
02
b1 6
#982590000000
1!
1%
1-
12
#982600000000
0!
0%
b10 *
0-
02
b10 6
#982610000000
1!
1%
1-
12
#982620000000
0!
0%
b11 *
0-
02
b11 6
#982630000000
1!
1%
1-
12
15
#982640000000
0!
0%
b100 *
0-
02
b100 6
#982650000000
1!
1%
1-
12
#982660000000
0!
0%
b101 *
0-
02
b101 6
#982670000000
1!
1%
1-
12
#982680000000
0!
0%
b110 *
0-
02
b110 6
#982690000000
1!
1%
1-
12
#982700000000
0!
0%
b111 *
0-
02
b111 6
#982710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#982720000000
0!
0%
b0 *
0-
02
b0 6
#982730000000
1!
1%
1-
12
#982740000000
0!
0%
b1 *
0-
02
b1 6
#982750000000
1!
1%
1-
12
#982760000000
0!
0%
b10 *
0-
02
b10 6
#982770000000
1!
1%
1-
12
#982780000000
0!
0%
b11 *
0-
02
b11 6
#982790000000
1!
1%
1-
12
15
#982800000000
0!
0%
b100 *
0-
02
b100 6
#982810000000
1!
1%
1-
12
#982820000000
0!
0%
b101 *
0-
02
b101 6
#982830000000
1!
1%
1-
12
#982840000000
0!
0%
b110 *
0-
02
b110 6
#982850000000
1!
1%
1-
12
#982860000000
0!
0%
b111 *
0-
02
b111 6
#982870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#982880000000
0!
0%
b0 *
0-
02
b0 6
#982890000000
1!
1%
1-
12
#982900000000
0!
0%
b1 *
0-
02
b1 6
#982910000000
1!
1%
1-
12
#982920000000
0!
0%
b10 *
0-
02
b10 6
#982930000000
1!
1%
1-
12
#982940000000
0!
0%
b11 *
0-
02
b11 6
#982950000000
1!
1%
1-
12
15
#982960000000
0!
0%
b100 *
0-
02
b100 6
#982970000000
1!
1%
1-
12
#982980000000
0!
0%
b101 *
0-
02
b101 6
#982990000000
1!
1%
1-
12
#983000000000
0!
0%
b110 *
0-
02
b110 6
#983010000000
1!
1%
1-
12
#983020000000
0!
0%
b111 *
0-
02
b111 6
#983030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#983040000000
0!
0%
b0 *
0-
02
b0 6
#983050000000
1!
1%
1-
12
#983060000000
0!
0%
b1 *
0-
02
b1 6
#983070000000
1!
1%
1-
12
#983080000000
0!
0%
b10 *
0-
02
b10 6
#983090000000
1!
1%
1-
12
#983100000000
0!
0%
b11 *
0-
02
b11 6
#983110000000
1!
1%
1-
12
15
#983120000000
0!
0%
b100 *
0-
02
b100 6
#983130000000
1!
1%
1-
12
#983140000000
0!
0%
b101 *
0-
02
b101 6
#983150000000
1!
1%
1-
12
#983160000000
0!
0%
b110 *
0-
02
b110 6
#983170000000
1!
1%
1-
12
#983180000000
0!
0%
b111 *
0-
02
b111 6
#983190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#983200000000
0!
0%
b0 *
0-
02
b0 6
#983210000000
1!
1%
1-
12
#983220000000
0!
0%
b1 *
0-
02
b1 6
#983230000000
1!
1%
1-
12
#983240000000
0!
0%
b10 *
0-
02
b10 6
#983250000000
1!
1%
1-
12
#983260000000
0!
0%
b11 *
0-
02
b11 6
#983270000000
1!
1%
1-
12
15
#983280000000
0!
0%
b100 *
0-
02
b100 6
#983290000000
1!
1%
1-
12
#983300000000
0!
0%
b101 *
0-
02
b101 6
#983310000000
1!
1%
1-
12
#983320000000
0!
0%
b110 *
0-
02
b110 6
#983330000000
1!
1%
1-
12
#983340000000
0!
0%
b111 *
0-
02
b111 6
#983350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#983360000000
0!
0%
b0 *
0-
02
b0 6
#983370000000
1!
1%
1-
12
#983380000000
0!
0%
b1 *
0-
02
b1 6
#983390000000
1!
1%
1-
12
#983400000000
0!
0%
b10 *
0-
02
b10 6
#983410000000
1!
1%
1-
12
#983420000000
0!
0%
b11 *
0-
02
b11 6
#983430000000
1!
1%
1-
12
15
#983440000000
0!
0%
b100 *
0-
02
b100 6
#983450000000
1!
1%
1-
12
#983460000000
0!
0%
b101 *
0-
02
b101 6
#983470000000
1!
1%
1-
12
#983480000000
0!
0%
b110 *
0-
02
b110 6
#983490000000
1!
1%
1-
12
#983500000000
0!
0%
b111 *
0-
02
b111 6
#983510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#983520000000
0!
0%
b0 *
0-
02
b0 6
#983530000000
1!
1%
1-
12
#983540000000
0!
0%
b1 *
0-
02
b1 6
#983550000000
1!
1%
1-
12
#983560000000
0!
0%
b10 *
0-
02
b10 6
#983570000000
1!
1%
1-
12
#983580000000
0!
0%
b11 *
0-
02
b11 6
#983590000000
1!
1%
1-
12
15
#983600000000
0!
0%
b100 *
0-
02
b100 6
#983610000000
1!
1%
1-
12
#983620000000
0!
0%
b101 *
0-
02
b101 6
#983630000000
1!
1%
1-
12
#983640000000
0!
0%
b110 *
0-
02
b110 6
#983650000000
1!
1%
1-
12
#983660000000
0!
0%
b111 *
0-
02
b111 6
#983670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#983680000000
0!
0%
b0 *
0-
02
b0 6
#983690000000
1!
1%
1-
12
#983700000000
0!
0%
b1 *
0-
02
b1 6
#983710000000
1!
1%
1-
12
#983720000000
0!
0%
b10 *
0-
02
b10 6
#983730000000
1!
1%
1-
12
#983740000000
0!
0%
b11 *
0-
02
b11 6
#983750000000
1!
1%
1-
12
15
#983760000000
0!
0%
b100 *
0-
02
b100 6
#983770000000
1!
1%
1-
12
#983780000000
0!
0%
b101 *
0-
02
b101 6
#983790000000
1!
1%
1-
12
#983800000000
0!
0%
b110 *
0-
02
b110 6
#983810000000
1!
1%
1-
12
#983820000000
0!
0%
b111 *
0-
02
b111 6
#983830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#983840000000
0!
0%
b0 *
0-
02
b0 6
#983850000000
1!
1%
1-
12
#983860000000
0!
0%
b1 *
0-
02
b1 6
#983870000000
1!
1%
1-
12
#983880000000
0!
0%
b10 *
0-
02
b10 6
#983890000000
1!
1%
1-
12
#983900000000
0!
0%
b11 *
0-
02
b11 6
#983910000000
1!
1%
1-
12
15
#983920000000
0!
0%
b100 *
0-
02
b100 6
#983930000000
1!
1%
1-
12
#983940000000
0!
0%
b101 *
0-
02
b101 6
#983950000000
1!
1%
1-
12
#983960000000
0!
0%
b110 *
0-
02
b110 6
#983970000000
1!
1%
1-
12
#983980000000
0!
0%
b111 *
0-
02
b111 6
#983990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#984000000000
0!
0%
b0 *
0-
02
b0 6
#984010000000
1!
1%
1-
12
#984020000000
0!
0%
b1 *
0-
02
b1 6
#984030000000
1!
1%
1-
12
#984040000000
0!
0%
b10 *
0-
02
b10 6
#984050000000
1!
1%
1-
12
#984060000000
0!
0%
b11 *
0-
02
b11 6
#984070000000
1!
1%
1-
12
15
#984080000000
0!
0%
b100 *
0-
02
b100 6
#984090000000
1!
1%
1-
12
#984100000000
0!
0%
b101 *
0-
02
b101 6
#984110000000
1!
1%
1-
12
#984120000000
0!
0%
b110 *
0-
02
b110 6
#984130000000
1!
1%
1-
12
#984140000000
0!
0%
b111 *
0-
02
b111 6
#984150000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#984160000000
0!
0%
b0 *
0-
02
b0 6
#984170000000
1!
1%
1-
12
#984180000000
0!
0%
b1 *
0-
02
b1 6
#984190000000
1!
1%
1-
12
#984200000000
0!
0%
b10 *
0-
02
b10 6
#984210000000
1!
1%
1-
12
#984220000000
0!
0%
b11 *
0-
02
b11 6
#984230000000
1!
1%
1-
12
15
#984240000000
0!
0%
b100 *
0-
02
b100 6
#984250000000
1!
1%
1-
12
#984260000000
0!
0%
b101 *
0-
02
b101 6
#984270000000
1!
1%
1-
12
#984280000000
0!
0%
b110 *
0-
02
b110 6
#984290000000
1!
1%
1-
12
#984300000000
0!
0%
b111 *
0-
02
b111 6
#984310000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#984320000000
0!
0%
b0 *
0-
02
b0 6
#984330000000
1!
1%
1-
12
#984340000000
0!
0%
b1 *
0-
02
b1 6
#984350000000
1!
1%
1-
12
#984360000000
0!
0%
b10 *
0-
02
b10 6
#984370000000
1!
1%
1-
12
#984380000000
0!
0%
b11 *
0-
02
b11 6
#984390000000
1!
1%
1-
12
15
#984400000000
0!
0%
b100 *
0-
02
b100 6
#984410000000
1!
1%
1-
12
#984420000000
0!
0%
b101 *
0-
02
b101 6
#984430000000
1!
1%
1-
12
#984440000000
0!
0%
b110 *
0-
02
b110 6
#984450000000
1!
1%
1-
12
#984460000000
0!
0%
b111 *
0-
02
b111 6
#984470000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#984480000000
0!
0%
b0 *
0-
02
b0 6
#984490000000
1!
1%
1-
12
#984500000000
0!
0%
b1 *
0-
02
b1 6
#984510000000
1!
1%
1-
12
#984520000000
0!
0%
b10 *
0-
02
b10 6
#984530000000
1!
1%
1-
12
#984540000000
0!
0%
b11 *
0-
02
b11 6
#984550000000
1!
1%
1-
12
15
#984560000000
0!
0%
b100 *
0-
02
b100 6
#984570000000
1!
1%
1-
12
#984580000000
0!
0%
b101 *
0-
02
b101 6
#984590000000
1!
1%
1-
12
#984600000000
0!
0%
b110 *
0-
02
b110 6
#984610000000
1!
1%
1-
12
#984620000000
0!
0%
b111 *
0-
02
b111 6
#984630000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#984640000000
0!
0%
b0 *
0-
02
b0 6
#984650000000
1!
1%
1-
12
#984660000000
0!
0%
b1 *
0-
02
b1 6
#984670000000
1!
1%
1-
12
#984680000000
0!
0%
b10 *
0-
02
b10 6
#984690000000
1!
1%
1-
12
#984700000000
0!
0%
b11 *
0-
02
b11 6
#984710000000
1!
1%
1-
12
15
#984720000000
0!
0%
b100 *
0-
02
b100 6
#984730000000
1!
1%
1-
12
#984740000000
0!
0%
b101 *
0-
02
b101 6
#984750000000
1!
1%
1-
12
#984760000000
0!
0%
b110 *
0-
02
b110 6
#984770000000
1!
1%
1-
12
#984780000000
0!
0%
b111 *
0-
02
b111 6
#984790000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#984800000000
0!
0%
b0 *
0-
02
b0 6
#984810000000
1!
1%
1-
12
#984820000000
0!
0%
b1 *
0-
02
b1 6
#984830000000
1!
1%
1-
12
#984840000000
0!
0%
b10 *
0-
02
b10 6
#984850000000
1!
1%
1-
12
#984860000000
0!
0%
b11 *
0-
02
b11 6
#984870000000
1!
1%
1-
12
15
#984880000000
0!
0%
b100 *
0-
02
b100 6
#984890000000
1!
1%
1-
12
#984900000000
0!
0%
b101 *
0-
02
b101 6
#984910000000
1!
1%
1-
12
#984920000000
0!
0%
b110 *
0-
02
b110 6
#984930000000
1!
1%
1-
12
#984940000000
0!
0%
b111 *
0-
02
b111 6
#984950000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#984960000000
0!
0%
b0 *
0-
02
b0 6
#984970000000
1!
1%
1-
12
#984980000000
0!
0%
b1 *
0-
02
b1 6
#984990000000
1!
1%
1-
12
#985000000000
0!
0%
b10 *
0-
02
b10 6
#985010000000
1!
1%
1-
12
#985020000000
0!
0%
b11 *
0-
02
b11 6
#985030000000
1!
1%
1-
12
15
#985040000000
0!
0%
b100 *
0-
02
b100 6
#985050000000
1!
1%
1-
12
#985060000000
0!
0%
b101 *
0-
02
b101 6
#985070000000
1!
1%
1-
12
#985080000000
0!
0%
b110 *
0-
02
b110 6
#985090000000
1!
1%
1-
12
#985100000000
0!
0%
b111 *
0-
02
b111 6
#985110000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#985120000000
0!
0%
b0 *
0-
02
b0 6
#985130000000
1!
1%
1-
12
#985140000000
0!
0%
b1 *
0-
02
b1 6
#985150000000
1!
1%
1-
12
#985160000000
0!
0%
b10 *
0-
02
b10 6
#985170000000
1!
1%
1-
12
#985180000000
0!
0%
b11 *
0-
02
b11 6
#985190000000
1!
1%
1-
12
15
#985200000000
0!
0%
b100 *
0-
02
b100 6
#985210000000
1!
1%
1-
12
#985220000000
0!
0%
b101 *
0-
02
b101 6
#985230000000
1!
1%
1-
12
#985240000000
0!
0%
b110 *
0-
02
b110 6
#985250000000
1!
1%
1-
12
#985260000000
0!
0%
b111 *
0-
02
b111 6
#985270000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#985280000000
0!
0%
b0 *
0-
02
b0 6
#985290000000
1!
1%
1-
12
#985300000000
0!
0%
b1 *
0-
02
b1 6
#985310000000
1!
1%
1-
12
#985320000000
0!
0%
b10 *
0-
02
b10 6
#985330000000
1!
1%
1-
12
#985340000000
0!
0%
b11 *
0-
02
b11 6
#985350000000
1!
1%
1-
12
15
#985360000000
0!
0%
b100 *
0-
02
b100 6
#985370000000
1!
1%
1-
12
#985380000000
0!
0%
b101 *
0-
02
b101 6
#985390000000
1!
1%
1-
12
#985400000000
0!
0%
b110 *
0-
02
b110 6
#985410000000
1!
1%
1-
12
#985420000000
0!
0%
b111 *
0-
02
b111 6
#985430000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#985440000000
0!
0%
b0 *
0-
02
b0 6
#985450000000
1!
1%
1-
12
#985460000000
0!
0%
b1 *
0-
02
b1 6
#985470000000
1!
1%
1-
12
#985480000000
0!
0%
b10 *
0-
02
b10 6
#985490000000
1!
1%
1-
12
#985500000000
0!
0%
b11 *
0-
02
b11 6
#985510000000
1!
1%
1-
12
15
#985520000000
0!
0%
b100 *
0-
02
b100 6
#985530000000
1!
1%
1-
12
#985540000000
0!
0%
b101 *
0-
02
b101 6
#985550000000
1!
1%
1-
12
#985560000000
0!
0%
b110 *
0-
02
b110 6
#985570000000
1!
1%
1-
12
#985580000000
0!
0%
b111 *
0-
02
b111 6
#985590000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#985600000000
0!
0%
b0 *
0-
02
b0 6
#985610000000
1!
1%
1-
12
#985620000000
0!
0%
b1 *
0-
02
b1 6
#985630000000
1!
1%
1-
12
#985640000000
0!
0%
b10 *
0-
02
b10 6
#985650000000
1!
1%
1-
12
#985660000000
0!
0%
b11 *
0-
02
b11 6
#985670000000
1!
1%
1-
12
15
#985680000000
0!
0%
b100 *
0-
02
b100 6
#985690000000
1!
1%
1-
12
#985700000000
0!
0%
b101 *
0-
02
b101 6
#985710000000
1!
1%
1-
12
#985720000000
0!
0%
b110 *
0-
02
b110 6
#985730000000
1!
1%
1-
12
#985740000000
0!
0%
b111 *
0-
02
b111 6
#985750000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#985760000000
0!
0%
b0 *
0-
02
b0 6
#985770000000
1!
1%
1-
12
#985780000000
0!
0%
b1 *
0-
02
b1 6
#985790000000
1!
1%
1-
12
#985800000000
0!
0%
b10 *
0-
02
b10 6
#985810000000
1!
1%
1-
12
#985820000000
0!
0%
b11 *
0-
02
b11 6
#985830000000
1!
1%
1-
12
15
#985840000000
0!
0%
b100 *
0-
02
b100 6
#985850000000
1!
1%
1-
12
#985860000000
0!
0%
b101 *
0-
02
b101 6
#985870000000
1!
1%
1-
12
#985880000000
0!
0%
b110 *
0-
02
b110 6
#985890000000
1!
1%
1-
12
#985900000000
0!
0%
b111 *
0-
02
b111 6
#985910000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#985920000000
0!
0%
b0 *
0-
02
b0 6
#985930000000
1!
1%
1-
12
#985940000000
0!
0%
b1 *
0-
02
b1 6
#985950000000
1!
1%
1-
12
#985960000000
0!
0%
b10 *
0-
02
b10 6
#985970000000
1!
1%
1-
12
#985980000000
0!
0%
b11 *
0-
02
b11 6
#985990000000
1!
1%
1-
12
15
#986000000000
0!
0%
b100 *
0-
02
b100 6
#986010000000
1!
1%
1-
12
#986020000000
0!
0%
b101 *
0-
02
b101 6
#986030000000
1!
1%
1-
12
#986040000000
0!
0%
b110 *
0-
02
b110 6
#986050000000
1!
1%
1-
12
#986060000000
0!
0%
b111 *
0-
02
b111 6
#986070000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#986080000000
0!
0%
b0 *
0-
02
b0 6
#986090000000
1!
1%
1-
12
#986100000000
0!
0%
b1 *
0-
02
b1 6
#986110000000
1!
1%
1-
12
#986120000000
0!
0%
b10 *
0-
02
b10 6
#986130000000
1!
1%
1-
12
#986140000000
0!
0%
b11 *
0-
02
b11 6
#986150000000
1!
1%
1-
12
15
#986160000000
0!
0%
b100 *
0-
02
b100 6
#986170000000
1!
1%
1-
12
#986180000000
0!
0%
b101 *
0-
02
b101 6
#986190000000
1!
1%
1-
12
#986200000000
0!
0%
b110 *
0-
02
b110 6
#986210000000
1!
1%
1-
12
#986220000000
0!
0%
b111 *
0-
02
b111 6
#986230000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#986240000000
0!
0%
b0 *
0-
02
b0 6
#986250000000
1!
1%
1-
12
#986260000000
0!
0%
b1 *
0-
02
b1 6
#986270000000
1!
1%
1-
12
#986280000000
0!
0%
b10 *
0-
02
b10 6
#986290000000
1!
1%
1-
12
#986300000000
0!
0%
b11 *
0-
02
b11 6
#986310000000
1!
1%
1-
12
15
#986320000000
0!
0%
b100 *
0-
02
b100 6
#986330000000
1!
1%
1-
12
#986340000000
0!
0%
b101 *
0-
02
b101 6
#986350000000
1!
1%
1-
12
#986360000000
0!
0%
b110 *
0-
02
b110 6
#986370000000
1!
1%
1-
12
#986380000000
0!
0%
b111 *
0-
02
b111 6
#986390000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#986400000000
0!
0%
b0 *
0-
02
b0 6
#986410000000
1!
1%
1-
12
#986420000000
0!
0%
b1 *
0-
02
b1 6
#986430000000
1!
1%
1-
12
#986440000000
0!
0%
b10 *
0-
02
b10 6
#986450000000
1!
1%
1-
12
#986460000000
0!
0%
b11 *
0-
02
b11 6
#986470000000
1!
1%
1-
12
15
#986480000000
0!
0%
b100 *
0-
02
b100 6
#986490000000
1!
1%
1-
12
#986500000000
0!
0%
b101 *
0-
02
b101 6
#986510000000
1!
1%
1-
12
#986520000000
0!
0%
b110 *
0-
02
b110 6
#986530000000
1!
1%
1-
12
#986540000000
0!
0%
b111 *
0-
02
b111 6
#986550000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#986560000000
0!
0%
b0 *
0-
02
b0 6
#986570000000
1!
1%
1-
12
#986580000000
0!
0%
b1 *
0-
02
b1 6
#986590000000
1!
1%
1-
12
#986600000000
0!
0%
b10 *
0-
02
b10 6
#986610000000
1!
1%
1-
12
#986620000000
0!
0%
b11 *
0-
02
b11 6
#986630000000
1!
1%
1-
12
15
#986640000000
0!
0%
b100 *
0-
02
b100 6
#986650000000
1!
1%
1-
12
#986660000000
0!
0%
b101 *
0-
02
b101 6
#986670000000
1!
1%
1-
12
#986680000000
0!
0%
b110 *
0-
02
b110 6
#986690000000
1!
1%
1-
12
#986700000000
0!
0%
b111 *
0-
02
b111 6
#986710000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#986720000000
0!
0%
b0 *
0-
02
b0 6
#986730000000
1!
1%
1-
12
#986740000000
0!
0%
b1 *
0-
02
b1 6
#986750000000
1!
1%
1-
12
#986760000000
0!
0%
b10 *
0-
02
b10 6
#986770000000
1!
1%
1-
12
#986780000000
0!
0%
b11 *
0-
02
b11 6
#986790000000
1!
1%
1-
12
15
#986800000000
0!
0%
b100 *
0-
02
b100 6
#986810000000
1!
1%
1-
12
#986820000000
0!
0%
b101 *
0-
02
b101 6
#986830000000
1!
1%
1-
12
#986840000000
0!
0%
b110 *
0-
02
b110 6
#986850000000
1!
1%
1-
12
#986860000000
0!
0%
b111 *
0-
02
b111 6
#986870000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#986880000000
0!
0%
b0 *
0-
02
b0 6
#986890000000
1!
1%
1-
12
#986900000000
0!
0%
b1 *
0-
02
b1 6
#986910000000
1!
1%
1-
12
#986920000000
0!
0%
b10 *
0-
02
b10 6
#986930000000
1!
1%
1-
12
#986940000000
0!
0%
b11 *
0-
02
b11 6
#986950000000
1!
1%
1-
12
15
#986960000000
0!
0%
b100 *
0-
02
b100 6
#986970000000
1!
1%
1-
12
#986980000000
0!
0%
b101 *
0-
02
b101 6
#986990000000
1!
1%
1-
12
#987000000000
0!
0%
b110 *
0-
02
b110 6
#987010000000
1!
1%
1-
12
#987020000000
0!
0%
b111 *
0-
02
b111 6
#987030000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#987040000000
0!
0%
b0 *
0-
02
b0 6
#987050000000
1!
1%
1-
12
#987060000000
0!
0%
b1 *
0-
02
b1 6
#987070000000
1!
1%
1-
12
#987080000000
0!
0%
b10 *
0-
02
b10 6
#987090000000
1!
1%
1-
12
#987100000000
0!
0%
b11 *
0-
02
b11 6
#987110000000
1!
1%
1-
12
15
#987120000000
0!
0%
b100 *
0-
02
b100 6
#987130000000
1!
1%
1-
12
#987140000000
0!
0%
b101 *
0-
02
b101 6
#987150000000
1!
1%
1-
12
#987160000000
0!
0%
b110 *
0-
02
b110 6
#987170000000
1!
1%
1-
12
#987180000000
0!
0%
b111 *
0-
02
b111 6
#987190000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#987200000000
0!
0%
b0 *
0-
02
b0 6
#987210000000
1!
1%
1-
12
#987220000000
0!
0%
b1 *
0-
02
b1 6
#987230000000
1!
1%
1-
12
#987240000000
0!
0%
b10 *
0-
02
b10 6
#987250000000
1!
1%
1-
12
#987260000000
0!
0%
b11 *
0-
02
b11 6
#987270000000
1!
1%
1-
12
15
#987280000000
0!
0%
b100 *
0-
02
b100 6
#987290000000
1!
1%
1-
12
#987300000000
0!
0%
b101 *
0-
02
b101 6
#987310000000
1!
1%
1-
12
#987320000000
0!
0%
b110 *
0-
02
b110 6
#987330000000
1!
1%
1-
12
#987340000000
0!
0%
b111 *
0-
02
b111 6
#987350000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#987360000000
0!
0%
b0 *
0-
02
b0 6
#987370000000
1!
1%
1-
12
#987380000000
0!
0%
b1 *
0-
02
b1 6
#987390000000
1!
1%
1-
12
#987400000000
0!
0%
b10 *
0-
02
b10 6
#987410000000
1!
1%
1-
12
#987420000000
0!
0%
b11 *
0-
02
b11 6
#987430000000
1!
1%
1-
12
15
#987440000000
0!
0%
b100 *
0-
02
b100 6
#987450000000
1!
1%
1-
12
#987460000000
0!
0%
b101 *
0-
02
b101 6
#987470000000
1!
1%
1-
12
#987480000000
0!
0%
b110 *
0-
02
b110 6
#987490000000
1!
1%
1-
12
#987500000000
0!
0%
b111 *
0-
02
b111 6
#987510000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#987520000000
0!
0%
b0 *
0-
02
b0 6
#987530000000
1!
1%
1-
12
#987540000000
0!
0%
b1 *
0-
02
b1 6
#987550000000
1!
1%
1-
12
#987560000000
0!
0%
b10 *
0-
02
b10 6
#987570000000
1!
1%
1-
12
#987580000000
0!
0%
b11 *
0-
02
b11 6
#987590000000
1!
1%
1-
12
15
#987600000000
0!
0%
b100 *
0-
02
b100 6
#987610000000
1!
1%
1-
12
#987620000000
0!
0%
b101 *
0-
02
b101 6
#987630000000
1!
1%
1-
12
#987640000000
0!
0%
b110 *
0-
02
b110 6
#987650000000
1!
1%
1-
12
#987660000000
0!
0%
b111 *
0-
02
b111 6
#987670000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#987680000000
0!
0%
b0 *
0-
02
b0 6
#987690000000
1!
1%
1-
12
#987700000000
0!
0%
b1 *
0-
02
b1 6
#987710000000
1!
1%
1-
12
#987720000000
0!
0%
b10 *
0-
02
b10 6
#987730000000
1!
1%
1-
12
#987740000000
0!
0%
b11 *
0-
02
b11 6
#987750000000
1!
1%
1-
12
15
#987760000000
0!
0%
b100 *
0-
02
b100 6
#987770000000
1!
1%
1-
12
#987780000000
0!
0%
b101 *
0-
02
b101 6
#987790000000
1!
1%
1-
12
#987800000000
0!
0%
b110 *
0-
02
b110 6
#987810000000
1!
1%
1-
12
#987820000000
0!
0%
b111 *
0-
02
b111 6
#987830000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#987840000000
0!
0%
b0 *
0-
02
b0 6
#987850000000
1!
1%
1-
12
#987860000000
0!
0%
b1 *
0-
02
b1 6
#987870000000
1!
1%
1-
12
#987880000000
0!
0%
b10 *
0-
02
b10 6
#987890000000
1!
1%
1-
12
#987900000000
0!
0%
b11 *
0-
02
b11 6
#987910000000
1!
1%
1-
12
15
#987920000000
0!
0%
b100 *
0-
02
b100 6
#987930000000
1!
1%
1-
12
#987940000000
0!
0%
b101 *
0-
02
b101 6
#987950000000
1!
1%
1-
12
#987960000000
0!
0%
b110 *
0-
02
b110 6
#987970000000
1!
1%
1-
12
#987980000000
0!
0%
b111 *
0-
02
b111 6
#987990000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#988000000000
0!
0%
b0 *
0-
02
b0 6
#988010000000
1!
1%
1-
12
#988020000000
0!
0%
b1 *
0-
02
b1 6
#988030000000
1!
1%
1-
12
#988040000000
0!
0%
b10 *
0-
02
b10 6
#988050000000
1!
1%
1-
12
#988060000000
0!
0%
b11 *
0-
02
b11 6
#988070000000
1!
1%
1-
12
15
#988080000000
0!
0%
b100 *
0-
02
b100 6
#988090000000
1!
1%
1-
12
#988100000000
0!
0%
b101 *
0-
02
b101 6
#988110000000
1!
1%
1-
12
#988120000000
0!
0%
b110 *
0-
02
b110 6
#988130000000
1!
1%
1-
12
#988140000000
0!
0%
b111 *
0-
02
b111 6
#988150000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#988160000000
0!
0%
b0 *
0-
02
b0 6
#988170000000
1!
1%
1-
12
#988180000000
0!
0%
b1 *
0-
02
b1 6
#988190000000
1!
1%
1-
12
#988200000000
0!
0%
b10 *
0-
02
b10 6
#988210000000
1!
1%
1-
12
#988220000000
0!
0%
b11 *
0-
02
b11 6
#988230000000
1!
1%
1-
12
15
#988240000000
0!
0%
b100 *
0-
02
b100 6
#988250000000
1!
1%
1-
12
#988260000000
0!
0%
b101 *
0-
02
b101 6
#988270000000
1!
1%
1-
12
#988280000000
0!
0%
b110 *
0-
02
b110 6
#988290000000
1!
1%
1-
12
#988300000000
0!
0%
b111 *
0-
02
b111 6
#988310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#988320000000
0!
0%
b0 *
0-
02
b0 6
#988330000000
1!
1%
1-
12
#988340000000
0!
0%
b1 *
0-
02
b1 6
#988350000000
1!
1%
1-
12
#988360000000
0!
0%
b10 *
0-
02
b10 6
#988370000000
1!
1%
1-
12
#988380000000
0!
0%
b11 *
0-
02
b11 6
#988390000000
1!
1%
1-
12
15
#988400000000
0!
0%
b100 *
0-
02
b100 6
#988410000000
1!
1%
1-
12
#988420000000
0!
0%
b101 *
0-
02
b101 6
#988430000000
1!
1%
1-
12
#988440000000
0!
0%
b110 *
0-
02
b110 6
#988450000000
1!
1%
1-
12
#988460000000
0!
0%
b111 *
0-
02
b111 6
#988470000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#988480000000
0!
0%
b0 *
0-
02
b0 6
#988490000000
1!
1%
1-
12
#988500000000
0!
0%
b1 *
0-
02
b1 6
#988510000000
1!
1%
1-
12
#988520000000
0!
0%
b10 *
0-
02
b10 6
#988530000000
1!
1%
1-
12
#988540000000
0!
0%
b11 *
0-
02
b11 6
#988550000000
1!
1%
1-
12
15
#988560000000
0!
0%
b100 *
0-
02
b100 6
#988570000000
1!
1%
1-
12
#988580000000
0!
0%
b101 *
0-
02
b101 6
#988590000000
1!
1%
1-
12
#988600000000
0!
0%
b110 *
0-
02
b110 6
#988610000000
1!
1%
1-
12
#988620000000
0!
0%
b111 *
0-
02
b111 6
#988630000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#988640000000
0!
0%
b0 *
0-
02
b0 6
#988650000000
1!
1%
1-
12
#988660000000
0!
0%
b1 *
0-
02
b1 6
#988670000000
1!
1%
1-
12
#988680000000
0!
0%
b10 *
0-
02
b10 6
#988690000000
1!
1%
1-
12
#988700000000
0!
0%
b11 *
0-
02
b11 6
#988710000000
1!
1%
1-
12
15
#988720000000
0!
0%
b100 *
0-
02
b100 6
#988730000000
1!
1%
1-
12
#988740000000
0!
0%
b101 *
0-
02
b101 6
#988750000000
1!
1%
1-
12
#988760000000
0!
0%
b110 *
0-
02
b110 6
#988770000000
1!
1%
1-
12
#988780000000
0!
0%
b111 *
0-
02
b111 6
#988790000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#988800000000
0!
0%
b0 *
0-
02
b0 6
#988810000000
1!
1%
1-
12
#988820000000
0!
0%
b1 *
0-
02
b1 6
#988830000000
1!
1%
1-
12
#988840000000
0!
0%
b10 *
0-
02
b10 6
#988850000000
1!
1%
1-
12
#988860000000
0!
0%
b11 *
0-
02
b11 6
#988870000000
1!
1%
1-
12
15
#988880000000
0!
0%
b100 *
0-
02
b100 6
#988890000000
1!
1%
1-
12
#988900000000
0!
0%
b101 *
0-
02
b101 6
#988910000000
1!
1%
1-
12
#988920000000
0!
0%
b110 *
0-
02
b110 6
#988930000000
1!
1%
1-
12
#988940000000
0!
0%
b111 *
0-
02
b111 6
#988950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#988960000000
0!
0%
b0 *
0-
02
b0 6
#988970000000
1!
1%
1-
12
#988980000000
0!
0%
b1 *
0-
02
b1 6
#988990000000
1!
1%
1-
12
#989000000000
0!
0%
b10 *
0-
02
b10 6
#989010000000
1!
1%
1-
12
#989020000000
0!
0%
b11 *
0-
02
b11 6
#989030000000
1!
1%
1-
12
15
#989040000000
0!
0%
b100 *
0-
02
b100 6
#989050000000
1!
1%
1-
12
#989060000000
0!
0%
b101 *
0-
02
b101 6
#989070000000
1!
1%
1-
12
#989080000000
0!
0%
b110 *
0-
02
b110 6
#989090000000
1!
1%
1-
12
#989100000000
0!
0%
b111 *
0-
02
b111 6
#989110000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#989120000000
0!
0%
b0 *
0-
02
b0 6
#989130000000
1!
1%
1-
12
#989140000000
0!
0%
b1 *
0-
02
b1 6
#989150000000
1!
1%
1-
12
#989160000000
0!
0%
b10 *
0-
02
b10 6
#989170000000
1!
1%
1-
12
#989180000000
0!
0%
b11 *
0-
02
b11 6
#989190000000
1!
1%
1-
12
15
#989200000000
0!
0%
b100 *
0-
02
b100 6
#989210000000
1!
1%
1-
12
#989220000000
0!
0%
b101 *
0-
02
b101 6
#989230000000
1!
1%
1-
12
#989240000000
0!
0%
b110 *
0-
02
b110 6
#989250000000
1!
1%
1-
12
#989260000000
0!
0%
b111 *
0-
02
b111 6
#989270000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#989280000000
0!
0%
b0 *
0-
02
b0 6
#989290000000
1!
1%
1-
12
#989300000000
0!
0%
b1 *
0-
02
b1 6
#989310000000
1!
1%
1-
12
#989320000000
0!
0%
b10 *
0-
02
b10 6
#989330000000
1!
1%
1-
12
#989340000000
0!
0%
b11 *
0-
02
b11 6
#989350000000
1!
1%
1-
12
15
#989360000000
0!
0%
b100 *
0-
02
b100 6
#989370000000
1!
1%
1-
12
#989380000000
0!
0%
b101 *
0-
02
b101 6
#989390000000
1!
1%
1-
12
#989400000000
0!
0%
b110 *
0-
02
b110 6
#989410000000
1!
1%
1-
12
#989420000000
0!
0%
b111 *
0-
02
b111 6
#989430000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#989440000000
0!
0%
b0 *
0-
02
b0 6
#989450000000
1!
1%
1-
12
#989460000000
0!
0%
b1 *
0-
02
b1 6
#989470000000
1!
1%
1-
12
#989480000000
0!
0%
b10 *
0-
02
b10 6
#989490000000
1!
1%
1-
12
#989500000000
0!
0%
b11 *
0-
02
b11 6
#989510000000
1!
1%
1-
12
15
#989520000000
0!
0%
b100 *
0-
02
b100 6
#989530000000
1!
1%
1-
12
#989540000000
0!
0%
b101 *
0-
02
b101 6
#989550000000
1!
1%
1-
12
#989560000000
0!
0%
b110 *
0-
02
b110 6
#989570000000
1!
1%
1-
12
#989580000000
0!
0%
b111 *
0-
02
b111 6
#989590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#989600000000
0!
0%
b0 *
0-
02
b0 6
#989610000000
1!
1%
1-
12
#989620000000
0!
0%
b1 *
0-
02
b1 6
#989630000000
1!
1%
1-
12
#989640000000
0!
0%
b10 *
0-
02
b10 6
#989650000000
1!
1%
1-
12
#989660000000
0!
0%
b11 *
0-
02
b11 6
#989670000000
1!
1%
1-
12
15
#989680000000
0!
0%
b100 *
0-
02
b100 6
#989690000000
1!
1%
1-
12
#989700000000
0!
0%
b101 *
0-
02
b101 6
#989710000000
1!
1%
1-
12
#989720000000
0!
0%
b110 *
0-
02
b110 6
#989730000000
1!
1%
1-
12
#989740000000
0!
0%
b111 *
0-
02
b111 6
#989750000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#989760000000
0!
0%
b0 *
0-
02
b0 6
#989770000000
1!
1%
1-
12
#989780000000
0!
0%
b1 *
0-
02
b1 6
#989790000000
1!
1%
1-
12
#989800000000
0!
0%
b10 *
0-
02
b10 6
#989810000000
1!
1%
1-
12
#989820000000
0!
0%
b11 *
0-
02
b11 6
#989830000000
1!
1%
1-
12
15
#989840000000
0!
0%
b100 *
0-
02
b100 6
#989850000000
1!
1%
1-
12
#989860000000
0!
0%
b101 *
0-
02
b101 6
#989870000000
1!
1%
1-
12
#989880000000
0!
0%
b110 *
0-
02
b110 6
#989890000000
1!
1%
1-
12
#989900000000
0!
0%
b111 *
0-
02
b111 6
#989910000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#989920000000
0!
0%
b0 *
0-
02
b0 6
#989930000000
1!
1%
1-
12
#989940000000
0!
0%
b1 *
0-
02
b1 6
#989950000000
1!
1%
1-
12
#989960000000
0!
0%
b10 *
0-
02
b10 6
#989970000000
1!
1%
1-
12
#989980000000
0!
0%
b11 *
0-
02
b11 6
#989990000000
1!
1%
1-
12
15
#990000000000
0!
0%
b100 *
0-
02
b100 6
#990010000000
1!
1%
1-
12
#990020000000
0!
0%
b101 *
0-
02
b101 6
#990030000000
1!
1%
1-
12
#990040000000
0!
0%
b110 *
0-
02
b110 6
#990050000000
1!
1%
1-
12
#990060000000
0!
0%
b111 *
0-
02
b111 6
#990070000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#990080000000
0!
0%
b0 *
0-
02
b0 6
#990090000000
1!
1%
1-
12
#990100000000
0!
0%
b1 *
0-
02
b1 6
#990110000000
1!
1%
1-
12
#990120000000
0!
0%
b10 *
0-
02
b10 6
#990130000000
1!
1%
1-
12
#990140000000
0!
0%
b11 *
0-
02
b11 6
#990150000000
1!
1%
1-
12
15
#990160000000
0!
0%
b100 *
0-
02
b100 6
#990170000000
1!
1%
1-
12
#990180000000
0!
0%
b101 *
0-
02
b101 6
#990190000000
1!
1%
1-
12
#990200000000
0!
0%
b110 *
0-
02
b110 6
#990210000000
1!
1%
1-
12
#990220000000
0!
0%
b111 *
0-
02
b111 6
#990230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#990240000000
0!
0%
b0 *
0-
02
b0 6
#990250000000
1!
1%
1-
12
#990260000000
0!
0%
b1 *
0-
02
b1 6
#990270000000
1!
1%
1-
12
#990280000000
0!
0%
b10 *
0-
02
b10 6
#990290000000
1!
1%
1-
12
#990300000000
0!
0%
b11 *
0-
02
b11 6
#990310000000
1!
1%
1-
12
15
#990320000000
0!
0%
b100 *
0-
02
b100 6
#990330000000
1!
1%
1-
12
#990340000000
0!
0%
b101 *
0-
02
b101 6
#990350000000
1!
1%
1-
12
#990360000000
0!
0%
b110 *
0-
02
b110 6
#990370000000
1!
1%
1-
12
#990380000000
0!
0%
b111 *
0-
02
b111 6
#990390000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#990400000000
0!
0%
b0 *
0-
02
b0 6
#990410000000
1!
1%
1-
12
#990420000000
0!
0%
b1 *
0-
02
b1 6
#990430000000
1!
1%
1-
12
#990440000000
0!
0%
b10 *
0-
02
b10 6
#990450000000
1!
1%
1-
12
#990460000000
0!
0%
b11 *
0-
02
b11 6
#990470000000
1!
1%
1-
12
15
#990480000000
0!
0%
b100 *
0-
02
b100 6
#990490000000
1!
1%
1-
12
#990500000000
0!
0%
b101 *
0-
02
b101 6
#990510000000
1!
1%
1-
12
#990520000000
0!
0%
b110 *
0-
02
b110 6
#990530000000
1!
1%
1-
12
#990540000000
0!
0%
b111 *
0-
02
b111 6
#990550000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#990560000000
0!
0%
b0 *
0-
02
b0 6
#990570000000
1!
1%
1-
12
#990580000000
0!
0%
b1 *
0-
02
b1 6
#990590000000
1!
1%
1-
12
#990600000000
0!
0%
b10 *
0-
02
b10 6
#990610000000
1!
1%
1-
12
#990620000000
0!
0%
b11 *
0-
02
b11 6
#990630000000
1!
1%
1-
12
15
#990640000000
0!
0%
b100 *
0-
02
b100 6
#990650000000
1!
1%
1-
12
#990660000000
0!
0%
b101 *
0-
02
b101 6
#990670000000
1!
1%
1-
12
#990680000000
0!
0%
b110 *
0-
02
b110 6
#990690000000
1!
1%
1-
12
#990700000000
0!
0%
b111 *
0-
02
b111 6
#990710000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#990720000000
0!
0%
b0 *
0-
02
b0 6
#990730000000
1!
1%
1-
12
#990740000000
0!
0%
b1 *
0-
02
b1 6
#990750000000
1!
1%
1-
12
#990760000000
0!
0%
b10 *
0-
02
b10 6
#990770000000
1!
1%
1-
12
#990780000000
0!
0%
b11 *
0-
02
b11 6
#990790000000
1!
1%
1-
12
15
#990800000000
0!
0%
b100 *
0-
02
b100 6
#990810000000
1!
1%
1-
12
#990820000000
0!
0%
b101 *
0-
02
b101 6
#990830000000
1!
1%
1-
12
#990840000000
0!
0%
b110 *
0-
02
b110 6
#990850000000
1!
1%
1-
12
#990860000000
0!
0%
b111 *
0-
02
b111 6
#990870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#990880000000
0!
0%
b0 *
0-
02
b0 6
#990890000000
1!
1%
1-
12
#990900000000
0!
0%
b1 *
0-
02
b1 6
#990910000000
1!
1%
1-
12
#990920000000
0!
0%
b10 *
0-
02
b10 6
#990930000000
1!
1%
1-
12
#990940000000
0!
0%
b11 *
0-
02
b11 6
#990950000000
1!
1%
1-
12
15
#990960000000
0!
0%
b100 *
0-
02
b100 6
#990970000000
1!
1%
1-
12
#990980000000
0!
0%
b101 *
0-
02
b101 6
#990990000000
1!
1%
1-
12
#991000000000
0!
0%
b110 *
0-
02
b110 6
#991010000000
1!
1%
1-
12
#991020000000
0!
0%
b111 *
0-
02
b111 6
#991030000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#991040000000
0!
0%
b0 *
0-
02
b0 6
#991050000000
1!
1%
1-
12
#991060000000
0!
0%
b1 *
0-
02
b1 6
#991070000000
1!
1%
1-
12
#991080000000
0!
0%
b10 *
0-
02
b10 6
#991090000000
1!
1%
1-
12
#991100000000
0!
0%
b11 *
0-
02
b11 6
#991110000000
1!
1%
1-
12
15
#991120000000
0!
0%
b100 *
0-
02
b100 6
#991130000000
1!
1%
1-
12
#991140000000
0!
0%
b101 *
0-
02
b101 6
#991150000000
1!
1%
1-
12
#991160000000
0!
0%
b110 *
0-
02
b110 6
#991170000000
1!
1%
1-
12
#991180000000
0!
0%
b111 *
0-
02
b111 6
#991190000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#991200000000
0!
0%
b0 *
0-
02
b0 6
#991210000000
1!
1%
1-
12
#991220000000
0!
0%
b1 *
0-
02
b1 6
#991230000000
1!
1%
1-
12
#991240000000
0!
0%
b10 *
0-
02
b10 6
#991250000000
1!
1%
1-
12
#991260000000
0!
0%
b11 *
0-
02
b11 6
#991270000000
1!
1%
1-
12
15
#991280000000
0!
0%
b100 *
0-
02
b100 6
#991290000000
1!
1%
1-
12
#991300000000
0!
0%
b101 *
0-
02
b101 6
#991310000000
1!
1%
1-
12
#991320000000
0!
0%
b110 *
0-
02
b110 6
#991330000000
1!
1%
1-
12
#991340000000
0!
0%
b111 *
0-
02
b111 6
#991350000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#991360000000
0!
0%
b0 *
0-
02
b0 6
#991370000000
1!
1%
1-
12
#991380000000
0!
0%
b1 *
0-
02
b1 6
#991390000000
1!
1%
1-
12
#991400000000
0!
0%
b10 *
0-
02
b10 6
#991410000000
1!
1%
1-
12
#991420000000
0!
0%
b11 *
0-
02
b11 6
#991430000000
1!
1%
1-
12
15
#991440000000
0!
0%
b100 *
0-
02
b100 6
#991450000000
1!
1%
1-
12
#991460000000
0!
0%
b101 *
0-
02
b101 6
#991470000000
1!
1%
1-
12
#991480000000
0!
0%
b110 *
0-
02
b110 6
#991490000000
1!
1%
1-
12
#991500000000
0!
0%
b111 *
0-
02
b111 6
#991510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#991520000000
0!
0%
b0 *
0-
02
b0 6
#991530000000
1!
1%
1-
12
#991540000000
0!
0%
b1 *
0-
02
b1 6
#991550000000
1!
1%
1-
12
#991560000000
0!
0%
b10 *
0-
02
b10 6
#991570000000
1!
1%
1-
12
#991580000000
0!
0%
b11 *
0-
02
b11 6
#991590000000
1!
1%
1-
12
15
#991600000000
0!
0%
b100 *
0-
02
b100 6
#991610000000
1!
1%
1-
12
#991620000000
0!
0%
b101 *
0-
02
b101 6
#991630000000
1!
1%
1-
12
#991640000000
0!
0%
b110 *
0-
02
b110 6
#991650000000
1!
1%
1-
12
#991660000000
0!
0%
b111 *
0-
02
b111 6
#991670000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#991680000000
0!
0%
b0 *
0-
02
b0 6
#991690000000
1!
1%
1-
12
#991700000000
0!
0%
b1 *
0-
02
b1 6
#991710000000
1!
1%
1-
12
#991720000000
0!
0%
b10 *
0-
02
b10 6
#991730000000
1!
1%
1-
12
#991740000000
0!
0%
b11 *
0-
02
b11 6
#991750000000
1!
1%
1-
12
15
#991760000000
0!
0%
b100 *
0-
02
b100 6
#991770000000
1!
1%
1-
12
#991780000000
0!
0%
b101 *
0-
02
b101 6
#991790000000
1!
1%
1-
12
#991800000000
0!
0%
b110 *
0-
02
b110 6
#991810000000
1!
1%
1-
12
#991820000000
0!
0%
b111 *
0-
02
b111 6
#991830000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#991840000000
0!
0%
b0 *
0-
02
b0 6
#991850000000
1!
1%
1-
12
#991860000000
0!
0%
b1 *
0-
02
b1 6
#991870000000
1!
1%
1-
12
#991880000000
0!
0%
b10 *
0-
02
b10 6
#991890000000
1!
1%
1-
12
#991900000000
0!
0%
b11 *
0-
02
b11 6
#991910000000
1!
1%
1-
12
15
#991920000000
0!
0%
b100 *
0-
02
b100 6
#991930000000
1!
1%
1-
12
#991940000000
0!
0%
b101 *
0-
02
b101 6
#991950000000
1!
1%
1-
12
#991960000000
0!
0%
b110 *
0-
02
b110 6
#991970000000
1!
1%
1-
12
#991980000000
0!
0%
b111 *
0-
02
b111 6
#991990000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#992000000000
0!
0%
b0 *
0-
02
b0 6
#992010000000
1!
1%
1-
12
#992020000000
0!
0%
b1 *
0-
02
b1 6
#992030000000
1!
1%
1-
12
#992040000000
0!
0%
b10 *
0-
02
b10 6
#992050000000
1!
1%
1-
12
#992060000000
0!
0%
b11 *
0-
02
b11 6
#992070000000
1!
1%
1-
12
15
#992080000000
0!
0%
b100 *
0-
02
b100 6
#992090000000
1!
1%
1-
12
#992100000000
0!
0%
b101 *
0-
02
b101 6
#992110000000
1!
1%
1-
12
#992120000000
0!
0%
b110 *
0-
02
b110 6
#992130000000
1!
1%
1-
12
#992140000000
0!
0%
b111 *
0-
02
b111 6
#992150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#992160000000
0!
0%
b0 *
0-
02
b0 6
#992170000000
1!
1%
1-
12
#992180000000
0!
0%
b1 *
0-
02
b1 6
#992190000000
1!
1%
1-
12
#992200000000
0!
0%
b10 *
0-
02
b10 6
#992210000000
1!
1%
1-
12
#992220000000
0!
0%
b11 *
0-
02
b11 6
#992230000000
1!
1%
1-
12
15
#992240000000
0!
0%
b100 *
0-
02
b100 6
#992250000000
1!
1%
1-
12
#992260000000
0!
0%
b101 *
0-
02
b101 6
#992270000000
1!
1%
1-
12
#992280000000
0!
0%
b110 *
0-
02
b110 6
#992290000000
1!
1%
1-
12
#992300000000
0!
0%
b111 *
0-
02
b111 6
#992310000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#992320000000
0!
0%
b0 *
0-
02
b0 6
#992330000000
1!
1%
1-
12
#992340000000
0!
0%
b1 *
0-
02
b1 6
#992350000000
1!
1%
1-
12
#992360000000
0!
0%
b10 *
0-
02
b10 6
#992370000000
1!
1%
1-
12
#992380000000
0!
0%
b11 *
0-
02
b11 6
#992390000000
1!
1%
1-
12
15
#992400000000
0!
0%
b100 *
0-
02
b100 6
#992410000000
1!
1%
1-
12
#992420000000
0!
0%
b101 *
0-
02
b101 6
#992430000000
1!
1%
1-
12
#992440000000
0!
0%
b110 *
0-
02
b110 6
#992450000000
1!
1%
1-
12
#992460000000
0!
0%
b111 *
0-
02
b111 6
#992470000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#992480000000
0!
0%
b0 *
0-
02
b0 6
#992490000000
1!
1%
1-
12
#992500000000
0!
0%
b1 *
0-
02
b1 6
#992510000000
1!
1%
1-
12
#992520000000
0!
0%
b10 *
0-
02
b10 6
#992530000000
1!
1%
1-
12
#992540000000
0!
0%
b11 *
0-
02
b11 6
#992550000000
1!
1%
1-
12
15
#992560000000
0!
0%
b100 *
0-
02
b100 6
#992570000000
1!
1%
1-
12
#992580000000
0!
0%
b101 *
0-
02
b101 6
#992590000000
1!
1%
1-
12
#992600000000
0!
0%
b110 *
0-
02
b110 6
#992610000000
1!
1%
1-
12
#992620000000
0!
0%
b111 *
0-
02
b111 6
#992630000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#992640000000
0!
0%
b0 *
0-
02
b0 6
#992650000000
1!
1%
1-
12
#992660000000
0!
0%
b1 *
0-
02
b1 6
#992670000000
1!
1%
1-
12
#992680000000
0!
0%
b10 *
0-
02
b10 6
#992690000000
1!
1%
1-
12
#992700000000
0!
0%
b11 *
0-
02
b11 6
#992710000000
1!
1%
1-
12
15
#992720000000
0!
0%
b100 *
0-
02
b100 6
#992730000000
1!
1%
1-
12
#992740000000
0!
0%
b101 *
0-
02
b101 6
#992750000000
1!
1%
1-
12
#992760000000
0!
0%
b110 *
0-
02
b110 6
#992770000000
1!
1%
1-
12
#992780000000
0!
0%
b111 *
0-
02
b111 6
#992790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#992800000000
0!
0%
b0 *
0-
02
b0 6
#992810000000
1!
1%
1-
12
#992820000000
0!
0%
b1 *
0-
02
b1 6
#992830000000
1!
1%
1-
12
#992840000000
0!
0%
b10 *
0-
02
b10 6
#992850000000
1!
1%
1-
12
#992860000000
0!
0%
b11 *
0-
02
b11 6
#992870000000
1!
1%
1-
12
15
#992880000000
0!
0%
b100 *
0-
02
b100 6
#992890000000
1!
1%
1-
12
#992900000000
0!
0%
b101 *
0-
02
b101 6
#992910000000
1!
1%
1-
12
#992920000000
0!
0%
b110 *
0-
02
b110 6
#992930000000
1!
1%
1-
12
#992940000000
0!
0%
b111 *
0-
02
b111 6
#992950000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#992960000000
0!
0%
b0 *
0-
02
b0 6
#992970000000
1!
1%
1-
12
#992980000000
0!
0%
b1 *
0-
02
b1 6
#992990000000
1!
1%
1-
12
#993000000000
0!
0%
b10 *
0-
02
b10 6
#993010000000
1!
1%
1-
12
#993020000000
0!
0%
b11 *
0-
02
b11 6
#993030000000
1!
1%
1-
12
15
#993040000000
0!
0%
b100 *
0-
02
b100 6
#993050000000
1!
1%
1-
12
#993060000000
0!
0%
b101 *
0-
02
b101 6
#993070000000
1!
1%
1-
12
#993080000000
0!
0%
b110 *
0-
02
b110 6
#993090000000
1!
1%
1-
12
#993100000000
0!
0%
b111 *
0-
02
b111 6
#993110000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#993120000000
0!
0%
b0 *
0-
02
b0 6
#993130000000
1!
1%
1-
12
#993140000000
0!
0%
b1 *
0-
02
b1 6
#993150000000
1!
1%
1-
12
#993160000000
0!
0%
b10 *
0-
02
b10 6
#993170000000
1!
1%
1-
12
#993180000000
0!
0%
b11 *
0-
02
b11 6
#993190000000
1!
1%
1-
12
15
#993200000000
0!
0%
b100 *
0-
02
b100 6
#993210000000
1!
1%
1-
12
#993220000000
0!
0%
b101 *
0-
02
b101 6
#993230000000
1!
1%
1-
12
#993240000000
0!
0%
b110 *
0-
02
b110 6
#993250000000
1!
1%
1-
12
#993260000000
0!
0%
b111 *
0-
02
b111 6
#993270000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#993280000000
0!
0%
b0 *
0-
02
b0 6
#993290000000
1!
1%
1-
12
#993300000000
0!
0%
b1 *
0-
02
b1 6
#993310000000
1!
1%
1-
12
#993320000000
0!
0%
b10 *
0-
02
b10 6
#993330000000
1!
1%
1-
12
#993340000000
0!
0%
b11 *
0-
02
b11 6
#993350000000
1!
1%
1-
12
15
#993360000000
0!
0%
b100 *
0-
02
b100 6
#993370000000
1!
1%
1-
12
#993380000000
0!
0%
b101 *
0-
02
b101 6
#993390000000
1!
1%
1-
12
#993400000000
0!
0%
b110 *
0-
02
b110 6
#993410000000
1!
1%
1-
12
#993420000000
0!
0%
b111 *
0-
02
b111 6
#993430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#993440000000
0!
0%
b0 *
0-
02
b0 6
#993450000000
1!
1%
1-
12
#993460000000
0!
0%
b1 *
0-
02
b1 6
#993470000000
1!
1%
1-
12
#993480000000
0!
0%
b10 *
0-
02
b10 6
#993490000000
1!
1%
1-
12
#993500000000
0!
0%
b11 *
0-
02
b11 6
#993510000000
1!
1%
1-
12
15
#993520000000
0!
0%
b100 *
0-
02
b100 6
#993530000000
1!
1%
1-
12
#993540000000
0!
0%
b101 *
0-
02
b101 6
#993550000000
1!
1%
1-
12
#993560000000
0!
0%
b110 *
0-
02
b110 6
#993570000000
1!
1%
1-
12
#993580000000
0!
0%
b111 *
0-
02
b111 6
#993590000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#993600000000
0!
0%
b0 *
0-
02
b0 6
#993610000000
1!
1%
1-
12
#993620000000
0!
0%
b1 *
0-
02
b1 6
#993630000000
1!
1%
1-
12
#993640000000
0!
0%
b10 *
0-
02
b10 6
#993650000000
1!
1%
1-
12
#993660000000
0!
0%
b11 *
0-
02
b11 6
#993670000000
1!
1%
1-
12
15
#993680000000
0!
0%
b100 *
0-
02
b100 6
#993690000000
1!
1%
1-
12
#993700000000
0!
0%
b101 *
0-
02
b101 6
#993710000000
1!
1%
1-
12
#993720000000
0!
0%
b110 *
0-
02
b110 6
#993730000000
1!
1%
1-
12
#993740000000
0!
0%
b111 *
0-
02
b111 6
#993750000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#993760000000
0!
0%
b0 *
0-
02
b0 6
#993770000000
1!
1%
1-
12
#993780000000
0!
0%
b1 *
0-
02
b1 6
#993790000000
1!
1%
1-
12
#993800000000
0!
0%
b10 *
0-
02
b10 6
#993810000000
1!
1%
1-
12
#993820000000
0!
0%
b11 *
0-
02
b11 6
#993830000000
1!
1%
1-
12
15
#993840000000
0!
0%
b100 *
0-
02
b100 6
#993850000000
1!
1%
1-
12
#993860000000
0!
0%
b101 *
0-
02
b101 6
#993870000000
1!
1%
1-
12
#993880000000
0!
0%
b110 *
0-
02
b110 6
#993890000000
1!
1%
1-
12
#993900000000
0!
0%
b111 *
0-
02
b111 6
#993910000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#993920000000
0!
0%
b0 *
0-
02
b0 6
#993930000000
1!
1%
1-
12
#993940000000
0!
0%
b1 *
0-
02
b1 6
#993950000000
1!
1%
1-
12
#993960000000
0!
0%
b10 *
0-
02
b10 6
#993970000000
1!
1%
1-
12
#993980000000
0!
0%
b11 *
0-
02
b11 6
#993990000000
1!
1%
1-
12
15
#994000000000
0!
0%
b100 *
0-
02
b100 6
#994010000000
1!
1%
1-
12
#994020000000
0!
0%
b101 *
0-
02
b101 6
#994030000000
1!
1%
1-
12
#994040000000
0!
0%
b110 *
0-
02
b110 6
#994050000000
1!
1%
1-
12
#994060000000
0!
0%
b111 *
0-
02
b111 6
#994070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#994080000000
0!
0%
b0 *
0-
02
b0 6
#994090000000
1!
1%
1-
12
#994100000000
0!
0%
b1 *
0-
02
b1 6
#994110000000
1!
1%
1-
12
#994120000000
0!
0%
b10 *
0-
02
b10 6
#994130000000
1!
1%
1-
12
#994140000000
0!
0%
b11 *
0-
02
b11 6
#994150000000
1!
1%
1-
12
15
#994160000000
0!
0%
b100 *
0-
02
b100 6
#994170000000
1!
1%
1-
12
#994180000000
0!
0%
b101 *
0-
02
b101 6
#994190000000
1!
1%
1-
12
#994200000000
0!
0%
b110 *
0-
02
b110 6
#994210000000
1!
1%
1-
12
#994220000000
0!
0%
b111 *
0-
02
b111 6
#994230000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#994240000000
0!
0%
b0 *
0-
02
b0 6
#994250000000
1!
1%
1-
12
#994260000000
0!
0%
b1 *
0-
02
b1 6
#994270000000
1!
1%
1-
12
#994280000000
0!
0%
b10 *
0-
02
b10 6
#994290000000
1!
1%
1-
12
#994300000000
0!
0%
b11 *
0-
02
b11 6
#994310000000
1!
1%
1-
12
15
#994320000000
0!
0%
b100 *
0-
02
b100 6
#994330000000
1!
1%
1-
12
#994340000000
0!
0%
b101 *
0-
02
b101 6
#994350000000
1!
1%
1-
12
#994360000000
0!
0%
b110 *
0-
02
b110 6
#994370000000
1!
1%
1-
12
#994380000000
0!
0%
b111 *
0-
02
b111 6
#994390000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#994400000000
0!
0%
b0 *
0-
02
b0 6
#994410000000
1!
1%
1-
12
#994420000000
0!
0%
b1 *
0-
02
b1 6
#994430000000
1!
1%
1-
12
#994440000000
0!
0%
b10 *
0-
02
b10 6
#994450000000
1!
1%
1-
12
#994460000000
0!
0%
b11 *
0-
02
b11 6
#994470000000
1!
1%
1-
12
15
#994480000000
0!
0%
b100 *
0-
02
b100 6
#994490000000
1!
1%
1-
12
#994500000000
0!
0%
b101 *
0-
02
b101 6
#994510000000
1!
1%
1-
12
#994520000000
0!
0%
b110 *
0-
02
b110 6
#994530000000
1!
1%
1-
12
#994540000000
0!
0%
b111 *
0-
02
b111 6
#994550000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#994560000000
0!
0%
b0 *
0-
02
b0 6
#994570000000
1!
1%
1-
12
#994580000000
0!
0%
b1 *
0-
02
b1 6
#994590000000
1!
1%
1-
12
#994600000000
0!
0%
b10 *
0-
02
b10 6
#994610000000
1!
1%
1-
12
#994620000000
0!
0%
b11 *
0-
02
b11 6
#994630000000
1!
1%
1-
12
15
#994640000000
0!
0%
b100 *
0-
02
b100 6
#994650000000
1!
1%
1-
12
#994660000000
0!
0%
b101 *
0-
02
b101 6
#994670000000
1!
1%
1-
12
#994680000000
0!
0%
b110 *
0-
02
b110 6
#994690000000
1!
1%
1-
12
#994700000000
0!
0%
b111 *
0-
02
b111 6
#994710000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#994720000000
0!
0%
b0 *
0-
02
b0 6
#994730000000
1!
1%
1-
12
#994740000000
0!
0%
b1 *
0-
02
b1 6
#994750000000
1!
1%
1-
12
#994760000000
0!
0%
b10 *
0-
02
b10 6
#994770000000
1!
1%
1-
12
#994780000000
0!
0%
b11 *
0-
02
b11 6
#994790000000
1!
1%
1-
12
15
#994800000000
0!
0%
b100 *
0-
02
b100 6
#994810000000
1!
1%
1-
12
#994820000000
0!
0%
b101 *
0-
02
b101 6
#994830000000
1!
1%
1-
12
#994840000000
0!
0%
b110 *
0-
02
b110 6
#994850000000
1!
1%
1-
12
#994860000000
0!
0%
b111 *
0-
02
b111 6
#994870000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#994880000000
0!
0%
b0 *
0-
02
b0 6
#994890000000
1!
1%
1-
12
#994900000000
0!
0%
b1 *
0-
02
b1 6
#994910000000
1!
1%
1-
12
#994920000000
0!
0%
b10 *
0-
02
b10 6
#994930000000
1!
1%
1-
12
#994940000000
0!
0%
b11 *
0-
02
b11 6
#994950000000
1!
1%
1-
12
15
#994960000000
0!
0%
b100 *
0-
02
b100 6
#994970000000
1!
1%
1-
12
#994980000000
0!
0%
b101 *
0-
02
b101 6
#994990000000
1!
1%
1-
12
#995000000000
0!
0%
b110 *
0-
02
b110 6
#995010000000
1!
1%
1-
12
#995020000000
0!
0%
b111 *
0-
02
b111 6
#995030000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#995040000000
0!
0%
b0 *
0-
02
b0 6
#995050000000
1!
1%
1-
12
#995060000000
0!
0%
b1 *
0-
02
b1 6
#995070000000
1!
1%
1-
12
#995080000000
0!
0%
b10 *
0-
02
b10 6
#995090000000
1!
1%
1-
12
#995100000000
0!
0%
b11 *
0-
02
b11 6
#995110000000
1!
1%
1-
12
15
#995120000000
0!
0%
b100 *
0-
02
b100 6
#995130000000
1!
1%
1-
12
#995140000000
0!
0%
b101 *
0-
02
b101 6
#995150000000
1!
1%
1-
12
#995160000000
0!
0%
b110 *
0-
02
b110 6
#995170000000
1!
1%
1-
12
#995180000000
0!
0%
b111 *
0-
02
b111 6
#995190000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#995200000000
0!
0%
b0 *
0-
02
b0 6
#995210000000
1!
1%
1-
12
#995220000000
0!
0%
b1 *
0-
02
b1 6
#995230000000
1!
1%
1-
12
#995240000000
0!
0%
b10 *
0-
02
b10 6
#995250000000
1!
1%
1-
12
#995260000000
0!
0%
b11 *
0-
02
b11 6
#995270000000
1!
1%
1-
12
15
#995280000000
0!
0%
b100 *
0-
02
b100 6
#995290000000
1!
1%
1-
12
#995300000000
0!
0%
b101 *
0-
02
b101 6
#995310000000
1!
1%
1-
12
#995320000000
0!
0%
b110 *
0-
02
b110 6
#995330000000
1!
1%
1-
12
#995340000000
0!
0%
b111 *
0-
02
b111 6
#995350000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#995360000000
0!
0%
b0 *
0-
02
b0 6
#995370000000
1!
1%
1-
12
#995380000000
0!
0%
b1 *
0-
02
b1 6
#995390000000
1!
1%
1-
12
#995400000000
0!
0%
b10 *
0-
02
b10 6
#995410000000
1!
1%
1-
12
#995420000000
0!
0%
b11 *
0-
02
b11 6
#995430000000
1!
1%
1-
12
15
#995440000000
0!
0%
b100 *
0-
02
b100 6
#995450000000
1!
1%
1-
12
#995460000000
0!
0%
b101 *
0-
02
b101 6
#995470000000
1!
1%
1-
12
#995480000000
0!
0%
b110 *
0-
02
b110 6
#995490000000
1!
1%
1-
12
#995500000000
0!
0%
b111 *
0-
02
b111 6
#995510000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#995520000000
0!
0%
b0 *
0-
02
b0 6
#995530000000
1!
1%
1-
12
#995540000000
0!
0%
b1 *
0-
02
b1 6
#995550000000
1!
1%
1-
12
#995560000000
0!
0%
b10 *
0-
02
b10 6
#995570000000
1!
1%
1-
12
#995580000000
0!
0%
b11 *
0-
02
b11 6
#995590000000
1!
1%
1-
12
15
#995600000000
0!
0%
b100 *
0-
02
b100 6
#995610000000
1!
1%
1-
12
#995620000000
0!
0%
b101 *
0-
02
b101 6
#995630000000
1!
1%
1-
12
#995640000000
0!
0%
b110 *
0-
02
b110 6
#995650000000
1!
1%
1-
12
#995660000000
0!
0%
b111 *
0-
02
b111 6
#995670000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#995680000000
0!
0%
b0 *
0-
02
b0 6
#995690000000
1!
1%
1-
12
#995700000000
0!
0%
b1 *
0-
02
b1 6
#995710000000
1!
1%
1-
12
#995720000000
0!
0%
b10 *
0-
02
b10 6
#995730000000
1!
1%
1-
12
#995740000000
0!
0%
b11 *
0-
02
b11 6
#995750000000
1!
1%
1-
12
15
#995760000000
0!
0%
b100 *
0-
02
b100 6
#995770000000
1!
1%
1-
12
#995780000000
0!
0%
b101 *
0-
02
b101 6
#995790000000
1!
1%
1-
12
#995800000000
0!
0%
b110 *
0-
02
b110 6
#995810000000
1!
1%
1-
12
#995820000000
0!
0%
b111 *
0-
02
b111 6
#995830000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#995840000000
0!
0%
b0 *
0-
02
b0 6
#995850000000
1!
1%
1-
12
#995860000000
0!
0%
b1 *
0-
02
b1 6
#995870000000
1!
1%
1-
12
#995880000000
0!
0%
b10 *
0-
02
b10 6
#995890000000
1!
1%
1-
12
#995900000000
0!
0%
b11 *
0-
02
b11 6
#995910000000
1!
1%
1-
12
15
#995920000000
0!
0%
b100 *
0-
02
b100 6
#995930000000
1!
1%
1-
12
#995940000000
0!
0%
b101 *
0-
02
b101 6
#995950000000
1!
1%
1-
12
#995960000000
0!
0%
b110 *
0-
02
b110 6
#995970000000
1!
1%
1-
12
#995980000000
0!
0%
b111 *
0-
02
b111 6
#995990000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#996000000000
0!
0%
b0 *
0-
02
b0 6
#996010000000
1!
1%
1-
12
#996020000000
0!
0%
b1 *
0-
02
b1 6
#996030000000
1!
1%
1-
12
#996040000000
0!
0%
b10 *
0-
02
b10 6
#996050000000
1!
1%
1-
12
#996060000000
0!
0%
b11 *
0-
02
b11 6
#996070000000
1!
1%
1-
12
15
#996080000000
0!
0%
b100 *
0-
02
b100 6
#996090000000
1!
1%
1-
12
#996100000000
0!
0%
b101 *
0-
02
b101 6
#996110000000
1!
1%
1-
12
#996120000000
0!
0%
b110 *
0-
02
b110 6
#996130000000
1!
1%
1-
12
#996140000000
0!
0%
b111 *
0-
02
b111 6
#996150000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#996160000000
0!
0%
b0 *
0-
02
b0 6
#996170000000
1!
1%
1-
12
#996180000000
0!
0%
b1 *
0-
02
b1 6
#996190000000
1!
1%
1-
12
#996200000000
0!
0%
b10 *
0-
02
b10 6
#996210000000
1!
1%
1-
12
#996220000000
0!
0%
b11 *
0-
02
b11 6
#996230000000
1!
1%
1-
12
15
#996240000000
0!
0%
b100 *
0-
02
b100 6
#996250000000
1!
1%
1-
12
#996260000000
0!
0%
b101 *
0-
02
b101 6
#996270000000
1!
1%
1-
12
#996280000000
0!
0%
b110 *
0-
02
b110 6
#996290000000
1!
1%
1-
12
#996300000000
0!
0%
b111 *
0-
02
b111 6
#996310000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#996320000000
0!
0%
b0 *
0-
02
b0 6
#996330000000
1!
1%
1-
12
#996340000000
0!
0%
b1 *
0-
02
b1 6
#996350000000
1!
1%
1-
12
#996360000000
0!
0%
b10 *
0-
02
b10 6
#996370000000
1!
1%
1-
12
#996380000000
0!
0%
b11 *
0-
02
b11 6
#996390000000
1!
1%
1-
12
15
#996400000000
0!
0%
b100 *
0-
02
b100 6
#996410000000
1!
1%
1-
12
#996420000000
0!
0%
b101 *
0-
02
b101 6
#996430000000
1!
1%
1-
12
#996440000000
0!
0%
b110 *
0-
02
b110 6
#996450000000
1!
1%
1-
12
#996460000000
0!
0%
b111 *
0-
02
b111 6
#996470000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#996480000000
0!
0%
b0 *
0-
02
b0 6
#996490000000
1!
1%
1-
12
#996500000000
0!
0%
b1 *
0-
02
b1 6
#996510000000
1!
1%
1-
12
#996520000000
0!
0%
b10 *
0-
02
b10 6
#996530000000
1!
1%
1-
12
#996540000000
0!
0%
b11 *
0-
02
b11 6
#996550000000
1!
1%
1-
12
15
#996560000000
0!
0%
b100 *
0-
02
b100 6
#996570000000
1!
1%
1-
12
#996580000000
0!
0%
b101 *
0-
02
b101 6
#996590000000
1!
1%
1-
12
#996600000000
0!
0%
b110 *
0-
02
b110 6
#996610000000
1!
1%
1-
12
#996620000000
0!
0%
b111 *
0-
02
b111 6
#996630000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#996640000000
0!
0%
b0 *
0-
02
b0 6
#996650000000
1!
1%
1-
12
#996660000000
0!
0%
b1 *
0-
02
b1 6
#996670000000
1!
1%
1-
12
#996680000000
0!
0%
b10 *
0-
02
b10 6
#996690000000
1!
1%
1-
12
#996700000000
0!
0%
b11 *
0-
02
b11 6
#996710000000
1!
1%
1-
12
15
#996720000000
0!
0%
b100 *
0-
02
b100 6
#996730000000
1!
1%
1-
12
#996740000000
0!
0%
b101 *
0-
02
b101 6
#996750000000
1!
1%
1-
12
#996760000000
0!
0%
b110 *
0-
02
b110 6
#996770000000
1!
1%
1-
12
#996780000000
0!
0%
b111 *
0-
02
b111 6
#996790000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#996800000000
0!
0%
b0 *
0-
02
b0 6
#996810000000
1!
1%
1-
12
#996820000000
0!
0%
b1 *
0-
02
b1 6
#996830000000
1!
1%
1-
12
#996840000000
0!
0%
b10 *
0-
02
b10 6
#996850000000
1!
1%
1-
12
#996860000000
0!
0%
b11 *
0-
02
b11 6
#996870000000
1!
1%
1-
12
15
#996880000000
0!
0%
b100 *
0-
02
b100 6
#996890000000
1!
1%
1-
12
#996900000000
0!
0%
b101 *
0-
02
b101 6
#996910000000
1!
1%
1-
12
#996920000000
0!
0%
b110 *
0-
02
b110 6
#996930000000
1!
1%
1-
12
#996940000000
0!
0%
b111 *
0-
02
b111 6
#996950000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#996960000000
0!
0%
b0 *
0-
02
b0 6
#996970000000
1!
1%
1-
12
#996980000000
0!
0%
b1 *
0-
02
b1 6
#996990000000
1!
1%
1-
12
#997000000000
0!
0%
b10 *
0-
02
b10 6
#997010000000
1!
1%
1-
12
#997020000000
0!
0%
b11 *
0-
02
b11 6
#997030000000
1!
1%
1-
12
15
#997040000000
0!
0%
b100 *
0-
02
b100 6
#997050000000
1!
1%
1-
12
#997060000000
0!
0%
b101 *
0-
02
b101 6
#997070000000
1!
1%
1-
12
#997080000000
0!
0%
b110 *
0-
02
b110 6
#997090000000
1!
1%
1-
12
#997100000000
0!
0%
b111 *
0-
02
b111 6
#997110000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#997120000000
0!
0%
b0 *
0-
02
b0 6
#997130000000
1!
1%
1-
12
#997140000000
0!
0%
b1 *
0-
02
b1 6
#997150000000
1!
1%
1-
12
#997160000000
0!
0%
b10 *
0-
02
b10 6
#997170000000
1!
1%
1-
12
#997180000000
0!
0%
b11 *
0-
02
b11 6
#997190000000
1!
1%
1-
12
15
#997200000000
0!
0%
b100 *
0-
02
b100 6
#997210000000
1!
1%
1-
12
#997220000000
0!
0%
b101 *
0-
02
b101 6
#997230000000
1!
1%
1-
12
#997240000000
0!
0%
b110 *
0-
02
b110 6
#997250000000
1!
1%
1-
12
#997260000000
0!
0%
b111 *
0-
02
b111 6
#997270000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#997280000000
0!
0%
b0 *
0-
02
b0 6
#997290000000
1!
1%
1-
12
#997300000000
0!
0%
b1 *
0-
02
b1 6
#997310000000
1!
1%
1-
12
#997320000000
0!
0%
b10 *
0-
02
b10 6
#997330000000
1!
1%
1-
12
#997340000000
0!
0%
b11 *
0-
02
b11 6
#997350000000
1!
1%
1-
12
15
#997360000000
0!
0%
b100 *
0-
02
b100 6
#997370000000
1!
1%
1-
12
#997380000000
0!
0%
b101 *
0-
02
b101 6
#997390000000
1!
1%
1-
12
#997400000000
0!
0%
b110 *
0-
02
b110 6
#997410000000
1!
1%
1-
12
#997420000000
0!
0%
b111 *
0-
02
b111 6
#997430000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#997440000000
0!
0%
b0 *
0-
02
b0 6
#997450000000
1!
1%
1-
12
#997460000000
0!
0%
b1 *
0-
02
b1 6
#997470000000
1!
1%
1-
12
#997480000000
0!
0%
b10 *
0-
02
b10 6
#997490000000
1!
1%
1-
12
#997500000000
0!
0%
b11 *
0-
02
b11 6
#997510000000
1!
1%
1-
12
15
#997520000000
0!
0%
b100 *
0-
02
b100 6
#997530000000
1!
1%
1-
12
#997540000000
0!
0%
b101 *
0-
02
b101 6
#997550000000
1!
1%
1-
12
#997560000000
0!
0%
b110 *
0-
02
b110 6
#997570000000
1!
1%
1-
12
#997580000000
0!
0%
b111 *
0-
02
b111 6
#997590000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#997600000000
0!
0%
b0 *
0-
02
b0 6
#997610000000
1!
1%
1-
12
#997620000000
0!
0%
b1 *
0-
02
b1 6
#997630000000
1!
1%
1-
12
#997640000000
0!
0%
b10 *
0-
02
b10 6
#997650000000
1!
1%
1-
12
#997660000000
0!
0%
b11 *
0-
02
b11 6
#997670000000
1!
1%
1-
12
15
#997680000000
0!
0%
b100 *
0-
02
b100 6
#997690000000
1!
1%
1-
12
#997700000000
0!
0%
b101 *
0-
02
b101 6
#997710000000
1!
1%
1-
12
#997720000000
0!
0%
b110 *
0-
02
b110 6
#997730000000
1!
1%
1-
12
#997740000000
0!
0%
b111 *
0-
02
b111 6
#997750000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#997760000000
0!
0%
b0 *
0-
02
b0 6
#997770000000
1!
1%
1-
12
#997780000000
0!
0%
b1 *
0-
02
b1 6
#997790000000
1!
1%
1-
12
#997800000000
0!
0%
b10 *
0-
02
b10 6
#997810000000
1!
1%
1-
12
#997820000000
0!
0%
b11 *
0-
02
b11 6
#997830000000
1!
1%
1-
12
15
#997840000000
0!
0%
b100 *
0-
02
b100 6
#997850000000
1!
1%
1-
12
#997860000000
0!
0%
b101 *
0-
02
b101 6
#997870000000
1!
1%
1-
12
#997880000000
0!
0%
b110 *
0-
02
b110 6
#997890000000
1!
1%
1-
12
#997900000000
0!
0%
b111 *
0-
02
b111 6
#997910000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#997920000000
0!
0%
b0 *
0-
02
b0 6
#997930000000
1!
1%
1-
12
#997940000000
0!
0%
b1 *
0-
02
b1 6
#997950000000
1!
1%
1-
12
#997960000000
0!
0%
b10 *
0-
02
b10 6
#997970000000
1!
1%
1-
12
#997980000000
0!
0%
b11 *
0-
02
b11 6
#997990000000
1!
1%
1-
12
15
#998000000000
0!
0%
b100 *
0-
02
b100 6
#998010000000
1!
1%
1-
12
#998020000000
0!
0%
b101 *
0-
02
b101 6
#998030000000
1!
1%
1-
12
#998040000000
0!
0%
b110 *
0-
02
b110 6
#998050000000
1!
1%
1-
12
#998060000000
0!
0%
b111 *
0-
02
b111 6
#998070000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#998080000000
0!
0%
b0 *
0-
02
b0 6
#998090000000
1!
1%
1-
12
#998100000000
0!
0%
b1 *
0-
02
b1 6
#998110000000
1!
1%
1-
12
#998120000000
0!
0%
b10 *
0-
02
b10 6
#998130000000
1!
1%
1-
12
#998140000000
0!
0%
b11 *
0-
02
b11 6
#998150000000
1!
1%
1-
12
15
#998160000000
0!
0%
b100 *
0-
02
b100 6
#998170000000
1!
1%
1-
12
#998180000000
0!
0%
b101 *
0-
02
b101 6
#998190000000
1!
1%
1-
12
#998200000000
0!
0%
b110 *
0-
02
b110 6
#998210000000
1!
1%
1-
12
#998220000000
0!
0%
b111 *
0-
02
b111 6
#998230000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#998240000000
0!
0%
b0 *
0-
02
b0 6
#998250000000
1!
1%
1-
12
#998260000000
0!
0%
b1 *
0-
02
b1 6
#998270000000
1!
1%
1-
12
#998280000000
0!
0%
b10 *
0-
02
b10 6
#998290000000
1!
1%
1-
12
#998300000000
0!
0%
b11 *
0-
02
b11 6
#998310000000
1!
1%
1-
12
15
#998320000000
0!
0%
b100 *
0-
02
b100 6
#998330000000
1!
1%
1-
12
#998340000000
0!
0%
b101 *
0-
02
b101 6
#998350000000
1!
1%
1-
12
#998360000000
0!
0%
b110 *
0-
02
b110 6
#998370000000
1!
1%
1-
12
#998380000000
0!
0%
b111 *
0-
02
b111 6
#998390000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#998400000000
0!
0%
b0 *
0-
02
b0 6
#998410000000
1!
1%
1-
12
#998420000000
0!
0%
b1 *
0-
02
b1 6
#998430000000
1!
1%
1-
12
#998440000000
0!
0%
b10 *
0-
02
b10 6
#998450000000
1!
1%
1-
12
#998460000000
0!
0%
b11 *
0-
02
b11 6
#998470000000
1!
1%
1-
12
15
#998480000000
0!
0%
b100 *
0-
02
b100 6
#998490000000
1!
1%
1-
12
#998500000000
0!
0%
b101 *
0-
02
b101 6
#998510000000
1!
1%
1-
12
#998520000000
0!
0%
b110 *
0-
02
b110 6
#998530000000
1!
1%
1-
12
#998540000000
0!
0%
b111 *
0-
02
b111 6
#998550000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#998560000000
0!
0%
b0 *
0-
02
b0 6
#998570000000
1!
1%
1-
12
#998580000000
0!
0%
b1 *
0-
02
b1 6
#998590000000
1!
1%
1-
12
#998600000000
0!
0%
b10 *
0-
02
b10 6
#998610000000
1!
1%
1-
12
#998620000000
0!
0%
b11 *
0-
02
b11 6
#998630000000
1!
1%
1-
12
15
#998640000000
0!
0%
b100 *
0-
02
b100 6
#998650000000
1!
1%
1-
12
#998660000000
0!
0%
b101 *
0-
02
b101 6
#998670000000
1!
1%
1-
12
#998680000000
0!
0%
b110 *
0-
02
b110 6
#998690000000
1!
1%
1-
12
#998700000000
0!
0%
b111 *
0-
02
b111 6
#998710000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#998720000000
0!
0%
b0 *
0-
02
b0 6
#998730000000
1!
1%
1-
12
#998740000000
0!
0%
b1 *
0-
02
b1 6
#998750000000
1!
1%
1-
12
#998760000000
0!
0%
b10 *
0-
02
b10 6
#998770000000
1!
1%
1-
12
#998780000000
0!
0%
b11 *
0-
02
b11 6
#998790000000
1!
1%
1-
12
15
#998800000000
0!
0%
b100 *
0-
02
b100 6
#998810000000
1!
1%
1-
12
#998820000000
0!
0%
b101 *
0-
02
b101 6
#998830000000
1!
1%
1-
12
#998840000000
0!
0%
b110 *
0-
02
b110 6
#998850000000
1!
1%
1-
12
#998860000000
0!
0%
b111 *
0-
02
b111 6
#998870000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#998880000000
0!
0%
b0 *
0-
02
b0 6
#998890000000
1!
1%
1-
12
#998900000000
0!
0%
b1 *
0-
02
b1 6
#998910000000
1!
1%
1-
12
#998920000000
0!
0%
b10 *
0-
02
b10 6
#998930000000
1!
1%
1-
12
#998940000000
0!
0%
b11 *
0-
02
b11 6
#998950000000
1!
1%
1-
12
15
#998960000000
0!
0%
b100 *
0-
02
b100 6
#998970000000
1!
1%
1-
12
#998980000000
0!
0%
b101 *
0-
02
b101 6
#998990000000
1!
1%
1-
12
#999000000000
0!
0%
b110 *
0-
02
b110 6
#999010000000
1!
1%
1-
12
#999020000000
0!
0%
b111 *
0-
02
b111 6
#999030000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#999040000000
0!
0%
b0 *
0-
02
b0 6
#999050000000
1!
1%
1-
12
#999060000000
0!
0%
b1 *
0-
02
b1 6
#999070000000
1!
1%
1-
12
#999080000000
0!
0%
b10 *
0-
02
b10 6
#999090000000
1!
1%
1-
12
#999100000000
0!
0%
b11 *
0-
02
b11 6
#999110000000
1!
1%
1-
12
15
#999120000000
0!
0%
b100 *
0-
02
b100 6
#999130000000
1!
1%
1-
12
#999140000000
0!
0%
b101 *
0-
02
b101 6
#999150000000
1!
1%
1-
12
#999160000000
0!
0%
b110 *
0-
02
b110 6
#999170000000
1!
1%
1-
12
#999180000000
0!
0%
b111 *
0-
02
b111 6
#999190000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#999200000000
0!
0%
b0 *
0-
02
b0 6
#999210000000
1!
1%
1-
12
#999220000000
0!
0%
b1 *
0-
02
b1 6
#999230000000
1!
1%
1-
12
#999240000000
0!
0%
b10 *
0-
02
b10 6
#999250000000
1!
1%
1-
12
#999260000000
0!
0%
b11 *
0-
02
b11 6
#999270000000
1!
1%
1-
12
15
#999280000000
0!
0%
b100 *
0-
02
b100 6
#999290000000
1!
1%
1-
12
#999300000000
0!
0%
b101 *
0-
02
b101 6
#999310000000
1!
1%
1-
12
#999320000000
0!
0%
b110 *
0-
02
b110 6
#999330000000
1!
1%
1-
12
#999340000000
0!
0%
b111 *
0-
02
b111 6
#999350000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#999360000000
0!
0%
b0 *
0-
02
b0 6
#999370000000
1!
1%
1-
12
#999380000000
0!
0%
b1 *
0-
02
b1 6
#999390000000
1!
1%
1-
12
#999400000000
0!
0%
b10 *
0-
02
b10 6
#999410000000
1!
1%
1-
12
#999420000000
0!
0%
b11 *
0-
02
b11 6
#999430000000
1!
1%
1-
12
15
#999440000000
0!
0%
b100 *
0-
02
b100 6
#999450000000
1!
1%
1-
12
#999460000000
0!
0%
b101 *
0-
02
b101 6
#999470000000
1!
1%
1-
12
#999480000000
0!
0%
b110 *
0-
02
b110 6
#999490000000
1!
1%
1-
12
#999500000000
0!
0%
b111 *
0-
02
b111 6
#999510000000
1!
b0001 #
b0110011 $
1%
b0001 '
b0110011 (
b0100 )
1-
12
05
b0110011 7
b0100 8
#999520000000
0!
0%
b0 *
0-
02
b0 6
#999530000000
1!
1%
1-
12
#999540000000
0!
0%
b1 *
0-
02
b1 6
#999550000000
1!
1%
1-
12
#999560000000
0!
0%
b10 *
0-
02
b10 6
#999570000000
1!
1%
1-
12
#999580000000
0!
0%
b11 *
0-
02
b11 6
#999590000000
1!
1%
1-
12
15
#999600000000
0!
0%
b100 *
0-
02
b100 6
#999610000000
1!
1%
1-
12
#999620000000
0!
0%
b101 *
0-
02
b101 6
#999630000000
1!
1%
1-
12
#999640000000
0!
0%
b110 *
0-
02
b110 6
#999650000000
1!
1%
1-
12
#999660000000
0!
0%
b111 *
0-
02
b111 6
#999670000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
1-
12
05
b0110000 7
b0001 8
#999680000000
0!
0%
b0 *
0-
02
b0 6
#999690000000
1!
1%
1-
12
#999700000000
0!
0%
b1 *
0-
02
b1 6
#999710000000
1!
1%
1-
12
#999720000000
0!
0%
b10 *
0-
02
b10 6
#999730000000
1!
1%
1-
12
#999740000000
0!
0%
b11 *
0-
02
b11 6
#999750000000
1!
1%
1-
12
15
#999760000000
0!
0%
b100 *
0-
02
b100 6
#999770000000
1!
1%
1-
12
#999780000000
0!
0%
b101 *
0-
02
b101 6
#999790000000
1!
1%
1-
12
#999800000000
0!
0%
b110 *
0-
02
b110 6
#999810000000
1!
1%
1-
12
#999820000000
0!
0%
b111 *
0-
02
b111 6
#999830000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1-
12
05
b1101101 7
b0010 8
#999840000000
0!
0%
b0 *
0-
02
b0 6
#999850000000
1!
1%
1-
12
#999860000000
0!
0%
b1 *
0-
02
b1 6
#999870000000
1!
1%
1-
12
#999880000000
0!
0%
b10 *
0-
02
b10 6
#999890000000
1!
1%
1-
12
#999900000000
0!
0%
b11 *
0-
02
b11 6
#999910000000
1!
1%
1-
12
15
#999920000000
0!
0%
b100 *
0-
02
b100 6
#999930000000
1!
1%
1-
12
#999940000000
0!
0%
b101 *
0-
02
b101 6
#999950000000
1!
1%
1-
12
#999960000000
0!
0%
b110 *
0-
02
b110 6
#999970000000
1!
1%
1-
12
#999980000000
0!
0%
b111 *
0-
02
b111 6
#999990000000
1!
b0010 #
b1111001 $
1%
b0010 '
b1111001 (
b0011 )
1-
12
05
b1111001 7
b0011 8
#1000000000000
0!
0%
b0 *
0-
02
b0 6
