$date
  Tue May 14 14:42:28 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_motor $end
$var reg 1 ! clk $end
$var reg 1 " key_asc $end
$var reg 1 # key_desc $end
$var reg 1 $ key_frec $end
$var reg 1 % enable_disp $end
$var reg 7 & segmentos[6:0] $end
$var reg 4 ' salida[3:0] $end
$scope module uut $end
$var reg 1 ( clk $end
$var reg 1 ) key_asc $end
$var reg 1 * key_desc $end
$var reg 1 + key_frec $end
$var reg 1 , enable_disp $end
$var reg 7 - segmentos[6:0] $end
$var reg 4 . salida[3:0] $end
$comment state is not handled $end
$var integer 32 / cuenta $end
$var integer 32 0 cuenta_maxima $end
$var integer 32 1 aux $end
$var integer 32 2 cuenta2 $end
$var reg 4 3 bcd_disp[3:0] $end
$scope module a $end
$var reg 1 4 clk $end
$var reg 1 5 reset $end
$var reg 1 6 enable $end
$var reg 1 7 cout $end
$var integer 32 8 q $end
$upscope $end
$scope module a2 $end
$var reg 1 9 clk $end
$var reg 1 : reset $end
$var reg 1 ; enable $end
$var reg 1 < cout $end
$var integer 32 = q $end
$upscope $end
$scope module b $end
$var reg 7 > segmentos[6:0] $end
$var reg 4 ? bcd[3:0] $end
$var reg 1 @ enable $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
0#
0$
0%
b0000001 &
b1000 '
0(
0)
0*
0+
0,
b0000001 -
b1000 .
b0 /
b101 0
b0 1
b0 2
b0000 3
04
05
16
U7
b0 8
09
0:
1;
U<
b0 =
b0000001 >
b0000 ?
0@
#10000000
1!
1(
14
07
19
0<
#20000000
0!
0(
b1 /
04
b1 8
09
#30000000
1!
1(
b1 1
14
17
19
0<
#40000000
0!
0(
b10 /
04
b10 8
09
#50000000
1!
1(
b10 1
14
19
0<
#60000000
0!
0(
b11 /
04
b11 8
09
#70000000
1!
1(
b11 1
14
19
0<
#80000000
0!
0(
b100 /
04
b100 8
09
#90000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b100 1
b0001 3
14
07
19
0<
b1001111 >
b0001 ?
#100000000
0!
0(
b0 /
04
b0 8
09
#110000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
0<
#120000000
0!
0(
b1 /
04
b1 8
09
#130000000
1!
1(
b1 1
14
17
19
0<
#140000000
0!
0(
b10 /
04
b10 8
09
#150000000
1!
1(
b10 1
14
19
0<
#160000000
0!
0(
b11 /
04
b11 8
09
#170000000
1!
1(
b11 1
14
19
0<
#180000000
0!
0(
b100 /
04
b100 8
09
#190000000
1!
1(
b100 1
14
07
19
0<
#200000000
0!
0(
b0 /
04
b0 8
09
#210000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
0<
#220000000
0!
0(
b1 /
04
b1 8
09
#230000000
1!
1(
b1 1
14
17
19
0<
#240000000
0!
0(
b10 /
04
b10 8
09
#250000000
1!
1(
b10 1
14
19
0<
#260000000
0!
0(
b11 /
04
b11 8
09
#270000000
1!
1(
b11 1
14
19
0<
#280000000
0!
0(
b100 /
04
b100 8
09
#290000000
1!
1(
b100 1
14
07
19
0<
#300000000
0!
0(
b0 /
04
b0 8
09
#310000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
0<
#320000000
0!
0(
b1 /
04
b1 8
09
#330000000
1!
1(
b1 1
14
17
19
0<
#340000000
0!
0(
b10 /
04
b10 8
09
#350000000
1!
1(
b10 1
14
19
0<
#360000000
0!
0(
b11 /
04
b11 8
09
#370000000
1!
1(
b11 1
14
19
0<
#380000000
0!
0(
b100 /
04
b100 8
09
#390000000
1!
1(
b100 1
14
07
19
0<
#400000000
0!
0(
b0 /
04
b0 8
09
#410000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
0<
#420000000
0!
0(
b1 /
04
b1 8
09
#430000000
1!
1(
b1 1
14
17
19
0<
#440000000
0!
0(
b10 /
04
b10 8
09
#450000000
1!
1(
b10 1
14
19
0<
#460000000
0!
0(
b11 /
04
b11 8
09
#470000000
1!
1(
b11 1
14
19
0<
#480000000
0!
0(
b100 /
04
b100 8
09
#490000000
1!
1$
1(
1+
b1 0
b0 1
14
07
19
0<
#500000000
0!
0(
b0 /
04
b0 8
09
#510000000
1!
b0011 '
1(
b0011 .
14
19
0<
#520000000
0!
0(
b1 /
04
b1 8
09
#530000000
1!
b0001 '
1(
b0001 .
14
17
19
0<
#540000000
0!
0(
b10 /
04
b10 8
09
#550000000
1!
b1001 '
1(
b1001 .
14
19
0<
#560000000
0!
0(
b11 /
04
b11 8
09
#570000000
1!
0$
b1000 '
1(
0+
b1000 .
b101 0
b11 1
14
19
0<
#580000000
0!
0(
b100 /
04
b100 8
09
#590000000
1!
1(
b100 1
14
07
19
0<
#600000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b0 /
b0000 3
04
b0 8
09
b0000001 >
b0000 ?
#610000000
1!
1(
b0 1
14
19
0<
#620000000
0!
0(
b1 /
04
b1 8
09
#630000000
1!
1(
b1 1
14
17
19
0<
#640000000
0!
0(
b10 /
04
b10 8
09
#650000000
1!
1(
b10 1
14
19
0<
#660000000
0!
0(
b11 /
04
b11 8
09
#670000000
1!
1(
b11 1
14
19
0<
#680000000
0!
0(
b100 /
04
b100 8
09
#690000000
1!
1(
b100 1
14
07
19
0<
#700000000
0!
0(
b0 /
04
b0 8
09
#710000000
1!
1(
b0 1
14
19
0<
#720000000
0!
0(
b1 /
04
b1 8
09
#730000000
1!
1(
b1 1
14
17
19
0<
#740000000
0!
0(
b10 /
04
b10 8
09
#750000000
1!
1(
b10 1
14
19
0<
#760000000
0!
0(
b11 /
04
b11 8
09
#770000000
1!
1#
b0010010 &
1(
1*
b0010010 -
b11 1
b0010 3
14
19
0<
b0010010 >
b0010 ?
#780000000
0!
0(
b100 /
04
b100 8
09
#790000000
1!
1(
b100 1
14
07
19
0<
#800000000
0!
0(
b0 /
04
b0 8
09
#810000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
0<
#820000000
0!
0(
b1 /
04
b1 8
09
#830000000
1!
1(
b1 1
14
17
19
0<
#840000000
0!
0(
b10 /
04
b10 8
09
#850000000
1!
1(
b10 1
14
19
0<
#860000000
0!
0(
b11 /
04
b11 8
09
#870000000
1!
1(
b11 1
14
19
0<
#880000000
0!
0(
b100 /
04
b100 8
09
#890000000
1!
1(
b100 1
14
07
19
0<
#900000000
0!
0(
b0 /
04
b0 8
09
#910000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
0<
#920000000
0!
0(
b1 /
04
b1 8
09
#930000000
1!
1(
b1 1
14
17
19
0<
#940000000
0!
0(
b10 /
04
b10 8
09
#950000000
1!
1(
b10 1
14
19
0<
#960000000
0!
0(
b11 /
04
b11 8
09
#970000000
1!
1(
b11 1
14
19
0<
#980000000
0!
0(
b100 /
04
b100 8
09
#990000000
1!
1(
b100 1
14
07
19
0<
#1000000000
0!
0(
b0 /
04
b0 8
09
#1010000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
0<
#1020000000
0!
0(
b1 /
04
b1 8
09
#1030000000
1!
1(
b1 1
14
17
19
0<
#1040000000
0!
0(
b10 /
04
b10 8
09
#1050000000
1!
1(
b10 1
14
19
0<
#1060000000
0!
0(
b11 /
04
b11 8
09
#1070000000
1!
1(
b11 1
14
19
0<
#1080000000
0!
0(
b100 /
04
b100 8
09
#1090000000
1!
1(
b100 1
14
07
19
0<
#1100000000
0!
0(
b0 /
04
b0 8
09
#1110000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
0<
#1120000000
0!
0(
b1 /
04
b1 8
09
#1130000000
1!
1(
b1 1
14
17
19
0<
#1140000000
0!
0(
b10 /
04
b10 8
09
#1150000000
1!
1(
b10 1
14
19
0<
#1160000000
0!
0(
b11 /
04
b11 8
09
#1170000000
1!
1(
b11 1
14
19
0<
#1180000000
0!
0(
b100 /
04
b100 8
09
#1190000000
1!
1(
b100 1
14
07
19
0<
#1200000000
0!
1$
0(
1+
b0 /
b1 0
b0 1
04
b0 8
09
#1210000000
1!
b0110 '
1(
b0110 .
14
19
0<
#1220000000
0!
0(
b1 /
04
b1 8
09
#1230000000
1!
b0100 '
1(
b0100 .
14
17
19
0<
#1240000000
0!
0(
b10 /
04
b10 8
09
#1250000000
1!
0$
b1100 '
1(
0+
b1100 .
b101 0
b10 1
14
19
0<
#1260000000
0!
0(
b11 /
04
b11 8
09
#1270000000
1!
1(
b11 1
14
19
0<
#1280000000
0!
0#
b0000001 &
0(
0*
b0000001 -
b100 /
b0000 3
04
b100 8
09
b0000001 >
b0000 ?
#1290000000
1!
1(
b100 1
14
07
19
0<
#1300000000
0!
0(
b0 /
04
b0 8
09
#1310000000
1!
1(
b0 1
14
19
0<
#1320000000
0!
0(
b1 /
04
b1 8
09
#1330000000
1!
1(
b1 1
14
17
19
0<
#1340000000
0!
0(
b10 /
04
b10 8
09
#1350000000
1!
1(
b10 1
14
19
0<
#1360000000
0!
0(
b11 /
04
b11 8
09
#1370000000
1!
1(
b11 1
14
19
0<
#1380000000
0!
0(
b100 /
04
b100 8
09
#1390000000
1!
1(
b100 1
14
07
19
0<
#1400000000
0!
0(
b0 /
04
b0 8
09
#1410000000
1!
1(
b0 1
14
19
0<
#1420000000
0!
0(
b1 /
04
b1 8
09
#1430000000
1!
1(
b1 1
14
17
19
0<
#1440000000
0!
0(
b10 /
04
b10 8
09
#1450000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b10 1
b0001 3
14
19
0<
b1001111 >
b0001 ?
#1460000000
0!
0(
b11 /
04
b11 8
09
#1470000000
1!
1(
b11 1
14
19
0<
#1480000000
0!
0(
b100 /
04
b100 8
09
#1490000000
1!
1(
b100 1
14
07
19
0<
#1500000000
0!
0(
b0 /
04
b0 8
09
#1510000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
0<
#1520000000
0!
0(
b1 /
04
b1 8
09
#1530000000
1!
1(
b1 1
14
17
19
0<
#1540000000
0!
0(
b10 /
04
b10 8
09
#1550000000
1!
1(
b10 1
14
19
0<
#1560000000
0!
0(
b11 /
04
b11 8
09
#1570000000
1!
1(
b11 1
14
19
0<
#1580000000
0!
0(
b100 /
04
b100 8
09
#1590000000
1!
1(
b100 1
14
07
19
0<
#1600000000
0!
0(
b0 /
04
b0 8
09
#1610000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
0<
#1620000000
0!
0(
b1 /
04
b1 8
09
#1630000000
1!
1(
b1 1
14
17
19
0<
#1640000000
0!
0(
b10 /
04
b10 8
09
#1650000000
1!
1(
b10 1
14
19
0<
#1660000000
0!
0(
b11 /
04
b11 8
09
#1670000000
1!
1(
b11 1
14
19
0<
#1680000000
0!
0(
b100 /
04
b100 8
09
#1690000000
1!
1(
b100 1
14
07
19
0<
#1700000000
0!
0(
b0 /
04
b0 8
09
#1710000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
0<
#1720000000
0!
0(
b1 /
04
b1 8
09
#1730000000
1!
1(
b1 1
14
17
19
0<
#1740000000
0!
0(
b10 /
04
b10 8
09
#1750000000
1!
1(
b10 1
14
19
0<
#1760000000
0!
0(
b11 /
04
b11 8
09
#1770000000
1!
1(
b11 1
14
19
0<
#1780000000
0!
0(
b100 /
04
b100 8
09
#1790000000
1!
1(
b100 1
14
07
19
0<
#1800000000
0!
0(
b0 /
04
b0 8
09
#1810000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
0<
#1820000000
0!
0(
b1 /
04
b1 8
09
#1830000000
1!
1(
b1 1
14
17
19
0<
#1840000000
0!
0(
b10 /
04
b10 8
09
#1850000000
1!
1$
1(
1+
b1 0
b0 1
14
19
0<
#1860000000
0!
0(
b11 /
04
b11 8
09
#1870000000
1!
b0001 '
1(
b0001 .
14
19
0<
#1880000000
0!
0(
b100 /
04
b100 8
09
#1890000000
1!
b1001 '
1(
b1001 .
14
07
19
0<
#1900000000
0!
0(
b0 /
04
b0 8
09
#1910000000
1!
b1000 '
1(
b1000 .
14
19
0<
#1920000000
0!
0(
b1 /
04
b1 8
09
#1930000000
1!
0$
b1100 '
1(
0+
b1100 .
b101 0
b1 1
14
17
19
0<
#1940000000
0!
0(
b10 /
04
b10 8
09
#1950000000
1!
1(
b10 1
14
19
0<
#1960000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b11 /
b0000 3
04
b11 8
09
b0000001 >
b0000 ?
#1970000000
1!
1(
b11 1
14
19
0<
#1980000000
0!
0(
b100 /
04
b100 8
09
#1990000000
1!
1(
b100 1
14
07
19
0<
#2000000000
0!
0(
b0 /
04
b0 8
09
#2010000000
1!
1(
b0 1
14
19
0<
#2020000000
0!
0(
b1 /
04
b1 8
09
#2030000000
1!
1(
b1 1
14
17
19
0<
#2040000000
0!
0(
b10 /
04
b10 8
09
#2050000000
1!
1(
b10 1
14
19
0<
#2060000000
0!
0(
b11 /
04
b11 8
09
#2070000000
1!
1(
b11 1
14
19
0<
#2080000000
0!
0(
b100 /
04
b100 8
09
#2090000000
1!
1(
b100 1
14
07
19
0<
#2100000000
0!
0(
b0 /
04
b0 8
09
#2110000000
1!
1(
b0 1
14
19
0<
#2120000000
0!
0(
b1 /
04
b1 8
09
#2130000000
1!
1#
b0010010 &
1(
1*
b0010010 -
b1 1
b0010 3
14
17
19
0<
b0010010 >
b0010 ?
#2140000000
0!
0(
b10 /
04
b10 8
09
#2150000000
1!
1(
b10 1
14
19
0<
#2160000000
0!
0(
b11 /
04
b11 8
09
#2170000000
1!
1(
b11 1
14
19
0<
#2180000000
0!
0(
b100 /
04
b100 8
09
#2190000000
1!
1(
b100 1
14
07
19
0<
#2200000000
0!
0(
b0 /
04
b0 8
09
#2210000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#2220000000
0!
0(
b1 /
04
b1 8
09
#2230000000
1!
1(
b1 1
14
17
19
0<
#2240000000
0!
0(
b10 /
04
b10 8
09
#2250000000
1!
1(
b10 1
14
19
0<
#2260000000
0!
0(
b11 /
04
b11 8
09
#2270000000
1!
1(
b11 1
14
19
0<
#2280000000
0!
0(
b100 /
04
b100 8
09
#2290000000
1!
1(
b100 1
14
07
19
0<
#2300000000
0!
0(
b0 /
04
b0 8
09
#2310000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
0<
#2320000000
0!
0(
b1 /
04
b1 8
09
#2330000000
1!
1(
b1 1
14
17
19
0<
#2340000000
0!
0(
b10 /
04
b10 8
09
#2350000000
1!
1(
b10 1
14
19
0<
#2360000000
0!
0(
b11 /
04
b11 8
09
#2370000000
1!
1(
b11 1
14
19
0<
#2380000000
0!
0(
b100 /
04
b100 8
09
#2390000000
1!
1(
b100 1
14
07
19
0<
#2400000000
0!
0(
b0 /
04
b0 8
09
#2410000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
0<
#2420000000
0!
0(
b1 /
04
b1 8
09
#2430000000
1!
1(
b1 1
14
17
19
0<
#2440000000
0!
0(
b10 /
04
b10 8
09
#2450000000
1!
1(
b10 1
14
19
0<
#2460000000
0!
0(
b11 /
04
b11 8
09
#2470000000
1!
1(
b11 1
14
19
0<
#2480000000
0!
0(
b100 /
04
b100 8
09
#2490000000
1!
1(
b100 1
14
07
19
0<
#2500000000
0!
0(
b0 /
04
b0 8
09
#2510000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
0<
#2520000000
0!
0(
b1 /
04
b1 8
09
#2530000000
1!
1(
b1 1
14
17
19
0<
#2540000000
0!
0(
b10 /
04
b10 8
09
#2550000000
1!
1(
b10 1
14
19
0<
#2560000000
0!
1$
0(
1+
b11 /
b1 0
b0 1
04
b11 8
09
#2570000000
1!
b0010 '
1(
b0010 .
14
19
0<
#2580000000
0!
0(
b100 /
04
b100 8
09
#2590000000
1!
b0110 '
1(
b0110 .
14
07
19
0<
#2600000000
0!
0(
b0 /
04
b0 8
09
#2610000000
1!
0$
b0100 '
1(
0+
b0100 .
b101 0
14
19
0<
#2620000000
0!
0(
b1 /
04
b1 8
09
#2630000000
1!
1(
b1 1
14
17
19
0<
#2640000000
0!
0#
b0000001 &
0(
0*
b0000001 -
b10 /
b0000 3
04
b10 8
09
b0000001 >
b0000 ?
#2650000000
1!
1(
b10 1
14
19
0<
#2660000000
0!
0(
b11 /
04
b11 8
09
#2670000000
1!
1(
b11 1
14
19
0<
#2680000000
0!
0(
b100 /
04
b100 8
09
#2690000000
1!
1(
b100 1
14
07
19
0<
#2700000000
0!
0(
b0 /
04
b0 8
09
#2710000000
1!
1(
b0 1
14
19
0<
#2720000000
0!
0(
b1 /
04
b1 8
09
#2730000000
1!
1(
b1 1
14
17
19
0<
#2740000000
0!
0(
b10 /
04
b10 8
09
#2750000000
1!
1(
b10 1
14
19
0<
#2760000000
0!
0(
b11 /
04
b11 8
09
#2770000000
1!
1(
b11 1
14
19
0<
#2780000000
0!
0(
b100 /
04
b100 8
09
#2790000000
1!
1(
b100 1
14
07
19
0<
#2800000000
0!
0(
b0 /
04
b0 8
09
#2810000000
1!
1"
b1001111 &
b0110 '
1(
1)
b1001111 -
b0110 .
b0 1
b0001 3
14
19
0<
b1001111 >
b0001 ?
#2820000000
0!
0(
b1 /
04
b1 8
09
#2830000000
1!
1(
b1 1
14
17
19
0<
#2840000000
0!
0(
b10 /
04
b10 8
09
#2850000000
1!
1(
b10 1
14
19
0<
#2860000000
0!
0(
b11 /
04
b11 8
09
#2870000000
1!
1(
b11 1
14
19
0<
#2880000000
0!
0(
b100 /
04
b100 8
09
#2890000000
1!
1(
b100 1
14
07
19
0<
#2900000000
0!
0(
b0 /
04
b0 8
09
#2910000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
0<
#2920000000
0!
0(
b1 /
04
b1 8
09
#2930000000
1!
1(
b1 1
14
17
19
0<
#2940000000
0!
0(
b10 /
04
b10 8
09
#2950000000
1!
1(
b10 1
14
19
0<
#2960000000
0!
0(
b11 /
04
b11 8
09
#2970000000
1!
1(
b11 1
14
19
0<
#2980000000
0!
0(
b100 /
04
b100 8
09
#2990000000
1!
1(
b100 1
14
07
19
0<
#3000000000
0!
0(
b0 /
04
b0 8
09
#3010000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
0<
#3020000000
0!
0(
b1 /
04
b1 8
09
#3030000000
1!
1(
b1 1
14
17
19
0<
#3040000000
0!
0(
b10 /
04
b10 8
09
#3050000000
1!
1(
b10 1
14
19
0<
#3060000000
0!
0(
b11 /
04
b11 8
09
#3070000000
1!
1(
b11 1
14
19
0<
#3080000000
0!
0(
b100 /
04
b100 8
09
#3090000000
1!
1(
b100 1
14
07
19
0<
#3100000000
0!
0(
b0 /
04
b0 8
09
#3110000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
0<
#3120000000
0!
0(
b1 /
04
b1 8
09
#3130000000
1!
1(
b1 1
14
17
19
0<
#3140000000
0!
0(
b10 /
04
b10 8
09
#3150000000
1!
1(
b10 1
14
19
0<
#3160000000
0!
0(
b11 /
04
b11 8
09
#3170000000
1!
1(
b11 1
14
19
0<
#3180000000
0!
0(
b100 /
04
b100 8
09
#3190000000
1!
1(
b100 1
14
07
19
0<
#3200000000
0!
0(
b0 /
04
b0 8
09
#3210000000
1!
1$
b1001 '
1(
1+
b1001 .
b1 0
b0 1
14
19
0<
#3220000000
0!
0(
b1 /
04
b1 8
09
#3230000000
1!
b1000 '
1(
b1000 .
14
17
19
0<
#3240000000
0!
0(
b10 /
04
b10 8
09
#3250000000
1!
b1100 '
1(
b1100 .
14
19
0<
#3260000000
0!
0(
b11 /
04
b11 8
09
#3270000000
1!
b0100 '
1(
b0100 .
14
19
0<
#3280000000
0!
0(
b100 /
04
b100 8
09
#3290000000
1!
0$
b0110 '
1(
0+
b0110 .
b101 0
b100 1
14
07
19
0<
#3300000000
0!
0(
b0 /
04
b0 8
09
#3310000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
0<
#3320000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b1 /
b0000 3
04
b1 8
09
b0000001 >
b0000 ?
#3330000000
1!
1(
b1 1
14
17
19
0<
#3340000000
0!
0(
b10 /
04
b10 8
09
#3350000000
1!
1(
b10 1
14
19
0<
#3360000000
0!
0(
b11 /
04
b11 8
09
#3370000000
1!
1(
b11 1
14
19
0<
#3380000000
0!
0(
b100 /
04
b100 8
09
#3390000000
1!
1(
b100 1
14
07
19
0<
#3400000000
0!
0(
b0 /
04
b0 8
09
#3410000000
1!
1(
b0 1
14
19
0<
#3420000000
0!
0(
b1 /
04
b1 8
09
#3430000000
1!
1(
b1 1
14
17
19
0<
#3440000000
0!
0(
b10 /
04
b10 8
09
#3450000000
1!
1(
b10 1
14
19
0<
#3460000000
0!
0(
b11 /
04
b11 8
09
#3470000000
1!
1(
b11 1
14
19
0<
#3480000000
0!
0(
b100 /
04
b100 8
09
#3490000000
1!
1#
b0010010 &
1(
1*
b0010010 -
b100 1
b0010 3
14
07
19
0<
b0010010 >
b0010 ?
#3500000000
0!
0(
b0 /
04
b0 8
09
#3510000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
0<
#3520000000
0!
0(
b1 /
04
b1 8
09
#3530000000
1!
1(
b1 1
14
17
19
0<
#3540000000
0!
0(
b10 /
04
b10 8
09
#3550000000
1!
1(
b10 1
14
19
0<
#3560000000
0!
0(
b11 /
04
b11 8
09
#3570000000
1!
1(
b11 1
14
19
0<
#3580000000
0!
0(
b100 /
04
b100 8
09
#3590000000
1!
1(
b100 1
14
07
19
0<
#3600000000
0!
0(
b0 /
04
b0 8
09
#3610000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
0<
#3620000000
0!
0(
b1 /
04
b1 8
09
#3630000000
1!
1(
b1 1
14
17
19
0<
#3640000000
0!
0(
b10 /
04
b10 8
09
#3650000000
1!
1(
b10 1
14
19
0<
#3660000000
0!
0(
b11 /
04
b11 8
09
#3670000000
1!
1(
b11 1
14
19
0<
#3680000000
0!
0(
b100 /
04
b100 8
09
#3690000000
1!
1(
b100 1
14
07
19
0<
#3700000000
0!
0(
b0 /
04
b0 8
09
#3710000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
0<
#3720000000
0!
0(
b1 /
04
b1 8
09
#3730000000
1!
1(
b1 1
14
17
19
0<
#3740000000
0!
0(
b10 /
04
b10 8
09
#3750000000
1!
1(
b10 1
14
19
0<
#3760000000
0!
0(
b11 /
04
b11 8
09
#3770000000
1!
1(
b11 1
14
19
0<
#3780000000
0!
0(
b100 /
04
b100 8
09
#3790000000
1!
1(
b100 1
14
07
19
0<
#3800000000
0!
0(
b0 /
04
b0 8
09
#3810000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#3820000000
0!
0(
b1 /
04
b1 8
09
#3830000000
1!
1(
b1 1
14
17
19
0<
#3840000000
0!
0(
b10 /
04
b10 8
09
#3850000000
1!
1(
b10 1
14
19
0<
#3860000000
0!
0(
b11 /
04
b11 8
09
#3870000000
1!
1(
b11 1
14
19
0<
#3880000000
0!
0(
b100 /
04
b100 8
09
#3890000000
1!
1(
b100 1
14
07
19
0<
#3900000000
0!
0(
b0 /
04
b0 8
09
#3910000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
0<
#3920000000
0!
1$
0(
1+
b1 /
b1 0
04
b1 8
09
#3930000000
1!
b0001 '
1(
b0001 .
14
17
19
0<
#3940000000
0!
0(
b10 /
04
b10 8
09
#3950000000
1!
b0011 '
1(
b0011 .
14
19
0<
#3960000000
0!
0(
b11 /
04
b11 8
09
#3970000000
1!
0$
b0010 '
1(
0+
b0010 .
b101 0
b11 1
14
19
0<
#3980000000
0!
0(
b100 /
04
b100 8
09
#3990000000
1!
1(
b100 1
14
07
19
0<
#4000000000
0!
0#
b0000001 &
0(
0*
b0000001 -
b0 /
b0000 3
04
b0 8
09
b0000001 >
b0000 ?
#4010000000
1!
1(
b0 1
14
19
0<
#4020000000
0!
0(
b1 /
04
b1 8
09
#4030000000
1!
1(
b1 1
14
17
19
0<
#4040000000
0!
0(
b10 /
04
b10 8
09
#4050000000
1!
1(
b10 1
14
19
0<
#4060000000
0!
0(
b11 /
04
b11 8
09
#4070000000
1!
1(
b11 1
14
19
0<
#4080000000
0!
0(
b100 /
04
b100 8
09
#4090000000
1!
1(
b100 1
14
07
19
0<
#4100000000
0!
0(
b0 /
04
b0 8
09
#4110000000
1!
1(
b0 1
14
19
0<
#4120000000
0!
0(
b1 /
04
b1 8
09
#4130000000
1!
1(
b1 1
14
17
19
0<
#4140000000
0!
0(
b10 /
04
b10 8
09
#4150000000
1!
1(
b10 1
14
19
0<
#4160000000
0!
0(
b11 /
04
b11 8
09
#4170000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b11 1
b0001 3
14
19
0<
b1001111 >
b0001 ?
#4180000000
0!
0(
b100 /
04
b100 8
09
#4190000000
1!
1(
b100 1
14
07
19
0<
#4200000000
0!
0(
b0 /
04
b0 8
09
#4210000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
0<
#4220000000
0!
0(
b1 /
04
b1 8
09
#4230000000
1!
1(
b1 1
14
17
19
0<
#4240000000
0!
0(
b10 /
04
b10 8
09
#4250000000
1!
1(
b10 1
14
19
0<
#4260000000
0!
0(
b11 /
04
b11 8
09
#4270000000
1!
1(
b11 1
14
19
0<
#4280000000
0!
0(
b100 /
04
b100 8
09
#4290000000
1!
1(
b100 1
14
07
19
0<
#4300000000
0!
0(
b0 /
04
b0 8
09
#4310000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
0<
#4320000000
0!
0(
b1 /
04
b1 8
09
#4330000000
1!
1(
b1 1
14
17
19
0<
#4340000000
0!
0(
b10 /
04
b10 8
09
#4350000000
1!
1(
b10 1
14
19
0<
#4360000000
0!
0(
b11 /
04
b11 8
09
#4370000000
1!
1(
b11 1
14
19
0<
#4380000000
0!
0(
b100 /
04
b100 8
09
#4390000000
1!
1(
b100 1
14
07
19
0<
#4400000000
0!
0(
b0 /
04
b0 8
09
#4410000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
0<
#4420000000
0!
0(
b1 /
04
b1 8
09
#4430000000
1!
1(
b1 1
14
17
19
0<
#4440000000
0!
0(
b10 /
04
b10 8
09
#4450000000
1!
1(
b10 1
14
19
0<
#4460000000
0!
0(
b11 /
04
b11 8
09
#4470000000
1!
1(
b11 1
14
19
0<
#4480000000
0!
0(
b100 /
04
b100 8
09
#4490000000
1!
1(
b100 1
14
07
19
0<
#4500000000
0!
0(
b0 /
04
b0 8
09
#4510000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#4520000000
0!
0(
b1 /
04
b1 8
09
#4530000000
1!
1(
b1 1
14
17
19
0<
#4540000000
0!
0(
b10 /
04
b10 8
09
#4550000000
1!
1(
b10 1
14
19
0<
#4560000000
0!
0(
b11 /
04
b11 8
09
#4570000000
1!
1$
1(
1+
b1 0
b0 1
14
19
0<
#4580000000
0!
0(
b100 /
04
b100 8
09
#4590000000
1!
b1100 '
1(
b1100 .
14
07
19
0<
#4600000000
0!
0(
b0 /
04
b0 8
09
#4610000000
1!
b0100 '
1(
b0100 .
14
19
0<
#4620000000
0!
0(
b1 /
04
b1 8
09
#4630000000
1!
b0110 '
1(
b0110 .
14
17
19
0<
#4640000000
0!
0(
b10 /
04
b10 8
09
#4650000000
1!
0$
b0010 '
1(
0+
b0010 .
b101 0
b10 1
14
19
0<
#4660000000
0!
0(
b11 /
04
b11 8
09
#4670000000
1!
1(
b11 1
14
19
0<
#4680000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b100 /
b0000 3
04
b100 8
09
b0000001 >
b0000 ?
#4690000000
1!
1(
b100 1
14
07
19
0<
#4700000000
0!
0(
b0 /
04
b0 8
09
#4710000000
1!
1(
b0 1
14
19
0<
#4720000000
0!
0(
b1 /
04
b1 8
09
#4730000000
1!
1(
b1 1
14
17
19
0<
#4740000000
0!
0(
b10 /
04
b10 8
09
#4750000000
1!
1(
b10 1
14
19
0<
#4760000000
0!
0(
b11 /
04
b11 8
09
#4770000000
1!
1(
b11 1
14
19
0<
#4780000000
0!
0(
b100 /
04
b100 8
09
#4790000000
1!
1(
b100 1
14
07
19
0<
#4800000000
0!
0(
b0 /
04
b0 8
09
#4810000000
1!
1(
b0 1
14
19
0<
#4820000000
0!
0(
b1 /
04
b1 8
09
#4830000000
1!
1(
b1 1
14
17
19
0<
#4840000000
0!
0(
b10 /
04
b10 8
09
#4850000000
1!
1#
b0010010 &
1(
1*
b0010010 -
b10 1
b0010 3
14
19
0<
b0010010 >
b0010 ?
#4860000000
0!
0(
b11 /
04
b11 8
09
#4870000000
1!
1(
b11 1
14
19
0<
#4880000000
0!
0(
b100 /
04
b100 8
09
#4890000000
1!
1(
b100 1
14
07
19
0<
#4900000000
0!
0(
b0 /
04
b0 8
09
#4910000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
0<
#4920000000
0!
0(
b1 /
04
b1 8
09
#4930000000
1!
1(
b1 1
14
17
19
0<
#4940000000
0!
0(
b10 /
04
b10 8
09
#4950000000
1!
1(
b10 1
14
19
0<
#4960000000
0!
0(
b11 /
04
b11 8
09
#4970000000
1!
1(
b11 1
14
19
0<
#4980000000
0!
0(
b100 /
04
b100 8
09
#4990000000
1!
1(
b100 1
14
07
19
0<
#5000000000
0!
0(
b0 /
04
b0 8
09
#5010000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
0<
#5020000000
0!
0(
b1 /
04
b1 8
09
#5030000000
1!
1(
b1 1
14
17
19
0<
#5040000000
0!
0(
b10 /
04
b10 8
09
#5050000000
1!
1(
b10 1
14
19
0<
#5060000000
0!
0(
b11 /
04
b11 8
09
#5070000000
1!
1(
b11 1
14
19
0<
#5080000000
0!
0(
b100 /
04
b100 8
09
#5090000000
1!
1(
b100 1
14
07
19
0<
#5100000000
0!
0(
b0 /
04
b0 8
09
#5110000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
0<
#5120000000
0!
0(
b1 /
04
b1 8
09
#5130000000
1!
1(
b1 1
14
17
19
0<
#5140000000
0!
0(
b10 /
04
b10 8
09
#5150000000
1!
1(
b10 1
14
19
0<
#5160000000
0!
0(
b11 /
04
b11 8
09
#5170000000
1!
1(
b11 1
14
19
0<
#5180000000
0!
0(
b100 /
04
b100 8
09
#5190000000
1!
1(
b100 1
14
07
19
0<
#5200000000
0!
0(
b0 /
04
b0 8
09
#5210000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#5220000000
0!
0(
b1 /
04
b1 8
09
#5230000000
1!
1(
b1 1
14
17
19
0<
#5240000000
0!
0(
b10 /
04
b10 8
09
#5250000000
1!
1(
b10 1
14
19
0<
#5260000000
0!
0(
b11 /
04
b11 8
09
#5270000000
1!
1(
b11 1
14
19
0<
#5280000000
0!
1$
0(
1+
b100 /
b1 0
b0 1
04
b100 8
09
#5290000000
1!
b1001 '
1(
b1001 .
14
07
19
0<
#5300000000
0!
0(
b0 /
04
b0 8
09
#5310000000
1!
b0001 '
1(
b0001 .
14
19
0<
#5320000000
0!
0(
b1 /
04
b1 8
09
#5330000000
1!
0$
b0011 '
1(
0+
b0011 .
b101 0
b1 1
14
17
19
0<
#5340000000
0!
0(
b10 /
04
b10 8
09
#5350000000
1!
1(
b10 1
14
19
0<
#5360000000
0!
0#
b0000001 &
0(
0*
b0000001 -
b11 /
b0000 3
04
b11 8
09
b0000001 >
b0000 ?
#5370000000
1!
1(
b11 1
14
19
0<
#5380000000
0!
0(
b100 /
04
b100 8
09
#5390000000
1!
1(
b100 1
14
07
19
0<
#5400000000
0!
0(
b0 /
04
b0 8
09
#5410000000
1!
1(
b0 1
14
19
0<
#5420000000
0!
0(
b1 /
04
b1 8
09
#5430000000
1!
1(
b1 1
14
17
19
0<
#5440000000
0!
0(
b10 /
04
b10 8
09
#5450000000
1!
1(
b10 1
14
19
0<
#5460000000
0!
0(
b11 /
04
b11 8
09
#5470000000
1!
1(
b11 1
14
19
0<
#5480000000
0!
0(
b100 /
04
b100 8
09
#5490000000
1!
1(
b100 1
14
07
19
0<
#5500000000
0!
0(
b0 /
04
b0 8
09
#5510000000
1!
1(
b0 1
14
19
0<
#5520000000
0!
0(
b1 /
04
b1 8
09
#5530000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b1 1
b0001 3
14
17
19
0<
b1001111 >
b0001 ?
#5540000000
0!
0(
b10 /
04
b10 8
09
#5550000000
1!
1(
b10 1
14
19
0<
#5560000000
0!
0(
b11 /
04
b11 8
09
#5570000000
1!
1(
b11 1
14
19
0<
#5580000000
0!
0(
b100 /
04
b100 8
09
#5590000000
1!
1(
b100 1
14
07
19
0<
#5600000000
0!
0(
b0 /
04
b0 8
09
#5610000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
0<
#5620000000
0!
0(
b1 /
04
b1 8
09
#5630000000
1!
1(
b1 1
14
17
19
0<
#5640000000
0!
0(
b10 /
04
b10 8
09
#5650000000
1!
1(
b10 1
14
19
0<
#5660000000
0!
0(
b11 /
04
b11 8
09
#5670000000
1!
1(
b11 1
14
19
0<
#5680000000
0!
0(
b100 /
04
b100 8
09
#5690000000
1!
1(
b100 1
14
07
19
0<
#5700000000
0!
0(
b0 /
04
b0 8
09
#5710000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
0<
#5720000000
0!
0(
b1 /
04
b1 8
09
#5730000000
1!
1(
b1 1
14
17
19
0<
#5740000000
0!
0(
b10 /
04
b10 8
09
#5750000000
1!
1(
b10 1
14
19
0<
#5760000000
0!
0(
b11 /
04
b11 8
09
#5770000000
1!
1(
b11 1
14
19
0<
#5780000000
0!
0(
b100 /
04
b100 8
09
#5790000000
1!
1(
b100 1
14
07
19
0<
#5800000000
0!
0(
b0 /
04
b0 8
09
#5810000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#5820000000
0!
0(
b1 /
04
b1 8
09
#5830000000
1!
1(
b1 1
14
17
19
0<
#5840000000
0!
0(
b10 /
04
b10 8
09
#5850000000
1!
1(
b10 1
14
19
0<
#5860000000
0!
0(
b11 /
04
b11 8
09
#5870000000
1!
1(
b11 1
14
19
0<
#5880000000
0!
0(
b100 /
04
b100 8
09
#5890000000
1!
1(
b100 1
14
07
19
0<
#5900000000
0!
0(
b0 /
04
b0 8
09
#5910000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
0<
#5920000000
0!
0(
b1 /
04
b1 8
09
#5930000000
1!
1$
1(
1+
b1 0
14
17
19
0<
#5940000000
0!
0(
b10 /
04
b10 8
09
#5950000000
1!
b0100 '
1(
b0100 .
14
19
0<
#5960000000
0!
0(
b11 /
04
b11 8
09
#5970000000
1!
b0110 '
1(
b0110 .
14
19
0<
#5980000000
0!
0(
b100 /
04
b100 8
09
#5990000000
1!
b0010 '
1(
b0010 .
14
07
19
0<
#6000000000
0!
0(
b0 /
04
b0 8
09
#6010000000
1!
0$
b0011 '
1(
0+
b0011 .
b101 0
14
19
0<
#6020000000
0!
0(
b1 /
04
b1 8
09
#6030000000
1!
1(
b1 1
14
17
19
0<
#6040000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b10 /
b0000 3
04
b10 8
09
b0000001 >
b0000 ?
#6050000000
1!
1(
b10 1
14
19
0<
#6060000000
0!
0(
b11 /
04
b11 8
09
#6070000000
1!
1(
b11 1
14
19
0<
#6080000000
0!
0(
b100 /
04
b100 8
09
#6090000000
1!
1(
b100 1
14
07
19
0<
#6100000000
0!
0(
b0 /
04
b0 8
09
#6110000000
1!
1(
b0 1
14
19
0<
#6120000000
0!
0(
b1 /
04
b1 8
09
#6130000000
1!
1(
b1 1
14
17
19
0<
#6140000000
0!
0(
b10 /
04
b10 8
09
#6150000000
1!
1(
b10 1
14
19
0<
#6160000000
0!
0(
b11 /
04
b11 8
09
#6170000000
1!
1(
b11 1
14
19
0<
#6180000000
0!
0(
b100 /
04
b100 8
09
#6190000000
1!
1(
b100 1
14
07
19
0<
#6200000000
0!
0(
b0 /
04
b0 8
09
#6210000000
1!
1#
b0010010 &
b0010 '
1(
1*
b0010010 -
b0010 .
b0 1
b0010 3
14
19
0<
b0010010 >
b0010 ?
#6220000000
0!
0(
b1 /
04
b1 8
09
#6230000000
1!
1(
b1 1
14
17
19
0<
#6240000000
0!
0(
b10 /
04
b10 8
09
#6250000000
1!
1(
b10 1
14
19
0<
#6260000000
0!
0(
b11 /
04
b11 8
09
#6270000000
1!
1(
b11 1
14
19
0<
#6280000000
0!
0(
b100 /
04
b100 8
09
#6290000000
1!
1(
b100 1
14
07
19
0<
#6300000000
0!
0(
b0 /
04
b0 8
09
#6310000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
0<
#6320000000
0!
0(
b1 /
04
b1 8
09
#6330000000
1!
1(
b1 1
14
17
19
0<
#6340000000
0!
0(
b10 /
04
b10 8
09
#6350000000
1!
1(
b10 1
14
19
0<
#6360000000
0!
0(
b11 /
04
b11 8
09
#6370000000
1!
1(
b11 1
14
19
0<
#6380000000
0!
0(
b100 /
04
b100 8
09
#6390000000
1!
1(
b100 1
14
07
19
0<
#6400000000
0!
0(
b0 /
04
b0 8
09
#6410000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
0<
#6420000000
0!
0(
b1 /
04
b1 8
09
#6430000000
1!
1(
b1 1
14
17
19
0<
#6440000000
0!
0(
b10 /
04
b10 8
09
#6450000000
1!
1(
b10 1
14
19
0<
#6460000000
0!
0(
b11 /
04
b11 8
09
#6470000000
1!
1(
b11 1
14
19
0<
#6480000000
0!
0(
b100 /
04
b100 8
09
#6490000000
1!
1(
b100 1
14
07
19
0<
#6500000000
0!
0(
b0 /
04
b0 8
09
#6510000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
0<
#6520000000
0!
0(
b1 /
04
b1 8
09
#6530000000
1!
1(
b1 1
14
17
19
0<
#6540000000
0!
0(
b10 /
04
b10 8
09
#6550000000
1!
1(
b10 1
14
19
0<
#6560000000
0!
0(
b11 /
04
b11 8
09
#6570000000
1!
1(
b11 1
14
19
0<
#6580000000
0!
0(
b100 /
04
b100 8
09
#6590000000
1!
1(
b100 1
14
07
19
0<
#6600000000
0!
0(
b0 /
04
b0 8
09
#6610000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#6620000000
0!
0(
b1 /
04
b1 8
09
#6630000000
1!
1(
b1 1
14
17
19
0<
#6640000000
0!
1$
0(
1+
b10 /
b1 0
b0 1
04
b10 8
09
#6650000000
1!
b1001 '
1(
b1001 .
14
19
0<
#6660000000
0!
0(
b11 /
04
b11 8
09
#6670000000
1!
b0001 '
1(
b0001 .
14
19
0<
#6680000000
0!
0(
b100 /
04
b100 8
09
#6690000000
1!
0$
b0011 '
1(
0+
b0011 .
b101 0
b100 1
14
07
19
0<
#6700000000
0!
0(
b0 /
04
b0 8
09
#6710000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
0<
#6720000000
0!
0#
b0000001 &
0(
0*
b0000001 -
b1 /
b0000 3
04
b1 8
09
b0000001 >
b0000 ?
#6730000000
1!
1(
b1 1
14
17
19
0<
#6740000000
0!
0(
b10 /
04
b10 8
09
#6750000000
1!
1(
b10 1
14
19
0<
#6760000000
0!
0(
b11 /
04
b11 8
09
#6770000000
1!
1(
b11 1
14
19
0<
#6780000000
0!
0(
b100 /
04
b100 8
09
#6790000000
1!
1(
b100 1
14
07
19
0<
#6800000000
0!
0(
b0 /
04
b0 8
09
#6810000000
1!
1(
b0 1
14
19
0<
#6820000000
0!
0(
b1 /
04
b1 8
09
#6830000000
1!
1(
b1 1
14
17
19
0<
#6840000000
0!
0(
b10 /
04
b10 8
09
#6850000000
1!
1(
b10 1
14
19
0<
#6860000000
0!
0(
b11 /
04
b11 8
09
#6870000000
1!
1(
b11 1
14
19
0<
#6880000000
0!
0(
b100 /
04
b100 8
09
#6890000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b100 1
b0001 3
14
07
19
0<
b1001111 >
b0001 ?
#6900000000
0!
0(
b0 /
04
b0 8
09
#6910000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
0<
#6920000000
0!
0(
b1 /
04
b1 8
09
#6930000000
1!
1(
b1 1
14
17
19
0<
#6940000000
0!
0(
b10 /
04
b10 8
09
#6950000000
1!
1(
b10 1
14
19
0<
#6960000000
0!
0(
b11 /
04
b11 8
09
#6970000000
1!
1(
b11 1
14
19
0<
#6980000000
0!
0(
b100 /
04
b100 8
09
#6990000000
1!
1(
b100 1
14
07
19
0<
#7000000000
0!
0(
b0 /
04
b0 8
09
#7010000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
0<
#7020000000
0!
0(
b1 /
04
b1 8
09
#7030000000
1!
1(
b1 1
14
17
19
0<
#7040000000
0!
0(
b10 /
04
b10 8
09
#7050000000
1!
1(
b10 1
14
19
0<
#7060000000
0!
0(
b11 /
04
b11 8
09
#7070000000
1!
1(
b11 1
14
19
0<
#7080000000
0!
0(
b100 /
04
b100 8
09
#7090000000
1!
1(
b100 1
14
07
19
0<
#7100000000
0!
0(
b0 /
04
b0 8
09
#7110000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
0<
#7120000000
0!
0(
b1 /
04
b1 8
09
#7130000000
1!
1(
b1 1
14
17
19
0<
#7140000000
0!
0(
b10 /
04
b10 8
09
#7150000000
1!
1(
b10 1
14
19
0<
#7160000000
0!
0(
b11 /
04
b11 8
09
#7170000000
1!
1(
b11 1
14
19
0<
#7180000000
0!
0(
b100 /
04
b100 8
09
#7190000000
1!
1(
b100 1
14
07
19
0<
#7200000000
0!
0(
b0 /
04
b0 8
09
#7210000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#7220000000
0!
0(
b1 /
04
b1 8
09
#7230000000
1!
1(
b1 1
14
17
19
0<
#7240000000
0!
0(
b10 /
04
b10 8
09
#7250000000
1!
1(
b10 1
14
19
0<
#7260000000
0!
0(
b11 /
04
b11 8
09
#7270000000
1!
1(
b11 1
14
19
0<
#7280000000
0!
0(
b100 /
04
b100 8
09
#7290000000
1!
1$
1(
1+
b1 0
b0 1
14
07
19
0<
#7300000000
0!
0(
b0 /
04
b0 8
09
#7310000000
1!
b1100 '
1(
b1100 .
14
19
0<
#7320000000
0!
0(
b1 /
04
b1 8
09
#7330000000
1!
b0100 '
1(
b0100 .
14
17
19
0<
#7340000000
0!
0(
b10 /
04
b10 8
09
#7350000000
1!
b0110 '
1(
b0110 .
14
19
0<
#7360000000
0!
0(
b11 /
04
b11 8
09
#7370000000
1!
0$
b0010 '
1(
0+
b0010 .
b101 0
b11 1
14
19
0<
#7380000000
0!
0(
b100 /
04
b100 8
09
#7390000000
1!
1(
b100 1
14
07
19
0<
#7400000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b0 /
b0000 3
04
b0 8
09
b0000001 >
b0000 ?
#7410000000
1!
1(
b0 1
14
19
0<
#7420000000
0!
0(
b1 /
04
b1 8
09
#7430000000
1!
1(
b1 1
14
17
19
0<
#7440000000
0!
0(
b10 /
04
b10 8
09
#7450000000
1!
1(
b10 1
14
19
0<
#7460000000
0!
0(
b11 /
04
b11 8
09
#7470000000
1!
1(
b11 1
14
19
0<
#7480000000
0!
0(
b100 /
04
b100 8
09
#7490000000
1!
1(
b100 1
14
07
19
0<
#7500000000
0!
0(
b0 /
04
b0 8
09
#7510000000
1!
1(
b0 1
14
19
0<
#7520000000
0!
0(
b1 /
04
b1 8
09
#7530000000
1!
1(
b1 1
14
17
19
0<
#7540000000
0!
0(
b10 /
04
b10 8
09
#7550000000
1!
1(
b10 1
14
19
0<
#7560000000
0!
0(
b11 /
04
b11 8
09
#7570000000
1!
1#
b0010010 &
1(
1*
b0010010 -
b11 1
b0010 3
14
19
0<
b0010010 >
b0010 ?
#7580000000
0!
0(
b100 /
04
b100 8
09
#7590000000
1!
1(
b100 1
14
07
19
0<
#7600000000
0!
0(
b0 /
04
b0 8
09
#7610000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
0<
#7620000000
0!
0(
b1 /
04
b1 8
09
#7630000000
1!
1(
b1 1
14
17
19
0<
#7640000000
0!
0(
b10 /
04
b10 8
09
#7650000000
1!
1(
b10 1
14
19
0<
#7660000000
0!
0(
b11 /
04
b11 8
09
#7670000000
1!
1(
b11 1
14
19
0<
#7680000000
0!
0(
b100 /
04
b100 8
09
#7690000000
1!
1(
b100 1
14
07
19
0<
#7700000000
0!
0(
b0 /
04
b0 8
09
#7710000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
0<
#7720000000
0!
0(
b1 /
04
b1 8
09
#7730000000
1!
1(
b1 1
14
17
19
0<
#7740000000
0!
0(
b10 /
04
b10 8
09
#7750000000
1!
1(
b10 1
14
19
0<
#7760000000
0!
0(
b11 /
04
b11 8
09
#7770000000
1!
1(
b11 1
14
19
0<
#7780000000
0!
0(
b100 /
04
b100 8
09
#7790000000
1!
1(
b100 1
14
07
19
0<
#7800000000
0!
0(
b0 /
04
b0 8
09
#7810000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
0<
#7820000000
0!
0(
b1 /
04
b1 8
09
#7830000000
1!
1(
b1 1
14
17
19
0<
#7840000000
0!
0(
b10 /
04
b10 8
09
#7850000000
1!
1(
b10 1
14
19
0<
#7860000000
0!
0(
b11 /
04
b11 8
09
#7870000000
1!
1(
b11 1
14
19
0<
#7880000000
0!
0(
b100 /
04
b100 8
09
#7890000000
1!
1(
b100 1
14
07
19
0<
#7900000000
0!
0(
b0 /
04
b0 8
09
#7910000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#7920000000
0!
0(
b1 /
04
b1 8
09
#7930000000
1!
1(
b1 1
14
17
19
0<
#7940000000
0!
0(
b10 /
04
b10 8
09
#7950000000
1!
1(
b10 1
14
19
0<
#7960000000
0!
0(
b11 /
04
b11 8
09
#7970000000
1!
1(
b11 1
14
19
0<
#7980000000
0!
0(
b100 /
04
b100 8
09
#7990000000
1!
1(
b100 1
14
07
19
0<
#8000000000
0!
1$
0(
1+
b0 /
b1 0
b0 1
04
b0 8
09
#8010000000
1!
b1001 '
1(
b1001 .
14
19
0<
#8020000000
0!
0(
b1 /
04
b1 8
09
#8030000000
1!
b0001 '
1(
b0001 .
14
17
19
0<
#8040000000
0!
0(
b10 /
04
b10 8
09
#8050000000
1!
0$
b0011 '
1(
0+
b0011 .
b101 0
b10 1
14
19
0<
#8060000000
0!
0(
b11 /
04
b11 8
09
#8070000000
1!
1(
b11 1
14
19
0<
#8080000000
0!
0#
b0000001 &
0(
0*
b0000001 -
b100 /
b0000 3
04
b100 8
09
b0000001 >
b0000 ?
#8090000000
1!
1(
b100 1
14
07
19
0<
#8100000000
0!
0(
b0 /
04
b0 8
09
#8110000000
1!
1(
b0 1
14
19
0<
#8120000000
0!
0(
b1 /
04
b1 8
09
#8130000000
1!
1(
b1 1
14
17
19
0<
#8140000000
0!
0(
b10 /
04
b10 8
09
#8150000000
1!
1(
b10 1
14
19
0<
#8160000000
0!
0(
b11 /
04
b11 8
09
#8170000000
1!
1(
b11 1
14
19
0<
#8180000000
0!
0(
b100 /
04
b100 8
09
#8190000000
1!
1(
b100 1
14
07
19
0<
#8200000000
0!
0(
b0 /
04
b0 8
09
#8210000000
1!
1(
b0 1
14
19
0<
#8220000000
0!
0(
b1 /
04
b1 8
09
#8230000000
1!
1(
b1 1
14
17
19
0<
#8240000000
0!
0(
b10 /
04
b10 8
09
#8250000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b10 1
b0001 3
14
19
0<
b1001111 >
b0001 ?
#8260000000
0!
0(
b11 /
04
b11 8
09
#8270000000
1!
1(
b11 1
14
19
0<
#8280000000
0!
0(
b100 /
04
b100 8
09
#8290000000
1!
1(
b100 1
14
07
19
0<
#8300000000
0!
0(
b0 /
04
b0 8
09
#8310000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
0<
#8320000000
0!
0(
b1 /
04
b1 8
09
#8330000000
1!
1(
b1 1
14
17
19
0<
#8340000000
0!
0(
b10 /
04
b10 8
09
#8350000000
1!
1(
b10 1
14
19
0<
#8360000000
0!
0(
b11 /
04
b11 8
09
#8370000000
1!
1(
b11 1
14
19
0<
#8380000000
0!
0(
b100 /
04
b100 8
09
#8390000000
1!
1(
b100 1
14
07
19
0<
#8400000000
0!
0(
b0 /
04
b0 8
09
#8410000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
0<
#8420000000
0!
0(
b1 /
04
b1 8
09
#8430000000
1!
1(
b1 1
14
17
19
0<
#8440000000
0!
0(
b10 /
04
b10 8
09
#8450000000
1!
1(
b10 1
14
19
0<
#8460000000
0!
0(
b11 /
04
b11 8
09
#8470000000
1!
1(
b11 1
14
19
0<
#8480000000
0!
0(
b100 /
04
b100 8
09
#8490000000
1!
1(
b100 1
14
07
19
0<
#8500000000
0!
0(
b0 /
04
b0 8
09
#8510000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#8520000000
0!
0(
b1 /
04
b1 8
09
#8530000000
1!
1(
b1 1
14
17
19
0<
#8540000000
0!
0(
b10 /
04
b10 8
09
#8550000000
1!
1(
b10 1
14
19
0<
#8560000000
0!
0(
b11 /
04
b11 8
09
#8570000000
1!
1(
b11 1
14
19
0<
#8580000000
0!
0(
b100 /
04
b100 8
09
#8590000000
1!
1(
b100 1
14
07
19
0<
#8600000000
0!
0(
b0 /
04
b0 8
09
#8610000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
0<
#8620000000
0!
0(
b1 /
04
b1 8
09
#8630000000
1!
1(
b1 1
14
17
19
0<
#8640000000
0!
0(
b10 /
04
b10 8
09
#8650000000
1!
1$
1(
1+
b1 0
b0 1
14
19
0<
#8660000000
0!
0(
b11 /
04
b11 8
09
#8670000000
1!
b0100 '
1(
b0100 .
14
19
0<
#8680000000
0!
0(
b100 /
04
b100 8
09
#8690000000
1!
b0110 '
1(
b0110 .
14
07
19
0<
#8700000000
0!
0(
b0 /
04
b0 8
09
#8710000000
1!
b0010 '
1(
b0010 .
14
19
0<
#8720000000
0!
0(
b1 /
04
b1 8
09
#8730000000
1!
0$
b0011 '
1(
0+
b0011 .
b101 0
b1 1
14
17
19
0<
#8740000000
0!
0(
b10 /
04
b10 8
09
#8750000000
1!
1(
b10 1
14
19
0<
#8760000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b11 /
b0000 3
04
b11 8
09
b0000001 >
b0000 ?
#8770000000
1!
1(
b11 1
14
19
0<
#8780000000
0!
0(
b100 /
04
b100 8
09
#8790000000
1!
1(
b100 1
14
07
19
0<
#8800000000
0!
0(
b0 /
04
b0 8
09
#8810000000
1!
1(
b0 1
14
19
0<
#8820000000
0!
0(
b1 /
04
b1 8
09
#8830000000
1!
1(
b1 1
14
17
19
0<
#8840000000
0!
0(
b10 /
04
b10 8
09
#8850000000
1!
1(
b10 1
14
19
0<
#8860000000
0!
0(
b11 /
04
b11 8
09
#8870000000
1!
1(
b11 1
14
19
0<
#8880000000
0!
0(
b100 /
04
b100 8
09
#8890000000
1!
1(
b100 1
14
07
19
0<
#8900000000
0!
0(
b0 /
04
b0 8
09
#8910000000
1!
1(
b0 1
14
19
0<
#8920000000
0!
0(
b1 /
04
b1 8
09
#8930000000
1!
1#
b0010010 &
1(
1*
b0010010 -
b1 1
b0010 3
14
17
19
0<
b0010010 >
b0010 ?
#8940000000
0!
0(
b10 /
04
b10 8
09
#8950000000
1!
1(
b10 1
14
19
0<
#8960000000
0!
0(
b11 /
04
b11 8
09
#8970000000
1!
1(
b11 1
14
19
0<
#8980000000
0!
0(
b100 /
04
b100 8
09
#8990000000
1!
1(
b100 1
14
07
19
0<
#9000000000
0!
0(
b0 /
04
b0 8
09
#9010000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
0<
#9020000000
0!
0(
b1 /
04
b1 8
09
#9030000000
1!
1(
b1 1
14
17
19
0<
#9040000000
0!
0(
b10 /
04
b10 8
09
#9050000000
1!
1(
b10 1
14
19
0<
#9060000000
0!
0(
b11 /
04
b11 8
09
#9070000000
1!
1(
b11 1
14
19
0<
#9080000000
0!
0(
b100 /
04
b100 8
09
#9090000000
1!
1(
b100 1
14
07
19
0<
#9100000000
0!
0(
b0 /
04
b0 8
09
#9110000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
0<
#9120000000
0!
0(
b1 /
04
b1 8
09
#9130000000
1!
1(
b1 1
14
17
19
0<
#9140000000
0!
0(
b10 /
04
b10 8
09
#9150000000
1!
1(
b10 1
14
19
0<
#9160000000
0!
0(
b11 /
04
b11 8
09
#9170000000
1!
1(
b11 1
14
19
0<
#9180000000
0!
0(
b100 /
04
b100 8
09
#9190000000
1!
1(
b100 1
14
07
19
0<
#9200000000
0!
0(
b0 /
04
b0 8
09
#9210000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
0<
#9220000000
0!
0(
b1 /
04
b1 8
09
#9230000000
1!
1(
b1 1
14
17
19
0<
#9240000000
0!
0(
b10 /
04
b10 8
09
#9250000000
1!
1(
b10 1
14
19
0<
#9260000000
0!
0(
b11 /
04
b11 8
09
#9270000000
1!
1(
b11 1
14
19
0<
#9280000000
0!
0(
b100 /
04
b100 8
09
#9290000000
1!
1(
b100 1
14
07
19
0<
#9300000000
0!
0(
b0 /
04
b0 8
09
#9310000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
0<
#9320000000
0!
0(
b1 /
04
b1 8
09
#9330000000
1!
1(
b1 1
14
17
19
0<
#9340000000
0!
0(
b10 /
04
b10 8
09
#9350000000
1!
1(
b10 1
14
19
0<
#9360000000
0!
1$
0(
1+
b11 /
b1 0
b0 1
04
b11 8
09
#9370000000
1!
b1000 '
1(
b1000 .
14
19
0<
#9380000000
0!
0(
b100 /
04
b100 8
09
#9390000000
1!
b1001 '
1(
b1001 .
14
07
19
0<
#9400000000
0!
0(
b0 /
04
b0 8
09
#9410000000
1!
0$
b0001 '
1(
0+
b0001 .
b101 0
14
19
0<
#9420000000
0!
0(
b1 /
04
b1 8
09
#9430000000
1!
1(
b1 1
14
17
19
0<
#9440000000
0!
0#
b0000001 &
0(
0*
b0000001 -
b10 /
b0000 3
04
b10 8
09
b0000001 >
b0000 ?
#9450000000
1!
1(
b10 1
14
19
0<
#9460000000
0!
0(
b11 /
04
b11 8
09
#9470000000
1!
1(
b11 1
14
19
0<
#9480000000
0!
0(
b100 /
04
b100 8
09
#9490000000
1!
1(
b100 1
14
07
19
0<
#9500000000
0!
0(
b0 /
04
b0 8
09
#9510000000
1!
1(
b0 1
14
19
0<
#9520000000
0!
0(
b1 /
04
b1 8
09
#9530000000
1!
1(
b1 1
14
17
19
0<
#9540000000
0!
0(
b10 /
04
b10 8
09
#9550000000
1!
1(
b10 1
14
19
0<
#9560000000
0!
0(
b11 /
04
b11 8
09
#9570000000
1!
1(
b11 1
14
19
0<
#9580000000
0!
0(
b100 /
04
b100 8
09
#9590000000
1!
1(
b100 1
14
07
19
0<
#9600000000
0!
0(
b0 /
04
b0 8
09
#9610000000
1!
1"
b1001111 &
b1001 '
1(
1)
b1001111 -
b1001 .
b0 1
b0001 3
14
19
0<
b1001111 >
b0001 ?
#9620000000
0!
0(
b1 /
04
b1 8
09
#9630000000
1!
1(
b1 1
14
17
19
0<
#9640000000
0!
0(
b10 /
04
b10 8
09
#9650000000
1!
1(
b10 1
14
19
0<
#9660000000
0!
0(
b11 /
04
b11 8
09
#9670000000
1!
1(
b11 1
14
19
0<
#9680000000
0!
0(
b100 /
04
b100 8
09
#9690000000
1!
1(
b100 1
14
07
19
0<
#9700000000
0!
0(
b0 /
04
b0 8
09
#9710000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
0<
#9720000000
0!
0(
b1 /
04
b1 8
09
#9730000000
1!
1(
b1 1
14
17
19
0<
#9740000000
0!
0(
b10 /
04
b10 8
09
#9750000000
1!
1(
b10 1
14
19
0<
#9760000000
0!
0(
b11 /
04
b11 8
09
#9770000000
1!
1(
b11 1
14
19
0<
#9780000000
0!
0(
b100 /
04
b100 8
09
#9790000000
1!
1(
b100 1
14
07
19
0<
#9800000000
0!
0(
b0 /
04
b0 8
09
#9810000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
0<
#9820000000
0!
0(
b1 /
04
b1 8
09
#9830000000
1!
1(
b1 1
14
17
19
0<
#9840000000
0!
0(
b10 /
04
b10 8
09
#9850000000
1!
1(
b10 1
14
19
0<
#9860000000
0!
0(
b11 /
04
b11 8
09
#9870000000
1!
1(
b11 1
14
19
0<
#9880000000
0!
0(
b100 /
04
b100 8
09
#9890000000
1!
1(
b100 1
14
07
19
0<
#9900000000
0!
0(
b0 /
04
b0 8
09
#9910000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
0<
#9920000000
0!
0(
b1 /
04
b1 8
09
#9930000000
1!
1(
b1 1
14
17
19
0<
#9940000000
0!
0(
b10 /
04
b10 8
09
#9950000000
1!
1(
b10 1
14
19
0<
#9960000000
0!
0(
b11 /
04
b11 8
09
#9970000000
1!
1(
b11 1
14
19
0<
#9980000000
0!
0(
b100 /
04
b100 8
09
#9990000000
1!
1(
b100 1
14
07
19
0<
#10000000000
0!
0(
b0 /
04
b0 8
09
