$date
  Wed May 22 22:33:24 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module math_real $end
$upscope $end
$scope module tb_transmisor_uart $end
$var reg 1 ! clk $end
$var reg 1 " key $end
$var reg 1 # reset $end
$scope module uut $end
$var reg 1 $ clk $end
$var reg 1 % key $end
$var reg 1 & reset $end
$comment state is not handled $end
$var reg 8 ' cadena[7:0] $end
$var reg 1 ( clk_tx $end
$var reg 1 ) clk_11tx $end
$var reg 1 * tx $end
$var reg 1 + done $end
$var reg 1 , send $end
$scope module a $end
$var reg 1 - clk $end
$var reg 1 . reset $end
$var reg 1 / enable $end
$var reg 1 0 cout $end
$var integer 32 1 q $end
$upscope $end
$scope module b $end
$var reg 1 2 clk $end
$var reg 1 3 reset $end
$var reg 1 4 enable $end
$var reg 1 5 cout $end
$var integer 32 6 q $end
$upscope $end
$scope module c $end
$var reg 1 7 clk $end
$var reg 1 8 reset $end
$var reg 1 9 enable $end
$var reg 1 : send $end
$var reg 8 ; cadena[7:0] $end
$var reg 1 < tx $end
$var reg 1 = done $end
$var reg 1 > clkss $end
$var reg 1 ? clkis $end
$var reg 1 @ rst1s $end
$var reg 8 A ds[7:0] $end
$comment estado is not handled $end
$var integer 32 B cnt $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
U"
0#
0$
U%
0&
bUUUUUUUU '
U(
U)
1*
0+
1,
0-
0.
1/
U0
b0 1
02
03
14
U5
b0 6
U7
08
19
1:
bUUUUUUUU ;
1<
0=
0>
0?
0@
bUUUUUUUU A
b1 B
#10000000
1!
1$
0(
0)
1-
00
b1 1
12
05
b1 6
07
#20000000
0!
0$
0-
02
#30000000
1!
1$
1-
b10 1
12
b10 6
#40000000
0!
0$
0-
02
#50000000
1!
1$
1-
b11 1
12
b11 6
#60000000
0!
1"
0$
1%
0-
02
#70000000
1!
1$
1-
b100 1
12
b100 6
#80000000
0!
0$
0-
02
#90000000
1!
1$
1-
b101 1
12
b101 6
#100000000
0!
0$
0-
02
#110000000
1!
1$
1-
b110 1
12
b110 6
#120000000
0!
0$
0-
02
#130000000
1!
1$
1-
b111 1
12
b111 6
#140000000
0!
0$
0-
02
#150000000
1!
1$
1-
b1000 1
12
b1000 6
#160000000
0!
0$
0-
02
#170000000
1!
1$
1-
b1001 1
12
b1001 6
#180000000
0!
0$
0-
02
#190000000
1!
1$
1-
b1010 1
12
b1010 6
#200000000
0!
0$
0-
02
#210000000
1!
1$
1-
b1011 1
12
b1011 6
#220000000
0!
0$
0-
02
#230000000
1!
1$
1-
b1100 1
12
b1100 6
#240000000
0!
0$
0-
02
#250000000
1!
1$
1-
b1101 1
12
b1101 6
#260000000
0!
0$
0-
02
#270000000
1!
1$
1-
b1110 1
12
b1110 6
#280000000
0!
0$
0-
02
#290000000
1!
1$
1-
b1111 1
12
b1111 6
#300000000
0!
0$
0-
02
#310000000
1!
1$
1-
b10000 1
12
b10000 6
#320000000
0!
0$
0-
02
#330000000
1!
1$
1-
b10001 1
12
b10001 6
#340000000
0!
0$
0-
02
#350000000
1!
1$
1-
b10010 1
12
b10010 6
#360000000
0!
0$
0-
02
#370000000
1!
1$
1-
b10011 1
12
b10011 6
#380000000
0!
0"
0$
0%
0-
02
#390000000
1!
1$
1-
b10100 1
12
b10100 6
#400000000
0!
0$
0-
02
#410000000
1!
1$
1-
b10101 1
12
b10101 6
#420000000
0!
0$
0-
02
#430000000
1!
1$
1-
b10110 1
12
b10110 6
#440000000
0!
0$
0-
02
#450000000
1!
1$
1-
b10111 1
12
b10111 6
#460000000
0!
0$
0-
02
#470000000
1!
1$
1-
b11000 1
12
b11000 6
#480000000
0!
0$
0-
02
#490000000
1!
1$
1-
b11001 1
12
b11001 6
#500000000
0!
0$
0-
02
#510000000
1!
1$
1-
b11010 1
12
b11010 6
#520000000
0!
0$
0-
02
#530000000
1!
1$
1-
b11011 1
12
b11011 6
#540000000
0!
0$
0-
02
#550000000
1!
1$
1-
b11100 1
12
b11100 6
#560000000
0!
0$
0-
02
#570000000
1!
1$
1-
b11101 1
12
b11101 6
#580000000
0!
0$
0-
02
#590000000
1!
1$
1-
b11110 1
12
b11110 6
#600000000
0!
0$
0-
02
#610000000
1!
1$
1-
b11111 1
12
b11111 6
#620000000
0!
0$
0-
02
#630000000
1!
1$
1-
b100000 1
12
b100000 6
#640000000
0!
0$
0-
02
#650000000
1!
1$
1-
b100001 1
12
b100001 6
#660000000
0!
0$
0-
02
#670000000
1!
1$
1-
b100010 1
12
b100010 6
#680000000
0!
0$
0-
02
#690000000
1!
1$
1-
b100011 1
12
b100011 6
#700000000
0!
0$
0-
02
#710000000
1!
1$
1-
b100100 1
12
b100100 6
#720000000
0!
0$
0-
02
#730000000
1!
1$
1-
b100101 1
12
b100101 6
#740000000
0!
0$
0-
02
#750000000
1!
1$
1-
b100110 1
12
b100110 6
#760000000
0!
0$
0-
02
#770000000
1!
1$
1-
b100111 1
12
b100111 6
#780000000
0!
0$
0-
02
#790000000
1!
1$
1-
b101000 1
12
b101000 6
#800000000
0!
0$
0-
02
#810000000
1!
1$
1-
b101001 1
12
b101001 6
#820000000
0!
0$
0-
02
#830000000
1!
1$
1-
b101010 1
12
b101010 6
#840000000
0!
0$
0-
02
#850000000
1!
1$
1-
b101011 1
12
b101011 6
#860000000
0!
0$
0-
02
#870000000
1!
1$
1-
b101100 1
12
b101100 6
#880000000
0!
0$
0-
02
#890000000
1!
1$
1-
b101101 1
12
b101101 6
#900000000
0!
0$
0-
02
#910000000
1!
1$
1-
b101110 1
12
b101110 6
#920000000
0!
0$
0-
02
#930000000
1!
1$
1-
b101111 1
12
b101111 6
#940000000
0!
0$
0-
02
#950000000
1!
1$
1-
b110000 1
12
b110000 6
#960000000
0!
0$
0-
02
#970000000
1!
1$
1-
b110001 1
12
b110001 6
#980000000
0!
0$
0-
02
#990000000
1!
1$
1-
b110010 1
12
b110010 6
#1000000000
0!
0$
0-
02
#1010000000
1!
1$
1-
b110011 1
12
b110011 6
#1020000000
0!
0$
0-
02
#1030000000
1!
1$
1-
b110100 1
12
b110100 6
#1040000000
0!
0$
0-
02
#1050000000
1!
1$
1-
b110101 1
12
b110101 6
#1060000000
0!
0$
0-
02
#1070000000
1!
1$
1-
b110110 1
12
b110110 6
#1080000000
0!
0$
0-
02
#1090000000
1!
1$
1-
b110111 1
12
b110111 6
#1100000000
0!
0$
0-
02
#1110000000
1!
1$
1-
b111000 1
12
b111000 6
#1120000000
0!
0$
0-
02
#1130000000
1!
1$
1-
b111001 1
12
b111001 6
#1140000000
0!
0$
0-
02
#1150000000
1!
1$
1-
b111010 1
12
b111010 6
#1160000000
0!
0$
0-
02
#1170000000
1!
1$
1-
b111011 1
12
b111011 6
#1180000000
0!
0$
0-
02
#1190000000
1!
1$
1-
b111100 1
12
b111100 6
#1200000000
0!
0$
0-
02
#1210000000
1!
1$
1-
b111101 1
12
b111101 6
#1220000000
0!
0$
0-
02
#1230000000
1!
1$
1-
b111110 1
12
b111110 6
#1240000000
0!
0$
0-
02
#1250000000
1!
1$
1-
b111111 1
12
b111111 6
#1260000000
0!
0$
0-
02
#1270000000
1!
1$
1-
b1000000 1
12
b1000000 6
#1280000000
0!
0$
0-
02
#1290000000
1!
1$
1-
b1000001 1
12
b1000001 6
#1300000000
0!
0$
0-
02
#1310000000
1!
1$
1-
b1000010 1
12
b1000010 6
#1320000000
0!
0$
0-
02
#1330000000
1!
1$
1-
b1000011 1
12
b1000011 6
#1340000000
0!
0$
0-
02
#1350000000
1!
1$
1-
b1000100 1
12
b1000100 6
#1360000000
0!
0$
0-
02
#1370000000
1!
1$
1-
b1000101 1
12
b1000101 6
#1380000000
0!
0$
0-
02
#1390000000
1!
1$
1-
b1000110 1
12
b1000110 6
#1400000000
0!
0$
0-
02
#1410000000
1!
1$
1-
b1000111 1
12
b1000111 6
#1420000000
0!
1"
0$
1%
0-
02
#1430000000
1!
1$
1-
b1001000 1
12
b1001000 6
#1440000000
0!
0$
0-
02
#1450000000
1!
1$
1-
b1001001 1
12
b1001001 6
#1460000000
0!
0$
0-
02
#1470000000
1!
1$
1-
b1001010 1
12
b1001010 6
#1480000000
0!
0$
0-
02
#1490000000
1!
1$
1-
b1001011 1
12
b1001011 6
#1500000000
0!
0$
0-
02
#1510000000
1!
1$
1-
b1001100 1
12
b1001100 6
#1520000000
0!
0$
0-
02
#1530000000
1!
1$
1-
b1001101 1
12
b1001101 6
#1540000000
0!
0$
0-
02
#1550000000
1!
1$
1-
b1001110 1
12
b1001110 6
#1560000000
0!
0$
0-
02
#1570000000
1!
1$
1-
b1001111 1
12
b1001111 6
#1580000000
0!
0$
0-
02
#1590000000
1!
1$
1-
b1010000 1
12
b1010000 6
#1600000000
0!
0$
0-
02
#1610000000
1!
1$
1-
b1010001 1
12
b1010001 6
#1620000000
0!
0$
0-
02
#1630000000
1!
1$
1-
b1010010 1
12
b1010010 6
#1640000000
0!
0$
0-
02
#1650000000
1!
1$
1-
b1010011 1
12
b1010011 6
#1660000000
0!
0$
0-
02
#1670000000
1!
1$
1-
b1010100 1
12
b1010100 6
#1680000000
0!
0$
0-
02
#1690000000
1!
1$
1-
b1010101 1
12
b1010101 6
#1700000000
0!
0$
0-
02
#1710000000
1!
1$
1-
b1010110 1
12
b1010110 6
#1720000000
0!
0$
0-
02
#1730000000
1!
1$
1-
b1010111 1
12
b1010111 6
#1740000000
0!
0"
0$
0%
0-
02
#1750000000
1!
1$
1-
b1011000 1
12
b1011000 6
#1760000000
0!
0$
0-
02
#1770000000
1!
1$
1-
b1011001 1
12
b1011001 6
#1780000000
0!
0$
0-
02
#1790000000
1!
1$
1-
b1011010 1
12
b1011010 6
#1800000000
0!
0$
0-
02
#1810000000
1!
1$
1-
b1011011 1
12
b1011011 6
#1820000000
0!
0$
0-
02
#1830000000
1!
1$
1-
b1011100 1
12
b1011100 6
#1840000000
0!
0$
0-
02
#1850000000
1!
1$
1-
b1011101 1
12
b1011101 6
#1860000000
0!
0$
0-
02
#1870000000
1!
1$
1-
b1011110 1
12
b1011110 6
#1880000000
0!
0$
0-
02
#1890000000
1!
1$
1-
b1011111 1
12
b1011111 6
#1900000000
0!
0$
0-
02
#1910000000
1!
1$
1-
b1100000 1
12
b1100000 6
#1920000000
0!
0$
0-
02
#1930000000
1!
1$
1-
b1100001 1
12
b1100001 6
#1940000000
0!
0$
0-
02
#1950000000
1!
1$
1-
b1100010 1
12
b1100010 6
#1960000000
0!
0$
0-
02
#1970000000
1!
1$
1-
b1100011 1
12
b1100011 6
#1980000000
0!
0$
0-
02
#1990000000
1!
1$
1-
b1100100 1
12
b1100100 6
#2000000000
0!
0$
0-
02
#2010000000
1!
1$
1-
b1100101 1
12
b1100101 6
#2020000000
0!
0$
0-
02
#2030000000
1!
1$
1-
b1100110 1
12
b1100110 6
#2040000000
0!
0$
0-
02
#2050000000
1!
1$
1-
b1100111 1
12
b1100111 6
#2060000000
0!
0$
0-
02
#2070000000
1!
1$
1-
b1101000 1
12
b1101000 6
#2080000000
0!
0$
0-
02
#2090000000
1!
1$
1-
b1101001 1
12
b1101001 6
#2100000000
0!
0$
0-
02
#2110000000
1!
1$
1-
b1101010 1
12
b1101010 6
#2120000000
0!
0$
0-
02
#2130000000
1!
1$
1-
b1101011 1
12
b1101011 6
#2140000000
0!
0$
0-
02
#2150000000
1!
1$
1-
b1101100 1
12
b1101100 6
#2160000000
0!
0$
0-
02
#2170000000
1!
1$
1-
b1101101 1
12
b1101101 6
#2180000000
0!
0$
0-
02
#2190000000
1!
1$
1-
b1101110 1
12
b1101110 6
#2200000000
0!
0$
0-
02
#2210000000
1!
1$
1-
b1101111 1
12
b1101111 6
#2220000000
0!
0$
0-
02
#2230000000
1!
1$
1-
b1110000 1
12
b1110000 6
#2240000000
0!
0$
0-
02
#2250000000
1!
1$
1-
b1110001 1
12
b1110001 6
#2260000000
0!
0$
0-
02
#2270000000
1!
1$
1-
b1110010 1
12
b1110010 6
#2280000000
0!
0$
0-
02
#2290000000
1!
1$
1-
b1110011 1
12
b1110011 6
#2300000000
0!
0$
0-
02
#2310000000
1!
1$
1-
b1110100 1
12
b1110100 6
#2320000000
0!
0$
0-
02
#2330000000
1!
1$
1-
b1110101 1
12
b1110101 6
#2340000000
0!
0$
0-
02
#2350000000
1!
1$
1-
b1110110 1
12
b1110110 6
#2360000000
0!
0$
0-
02
#2370000000
1!
1$
1-
b1110111 1
12
b1110111 6
#2380000000
0!
0$
0-
02
#2390000000
1!
1$
1-
b1111000 1
12
b1111000 6
#2400000000
0!
0$
0-
02
#2410000000
1!
1$
1-
b1111001 1
12
b1111001 6
#2420000000
0!
0$
0-
02
#2430000000
1!
1$
1-
b1111010 1
12
b1111010 6
#2440000000
0!
0$
0-
02
#2450000000
1!
1$
1-
b1111011 1
12
b1111011 6
#2460000000
0!
0$
0-
02
#2470000000
1!
1$
1-
b1111100 1
12
b1111100 6
#2480000000
0!
0$
0-
02
#2490000000
1!
1$
1-
b1111101 1
12
b1111101 6
#2500000000
0!
0$
0-
02
#2510000000
1!
1$
1-
b1111110 1
12
b1111110 6
#2520000000
0!
0$
0-
02
#2530000000
1!
1$
1-
b1111111 1
12
b1111111 6
#2540000000
0!
0$
0-
02
#2550000000
1!
1$
1-
b10000000 1
12
b10000000 6
#2560000000
0!
0$
0-
02
#2570000000
1!
1$
1-
b10000001 1
12
b10000001 6
#2580000000
0!
0$
0-
02
#2590000000
1!
1$
1-
b10000010 1
12
b10000010 6
#2600000000
0!
0$
0-
02
#2610000000
1!
1$
1-
b10000011 1
12
b10000011 6
#2620000000
0!
0$
0-
02
#2630000000
1!
1$
1-
b10000100 1
12
b10000100 6
#2640000000
0!
0$
0-
02
#2650000000
1!
1$
1-
b10000101 1
12
b10000101 6
#2660000000
0!
0$
0-
02
#2670000000
1!
1$
1-
b10000110 1
12
b10000110 6
#2680000000
0!
0$
0-
02
#2690000000
1!
1$
1-
b10000111 1
12
b10000111 6
#2700000000
0!
0$
0-
02
#2710000000
1!
1$
1-
b10001000 1
12
b10001000 6
#2720000000
0!
0$
0-
02
#2730000000
1!
1$
1-
b10001001 1
12
b10001001 6
#2740000000
0!
0$
0-
02
#2750000000
1!
1$
1-
b10001010 1
12
b10001010 6
#2760000000
0!
0$
0-
02
#2770000000
1!
1$
1-
b10001011 1
12
b10001011 6
#2780000000
0!
1"
0$
1%
0-
02
#2790000000
1!
1$
1-
b10001100 1
12
b10001100 6
#2800000000
0!
0$
0-
02
#2810000000
1!
1$
1-
b10001101 1
12
b10001101 6
#2820000000
0!
0$
0-
02
#2830000000
1!
1$
1-
b10001110 1
12
b10001110 6
#2840000000
0!
0$
0-
02
#2850000000
1!
1$
1-
b10001111 1
12
b10001111 6
#2860000000
0!
0$
0-
02
#2870000000
1!
1$
1-
b10010000 1
12
b10010000 6
#2880000000
0!
0$
0-
02
#2890000000
1!
1$
1-
b10010001 1
12
b10010001 6
#2900000000
0!
0$
0-
02
#2910000000
1!
1$
1-
b10010010 1
12
b10010010 6
#2920000000
0!
0$
0-
02
#2930000000
1!
1$
1-
b10010011 1
12
b10010011 6
#2940000000
0!
0$
0-
02
#2950000000
1!
1$
1-
b10010100 1
12
b10010100 6
#2960000000
0!
0$
0-
02
#2970000000
1!
1$
1-
b10010101 1
12
b10010101 6
#2980000000
0!
0$
0-
02
#2990000000
1!
1$
1-
b10010110 1
12
b10010110 6
#3000000000
0!
0$
0-
02
#3010000000
1!
1$
1-
b10010111 1
12
b10010111 6
#3020000000
0!
0$
0-
02
#3030000000
1!
1$
1-
b10011000 1
12
b10011000 6
#3040000000
0!
0$
0-
02
#3050000000
1!
1$
1-
b10011001 1
12
b10011001 6
#3060000000
0!
0$
0-
02
#3070000000
1!
1$
1-
b10011010 1
12
b10011010 6
#3080000000
0!
0$
0-
02
#3090000000
1!
1$
1-
b10011011 1
12
b10011011 6
#3100000000
0!
0"
0$
0%
0-
02
#3110000000
1!
1$
1-
b10011100 1
12
b10011100 6
#3120000000
0!
0$
0-
02
#3130000000
1!
1$
1-
b10011101 1
12
b10011101 6
#3140000000
0!
0$
0-
02
#3150000000
1!
1$
1-
b10011110 1
12
b10011110 6
#3160000000
0!
0$
0-
02
#3170000000
1!
1$
1-
b10011111 1
12
b10011111 6
#3180000000
0!
0$
0-
02
#3190000000
1!
1$
1-
b10100000 1
12
b10100000 6
#3200000000
0!
0$
0-
02
#3210000000
1!
1$
1-
b10100001 1
12
b10100001 6
#3220000000
0!
0$
0-
02
#3230000000
1!
1$
1-
b10100010 1
12
b10100010 6
#3240000000
0!
0$
0-
02
#3250000000
1!
1$
1-
b10100011 1
12
b10100011 6
#3260000000
0!
0$
0-
02
#3270000000
1!
1$
1-
b10100100 1
12
b10100100 6
#3280000000
0!
0$
0-
02
#3290000000
1!
1$
1-
b10100101 1
12
b10100101 6
#3300000000
0!
0$
0-
02
#3310000000
1!
1$
1-
b10100110 1
12
b10100110 6
#3320000000
0!
0$
0-
02
#3330000000
1!
1$
1-
b10100111 1
12
b10100111 6
#3340000000
0!
0$
0-
02
#3350000000
1!
1$
1-
b10101000 1
12
b10101000 6
#3360000000
0!
0$
0-
02
#3370000000
1!
1$
1-
b10101001 1
12
b10101001 6
#3380000000
0!
0$
0-
02
#3390000000
1!
1$
1-
b10101010 1
12
b10101010 6
#3400000000
0!
0$
0-
02
#3410000000
1!
1$
1-
b10101011 1
12
b10101011 6
#3420000000
0!
0$
0-
02
#3430000000
1!
1$
1-
b10101100 1
12
b10101100 6
#3440000000
0!
0$
0-
02
#3450000000
1!
1$
1-
b10101101 1
12
b10101101 6
#3460000000
0!
0$
0-
02
#3470000000
1!
1$
1-
b10101110 1
12
b10101110 6
#3480000000
0!
0$
0-
02
#3490000000
1!
1$
1-
b10101111 1
12
b10101111 6
#3500000000
0!
0$
0-
02
#3510000000
1!
1$
1-
b10110000 1
12
b10110000 6
#3520000000
0!
0$
0-
02
#3530000000
1!
1$
1-
b10110001 1
12
b10110001 6
#3540000000
0!
0$
0-
02
#3550000000
1!
1$
1-
b10110010 1
12
b10110010 6
#3560000000
0!
0$
0-
02
#3570000000
1!
1$
1-
b10110011 1
12
b10110011 6
#3580000000
0!
0$
0-
02
#3590000000
1!
1$
1-
b10110100 1
12
b10110100 6
#3600000000
0!
0$
0-
02
#3610000000
1!
1$
1-
b10110101 1
12
b10110101 6
#3620000000
0!
0$
0-
02
#3630000000
1!
1$
1-
b10110110 1
12
b10110110 6
#3640000000
0!
0$
0-
02
#3650000000
1!
1$
1-
b10110111 1
12
b10110111 6
#3660000000
0!
0$
0-
02
#3670000000
1!
1$
1-
b10111000 1
12
b10111000 6
#3680000000
0!
0$
0-
02
#3690000000
1!
1$
1-
b10111001 1
12
b10111001 6
#3700000000
0!
0$
0-
02
#3710000000
1!
1$
1-
b10111010 1
12
b10111010 6
#3720000000
0!
0$
0-
02
#3730000000
1!
1$
1-
b10111011 1
12
b10111011 6
#3740000000
0!
0$
0-
02
#3750000000
1!
1$
1-
b10111100 1
12
b10111100 6
#3760000000
0!
0$
0-
02
#3770000000
1!
1$
1-
b10111101 1
12
b10111101 6
#3780000000
0!
0$
0-
02
#3790000000
1!
1$
1-
b10111110 1
12
b10111110 6
#3800000000
0!
0$
0-
02
#3810000000
1!
1$
1-
b10111111 1
12
b10111111 6
#3820000000
0!
0$
0-
02
#3830000000
1!
1$
1-
b11000000 1
12
b11000000 6
#3840000000
0!
0$
0-
02
#3850000000
1!
1$
1-
b11000001 1
12
b11000001 6
#3860000000
0!
0$
0-
02
#3870000000
1!
1$
1-
b11000010 1
12
b11000010 6
#3880000000
0!
0$
0-
02
#3890000000
1!
1$
1-
b11000011 1
12
b11000011 6
#3900000000
0!
0$
0-
02
#3910000000
1!
1$
1-
b11000100 1
12
b11000100 6
#3920000000
0!
0$
0-
02
#3930000000
1!
1$
1-
b11000101 1
12
b11000101 6
#3940000000
0!
0$
0-
02
#3950000000
1!
1$
1-
b11000110 1
12
b11000110 6
#3960000000
0!
0$
0-
02
#3970000000
1!
1$
1-
b11000111 1
12
b11000111 6
#3980000000
0!
0$
0-
02
#3990000000
1!
1$
1-
b11001000 1
12
b11001000 6
#4000000000
0!
0$
0-
02
#4010000000
1!
1$
1-
b11001001 1
12
b11001001 6
#4020000000
0!
0$
0-
02
#4030000000
1!
1$
1-
b11001010 1
12
b11001010 6
#4040000000
0!
0$
0-
02
#4050000000
1!
1$
1-
b11001011 1
12
b11001011 6
#4060000000
0!
0$
0-
02
#4070000000
1!
1$
1-
b11001100 1
12
b11001100 6
#4080000000
0!
0$
0-
02
#4090000000
1!
1$
1-
b11001101 1
12
b11001101 6
#4100000000
0!
0$
0-
02
#4110000000
1!
1$
1-
b11001110 1
12
b11001110 6
#4120000000
0!
0$
0-
02
#4130000000
1!
1$
1-
b11001111 1
12
b11001111 6
#4140000000
0!
1"
0$
1%
0-
02
#4150000000
1!
1$
1-
b11010000 1
12
b11010000 6
#4160000000
0!
0$
0-
02
#4170000000
1!
1$
1-
b11010001 1
12
b11010001 6
#4180000000
0!
0$
0-
02
#4190000000
1!
1$
1-
b11010010 1
12
b11010010 6
#4200000000
0!
0$
0-
02
#4210000000
1!
1$
1-
b11010011 1
12
b11010011 6
#4220000000
0!
0$
0-
02
#4230000000
1!
1$
1-
b11010100 1
12
b11010100 6
#4240000000
0!
0$
0-
02
#4250000000
1!
1$
1-
b11010101 1
12
b11010101 6
#4260000000
0!
0$
0-
02
#4270000000
1!
1$
1-
b11010110 1
12
b11010110 6
#4280000000
0!
0$
0-
02
#4290000000
1!
1$
1-
b11010111 1
12
b11010111 6
#4300000000
0!
0$
0-
02
#4310000000
1!
1$
1-
b11011000 1
12
b11011000 6
#4320000000
0!
0$
0-
02
#4330000000
1!
1$
1-
b11011001 1
12
b11011001 6
#4340000000
0!
0$
0-
02
#4350000000
1!
1$
1-
b11011010 1
12
b11011010 6
#4360000000
0!
0$
0-
02
#4370000000
1!
1$
1-
b11011011 1
12
b11011011 6
#4380000000
0!
0$
0-
02
#4390000000
1!
1$
1-
b11011100 1
12
b11011100 6
#4400000000
0!
0$
0-
02
#4410000000
1!
1$
1-
b11011101 1
12
b11011101 6
#4420000000
0!
0$
0-
02
#4430000000
1!
1$
1-
b11011110 1
12
b11011110 6
#4440000000
0!
0$
0-
02
#4450000000
1!
1$
1-
b11011111 1
12
b11011111 6
#4460000000
0!
0"
0$
0%
0-
02
#4470000000
1!
1$
1-
b11100000 1
12
b11100000 6
#4480000000
0!
0$
0-
02
#4490000000
1!
1$
1-
b11100001 1
12
b11100001 6
#4500000000
0!
0$
0-
02
#4510000000
1!
1$
1-
b11100010 1
12
b11100010 6
#4520000000
0!
0$
0-
02
#4530000000
1!
1$
1-
b11100011 1
12
b11100011 6
#4540000000
0!
0$
0-
02
#4550000000
1!
1$
1-
b11100100 1
12
b11100100 6
#4560000000
0!
0$
0-
02
#4570000000
1!
1$
1-
b11100101 1
12
b11100101 6
#4580000000
0!
0$
0-
02
#4590000000
1!
1$
1-
b11100110 1
12
b11100110 6
#4600000000
0!
0$
0-
02
#4610000000
1!
1$
1-
b11100111 1
12
b11100111 6
#4620000000
0!
0$
0-
02
#4630000000
1!
1$
1-
b11101000 1
12
b11101000 6
#4640000000
0!
0$
0-
02
#4650000000
1!
1$
1-
b11101001 1
12
b11101001 6
#4660000000
0!
0$
0-
02
#4670000000
1!
1$
1-
b11101010 1
12
b11101010 6
#4680000000
0!
0$
0-
02
#4690000000
1!
1$
1-
b11101011 1
12
b11101011 6
#4700000000
0!
0$
0-
02
#4710000000
1!
1$
1-
b11101100 1
12
b11101100 6
#4720000000
0!
0$
0-
02
#4730000000
1!
1$
1-
b11101101 1
12
b11101101 6
#4740000000
0!
0$
0-
02
#4750000000
1!
1$
1-
b11101110 1
12
b11101110 6
#4760000000
0!
0$
0-
02
#4770000000
1!
1$
1-
b11101111 1
12
b11101111 6
#4780000000
0!
0$
0-
02
#4790000000
1!
1$
1-
b11110000 1
12
b11110000 6
#4800000000
0!
0$
0-
02
#4810000000
1!
1$
1-
b11110001 1
12
b11110001 6
#4820000000
0!
0$
0-
02
#4830000000
1!
1$
1-
b11110010 1
12
b11110010 6
#4840000000
0!
0$
0-
02
#4850000000
1!
1$
1-
b11110011 1
12
b11110011 6
#4860000000
0!
0$
0-
02
#4870000000
1!
1$
1-
b11110100 1
12
b11110100 6
#4880000000
0!
0$
0-
02
#4890000000
1!
1$
1-
b11110101 1
12
b11110101 6
#4900000000
0!
0$
0-
02
#4910000000
1!
1$
1-
b11110110 1
12
b11110110 6
#4920000000
0!
0$
0-
02
#4930000000
1!
1$
1-
b11110111 1
12
b11110111 6
#4940000000
0!
0$
0-
02
#4950000000
1!
1$
1-
b11111000 1
12
b11111000 6
#4960000000
0!
0$
0-
02
#4970000000
1!
1$
1-
b11111001 1
12
b11111001 6
#4980000000
0!
0$
0-
02
#4990000000
1!
1$
1-
b11111010 1
12
b11111010 6
#5000000000
0!
0$
0-
02
#5010000000
1!
1$
1-
b11111011 1
12
b11111011 6
#5020000000
0!
0$
0-
02
#5030000000
1!
1$
1-
b11111100 1
12
b11111100 6
#5040000000
0!
0$
0-
02
#5050000000
1!
1$
1-
b11111101 1
12
b11111101 6
#5060000000
0!
0$
0-
02
#5070000000
1!
1$
1-
b11111110 1
12
b11111110 6
#5080000000
0!
0$
0-
02
#5090000000
1!
1$
1-
b11111111 1
12
b11111111 6
#5100000000
0!
0$
0-
02
#5110000000
1!
1$
1-
b100000000 1
12
b100000000 6
#5120000000
0!
0$
0-
02
#5130000000
1!
1$
1-
b100000001 1
12
b100000001 6
#5140000000
0!
0$
0-
02
#5150000000
1!
1$
1-
b100000010 1
12
b100000010 6
#5160000000
0!
0$
0-
02
#5170000000
1!
1$
1-
b100000011 1
12
b100000011 6
#5180000000
0!
0$
0-
02
#5190000000
1!
1$
1-
b100000100 1
12
b100000100 6
#5200000000
0!
0$
0-
02
#5210000000
1!
1$
1-
b100000101 1
12
b100000101 6
#5220000000
0!
0$
0-
02
#5230000000
1!
1$
1-
b100000110 1
12
b100000110 6
#5240000000
0!
0$
0-
02
#5250000000
1!
1$
1-
b100000111 1
12
b100000111 6
#5260000000
0!
0$
0-
02
#5270000000
1!
1$
1-
b100001000 1
12
b100001000 6
#5280000000
0!
0$
0-
02
#5290000000
1!
1$
1-
b100001001 1
12
b100001001 6
#5300000000
0!
0$
0-
02
#5310000000
1!
1$
1-
b100001010 1
12
b100001010 6
#5320000000
0!
0$
0-
02
#5330000000
1!
1$
1-
b100001011 1
12
b100001011 6
#5340000000
0!
0$
0-
02
#5350000000
1!
1$
1-
b100001100 1
12
b100001100 6
#5360000000
0!
0$
0-
02
#5370000000
1!
1$
1-
b100001101 1
12
b100001101 6
#5380000000
0!
0$
0-
02
#5390000000
1!
1$
1-
b100001110 1
12
b100001110 6
#5400000000
0!
0$
0-
02
#5410000000
1!
1$
1-
b100001111 1
12
b100001111 6
#5420000000
0!
0$
0-
02
#5430000000
1!
1$
1-
b100010000 1
12
b100010000 6
#5440000000
0!
0$
0-
02
#5450000000
1!
1$
1-
b100010001 1
12
b100010001 6
#5460000000
0!
0$
0-
02
#5470000000
1!
1$
1-
b100010010 1
12
b100010010 6
#5480000000
0!
0$
0-
02
#5490000000
1!
1$
1-
b100010011 1
12
b100010011 6
#5500000000
0!
1"
0$
1%
0-
02
#5510000000
1!
1$
1-
b100010100 1
12
b100010100 6
#5520000000
0!
0$
0-
02
#5530000000
1!
1$
1-
b100010101 1
12
b100010101 6
#5540000000
0!
0$
0-
02
#5550000000
1!
1$
1-
b100010110 1
12
b100010110 6
#5560000000
0!
0$
0-
02
#5570000000
1!
1$
1-
b100010111 1
12
b100010111 6
#5580000000
0!
0$
0-
02
#5590000000
1!
1$
1-
b100011000 1
12
b100011000 6
#5600000000
0!
0$
0-
02
#5610000000
1!
1$
1-
b100011001 1
12
b100011001 6
#5620000000
0!
0$
0-
02
#5630000000
1!
1$
1-
b100011010 1
12
b100011010 6
#5640000000
0!
0$
0-
02
#5650000000
1!
1$
1-
b100011011 1
12
b100011011 6
#5660000000
0!
0$
0-
02
#5670000000
1!
1$
1-
b100011100 1
12
b100011100 6
#5680000000
0!
0$
0-
02
#5690000000
1!
1$
1-
b100011101 1
12
b100011101 6
#5700000000
0!
0$
0-
02
#5710000000
1!
1$
1-
b100011110 1
12
b100011110 6
#5720000000
0!
0$
0-
02
#5730000000
1!
1$
1-
b100011111 1
12
b100011111 6
#5740000000
0!
0$
0-
02
#5750000000
1!
1$
1-
b100100000 1
12
b100100000 6
#5760000000
0!
0$
0-
02
#5770000000
1!
1$
1-
b100100001 1
12
b100100001 6
#5780000000
0!
0$
0-
02
#5790000000
1!
1$
1-
b100100010 1
12
b100100010 6
#5800000000
0!
0$
0-
02
#5810000000
1!
1$
1-
b100100011 1
12
b100100011 6
#5820000000
0!
0"
0$
0%
0-
02
#5830000000
1!
1$
1-
b100100100 1
12
b100100100 6
#5840000000
0!
0$
0-
02
#5850000000
1!
1$
1-
b100100101 1
12
b100100101 6
#5860000000
0!
0$
0-
02
#5870000000
1!
1$
1-
b100100110 1
12
b100100110 6
#5880000000
0!
0$
0-
02
#5890000000
1!
1$
1-
b100100111 1
12
b100100111 6
#5900000000
0!
0$
0-
02
#5910000000
1!
1$
1-
b100101000 1
12
b100101000 6
#5920000000
0!
0$
0-
02
#5930000000
1!
1$
1-
b100101001 1
12
b100101001 6
#5940000000
0!
0$
0-
02
#5950000000
1!
1$
1-
b100101010 1
12
b100101010 6
#5960000000
0!
0$
0-
02
#5970000000
1!
1$
1-
b100101011 1
12
b100101011 6
#5980000000
0!
0$
0-
02
#5990000000
1!
1$
1-
b100101100 1
12
b100101100 6
#6000000000
0!
0$
0-
02
#6010000000
1!
1$
1-
b100101101 1
12
b100101101 6
#6020000000
0!
0$
0-
02
#6030000000
1!
1$
1-
b100101110 1
12
b100101110 6
#6040000000
0!
0$
0-
02
#6050000000
1!
1$
1-
b100101111 1
12
b100101111 6
#6060000000
0!
0$
0-
02
#6070000000
1!
1$
1-
b100110000 1
12
b100110000 6
#6080000000
0!
0$
0-
02
#6090000000
1!
1$
1-
b100110001 1
12
b100110001 6
#6100000000
0!
0$
0-
02
#6110000000
1!
1$
1-
b100110010 1
12
b100110010 6
#6120000000
0!
0$
0-
02
#6130000000
1!
1$
1-
b100110011 1
12
b100110011 6
#6140000000
0!
0$
0-
02
#6150000000
1!
1$
1-
b100110100 1
12
b100110100 6
#6160000000
0!
0$
0-
02
#6170000000
1!
1$
1-
b100110101 1
12
b100110101 6
#6180000000
0!
0$
0-
02
#6190000000
1!
1$
1-
b100110110 1
12
b100110110 6
#6200000000
0!
0$
0-
02
#6210000000
1!
1$
1-
b100110111 1
12
b100110111 6
#6220000000
0!
0$
0-
02
#6230000000
1!
1$
1-
b100111000 1
12
b100111000 6
#6240000000
0!
0$
0-
02
#6250000000
1!
1$
1-
b100111001 1
12
b100111001 6
#6260000000
0!
0$
0-
02
#6270000000
1!
1$
1-
b100111010 1
12
b100111010 6
#6280000000
0!
0$
0-
02
#6290000000
1!
1$
1-
b100111011 1
12
b100111011 6
#6300000000
0!
0$
0-
02
#6310000000
1!
1$
1-
b100111100 1
12
b100111100 6
#6320000000
0!
0$
0-
02
#6330000000
1!
1$
1-
b100111101 1
12
b100111101 6
#6340000000
0!
0$
0-
02
#6350000000
1!
1$
1-
b100111110 1
12
b100111110 6
#6360000000
0!
0$
0-
02
#6370000000
1!
1$
1-
b100111111 1
12
b100111111 6
#6380000000
0!
0$
0-
02
#6390000000
1!
1$
1-
b101000000 1
12
b101000000 6
#6400000000
0!
0$
0-
02
#6410000000
1!
1$
1-
b101000001 1
12
b101000001 6
#6420000000
0!
0$
0-
02
#6430000000
1!
1$
1-
b101000010 1
12
b101000010 6
#6440000000
0!
0$
0-
02
#6450000000
1!
1$
1-
b101000011 1
12
b101000011 6
#6460000000
0!
0$
0-
02
#6470000000
1!
1$
1-
b101000100 1
12
b101000100 6
#6480000000
0!
0$
0-
02
#6490000000
1!
1$
1-
b101000101 1
12
b101000101 6
#6500000000
0!
0$
0-
02
#6510000000
1!
1$
1-
b101000110 1
12
b101000110 6
#6520000000
0!
0$
0-
02
#6530000000
1!
1$
1-
b101000111 1
12
b101000111 6
#6540000000
0!
0$
0-
02
#6550000000
1!
1$
1-
b101001000 1
12
b101001000 6
#6560000000
0!
0$
0-
02
#6570000000
1!
1$
1-
b101001001 1
12
b101001001 6
#6580000000
0!
0$
0-
02
#6590000000
1!
1$
1-
b101001010 1
12
b101001010 6
#6600000000
0!
0$
0-
02
#6610000000
1!
1$
1-
b101001011 1
12
b101001011 6
#6620000000
0!
0$
0-
02
#6630000000
1!
1$
1-
b101001100 1
12
b101001100 6
#6640000000
0!
0$
0-
02
#6650000000
1!
1$
1-
b101001101 1
12
b101001101 6
#6660000000
0!
0$
0-
02
#6670000000
1!
1$
1-
b101001110 1
12
b101001110 6
#6680000000
0!
0$
0-
02
#6690000000
1!
1$
1-
b101001111 1
12
b101001111 6
#6700000000
0!
0$
0-
02
#6710000000
1!
1$
1-
b101010000 1
12
b101010000 6
#6720000000
0!
0$
0-
02
#6730000000
1!
1$
1-
b101010001 1
12
b101010001 6
#6740000000
0!
0$
0-
02
#6750000000
1!
1$
1-
b101010010 1
12
b101010010 6
#6760000000
0!
0$
0-
02
#6770000000
1!
1$
1-
b101010011 1
12
b101010011 6
#6780000000
0!
0$
0-
02
#6790000000
1!
1$
1-
b101010100 1
12
b101010100 6
#6800000000
0!
0$
0-
02
#6810000000
1!
1$
1-
b101010101 1
12
b101010101 6
#6820000000
0!
0$
0-
02
#6830000000
1!
1$
1-
b101010110 1
12
b101010110 6
#6840000000
0!
0$
0-
02
#6850000000
1!
1$
1-
b101010111 1
12
b101010111 6
#6860000000
0!
1"
0$
1%
0-
02
#6870000000
1!
1$
1-
b101011000 1
12
b101011000 6
#6880000000
0!
0$
0-
02
#6890000000
1!
1$
1-
b101011001 1
12
b101011001 6
#6900000000
0!
0$
0-
02
#6910000000
1!
1$
1-
b101011010 1
12
b101011010 6
#6920000000
0!
0$
0-
02
#6930000000
1!
1$
1-
b101011011 1
12
b101011011 6
#6940000000
0!
0$
0-
02
#6950000000
1!
1$
1-
b101011100 1
12
b101011100 6
#6960000000
0!
0$
0-
02
#6970000000
1!
1$
1-
b101011101 1
12
b101011101 6
#6980000000
0!
0$
0-
02
#6990000000
1!
1$
1-
b101011110 1
12
b101011110 6
#7000000000
0!
0$
0-
02
#7010000000
1!
1$
1-
b101011111 1
12
b101011111 6
#7020000000
0!
0$
0-
02
#7030000000
1!
1$
1-
b101100000 1
12
b101100000 6
#7040000000
0!
0$
0-
02
#7050000000
1!
1$
1-
b101100001 1
12
b101100001 6
#7060000000
0!
0$
0-
02
#7070000000
1!
1$
1-
b101100010 1
12
b101100010 6
#7080000000
0!
0$
0-
02
#7090000000
1!
1$
1-
b101100011 1
12
b101100011 6
#7100000000
0!
0$
0-
02
#7110000000
1!
1$
1-
b101100100 1
12
b101100100 6
#7120000000
0!
0$
0-
02
#7130000000
1!
1$
1-
b101100101 1
12
b101100101 6
#7140000000
0!
0$
0-
02
#7150000000
1!
1$
1-
b101100110 1
12
b101100110 6
#7160000000
0!
0$
0-
02
#7170000000
1!
1$
1-
b101100111 1
12
b101100111 6
#7180000000
0!
0"
0$
0%
0-
02
#7190000000
1!
1$
1-
b101101000 1
12
b101101000 6
#7200000000
0!
0$
0-
02
#7210000000
1!
1$
1-
b101101001 1
12
b101101001 6
#7220000000
0!
0$
0-
02
#7230000000
1!
1$
1-
b101101010 1
12
b101101010 6
#7240000000
0!
0$
0-
02
#7250000000
1!
1$
1-
b101101011 1
12
b101101011 6
#7260000000
0!
0$
0-
02
#7270000000
1!
1$
1-
b101101100 1
12
b101101100 6
#7280000000
0!
0$
0-
02
#7290000000
1!
1$
1-
b101101101 1
12
b101101101 6
#7300000000
0!
0$
0-
02
#7310000000
1!
1$
1-
b101101110 1
12
b101101110 6
#7320000000
0!
0$
0-
02
#7330000000
1!
1$
1-
b101101111 1
12
b101101111 6
#7340000000
0!
0$
0-
02
#7350000000
1!
1$
1-
b101110000 1
12
b101110000 6
#7360000000
0!
0$
0-
02
#7370000000
1!
1$
1-
b101110001 1
12
b101110001 6
#7380000000
0!
0$
0-
02
#7390000000
1!
1$
1-
b101110010 1
12
b101110010 6
#7400000000
0!
0$
0-
02
#7410000000
1!
1$
1-
b101110011 1
12
b101110011 6
#7420000000
0!
0$
0-
02
#7430000000
1!
1$
1-
b101110100 1
12
b101110100 6
#7440000000
0!
0$
0-
02
#7450000000
1!
1$
1-
b101110101 1
12
b101110101 6
#7460000000
0!
0$
0-
02
#7470000000
1!
1$
1-
b101110110 1
12
b101110110 6
#7480000000
0!
0$
0-
02
#7490000000
1!
1$
1-
b101110111 1
12
b101110111 6
#7500000000
0!
0$
0-
02
#7510000000
1!
1$
1-
b101111000 1
12
b101111000 6
#7520000000
0!
0$
0-
02
#7530000000
1!
1$
1-
b101111001 1
12
b101111001 6
#7540000000
0!
0$
0-
02
#7550000000
1!
1$
1-
b101111010 1
12
b101111010 6
#7560000000
0!
0$
0-
02
#7570000000
1!
1$
1-
b101111011 1
12
b101111011 6
#7580000000
0!
0$
0-
02
#7590000000
1!
1$
1-
b101111100 1
12
b101111100 6
#7600000000
0!
0$
0-
02
#7610000000
1!
1$
1-
b101111101 1
12
b101111101 6
#7620000000
0!
0$
0-
02
#7630000000
1!
1$
1-
b101111110 1
12
b101111110 6
#7640000000
0!
0$
0-
02
#7650000000
1!
1$
1-
b101111111 1
12
b101111111 6
#7660000000
0!
0$
0-
02
#7670000000
1!
1$
1-
b110000000 1
12
b110000000 6
#7680000000
0!
0$
0-
02
#7690000000
1!
1$
1-
b110000001 1
12
b110000001 6
#7700000000
0!
0$
0-
02
#7710000000
1!
1$
1-
b110000010 1
12
b110000010 6
#7720000000
0!
0$
0-
02
#7730000000
1!
1$
1-
b110000011 1
12
b110000011 6
#7740000000
0!
0$
0-
02
#7750000000
1!
1$
1-
b110000100 1
12
b110000100 6
#7760000000
0!
0$
0-
02
#7770000000
1!
1$
1-
b110000101 1
12
b110000101 6
#7780000000
0!
0$
0-
02
#7790000000
1!
1$
1-
b110000110 1
12
b110000110 6
#7800000000
0!
0$
0-
02
#7810000000
1!
1$
1-
b110000111 1
12
b110000111 6
#7820000000
0!
0$
0-
02
#7830000000
1!
1$
1-
b110001000 1
12
b110001000 6
#7840000000
0!
0$
0-
02
#7850000000
1!
1$
1-
b110001001 1
12
b110001001 6
#7860000000
0!
0$
0-
02
#7870000000
1!
1$
1-
b110001010 1
12
b110001010 6
#7880000000
0!
0$
0-
02
#7890000000
1!
1$
1-
b110001011 1
12
b110001011 6
#7900000000
0!
0$
0-
02
#7910000000
1!
1$
1-
b110001100 1
12
b110001100 6
#7920000000
0!
0$
0-
02
#7930000000
1!
1$
1-
b110001101 1
12
b110001101 6
#7940000000
0!
0$
0-
02
#7950000000
1!
1$
1-
b110001110 1
12
b110001110 6
#7960000000
0!
0$
0-
02
#7970000000
1!
1$
1-
b110001111 1
12
b110001111 6
#7980000000
0!
0$
0-
02
#7990000000
1!
1$
1-
b110010000 1
12
b110010000 6
#8000000000
0!
0$
0-
02
#8010000000
1!
1$
1-
b110010001 1
12
b110010001 6
#8020000000
0!
0$
0-
02
#8030000000
1!
1$
1-
b110010010 1
12
b110010010 6
#8040000000
0!
0$
0-
02
#8050000000
1!
1$
1-
b110010011 1
12
b110010011 6
#8060000000
0!
0$
0-
02
#8070000000
1!
1$
1-
b110010100 1
12
b110010100 6
#8080000000
0!
0$
0-
02
#8090000000
1!
1$
1-
b110010101 1
12
b110010101 6
#8100000000
0!
0$
0-
02
#8110000000
1!
1$
1-
b110010110 1
12
b110010110 6
#8120000000
0!
0$
0-
02
#8130000000
1!
1$
1-
b110010111 1
12
b110010111 6
#8140000000
0!
0$
0-
02
#8150000000
1!
1$
1-
b110011000 1
12
b110011000 6
#8160000000
0!
0$
0-
02
#8170000000
1!
1$
1-
b110011001 1
12
b110011001 6
#8180000000
0!
0$
0-
02
#8190000000
1!
1$
1-
b110011010 1
12
b110011010 6
#8200000000
0!
0$
0-
02
#8210000000
1!
1$
1-
b110011011 1
12
b110011011 6
#8220000000
0!
1"
0$
1%
0-
02
#8230000000
1!
1$
1-
b110011100 1
12
b110011100 6
#8240000000
0!
0$
0-
02
#8250000000
1!
1$
1-
b110011101 1
12
b110011101 6
#8260000000
0!
0$
0-
02
#8270000000
1!
1$
1-
b110011110 1
12
b110011110 6
#8280000000
0!
0$
0-
02
#8290000000
1!
1$
1-
b110011111 1
12
b110011111 6
#8300000000
0!
0$
0-
02
#8310000000
1!
1$
1-
b110100000 1
12
b110100000 6
#8320000000
0!
0$
0-
02
#8330000000
1!
1$
1-
b110100001 1
12
b110100001 6
#8340000000
0!
0$
0-
02
#8350000000
1!
1$
1-
b110100010 1
12
b110100010 6
#8360000000
0!
0$
0-
02
#8370000000
1!
1$
1-
b110100011 1
12
b110100011 6
#8380000000
0!
0$
0-
02
#8390000000
1!
1$
1-
b110100100 1
12
b110100100 6
#8400000000
0!
0$
0-
02
#8410000000
1!
1$
1-
b110100101 1
12
b110100101 6
#8420000000
0!
0$
0-
02
#8430000000
1!
1$
1-
b110100110 1
12
b110100110 6
#8440000000
0!
0$
0-
02
#8450000000
1!
1$
1-
b110100111 1
12
b110100111 6
#8460000000
0!
0$
0-
02
#8470000000
1!
1$
1-
b110101000 1
12
b110101000 6
#8480000000
0!
0$
0-
02
#8490000000
1!
1$
1-
b110101001 1
12
b110101001 6
#8500000000
0!
0$
0-
02
#8510000000
1!
1$
1-
b110101010 1
12
b110101010 6
#8520000000
0!
0$
0-
02
#8530000000
1!
1$
1-
b110101011 1
12
b110101011 6
#8540000000
0!
0"
0$
0%
0-
02
#8550000000
1!
1$
1-
b110101100 1
12
b110101100 6
#8560000000
0!
0$
0-
02
#8570000000
1!
1$
1-
b110101101 1
12
b110101101 6
#8580000000
0!
0$
0-
02
#8590000000
1!
1$
1-
b110101110 1
12
b110101110 6
#8600000000
0!
0$
0-
02
#8610000000
1!
1$
1-
b110101111 1
12
b110101111 6
#8620000000
0!
0$
0-
02
#8630000000
1!
1$
1-
b110110000 1
12
b110110000 6
#8640000000
0!
0$
0-
02
#8650000000
1!
1$
1-
b110110001 1
12
b110110001 6
#8660000000
0!
0$
0-
02
#8670000000
1!
1$
1-
b110110010 1
12
b110110010 6
#8680000000
0!
0$
0-
02
#8690000000
1!
1$
1-
b110110011 1
12
b110110011 6
#8700000000
0!
0$
0-
02
#8710000000
1!
1$
1-
b110110100 1
12
b110110100 6
#8720000000
0!
0$
0-
02
#8730000000
1!
1$
1-
b110110101 1
12
b110110101 6
#8740000000
0!
0$
0-
02
#8750000000
1!
1$
1-
b110110110 1
12
b110110110 6
#8760000000
0!
0$
0-
02
#8770000000
1!
1$
1-
b110110111 1
12
b110110111 6
#8780000000
0!
0$
0-
02
#8790000000
1!
1$
1-
b110111000 1
12
b110111000 6
#8800000000
0!
0$
0-
02
#8810000000
1!
1$
1-
b110111001 1
12
b110111001 6
#8820000000
0!
0$
0-
02
#8830000000
1!
1$
1-
b110111010 1
12
b110111010 6
#8840000000
0!
0$
0-
02
#8850000000
1!
1$
1-
b110111011 1
12
b110111011 6
#8860000000
0!
0$
0-
02
#8870000000
1!
1$
1-
b110111100 1
12
b110111100 6
#8880000000
0!
0$
0-
02
#8890000000
1!
1$
1-
b110111101 1
12
b110111101 6
#8900000000
0!
0$
0-
02
#8910000000
1!
1$
1-
b110111110 1
12
b110111110 6
#8920000000
0!
0$
0-
02
#8930000000
1!
1$
1-
b110111111 1
12
b110111111 6
#8940000000
0!
0$
0-
02
#8950000000
1!
1$
1-
b111000000 1
12
b111000000 6
#8960000000
0!
0$
0-
02
#8970000000
1!
1$
1-
b111000001 1
12
b111000001 6
#8980000000
0!
0$
0-
02
#8990000000
1!
1$
1-
b111000010 1
12
b111000010 6
#9000000000
0!
0$
0-
02
#9010000000
1!
1$
1-
b111000011 1
12
b111000011 6
#9020000000
0!
0$
0-
02
#9030000000
1!
1$
1-
b111000100 1
12
b111000100 6
#9040000000
0!
0$
0-
02
#9050000000
1!
1$
1-
b111000101 1
12
b111000101 6
#9060000000
0!
0$
0-
02
#9070000000
1!
1$
1-
b111000110 1
12
b111000110 6
#9080000000
0!
0$
0-
02
#9090000000
1!
1$
1-
b111000111 1
12
b111000111 6
#9100000000
0!
0$
0-
02
#9110000000
1!
1$
1-
b111001000 1
12
b111001000 6
#9120000000
0!
0$
0-
02
#9130000000
1!
1$
1-
b111001001 1
12
b111001001 6
#9140000000
0!
0$
0-
02
#9150000000
1!
1$
1-
b111001010 1
12
b111001010 6
#9160000000
0!
0$
0-
02
#9170000000
1!
1$
1-
b111001011 1
12
b111001011 6
#9180000000
0!
0$
0-
02
#9190000000
1!
1$
1-
b111001100 1
12
b111001100 6
#9200000000
0!
0$
0-
02
#9210000000
1!
1$
1-
b111001101 1
12
b111001101 6
#9220000000
0!
0$
0-
02
#9230000000
1!
1$
1-
b111001110 1
12
b111001110 6
#9240000000
0!
0$
0-
02
#9250000000
1!
1$
1-
b111001111 1
12
b111001111 6
#9260000000
0!
0$
0-
02
#9270000000
1!
1$
1-
b111010000 1
12
b111010000 6
#9280000000
0!
0$
0-
02
#9290000000
1!
1$
1-
b111010001 1
12
b111010001 6
#9300000000
0!
0$
0-
02
#9310000000
1!
1$
1-
b111010010 1
12
b111010010 6
#9320000000
0!
0$
0-
02
#9330000000
1!
1$
1-
b111010011 1
12
b111010011 6
#9340000000
0!
0$
0-
02
#9350000000
1!
1$
1-
b111010100 1
12
b111010100 6
#9360000000
0!
0$
0-
02
#9370000000
1!
1$
1-
b111010101 1
12
b111010101 6
#9380000000
0!
0$
0-
02
#9390000000
1!
1$
1-
b111010110 1
12
b111010110 6
#9400000000
0!
0$
0-
02
#9410000000
1!
1$
1-
b111010111 1
12
b111010111 6
#9420000000
0!
0$
0-
02
#9430000000
1!
1$
1-
b111011000 1
12
b111011000 6
#9440000000
0!
0$
0-
02
#9450000000
1!
1$
1-
b111011001 1
12
b111011001 6
#9460000000
0!
0$
0-
02
#9470000000
1!
1$
1-
b111011010 1
12
b111011010 6
#9480000000
0!
0$
0-
02
#9490000000
1!
1$
1-
b111011011 1
12
b111011011 6
#9500000000
0!
0$
0-
02
#9510000000
1!
1$
1-
b111011100 1
12
b111011100 6
#9520000000
0!
0$
0-
02
#9530000000
1!
1$
1-
b111011101 1
12
b111011101 6
#9540000000
0!
0$
0-
02
#9550000000
1!
1$
1-
b111011110 1
12
b111011110 6
#9560000000
0!
0$
0-
02
#9570000000
1!
1$
1-
b111011111 1
12
b111011111 6
#9580000000
0!
1"
0$
1%
0-
02
#9590000000
1!
1$
1-
b111100000 1
12
b111100000 6
#9600000000
0!
0$
0-
02
#9610000000
1!
1$
1-
b111100001 1
12
b111100001 6
#9620000000
0!
0$
0-
02
#9630000000
1!
1$
1-
b111100010 1
12
b111100010 6
#9640000000
0!
0$
0-
02
#9650000000
1!
1$
1-
b111100011 1
12
b111100011 6
#9660000000
0!
0$
0-
02
#9670000000
1!
1$
1-
b111100100 1
12
b111100100 6
#9680000000
0!
0$
0-
02
#9690000000
1!
1$
1-
b111100101 1
12
b111100101 6
#9700000000
0!
0$
0-
02
#9710000000
1!
1$
1-
b111100110 1
12
b111100110 6
#9720000000
0!
0$
0-
02
#9730000000
1!
1$
1-
b111100111 1
12
b111100111 6
#9740000000
0!
0$
0-
02
#9750000000
1!
1$
1-
b111101000 1
12
b111101000 6
#9760000000
0!
0$
0-
02
#9770000000
1!
1$
1-
b111101001 1
12
b111101001 6
#9780000000
0!
0$
0-
02
#9790000000
1!
1$
1-
b111101010 1
12
b111101010 6
#9800000000
0!
0$
0-
02
#9810000000
1!
1$
1-
b111101011 1
12
b111101011 6
#9820000000
0!
0$
0-
02
#9830000000
1!
1$
1-
b111101100 1
12
b111101100 6
#9840000000
0!
0$
0-
02
#9850000000
1!
1$
1-
b111101101 1
12
b111101101 6
#9860000000
0!
0$
0-
02
#9870000000
1!
1$
1-
b111101110 1
12
b111101110 6
#9880000000
0!
0$
0-
02
#9890000000
1!
1$
1-
b111101111 1
12
b111101111 6
#9900000000
0!
0"
0$
0%
0-
02
#9910000000
1!
1$
1-
b111110000 1
12
b111110000 6
#9920000000
0!
0$
0-
02
#9930000000
1!
1$
1-
b111110001 1
12
b111110001 6
#9940000000
0!
0$
0-
02
#9950000000
1!
1$
1-
b111110010 1
12
b111110010 6
#9960000000
0!
0$
0-
02
#9970000000
1!
1$
1-
b111110011 1
12
b111110011 6
#9980000000
0!
0$
0-
02
#9990000000
1!
1$
1-
b111110100 1
12
b111110100 6
#10000000000
0!
0$
0-
02
