$date
  Sun May 05 01:54:29 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp3_2 $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 1 # up $end
$var reg 1 $ down $end
$var reg 4 % enable_disp[3:0] $end
$var reg 7 & segmentos[6:0] $end
$scope module uut $end
$var reg 1 ' clk $end
$var reg 1 ( reset $end
$var reg 1 ) up $end
$var reg 1 * down $end
$var reg 4 + enable_disp[3:0] $end
$var reg 7 , segmentos[6:0] $end
$var reg 1 - debounced_reset $end
$var reg 1 . debounced_up $end
$var reg 1 / debounced_down $end
$var reg 4 0 dig3[3:0] $end
$var reg 4 1 dig2[3:0] $end
$var reg 4 2 dig1[3:0] $end
$var reg 4 3 dig0[3:0] $end
$scope module a $end
$var reg 1 4 clk $end
$var reg 1 5 key $end
$var reg 1 6 debounced_key $end
$var reg 1 7 key_stable $end
$var reg 1 8 last_key $end
$upscope $end
$scope module b $end
$var reg 1 9 clk $end
$var reg 1 : key $end
$var reg 1 ; debounced_key $end
$var reg 1 < key_stable $end
$var reg 1 = last_key $end
$upscope $end
$scope module c $end
$var reg 1 > clk $end
$var reg 1 ? key $end
$var reg 1 @ debounced_key $end
$var reg 1 A key_stable $end
$var reg 1 B last_key $end
$upscope $end
$scope module d $end
$var reg 1 C clk $end
$var reg 1 D reset $end
$var reg 4 E dig3[3:0] $end
$var reg 4 F dig2[3:0] $end
$var reg 4 G dig1[3:0] $end
$var reg 4 H dig0[3:0] $end
$var reg 4 I enable_disp[3:0] $end
$var reg 7 J segmentos[6:0] $end
$comment state is not handled $end
$var integer 32 K cuenta $end
$var reg 1 L debounced_reset $end
$var reg 1 M enable_conta $end
$var reg 4 N bcd[3:0] $end
$scope module a $end
$var reg 1 O clk $end
$var reg 1 P key $end
$var reg 1 Q debounced_key $end
$var reg 1 R key_stable $end
$var reg 1 S last_key $end
$upscope $end
$scope module b $end
$var reg 1 T clk $end
$var reg 1 U reset $end
$var reg 1 V enable $end
$var reg 1 W cout $end
$var integer 32 X q $end
$upscope $end
$scope module d $end
$var reg 7 Y segmentos[6:0] $end
$var reg 4 Z bcd[3:0] $end
$upscope $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
0#
0$
b0001 %
b0111000 &
0'
0(
0)
0*
b0001 +
b0111000 ,
U-
U.
U/
b0000 0
b0000 1
b0000 2
b0000 3
04
05
U6
U7
U8
09
0:
U;
U<
U=
0>
0?
U@
UA
UB
0C
UD
b0000 E
b0000 F
b0000 G
b0000 H
b0001 I
b0111000 J
b0 K
UL
1M
bUUUU N
0O
UP
UQ
UR
US
0T
UU
1V
UW
b0 X
b0111000 Y
bUUUU Z
#10000000
1!
1'
0-
0.
0/
14
06
07
08
19
0;
0<
0=
1>
0@
0A
0B
1C
0D
1O
0P
1T
0W
#20000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#30000000
1!
1'
14
19
1>
1C
0L
1O
0Q
0R
0S
1T
0U
#40000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#50000000
1!
1'
14
19
1>
1C
1O
1T
1W
#60000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#70000000
1!
1'
14
19
1>
1C
1O
1T
#80000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#90000000
1!
1'
14
19
1>
1C
1O
1T
#100000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#110000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#120000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#130000000
1!
1'
14
19
1>
1C
1O
1T
#140000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#150000000
1!
1'
14
19
1>
1C
1O
1T
#160000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#170000000
1!
1'
14
19
1>
1C
1O
1T
1W
#180000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#190000000
1!
1'
14
19
1>
1C
1O
1T
#200000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#210000000
1!
1'
14
19
1>
1C
1O
1T
#220000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#230000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#240000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#250000000
1!
1'
14
19
1>
1C
1O
1T
#260000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#270000000
1!
1'
14
19
1>
1C
1O
1T
#280000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#290000000
1!
1'
14
19
1>
1C
1O
1T
1W
#300000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#310000000
1!
1'
14
19
1>
1C
1O
1T
#320000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#330000000
1!
1'
14
19
1>
1C
1O
1T
#340000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#350000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#360000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#370000000
1!
1'
14
19
1>
1C
1O
1T
#380000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#390000000
1!
1'
14
19
1>
1C
1O
1T
#400000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#410000000
1!
1'
14
19
1>
1C
1O
1T
1W
#420000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#430000000
1!
1'
14
19
1>
1C
1O
1T
#440000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#450000000
1!
1'
14
19
1>
1C
1O
1T
#460000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#470000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#480000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#490000000
1!
1'
14
19
1>
1C
1O
1T
#500000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#510000000
1!
1'
14
19
1>
1C
1O
1T
#520000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#530000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
1W
#540000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#550000000
1!
1'
b0001 3
14
19
1>
1C
b0001 H
1O
1T
#560000000
0!
0#
0'
0)
04
09
0:
0>
0C
b100 K
0O
0T
b100 X
#570000000
#580000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#590000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#600000000
1!
b0010 %
1'
b0010 +
14
19
1>
1C
b0010 I
1O
1T
0W
#610000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#620000000
1!
1'
14
19
1>
1C
1O
1T
#630000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#640000000
1!
1'
14
19
1>
1C
1O
1T
#650000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#660000000
1!
1'
14
19
1>
1C
1O
1T
1W
#670000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#680000000
1!
1'
14
19
1>
1C
1O
1T
#690000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#700000000
1!
1'
14
19
1>
1C
1O
1T
#710000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#720000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#730000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#740000000
1!
1'
14
19
1>
1C
1O
1T
#750000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#760000000
1!
1'
14
19
1>
1C
1O
1T
#770000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#780000000
1!
1'
14
19
1>
1C
1O
1T
1W
#790000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#800000000
1!
1'
14
19
1>
1C
1O
1T
#810000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#820000000
1!
1'
14
19
1>
1C
1O
1T
#830000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#840000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#850000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#860000000
1!
1'
14
19
1>
1C
1O
1T
#870000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#880000000
1!
1'
14
19
1>
1C
1O
1T
#890000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#900000000
1!
1'
14
19
1>
1C
1O
1T
1W
#910000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#920000000
1!
1'
14
19
1>
1C
1O
1T
#930000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#940000000
1!
1'
14
19
1>
1C
1O
1T
#950000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#960000000
1!
b0001 %
b1001111 &
1'
b0001 +
b1001111 ,
14
19
1>
1C
b0001 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#970000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#980000000
1!
1'
14
19
1>
1C
1O
1T
#990000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#1000000000
1!
1'
14
19
1>
1C
1O
1T
#1010000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#1020000000
1!
1'
14
19
1>
1C
1O
1T
1W
#1030000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#1040000000
1!
1'
14
19
1>
1C
1O
1T
#1050000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#1060000000
1!
1'
14
19
1>
1C
1O
1T
#1070000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#1080000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#1090000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#1100000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#1110000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#1120000000
1!
1'
b0010 3
14
19
1>
1C
b0010 H
1O
1T
#1130000000
0!
0#
0'
0)
04
09
0:
0>
0C
b10 K
0O
0T
b10 X
#1140000000
#1150000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
1W
#1160000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#1170000000
1!
1'
14
19
1>
1C
1O
1T
#1180000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#1190000000
1!
1'
14
19
1>
1C
1O
1T
#1200000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#1210000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#1220000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#1230000000
1!
1'
14
19
1>
1C
1O
1T
#1240000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#1250000000
1!
1'
14
19
1>
1C
1O
1T
#1260000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#1270000000
1!
1'
14
19
1>
1C
1O
1T
1W
#1280000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#1290000000
1!
1'
14
19
1>
1C
1O
1T
#1300000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#1310000000
1!
1'
14
19
1>
1C
1O
1T
#1320000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#1330000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#1340000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#1350000000
1!
1'
14
19
1>
1C
1O
1T
#1360000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#1370000000
1!
1'
14
19
1>
1C
1O
1T
#1380000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#1390000000
1!
1'
14
19
1>
1C
1O
1T
1W
#1400000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#1410000000
1!
1'
14
19
1>
1C
1O
1T
#1420000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#1430000000
1!
1'
14
19
1>
1C
1O
1T
#1440000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#1450000000
1!
b0001 %
b0010010 &
1'
b0001 +
b0010010 ,
14
19
1>
1C
b0001 I
b0010010 J
b0010 N
1O
1T
0W
b0010010 Y
b0010 Z
#1460000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#1470000000
1!
1'
14
19
1>
1C
1O
1T
#1480000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#1490000000
1!
1'
14
19
1>
1C
1O
1T
#1500000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#1510000000
1!
1'
14
19
1>
1C
1O
1T
1W
#1520000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#1530000000
1!
1'
14
19
1>
1C
1O
1T
#1540000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#1550000000
1!
1'
14
19
1>
1C
1O
1T
#1560000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#1570000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#1580000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#1590000000
1!
1'
14
19
1>
1C
1O
1T
#1600000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#1610000000
1!
1'
14
19
1>
1C
1O
1T
#1620000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#1630000000
1!
1'
14
19
1>
1C
1O
1T
1W
#1640000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#1650000000
1!
1'
14
19
1>
1C
1O
1T
#1660000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#1670000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#1680000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#1690000000
1!
b0100 %
1'
b0100 +
b0011 3
14
19
1>
1C
b0011 H
b0100 I
1O
1T
0W
#1700000000
0!
0#
0'
0)
04
09
0:
0>
0C
b0 K
0O
0T
b0 X
#1710000000
#1720000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#1730000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#1740000000
1!
1'
14
19
1>
1C
1O
1T
#1750000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#1760000000
1!
1'
14
19
1>
1C
1O
1T
1W
#1770000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#1780000000
1!
1'
14
19
1>
1C
1O
1T
#1790000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#1800000000
1!
1'
14
19
1>
1C
1O
1T
#1810000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#1820000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#1830000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#1840000000
1!
1'
14
19
1>
1C
1O
1T
#1850000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#1860000000
1!
1'
14
19
1>
1C
1O
1T
#1870000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#1880000000
1!
1'
14
19
1>
1C
1O
1T
1W
#1890000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#1900000000
1!
1'
14
19
1>
1C
1O
1T
#1910000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#1920000000
1!
1'
14
19
1>
1C
1O
1T
#1930000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#1940000000
1!
b0001 %
b0000110 &
1'
b0001 +
b0000110 ,
14
19
1>
1C
b0001 I
b0000110 J
b0011 N
1O
1T
0W
b0000110 Y
b0011 Z
#1950000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#1960000000
1!
1'
14
19
1>
1C
1O
1T
#1970000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#1980000000
1!
1'
14
19
1>
1C
1O
1T
#1990000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#2000000000
1!
1'
14
19
1>
1C
1O
1T
1W
#2010000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#2020000000
1!
1'
14
19
1>
1C
1O
1T
#2030000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#2040000000
1!
1'
14
19
1>
1C
1O
1T
#2050000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#2060000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#2070000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#2080000000
1!
1'
14
19
1>
1C
1O
1T
#2090000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#2100000000
1!
1'
14
19
1>
1C
1O
1T
#2110000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#2120000000
1!
1'
14
19
1>
1C
1O
1T
1W
#2130000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#2140000000
1!
1'
14
19
1>
1C
1O
1T
#2150000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#2160000000
1!
1'
14
19
1>
1C
1O
1T
#2170000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#2180000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#2190000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#2200000000
1!
1'
14
19
1>
1C
1O
1T
#2210000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#2220000000
1!
1'
14
19
1>
1C
1O
1T
#2230000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#2240000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
1W
#2250000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#2260000000
1!
1'
b0100 3
14
19
1>
1C
b0100 H
1O
1T
#2270000000
0!
0#
0'
0)
04
09
0:
0>
0C
b100 K
0O
0T
b100 X
#2280000000
#2290000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#2300000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#2310000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#2320000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#2330000000
1!
1'
14
19
1>
1C
1O
1T
#2340000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#2350000000
1!
1'
14
19
1>
1C
1O
1T
#2360000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#2370000000
1!
1'
14
19
1>
1C
1O
1T
1W
#2380000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#2390000000
1!
1'
14
19
1>
1C
1O
1T
#2400000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#2410000000
1!
1'
14
19
1>
1C
1O
1T
#2420000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#2430000000
1!
b0001 %
b1001100 &
1'
b0001 +
b1001100 ,
14
19
1>
1C
b0001 I
b1001100 J
b0100 N
1O
1T
0W
b1001100 Y
b0100 Z
#2440000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#2450000000
1!
1'
14
19
1>
1C
1O
1T
#2460000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#2470000000
1!
1'
14
19
1>
1C
1O
1T
#2480000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#2490000000
1!
1'
14
19
1>
1C
1O
1T
1W
#2500000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#2510000000
1!
1'
14
19
1>
1C
1O
1T
#2520000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#2530000000
1!
1'
14
19
1>
1C
1O
1T
#2540000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#2550000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#2560000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#2570000000
1!
1'
14
19
1>
1C
1O
1T
#2580000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#2590000000
1!
1'
14
19
1>
1C
1O
1T
#2600000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#2610000000
1!
1'
14
19
1>
1C
1O
1T
1W
#2620000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#2630000000
1!
1'
14
19
1>
1C
1O
1T
#2640000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#2650000000
1!
1'
14
19
1>
1C
1O
1T
#2660000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#2670000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#2680000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#2690000000
1!
1'
14
19
1>
1C
1O
1T
#2700000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#2710000000
1!
1'
14
19
1>
1C
1O
1T
#2720000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#2730000000
1!
1'
14
19
1>
1C
1O
1T
1W
#2740000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#2750000000
1!
1'
14
19
1>
1C
1O
1T
#2760000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#2770000000
1!
1'
14
19
1>
1C
1O
1T
#2780000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#2790000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#2800000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#2810000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#2820000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#2830000000
1!
1'
b0101 3
14
19
1>
1C
b0101 H
1O
1T
#2840000000
0!
0#
0'
0)
04
09
0:
0>
0C
b10 K
0O
0T
b10 X
#2850000000
#2860000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
1W
#2870000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#2880000000
1!
1'
14
19
1>
1C
1O
1T
#2890000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#2900000000
1!
1'
14
19
1>
1C
1O
1T
#2910000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#2920000000
1!
b0001 %
b0100100 &
1'
b0001 +
b0100100 ,
14
19
1>
1C
b0001 I
b0100100 J
b0101 N
1O
1T
0W
b0100100 Y
b0101 Z
#2930000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#2940000000
1!
1'
14
19
1>
1C
1O
1T
#2950000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#2960000000
1!
1'
14
19
1>
1C
1O
1T
#2970000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#2980000000
1!
1'
14
19
1>
1C
1O
1T
1W
#2990000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#3000000000
1!
1'
14
19
1>
1C
1O
1T
#3010000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#3020000000
1!
1'
14
19
1>
1C
1O
1T
#3030000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#3040000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#3050000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#3060000000
1!
1'
14
19
1>
1C
1O
1T
#3070000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#3080000000
1!
1'
14
19
1>
1C
1O
1T
#3090000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#3100000000
1!
1'
14
19
1>
1C
1O
1T
1W
#3110000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#3120000000
1!
1'
14
19
1>
1C
1O
1T
#3130000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#3140000000
1!
1'
14
19
1>
1C
1O
1T
#3150000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#3160000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#3170000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#3180000000
1!
1'
14
19
1>
1C
1O
1T
#3190000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#3200000000
1!
1'
14
19
1>
1C
1O
1T
#3210000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#3220000000
1!
1'
14
19
1>
1C
1O
1T
1W
#3230000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#3240000000
1!
1'
14
19
1>
1C
1O
1T
#3250000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#3260000000
1!
1'
14
19
1>
1C
1O
1T
#3270000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#3280000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#3290000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#3300000000
1!
1'
14
19
1>
1C
1O
1T
#3310000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#3320000000
1!
1'
14
19
1>
1C
1O
1T
#3330000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#3340000000
1!
1'
14
19
1>
1C
1O
1T
1W
#3350000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#3360000000
1!
1'
14
19
1>
1C
1O
1T
#3370000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#3380000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#3390000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#3400000000
1!
b0001 %
b0100000 &
1'
b0001 +
b0100000 ,
b0110 3
14
19
1>
1C
b0110 H
b0001 I
b0100000 J
b0110 N
1O
1T
0W
b0100000 Y
b0110 Z
#3410000000
0!
0#
0'
0)
04
09
0:
0>
0C
b0 K
0O
0T
b0 X
#3420000000
#3430000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#3440000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#3450000000
1!
1'
14
19
1>
1C
1O
1T
#3460000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#3470000000
1!
1'
14
19
1>
1C
1O
1T
1W
#3480000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#3490000000
1!
1'
14
19
1>
1C
1O
1T
#3500000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#3510000000
1!
1'
14
19
1>
1C
1O
1T
#3520000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#3530000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#3540000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#3550000000
1!
1'
14
19
1>
1C
1O
1T
#3560000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#3570000000
1!
1'
14
19
1>
1C
1O
1T
#3580000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#3590000000
1!
1'
14
19
1>
1C
1O
1T
1W
#3600000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#3610000000
1!
1'
14
19
1>
1C
1O
1T
#3620000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#3630000000
1!
1'
14
19
1>
1C
1O
1T
#3640000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#3650000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#3660000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#3670000000
1!
1'
14
19
1>
1C
1O
1T
#3680000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#3690000000
1!
1'
14
19
1>
1C
1O
1T
#3700000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#3710000000
1!
1'
14
19
1>
1C
1O
1T
1W
#3720000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#3730000000
1!
1'
14
19
1>
1C
1O
1T
#3740000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#3750000000
1!
1'
14
19
1>
1C
1O
1T
#3760000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#3770000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#3780000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#3790000000
1!
1'
14
19
1>
1C
1O
1T
#3800000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#3810000000
1!
1'
14
19
1>
1C
1O
1T
#3820000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#3830000000
1!
1'
14
19
1>
1C
1O
1T
1W
#3840000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#3850000000
1!
1'
14
19
1>
1C
1O
1T
#3860000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#3870000000
1!
1'
14
19
1>
1C
1O
1T
#3880000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#3890000000
1!
b0001 %
b0100000 &
1'
b0001 +
b0100000 ,
14
19
1>
1C
b0001 I
b0100000 J
b0110 N
1O
1T
0W
b0100000 Y
b0110 Z
#3900000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#3910000000
1!
1'
14
19
1>
1C
1O
1T
#3920000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#3930000000
1!
1'
14
19
1>
1C
1O
1T
#3940000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#3950000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
1W
#3960000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#3970000000
1!
1'
b0111 3
14
19
1>
1C
b0111 H
1O
1T
#3980000000
0!
0#
0'
0)
04
09
0:
0>
0C
b100 K
0O
0T
b100 X
#3990000000
#4000000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#4010000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#4020000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#4030000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#4040000000
1!
1'
14
19
1>
1C
1O
1T
#4050000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#4060000000
1!
1'
14
19
1>
1C
1O
1T
#4070000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#4080000000
1!
1'
14
19
1>
1C
1O
1T
1W
#4090000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#4100000000
1!
1'
14
19
1>
1C
1O
1T
#4110000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#4120000000
1!
1'
14
19
1>
1C
1O
1T
#4130000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#4140000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#4150000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#4160000000
1!
1'
14
19
1>
1C
1O
1T
#4170000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#4180000000
1!
1'
14
19
1>
1C
1O
1T
#4190000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#4200000000
1!
1'
14
19
1>
1C
1O
1T
1W
#4210000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#4220000000
1!
1'
14
19
1>
1C
1O
1T
#4230000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#4240000000
1!
1'
14
19
1>
1C
1O
1T
#4250000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#4260000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#4270000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#4280000000
1!
1'
14
19
1>
1C
1O
1T
#4290000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#4300000000
1!
1'
14
19
1>
1C
1O
1T
#4310000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#4320000000
1!
1'
14
19
1>
1C
1O
1T
1W
#4330000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#4340000000
1!
1'
14
19
1>
1C
1O
1T
#4350000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#4360000000
1!
1'
14
19
1>
1C
1O
1T
#4370000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#4380000000
1!
b0001 %
b0001111 &
1'
b0001 +
b0001111 ,
14
19
1>
1C
b0001 I
b0001111 J
b0111 N
1O
1T
0W
b0001111 Y
b0111 Z
#4390000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#4400000000
1!
1'
14
19
1>
1C
1O
1T
#4410000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#4420000000
1!
1'
14
19
1>
1C
1O
1T
#4430000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#4440000000
1!
1'
14
19
1>
1C
1O
1T
1W
#4450000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#4460000000
1!
1'
14
19
1>
1C
1O
1T
#4470000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#4480000000
1!
1'
14
19
1>
1C
1O
1T
#4490000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#4500000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#4510000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#4520000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#4530000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#4540000000
1!
1'
b1000 3
14
19
1>
1C
b1000 H
1O
1T
#4550000000
0!
0#
0'
0)
04
09
0:
0>
0C
b10 K
0O
0T
b10 X
#4560000000
#4570000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
1W
#4580000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#4590000000
1!
1'
14
19
1>
1C
1O
1T
#4600000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#4610000000
1!
1'
14
19
1>
1C
1O
1T
#4620000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#4630000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#4640000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#4650000000
1!
1'
14
19
1>
1C
1O
1T
#4660000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#4670000000
1!
1'
14
19
1>
1C
1O
1T
#4680000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#4690000000
1!
1'
14
19
1>
1C
1O
1T
1W
#4700000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#4710000000
1!
1'
14
19
1>
1C
1O
1T
#4720000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#4730000000
1!
1'
14
19
1>
1C
1O
1T
#4740000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#4750000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#4760000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#4770000000
1!
1'
14
19
1>
1C
1O
1T
#4780000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#4790000000
1!
1'
14
19
1>
1C
1O
1T
#4800000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#4810000000
1!
1'
14
19
1>
1C
1O
1T
1W
#4820000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#4830000000
1!
1'
14
19
1>
1C
1O
1T
#4840000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#4850000000
1!
1'
14
19
1>
1C
1O
1T
#4860000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#4870000000
1!
b0001 %
b0000000 &
1'
b0001 +
b0000000 ,
14
19
1>
1C
b0001 I
b0000000 J
b1000 N
1O
1T
0W
b0000000 Y
b1000 Z
#4880000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#4890000000
1!
1'
14
19
1>
1C
1O
1T
#4900000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#4910000000
1!
1'
14
19
1>
1C
1O
1T
#4920000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#4930000000
1!
1'
14
19
1>
1C
1O
1T
1W
#4940000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#4950000000
1!
1'
14
19
1>
1C
1O
1T
#4960000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#4970000000
1!
1'
14
19
1>
1C
1O
1T
#4980000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#4990000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#5000000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#5010000000
1!
1'
14
19
1>
1C
1O
1T
#5020000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#5030000000
1!
1'
14
19
1>
1C
1O
1T
#5040000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#5050000000
1!
1'
14
19
1>
1C
1O
1T
1W
#5060000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#5070000000
1!
1'
14
19
1>
1C
1O
1T
#5080000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#5090000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#5100000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#5110000000
1!
b0100 %
1'
b0100 +
b1001 3
14
19
1>
1C
b1001 H
b0100 I
1O
1T
0W
#5120000000
0!
0#
0'
0)
04
09
0:
0>
0C
b0 K
0O
0T
b0 X
#5130000000
#5140000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#5150000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#5160000000
1!
1'
14
19
1>
1C
1O
1T
#5170000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#5180000000
1!
1'
14
19
1>
1C
1O
1T
1W
#5190000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#5200000000
1!
1'
14
19
1>
1C
1O
1T
#5210000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#5220000000
1!
1'
14
19
1>
1C
1O
1T
#5230000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#5240000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#5250000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#5260000000
1!
1'
14
19
1>
1C
1O
1T
#5270000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#5280000000
1!
1'
14
19
1>
1C
1O
1T
#5290000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#5300000000
1!
1'
14
19
1>
1C
1O
1T
1W
#5310000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#5320000000
1!
1'
14
19
1>
1C
1O
1T
#5330000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#5340000000
1!
1'
14
19
1>
1C
1O
1T
#5350000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#5360000000
1!
b0001 %
b0000100 &
1'
b0001 +
b0000100 ,
14
19
1>
1C
b0001 I
b0000100 J
b1001 N
1O
1T
0W
b0000100 Y
b1001 Z
#5370000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#5380000000
1!
1'
14
19
1>
1C
1O
1T
#5390000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#5400000000
1!
1'
14
19
1>
1C
1O
1T
#5410000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#5420000000
1!
1'
14
19
1>
1C
1O
1T
1W
#5430000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#5440000000
1!
1'
14
19
1>
1C
1O
1T
#5450000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#5460000000
1!
1'
14
19
1>
1C
1O
1T
#5470000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#5480000000
1!
b0010 %
b0000001 &
1'
b0010 +
b0000001 ,
14
19
1>
1C
b0010 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#5490000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#5500000000
1!
1'
14
19
1>
1C
1O
1T
#5510000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#5520000000
1!
1'
14
19
1>
1C
1O
1T
#5530000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#5540000000
1!
1'
14
19
1>
1C
1O
1T
1W
#5550000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#5560000000
1!
1'
14
19
1>
1C
1O
1T
#5570000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#5580000000
1!
1'
14
19
1>
1C
1O
1T
#5590000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#5600000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1O
1T
0W
#5610000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#5620000000
1!
1'
14
19
1>
1C
1O
1T
#5630000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#5640000000
1!
1'
14
19
1>
1C
1O
1T
#5650000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#5660000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
1W
#5670000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#5680000000
1!
1'
b0001 2
b0000 3
14
19
1>
1C
b0001 G
b0000 H
1O
1T
#5690000000
0!
0#
0'
0)
04
09
0:
0>
0C
b100 K
0O
0T
b100 X
#5700000000
#5710000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#5720000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#5730000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#5740000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#5750000000
1!
1'
14
19
1>
1C
1O
1T
#5760000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#5770000000
1!
1'
14
19
1>
1C
1O
1T
#5780000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#5790000000
1!
1'
14
19
1>
1C
1O
1T
1W
#5800000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#5810000000
1!
1'
14
19
1>
1C
1O
1T
#5820000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#5830000000
1!
1'
14
19
1>
1C
1O
1T
#5840000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#5850000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#5860000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#5870000000
1!
1'
14
19
1>
1C
1O
1T
#5880000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#5890000000
1!
1'
14
19
1>
1C
1O
1T
#5900000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#5910000000
1!
1'
14
19
1>
1C
1O
1T
1W
#5920000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#5930000000
1!
1'
14
19
1>
1C
1O
1T
#5940000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#5950000000
1!
1'
14
19
1>
1C
1O
1T
#5960000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#5970000000
1!
b0010 %
b1001111 &
1'
b0010 +
b1001111 ,
14
19
1>
1C
b0010 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#5980000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#5990000000
1!
1'
14
19
1>
1C
1O
1T
#6000000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#6010000000
1!
1'
14
19
1>
1C
1O
1T
#6020000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#6030000000
1!
1'
14
19
1>
1C
1O
1T
1W
#6040000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#6050000000
1!
1'
14
19
1>
1C
1O
1T
#6060000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#6070000000
1!
1'
14
19
1>
1C
1O
1T
#6080000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#6090000000
1!
b0100 %
b0000001 &
1'
b0100 +
b0000001 ,
14
19
1>
1C
b0100 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#6100000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#6110000000
1!
1'
14
19
1>
1C
1O
1T
#6120000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#6130000000
1!
1'
14
19
1>
1C
1O
1T
#6140000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#6150000000
1!
1'
14
19
1>
1C
1O
1T
1W
#6160000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#6170000000
1!
1'
14
19
1>
1C
1O
1T
#6180000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#6190000000
1!
1'
14
19
1>
1C
1O
1T
#6200000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#6210000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#6220000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#6230000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#6240000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#6250000000
1!
1'
14
19
1>
1C
1O
1T
#6260000000
0!
0#
0'
0)
04
09
0:
0>
0C
b10 K
0O
0T
b10 X
#6270000000
#6280000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
1W
#6290000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#6300000000
1!
1'
14
19
1>
1C
1O
1T
#6310000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#6320000000
1!
1'
14
19
1>
1C
1O
1T
#6330000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#6340000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#6350000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#6360000000
1!
1'
14
19
1>
1C
1O
1T
#6370000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#6380000000
1!
1'
14
19
1>
1C
1O
1T
#6390000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#6400000000
1!
1'
14
19
1>
1C
1O
1T
1W
#6410000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#6420000000
1!
1'
14
19
1>
1C
1O
1T
#6430000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#6440000000
1!
1'
14
19
1>
1C
1O
1T
#6450000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#6460000000
1!
b0010 %
b1001111 &
1'
b0010 +
b1001111 ,
14
19
1>
1C
b0010 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#6470000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#6480000000
1!
1'
14
19
1>
1C
1O
1T
#6490000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#6500000000
1!
1'
14
19
1>
1C
1O
1T
#6510000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#6520000000
1!
1'
14
19
1>
1C
1O
1T
1W
#6530000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#6540000000
1!
1'
14
19
1>
1C
1O
1T
#6550000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#6560000000
1!
1'
14
19
1>
1C
1O
1T
#6570000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#6580000000
1!
b0100 %
b0000001 &
1'
b0100 +
b0000001 ,
14
19
1>
1C
b0100 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#6590000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#6600000000
1!
1'
14
19
1>
1C
1O
1T
#6610000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#6620000000
1!
1'
14
19
1>
1C
1O
1T
#6630000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#6640000000
1!
1'
14
19
1>
1C
1O
1T
1W
#6650000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#6660000000
1!
1'
14
19
1>
1C
1O
1T
#6670000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#6680000000
1!
1'
14
19
1>
1C
1O
1T
#6690000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#6700000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#6710000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#6720000000
1!
1'
14
19
1>
1C
1O
1T
#6730000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#6740000000
1!
1'
14
19
1>
1C
1O
1T
#6750000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#6760000000
1!
1'
14
19
1>
1C
1O
1T
1W
#6770000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#6780000000
1!
1'
14
19
1>
1C
1O
1T
#6790000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#6800000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#6810000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#6820000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#6830000000
0!
0#
0'
0)
04
09
0:
0>
0C
b0 K
0O
0T
b0 X
#6840000000
#6850000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#6860000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#6870000000
1!
1'
14
19
1>
1C
1O
1T
#6880000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#6890000000
1!
1'
14
19
1>
1C
1O
1T
1W
#6900000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#6910000000
1!
1'
14
19
1>
1C
1O
1T
#6920000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#6930000000
1!
1'
14
19
1>
1C
1O
1T
#6940000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#6950000000
1!
b0010 %
b1001111 &
1'
b0010 +
b1001111 ,
14
19
1>
1C
b0010 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#6960000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#6970000000
1!
1'
14
19
1>
1C
1O
1T
#6980000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#6990000000
1!
1'
14
19
1>
1C
1O
1T
#7000000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#7010000000
1!
1'
14
19
1>
1C
1O
1T
1W
#7020000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#7030000000
1!
1'
14
19
1>
1C
1O
1T
#7040000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#7050000000
1!
1'
14
19
1>
1C
1O
1T
#7060000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#7070000000
1!
b0100 %
b0000001 &
1'
b0100 +
b0000001 ,
14
19
1>
1C
b0100 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#7080000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#7090000000
1!
1'
14
19
1>
1C
1O
1T
#7100000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#7110000000
1!
1'
14
19
1>
1C
1O
1T
#7120000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#7130000000
1!
1'
14
19
1>
1C
1O
1T
1W
#7140000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#7150000000
1!
1'
14
19
1>
1C
1O
1T
#7160000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#7170000000
1!
1'
14
19
1>
1C
1O
1T
#7180000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#7190000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#7200000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#7210000000
1!
1'
14
19
1>
1C
1O
1T
#7220000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#7230000000
1!
1'
14
19
1>
1C
1O
1T
#7240000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#7250000000
1!
1'
14
19
1>
1C
1O
1T
1W
#7260000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#7270000000
1!
1'
14
19
1>
1C
1O
1T
#7280000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#7290000000
1!
1'
14
19
1>
1C
1O
1T
#7300000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#7310000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#7320000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#7330000000
1!
1'
14
19
1>
1C
1O
1T
#7340000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#7350000000
1!
1'
14
19
1>
1C
1O
1T
#7360000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#7370000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
1W
#7380000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#7390000000
1!
1'
14
19
1>
1C
1O
1T
#7400000000
0!
0#
0'
0)
04
09
0:
0>
0C
b100 K
0O
0T
b100 X
#7410000000
#7420000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#7430000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#7440000000
1!
b0010 %
b1001111 &
1'
b0010 +
b1001111 ,
14
19
1>
1C
b0010 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#7450000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#7460000000
1!
1'
14
19
1>
1C
1O
1T
#7470000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#7480000000
1!
1'
14
19
1>
1C
1O
1T
#7490000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#7500000000
1!
1'
14
19
1>
1C
1O
1T
1W
#7510000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#7520000000
1!
1'
14
19
1>
1C
1O
1T
#7530000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#7540000000
1!
1'
14
19
1>
1C
1O
1T
#7550000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#7560000000
1!
b0100 %
b0000001 &
1'
b0100 +
b0000001 ,
14
19
1>
1C
b0100 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#7570000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#7580000000
1!
1'
14
19
1>
1C
1O
1T
#7590000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#7600000000
1!
1'
14
19
1>
1C
1O
1T
#7610000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#7620000000
1!
1'
14
19
1>
1C
1O
1T
1W
#7630000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#7640000000
1!
1'
14
19
1>
1C
1O
1T
#7650000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#7660000000
1!
1'
14
19
1>
1C
1O
1T
#7670000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#7680000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#7690000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#7700000000
1!
1'
14
19
1>
1C
1O
1T
#7710000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#7720000000
1!
1'
14
19
1>
1C
1O
1T
#7730000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#7740000000
1!
1'
14
19
1>
1C
1O
1T
1W
#7750000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#7760000000
1!
1'
14
19
1>
1C
1O
1T
#7770000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#7780000000
1!
1'
14
19
1>
1C
1O
1T
#7790000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#7800000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#7810000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#7820000000
1!
1'
14
19
1>
1C
1O
1T
#7830000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#7840000000
1!
1'
14
19
1>
1C
1O
1T
#7850000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#7860000000
1!
1'
14
19
1>
1C
1O
1T
1W
#7870000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#7880000000
1!
1'
14
19
1>
1C
1O
1T
#7890000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#7900000000
1!
1'
14
19
1>
1C
1O
1T
#7910000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#7920000000
1!
b0010 %
b1001111 &
1'
b0010 +
b1001111 ,
14
19
1>
1C
b0010 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#7930000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#7940000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#7950000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#7960000000
1!
1'
14
19
1>
1C
1O
1T
#7970000000
0!
0#
0'
0)
04
09
0:
0>
0C
b10 K
0O
0T
b10 X
#7980000000
#7990000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
1W
#8000000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#8010000000
1!
1'
14
19
1>
1C
1O
1T
#8020000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#8030000000
1!
1'
14
19
1>
1C
1O
1T
#8040000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#8050000000
1!
b0100 %
b0000001 &
1'
b0100 +
b0000001 ,
14
19
1>
1C
b0100 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#8060000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#8070000000
1!
1'
14
19
1>
1C
1O
1T
#8080000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#8090000000
1!
1'
14
19
1>
1C
1O
1T
#8100000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#8110000000
1!
1'
14
19
1>
1C
1O
1T
1W
#8120000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#8130000000
1!
1'
14
19
1>
1C
1O
1T
#8140000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#8150000000
1!
1'
14
19
1>
1C
1O
1T
#8160000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#8170000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#8180000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#8190000000
1!
1'
14
19
1>
1C
1O
1T
#8200000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#8210000000
1!
1'
14
19
1>
1C
1O
1T
#8220000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#8230000000
1!
1'
14
19
1>
1C
1O
1T
1W
#8240000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#8250000000
1!
1'
14
19
1>
1C
1O
1T
#8260000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#8270000000
1!
1'
14
19
1>
1C
1O
1T
#8280000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#8290000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#8300000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#8310000000
1!
1'
14
19
1>
1C
1O
1T
#8320000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#8330000000
1!
1'
14
19
1>
1C
1O
1T
#8340000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#8350000000
1!
1'
14
19
1>
1C
1O
1T
1W
#8360000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#8370000000
1!
1'
14
19
1>
1C
1O
1T
#8380000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#8390000000
1!
1'
14
19
1>
1C
1O
1T
#8400000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#8410000000
1!
b0010 %
b1001111 &
1'
b0010 +
b1001111 ,
14
19
1>
1C
b0010 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#8420000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#8430000000
1!
1'
14
19
1>
1C
1O
1T
#8440000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#8450000000
1!
1'
14
19
1>
1C
1O
1T
#8460000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#8470000000
1!
1'
14
19
1>
1C
1O
1T
1W
#8480000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#8490000000
1!
1'
14
19
1>
1C
1O
1T
#8500000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#8510000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#8520000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#8530000000
1!
b0100 %
b0000001 &
1'
b0100 +
b0000001 ,
14
19
1>
1C
b0100 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#8540000000
0!
0#
0'
0)
04
09
0:
0>
0C
b0 K
0O
0T
b0 X
#8550000000
#8560000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#8570000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#8580000000
1!
1'
14
19
1>
1C
1O
1T
#8590000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#8600000000
1!
1'
14
19
1>
1C
1O
1T
1W
#8610000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#8620000000
1!
1'
14
19
1>
1C
1O
1T
#8630000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#8640000000
1!
1'
14
19
1>
1C
1O
1T
#8650000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#8660000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#8670000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#8680000000
1!
1'
14
19
1>
1C
1O
1T
#8690000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#8700000000
1!
1'
14
19
1>
1C
1O
1T
#8710000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#8720000000
1!
1'
14
19
1>
1C
1O
1T
1W
#8730000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#8740000000
1!
1'
14
19
1>
1C
1O
1T
#8750000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#8760000000
1!
1'
14
19
1>
1C
1O
1T
#8770000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#8780000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#8790000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#8800000000
1!
1'
14
19
1>
1C
1O
1T
#8810000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#8820000000
1!
1'
14
19
1>
1C
1O
1T
#8830000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#8840000000
1!
1'
14
19
1>
1C
1O
1T
1W
#8850000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#8860000000
1!
1'
14
19
1>
1C
1O
1T
#8870000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#8880000000
1!
1'
14
19
1>
1C
1O
1T
#8890000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#8900000000
1!
b0010 %
b1001111 &
1'
b0010 +
b1001111 ,
14
19
1>
1C
b0010 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#8910000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#8920000000
1!
1'
14
19
1>
1C
1O
1T
#8930000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#8940000000
1!
1'
14
19
1>
1C
1O
1T
#8950000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#8960000000
1!
1'
14
19
1>
1C
1O
1T
1W
#8970000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#8980000000
1!
1'
14
19
1>
1C
1O
1T
#8990000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#9000000000
1!
1'
14
19
1>
1C
1O
1T
#9010000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#9020000000
1!
b0100 %
b0000001 &
1'
b0100 +
b0000001 ,
14
19
1>
1C
b0100 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#9030000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#9040000000
1!
1'
14
19
1>
1C
1O
1T
#9050000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#9060000000
1!
1'
14
19
1>
1C
1O
1T
#9070000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#9080000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
1W
#9090000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#9100000000
1!
1'
14
19
1>
1C
1O
1T
#9110000000
0!
0#
0'
0)
04
09
0:
0>
0C
b100 K
0O
0T
b100 X
#9120000000
#9130000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
#9140000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#9150000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#9160000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#9170000000
1!
1'
14
19
1>
1C
1O
1T
#9180000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#9190000000
1!
1'
14
19
1>
1C
1O
1T
#9200000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#9210000000
1!
1'
14
19
1>
1C
1O
1T
1W
#9220000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#9230000000
1!
1'
14
19
1>
1C
1O
1T
#9240000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#9250000000
1!
1'
14
19
1>
1C
1O
1T
#9260000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#9270000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#9280000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#9290000000
1!
1'
14
19
1>
1C
1O
1T
#9300000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#9310000000
1!
1'
14
19
1>
1C
1O
1T
#9320000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#9330000000
1!
1'
14
19
1>
1C
1O
1T
1W
#9340000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#9350000000
1!
1'
14
19
1>
1C
1O
1T
#9360000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#9370000000
1!
1'
14
19
1>
1C
1O
1T
#9380000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#9390000000
1!
b0010 %
b1001111 &
1'
b0010 +
b1001111 ,
14
19
1>
1C
b0010 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#9400000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#9410000000
1!
1'
14
19
1>
1C
1O
1T
#9420000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#9430000000
1!
1'
14
19
1>
1C
1O
1T
#9440000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#9450000000
1!
1'
14
19
1>
1C
1O
1T
1W
#9460000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#9470000000
1!
1'
14
19
1>
1C
1O
1T
#9480000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#9490000000
1!
1'
14
19
1>
1C
1O
1T
#9500000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#9510000000
1!
b0100 %
b0000001 &
1'
b0100 +
b0000001 ,
14
19
1>
1C
b0100 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
#9520000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#9530000000
1!
1'
14
19
1>
1C
1O
1T
#9540000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#9550000000
1!
1'
14
19
1>
1C
1O
1T
#9560000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#9570000000
1!
1'
14
19
1>
1C
1O
1T
1W
#9580000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#9590000000
1!
1'
14
19
1>
1C
1O
1T
#9600000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#9610000000
1!
1'
14
19
1>
1C
1O
1T
#9620000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#9630000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1O
1T
0W
#9640000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#9650000000
1!
1#
1'
1)
1.
14
19
1:
1;
1<
1=
1>
1C
1O
1T
#9660000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#9670000000
1!
1'
14
19
1>
1C
1O
1T
#9680000000
0!
0#
0'
0)
04
09
0:
0>
0C
b10 K
0O
0T
b10 X
#9690000000
#9700000000
1!
1'
0.
14
19
0;
0<
0=
1>
1C
1O
1T
1W
#9710000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#9720000000
1!
1'
14
19
1>
1C
1O
1T
#9730000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#9740000000
1!
1'
14
19
1>
1C
1O
1T
#9750000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#9760000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1O
1T
0W
#9770000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#9780000000
1!
1'
14
19
1>
1C
1O
1T
#9790000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#9800000000
1!
1'
14
19
1>
1C
1O
1T
#9810000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#9820000000
1!
1'
14
19
1>
1C
1O
1T
1W
#9830000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#9840000000
1!
1'
14
19
1>
1C
1O
1T
#9850000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#9860000000
1!
1'
14
19
1>
1C
1O
1T
#9870000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#9880000000
1!
b0010 %
b1001111 &
1'
b0010 +
b1001111 ,
14
19
1>
1C
b0010 I
b1001111 J
b0001 N
1O
1T
0W
b1001111 Y
b0001 Z
#9890000000
0!
0'
04
09
0>
0C
b0 K
0O
0T
b0 X
#9900000000
1!
1'
14
19
1>
1C
1O
1T
#9910000000
0!
0'
04
09
0>
0C
b1 K
0O
0T
b1 X
#9920000000
1!
1'
14
19
1>
1C
1O
1T
#9930000000
0!
0'
04
09
0>
0C
b10 K
0O
0T
b10 X
#9940000000
1!
1'
14
19
1>
1C
1O
1T
1W
#9950000000
0!
0'
04
09
0>
0C
b11 K
0O
0T
b11 X
#9960000000
1!
1'
14
19
1>
1C
1O
1T
#9970000000
0!
0'
04
09
0>
0C
b100 K
0O
0T
b100 X
#9980000000
1!
1'
14
19
1>
1C
1O
1T
#9990000000
0!
0'
04
09
0>
0C
b101 K
0O
0T
b101 X
#10000000000
1!
b0100 %
b0000001 &
1'
b0100 +
b0000001 ,
14
19
1>
1C
b0100 I
b0000001 J
b0000 N
1O
1T
0W
b0000001 Y
b0000 Z
