$date
  Fri Apr 05 21:14:17 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp1_1 $end
$var reg 1 ! in1 $end
$var reg 1 " in2 $end
$var reg 1 # in3 $end
$var reg 1 $ salida $end
$scope module uut $end
$var reg 1 % z $end
$var reg 1 & a $end
$var reg 1 ' b $end
$var reg 1 ( c $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
U"
U#
0$
0%
0&
U'
U(
#10000000
0"
0'
#20000000
0#
0(
#30000000
1#
1(
#40000000
1"
1'
#50000000
0#
0(
#60000000
#70000000
1#
1(
#80000000
1!
1$
1%
1&
#90000000
0"
0'
#100000000
0#
0$
0%
0(
#110000000
1#
1$
1%
1(
#120000000
1"
1'
#130000000
0#
0(
#140000000
#150000000
1#
1(
#160000000
0!
0$
0%
0&
#170000000
0"
0'
#180000000
0#
0(
#190000000
1#
1(
#200000000
1"
1'
#210000000
0#
0(
#220000000
#230000000
1#
1(
#240000000
1!
1$
1%
1&
#250000000
0"
0'
#260000000
0#
0$
0%
0(
#270000000
1#
1$
1%
1(
#280000000
1"
1'
#290000000
0#
0(
#300000000
#310000000
1#
1(
#320000000
0!
0$
0%
0&
#330000000
0"
0'
#340000000
0#
0(
#350000000
1#
1(
#360000000
1"
1'
#370000000
0#
0(
#380000000
#390000000
1#
1(
#400000000
1!
1$
1%
1&
#410000000
0"
0'
#420000000
0#
0$
0%
0(
#430000000
1#
1$
1%
1(
#440000000
1"
1'
#450000000
0#
0(
#460000000
#470000000
1#
1(
#480000000
0!
0$
0%
0&
#490000000
0"
0'
#500000000
0#
0(
#510000000
1#
1(
#520000000
1"
1'
#530000000
0#
0(
#540000000
#550000000
1#
1(
#560000000
1!
1$
1%
1&
#570000000
0"
0'
#580000000
0#
0$
0%
0(
#590000000
1#
1$
1%
1(
#600000000
1"
1'
#610000000
0#
0(
#620000000
#630000000
1#
1(
#640000000
0!
0$
0%
0&
#650000000
0"
0'
#660000000
0#
0(
#670000000
1#
1(
#680000000
1"
1'
#690000000
0#
0(
#700000000
#710000000
1#
1(
#720000000
1!
1$
1%
1&
#730000000
0"
0'
#740000000
0#
0$
0%
0(
#750000000
1#
1$
1%
1(
#760000000
1"
1'
#770000000
0#
0(
#780000000
#790000000
1#
1(
#800000000
0!
0$
0%
0&
#810000000
0"
0'
#820000000
0#
0(
#830000000
1#
1(
#840000000
1"
1'
#850000000
0#
0(
#860000000
#870000000
1#
1(
#880000000
1!
1$
1%
1&
#890000000
0"
0'
#900000000
0#
0$
0%
0(
#910000000
1#
1$
1%
1(
#920000000
1"
1'
#930000000
0#
0(
#940000000
#950000000
1#
1(
#960000000
0!
0$
0%
0&
#970000000
0"
0'
#980000000
0#
0(
#990000000
1#
1(
#1000000000
1"
1'
#1010000000
0#
0(
#1020000000
#1030000000
1#
1(
#1040000000
1!
1$
1%
1&
#1050000000
0"
0'
#1060000000
0#
0$
0%
0(
#1070000000
1#
1$
1%
1(
#1080000000
1"
1'
#1090000000
0#
0(
#1100000000
#1110000000
1#
1(
#1120000000
0!
0$
0%
0&
#1130000000
0"
0'
#1140000000
0#
0(
#1150000000
1#
1(
#1160000000
1"
1'
#1170000000
0#
0(
#1180000000
#1190000000
1#
1(
#1200000000
1!
1$
1%
1&
#1210000000
0"
0'
#1220000000
0#
0$
0%
0(
#1230000000
1#
1$
1%
1(
#1240000000
1"
1'
#1250000000
0#
0(
#1260000000
#1270000000
1#
1(
#1280000000
0!
0$
0%
0&
#1290000000
0"
0'
#1300000000
0#
0(
#1310000000
1#
1(
#1320000000
1"
1'
#1330000000
0#
0(
#1340000000
#1350000000
1#
1(
#1360000000
1!
1$
1%
1&
#1370000000
0"
0'
#1380000000
0#
0$
0%
0(
#1390000000
1#
1$
1%
1(
#1400000000
1"
1'
#1410000000
0#
0(
#1420000000
#1430000000
1#
1(
#1440000000
0!
0$
0%
0&
#1450000000
0"
0'
#1460000000
0#
0(
#1470000000
1#
1(
#1480000000
1"
1'
#1490000000
0#
0(
#1500000000
#1510000000
1#
1(
#1520000000
1!
1$
1%
1&
#1530000000
0"
0'
#1540000000
0#
0$
0%
0(
#1550000000
1#
1$
1%
1(
#1560000000
1"
1'
#1570000000
0#
0(
#1580000000
#1590000000
1#
1(
#1600000000
0!
0$
0%
0&
#1610000000
0"
0'
#1620000000
0#
0(
#1630000000
1#
1(
#1640000000
1"
1'
#1650000000
0#
0(
#1660000000
#1670000000
1#
1(
#1680000000
1!
1$
1%
1&
#1690000000
0"
0'
#1700000000
0#
0$
0%
0(
#1710000000
1#
1$
1%
1(
#1720000000
1"
1'
#1730000000
0#
0(
#1740000000
#1750000000
1#
1(
#1760000000
0!
0$
0%
0&
#1770000000
0"
0'
#1780000000
0#
0(
#1790000000
1#
1(
#1800000000
1"
1'
#1810000000
0#
0(
#1820000000
#1830000000
1#
1(
#1840000000
1!
1$
1%
1&
#1850000000
0"
0'
#1860000000
0#
0$
0%
0(
#1870000000
1#
1$
1%
1(
#1880000000
1"
1'
#1890000000
0#
0(
#1900000000
#1910000000
1#
1(
#1920000000
0!
0$
0%
0&
#1930000000
0"
0'
#1940000000
0#
0(
#1950000000
1#
1(
#1960000000
1"
1'
#1970000000
0#
0(
#1980000000
#1990000000
1#
1(
#2000000000
1!
1$
1%
1&
#2010000000
0"
0'
#2020000000
0#
0$
0%
0(
#2030000000
1#
1$
1%
1(
#2040000000
1"
1'
#2050000000
0#
0(
#2060000000
#2070000000
1#
1(
#2080000000
0!
0$
0%
0&
#2090000000
0"
0'
#2100000000
0#
0(
#2110000000
1#
1(
#2120000000
1"
1'
#2130000000
0#
0(
#2140000000
#2150000000
1#
1(
#2160000000
1!
1$
1%
1&
#2170000000
0"
0'
#2180000000
0#
0$
0%
0(
#2190000000
1#
1$
1%
1(
#2200000000
1"
1'
#2210000000
0#
0(
#2220000000
#2230000000
1#
1(
#2240000000
0!
0$
0%
0&
#2250000000
0"
0'
#2260000000
0#
0(
#2270000000
1#
1(
#2280000000
1"
1'
#2290000000
0#
0(
#2300000000
#2310000000
1#
1(
#2320000000
1!
1$
1%
1&
#2330000000
0"
0'
#2340000000
0#
0$
0%
0(
#2350000000
1#
1$
1%
1(
#2360000000
1"
1'
#2370000000
0#
0(
#2380000000
#2390000000
1#
1(
#2400000000
0!
0$
0%
0&
#2410000000
0"
0'
#2420000000
0#
0(
#2430000000
1#
1(
#2440000000
1"
1'
#2450000000
0#
0(
#2460000000
#2470000000
1#
1(
#2480000000
1!
1$
1%
1&
#2490000000
0"
0'
#2500000000
0#
0$
0%
0(
#2510000000
1#
1$
1%
1(
#2520000000
1"
1'
#2530000000
0#
0(
#2540000000
#2550000000
1#
1(
#2560000000
0!
0$
0%
0&
#2570000000
0"
0'
#2580000000
0#
0(
#2590000000
1#
1(
#2600000000
1"
1'
#2610000000
0#
0(
#2620000000
#2630000000
1#
1(
#2640000000
1!
1$
1%
1&
#2650000000
0"
0'
#2660000000
0#
0$
0%
0(
#2670000000
1#
1$
1%
1(
#2680000000
1"
1'
#2690000000
0#
0(
#2700000000
#2710000000
1#
1(
#2720000000
0!
0$
0%
0&
#2730000000
0"
0'
#2740000000
0#
0(
#2750000000
1#
1(
#2760000000
1"
1'
#2770000000
0#
0(
#2780000000
#2790000000
1#
1(
#2800000000
1!
1$
1%
1&
#2810000000
0"
0'
#2820000000
0#
0$
0%
0(
#2830000000
1#
1$
1%
1(
#2840000000
1"
1'
#2850000000
0#
0(
#2860000000
#2870000000
1#
1(
#2880000000
0!
0$
0%
0&
#2890000000
0"
0'
#2900000000
0#
0(
#2910000000
1#
1(
#2920000000
1"
1'
#2930000000
0#
0(
#2940000000
#2950000000
1#
1(
#2960000000
1!
1$
1%
1&
#2970000000
0"
0'
#2980000000
0#
0$
0%
0(
#2990000000
1#
1$
1%
1(
#3000000000
1"
1'
#3010000000
0#
0(
#3020000000
#3030000000
1#
1(
#3040000000
0!
0$
0%
0&
#3050000000
0"
0'
#3060000000
0#
0(
#3070000000
1#
1(
#3080000000
1"
1'
#3090000000
0#
0(
#3100000000
#3110000000
1#
1(
#3120000000
1!
1$
1%
1&
#3130000000
0"
0'
#3140000000
0#
0$
0%
0(
#3150000000
1#
1$
1%
1(
#3160000000
1"
1'
#3170000000
0#
0(
#3180000000
#3190000000
1#
1(
#3200000000
0!
0$
0%
0&
#3210000000
0"
0'
#3220000000
0#
0(
#3230000000
1#
1(
#3240000000
1"
1'
#3250000000
0#
0(
#3260000000
#3270000000
1#
1(
#3280000000
1!
1$
1%
1&
#3290000000
0"
0'
#3300000000
0#
0$
0%
0(
#3310000000
1#
1$
1%
1(
#3320000000
1"
1'
#3330000000
0#
0(
#3340000000
#3350000000
1#
1(
#3360000000
0!
0$
0%
0&
#3370000000
0"
0'
#3380000000
0#
0(
#3390000000
1#
1(
#3400000000
1"
1'
#3410000000
0#
0(
#3420000000
#3430000000
1#
1(
#3440000000
1!
1$
1%
1&
#3450000000
0"
0'
#3460000000
0#
0$
0%
0(
#3470000000
1#
1$
1%
1(
#3480000000
1"
1'
#3490000000
0#
0(
#3500000000
#3510000000
1#
1(
#3520000000
0!
0$
0%
0&
#3530000000
0"
0'
#3540000000
0#
0(
#3550000000
1#
1(
#3560000000
1"
1'
#3570000000
0#
0(
#3580000000
#3590000000
1#
1(
#3600000000
1!
1$
1%
1&
#3610000000
0"
0'
#3620000000
0#
0$
0%
0(
#3630000000
1#
1$
1%
1(
#3640000000
1"
1'
#3650000000
0#
0(
#3660000000
#3670000000
1#
1(
#3680000000
0!
0$
0%
0&
#3690000000
0"
0'
#3700000000
0#
0(
#3710000000
1#
1(
#3720000000
1"
1'
#3730000000
0#
0(
#3740000000
#3750000000
1#
1(
#3760000000
1!
1$
1%
1&
#3770000000
0"
0'
#3780000000
0#
0$
0%
0(
#3790000000
1#
1$
1%
1(
#3800000000
1"
1'
#3810000000
0#
0(
#3820000000
#3830000000
1#
1(
#3840000000
0!
0$
0%
0&
#3850000000
0"
0'
#3860000000
0#
0(
#3870000000
1#
1(
#3880000000
1"
1'
#3890000000
0#
0(
#3900000000
#3910000000
1#
1(
#3920000000
1!
1$
1%
1&
#3930000000
0"
0'
#3940000000
0#
0$
0%
0(
#3950000000
1#
1$
1%
1(
#3960000000
1"
1'
#3970000000
0#
0(
#3980000000
#3990000000
1#
1(
#4000000000
0!
0$
0%
0&
#4010000000
0"
0'
#4020000000
0#
0(
#4030000000
1#
1(
#4040000000
1"
1'
#4050000000
0#
0(
#4060000000
#4070000000
1#
1(
#4080000000
1!
1$
1%
1&
#4090000000
0"
0'
#4100000000
0#
0$
0%
0(
#4110000000
1#
1$
1%
1(
#4120000000
1"
1'
#4130000000
0#
0(
#4140000000
#4150000000
1#
1(
#4160000000
0!
0$
0%
0&
#4170000000
0"
0'
#4180000000
0#
0(
#4190000000
1#
1(
#4200000000
1"
1'
#4210000000
0#
0(
#4220000000
#4230000000
1#
1(
#4240000000
1!
1$
1%
1&
#4250000000
0"
0'
#4260000000
0#
0$
0%
0(
#4270000000
1#
1$
1%
1(
#4280000000
1"
1'
#4290000000
0#
0(
#4300000000
#4310000000
1#
1(
#4320000000
0!
0$
0%
0&
#4330000000
0"
0'
#4340000000
0#
0(
#4350000000
1#
1(
#4360000000
1"
1'
#4370000000
0#
0(
#4380000000
#4390000000
1#
1(
#4400000000
1!
1$
1%
1&
#4410000000
0"
0'
#4420000000
0#
0$
0%
0(
#4430000000
1#
1$
1%
1(
#4440000000
1"
1'
#4450000000
0#
0(
#4460000000
#4470000000
1#
1(
#4480000000
0!
0$
0%
0&
#4490000000
0"
0'
#4500000000
0#
0(
#4510000000
1#
1(
#4520000000
1"
1'
#4530000000
0#
0(
#4540000000
#4550000000
1#
1(
#4560000000
1!
1$
1%
1&
#4570000000
0"
0'
#4580000000
0#
0$
0%
0(
#4590000000
1#
1$
1%
1(
#4600000000
1"
1'
#4610000000
0#
0(
#4620000000
#4630000000
1#
1(
#4640000000
0!
0$
0%
0&
#4650000000
0"
0'
#4660000000
0#
0(
#4670000000
1#
1(
#4680000000
1"
1'
#4690000000
0#
0(
#4700000000
#4710000000
1#
1(
#4720000000
1!
1$
1%
1&
#4730000000
0"
0'
#4740000000
0#
0$
0%
0(
#4750000000
1#
1$
1%
1(
#4760000000
1"
1'
#4770000000
0#
0(
#4780000000
#4790000000
1#
1(
#4800000000
0!
0$
0%
0&
#4810000000
0"
0'
#4820000000
0#
0(
#4830000000
1#
1(
#4840000000
1"
1'
#4850000000
0#
0(
#4860000000
#4870000000
1#
1(
#4880000000
1!
1$
1%
1&
#4890000000
0"
0'
#4900000000
0#
0$
0%
0(
#4910000000
1#
1$
1%
1(
#4920000000
1"
1'
#4930000000
0#
0(
#4940000000
#4950000000
1#
1(
#4960000000
0!
0$
0%
0&
#4970000000
0"
0'
#4980000000
0#
0(
#4990000000
1#
1(
#5000000000
1"
1'
#5010000000
0#
0(
#5020000000
#5030000000
1#
1(
#5040000000
1!
1$
1%
1&
#5050000000
0"
0'
#5060000000
0#
0$
0%
0(
#5070000000
1#
1$
1%
1(
#5080000000
1"
1'
#5090000000
0#
0(
#5100000000
#5110000000
1#
1(
#5120000000
0!
0$
0%
0&
#5130000000
0"
0'
#5140000000
0#
0(
#5150000000
1#
1(
#5160000000
1"
1'
#5170000000
0#
0(
#5180000000
#5190000000
1#
1(
#5200000000
1!
1$
1%
1&
#5210000000
0"
0'
#5220000000
0#
0$
0%
0(
#5230000000
1#
1$
1%
1(
#5240000000
1"
1'
#5250000000
0#
0(
#5260000000
#5270000000
1#
1(
#5280000000
0!
0$
0%
0&
#5290000000
0"
0'
#5300000000
0#
0(
#5310000000
1#
1(
#5320000000
1"
1'
#5330000000
0#
0(
#5340000000
#5350000000
1#
1(
#5360000000
1!
1$
1%
1&
#5370000000
0"
0'
#5380000000
0#
0$
0%
0(
#5390000000
1#
1$
1%
1(
#5400000000
1"
1'
#5410000000
0#
0(
#5420000000
#5430000000
1#
1(
#5440000000
0!
0$
0%
0&
#5450000000
0"
0'
#5460000000
0#
0(
#5470000000
1#
1(
#5480000000
1"
1'
#5490000000
0#
0(
#5500000000
#5510000000
1#
1(
#5520000000
1!
1$
1%
1&
#5530000000
0"
0'
#5540000000
0#
0$
0%
0(
#5550000000
1#
1$
1%
1(
#5560000000
1"
1'
#5570000000
0#
0(
#5580000000
#5590000000
1#
1(
#5600000000
0!
0$
0%
0&
#5610000000
0"
0'
#5620000000
0#
0(
#5630000000
1#
1(
#5640000000
1"
1'
#5650000000
0#
0(
#5660000000
#5670000000
1#
1(
#5680000000
1!
1$
1%
1&
#5690000000
0"
0'
#5700000000
0#
0$
0%
0(
#5710000000
1#
1$
1%
1(
#5720000000
1"
1'
#5730000000
0#
0(
#5740000000
#5750000000
1#
1(
#5760000000
0!
0$
0%
0&
#5770000000
0"
0'
#5780000000
0#
0(
#5790000000
1#
1(
#5800000000
1"
1'
#5810000000
0#
0(
#5820000000
#5830000000
1#
1(
#5840000000
1!
1$
1%
1&
#5850000000
0"
0'
#5860000000
0#
0$
0%
0(
#5870000000
1#
1$
1%
1(
#5880000000
1"
1'
#5890000000
0#
0(
#5900000000
#5910000000
1#
1(
#5920000000
0!
0$
0%
0&
#5930000000
0"
0'
#5940000000
0#
0(
#5950000000
1#
1(
#5960000000
1"
1'
#5970000000
0#
0(
#5980000000
#5990000000
1#
1(
#6000000000
1!
1$
1%
1&
#6010000000
0"
0'
#6020000000
0#
0$
0%
0(
#6030000000
1#
1$
1%
1(
#6040000000
1"
1'
#6050000000
0#
0(
#6060000000
#6070000000
1#
1(
#6080000000
0!
0$
0%
0&
#6090000000
0"
0'
#6100000000
0#
0(
#6110000000
1#
1(
#6120000000
1"
1'
#6130000000
0#
0(
#6140000000
#6150000000
1#
1(
#6160000000
1!
1$
1%
1&
#6170000000
0"
0'
#6180000000
0#
0$
0%
0(
#6190000000
1#
1$
1%
1(
#6200000000
1"
1'
#6210000000
0#
0(
#6220000000
#6230000000
1#
1(
#6240000000
0!
0$
0%
0&
#6250000000
0"
0'
#6260000000
0#
0(
#6270000000
1#
1(
#6280000000
1"
1'
#6290000000
0#
0(
#6300000000
#6310000000
1#
1(
#6320000000
1!
1$
1%
1&
#6330000000
0"
0'
#6340000000
0#
0$
0%
0(
#6350000000
1#
1$
1%
1(
#6360000000
1"
1'
#6370000000
0#
0(
#6380000000
#6390000000
1#
1(
#6400000000
0!
0$
0%
0&
#6410000000
0"
0'
#6420000000
0#
0(
#6430000000
1#
1(
#6440000000
1"
1'
#6450000000
0#
0(
#6460000000
#6470000000
1#
1(
#6480000000
1!
1$
1%
1&
#6490000000
0"
0'
#6500000000
0#
0$
0%
0(
#6510000000
1#
1$
1%
1(
#6520000000
1"
1'
#6530000000
0#
0(
#6540000000
#6550000000
1#
1(
#6560000000
0!
0$
0%
0&
#6570000000
0"
0'
#6580000000
0#
0(
#6590000000
1#
1(
#6600000000
1"
1'
#6610000000
0#
0(
#6620000000
#6630000000
1#
1(
#6640000000
1!
1$
1%
1&
#6650000000
0"
0'
#6660000000
0#
0$
0%
0(
#6670000000
1#
1$
1%
1(
#6680000000
1"
1'
#6690000000
0#
0(
#6700000000
#6710000000
1#
1(
#6720000000
0!
0$
0%
0&
#6730000000
0"
0'
#6740000000
0#
0(
#6750000000
1#
1(
#6760000000
1"
1'
#6770000000
0#
0(
#6780000000
#6790000000
1#
1(
#6800000000
1!
1$
1%
1&
#6810000000
0"
0'
#6820000000
0#
0$
0%
0(
#6830000000
1#
1$
1%
1(
#6840000000
1"
1'
#6850000000
0#
0(
#6860000000
#6870000000
1#
1(
#6880000000
0!
0$
0%
0&
#6890000000
0"
0'
#6900000000
0#
0(
#6910000000
1#
1(
#6920000000
1"
1'
#6930000000
0#
0(
#6940000000
#6950000000
1#
1(
#6960000000
1!
1$
1%
1&
#6970000000
0"
0'
#6980000000
0#
0$
0%
0(
#6990000000
1#
1$
1%
1(
#7000000000
1"
1'
#7010000000
0#
0(
#7020000000
#7030000000
1#
1(
#7040000000
0!
0$
0%
0&
#7050000000
0"
0'
#7060000000
0#
0(
#7070000000
1#
1(
#7080000000
1"
1'
#7090000000
0#
0(
#7100000000
#7110000000
1#
1(
#7120000000
1!
1$
1%
1&
#7130000000
0"
0'
#7140000000
0#
0$
0%
0(
#7150000000
1#
1$
1%
1(
#7160000000
1"
1'
#7170000000
0#
0(
#7180000000
#7190000000
1#
1(
#7200000000
0!
0$
0%
0&
#7210000000
0"
0'
#7220000000
0#
0(
#7230000000
1#
1(
#7240000000
1"
1'
#7250000000
0#
0(
#7260000000
#7270000000
1#
1(
#7280000000
1!
1$
1%
1&
#7290000000
0"
0'
#7300000000
0#
0$
0%
0(
#7310000000
1#
1$
1%
1(
#7320000000
1"
1'
#7330000000
0#
0(
#7340000000
#7350000000
1#
1(
#7360000000
0!
0$
0%
0&
#7370000000
0"
0'
#7380000000
0#
0(
#7390000000
1#
1(
#7400000000
1"
1'
#7410000000
0#
0(
#7420000000
#7430000000
1#
1(
#7440000000
1!
1$
1%
1&
#7450000000
0"
0'
#7460000000
0#
0$
0%
0(
#7470000000
1#
1$
1%
1(
#7480000000
1"
1'
#7490000000
0#
0(
#7500000000
#7510000000
1#
1(
#7520000000
0!
0$
0%
0&
#7530000000
0"
0'
#7540000000
0#
0(
#7550000000
1#
1(
#7560000000
1"
1'
#7570000000
0#
0(
#7580000000
#7590000000
1#
1(
#7600000000
1!
1$
1%
1&
#7610000000
0"
0'
#7620000000
0#
0$
0%
0(
#7630000000
1#
1$
1%
1(
#7640000000
1"
1'
#7650000000
0#
0(
#7660000000
#7670000000
1#
1(
#7680000000
0!
0$
0%
0&
#7690000000
0"
0'
#7700000000
0#
0(
#7710000000
1#
1(
#7720000000
1"
1'
#7730000000
0#
0(
#7740000000
#7750000000
1#
1(
#7760000000
1!
1$
1%
1&
#7770000000
0"
0'
#7780000000
0#
0$
0%
0(
#7790000000
1#
1$
1%
1(
#7800000000
1"
1'
#7810000000
0#
0(
#7820000000
#7830000000
1#
1(
#7840000000
0!
0$
0%
0&
#7850000000
0"
0'
#7860000000
0#
0(
#7870000000
1#
1(
#7880000000
1"
1'
#7890000000
0#
0(
#7900000000
#7910000000
1#
1(
#7920000000
1!
1$
1%
1&
#7930000000
0"
0'
#7940000000
0#
0$
0%
0(
#7950000000
1#
1$
1%
1(
#7960000000
1"
1'
#7970000000
0#
0(
#7980000000
#7990000000
1#
1(
#8000000000
0!
0$
0%
0&
#8010000000
0"
0'
#8020000000
0#
0(
#8030000000
1#
1(
#8040000000
1"
1'
#8050000000
0#
0(
#8060000000
#8070000000
1#
1(
#8080000000
1!
1$
1%
1&
#8090000000
0"
0'
#8100000000
0#
0$
0%
0(
#8110000000
1#
1$
1%
1(
#8120000000
1"
1'
#8130000000
0#
0(
#8140000000
#8150000000
1#
1(
#8160000000
0!
0$
0%
0&
#8170000000
0"
0'
#8180000000
0#
0(
#8190000000
1#
1(
#8200000000
1"
1'
#8210000000
0#
0(
#8220000000
#8230000000
1#
1(
#8240000000
1!
1$
1%
1&
#8250000000
0"
0'
#8260000000
0#
0$
0%
0(
#8270000000
1#
1$
1%
1(
#8280000000
1"
1'
#8290000000
0#
0(
#8300000000
#8310000000
1#
1(
#8320000000
0!
0$
0%
0&
#8330000000
0"
0'
#8340000000
0#
0(
#8350000000
1#
1(
#8360000000
1"
1'
#8370000000
0#
0(
#8380000000
#8390000000
1#
1(
#8400000000
1!
1$
1%
1&
#8410000000
0"
0'
#8420000000
0#
0$
0%
0(
#8430000000
1#
1$
1%
1(
#8440000000
1"
1'
#8450000000
0#
0(
#8460000000
#8470000000
1#
1(
#8480000000
0!
0$
0%
0&
#8490000000
0"
0'
#8500000000
0#
0(
#8510000000
1#
1(
#8520000000
1"
1'
#8530000000
0#
0(
#8540000000
#8550000000
1#
1(
#8560000000
1!
1$
1%
1&
#8570000000
0"
0'
#8580000000
0#
0$
0%
0(
#8590000000
1#
1$
1%
1(
#8600000000
1"
1'
#8610000000
0#
0(
#8620000000
#8630000000
1#
1(
#8640000000
0!
0$
0%
0&
#8650000000
0"
0'
#8660000000
0#
0(
#8670000000
1#
1(
#8680000000
1"
1'
#8690000000
0#
0(
#8700000000
#8710000000
1#
1(
#8720000000
1!
1$
1%
1&
#8730000000
0"
0'
#8740000000
0#
0$
0%
0(
#8750000000
1#
1$
1%
1(
#8760000000
1"
1'
#8770000000
0#
0(
#8780000000
#8790000000
1#
1(
#8800000000
0!
0$
0%
0&
#8810000000
0"
0'
#8820000000
0#
0(
#8830000000
1#
1(
#8840000000
1"
1'
#8850000000
0#
0(
#8860000000
#8870000000
1#
1(
#8880000000
1!
1$
1%
1&
#8890000000
0"
0'
#8900000000
0#
0$
0%
0(
#8910000000
1#
1$
1%
1(
#8920000000
1"
1'
#8930000000
0#
0(
#8940000000
#8950000000
1#
1(
#8960000000
0!
0$
0%
0&
#8970000000
0"
0'
#8980000000
0#
0(
#8990000000
1#
1(
#9000000000
1"
1'
#9010000000
0#
0(
#9020000000
#9030000000
1#
1(
#9040000000
1!
1$
1%
1&
#9050000000
0"
0'
#9060000000
0#
0$
0%
0(
#9070000000
1#
1$
1%
1(
#9080000000
1"
1'
#9090000000
0#
0(
#9100000000
#9110000000
1#
1(
#9120000000
0!
0$
0%
0&
#9130000000
0"
0'
#9140000000
0#
0(
#9150000000
1#
1(
#9160000000
1"
1'
#9170000000
0#
0(
#9180000000
#9190000000
1#
1(
#9200000000
1!
1$
1%
1&
#9210000000
0"
0'
#9220000000
0#
0$
0%
0(
#9230000000
1#
1$
1%
1(
#9240000000
1"
1'
#9250000000
0#
0(
#9260000000
#9270000000
1#
1(
#9280000000
0!
0$
0%
0&
#9290000000
0"
0'
#9300000000
0#
0(
#9310000000
1#
1(
#9320000000
1"
1'
#9330000000
0#
0(
#9340000000
#9350000000
1#
1(
#9360000000
1!
1$
1%
1&
#9370000000
0"
0'
#9380000000
0#
0$
0%
0(
#9390000000
1#
1$
1%
1(
#9400000000
1"
1'
#9410000000
0#
0(
#9420000000
#9430000000
1#
1(
#9440000000
0!
0$
0%
0&
#9450000000
0"
0'
#9460000000
0#
0(
#9470000000
1#
1(
#9480000000
1"
1'
#9490000000
0#
0(
#9500000000
#9510000000
1#
1(
#9520000000
1!
1$
1%
1&
#9530000000
0"
0'
#9540000000
0#
0$
0%
0(
#9550000000
1#
1$
1%
1(
#9560000000
1"
1'
#9570000000
0#
0(
#9580000000
#9590000000
1#
1(
#9600000000
0!
0$
0%
0&
#9610000000
0"
0'
#9620000000
0#
0(
#9630000000
1#
1(
#9640000000
1"
1'
#9650000000
0#
0(
#9660000000
#9670000000
1#
1(
#9680000000
1!
1$
1%
1&
#9690000000
0"
0'
#9700000000
0#
0$
0%
0(
#9710000000
1#
1$
1%
1(
#9720000000
1"
1'
#9730000000
0#
0(
#9740000000
#9750000000
1#
1(
#9760000000
0!
0$
0%
0&
#9770000000
0"
0'
#9780000000
0#
0(
#9790000000
1#
1(
#9800000000
1"
1'
#9810000000
0#
0(
#9820000000
#9830000000
1#
1(
#9840000000
1!
1$
1%
1&
#9850000000
0"
0'
#9860000000
0#
0$
0%
0(
#9870000000
1#
1$
1%
1(
#9880000000
1"
1'
#9890000000
0#
0(
#9900000000
#9910000000
1#
1(
#9920000000
0!
0$
0%
0&
#9930000000
0"
0'
#9940000000
0#
0(
#9950000000
1#
1(
#9960000000
1"
1'
#9970000000
0#
0(
#9980000000
#9990000000
1#
1(
#10000000000
1!
1$
1%
1&
