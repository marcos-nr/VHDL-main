$date
  Tue Apr 30 10:55:26 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp2_2 $end
$var reg 1 ! clk $end
$var reg 1 " start $end
$var reg 1 # reset $end
$var reg 1 $ led_uv $end
$var reg 1 % led_rojo $end
$var reg 1 & led_conta $end
$var reg 7 ' segmentos[6:0] $end
$var integer 32 ( min_count $end
$var integer 32 ) max_count $end
$scope module uut $end
$var reg 1 * clk $end
$var reg 1 + start $end
$var reg 1 , reset $end
$var reg 1 - led_uv $end
$var reg 1 . led_rojo $end
$var reg 1 / led_conta $end
$var reg 7 0 segmentos[6:0] $end
$var reg 1 1 debounced_start $end
$var reg 1 2 debounced_recet $end
$var reg 1 3 enable_conta $end
$var reg 1 4 reset_conta $end
$var reg 4 5 bcd[3:0] $end
$var integer 32 6 cuenta $end
$var reg 1 7 enable_display $end
$var integer 32 8 segundos $end
$scope module a $end
$var reg 1 9 clk $end
$var reg 1 : key $end
$var reg 1 ; debounced_key $end
$var reg 1 < key_stable $end
$var reg 1 = last_key $end
$upscope $end
$scope module b $end
$var reg 1 > clk $end
$var reg 1 ? key $end
$var reg 1 @ debounced_key $end
$var reg 1 A key_stable $end
$var reg 1 B last_key $end
$upscope $end
$scope module c $end
$var reg 1 C clk $end
$var reg 1 D reset $end
$var reg 1 E enable $end
$var reg 1 F cout $end
$var integer 32 G q $end
$upscope $end
$scope module d $end
$var reg 7 H segmentos[6:0] $end
$var reg 4 I bcd[3:0] $end
$var reg 1 J enable $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
0#
0$
0%
U&
b1111110 '
b0 (
b0 )
0*
0+
0,
0-
0.
U/
b1111110 0
U1
U2
U3
U4
b0000 5
b0 6
17
b0 8
09
0:
U;
U<
U=
0>
0?
U@
UA
UB
0C
UD
UE
UF
b0 G
b1111110 H
b0000 I
1J
#10000000
1!
U$
U%
0&
1*
U-
U.
0/
01
02
19
0;
0<
0=
1>
0@
0A
0B
1C
0F
#20000000
0!
0*
09
0>
0C
#30000000
1!
1*
19
1>
1C
#40000000
0!
1"
0*
1+
09
1:
0>
0C
#50000000
1!
1*
11
19
1;
1<
1=
1>
1C
#60000000
0!
0*
09
0>
0C
#70000000
1!
1*
13
04
19
1>
1C
0D
1E
#80000000
0!
0*
09
0>
0C
#90000000
1!
0"
1$
0%
1*
0+
1-
0.
01
b1 6
19
0:
0;
0<
0=
1>
1C
b1 G
#100000000
0!
0*
09
0>
0C
#110000000
1!
1#
1*
1,
12
b10 6
19
1>
1?
1@
1A
1B
1C
b10 G
#120000000
0!
0*
09
0>
0C
#130000000
1!
1*
03
14
b11 6
19
1>
1C
1D
0E
b11 G
#140000000
0!
0*
09
0>
0C
#150000000
1!
0$
1%
1*
0-
1.
b0 6
19
1>
1C
b0 G
#160000000
0!
0#
0*
0,
09
0>
0?
0C
#170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#180000000
0!
0*
09
0>
0C
#190000000
1!
1*
19
1>
1C
#200000000
0!
0*
09
0>
0C
#210000000
1!
1*
19
1>
1C
#220000000
0!
0*
09
0>
0C
#230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#240000000
0!
0*
09
0>
0C
#250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#260000000
0!
0*
09
0>
0C
#270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#280000000
0!
0*
09
0>
0C
#290000000
1!
1*
b10 6
19
1>
1C
b10 G
#300000000
0!
0*
09
0>
0C
#310000000
1!
1*
b11 6
19
1>
1C
b11 G
#320000000
0!
0*
09
0>
0C
#330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#340000000
0!
0*
09
0>
0C
#350000000
1!
1*
b101 6
19
1>
1C
b101 G
#360000000
0!
0*
09
0>
0C
#370000000
1!
1*
b110 6
19
1>
1C
b110 G
#380000000
0!
0*
09
0>
0C
#390000000
1!
1*
b111 6
19
1>
1C
b111 G
#400000000
0!
0*
09
0>
0C
#410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#420000000
0!
0*
09
0>
0C
#430000000
1!
1*
b1 6
19
1>
1C
b1 G
#440000000
0!
0*
09
0>
0C
#450000000
1!
1*
b10 6
19
1>
1C
b10 G
#460000000
0!
0*
09
0>
0C
#470000000
1!
1*
b11 6
19
1>
1C
b11 G
#480000000
0!
0*
09
0>
0C
#490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#500000000
0!
0*
09
0>
0C
#510000000
1!
1*
b101 6
19
1>
1C
b101 G
#520000000
0!
0*
09
0>
0C
#530000000
1!
1*
b110 6
19
1>
1C
b110 G
#540000000
0!
0*
09
0>
0C
#550000000
1!
1*
b111 6
19
1>
1C
b111 G
#560000000
0!
0*
09
0>
0C
#570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#580000000
0!
0*
09
0>
0C
#590000000
1!
1*
b1 6
19
1>
1C
b1 G
#600000000
0!
0*
09
0>
0C
#610000000
1!
1*
b10 6
19
1>
1C
b10 G
#620000000
0!
0*
09
0>
0C
#630000000
1!
1*
b11 6
19
1>
1C
b11 G
#640000000
0!
0*
09
0>
0C
#650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#660000000
0!
0*
09
0>
0C
#670000000
1!
1*
b101 6
19
1>
1C
b101 G
#680000000
0!
0*
09
0>
0C
#690000000
1!
1*
b110 6
19
1>
1C
b110 G
#700000000
0!
0*
09
0>
0C
#710000000
1!
1*
b111 6
19
1>
1C
b111 G
#720000000
0!
1"
0*
1+
09
1:
0>
0C
#730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#740000000
0!
0*
09
0>
0C
#750000000
1!
1*
b1 6
19
1>
1C
b1 G
#760000000
0!
0*
09
0>
0C
#770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#780000000
0!
0*
09
0>
0C
#790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#800000000
0!
0*
09
0>
0C
#810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#820000000
0!
0*
09
0>
0C
#830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#840000000
0!
0#
0*
0,
09
0>
0?
0C
#850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#860000000
0!
0*
09
0>
0C
#870000000
1!
1*
19
1>
1C
#880000000
0!
0*
09
0>
0C
#890000000
1!
1*
19
1>
1C
#900000000
0!
0*
09
0>
0C
#910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#920000000
0!
0*
09
0>
0C
#930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#940000000
0!
0*
09
0>
0C
#950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#960000000
0!
0*
09
0>
0C
#970000000
1!
1*
b10 6
19
1>
1C
b10 G
#980000000
0!
0*
09
0>
0C
#990000000
1!
1*
b11 6
19
1>
1C
b11 G
#1000000000
0!
0*
09
0>
0C
#1010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1020000000
0!
0*
09
0>
0C
#1030000000
1!
1*
b101 6
19
1>
1C
b101 G
#1040000000
0!
0*
09
0>
0C
#1050000000
1!
1*
b110 6
19
1>
1C
b110 G
#1060000000
0!
0*
09
0>
0C
#1070000000
1!
1*
b111 6
19
1>
1C
b111 G
#1080000000
0!
0*
09
0>
0C
#1090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#1100000000
0!
0*
09
0>
0C
#1110000000
1!
1*
b1 6
19
1>
1C
b1 G
#1120000000
0!
0*
09
0>
0C
#1130000000
1!
1*
b10 6
19
1>
1C
b10 G
#1140000000
0!
0*
09
0>
0C
#1150000000
1!
1*
b11 6
19
1>
1C
b11 G
#1160000000
0!
0*
09
0>
0C
#1170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1180000000
0!
0*
09
0>
0C
#1190000000
1!
1*
b101 6
19
1>
1C
b101 G
#1200000000
0!
0*
09
0>
0C
#1210000000
1!
1*
b110 6
19
1>
1C
b110 G
#1220000000
0!
0*
09
0>
0C
#1230000000
1!
1*
b111 6
19
1>
1C
b111 G
#1240000000
0!
0*
09
0>
0C
#1250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#1260000000
0!
0*
09
0>
0C
#1270000000
1!
1*
b1 6
19
1>
1C
b1 G
#1280000000
0!
0*
09
0>
0C
#1290000000
1!
1*
b10 6
19
1>
1C
b10 G
#1300000000
0!
0*
09
0>
0C
#1310000000
1!
1*
b11 6
19
1>
1C
b11 G
#1320000000
0!
0*
09
0>
0C
#1330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1340000000
0!
0*
09
0>
0C
#1350000000
1!
1*
b101 6
19
1>
1C
b101 G
#1360000000
0!
0*
09
0>
0C
#1370000000
1!
1*
b110 6
19
1>
1C
b110 G
#1380000000
0!
0*
09
0>
0C
#1390000000
1!
1*
b111 6
19
1>
1C
b111 G
#1400000000
0!
1"
0*
1+
09
1:
0>
0C
#1410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#1420000000
0!
0*
09
0>
0C
#1430000000
1!
1*
b1 6
19
1>
1C
b1 G
#1440000000
0!
0*
09
0>
0C
#1450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#1460000000
0!
0*
09
0>
0C
#1470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#1480000000
0!
0*
09
0>
0C
#1490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#1500000000
0!
0*
09
0>
0C
#1510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#1520000000
0!
0#
0*
0,
09
0>
0?
0C
#1530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#1540000000
0!
0*
09
0>
0C
#1550000000
1!
1*
19
1>
1C
#1560000000
0!
0*
09
0>
0C
#1570000000
1!
1*
19
1>
1C
#1580000000
0!
0*
09
0>
0C
#1590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#1600000000
0!
0*
09
0>
0C
#1610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#1620000000
0!
0*
09
0>
0C
#1630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#1640000000
0!
0*
09
0>
0C
#1650000000
1!
1*
b10 6
19
1>
1C
b10 G
#1660000000
0!
0*
09
0>
0C
#1670000000
1!
1*
b11 6
19
1>
1C
b11 G
#1680000000
0!
0*
09
0>
0C
#1690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1700000000
0!
0*
09
0>
0C
#1710000000
1!
1*
b101 6
19
1>
1C
b101 G
#1720000000
0!
0*
09
0>
0C
#1730000000
1!
1*
b110 6
19
1>
1C
b110 G
#1740000000
0!
0*
09
0>
0C
#1750000000
1!
1*
b111 6
19
1>
1C
b111 G
#1760000000
0!
0*
09
0>
0C
#1770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#1780000000
0!
0*
09
0>
0C
#1790000000
1!
1*
b1 6
19
1>
1C
b1 G
#1800000000
0!
0*
09
0>
0C
#1810000000
1!
1*
b10 6
19
1>
1C
b10 G
#1820000000
0!
0*
09
0>
0C
#1830000000
1!
1*
b11 6
19
1>
1C
b11 G
#1840000000
0!
0*
09
0>
0C
#1850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1860000000
0!
0*
09
0>
0C
#1870000000
1!
1*
b101 6
19
1>
1C
b101 G
#1880000000
0!
0*
09
0>
0C
#1890000000
1!
1*
b110 6
19
1>
1C
b110 G
#1900000000
0!
0*
09
0>
0C
#1910000000
1!
1*
b111 6
19
1>
1C
b111 G
#1920000000
0!
0*
09
0>
0C
#1930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#1940000000
0!
0*
09
0>
0C
#1950000000
1!
1*
b1 6
19
1>
1C
b1 G
#1960000000
0!
0*
09
0>
0C
#1970000000
1!
1*
b10 6
19
1>
1C
b10 G
#1980000000
0!
0*
09
0>
0C
#1990000000
1!
1*
b11 6
19
1>
1C
b11 G
#2000000000
0!
0*
09
0>
0C
#2010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2020000000
0!
0*
09
0>
0C
#2030000000
1!
1*
b101 6
19
1>
1C
b101 G
#2040000000
0!
0*
09
0>
0C
#2050000000
1!
1*
b110 6
19
1>
1C
b110 G
#2060000000
0!
0*
09
0>
0C
#2070000000
1!
1*
b111 6
19
1>
1C
b111 G
#2080000000
0!
1"
0*
1+
09
1:
0>
0C
#2090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#2100000000
0!
0*
09
0>
0C
#2110000000
1!
1*
b1 6
19
1>
1C
b1 G
#2120000000
0!
0*
09
0>
0C
#2130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#2140000000
0!
0*
09
0>
0C
#2150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#2160000000
0!
0*
09
0>
0C
#2170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#2180000000
0!
0*
09
0>
0C
#2190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#2200000000
0!
0#
0*
0,
09
0>
0?
0C
#2210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#2220000000
0!
0*
09
0>
0C
#2230000000
1!
1*
19
1>
1C
#2240000000
0!
0*
09
0>
0C
#2250000000
1!
1*
19
1>
1C
#2260000000
0!
0*
09
0>
0C
#2270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#2280000000
0!
0*
09
0>
0C
#2290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#2300000000
0!
0*
09
0>
0C
#2310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#2320000000
0!
0*
09
0>
0C
#2330000000
1!
1*
b10 6
19
1>
1C
b10 G
#2340000000
0!
0*
09
0>
0C
#2350000000
1!
1*
b11 6
19
1>
1C
b11 G
#2360000000
0!
0*
09
0>
0C
#2370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2380000000
0!
0*
09
0>
0C
#2390000000
1!
1*
b101 6
19
1>
1C
b101 G
#2400000000
0!
0*
09
0>
0C
#2410000000
1!
1*
b110 6
19
1>
1C
b110 G
#2420000000
0!
0*
09
0>
0C
#2430000000
1!
1*
b111 6
19
1>
1C
b111 G
#2440000000
0!
0*
09
0>
0C
#2450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#2460000000
0!
0*
09
0>
0C
#2470000000
1!
1*
b1 6
19
1>
1C
b1 G
#2480000000
0!
0*
09
0>
0C
#2490000000
1!
1*
b10 6
19
1>
1C
b10 G
#2500000000
0!
0*
09
0>
0C
#2510000000
1!
1*
b11 6
19
1>
1C
b11 G
#2520000000
0!
0*
09
0>
0C
#2530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2540000000
0!
0*
09
0>
0C
#2550000000
1!
1*
b101 6
19
1>
1C
b101 G
#2560000000
0!
0*
09
0>
0C
#2570000000
1!
1*
b110 6
19
1>
1C
b110 G
#2580000000
0!
0*
09
0>
0C
#2590000000
1!
1*
b111 6
19
1>
1C
b111 G
#2600000000
0!
0*
09
0>
0C
#2610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#2620000000
0!
0*
09
0>
0C
#2630000000
1!
1*
b1 6
19
1>
1C
b1 G
#2640000000
0!
0*
09
0>
0C
#2650000000
1!
1*
b10 6
19
1>
1C
b10 G
#2660000000
0!
0*
09
0>
0C
#2670000000
1!
1*
b11 6
19
1>
1C
b11 G
#2680000000
0!
0*
09
0>
0C
#2690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2700000000
0!
0*
09
0>
0C
#2710000000
1!
1*
b101 6
19
1>
1C
b101 G
#2720000000
0!
0*
09
0>
0C
#2730000000
1!
1*
b110 6
19
1>
1C
b110 G
#2740000000
0!
0*
09
0>
0C
#2750000000
1!
1*
b111 6
19
1>
1C
b111 G
#2760000000
0!
1"
0*
1+
09
1:
0>
0C
#2770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#2780000000
0!
0*
09
0>
0C
#2790000000
1!
1*
b1 6
19
1>
1C
b1 G
#2800000000
0!
0*
09
0>
0C
#2810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#2820000000
0!
0*
09
0>
0C
#2830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#2840000000
0!
0*
09
0>
0C
#2850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#2860000000
0!
0*
09
0>
0C
#2870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#2880000000
0!
0#
0*
0,
09
0>
0?
0C
#2890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#2900000000
0!
0*
09
0>
0C
#2910000000
1!
1*
19
1>
1C
#2920000000
0!
0*
09
0>
0C
#2930000000
1!
1*
19
1>
1C
#2940000000
0!
0*
09
0>
0C
#2950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#2960000000
0!
0*
09
0>
0C
#2970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#2980000000
0!
0*
09
0>
0C
#2990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#3000000000
0!
0*
09
0>
0C
#3010000000
1!
1*
b10 6
19
1>
1C
b10 G
#3020000000
0!
0*
09
0>
0C
#3030000000
1!
1*
b11 6
19
1>
1C
b11 G
#3040000000
0!
0*
09
0>
0C
#3050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3060000000
0!
0*
09
0>
0C
#3070000000
1!
1*
b101 6
19
1>
1C
b101 G
#3080000000
0!
0*
09
0>
0C
#3090000000
1!
1*
b110 6
19
1>
1C
b110 G
#3100000000
0!
0*
09
0>
0C
#3110000000
1!
1*
b111 6
19
1>
1C
b111 G
#3120000000
0!
0*
09
0>
0C
#3130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#3140000000
0!
0*
09
0>
0C
#3150000000
1!
1*
b1 6
19
1>
1C
b1 G
#3160000000
0!
0*
09
0>
0C
#3170000000
1!
1*
b10 6
19
1>
1C
b10 G
#3180000000
0!
0*
09
0>
0C
#3190000000
1!
1*
b11 6
19
1>
1C
b11 G
#3200000000
0!
0*
09
0>
0C
#3210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3220000000
0!
0*
09
0>
0C
#3230000000
1!
1*
b101 6
19
1>
1C
b101 G
#3240000000
0!
0*
09
0>
0C
#3250000000
1!
1*
b110 6
19
1>
1C
b110 G
#3260000000
0!
0*
09
0>
0C
#3270000000
1!
1*
b111 6
19
1>
1C
b111 G
#3280000000
0!
0*
09
0>
0C
#3290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#3300000000
0!
0*
09
0>
0C
#3310000000
1!
1*
b1 6
19
1>
1C
b1 G
#3320000000
0!
0*
09
0>
0C
#3330000000
1!
1*
b10 6
19
1>
1C
b10 G
#3340000000
0!
0*
09
0>
0C
#3350000000
1!
1*
b11 6
19
1>
1C
b11 G
#3360000000
0!
0*
09
0>
0C
#3370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3380000000
0!
0*
09
0>
0C
#3390000000
1!
1*
b101 6
19
1>
1C
b101 G
#3400000000
0!
0*
09
0>
0C
#3410000000
1!
1*
b110 6
19
1>
1C
b110 G
#3420000000
0!
0*
09
0>
0C
#3430000000
1!
1*
b111 6
19
1>
1C
b111 G
#3440000000
0!
1"
0*
1+
09
1:
0>
0C
#3450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#3460000000
0!
0*
09
0>
0C
#3470000000
1!
1*
b1 6
19
1>
1C
b1 G
#3480000000
0!
0*
09
0>
0C
#3490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#3500000000
0!
0*
09
0>
0C
#3510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#3520000000
0!
0*
09
0>
0C
#3530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#3540000000
0!
0*
09
0>
0C
#3550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#3560000000
0!
0#
0*
0,
09
0>
0?
0C
#3570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#3580000000
0!
0*
09
0>
0C
#3590000000
1!
1*
19
1>
1C
#3600000000
0!
0*
09
0>
0C
#3610000000
1!
1*
19
1>
1C
#3620000000
0!
0*
09
0>
0C
#3630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#3640000000
0!
0*
09
0>
0C
#3650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#3660000000
0!
0*
09
0>
0C
#3670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#3680000000
0!
0*
09
0>
0C
#3690000000
1!
1*
b10 6
19
1>
1C
b10 G
#3700000000
0!
0*
09
0>
0C
#3710000000
1!
1*
b11 6
19
1>
1C
b11 G
#3720000000
0!
0*
09
0>
0C
#3730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3740000000
0!
0*
09
0>
0C
#3750000000
1!
1*
b101 6
19
1>
1C
b101 G
#3760000000
0!
0*
09
0>
0C
#3770000000
1!
1*
b110 6
19
1>
1C
b110 G
#3780000000
0!
0*
09
0>
0C
#3790000000
1!
1*
b111 6
19
1>
1C
b111 G
#3800000000
0!
0*
09
0>
0C
#3810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#3820000000
0!
0*
09
0>
0C
#3830000000
1!
1*
b1 6
19
1>
1C
b1 G
#3840000000
0!
0*
09
0>
0C
#3850000000
1!
1*
b10 6
19
1>
1C
b10 G
#3860000000
0!
0*
09
0>
0C
#3870000000
1!
1*
b11 6
19
1>
1C
b11 G
#3880000000
0!
0*
09
0>
0C
#3890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3900000000
0!
0*
09
0>
0C
#3910000000
1!
1*
b101 6
19
1>
1C
b101 G
#3920000000
0!
0*
09
0>
0C
#3930000000
1!
1*
b110 6
19
1>
1C
b110 G
#3940000000
0!
0*
09
0>
0C
#3950000000
1!
1*
b111 6
19
1>
1C
b111 G
#3960000000
0!
0*
09
0>
0C
#3970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#3980000000
0!
0*
09
0>
0C
#3990000000
1!
1*
b1 6
19
1>
1C
b1 G
#4000000000
0!
0*
09
0>
0C
#4010000000
1!
1*
b10 6
19
1>
1C
b10 G
#4020000000
0!
0*
09
0>
0C
#4030000000
1!
1*
b11 6
19
1>
1C
b11 G
#4040000000
0!
0*
09
0>
0C
#4050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4060000000
0!
0*
09
0>
0C
#4070000000
1!
1*
b101 6
19
1>
1C
b101 G
#4080000000
0!
0*
09
0>
0C
#4090000000
1!
1*
b110 6
19
1>
1C
b110 G
#4100000000
0!
0*
09
0>
0C
#4110000000
1!
1*
b111 6
19
1>
1C
b111 G
#4120000000
0!
1"
0*
1+
09
1:
0>
0C
#4130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#4140000000
0!
0*
09
0>
0C
#4150000000
1!
1*
b1 6
19
1>
1C
b1 G
#4160000000
0!
0*
09
0>
0C
#4170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#4180000000
0!
0*
09
0>
0C
#4190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#4200000000
0!
0*
09
0>
0C
#4210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#4220000000
0!
0*
09
0>
0C
#4230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#4240000000
0!
0#
0*
0,
09
0>
0?
0C
#4250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#4260000000
0!
0*
09
0>
0C
#4270000000
1!
1*
19
1>
1C
#4280000000
0!
0*
09
0>
0C
#4290000000
1!
1*
19
1>
1C
#4300000000
0!
0*
09
0>
0C
#4310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#4320000000
0!
0*
09
0>
0C
#4330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#4340000000
0!
0*
09
0>
0C
#4350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#4360000000
0!
0*
09
0>
0C
#4370000000
1!
1*
b10 6
19
1>
1C
b10 G
#4380000000
0!
0*
09
0>
0C
#4390000000
1!
1*
b11 6
19
1>
1C
b11 G
#4400000000
0!
0*
09
0>
0C
#4410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4420000000
0!
0*
09
0>
0C
#4430000000
1!
1*
b101 6
19
1>
1C
b101 G
#4440000000
0!
0*
09
0>
0C
#4450000000
1!
1*
b110 6
19
1>
1C
b110 G
#4460000000
0!
0*
09
0>
0C
#4470000000
1!
1*
b111 6
19
1>
1C
b111 G
#4480000000
0!
0*
09
0>
0C
#4490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#4500000000
0!
0*
09
0>
0C
#4510000000
1!
1*
b1 6
19
1>
1C
b1 G
#4520000000
0!
0*
09
0>
0C
#4530000000
1!
1*
b10 6
19
1>
1C
b10 G
#4540000000
0!
0*
09
0>
0C
#4550000000
1!
1*
b11 6
19
1>
1C
b11 G
#4560000000
0!
0*
09
0>
0C
#4570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4580000000
0!
0*
09
0>
0C
#4590000000
1!
1*
b101 6
19
1>
1C
b101 G
#4600000000
0!
0*
09
0>
0C
#4610000000
1!
1*
b110 6
19
1>
1C
b110 G
#4620000000
0!
0*
09
0>
0C
#4630000000
1!
1*
b111 6
19
1>
1C
b111 G
#4640000000
0!
0*
09
0>
0C
#4650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#4660000000
0!
0*
09
0>
0C
#4670000000
1!
1*
b1 6
19
1>
1C
b1 G
#4680000000
0!
0*
09
0>
0C
#4690000000
1!
1*
b10 6
19
1>
1C
b10 G
#4700000000
0!
0*
09
0>
0C
#4710000000
1!
1*
b11 6
19
1>
1C
b11 G
#4720000000
0!
0*
09
0>
0C
#4730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4740000000
0!
0*
09
0>
0C
#4750000000
1!
1*
b101 6
19
1>
1C
b101 G
#4760000000
0!
0*
09
0>
0C
#4770000000
1!
1*
b110 6
19
1>
1C
b110 G
#4780000000
0!
0*
09
0>
0C
#4790000000
1!
1*
b111 6
19
1>
1C
b111 G
#4800000000
0!
1"
0*
1+
09
1:
0>
0C
#4810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#4820000000
0!
0*
09
0>
0C
#4830000000
1!
1*
b1 6
19
1>
1C
b1 G
#4840000000
0!
0*
09
0>
0C
#4850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#4860000000
0!
0*
09
0>
0C
#4870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#4880000000
0!
0*
09
0>
0C
#4890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#4900000000
0!
0*
09
0>
0C
#4910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#4920000000
0!
0#
0*
0,
09
0>
0?
0C
#4930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#4940000000
0!
0*
09
0>
0C
#4950000000
1!
1*
19
1>
1C
#4960000000
0!
0*
09
0>
0C
#4970000000
1!
1*
19
1>
1C
#4980000000
0!
0*
09
0>
0C
#4990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#5000000000
0!
0*
09
0>
0C
#5010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#5020000000
0!
0*
09
0>
0C
#5030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#5040000000
0!
0*
09
0>
0C
#5050000000
1!
1*
b10 6
19
1>
1C
b10 G
#5060000000
0!
0*
09
0>
0C
#5070000000
1!
1*
b11 6
19
1>
1C
b11 G
#5080000000
0!
0*
09
0>
0C
#5090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5100000000
0!
0*
09
0>
0C
#5110000000
1!
1*
b101 6
19
1>
1C
b101 G
#5120000000
0!
0*
09
0>
0C
#5130000000
1!
1*
b110 6
19
1>
1C
b110 G
#5140000000
0!
0*
09
0>
0C
#5150000000
1!
1*
b111 6
19
1>
1C
b111 G
#5160000000
0!
0*
09
0>
0C
#5170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#5180000000
0!
0*
09
0>
0C
#5190000000
1!
1*
b1 6
19
1>
1C
b1 G
#5200000000
0!
0*
09
0>
0C
#5210000000
1!
1*
b10 6
19
1>
1C
b10 G
#5220000000
0!
0*
09
0>
0C
#5230000000
1!
1*
b11 6
19
1>
1C
b11 G
#5240000000
0!
0*
09
0>
0C
#5250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5260000000
0!
0*
09
0>
0C
#5270000000
1!
1*
b101 6
19
1>
1C
b101 G
#5280000000
0!
0*
09
0>
0C
#5290000000
1!
1*
b110 6
19
1>
1C
b110 G
#5300000000
0!
0*
09
0>
0C
#5310000000
1!
1*
b111 6
19
1>
1C
b111 G
#5320000000
0!
0*
09
0>
0C
#5330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#5340000000
0!
0*
09
0>
0C
#5350000000
1!
1*
b1 6
19
1>
1C
b1 G
#5360000000
0!
0*
09
0>
0C
#5370000000
1!
1*
b10 6
19
1>
1C
b10 G
#5380000000
0!
0*
09
0>
0C
#5390000000
1!
1*
b11 6
19
1>
1C
b11 G
#5400000000
0!
0*
09
0>
0C
#5410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5420000000
0!
0*
09
0>
0C
#5430000000
1!
1*
b101 6
19
1>
1C
b101 G
#5440000000
0!
0*
09
0>
0C
#5450000000
1!
1*
b110 6
19
1>
1C
b110 G
#5460000000
0!
0*
09
0>
0C
#5470000000
1!
1*
b111 6
19
1>
1C
b111 G
#5480000000
0!
1"
0*
1+
09
1:
0>
0C
#5490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#5500000000
0!
0*
09
0>
0C
#5510000000
1!
1*
b1 6
19
1>
1C
b1 G
#5520000000
0!
0*
09
0>
0C
#5530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#5540000000
0!
0*
09
0>
0C
#5550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#5560000000
0!
0*
09
0>
0C
#5570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#5580000000
0!
0*
09
0>
0C
#5590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#5600000000
0!
0#
0*
0,
09
0>
0?
0C
#5610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#5620000000
0!
0*
09
0>
0C
#5630000000
1!
1*
19
1>
1C
#5640000000
0!
0*
09
0>
0C
#5650000000
1!
1*
19
1>
1C
#5660000000
0!
0*
09
0>
0C
#5670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#5680000000
0!
0*
09
0>
0C
#5690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#5700000000
0!
0*
09
0>
0C
#5710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#5720000000
0!
0*
09
0>
0C
#5730000000
1!
1*
b10 6
19
1>
1C
b10 G
#5740000000
0!
0*
09
0>
0C
#5750000000
1!
1*
b11 6
19
1>
1C
b11 G
#5760000000
0!
0*
09
0>
0C
#5770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5780000000
0!
0*
09
0>
0C
#5790000000
1!
1*
b101 6
19
1>
1C
b101 G
#5800000000
0!
0*
09
0>
0C
#5810000000
1!
1*
b110 6
19
1>
1C
b110 G
#5820000000
0!
0*
09
0>
0C
#5830000000
1!
1*
b111 6
19
1>
1C
b111 G
#5840000000
0!
0*
09
0>
0C
#5850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#5860000000
0!
0*
09
0>
0C
#5870000000
1!
1*
b1 6
19
1>
1C
b1 G
#5880000000
0!
0*
09
0>
0C
#5890000000
1!
1*
b10 6
19
1>
1C
b10 G
#5900000000
0!
0*
09
0>
0C
#5910000000
1!
1*
b11 6
19
1>
1C
b11 G
#5920000000
0!
0*
09
0>
0C
#5930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5940000000
0!
0*
09
0>
0C
#5950000000
1!
1*
b101 6
19
1>
1C
b101 G
#5960000000
0!
0*
09
0>
0C
#5970000000
1!
1*
b110 6
19
1>
1C
b110 G
#5980000000
0!
0*
09
0>
0C
#5990000000
1!
1*
b111 6
19
1>
1C
b111 G
#6000000000
0!
0*
09
0>
0C
#6010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#6020000000
0!
0*
09
0>
0C
#6030000000
1!
1*
b1 6
19
1>
1C
b1 G
#6040000000
0!
0*
09
0>
0C
#6050000000
1!
1*
b10 6
19
1>
1C
b10 G
#6060000000
0!
0*
09
0>
0C
#6070000000
1!
1*
b11 6
19
1>
1C
b11 G
#6080000000
0!
0*
09
0>
0C
#6090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6100000000
0!
0*
09
0>
0C
#6110000000
1!
1*
b101 6
19
1>
1C
b101 G
#6120000000
0!
0*
09
0>
0C
#6130000000
1!
1*
b110 6
19
1>
1C
b110 G
#6140000000
0!
0*
09
0>
0C
#6150000000
1!
1*
b111 6
19
1>
1C
b111 G
#6160000000
0!
1"
0*
1+
09
1:
0>
0C
#6170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#6180000000
0!
0*
09
0>
0C
#6190000000
1!
1*
b1 6
19
1>
1C
b1 G
#6200000000
0!
0*
09
0>
0C
#6210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#6220000000
0!
0*
09
0>
0C
#6230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#6240000000
0!
0*
09
0>
0C
#6250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#6260000000
0!
0*
09
0>
0C
#6270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#6280000000
0!
0#
0*
0,
09
0>
0?
0C
#6290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#6300000000
0!
0*
09
0>
0C
#6310000000
1!
1*
19
1>
1C
#6320000000
0!
0*
09
0>
0C
#6330000000
1!
1*
19
1>
1C
#6340000000
0!
0*
09
0>
0C
#6350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#6360000000
0!
0*
09
0>
0C
#6370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#6380000000
0!
0*
09
0>
0C
#6390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#6400000000
0!
0*
09
0>
0C
#6410000000
1!
1*
b10 6
19
1>
1C
b10 G
#6420000000
0!
0*
09
0>
0C
#6430000000
1!
1*
b11 6
19
1>
1C
b11 G
#6440000000
0!
0*
09
0>
0C
#6450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6460000000
0!
0*
09
0>
0C
#6470000000
1!
1*
b101 6
19
1>
1C
b101 G
#6480000000
0!
0*
09
0>
0C
#6490000000
1!
1*
b110 6
19
1>
1C
b110 G
#6500000000
0!
0*
09
0>
0C
#6510000000
1!
1*
b111 6
19
1>
1C
b111 G
#6520000000
0!
0*
09
0>
0C
#6530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#6540000000
0!
0*
09
0>
0C
#6550000000
1!
1*
b1 6
19
1>
1C
b1 G
#6560000000
0!
0*
09
0>
0C
#6570000000
1!
1*
b10 6
19
1>
1C
b10 G
#6580000000
0!
0*
09
0>
0C
#6590000000
1!
1*
b11 6
19
1>
1C
b11 G
#6600000000
0!
0*
09
0>
0C
#6610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6620000000
0!
0*
09
0>
0C
#6630000000
1!
1*
b101 6
19
1>
1C
b101 G
#6640000000
0!
0*
09
0>
0C
#6650000000
1!
1*
b110 6
19
1>
1C
b110 G
#6660000000
0!
0*
09
0>
0C
#6670000000
1!
1*
b111 6
19
1>
1C
b111 G
#6680000000
0!
0*
09
0>
0C
#6690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#6700000000
0!
0*
09
0>
0C
#6710000000
1!
1*
b1 6
19
1>
1C
b1 G
#6720000000
0!
0*
09
0>
0C
#6730000000
1!
1*
b10 6
19
1>
1C
b10 G
#6740000000
0!
0*
09
0>
0C
#6750000000
1!
1*
b11 6
19
1>
1C
b11 G
#6760000000
0!
0*
09
0>
0C
#6770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6780000000
0!
0*
09
0>
0C
#6790000000
1!
1*
b101 6
19
1>
1C
b101 G
#6800000000
0!
0*
09
0>
0C
#6810000000
1!
1*
b110 6
19
1>
1C
b110 G
#6820000000
0!
0*
09
0>
0C
#6830000000
1!
1*
b111 6
19
1>
1C
b111 G
#6840000000
0!
1"
0*
1+
09
1:
0>
0C
#6850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#6860000000
0!
0*
09
0>
0C
#6870000000
1!
1*
b1 6
19
1>
1C
b1 G
#6880000000
0!
0*
09
0>
0C
#6890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#6900000000
0!
0*
09
0>
0C
#6910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#6920000000
0!
0*
09
0>
0C
#6930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#6940000000
0!
0*
09
0>
0C
#6950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#6960000000
0!
0#
0*
0,
09
0>
0?
0C
#6970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#6980000000
0!
0*
09
0>
0C
#6990000000
1!
1*
19
1>
1C
#7000000000
0!
0*
09
0>
0C
#7010000000
1!
1*
19
1>
1C
#7020000000
0!
0*
09
0>
0C
#7030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#7040000000
0!
0*
09
0>
0C
#7050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#7060000000
0!
0*
09
0>
0C
#7070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#7080000000
0!
0*
09
0>
0C
#7090000000
1!
1*
b10 6
19
1>
1C
b10 G
#7100000000
0!
0*
09
0>
0C
#7110000000
1!
1*
b11 6
19
1>
1C
b11 G
#7120000000
0!
0*
09
0>
0C
#7130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7140000000
0!
0*
09
0>
0C
#7150000000
1!
1*
b101 6
19
1>
1C
b101 G
#7160000000
0!
0*
09
0>
0C
#7170000000
1!
1*
b110 6
19
1>
1C
b110 G
#7180000000
0!
0*
09
0>
0C
#7190000000
1!
1*
b111 6
19
1>
1C
b111 G
#7200000000
0!
0*
09
0>
0C
#7210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#7220000000
0!
0*
09
0>
0C
#7230000000
1!
1*
b1 6
19
1>
1C
b1 G
#7240000000
0!
0*
09
0>
0C
#7250000000
1!
1*
b10 6
19
1>
1C
b10 G
#7260000000
0!
0*
09
0>
0C
#7270000000
1!
1*
b11 6
19
1>
1C
b11 G
#7280000000
0!
0*
09
0>
0C
#7290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7300000000
0!
0*
09
0>
0C
#7310000000
1!
1*
b101 6
19
1>
1C
b101 G
#7320000000
0!
0*
09
0>
0C
#7330000000
1!
1*
b110 6
19
1>
1C
b110 G
#7340000000
0!
0*
09
0>
0C
#7350000000
1!
1*
b111 6
19
1>
1C
b111 G
#7360000000
0!
0*
09
0>
0C
#7370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#7380000000
0!
0*
09
0>
0C
#7390000000
1!
1*
b1 6
19
1>
1C
b1 G
#7400000000
0!
0*
09
0>
0C
#7410000000
1!
1*
b10 6
19
1>
1C
b10 G
#7420000000
0!
0*
09
0>
0C
#7430000000
1!
1*
b11 6
19
1>
1C
b11 G
#7440000000
0!
0*
09
0>
0C
#7450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7460000000
0!
0*
09
0>
0C
#7470000000
1!
1*
b101 6
19
1>
1C
b101 G
#7480000000
0!
0*
09
0>
0C
#7490000000
1!
1*
b110 6
19
1>
1C
b110 G
#7500000000
0!
0*
09
0>
0C
#7510000000
1!
1*
b111 6
19
1>
1C
b111 G
#7520000000
0!
1"
0*
1+
09
1:
0>
0C
#7530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#7540000000
0!
0*
09
0>
0C
#7550000000
1!
1*
b1 6
19
1>
1C
b1 G
#7560000000
0!
0*
09
0>
0C
#7570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#7580000000
0!
0*
09
0>
0C
#7590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#7600000000
0!
0*
09
0>
0C
#7610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#7620000000
0!
0*
09
0>
0C
#7630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#7640000000
0!
0#
0*
0,
09
0>
0?
0C
#7650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#7660000000
0!
0*
09
0>
0C
#7670000000
1!
1*
19
1>
1C
#7680000000
0!
0*
09
0>
0C
#7690000000
1!
1*
19
1>
1C
#7700000000
0!
0*
09
0>
0C
#7710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#7720000000
0!
0*
09
0>
0C
#7730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#7740000000
0!
0*
09
0>
0C
#7750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#7760000000
0!
0*
09
0>
0C
#7770000000
1!
1*
b10 6
19
1>
1C
b10 G
#7780000000
0!
0*
09
0>
0C
#7790000000
1!
1*
b11 6
19
1>
1C
b11 G
#7800000000
0!
0*
09
0>
0C
#7810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7820000000
0!
0*
09
0>
0C
#7830000000
1!
1*
b101 6
19
1>
1C
b101 G
#7840000000
0!
0*
09
0>
0C
#7850000000
1!
1*
b110 6
19
1>
1C
b110 G
#7860000000
0!
0*
09
0>
0C
#7870000000
1!
1*
b111 6
19
1>
1C
b111 G
#7880000000
0!
0*
09
0>
0C
#7890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#7900000000
0!
0*
09
0>
0C
#7910000000
1!
1*
b1 6
19
1>
1C
b1 G
#7920000000
0!
0*
09
0>
0C
#7930000000
1!
1*
b10 6
19
1>
1C
b10 G
#7940000000
0!
0*
09
0>
0C
#7950000000
1!
1*
b11 6
19
1>
1C
b11 G
#7960000000
0!
0*
09
0>
0C
#7970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7980000000
0!
0*
09
0>
0C
#7990000000
1!
1*
b101 6
19
1>
1C
b101 G
#8000000000
0!
0*
09
0>
0C
#8010000000
1!
1*
b110 6
19
1>
1C
b110 G
#8020000000
0!
0*
09
0>
0C
#8030000000
1!
1*
b111 6
19
1>
1C
b111 G
#8040000000
0!
0*
09
0>
0C
#8050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#8060000000
0!
0*
09
0>
0C
#8070000000
1!
1*
b1 6
19
1>
1C
b1 G
#8080000000
0!
0*
09
0>
0C
#8090000000
1!
1*
b10 6
19
1>
1C
b10 G
#8100000000
0!
0*
09
0>
0C
#8110000000
1!
1*
b11 6
19
1>
1C
b11 G
#8120000000
0!
0*
09
0>
0C
#8130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8140000000
0!
0*
09
0>
0C
#8150000000
1!
1*
b101 6
19
1>
1C
b101 G
#8160000000
0!
0*
09
0>
0C
#8170000000
1!
1*
b110 6
19
1>
1C
b110 G
#8180000000
0!
0*
09
0>
0C
#8190000000
1!
1*
b111 6
19
1>
1C
b111 G
#8200000000
0!
1"
0*
1+
09
1:
0>
0C
#8210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#8220000000
0!
0*
09
0>
0C
#8230000000
1!
1*
b1 6
19
1>
1C
b1 G
#8240000000
0!
0*
09
0>
0C
#8250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#8260000000
0!
0*
09
0>
0C
#8270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#8280000000
0!
0*
09
0>
0C
#8290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#8300000000
0!
0*
09
0>
0C
#8310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#8320000000
0!
0#
0*
0,
09
0>
0?
0C
#8330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#8340000000
0!
0*
09
0>
0C
#8350000000
1!
1*
19
1>
1C
#8360000000
0!
0*
09
0>
0C
#8370000000
1!
1*
19
1>
1C
#8380000000
0!
0*
09
0>
0C
#8390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#8400000000
0!
0*
09
0>
0C
#8410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#8420000000
0!
0*
09
0>
0C
#8430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#8440000000
0!
0*
09
0>
0C
#8450000000
1!
1*
b10 6
19
1>
1C
b10 G
#8460000000
0!
0*
09
0>
0C
#8470000000
1!
1*
b11 6
19
1>
1C
b11 G
#8480000000
0!
0*
09
0>
0C
#8490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8500000000
0!
0*
09
0>
0C
#8510000000
1!
1*
b101 6
19
1>
1C
b101 G
#8520000000
0!
0*
09
0>
0C
#8530000000
1!
1*
b110 6
19
1>
1C
b110 G
#8540000000
0!
0*
09
0>
0C
#8550000000
1!
1*
b111 6
19
1>
1C
b111 G
#8560000000
0!
0*
09
0>
0C
#8570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#8580000000
0!
0*
09
0>
0C
#8590000000
1!
1*
b1 6
19
1>
1C
b1 G
#8600000000
0!
0*
09
0>
0C
#8610000000
1!
1*
b10 6
19
1>
1C
b10 G
#8620000000
0!
0*
09
0>
0C
#8630000000
1!
1*
b11 6
19
1>
1C
b11 G
#8640000000
0!
0*
09
0>
0C
#8650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8660000000
0!
0*
09
0>
0C
#8670000000
1!
1*
b101 6
19
1>
1C
b101 G
#8680000000
0!
0*
09
0>
0C
#8690000000
1!
1*
b110 6
19
1>
1C
b110 G
#8700000000
0!
0*
09
0>
0C
#8710000000
1!
1*
b111 6
19
1>
1C
b111 G
#8720000000
0!
0*
09
0>
0C
#8730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#8740000000
0!
0*
09
0>
0C
#8750000000
1!
1*
b1 6
19
1>
1C
b1 G
#8760000000
0!
0*
09
0>
0C
#8770000000
1!
1*
b10 6
19
1>
1C
b10 G
#8780000000
0!
0*
09
0>
0C
#8790000000
1!
1*
b11 6
19
1>
1C
b11 G
#8800000000
0!
0*
09
0>
0C
#8810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8820000000
0!
0*
09
0>
0C
#8830000000
1!
1*
b101 6
19
1>
1C
b101 G
#8840000000
0!
0*
09
0>
0C
#8850000000
1!
1*
b110 6
19
1>
1C
b110 G
#8860000000
0!
0*
09
0>
0C
#8870000000
1!
1*
b111 6
19
1>
1C
b111 G
#8880000000
0!
1"
0*
1+
09
1:
0>
0C
#8890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#8900000000
0!
0*
09
0>
0C
#8910000000
1!
1*
b1 6
19
1>
1C
b1 G
#8920000000
0!
0*
09
0>
0C
#8930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#8940000000
0!
0*
09
0>
0C
#8950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#8960000000
0!
0*
09
0>
0C
#8970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#8980000000
0!
0*
09
0>
0C
#8990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#9000000000
0!
0#
0*
0,
09
0>
0?
0C
#9010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#9020000000
0!
0*
09
0>
0C
#9030000000
1!
1*
19
1>
1C
#9040000000
0!
0*
09
0>
0C
#9050000000
1!
1*
19
1>
1C
#9060000000
0!
0*
09
0>
0C
#9070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#9080000000
0!
0*
09
0>
0C
#9090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#9100000000
0!
0*
09
0>
0C
#9110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#9120000000
0!
0*
09
0>
0C
#9130000000
1!
1*
b10 6
19
1>
1C
b10 G
#9140000000
0!
0*
09
0>
0C
#9150000000
1!
1*
b11 6
19
1>
1C
b11 G
#9160000000
0!
0*
09
0>
0C
#9170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#9180000000
0!
0*
09
0>
0C
#9190000000
1!
1*
b101 6
19
1>
1C
b101 G
#9200000000
0!
0*
09
0>
0C
#9210000000
1!
1*
b110 6
19
1>
1C
b110 G
#9220000000
0!
0*
09
0>
0C
#9230000000
1!
1*
b111 6
19
1>
1C
b111 G
#9240000000
0!
0*
09
0>
0C
#9250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#9260000000
0!
0*
09
0>
0C
#9270000000
1!
1*
b1 6
19
1>
1C
b1 G
#9280000000
0!
0*
09
0>
0C
#9290000000
1!
1*
b10 6
19
1>
1C
b10 G
#9300000000
0!
0*
09
0>
0C
#9310000000
1!
1*
b11 6
19
1>
1C
b11 G
#9320000000
0!
0*
09
0>
0C
#9330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#9340000000
0!
0*
09
0>
0C
#9350000000
1!
1*
b101 6
19
1>
1C
b101 G
#9360000000
0!
0*
09
0>
0C
#9370000000
1!
1*
b110 6
19
1>
1C
b110 G
#9380000000
0!
0*
09
0>
0C
#9390000000
1!
1*
b111 6
19
1>
1C
b111 G
#9400000000
0!
0*
09
0>
0C
#9410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#9420000000
0!
0*
09
0>
0C
#9430000000
1!
1*
b1 6
19
1>
1C
b1 G
#9440000000
0!
0*
09
0>
0C
#9450000000
1!
1*
b10 6
19
1>
1C
b10 G
#9460000000
0!
0*
09
0>
0C
#9470000000
1!
1*
b11 6
19
1>
1C
b11 G
#9480000000
0!
0*
09
0>
0C
#9490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#9500000000
0!
0*
09
0>
0C
#9510000000
1!
1*
b101 6
19
1>
1C
b101 G
#9520000000
0!
0*
09
0>
0C
#9530000000
1!
1*
b110 6
19
1>
1C
b110 G
#9540000000
0!
0*
09
0>
0C
#9550000000
1!
1*
b111 6
19
1>
1C
b111 G
#9560000000
0!
1"
0*
1+
09
1:
0>
0C
#9570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#9580000000
0!
0*
09
0>
0C
#9590000000
1!
1*
b1 6
19
1>
1C
b1 G
#9600000000
0!
0*
09
0>
0C
#9610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#9620000000
0!
0*
09
0>
0C
#9630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#9640000000
0!
0*
09
0>
0C
#9650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#9660000000
0!
0*
09
0>
0C
#9670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#9680000000
0!
0#
0*
0,
09
0>
0?
0C
#9690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#9700000000
0!
0*
09
0>
0C
#9710000000
1!
1*
19
1>
1C
#9720000000
0!
0*
09
0>
0C
#9730000000
1!
1*
19
1>
1C
#9740000000
0!
0*
09
0>
0C
#9750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#9760000000
0!
0*
09
0>
0C
#9770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#9780000000
0!
0*
09
0>
0C
#9790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#9800000000
0!
0*
09
0>
0C
#9810000000
1!
1*
b10 6
19
1>
1C
b10 G
#9820000000
0!
0*
09
0>
0C
#9830000000
1!
1*
b11 6
19
1>
1C
b11 G
#9840000000
0!
0*
09
0>
0C
#9850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#9860000000
0!
0*
09
0>
0C
#9870000000
1!
1*
b101 6
19
1>
1C
b101 G
#9880000000
0!
0*
09
0>
0C
#9890000000
1!
1*
b110 6
19
1>
1C
b110 G
#9900000000
0!
0*
09
0>
0C
#9910000000
1!
1*
b111 6
19
1>
1C
b111 G
#9920000000
0!
0*
09
0>
0C
#9930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#9940000000
0!
0*
09
0>
0C
#9950000000
1!
1*
b1 6
19
1>
1C
b1 G
#9960000000
0!
0*
09
0>
0C
#9970000000
1!
1*
b10 6
19
1>
1C
b10 G
#9980000000
0!
0*
09
0>
0C
#9990000000
1!
1*
b11 6
19
1>
1C
b11 G
#10000000000
0!
0*
09
0>
0C
#10010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#10020000000
0!
0*
09
0>
0C
#10030000000
1!
1*
b101 6
19
1>
1C
b101 G
#10040000000
0!
0*
09
0>
0C
#10050000000
1!
1*
b110 6
19
1>
1C
b110 G
#10060000000
0!
0*
09
0>
0C
#10070000000
1!
1*
b111 6
19
1>
1C
b111 G
#10080000000
0!
0*
09
0>
0C
#10090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#10100000000
0!
0*
09
0>
0C
#10110000000
1!
1*
b1 6
19
1>
1C
b1 G
#10120000000
0!
0*
09
0>
0C
#10130000000
1!
1*
b10 6
19
1>
1C
b10 G
#10140000000
0!
0*
09
0>
0C
#10150000000
1!
1*
b11 6
19
1>
1C
b11 G
#10160000000
0!
0*
09
0>
0C
#10170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#10180000000
0!
0*
09
0>
0C
#10190000000
1!
1*
b101 6
19
1>
1C
b101 G
#10200000000
0!
0*
09
0>
0C
#10210000000
1!
1*
b110 6
19
1>
1C
b110 G
#10220000000
0!
0*
09
0>
0C
#10230000000
1!
1*
b111 6
19
1>
1C
b111 G
#10240000000
0!
1"
0*
1+
09
1:
0>
0C
#10250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#10260000000
0!
0*
09
0>
0C
#10270000000
1!
1*
b1 6
19
1>
1C
b1 G
#10280000000
0!
0*
09
0>
0C
#10290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#10300000000
0!
0*
09
0>
0C
#10310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#10320000000
0!
0*
09
0>
0C
#10330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#10340000000
0!
0*
09
0>
0C
#10350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#10360000000
0!
0#
0*
0,
09
0>
0?
0C
#10370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#10380000000
0!
0*
09
0>
0C
#10390000000
1!
1*
19
1>
1C
#10400000000
0!
0*
09
0>
0C
#10410000000
1!
1*
19
1>
1C
#10420000000
0!
0*
09
0>
0C
#10430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#10440000000
0!
0*
09
0>
0C
#10450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#10460000000
0!
0*
09
0>
0C
#10470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#10480000000
0!
0*
09
0>
0C
#10490000000
1!
1*
b10 6
19
1>
1C
b10 G
#10500000000
0!
0*
09
0>
0C
#10510000000
1!
1*
b11 6
19
1>
1C
b11 G
#10520000000
0!
0*
09
0>
0C
#10530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#10540000000
0!
0*
09
0>
0C
#10550000000
1!
1*
b101 6
19
1>
1C
b101 G
#10560000000
0!
0*
09
0>
0C
#10570000000
1!
1*
b110 6
19
1>
1C
b110 G
#10580000000
0!
0*
09
0>
0C
#10590000000
1!
1*
b111 6
19
1>
1C
b111 G
#10600000000
0!
0*
09
0>
0C
#10610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#10620000000
0!
0*
09
0>
0C
#10630000000
1!
1*
b1 6
19
1>
1C
b1 G
#10640000000
0!
0*
09
0>
0C
#10650000000
1!
1*
b10 6
19
1>
1C
b10 G
#10660000000
0!
0*
09
0>
0C
#10670000000
1!
1*
b11 6
19
1>
1C
b11 G
#10680000000
0!
0*
09
0>
0C
#10690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#10700000000
0!
0*
09
0>
0C
#10710000000
1!
1*
b101 6
19
1>
1C
b101 G
#10720000000
0!
0*
09
0>
0C
#10730000000
1!
1*
b110 6
19
1>
1C
b110 G
#10740000000
0!
0*
09
0>
0C
#10750000000
1!
1*
b111 6
19
1>
1C
b111 G
#10760000000
0!
0*
09
0>
0C
#10770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#10780000000
0!
0*
09
0>
0C
#10790000000
1!
1*
b1 6
19
1>
1C
b1 G
#10800000000
0!
0*
09
0>
0C
#10810000000
1!
1*
b10 6
19
1>
1C
b10 G
#10820000000
0!
0*
09
0>
0C
#10830000000
1!
1*
b11 6
19
1>
1C
b11 G
#10840000000
0!
0*
09
0>
0C
#10850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#10860000000
0!
0*
09
0>
0C
#10870000000
1!
1*
b101 6
19
1>
1C
b101 G
#10880000000
0!
0*
09
0>
0C
#10890000000
1!
1*
b110 6
19
1>
1C
b110 G
#10900000000
0!
0*
09
0>
0C
#10910000000
1!
1*
b111 6
19
1>
1C
b111 G
#10920000000
0!
1"
0*
1+
09
1:
0>
0C
#10930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#10940000000
0!
0*
09
0>
0C
#10950000000
1!
1*
b1 6
19
1>
1C
b1 G
#10960000000
0!
0*
09
0>
0C
#10970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#10980000000
0!
0*
09
0>
0C
#10990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#11000000000
0!
0*
09
0>
0C
#11010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#11020000000
0!
0*
09
0>
0C
#11030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#11040000000
0!
0#
0*
0,
09
0>
0?
0C
#11050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#11060000000
0!
0*
09
0>
0C
#11070000000
1!
1*
19
1>
1C
#11080000000
0!
0*
09
0>
0C
#11090000000
1!
1*
19
1>
1C
#11100000000
0!
0*
09
0>
0C
#11110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#11120000000
0!
0*
09
0>
0C
#11130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#11140000000
0!
0*
09
0>
0C
#11150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#11160000000
0!
0*
09
0>
0C
#11170000000
1!
1*
b10 6
19
1>
1C
b10 G
#11180000000
0!
0*
09
0>
0C
#11190000000
1!
1*
b11 6
19
1>
1C
b11 G
#11200000000
0!
0*
09
0>
0C
#11210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#11220000000
0!
0*
09
0>
0C
#11230000000
1!
1*
b101 6
19
1>
1C
b101 G
#11240000000
0!
0*
09
0>
0C
#11250000000
1!
1*
b110 6
19
1>
1C
b110 G
#11260000000
0!
0*
09
0>
0C
#11270000000
1!
1*
b111 6
19
1>
1C
b111 G
#11280000000
0!
0*
09
0>
0C
#11290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#11300000000
0!
0*
09
0>
0C
#11310000000
1!
1*
b1 6
19
1>
1C
b1 G
#11320000000
0!
0*
09
0>
0C
#11330000000
1!
1*
b10 6
19
1>
1C
b10 G
#11340000000
0!
0*
09
0>
0C
#11350000000
1!
1*
b11 6
19
1>
1C
b11 G
#11360000000
0!
0*
09
0>
0C
#11370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#11380000000
0!
0*
09
0>
0C
#11390000000
1!
1*
b101 6
19
1>
1C
b101 G
#11400000000
0!
0*
09
0>
0C
#11410000000
1!
1*
b110 6
19
1>
1C
b110 G
#11420000000
0!
0*
09
0>
0C
#11430000000
1!
1*
b111 6
19
1>
1C
b111 G
#11440000000
0!
0*
09
0>
0C
#11450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#11460000000
0!
0*
09
0>
0C
#11470000000
1!
1*
b1 6
19
1>
1C
b1 G
#11480000000
0!
0*
09
0>
0C
#11490000000
1!
1*
b10 6
19
1>
1C
b10 G
#11500000000
0!
0*
09
0>
0C
#11510000000
1!
1*
b11 6
19
1>
1C
b11 G
#11520000000
0!
0*
09
0>
0C
#11530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#11540000000
0!
0*
09
0>
0C
#11550000000
1!
1*
b101 6
19
1>
1C
b101 G
#11560000000
0!
0*
09
0>
0C
#11570000000
1!
1*
b110 6
19
1>
1C
b110 G
#11580000000
0!
0*
09
0>
0C
#11590000000
1!
1*
b111 6
19
1>
1C
b111 G
#11600000000
0!
1"
0*
1+
09
1:
0>
0C
#11610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#11620000000
0!
0*
09
0>
0C
#11630000000
1!
1*
b1 6
19
1>
1C
b1 G
#11640000000
0!
0*
09
0>
0C
#11650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#11660000000
0!
0*
09
0>
0C
#11670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#11680000000
0!
0*
09
0>
0C
#11690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#11700000000
0!
0*
09
0>
0C
#11710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#11720000000
0!
0#
0*
0,
09
0>
0?
0C
#11730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#11740000000
0!
0*
09
0>
0C
#11750000000
1!
1*
19
1>
1C
#11760000000
0!
0*
09
0>
0C
#11770000000
1!
1*
19
1>
1C
#11780000000
0!
0*
09
0>
0C
#11790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#11800000000
0!
0*
09
0>
0C
#11810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#11820000000
0!
0*
09
0>
0C
#11830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#11840000000
0!
0*
09
0>
0C
#11850000000
1!
1*
b10 6
19
1>
1C
b10 G
#11860000000
0!
0*
09
0>
0C
#11870000000
1!
1*
b11 6
19
1>
1C
b11 G
#11880000000
0!
0*
09
0>
0C
#11890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#11900000000
0!
0*
09
0>
0C
#11910000000
1!
1*
b101 6
19
1>
1C
b101 G
#11920000000
0!
0*
09
0>
0C
#11930000000
1!
1*
b110 6
19
1>
1C
b110 G
#11940000000
0!
0*
09
0>
0C
#11950000000
1!
1*
b111 6
19
1>
1C
b111 G
#11960000000
0!
0*
09
0>
0C
#11970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#11980000000
0!
0*
09
0>
0C
#11990000000
1!
1*
b1 6
19
1>
1C
b1 G
#12000000000
0!
0*
09
0>
0C
#12010000000
1!
1*
b10 6
19
1>
1C
b10 G
#12020000000
0!
0*
09
0>
0C
#12030000000
1!
1*
b11 6
19
1>
1C
b11 G
#12040000000
0!
0*
09
0>
0C
#12050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#12060000000
0!
0*
09
0>
0C
#12070000000
1!
1*
b101 6
19
1>
1C
b101 G
#12080000000
0!
0*
09
0>
0C
#12090000000
1!
1*
b110 6
19
1>
1C
b110 G
#12100000000
0!
0*
09
0>
0C
#12110000000
1!
1*
b111 6
19
1>
1C
b111 G
#12120000000
0!
0*
09
0>
0C
#12130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#12140000000
0!
0*
09
0>
0C
#12150000000
1!
1*
b1 6
19
1>
1C
b1 G
#12160000000
0!
0*
09
0>
0C
#12170000000
1!
1*
b10 6
19
1>
1C
b10 G
#12180000000
0!
0*
09
0>
0C
#12190000000
1!
1*
b11 6
19
1>
1C
b11 G
#12200000000
0!
0*
09
0>
0C
#12210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#12220000000
0!
0*
09
0>
0C
#12230000000
1!
1*
b101 6
19
1>
1C
b101 G
#12240000000
0!
0*
09
0>
0C
#12250000000
1!
1*
b110 6
19
1>
1C
b110 G
#12260000000
0!
0*
09
0>
0C
#12270000000
1!
1*
b111 6
19
1>
1C
b111 G
#12280000000
0!
1"
0*
1+
09
1:
0>
0C
#12290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#12300000000
0!
0*
09
0>
0C
#12310000000
1!
1*
b1 6
19
1>
1C
b1 G
#12320000000
0!
0*
09
0>
0C
#12330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#12340000000
0!
0*
09
0>
0C
#12350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#12360000000
0!
0*
09
0>
0C
#12370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#12380000000
0!
0*
09
0>
0C
#12390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#12400000000
0!
0#
0*
0,
09
0>
0?
0C
#12410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#12420000000
0!
0*
09
0>
0C
#12430000000
1!
1*
19
1>
1C
#12440000000
0!
0*
09
0>
0C
#12450000000
1!
1*
19
1>
1C
#12460000000
0!
0*
09
0>
0C
#12470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#12480000000
0!
0*
09
0>
0C
#12490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#12500000000
0!
0*
09
0>
0C
#12510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#12520000000
0!
0*
09
0>
0C
#12530000000
1!
1*
b10 6
19
1>
1C
b10 G
#12540000000
0!
0*
09
0>
0C
#12550000000
1!
1*
b11 6
19
1>
1C
b11 G
#12560000000
0!
0*
09
0>
0C
#12570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#12580000000
0!
0*
09
0>
0C
#12590000000
1!
1*
b101 6
19
1>
1C
b101 G
#12600000000
0!
0*
09
0>
0C
#12610000000
1!
1*
b110 6
19
1>
1C
b110 G
#12620000000
0!
0*
09
0>
0C
#12630000000
1!
1*
b111 6
19
1>
1C
b111 G
#12640000000
0!
0*
09
0>
0C
#12650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#12660000000
0!
0*
09
0>
0C
#12670000000
1!
1*
b1 6
19
1>
1C
b1 G
#12680000000
0!
0*
09
0>
0C
#12690000000
1!
1*
b10 6
19
1>
1C
b10 G
#12700000000
0!
0*
09
0>
0C
#12710000000
1!
1*
b11 6
19
1>
1C
b11 G
#12720000000
0!
0*
09
0>
0C
#12730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#12740000000
0!
0*
09
0>
0C
#12750000000
1!
1*
b101 6
19
1>
1C
b101 G
#12760000000
0!
0*
09
0>
0C
#12770000000
1!
1*
b110 6
19
1>
1C
b110 G
#12780000000
0!
0*
09
0>
0C
#12790000000
1!
1*
b111 6
19
1>
1C
b111 G
#12800000000
0!
0*
09
0>
0C
#12810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#12820000000
0!
0*
09
0>
0C
#12830000000
1!
1*
b1 6
19
1>
1C
b1 G
#12840000000
0!
0*
09
0>
0C
#12850000000
1!
1*
b10 6
19
1>
1C
b10 G
#12860000000
0!
0*
09
0>
0C
#12870000000
1!
1*
b11 6
19
1>
1C
b11 G
#12880000000
0!
0*
09
0>
0C
#12890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#12900000000
0!
0*
09
0>
0C
#12910000000
1!
1*
b101 6
19
1>
1C
b101 G
#12920000000
0!
0*
09
0>
0C
#12930000000
1!
1*
b110 6
19
1>
1C
b110 G
#12940000000
0!
0*
09
0>
0C
#12950000000
1!
1*
b111 6
19
1>
1C
b111 G
#12960000000
0!
1"
0*
1+
09
1:
0>
0C
#12970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#12980000000
0!
0*
09
0>
0C
#12990000000
1!
1*
b1 6
19
1>
1C
b1 G
#13000000000
0!
0*
09
0>
0C
#13010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#13020000000
0!
0*
09
0>
0C
#13030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#13040000000
0!
0*
09
0>
0C
#13050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#13060000000
0!
0*
09
0>
0C
#13070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#13080000000
0!
0#
0*
0,
09
0>
0?
0C
#13090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#13100000000
0!
0*
09
0>
0C
#13110000000
1!
1*
19
1>
1C
#13120000000
0!
0*
09
0>
0C
#13130000000
1!
1*
19
1>
1C
#13140000000
0!
0*
09
0>
0C
#13150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#13160000000
0!
0*
09
0>
0C
#13170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#13180000000
0!
0*
09
0>
0C
#13190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#13200000000
0!
0*
09
0>
0C
#13210000000
1!
1*
b10 6
19
1>
1C
b10 G
#13220000000
0!
0*
09
0>
0C
#13230000000
1!
1*
b11 6
19
1>
1C
b11 G
#13240000000
0!
0*
09
0>
0C
#13250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#13260000000
0!
0*
09
0>
0C
#13270000000
1!
1*
b101 6
19
1>
1C
b101 G
#13280000000
0!
0*
09
0>
0C
#13290000000
1!
1*
b110 6
19
1>
1C
b110 G
#13300000000
0!
0*
09
0>
0C
#13310000000
1!
1*
b111 6
19
1>
1C
b111 G
#13320000000
0!
0*
09
0>
0C
#13330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#13340000000
0!
0*
09
0>
0C
#13350000000
1!
1*
b1 6
19
1>
1C
b1 G
#13360000000
0!
0*
09
0>
0C
#13370000000
1!
1*
b10 6
19
1>
1C
b10 G
#13380000000
0!
0*
09
0>
0C
#13390000000
1!
1*
b11 6
19
1>
1C
b11 G
#13400000000
0!
0*
09
0>
0C
#13410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#13420000000
0!
0*
09
0>
0C
#13430000000
1!
1*
b101 6
19
1>
1C
b101 G
#13440000000
0!
0*
09
0>
0C
#13450000000
1!
1*
b110 6
19
1>
1C
b110 G
#13460000000
0!
0*
09
0>
0C
#13470000000
1!
1*
b111 6
19
1>
1C
b111 G
#13480000000
0!
0*
09
0>
0C
#13490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#13500000000
0!
0*
09
0>
0C
#13510000000
1!
1*
b1 6
19
1>
1C
b1 G
#13520000000
0!
0*
09
0>
0C
#13530000000
1!
1*
b10 6
19
1>
1C
b10 G
#13540000000
0!
0*
09
0>
0C
#13550000000
1!
1*
b11 6
19
1>
1C
b11 G
#13560000000
0!
0*
09
0>
0C
#13570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#13580000000
0!
0*
09
0>
0C
#13590000000
1!
1*
b101 6
19
1>
1C
b101 G
#13600000000
0!
0*
09
0>
0C
#13610000000
1!
1*
b110 6
19
1>
1C
b110 G
#13620000000
0!
0*
09
0>
0C
#13630000000
1!
1*
b111 6
19
1>
1C
b111 G
#13640000000
0!
1"
0*
1+
09
1:
0>
0C
#13650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#13660000000
0!
0*
09
0>
0C
#13670000000
1!
1*
b1 6
19
1>
1C
b1 G
#13680000000
0!
0*
09
0>
0C
#13690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#13700000000
0!
0*
09
0>
0C
#13710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#13720000000
0!
0*
09
0>
0C
#13730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#13740000000
0!
0*
09
0>
0C
#13750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#13760000000
0!
0#
0*
0,
09
0>
0?
0C
#13770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#13780000000
0!
0*
09
0>
0C
#13790000000
1!
1*
19
1>
1C
#13800000000
0!
0*
09
0>
0C
#13810000000
1!
1*
19
1>
1C
#13820000000
0!
0*
09
0>
0C
#13830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#13840000000
0!
0*
09
0>
0C
#13850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#13860000000
0!
0*
09
0>
0C
#13870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#13880000000
0!
0*
09
0>
0C
#13890000000
1!
1*
b10 6
19
1>
1C
b10 G
#13900000000
0!
0*
09
0>
0C
#13910000000
1!
1*
b11 6
19
1>
1C
b11 G
#13920000000
0!
0*
09
0>
0C
#13930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#13940000000
0!
0*
09
0>
0C
#13950000000
1!
1*
b101 6
19
1>
1C
b101 G
#13960000000
0!
0*
09
0>
0C
#13970000000
1!
1*
b110 6
19
1>
1C
b110 G
#13980000000
0!
0*
09
0>
0C
#13990000000
1!
1*
b111 6
19
1>
1C
b111 G
#14000000000
0!
0*
09
0>
0C
#14010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#14020000000
0!
0*
09
0>
0C
#14030000000
1!
1*
b1 6
19
1>
1C
b1 G
#14040000000
0!
0*
09
0>
0C
#14050000000
1!
1*
b10 6
19
1>
1C
b10 G
#14060000000
0!
0*
09
0>
0C
#14070000000
1!
1*
b11 6
19
1>
1C
b11 G
#14080000000
0!
0*
09
0>
0C
#14090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#14100000000
0!
0*
09
0>
0C
#14110000000
1!
1*
b101 6
19
1>
1C
b101 G
#14120000000
0!
0*
09
0>
0C
#14130000000
1!
1*
b110 6
19
1>
1C
b110 G
#14140000000
0!
0*
09
0>
0C
#14150000000
1!
1*
b111 6
19
1>
1C
b111 G
#14160000000
0!
0*
09
0>
0C
#14170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#14180000000
0!
0*
09
0>
0C
#14190000000
1!
1*
b1 6
19
1>
1C
b1 G
#14200000000
0!
0*
09
0>
0C
#14210000000
1!
1*
b10 6
19
1>
1C
b10 G
#14220000000
0!
0*
09
0>
0C
#14230000000
1!
1*
b11 6
19
1>
1C
b11 G
#14240000000
0!
0*
09
0>
0C
#14250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#14260000000
0!
0*
09
0>
0C
#14270000000
1!
1*
b101 6
19
1>
1C
b101 G
#14280000000
0!
0*
09
0>
0C
#14290000000
1!
1*
b110 6
19
1>
1C
b110 G
#14300000000
0!
0*
09
0>
0C
#14310000000
1!
1*
b111 6
19
1>
1C
b111 G
#14320000000
0!
1"
0*
1+
09
1:
0>
0C
#14330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#14340000000
0!
0*
09
0>
0C
#14350000000
1!
1*
b1 6
19
1>
1C
b1 G
#14360000000
0!
0*
09
0>
0C
#14370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#14380000000
0!
0*
09
0>
0C
#14390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#14400000000
0!
0*
09
0>
0C
#14410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#14420000000
0!
0*
09
0>
0C
#14430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#14440000000
0!
0#
0*
0,
09
0>
0?
0C
#14450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#14460000000
0!
0*
09
0>
0C
#14470000000
1!
1*
19
1>
1C
#14480000000
0!
0*
09
0>
0C
#14490000000
1!
1*
19
1>
1C
#14500000000
0!
0*
09
0>
0C
#14510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#14520000000
0!
0*
09
0>
0C
#14530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#14540000000
0!
0*
09
0>
0C
#14550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#14560000000
0!
0*
09
0>
0C
#14570000000
1!
1*
b10 6
19
1>
1C
b10 G
#14580000000
0!
0*
09
0>
0C
#14590000000
1!
1*
b11 6
19
1>
1C
b11 G
#14600000000
0!
0*
09
0>
0C
#14610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#14620000000
0!
0*
09
0>
0C
#14630000000
1!
1*
b101 6
19
1>
1C
b101 G
#14640000000
0!
0*
09
0>
0C
#14650000000
1!
1*
b110 6
19
1>
1C
b110 G
#14660000000
0!
0*
09
0>
0C
#14670000000
1!
1*
b111 6
19
1>
1C
b111 G
#14680000000
0!
0*
09
0>
0C
#14690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#14700000000
0!
0*
09
0>
0C
#14710000000
1!
1*
b1 6
19
1>
1C
b1 G
#14720000000
0!
0*
09
0>
0C
#14730000000
1!
1*
b10 6
19
1>
1C
b10 G
#14740000000
0!
0*
09
0>
0C
#14750000000
1!
1*
b11 6
19
1>
1C
b11 G
#14760000000
0!
0*
09
0>
0C
#14770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#14780000000
0!
0*
09
0>
0C
#14790000000
1!
1*
b101 6
19
1>
1C
b101 G
#14800000000
0!
0*
09
0>
0C
#14810000000
1!
1*
b110 6
19
1>
1C
b110 G
#14820000000
0!
0*
09
0>
0C
#14830000000
1!
1*
b111 6
19
1>
1C
b111 G
#14840000000
0!
0*
09
0>
0C
#14850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#14860000000
0!
0*
09
0>
0C
#14870000000
1!
1*
b1 6
19
1>
1C
b1 G
#14880000000
0!
0*
09
0>
0C
#14890000000
1!
1*
b10 6
19
1>
1C
b10 G
#14900000000
0!
0*
09
0>
0C
#14910000000
1!
1*
b11 6
19
1>
1C
b11 G
#14920000000
0!
0*
09
0>
0C
#14930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#14940000000
0!
0*
09
0>
0C
#14950000000
1!
1*
b101 6
19
1>
1C
b101 G
#14960000000
0!
0*
09
0>
0C
#14970000000
1!
1*
b110 6
19
1>
1C
b110 G
#14980000000
0!
0*
09
0>
0C
#14990000000
1!
1*
b111 6
19
1>
1C
b111 G
#15000000000
0!
1"
0*
1+
09
1:
0>
0C
#15010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#15020000000
0!
0*
09
0>
0C
#15030000000
1!
1*
b1 6
19
1>
1C
b1 G
#15040000000
0!
0*
09
0>
0C
#15050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#15060000000
0!
0*
09
0>
0C
#15070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#15080000000
0!
0*
09
0>
0C
#15090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#15100000000
0!
0*
09
0>
0C
#15110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#15120000000
0!
0#
0*
0,
09
0>
0?
0C
#15130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#15140000000
0!
0*
09
0>
0C
#15150000000
1!
1*
19
1>
1C
#15160000000
0!
0*
09
0>
0C
#15170000000
1!
1*
19
1>
1C
#15180000000
0!
0*
09
0>
0C
#15190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#15200000000
0!
0*
09
0>
0C
#15210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#15220000000
0!
0*
09
0>
0C
#15230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#15240000000
0!
0*
09
0>
0C
#15250000000
1!
1*
b10 6
19
1>
1C
b10 G
#15260000000
0!
0*
09
0>
0C
#15270000000
1!
1*
b11 6
19
1>
1C
b11 G
#15280000000
0!
0*
09
0>
0C
#15290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#15300000000
0!
0*
09
0>
0C
#15310000000
1!
1*
b101 6
19
1>
1C
b101 G
#15320000000
0!
0*
09
0>
0C
#15330000000
1!
1*
b110 6
19
1>
1C
b110 G
#15340000000
0!
0*
09
0>
0C
#15350000000
1!
1*
b111 6
19
1>
1C
b111 G
#15360000000
0!
0*
09
0>
0C
#15370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#15380000000
0!
0*
09
0>
0C
#15390000000
1!
1*
b1 6
19
1>
1C
b1 G
#15400000000
0!
0*
09
0>
0C
#15410000000
1!
1*
b10 6
19
1>
1C
b10 G
#15420000000
0!
0*
09
0>
0C
#15430000000
1!
1*
b11 6
19
1>
1C
b11 G
#15440000000
0!
0*
09
0>
0C
#15450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#15460000000
0!
0*
09
0>
0C
#15470000000
1!
1*
b101 6
19
1>
1C
b101 G
#15480000000
0!
0*
09
0>
0C
#15490000000
1!
1*
b110 6
19
1>
1C
b110 G
#15500000000
0!
0*
09
0>
0C
#15510000000
1!
1*
b111 6
19
1>
1C
b111 G
#15520000000
0!
0*
09
0>
0C
#15530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#15540000000
0!
0*
09
0>
0C
#15550000000
1!
1*
b1 6
19
1>
1C
b1 G
#15560000000
0!
0*
09
0>
0C
#15570000000
1!
1*
b10 6
19
1>
1C
b10 G
#15580000000
0!
0*
09
0>
0C
#15590000000
1!
1*
b11 6
19
1>
1C
b11 G
#15600000000
0!
0*
09
0>
0C
#15610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#15620000000
0!
0*
09
0>
0C
#15630000000
1!
1*
b101 6
19
1>
1C
b101 G
#15640000000
0!
0*
09
0>
0C
#15650000000
1!
1*
b110 6
19
1>
1C
b110 G
#15660000000
0!
0*
09
0>
0C
#15670000000
1!
1*
b111 6
19
1>
1C
b111 G
#15680000000
0!
1"
0*
1+
09
1:
0>
0C
#15690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#15700000000
0!
0*
09
0>
0C
#15710000000
1!
1*
b1 6
19
1>
1C
b1 G
#15720000000
0!
0*
09
0>
0C
#15730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#15740000000
0!
0*
09
0>
0C
#15750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#15760000000
0!
0*
09
0>
0C
#15770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#15780000000
0!
0*
09
0>
0C
#15790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#15800000000
0!
0#
0*
0,
09
0>
0?
0C
#15810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#15820000000
0!
0*
09
0>
0C
#15830000000
1!
1*
19
1>
1C
#15840000000
0!
0*
09
0>
0C
#15850000000
1!
1*
19
1>
1C
#15860000000
0!
0*
09
0>
0C
#15870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#15880000000
0!
0*
09
0>
0C
#15890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#15900000000
0!
0*
09
0>
0C
#15910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#15920000000
0!
0*
09
0>
0C
#15930000000
1!
1*
b10 6
19
1>
1C
b10 G
#15940000000
0!
0*
09
0>
0C
#15950000000
1!
1*
b11 6
19
1>
1C
b11 G
#15960000000
0!
0*
09
0>
0C
#15970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#15980000000
0!
0*
09
0>
0C
#15990000000
1!
1*
b101 6
19
1>
1C
b101 G
#16000000000
0!
0*
09
0>
0C
#16010000000
1!
1*
b110 6
19
1>
1C
b110 G
#16020000000
0!
0*
09
0>
0C
#16030000000
1!
1*
b111 6
19
1>
1C
b111 G
#16040000000
0!
0*
09
0>
0C
#16050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#16060000000
0!
0*
09
0>
0C
#16070000000
1!
1*
b1 6
19
1>
1C
b1 G
#16080000000
0!
0*
09
0>
0C
#16090000000
1!
1*
b10 6
19
1>
1C
b10 G
#16100000000
0!
0*
09
0>
0C
#16110000000
1!
1*
b11 6
19
1>
1C
b11 G
#16120000000
0!
0*
09
0>
0C
#16130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#16140000000
0!
0*
09
0>
0C
#16150000000
1!
1*
b101 6
19
1>
1C
b101 G
#16160000000
0!
0*
09
0>
0C
#16170000000
1!
1*
b110 6
19
1>
1C
b110 G
#16180000000
0!
0*
09
0>
0C
#16190000000
1!
1*
b111 6
19
1>
1C
b111 G
#16200000000
0!
0*
09
0>
0C
#16210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#16220000000
0!
0*
09
0>
0C
#16230000000
1!
1*
b1 6
19
1>
1C
b1 G
#16240000000
0!
0*
09
0>
0C
#16250000000
1!
1*
b10 6
19
1>
1C
b10 G
#16260000000
0!
0*
09
0>
0C
#16270000000
1!
1*
b11 6
19
1>
1C
b11 G
#16280000000
0!
0*
09
0>
0C
#16290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#16300000000
0!
0*
09
0>
0C
#16310000000
1!
1*
b101 6
19
1>
1C
b101 G
#16320000000
0!
0*
09
0>
0C
#16330000000
1!
1*
b110 6
19
1>
1C
b110 G
#16340000000
0!
0*
09
0>
0C
#16350000000
1!
1*
b111 6
19
1>
1C
b111 G
#16360000000
0!
1"
0*
1+
09
1:
0>
0C
#16370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#16380000000
0!
0*
09
0>
0C
#16390000000
1!
1*
b1 6
19
1>
1C
b1 G
#16400000000
0!
0*
09
0>
0C
#16410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#16420000000
0!
0*
09
0>
0C
#16430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#16440000000
0!
0*
09
0>
0C
#16450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#16460000000
0!
0*
09
0>
0C
#16470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#16480000000
0!
0#
0*
0,
09
0>
0?
0C
#16490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#16500000000
0!
0*
09
0>
0C
#16510000000
1!
1*
19
1>
1C
#16520000000
0!
0*
09
0>
0C
#16530000000
1!
1*
19
1>
1C
#16540000000
0!
0*
09
0>
0C
#16550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#16560000000
0!
0*
09
0>
0C
#16570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#16580000000
0!
0*
09
0>
0C
#16590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#16600000000
0!
0*
09
0>
0C
#16610000000
1!
1*
b10 6
19
1>
1C
b10 G
#16620000000
0!
0*
09
0>
0C
#16630000000
1!
1*
b11 6
19
1>
1C
b11 G
#16640000000
0!
0*
09
0>
0C
#16650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#16660000000
0!
0*
09
0>
0C
#16670000000
1!
1*
b101 6
19
1>
1C
b101 G
#16680000000
0!
0*
09
0>
0C
#16690000000
1!
1*
b110 6
19
1>
1C
b110 G
#16700000000
0!
0*
09
0>
0C
#16710000000
1!
1*
b111 6
19
1>
1C
b111 G
#16720000000
0!
0*
09
0>
0C
#16730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#16740000000
0!
0*
09
0>
0C
#16750000000
1!
1*
b1 6
19
1>
1C
b1 G
#16760000000
0!
0*
09
0>
0C
#16770000000
1!
1*
b10 6
19
1>
1C
b10 G
#16780000000
0!
0*
09
0>
0C
#16790000000
1!
1*
b11 6
19
1>
1C
b11 G
#16800000000
0!
0*
09
0>
0C
#16810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#16820000000
0!
0*
09
0>
0C
#16830000000
1!
1*
b101 6
19
1>
1C
b101 G
#16840000000
0!
0*
09
0>
0C
#16850000000
1!
1*
b110 6
19
1>
1C
b110 G
#16860000000
0!
0*
09
0>
0C
#16870000000
1!
1*
b111 6
19
1>
1C
b111 G
#16880000000
0!
0*
09
0>
0C
#16890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#16900000000
0!
0*
09
0>
0C
#16910000000
1!
1*
b1 6
19
1>
1C
b1 G
#16920000000
0!
0*
09
0>
0C
#16930000000
1!
1*
b10 6
19
1>
1C
b10 G
#16940000000
0!
0*
09
0>
0C
#16950000000
1!
1*
b11 6
19
1>
1C
b11 G
#16960000000
0!
0*
09
0>
0C
#16970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#16980000000
0!
0*
09
0>
0C
#16990000000
1!
1*
b101 6
19
1>
1C
b101 G
#17000000000
0!
0*
09
0>
0C
#17010000000
1!
1*
b110 6
19
1>
1C
b110 G
#17020000000
0!
0*
09
0>
0C
#17030000000
1!
1*
b111 6
19
1>
1C
b111 G
#17040000000
0!
1"
0*
1+
09
1:
0>
0C
#17050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#17060000000
0!
0*
09
0>
0C
#17070000000
1!
1*
b1 6
19
1>
1C
b1 G
#17080000000
0!
0*
09
0>
0C
#17090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#17100000000
0!
0*
09
0>
0C
#17110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#17120000000
0!
0*
09
0>
0C
#17130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#17140000000
0!
0*
09
0>
0C
#17150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#17160000000
0!
0#
0*
0,
09
0>
0?
0C
#17170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#17180000000
0!
0*
09
0>
0C
#17190000000
1!
1*
19
1>
1C
#17200000000
0!
0*
09
0>
0C
#17210000000
1!
1*
19
1>
1C
#17220000000
0!
0*
09
0>
0C
#17230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#17240000000
0!
0*
09
0>
0C
#17250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#17260000000
0!
0*
09
0>
0C
#17270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#17280000000
0!
0*
09
0>
0C
#17290000000
1!
1*
b10 6
19
1>
1C
b10 G
#17300000000
0!
0*
09
0>
0C
#17310000000
1!
1*
b11 6
19
1>
1C
b11 G
#17320000000
0!
0*
09
0>
0C
#17330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#17340000000
0!
0*
09
0>
0C
#17350000000
1!
1*
b101 6
19
1>
1C
b101 G
#17360000000
0!
0*
09
0>
0C
#17370000000
1!
1*
b110 6
19
1>
1C
b110 G
#17380000000
0!
0*
09
0>
0C
#17390000000
1!
1*
b111 6
19
1>
1C
b111 G
#17400000000
0!
0*
09
0>
0C
#17410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#17420000000
0!
0*
09
0>
0C
#17430000000
1!
1*
b1 6
19
1>
1C
b1 G
#17440000000
0!
0*
09
0>
0C
#17450000000
1!
1*
b10 6
19
1>
1C
b10 G
#17460000000
0!
0*
09
0>
0C
#17470000000
1!
1*
b11 6
19
1>
1C
b11 G
#17480000000
0!
0*
09
0>
0C
#17490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#17500000000
0!
0*
09
0>
0C
#17510000000
1!
1*
b101 6
19
1>
1C
b101 G
#17520000000
0!
0*
09
0>
0C
#17530000000
1!
1*
b110 6
19
1>
1C
b110 G
#17540000000
0!
0*
09
0>
0C
#17550000000
1!
1*
b111 6
19
1>
1C
b111 G
#17560000000
0!
0*
09
0>
0C
#17570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#17580000000
0!
0*
09
0>
0C
#17590000000
1!
1*
b1 6
19
1>
1C
b1 G
#17600000000
0!
0*
09
0>
0C
#17610000000
1!
1*
b10 6
19
1>
1C
b10 G
#17620000000
0!
0*
09
0>
0C
#17630000000
1!
1*
b11 6
19
1>
1C
b11 G
#17640000000
0!
0*
09
0>
0C
#17650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#17660000000
0!
0*
09
0>
0C
#17670000000
1!
1*
b101 6
19
1>
1C
b101 G
#17680000000
0!
0*
09
0>
0C
#17690000000
1!
1*
b110 6
19
1>
1C
b110 G
#17700000000
0!
0*
09
0>
0C
#17710000000
1!
1*
b111 6
19
1>
1C
b111 G
#17720000000
0!
1"
0*
1+
09
1:
0>
0C
#17730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#17740000000
0!
0*
09
0>
0C
#17750000000
1!
1*
b1 6
19
1>
1C
b1 G
#17760000000
0!
0*
09
0>
0C
#17770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#17780000000
0!
0*
09
0>
0C
#17790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#17800000000
0!
0*
09
0>
0C
#17810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#17820000000
0!
0*
09
0>
0C
#17830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#17840000000
0!
0#
0*
0,
09
0>
0?
0C
#17850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#17860000000
0!
0*
09
0>
0C
#17870000000
1!
1*
19
1>
1C
#17880000000
0!
0*
09
0>
0C
#17890000000
1!
1*
19
1>
1C
#17900000000
0!
0*
09
0>
0C
#17910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#17920000000
0!
0*
09
0>
0C
#17930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#17940000000
0!
0*
09
0>
0C
#17950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#17960000000
0!
0*
09
0>
0C
#17970000000
1!
1*
b10 6
19
1>
1C
b10 G
#17980000000
0!
0*
09
0>
0C
#17990000000
1!
1*
b11 6
19
1>
1C
b11 G
#18000000000
0!
0*
09
0>
0C
#18010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#18020000000
0!
0*
09
0>
0C
#18030000000
1!
1*
b101 6
19
1>
1C
b101 G
#18040000000
0!
0*
09
0>
0C
#18050000000
1!
1*
b110 6
19
1>
1C
b110 G
#18060000000
0!
0*
09
0>
0C
#18070000000
1!
1*
b111 6
19
1>
1C
b111 G
#18080000000
0!
0*
09
0>
0C
#18090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#18100000000
0!
0*
09
0>
0C
#18110000000
1!
1*
b1 6
19
1>
1C
b1 G
#18120000000
0!
0*
09
0>
0C
#18130000000
1!
1*
b10 6
19
1>
1C
b10 G
#18140000000
0!
0*
09
0>
0C
#18150000000
1!
1*
b11 6
19
1>
1C
b11 G
#18160000000
0!
0*
09
0>
0C
#18170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#18180000000
0!
0*
09
0>
0C
#18190000000
1!
1*
b101 6
19
1>
1C
b101 G
#18200000000
0!
0*
09
0>
0C
#18210000000
1!
1*
b110 6
19
1>
1C
b110 G
#18220000000
0!
0*
09
0>
0C
#18230000000
1!
1*
b111 6
19
1>
1C
b111 G
#18240000000
0!
0*
09
0>
0C
#18250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#18260000000
0!
0*
09
0>
0C
#18270000000
1!
1*
b1 6
19
1>
1C
b1 G
#18280000000
0!
0*
09
0>
0C
#18290000000
1!
1*
b10 6
19
1>
1C
b10 G
#18300000000
0!
0*
09
0>
0C
#18310000000
1!
1*
b11 6
19
1>
1C
b11 G
#18320000000
0!
0*
09
0>
0C
#18330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#18340000000
0!
0*
09
0>
0C
#18350000000
1!
1*
b101 6
19
1>
1C
b101 G
#18360000000
0!
0*
09
0>
0C
#18370000000
1!
1*
b110 6
19
1>
1C
b110 G
#18380000000
0!
0*
09
0>
0C
#18390000000
1!
1*
b111 6
19
1>
1C
b111 G
#18400000000
0!
1"
0*
1+
09
1:
0>
0C
#18410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#18420000000
0!
0*
09
0>
0C
#18430000000
1!
1*
b1 6
19
1>
1C
b1 G
#18440000000
0!
0*
09
0>
0C
#18450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#18460000000
0!
0*
09
0>
0C
#18470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#18480000000
0!
0*
09
0>
0C
#18490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#18500000000
0!
0*
09
0>
0C
#18510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#18520000000
0!
0#
0*
0,
09
0>
0?
0C
#18530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#18540000000
0!
0*
09
0>
0C
#18550000000
1!
1*
19
1>
1C
#18560000000
0!
0*
09
0>
0C
#18570000000
1!
1*
19
1>
1C
#18580000000
0!
0*
09
0>
0C
#18590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#18600000000
0!
0*
09
0>
0C
#18610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#18620000000
0!
0*
09
0>
0C
#18630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#18640000000
0!
0*
09
0>
0C
#18650000000
1!
1*
b10 6
19
1>
1C
b10 G
#18660000000
0!
0*
09
0>
0C
#18670000000
1!
1*
b11 6
19
1>
1C
b11 G
#18680000000
0!
0*
09
0>
0C
#18690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#18700000000
0!
0*
09
0>
0C
#18710000000
1!
1*
b101 6
19
1>
1C
b101 G
#18720000000
0!
0*
09
0>
0C
#18730000000
1!
1*
b110 6
19
1>
1C
b110 G
#18740000000
0!
0*
09
0>
0C
#18750000000
1!
1*
b111 6
19
1>
1C
b111 G
#18760000000
0!
0*
09
0>
0C
#18770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#18780000000
0!
0*
09
0>
0C
#18790000000
1!
1*
b1 6
19
1>
1C
b1 G
#18800000000
0!
0*
09
0>
0C
#18810000000
1!
1*
b10 6
19
1>
1C
b10 G
#18820000000
0!
0*
09
0>
0C
#18830000000
1!
1*
b11 6
19
1>
1C
b11 G
#18840000000
0!
0*
09
0>
0C
#18850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#18860000000
0!
0*
09
0>
0C
#18870000000
1!
1*
b101 6
19
1>
1C
b101 G
#18880000000
0!
0*
09
0>
0C
#18890000000
1!
1*
b110 6
19
1>
1C
b110 G
#18900000000
0!
0*
09
0>
0C
#18910000000
1!
1*
b111 6
19
1>
1C
b111 G
#18920000000
0!
0*
09
0>
0C
#18930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#18940000000
0!
0*
09
0>
0C
#18950000000
1!
1*
b1 6
19
1>
1C
b1 G
#18960000000
0!
0*
09
0>
0C
#18970000000
1!
1*
b10 6
19
1>
1C
b10 G
#18980000000
0!
0*
09
0>
0C
#18990000000
1!
1*
b11 6
19
1>
1C
b11 G
#19000000000
0!
0*
09
0>
0C
#19010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#19020000000
0!
0*
09
0>
0C
#19030000000
1!
1*
b101 6
19
1>
1C
b101 G
#19040000000
0!
0*
09
0>
0C
#19050000000
1!
1*
b110 6
19
1>
1C
b110 G
#19060000000
0!
0*
09
0>
0C
#19070000000
1!
1*
b111 6
19
1>
1C
b111 G
#19080000000
0!
1"
0*
1+
09
1:
0>
0C
#19090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#19100000000
0!
0*
09
0>
0C
#19110000000
1!
1*
b1 6
19
1>
1C
b1 G
#19120000000
0!
0*
09
0>
0C
#19130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#19140000000
0!
0*
09
0>
0C
#19150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#19160000000
0!
0*
09
0>
0C
#19170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#19180000000
0!
0*
09
0>
0C
#19190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#19200000000
0!
0#
0*
0,
09
0>
0?
0C
#19210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#19220000000
0!
0*
09
0>
0C
#19230000000
1!
1*
19
1>
1C
#19240000000
0!
0*
09
0>
0C
#19250000000
1!
1*
19
1>
1C
#19260000000
0!
0*
09
0>
0C
#19270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#19280000000
0!
0*
09
0>
0C
#19290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#19300000000
0!
0*
09
0>
0C
#19310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#19320000000
0!
0*
09
0>
0C
#19330000000
1!
1*
b10 6
19
1>
1C
b10 G
#19340000000
0!
0*
09
0>
0C
#19350000000
1!
1*
b11 6
19
1>
1C
b11 G
#19360000000
0!
0*
09
0>
0C
#19370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#19380000000
0!
0*
09
0>
0C
#19390000000
1!
1*
b101 6
19
1>
1C
b101 G
#19400000000
0!
0*
09
0>
0C
#19410000000
1!
1*
b110 6
19
1>
1C
b110 G
#19420000000
0!
0*
09
0>
0C
#19430000000
1!
1*
b111 6
19
1>
1C
b111 G
#19440000000
0!
0*
09
0>
0C
#19450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#19460000000
0!
0*
09
0>
0C
#19470000000
1!
1*
b1 6
19
1>
1C
b1 G
#19480000000
0!
0*
09
0>
0C
#19490000000
1!
1*
b10 6
19
1>
1C
b10 G
#19500000000
0!
0*
09
0>
0C
#19510000000
1!
1*
b11 6
19
1>
1C
b11 G
#19520000000
0!
0*
09
0>
0C
#19530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#19540000000
0!
0*
09
0>
0C
#19550000000
1!
1*
b101 6
19
1>
1C
b101 G
#19560000000
0!
0*
09
0>
0C
#19570000000
1!
1*
b110 6
19
1>
1C
b110 G
#19580000000
0!
0*
09
0>
0C
#19590000000
1!
1*
b111 6
19
1>
1C
b111 G
#19600000000
0!
0*
09
0>
0C
#19610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#19620000000
0!
0*
09
0>
0C
#19630000000
1!
1*
b1 6
19
1>
1C
b1 G
#19640000000
0!
0*
09
0>
0C
#19650000000
1!
1*
b10 6
19
1>
1C
b10 G
#19660000000
0!
0*
09
0>
0C
#19670000000
1!
1*
b11 6
19
1>
1C
b11 G
#19680000000
0!
0*
09
0>
0C
#19690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#19700000000
0!
0*
09
0>
0C
#19710000000
1!
1*
b101 6
19
1>
1C
b101 G
#19720000000
0!
0*
09
0>
0C
#19730000000
1!
1*
b110 6
19
1>
1C
b110 G
#19740000000
0!
0*
09
0>
0C
#19750000000
1!
1*
b111 6
19
1>
1C
b111 G
#19760000000
0!
1"
0*
1+
09
1:
0>
0C
#19770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#19780000000
0!
0*
09
0>
0C
#19790000000
1!
1*
b1 6
19
1>
1C
b1 G
#19800000000
0!
0*
09
0>
0C
#19810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#19820000000
0!
0*
09
0>
0C
#19830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#19840000000
0!
0*
09
0>
0C
#19850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#19860000000
0!
0*
09
0>
0C
#19870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#19880000000
0!
0#
0*
0,
09
0>
0?
0C
#19890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#19900000000
0!
0*
09
0>
0C
#19910000000
1!
1*
19
1>
1C
#19920000000
0!
0*
09
0>
0C
#19930000000
1!
1*
19
1>
1C
#19940000000
0!
0*
09
0>
0C
#19950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#19960000000
0!
0*
09
0>
0C
#19970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#19980000000
0!
0*
09
0>
0C
#19990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#20000000000
0!
0*
09
0>
0C
#20010000000
1!
1*
b10 6
19
1>
1C
b10 G
#20020000000
0!
0*
09
0>
0C
#20030000000
1!
1*
b11 6
19
1>
1C
b11 G
#20040000000
0!
0*
09
0>
0C
#20050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#20060000000
0!
0*
09
0>
0C
#20070000000
1!
1*
b101 6
19
1>
1C
b101 G
#20080000000
0!
0*
09
0>
0C
#20090000000
1!
1*
b110 6
19
1>
1C
b110 G
#20100000000
0!
0*
09
0>
0C
#20110000000
1!
1*
b111 6
19
1>
1C
b111 G
#20120000000
0!
0*
09
0>
0C
#20130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#20140000000
0!
0*
09
0>
0C
#20150000000
1!
1*
b1 6
19
1>
1C
b1 G
#20160000000
0!
0*
09
0>
0C
#20170000000
1!
1*
b10 6
19
1>
1C
b10 G
#20180000000
0!
0*
09
0>
0C
#20190000000
1!
1*
b11 6
19
1>
1C
b11 G
#20200000000
0!
0*
09
0>
0C
#20210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#20220000000
0!
0*
09
0>
0C
#20230000000
1!
1*
b101 6
19
1>
1C
b101 G
#20240000000
0!
0*
09
0>
0C
#20250000000
1!
1*
b110 6
19
1>
1C
b110 G
#20260000000
0!
0*
09
0>
0C
#20270000000
1!
1*
b111 6
19
1>
1C
b111 G
#20280000000
0!
0*
09
0>
0C
#20290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#20300000000
0!
0*
09
0>
0C
#20310000000
1!
1*
b1 6
19
1>
1C
b1 G
#20320000000
0!
0*
09
0>
0C
#20330000000
1!
1*
b10 6
19
1>
1C
b10 G
#20340000000
0!
0*
09
0>
0C
#20350000000
1!
1*
b11 6
19
1>
1C
b11 G
#20360000000
0!
0*
09
0>
0C
#20370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#20380000000
0!
0*
09
0>
0C
#20390000000
1!
1*
b101 6
19
1>
1C
b101 G
#20400000000
0!
0*
09
0>
0C
#20410000000
1!
1*
b110 6
19
1>
1C
b110 G
#20420000000
0!
0*
09
0>
0C
#20430000000
1!
1*
b111 6
19
1>
1C
b111 G
#20440000000
0!
1"
0*
1+
09
1:
0>
0C
#20450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#20460000000
0!
0*
09
0>
0C
#20470000000
1!
1*
b1 6
19
1>
1C
b1 G
#20480000000
0!
0*
09
0>
0C
#20490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#20500000000
0!
0*
09
0>
0C
#20510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#20520000000
0!
0*
09
0>
0C
#20530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#20540000000
0!
0*
09
0>
0C
#20550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#20560000000
0!
0#
0*
0,
09
0>
0?
0C
#20570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#20580000000
0!
0*
09
0>
0C
#20590000000
1!
1*
19
1>
1C
#20600000000
0!
0*
09
0>
0C
#20610000000
1!
1*
19
1>
1C
#20620000000
0!
0*
09
0>
0C
#20630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#20640000000
0!
0*
09
0>
0C
#20650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#20660000000
0!
0*
09
0>
0C
#20670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#20680000000
0!
0*
09
0>
0C
#20690000000
1!
1*
b10 6
19
1>
1C
b10 G
#20700000000
0!
0*
09
0>
0C
#20710000000
1!
1*
b11 6
19
1>
1C
b11 G
#20720000000
0!
0*
09
0>
0C
#20730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#20740000000
0!
0*
09
0>
0C
#20750000000
1!
1*
b101 6
19
1>
1C
b101 G
#20760000000
0!
0*
09
0>
0C
#20770000000
1!
1*
b110 6
19
1>
1C
b110 G
#20780000000
0!
0*
09
0>
0C
#20790000000
1!
1*
b111 6
19
1>
1C
b111 G
#20800000000
0!
0*
09
0>
0C
#20810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#20820000000
0!
0*
09
0>
0C
#20830000000
1!
1*
b1 6
19
1>
1C
b1 G
#20840000000
0!
0*
09
0>
0C
#20850000000
1!
1*
b10 6
19
1>
1C
b10 G
#20860000000
0!
0*
09
0>
0C
#20870000000
1!
1*
b11 6
19
1>
1C
b11 G
#20880000000
0!
0*
09
0>
0C
#20890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#20900000000
0!
0*
09
0>
0C
#20910000000
1!
1*
b101 6
19
1>
1C
b101 G
#20920000000
0!
0*
09
0>
0C
#20930000000
1!
1*
b110 6
19
1>
1C
b110 G
#20940000000
0!
0*
09
0>
0C
#20950000000
1!
1*
b111 6
19
1>
1C
b111 G
#20960000000
0!
0*
09
0>
0C
#20970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#20980000000
0!
0*
09
0>
0C
#20990000000
1!
1*
b1 6
19
1>
1C
b1 G
#21000000000
0!
0*
09
0>
0C
#21010000000
1!
1*
b10 6
19
1>
1C
b10 G
#21020000000
0!
0*
09
0>
0C
#21030000000
1!
1*
b11 6
19
1>
1C
b11 G
#21040000000
0!
0*
09
0>
0C
#21050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#21060000000
0!
0*
09
0>
0C
#21070000000
1!
1*
b101 6
19
1>
1C
b101 G
#21080000000
0!
0*
09
0>
0C
#21090000000
1!
1*
b110 6
19
1>
1C
b110 G
#21100000000
0!
0*
09
0>
0C
#21110000000
1!
1*
b111 6
19
1>
1C
b111 G
#21120000000
0!
1"
0*
1+
09
1:
0>
0C
#21130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#21140000000
0!
0*
09
0>
0C
#21150000000
1!
1*
b1 6
19
1>
1C
b1 G
#21160000000
0!
0*
09
0>
0C
#21170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#21180000000
0!
0*
09
0>
0C
#21190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#21200000000
0!
0*
09
0>
0C
#21210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#21220000000
0!
0*
09
0>
0C
#21230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#21240000000
0!
0#
0*
0,
09
0>
0?
0C
#21250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#21260000000
0!
0*
09
0>
0C
#21270000000
1!
1*
19
1>
1C
#21280000000
0!
0*
09
0>
0C
#21290000000
1!
1*
19
1>
1C
#21300000000
0!
0*
09
0>
0C
#21310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#21320000000
0!
0*
09
0>
0C
#21330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#21340000000
0!
0*
09
0>
0C
#21350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#21360000000
0!
0*
09
0>
0C
#21370000000
1!
1*
b10 6
19
1>
1C
b10 G
#21380000000
0!
0*
09
0>
0C
#21390000000
1!
1*
b11 6
19
1>
1C
b11 G
#21400000000
0!
0*
09
0>
0C
#21410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#21420000000
0!
0*
09
0>
0C
#21430000000
1!
1*
b101 6
19
1>
1C
b101 G
#21440000000
0!
0*
09
0>
0C
#21450000000
1!
1*
b110 6
19
1>
1C
b110 G
#21460000000
0!
0*
09
0>
0C
#21470000000
1!
1*
b111 6
19
1>
1C
b111 G
#21480000000
0!
0*
09
0>
0C
#21490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#21500000000
0!
0*
09
0>
0C
#21510000000
1!
1*
b1 6
19
1>
1C
b1 G
#21520000000
0!
0*
09
0>
0C
#21530000000
1!
1*
b10 6
19
1>
1C
b10 G
#21540000000
0!
0*
09
0>
0C
#21550000000
1!
1*
b11 6
19
1>
1C
b11 G
#21560000000
0!
0*
09
0>
0C
#21570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#21580000000
0!
0*
09
0>
0C
#21590000000
1!
1*
b101 6
19
1>
1C
b101 G
#21600000000
0!
0*
09
0>
0C
#21610000000
1!
1*
b110 6
19
1>
1C
b110 G
#21620000000
0!
0*
09
0>
0C
#21630000000
1!
1*
b111 6
19
1>
1C
b111 G
#21640000000
0!
0*
09
0>
0C
#21650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#21660000000
0!
0*
09
0>
0C
#21670000000
1!
1*
b1 6
19
1>
1C
b1 G
#21680000000
0!
0*
09
0>
0C
#21690000000
1!
1*
b10 6
19
1>
1C
b10 G
#21700000000
0!
0*
09
0>
0C
#21710000000
1!
1*
b11 6
19
1>
1C
b11 G
#21720000000
0!
0*
09
0>
0C
#21730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#21740000000
0!
0*
09
0>
0C
#21750000000
1!
1*
b101 6
19
1>
1C
b101 G
#21760000000
0!
0*
09
0>
0C
#21770000000
1!
1*
b110 6
19
1>
1C
b110 G
#21780000000
0!
0*
09
0>
0C
#21790000000
1!
1*
b111 6
19
1>
1C
b111 G
#21800000000
0!
1"
0*
1+
09
1:
0>
0C
#21810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#21820000000
0!
0*
09
0>
0C
#21830000000
1!
1*
b1 6
19
1>
1C
b1 G
#21840000000
0!
0*
09
0>
0C
#21850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#21860000000
0!
0*
09
0>
0C
#21870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#21880000000
0!
0*
09
0>
0C
#21890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#21900000000
0!
0*
09
0>
0C
#21910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#21920000000
0!
0#
0*
0,
09
0>
0?
0C
#21930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#21940000000
0!
0*
09
0>
0C
#21950000000
1!
1*
19
1>
1C
#21960000000
0!
0*
09
0>
0C
#21970000000
1!
1*
19
1>
1C
#21980000000
0!
0*
09
0>
0C
#21990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#22000000000
0!
0*
09
0>
0C
#22010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#22020000000
0!
0*
09
0>
0C
#22030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#22040000000
0!
0*
09
0>
0C
#22050000000
1!
1*
b10 6
19
1>
1C
b10 G
#22060000000
0!
0*
09
0>
0C
#22070000000
1!
1*
b11 6
19
1>
1C
b11 G
#22080000000
0!
0*
09
0>
0C
#22090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#22100000000
0!
0*
09
0>
0C
#22110000000
1!
1*
b101 6
19
1>
1C
b101 G
#22120000000
0!
0*
09
0>
0C
#22130000000
1!
1*
b110 6
19
1>
1C
b110 G
#22140000000
0!
0*
09
0>
0C
#22150000000
1!
1*
b111 6
19
1>
1C
b111 G
#22160000000
0!
0*
09
0>
0C
#22170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#22180000000
0!
0*
09
0>
0C
#22190000000
1!
1*
b1 6
19
1>
1C
b1 G
#22200000000
0!
0*
09
0>
0C
#22210000000
1!
1*
b10 6
19
1>
1C
b10 G
#22220000000
0!
0*
09
0>
0C
#22230000000
1!
1*
b11 6
19
1>
1C
b11 G
#22240000000
0!
0*
09
0>
0C
#22250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#22260000000
0!
0*
09
0>
0C
#22270000000
1!
1*
b101 6
19
1>
1C
b101 G
#22280000000
0!
0*
09
0>
0C
#22290000000
1!
1*
b110 6
19
1>
1C
b110 G
#22300000000
0!
0*
09
0>
0C
#22310000000
1!
1*
b111 6
19
1>
1C
b111 G
#22320000000
0!
0*
09
0>
0C
#22330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#22340000000
0!
0*
09
0>
0C
#22350000000
1!
1*
b1 6
19
1>
1C
b1 G
#22360000000
0!
0*
09
0>
0C
#22370000000
1!
1*
b10 6
19
1>
1C
b10 G
#22380000000
0!
0*
09
0>
0C
#22390000000
1!
1*
b11 6
19
1>
1C
b11 G
#22400000000
0!
0*
09
0>
0C
#22410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#22420000000
0!
0*
09
0>
0C
#22430000000
1!
1*
b101 6
19
1>
1C
b101 G
#22440000000
0!
0*
09
0>
0C
#22450000000
1!
1*
b110 6
19
1>
1C
b110 G
#22460000000
0!
0*
09
0>
0C
#22470000000
1!
1*
b111 6
19
1>
1C
b111 G
#22480000000
0!
1"
0*
1+
09
1:
0>
0C
#22490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#22500000000
0!
0*
09
0>
0C
#22510000000
1!
1*
b1 6
19
1>
1C
b1 G
#22520000000
0!
0*
09
0>
0C
#22530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#22540000000
0!
0*
09
0>
0C
#22550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#22560000000
0!
0*
09
0>
0C
#22570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#22580000000
0!
0*
09
0>
0C
#22590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#22600000000
0!
0#
0*
0,
09
0>
0?
0C
#22610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#22620000000
0!
0*
09
0>
0C
#22630000000
1!
1*
19
1>
1C
#22640000000
0!
0*
09
0>
0C
#22650000000
1!
1*
19
1>
1C
#22660000000
0!
0*
09
0>
0C
#22670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#22680000000
0!
0*
09
0>
0C
#22690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#22700000000
0!
0*
09
0>
0C
#22710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#22720000000
0!
0*
09
0>
0C
#22730000000
1!
1*
b10 6
19
1>
1C
b10 G
#22740000000
0!
0*
09
0>
0C
#22750000000
1!
1*
b11 6
19
1>
1C
b11 G
#22760000000
0!
0*
09
0>
0C
#22770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#22780000000
0!
0*
09
0>
0C
#22790000000
1!
1*
b101 6
19
1>
1C
b101 G
#22800000000
0!
0*
09
0>
0C
#22810000000
1!
1*
b110 6
19
1>
1C
b110 G
#22820000000
0!
0*
09
0>
0C
#22830000000
1!
1*
b111 6
19
1>
1C
b111 G
#22840000000
0!
0*
09
0>
0C
#22850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#22860000000
0!
0*
09
0>
0C
#22870000000
1!
1*
b1 6
19
1>
1C
b1 G
#22880000000
0!
0*
09
0>
0C
#22890000000
1!
1*
b10 6
19
1>
1C
b10 G
#22900000000
0!
0*
09
0>
0C
#22910000000
1!
1*
b11 6
19
1>
1C
b11 G
#22920000000
0!
0*
09
0>
0C
#22930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#22940000000
0!
0*
09
0>
0C
#22950000000
1!
1*
b101 6
19
1>
1C
b101 G
#22960000000
0!
0*
09
0>
0C
#22970000000
1!
1*
b110 6
19
1>
1C
b110 G
#22980000000
0!
0*
09
0>
0C
#22990000000
1!
1*
b111 6
19
1>
1C
b111 G
#23000000000
0!
0*
09
0>
0C
#23010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#23020000000
0!
0*
09
0>
0C
#23030000000
1!
1*
b1 6
19
1>
1C
b1 G
#23040000000
0!
0*
09
0>
0C
#23050000000
1!
1*
b10 6
19
1>
1C
b10 G
#23060000000
0!
0*
09
0>
0C
#23070000000
1!
1*
b11 6
19
1>
1C
b11 G
#23080000000
0!
0*
09
0>
0C
#23090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#23100000000
0!
0*
09
0>
0C
#23110000000
1!
1*
b101 6
19
1>
1C
b101 G
#23120000000
0!
0*
09
0>
0C
#23130000000
1!
1*
b110 6
19
1>
1C
b110 G
#23140000000
0!
0*
09
0>
0C
#23150000000
1!
1*
b111 6
19
1>
1C
b111 G
#23160000000
0!
1"
0*
1+
09
1:
0>
0C
#23170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#23180000000
0!
0*
09
0>
0C
#23190000000
1!
1*
b1 6
19
1>
1C
b1 G
#23200000000
0!
0*
09
0>
0C
#23210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#23220000000
0!
0*
09
0>
0C
#23230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#23240000000
0!
0*
09
0>
0C
#23250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#23260000000
0!
0*
09
0>
0C
#23270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#23280000000
0!
0#
0*
0,
09
0>
0?
0C
#23290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#23300000000
0!
0*
09
0>
0C
#23310000000
1!
1*
19
1>
1C
#23320000000
0!
0*
09
0>
0C
#23330000000
1!
1*
19
1>
1C
#23340000000
0!
0*
09
0>
0C
#23350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#23360000000
0!
0*
09
0>
0C
#23370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#23380000000
0!
0*
09
0>
0C
#23390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#23400000000
0!
0*
09
0>
0C
#23410000000
1!
1*
b10 6
19
1>
1C
b10 G
#23420000000
0!
0*
09
0>
0C
#23430000000
1!
1*
b11 6
19
1>
1C
b11 G
#23440000000
0!
0*
09
0>
0C
#23450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#23460000000
0!
0*
09
0>
0C
#23470000000
1!
1*
b101 6
19
1>
1C
b101 G
#23480000000
0!
0*
09
0>
0C
#23490000000
1!
1*
b110 6
19
1>
1C
b110 G
#23500000000
0!
0*
09
0>
0C
#23510000000
1!
1*
b111 6
19
1>
1C
b111 G
#23520000000
0!
0*
09
0>
0C
#23530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#23540000000
0!
0*
09
0>
0C
#23550000000
1!
1*
b1 6
19
1>
1C
b1 G
#23560000000
0!
0*
09
0>
0C
#23570000000
1!
1*
b10 6
19
1>
1C
b10 G
#23580000000
0!
0*
09
0>
0C
#23590000000
1!
1*
b11 6
19
1>
1C
b11 G
#23600000000
0!
0*
09
0>
0C
#23610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#23620000000
0!
0*
09
0>
0C
#23630000000
1!
1*
b101 6
19
1>
1C
b101 G
#23640000000
0!
0*
09
0>
0C
#23650000000
1!
1*
b110 6
19
1>
1C
b110 G
#23660000000
0!
0*
09
0>
0C
#23670000000
1!
1*
b111 6
19
1>
1C
b111 G
#23680000000
0!
0*
09
0>
0C
#23690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#23700000000
0!
0*
09
0>
0C
#23710000000
1!
1*
b1 6
19
1>
1C
b1 G
#23720000000
0!
0*
09
0>
0C
#23730000000
1!
1*
b10 6
19
1>
1C
b10 G
#23740000000
0!
0*
09
0>
0C
#23750000000
1!
1*
b11 6
19
1>
1C
b11 G
#23760000000
0!
0*
09
0>
0C
#23770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#23780000000
0!
0*
09
0>
0C
#23790000000
1!
1*
b101 6
19
1>
1C
b101 G
#23800000000
0!
0*
09
0>
0C
#23810000000
1!
1*
b110 6
19
1>
1C
b110 G
#23820000000
0!
0*
09
0>
0C
#23830000000
1!
1*
b111 6
19
1>
1C
b111 G
#23840000000
0!
1"
0*
1+
09
1:
0>
0C
#23850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#23860000000
0!
0*
09
0>
0C
#23870000000
1!
1*
b1 6
19
1>
1C
b1 G
#23880000000
0!
0*
09
0>
0C
#23890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#23900000000
0!
0*
09
0>
0C
#23910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#23920000000
0!
0*
09
0>
0C
#23930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#23940000000
0!
0*
09
0>
0C
#23950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#23960000000
0!
0#
0*
0,
09
0>
0?
0C
#23970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#23980000000
0!
0*
09
0>
0C
#23990000000
1!
1*
19
1>
1C
#24000000000
0!
0*
09
0>
0C
#24010000000
1!
1*
19
1>
1C
#24020000000
0!
0*
09
0>
0C
#24030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#24040000000
0!
0*
09
0>
0C
#24050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#24060000000
0!
0*
09
0>
0C
#24070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#24080000000
0!
0*
09
0>
0C
#24090000000
1!
1*
b10 6
19
1>
1C
b10 G
#24100000000
0!
0*
09
0>
0C
#24110000000
1!
1*
b11 6
19
1>
1C
b11 G
#24120000000
0!
0*
09
0>
0C
#24130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#24140000000
0!
0*
09
0>
0C
#24150000000
1!
1*
b101 6
19
1>
1C
b101 G
#24160000000
0!
0*
09
0>
0C
#24170000000
1!
1*
b110 6
19
1>
1C
b110 G
#24180000000
0!
0*
09
0>
0C
#24190000000
1!
1*
b111 6
19
1>
1C
b111 G
#24200000000
0!
0*
09
0>
0C
#24210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#24220000000
0!
0*
09
0>
0C
#24230000000
1!
1*
b1 6
19
1>
1C
b1 G
#24240000000
0!
0*
09
0>
0C
#24250000000
1!
1*
b10 6
19
1>
1C
b10 G
#24260000000
0!
0*
09
0>
0C
#24270000000
1!
1*
b11 6
19
1>
1C
b11 G
#24280000000
0!
0*
09
0>
0C
#24290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#24300000000
0!
0*
09
0>
0C
#24310000000
1!
1*
b101 6
19
1>
1C
b101 G
#24320000000
0!
0*
09
0>
0C
#24330000000
1!
1*
b110 6
19
1>
1C
b110 G
#24340000000
0!
0*
09
0>
0C
#24350000000
1!
1*
b111 6
19
1>
1C
b111 G
#24360000000
0!
0*
09
0>
0C
#24370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#24380000000
0!
0*
09
0>
0C
#24390000000
1!
1*
b1 6
19
1>
1C
b1 G
#24400000000
0!
0*
09
0>
0C
#24410000000
1!
1*
b10 6
19
1>
1C
b10 G
#24420000000
0!
0*
09
0>
0C
#24430000000
1!
1*
b11 6
19
1>
1C
b11 G
#24440000000
0!
0*
09
0>
0C
#24450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#24460000000
0!
0*
09
0>
0C
#24470000000
1!
1*
b101 6
19
1>
1C
b101 G
#24480000000
0!
0*
09
0>
0C
#24490000000
1!
1*
b110 6
19
1>
1C
b110 G
#24500000000
0!
0*
09
0>
0C
#24510000000
1!
1*
b111 6
19
1>
1C
b111 G
#24520000000
0!
1"
0*
1+
09
1:
0>
0C
#24530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#24540000000
0!
0*
09
0>
0C
#24550000000
1!
1*
b1 6
19
1>
1C
b1 G
#24560000000
0!
0*
09
0>
0C
#24570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#24580000000
0!
0*
09
0>
0C
#24590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#24600000000
0!
0*
09
0>
0C
#24610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#24620000000
0!
0*
09
0>
0C
#24630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#24640000000
0!
0#
0*
0,
09
0>
0?
0C
#24650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#24660000000
0!
0*
09
0>
0C
#24670000000
1!
1*
19
1>
1C
#24680000000
0!
0*
09
0>
0C
#24690000000
1!
1*
19
1>
1C
#24700000000
0!
0*
09
0>
0C
#24710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#24720000000
0!
0*
09
0>
0C
#24730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#24740000000
0!
0*
09
0>
0C
#24750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#24760000000
0!
0*
09
0>
0C
#24770000000
1!
1*
b10 6
19
1>
1C
b10 G
#24780000000
0!
0*
09
0>
0C
#24790000000
1!
1*
b11 6
19
1>
1C
b11 G
#24800000000
0!
0*
09
0>
0C
#24810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#24820000000
0!
0*
09
0>
0C
#24830000000
1!
1*
b101 6
19
1>
1C
b101 G
#24840000000
0!
0*
09
0>
0C
#24850000000
1!
1*
b110 6
19
1>
1C
b110 G
#24860000000
0!
0*
09
0>
0C
#24870000000
1!
1*
b111 6
19
1>
1C
b111 G
#24880000000
0!
0*
09
0>
0C
#24890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#24900000000
0!
0*
09
0>
0C
#24910000000
1!
1*
b1 6
19
1>
1C
b1 G
#24920000000
0!
0*
09
0>
0C
#24930000000
1!
1*
b10 6
19
1>
1C
b10 G
#24940000000
0!
0*
09
0>
0C
#24950000000
1!
1*
b11 6
19
1>
1C
b11 G
#24960000000
0!
0*
09
0>
0C
#24970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#24980000000
0!
0*
09
0>
0C
#24990000000
1!
1*
b101 6
19
1>
1C
b101 G
#25000000000
0!
0*
09
0>
0C
#25010000000
1!
1*
b110 6
19
1>
1C
b110 G
#25020000000
0!
0*
09
0>
0C
#25030000000
1!
1*
b111 6
19
1>
1C
b111 G
#25040000000
0!
0*
09
0>
0C
#25050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#25060000000
0!
0*
09
0>
0C
#25070000000
1!
1*
b1 6
19
1>
1C
b1 G
#25080000000
0!
0*
09
0>
0C
#25090000000
1!
1*
b10 6
19
1>
1C
b10 G
#25100000000
0!
0*
09
0>
0C
#25110000000
1!
1*
b11 6
19
1>
1C
b11 G
#25120000000
0!
0*
09
0>
0C
#25130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#25140000000
0!
0*
09
0>
0C
#25150000000
1!
1*
b101 6
19
1>
1C
b101 G
#25160000000
0!
0*
09
0>
0C
#25170000000
1!
1*
b110 6
19
1>
1C
b110 G
#25180000000
0!
0*
09
0>
0C
#25190000000
1!
1*
b111 6
19
1>
1C
b111 G
#25200000000
0!
1"
0*
1+
09
1:
0>
0C
#25210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#25220000000
0!
0*
09
0>
0C
#25230000000
1!
1*
b1 6
19
1>
1C
b1 G
#25240000000
0!
0*
09
0>
0C
#25250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#25260000000
0!
0*
09
0>
0C
#25270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#25280000000
0!
0*
09
0>
0C
#25290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#25300000000
0!
0*
09
0>
0C
#25310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#25320000000
0!
0#
0*
0,
09
0>
0?
0C
#25330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#25340000000
0!
0*
09
0>
0C
#25350000000
1!
1*
19
1>
1C
#25360000000
0!
0*
09
0>
0C
#25370000000
1!
1*
19
1>
1C
#25380000000
0!
0*
09
0>
0C
#25390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#25400000000
0!
0*
09
0>
0C
#25410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#25420000000
0!
0*
09
0>
0C
#25430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#25440000000
0!
0*
09
0>
0C
#25450000000
1!
1*
b10 6
19
1>
1C
b10 G
#25460000000
0!
0*
09
0>
0C
#25470000000
1!
1*
b11 6
19
1>
1C
b11 G
#25480000000
0!
0*
09
0>
0C
#25490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#25500000000
0!
0*
09
0>
0C
#25510000000
1!
1*
b101 6
19
1>
1C
b101 G
#25520000000
0!
0*
09
0>
0C
#25530000000
1!
1*
b110 6
19
1>
1C
b110 G
#25540000000
0!
0*
09
0>
0C
#25550000000
1!
1*
b111 6
19
1>
1C
b111 G
#25560000000
0!
0*
09
0>
0C
#25570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#25580000000
0!
0*
09
0>
0C
#25590000000
1!
1*
b1 6
19
1>
1C
b1 G
#25600000000
0!
0*
09
0>
0C
#25610000000
1!
1*
b10 6
19
1>
1C
b10 G
#25620000000
0!
0*
09
0>
0C
#25630000000
1!
1*
b11 6
19
1>
1C
b11 G
#25640000000
0!
0*
09
0>
0C
#25650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#25660000000
0!
0*
09
0>
0C
#25670000000
1!
1*
b101 6
19
1>
1C
b101 G
#25680000000
0!
0*
09
0>
0C
#25690000000
1!
1*
b110 6
19
1>
1C
b110 G
#25700000000
0!
0*
09
0>
0C
#25710000000
1!
1*
b111 6
19
1>
1C
b111 G
#25720000000
0!
0*
09
0>
0C
#25730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#25740000000
0!
0*
09
0>
0C
#25750000000
1!
1*
b1 6
19
1>
1C
b1 G
#25760000000
0!
0*
09
0>
0C
#25770000000
1!
1*
b10 6
19
1>
1C
b10 G
#25780000000
0!
0*
09
0>
0C
#25790000000
1!
1*
b11 6
19
1>
1C
b11 G
#25800000000
0!
0*
09
0>
0C
#25810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#25820000000
0!
0*
09
0>
0C
#25830000000
1!
1*
b101 6
19
1>
1C
b101 G
#25840000000
0!
0*
09
0>
0C
#25850000000
1!
1*
b110 6
19
1>
1C
b110 G
#25860000000
0!
0*
09
0>
0C
#25870000000
1!
1*
b111 6
19
1>
1C
b111 G
#25880000000
0!
1"
0*
1+
09
1:
0>
0C
#25890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#25900000000
0!
0*
09
0>
0C
#25910000000
1!
1*
b1 6
19
1>
1C
b1 G
#25920000000
0!
0*
09
0>
0C
#25930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#25940000000
0!
0*
09
0>
0C
#25950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#25960000000
0!
0*
09
0>
0C
#25970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#25980000000
0!
0*
09
0>
0C
#25990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#26000000000
0!
0#
0*
0,
09
0>
0?
0C
#26010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#26020000000
0!
0*
09
0>
0C
#26030000000
1!
1*
19
1>
1C
#26040000000
0!
0*
09
0>
0C
#26050000000
1!
1*
19
1>
1C
#26060000000
0!
0*
09
0>
0C
#26070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#26080000000
0!
0*
09
0>
0C
#26090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#26100000000
0!
0*
09
0>
0C
#26110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#26120000000
0!
0*
09
0>
0C
#26130000000
1!
1*
b10 6
19
1>
1C
b10 G
#26140000000
0!
0*
09
0>
0C
#26150000000
1!
1*
b11 6
19
1>
1C
b11 G
#26160000000
0!
0*
09
0>
0C
#26170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#26180000000
0!
0*
09
0>
0C
#26190000000
1!
1*
b101 6
19
1>
1C
b101 G
#26200000000
0!
0*
09
0>
0C
#26210000000
1!
1*
b110 6
19
1>
1C
b110 G
#26220000000
0!
0*
09
0>
0C
#26230000000
1!
1*
b111 6
19
1>
1C
b111 G
#26240000000
0!
0*
09
0>
0C
#26250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#26260000000
0!
0*
09
0>
0C
#26270000000
1!
1*
b1 6
19
1>
1C
b1 G
#26280000000
0!
0*
09
0>
0C
#26290000000
1!
1*
b10 6
19
1>
1C
b10 G
#26300000000
0!
0*
09
0>
0C
#26310000000
1!
1*
b11 6
19
1>
1C
b11 G
#26320000000
0!
0*
09
0>
0C
#26330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#26340000000
0!
0*
09
0>
0C
#26350000000
1!
1*
b101 6
19
1>
1C
b101 G
#26360000000
0!
0*
09
0>
0C
#26370000000
1!
1*
b110 6
19
1>
1C
b110 G
#26380000000
0!
0*
09
0>
0C
#26390000000
1!
1*
b111 6
19
1>
1C
b111 G
#26400000000
0!
0*
09
0>
0C
#26410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#26420000000
0!
0*
09
0>
0C
#26430000000
1!
1*
b1 6
19
1>
1C
b1 G
#26440000000
0!
0*
09
0>
0C
#26450000000
1!
1*
b10 6
19
1>
1C
b10 G
#26460000000
0!
0*
09
0>
0C
#26470000000
1!
1*
b11 6
19
1>
1C
b11 G
#26480000000
0!
0*
09
0>
0C
#26490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#26500000000
0!
0*
09
0>
0C
#26510000000
1!
1*
b101 6
19
1>
1C
b101 G
#26520000000
0!
0*
09
0>
0C
#26530000000
1!
1*
b110 6
19
1>
1C
b110 G
#26540000000
0!
0*
09
0>
0C
#26550000000
1!
1*
b111 6
19
1>
1C
b111 G
#26560000000
0!
1"
0*
1+
09
1:
0>
0C
#26570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#26580000000
0!
0*
09
0>
0C
#26590000000
1!
1*
b1 6
19
1>
1C
b1 G
#26600000000
0!
0*
09
0>
0C
#26610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#26620000000
0!
0*
09
0>
0C
#26630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#26640000000
0!
0*
09
0>
0C
#26650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#26660000000
0!
0*
09
0>
0C
#26670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#26680000000
0!
0#
0*
0,
09
0>
0?
0C
#26690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#26700000000
0!
0*
09
0>
0C
#26710000000
1!
1*
19
1>
1C
#26720000000
0!
0*
09
0>
0C
#26730000000
1!
1*
19
1>
1C
#26740000000
0!
0*
09
0>
0C
#26750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#26760000000
0!
0*
09
0>
0C
#26770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#26780000000
0!
0*
09
0>
0C
#26790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#26800000000
0!
0*
09
0>
0C
#26810000000
1!
1*
b10 6
19
1>
1C
b10 G
#26820000000
0!
0*
09
0>
0C
#26830000000
1!
1*
b11 6
19
1>
1C
b11 G
#26840000000
0!
0*
09
0>
0C
#26850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#26860000000
0!
0*
09
0>
0C
#26870000000
1!
1*
b101 6
19
1>
1C
b101 G
#26880000000
0!
0*
09
0>
0C
#26890000000
1!
1*
b110 6
19
1>
1C
b110 G
#26900000000
0!
0*
09
0>
0C
#26910000000
1!
1*
b111 6
19
1>
1C
b111 G
#26920000000
0!
0*
09
0>
0C
#26930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#26940000000
0!
0*
09
0>
0C
#26950000000
1!
1*
b1 6
19
1>
1C
b1 G
#26960000000
0!
0*
09
0>
0C
#26970000000
1!
1*
b10 6
19
1>
1C
b10 G
#26980000000
0!
0*
09
0>
0C
#26990000000
1!
1*
b11 6
19
1>
1C
b11 G
#27000000000
0!
0*
09
0>
0C
#27010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#27020000000
0!
0*
09
0>
0C
#27030000000
1!
1*
b101 6
19
1>
1C
b101 G
#27040000000
0!
0*
09
0>
0C
#27050000000
1!
1*
b110 6
19
1>
1C
b110 G
#27060000000
0!
0*
09
0>
0C
#27070000000
1!
1*
b111 6
19
1>
1C
b111 G
#27080000000
0!
0*
09
0>
0C
#27090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#27100000000
0!
0*
09
0>
0C
#27110000000
1!
1*
b1 6
19
1>
1C
b1 G
#27120000000
0!
0*
09
0>
0C
#27130000000
1!
1*
b10 6
19
1>
1C
b10 G
#27140000000
0!
0*
09
0>
0C
#27150000000
1!
1*
b11 6
19
1>
1C
b11 G
#27160000000
0!
0*
09
0>
0C
#27170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#27180000000
0!
0*
09
0>
0C
#27190000000
1!
1*
b101 6
19
1>
1C
b101 G
#27200000000
0!
0*
09
0>
0C
#27210000000
1!
1*
b110 6
19
1>
1C
b110 G
#27220000000
0!
0*
09
0>
0C
#27230000000
1!
1*
b111 6
19
1>
1C
b111 G
#27240000000
0!
1"
0*
1+
09
1:
0>
0C
#27250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#27260000000
0!
0*
09
0>
0C
#27270000000
1!
1*
b1 6
19
1>
1C
b1 G
#27280000000
0!
0*
09
0>
0C
#27290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#27300000000
0!
0*
09
0>
0C
#27310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#27320000000
0!
0*
09
0>
0C
#27330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#27340000000
0!
0*
09
0>
0C
#27350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#27360000000
0!
0#
0*
0,
09
0>
0?
0C
#27370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#27380000000
0!
0*
09
0>
0C
#27390000000
1!
1*
19
1>
1C
#27400000000
0!
0*
09
0>
0C
#27410000000
1!
1*
19
1>
1C
#27420000000
0!
0*
09
0>
0C
#27430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#27440000000
0!
0*
09
0>
0C
#27450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#27460000000
0!
0*
09
0>
0C
#27470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#27480000000
0!
0*
09
0>
0C
#27490000000
1!
1*
b10 6
19
1>
1C
b10 G
#27500000000
0!
0*
09
0>
0C
#27510000000
1!
1*
b11 6
19
1>
1C
b11 G
#27520000000
0!
0*
09
0>
0C
#27530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#27540000000
0!
0*
09
0>
0C
#27550000000
1!
1*
b101 6
19
1>
1C
b101 G
#27560000000
0!
0*
09
0>
0C
#27570000000
1!
1*
b110 6
19
1>
1C
b110 G
#27580000000
0!
0*
09
0>
0C
#27590000000
1!
1*
b111 6
19
1>
1C
b111 G
#27600000000
0!
0*
09
0>
0C
#27610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#27620000000
0!
0*
09
0>
0C
#27630000000
1!
1*
b1 6
19
1>
1C
b1 G
#27640000000
0!
0*
09
0>
0C
#27650000000
1!
1*
b10 6
19
1>
1C
b10 G
#27660000000
0!
0*
09
0>
0C
#27670000000
1!
1*
b11 6
19
1>
1C
b11 G
#27680000000
0!
0*
09
0>
0C
#27690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#27700000000
0!
0*
09
0>
0C
#27710000000
1!
1*
b101 6
19
1>
1C
b101 G
#27720000000
0!
0*
09
0>
0C
#27730000000
1!
1*
b110 6
19
1>
1C
b110 G
#27740000000
0!
0*
09
0>
0C
#27750000000
1!
1*
b111 6
19
1>
1C
b111 G
#27760000000
0!
0*
09
0>
0C
#27770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#27780000000
0!
0*
09
0>
0C
#27790000000
1!
1*
b1 6
19
1>
1C
b1 G
#27800000000
0!
0*
09
0>
0C
#27810000000
1!
1*
b10 6
19
1>
1C
b10 G
#27820000000
0!
0*
09
0>
0C
#27830000000
1!
1*
b11 6
19
1>
1C
b11 G
#27840000000
0!
0*
09
0>
0C
#27850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#27860000000
0!
0*
09
0>
0C
#27870000000
1!
1*
b101 6
19
1>
1C
b101 G
#27880000000
0!
0*
09
0>
0C
#27890000000
1!
1*
b110 6
19
1>
1C
b110 G
#27900000000
0!
0*
09
0>
0C
#27910000000
1!
1*
b111 6
19
1>
1C
b111 G
#27920000000
0!
1"
0*
1+
09
1:
0>
0C
#27930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#27940000000
0!
0*
09
0>
0C
#27950000000
1!
1*
b1 6
19
1>
1C
b1 G
#27960000000
0!
0*
09
0>
0C
#27970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#27980000000
0!
0*
09
0>
0C
#27990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#28000000000
0!
0*
09
0>
0C
#28010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#28020000000
0!
0*
09
0>
0C
#28030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#28040000000
0!
0#
0*
0,
09
0>
0?
0C
#28050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#28060000000
0!
0*
09
0>
0C
#28070000000
1!
1*
19
1>
1C
#28080000000
0!
0*
09
0>
0C
#28090000000
1!
1*
19
1>
1C
#28100000000
0!
0*
09
0>
0C
#28110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#28120000000
0!
0*
09
0>
0C
#28130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#28140000000
0!
0*
09
0>
0C
#28150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#28160000000
0!
0*
09
0>
0C
#28170000000
1!
1*
b10 6
19
1>
1C
b10 G
#28180000000
0!
0*
09
0>
0C
#28190000000
1!
1*
b11 6
19
1>
1C
b11 G
#28200000000
0!
0*
09
0>
0C
#28210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#28220000000
0!
0*
09
0>
0C
#28230000000
1!
1*
b101 6
19
1>
1C
b101 G
#28240000000
0!
0*
09
0>
0C
#28250000000
1!
1*
b110 6
19
1>
1C
b110 G
#28260000000
0!
0*
09
0>
0C
#28270000000
1!
1*
b111 6
19
1>
1C
b111 G
#28280000000
0!
0*
09
0>
0C
#28290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#28300000000
0!
0*
09
0>
0C
#28310000000
1!
1*
b1 6
19
1>
1C
b1 G
#28320000000
0!
0*
09
0>
0C
#28330000000
1!
1*
b10 6
19
1>
1C
b10 G
#28340000000
0!
0*
09
0>
0C
#28350000000
1!
1*
b11 6
19
1>
1C
b11 G
#28360000000
0!
0*
09
0>
0C
#28370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#28380000000
0!
0*
09
0>
0C
#28390000000
1!
1*
b101 6
19
1>
1C
b101 G
#28400000000
0!
0*
09
0>
0C
#28410000000
1!
1*
b110 6
19
1>
1C
b110 G
#28420000000
0!
0*
09
0>
0C
#28430000000
1!
1*
b111 6
19
1>
1C
b111 G
#28440000000
0!
0*
09
0>
0C
#28450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#28460000000
0!
0*
09
0>
0C
#28470000000
1!
1*
b1 6
19
1>
1C
b1 G
#28480000000
0!
0*
09
0>
0C
#28490000000
1!
1*
b10 6
19
1>
1C
b10 G
#28500000000
0!
0*
09
0>
0C
#28510000000
1!
1*
b11 6
19
1>
1C
b11 G
#28520000000
0!
0*
09
0>
0C
#28530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#28540000000
0!
0*
09
0>
0C
#28550000000
1!
1*
b101 6
19
1>
1C
b101 G
#28560000000
0!
0*
09
0>
0C
#28570000000
1!
1*
b110 6
19
1>
1C
b110 G
#28580000000
0!
0*
09
0>
0C
#28590000000
1!
1*
b111 6
19
1>
1C
b111 G
#28600000000
0!
1"
0*
1+
09
1:
0>
0C
#28610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#28620000000
0!
0*
09
0>
0C
#28630000000
1!
1*
b1 6
19
1>
1C
b1 G
#28640000000
0!
0*
09
0>
0C
#28650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#28660000000
0!
0*
09
0>
0C
#28670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#28680000000
0!
0*
09
0>
0C
#28690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#28700000000
0!
0*
09
0>
0C
#28710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#28720000000
0!
0#
0*
0,
09
0>
0?
0C
#28730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#28740000000
0!
0*
09
0>
0C
#28750000000
1!
1*
19
1>
1C
#28760000000
0!
0*
09
0>
0C
#28770000000
1!
1*
19
1>
1C
#28780000000
0!
0*
09
0>
0C
#28790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#28800000000
0!
0*
09
0>
0C
#28810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#28820000000
0!
0*
09
0>
0C
#28830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#28840000000
0!
0*
09
0>
0C
#28850000000
1!
1*
b10 6
19
1>
1C
b10 G
#28860000000
0!
0*
09
0>
0C
#28870000000
1!
1*
b11 6
19
1>
1C
b11 G
#28880000000
0!
0*
09
0>
0C
#28890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#28900000000
0!
0*
09
0>
0C
#28910000000
1!
1*
b101 6
19
1>
1C
b101 G
#28920000000
0!
0*
09
0>
0C
#28930000000
1!
1*
b110 6
19
1>
1C
b110 G
#28940000000
0!
0*
09
0>
0C
#28950000000
1!
1*
b111 6
19
1>
1C
b111 G
#28960000000
0!
0*
09
0>
0C
#28970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#28980000000
0!
0*
09
0>
0C
#28990000000
1!
1*
b1 6
19
1>
1C
b1 G
#29000000000
0!
0*
09
0>
0C
#29010000000
1!
1*
b10 6
19
1>
1C
b10 G
#29020000000
0!
0*
09
0>
0C
#29030000000
1!
1*
b11 6
19
1>
1C
b11 G
#29040000000
0!
0*
09
0>
0C
#29050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#29060000000
0!
0*
09
0>
0C
#29070000000
1!
1*
b101 6
19
1>
1C
b101 G
#29080000000
0!
0*
09
0>
0C
#29090000000
1!
1*
b110 6
19
1>
1C
b110 G
#29100000000
0!
0*
09
0>
0C
#29110000000
1!
1*
b111 6
19
1>
1C
b111 G
#29120000000
0!
0*
09
0>
0C
#29130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#29140000000
0!
0*
09
0>
0C
#29150000000
1!
1*
b1 6
19
1>
1C
b1 G
#29160000000
0!
0*
09
0>
0C
#29170000000
1!
1*
b10 6
19
1>
1C
b10 G
#29180000000
0!
0*
09
0>
0C
#29190000000
1!
1*
b11 6
19
1>
1C
b11 G
#29200000000
0!
0*
09
0>
0C
#29210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#29220000000
0!
0*
09
0>
0C
#29230000000
1!
1*
b101 6
19
1>
1C
b101 G
#29240000000
0!
0*
09
0>
0C
#29250000000
1!
1*
b110 6
19
1>
1C
b110 G
#29260000000
0!
0*
09
0>
0C
#29270000000
1!
1*
b111 6
19
1>
1C
b111 G
#29280000000
0!
1"
0*
1+
09
1:
0>
0C
#29290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#29300000000
0!
0*
09
0>
0C
#29310000000
1!
1*
b1 6
19
1>
1C
b1 G
#29320000000
0!
0*
09
0>
0C
#29330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#29340000000
0!
0*
09
0>
0C
#29350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#29360000000
0!
0*
09
0>
0C
#29370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#29380000000
0!
0*
09
0>
0C
#29390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#29400000000
0!
0#
0*
0,
09
0>
0?
0C
#29410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#29420000000
0!
0*
09
0>
0C
#29430000000
1!
1*
19
1>
1C
#29440000000
0!
0*
09
0>
0C
#29450000000
1!
1*
19
1>
1C
#29460000000
0!
0*
09
0>
0C
#29470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#29480000000
0!
0*
09
0>
0C
#29490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#29500000000
0!
0*
09
0>
0C
#29510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#29520000000
0!
0*
09
0>
0C
#29530000000
1!
1*
b10 6
19
1>
1C
b10 G
#29540000000
0!
0*
09
0>
0C
#29550000000
1!
1*
b11 6
19
1>
1C
b11 G
#29560000000
0!
0*
09
0>
0C
#29570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#29580000000
0!
0*
09
0>
0C
#29590000000
1!
1*
b101 6
19
1>
1C
b101 G
#29600000000
0!
0*
09
0>
0C
#29610000000
1!
1*
b110 6
19
1>
1C
b110 G
#29620000000
0!
0*
09
0>
0C
#29630000000
1!
1*
b111 6
19
1>
1C
b111 G
#29640000000
0!
0*
09
0>
0C
#29650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#29660000000
0!
0*
09
0>
0C
#29670000000
1!
1*
b1 6
19
1>
1C
b1 G
#29680000000
0!
0*
09
0>
0C
#29690000000
1!
1*
b10 6
19
1>
1C
b10 G
#29700000000
0!
0*
09
0>
0C
#29710000000
1!
1*
b11 6
19
1>
1C
b11 G
#29720000000
0!
0*
09
0>
0C
#29730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#29740000000
0!
0*
09
0>
0C
#29750000000
1!
1*
b101 6
19
1>
1C
b101 G
#29760000000
0!
0*
09
0>
0C
#29770000000
1!
1*
b110 6
19
1>
1C
b110 G
#29780000000
0!
0*
09
0>
0C
#29790000000
1!
1*
b111 6
19
1>
1C
b111 G
#29800000000
0!
0*
09
0>
0C
#29810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#29820000000
0!
0*
09
0>
0C
#29830000000
1!
1*
b1 6
19
1>
1C
b1 G
#29840000000
0!
0*
09
0>
0C
#29850000000
1!
1*
b10 6
19
1>
1C
b10 G
#29860000000
0!
0*
09
0>
0C
#29870000000
1!
1*
b11 6
19
1>
1C
b11 G
#29880000000
0!
0*
09
0>
0C
#29890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#29900000000
0!
0*
09
0>
0C
#29910000000
1!
1*
b101 6
19
1>
1C
b101 G
#29920000000
0!
0*
09
0>
0C
#29930000000
1!
1*
b110 6
19
1>
1C
b110 G
#29940000000
0!
0*
09
0>
0C
#29950000000
1!
1*
b111 6
19
1>
1C
b111 G
#29960000000
0!
1"
0*
1+
09
1:
0>
0C
#29970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#29980000000
0!
0*
09
0>
0C
#29990000000
1!
1*
b1 6
19
1>
1C
b1 G
#30000000000
0!
0*
09
0>
0C
#30010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#30020000000
0!
0*
09
0>
0C
#30030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#30040000000
0!
0*
09
0>
0C
#30050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#30060000000
0!
0*
09
0>
0C
#30070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#30080000000
0!
0#
0*
0,
09
0>
0?
0C
#30090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#30100000000
0!
0*
09
0>
0C
#30110000000
1!
1*
19
1>
1C
#30120000000
0!
0*
09
0>
0C
#30130000000
1!
1*
19
1>
1C
#30140000000
0!
0*
09
0>
0C
#30150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#30160000000
0!
0*
09
0>
0C
#30170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#30180000000
0!
0*
09
0>
0C
#30190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#30200000000
0!
0*
09
0>
0C
#30210000000
1!
1*
b10 6
19
1>
1C
b10 G
#30220000000
0!
0*
09
0>
0C
#30230000000
1!
1*
b11 6
19
1>
1C
b11 G
#30240000000
0!
0*
09
0>
0C
#30250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#30260000000
0!
0*
09
0>
0C
#30270000000
1!
1*
b101 6
19
1>
1C
b101 G
#30280000000
0!
0*
09
0>
0C
#30290000000
1!
1*
b110 6
19
1>
1C
b110 G
#30300000000
0!
0*
09
0>
0C
#30310000000
1!
1*
b111 6
19
1>
1C
b111 G
#30320000000
0!
0*
09
0>
0C
#30330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#30340000000
0!
0*
09
0>
0C
#30350000000
1!
1*
b1 6
19
1>
1C
b1 G
#30360000000
0!
0*
09
0>
0C
#30370000000
1!
1*
b10 6
19
1>
1C
b10 G
#30380000000
0!
0*
09
0>
0C
#30390000000
1!
1*
b11 6
19
1>
1C
b11 G
#30400000000
0!
0*
09
0>
0C
#30410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#30420000000
0!
0*
09
0>
0C
#30430000000
1!
1*
b101 6
19
1>
1C
b101 G
#30440000000
0!
0*
09
0>
0C
#30450000000
1!
1*
b110 6
19
1>
1C
b110 G
#30460000000
0!
0*
09
0>
0C
#30470000000
1!
1*
b111 6
19
1>
1C
b111 G
#30480000000
0!
0*
09
0>
0C
#30490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#30500000000
0!
0*
09
0>
0C
#30510000000
1!
1*
b1 6
19
1>
1C
b1 G
#30520000000
0!
0*
09
0>
0C
#30530000000
1!
1*
b10 6
19
1>
1C
b10 G
#30540000000
0!
0*
09
0>
0C
#30550000000
1!
1*
b11 6
19
1>
1C
b11 G
#30560000000
0!
0*
09
0>
0C
#30570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#30580000000
0!
0*
09
0>
0C
#30590000000
1!
1*
b101 6
19
1>
1C
b101 G
#30600000000
0!
0*
09
0>
0C
#30610000000
1!
1*
b110 6
19
1>
1C
b110 G
#30620000000
0!
0*
09
0>
0C
#30630000000
1!
1*
b111 6
19
1>
1C
b111 G
#30640000000
0!
1"
0*
1+
09
1:
0>
0C
#30650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#30660000000
0!
0*
09
0>
0C
#30670000000
1!
1*
b1 6
19
1>
1C
b1 G
#30680000000
0!
0*
09
0>
0C
#30690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#30700000000
0!
0*
09
0>
0C
#30710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#30720000000
0!
0*
09
0>
0C
#30730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#30740000000
0!
0*
09
0>
0C
#30750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#30760000000
0!
0#
0*
0,
09
0>
0?
0C
#30770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#30780000000
0!
0*
09
0>
0C
#30790000000
1!
1*
19
1>
1C
#30800000000
0!
0*
09
0>
0C
#30810000000
1!
1*
19
1>
1C
#30820000000
0!
0*
09
0>
0C
#30830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#30840000000
0!
0*
09
0>
0C
#30850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#30860000000
0!
0*
09
0>
0C
#30870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#30880000000
0!
0*
09
0>
0C
#30890000000
1!
1*
b10 6
19
1>
1C
b10 G
#30900000000
0!
0*
09
0>
0C
#30910000000
1!
1*
b11 6
19
1>
1C
b11 G
#30920000000
0!
0*
09
0>
0C
#30930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#30940000000
0!
0*
09
0>
0C
#30950000000
1!
1*
b101 6
19
1>
1C
b101 G
#30960000000
0!
0*
09
0>
0C
#30970000000
1!
1*
b110 6
19
1>
1C
b110 G
#30980000000
0!
0*
09
0>
0C
#30990000000
1!
1*
b111 6
19
1>
1C
b111 G
#31000000000
0!
0*
09
0>
0C
#31010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#31020000000
0!
0*
09
0>
0C
#31030000000
1!
1*
b1 6
19
1>
1C
b1 G
#31040000000
0!
0*
09
0>
0C
#31050000000
1!
1*
b10 6
19
1>
1C
b10 G
#31060000000
0!
0*
09
0>
0C
#31070000000
1!
1*
b11 6
19
1>
1C
b11 G
#31080000000
0!
0*
09
0>
0C
#31090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#31100000000
0!
0*
09
0>
0C
#31110000000
1!
1*
b101 6
19
1>
1C
b101 G
#31120000000
0!
0*
09
0>
0C
#31130000000
1!
1*
b110 6
19
1>
1C
b110 G
#31140000000
0!
0*
09
0>
0C
#31150000000
1!
1*
b111 6
19
1>
1C
b111 G
#31160000000
0!
0*
09
0>
0C
#31170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#31180000000
0!
0*
09
0>
0C
#31190000000
1!
1*
b1 6
19
1>
1C
b1 G
#31200000000
0!
0*
09
0>
0C
#31210000000
1!
1*
b10 6
19
1>
1C
b10 G
#31220000000
0!
0*
09
0>
0C
#31230000000
1!
1*
b11 6
19
1>
1C
b11 G
#31240000000
0!
0*
09
0>
0C
#31250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#31260000000
0!
0*
09
0>
0C
#31270000000
1!
1*
b101 6
19
1>
1C
b101 G
#31280000000
0!
0*
09
0>
0C
#31290000000
1!
1*
b110 6
19
1>
1C
b110 G
#31300000000
0!
0*
09
0>
0C
#31310000000
1!
1*
b111 6
19
1>
1C
b111 G
#31320000000
0!
1"
0*
1+
09
1:
0>
0C
#31330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#31340000000
0!
0*
09
0>
0C
#31350000000
1!
1*
b1 6
19
1>
1C
b1 G
#31360000000
0!
0*
09
0>
0C
#31370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#31380000000
0!
0*
09
0>
0C
#31390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#31400000000
0!
0*
09
0>
0C
#31410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#31420000000
0!
0*
09
0>
0C
#31430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#31440000000
0!
0#
0*
0,
09
0>
0?
0C
#31450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#31460000000
0!
0*
09
0>
0C
#31470000000
1!
1*
19
1>
1C
#31480000000
0!
0*
09
0>
0C
#31490000000
1!
1*
19
1>
1C
#31500000000
0!
0*
09
0>
0C
#31510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#31520000000
0!
0*
09
0>
0C
#31530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#31540000000
0!
0*
09
0>
0C
#31550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#31560000000
0!
0*
09
0>
0C
#31570000000
1!
1*
b10 6
19
1>
1C
b10 G
#31580000000
0!
0*
09
0>
0C
#31590000000
1!
1*
b11 6
19
1>
1C
b11 G
#31600000000
0!
0*
09
0>
0C
#31610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#31620000000
0!
0*
09
0>
0C
#31630000000
1!
1*
b101 6
19
1>
1C
b101 G
#31640000000
0!
0*
09
0>
0C
#31650000000
1!
1*
b110 6
19
1>
1C
b110 G
#31660000000
0!
0*
09
0>
0C
#31670000000
1!
1*
b111 6
19
1>
1C
b111 G
#31680000000
0!
0*
09
0>
0C
#31690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#31700000000
0!
0*
09
0>
0C
#31710000000
1!
1*
b1 6
19
1>
1C
b1 G
#31720000000
0!
0*
09
0>
0C
#31730000000
1!
1*
b10 6
19
1>
1C
b10 G
#31740000000
0!
0*
09
0>
0C
#31750000000
1!
1*
b11 6
19
1>
1C
b11 G
#31760000000
0!
0*
09
0>
0C
#31770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#31780000000
0!
0*
09
0>
0C
#31790000000
1!
1*
b101 6
19
1>
1C
b101 G
#31800000000
0!
0*
09
0>
0C
#31810000000
1!
1*
b110 6
19
1>
1C
b110 G
#31820000000
0!
0*
09
0>
0C
#31830000000
1!
1*
b111 6
19
1>
1C
b111 G
#31840000000
0!
0*
09
0>
0C
#31850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#31860000000
0!
0*
09
0>
0C
#31870000000
1!
1*
b1 6
19
1>
1C
b1 G
#31880000000
0!
0*
09
0>
0C
#31890000000
1!
1*
b10 6
19
1>
1C
b10 G
#31900000000
0!
0*
09
0>
0C
#31910000000
1!
1*
b11 6
19
1>
1C
b11 G
#31920000000
0!
0*
09
0>
0C
#31930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#31940000000
0!
0*
09
0>
0C
#31950000000
1!
1*
b101 6
19
1>
1C
b101 G
#31960000000
0!
0*
09
0>
0C
#31970000000
1!
1*
b110 6
19
1>
1C
b110 G
#31980000000
0!
0*
09
0>
0C
#31990000000
1!
1*
b111 6
19
1>
1C
b111 G
#32000000000
0!
1"
0*
1+
09
1:
0>
0C
#32010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#32020000000
0!
0*
09
0>
0C
#32030000000
1!
1*
b1 6
19
1>
1C
b1 G
#32040000000
0!
0*
09
0>
0C
#32050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#32060000000
0!
0*
09
0>
0C
#32070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#32080000000
0!
0*
09
0>
0C
#32090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#32100000000
0!
0*
09
0>
0C
#32110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#32120000000
0!
0#
0*
0,
09
0>
0?
0C
#32130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#32140000000
0!
0*
09
0>
0C
#32150000000
1!
1*
19
1>
1C
#32160000000
0!
0*
09
0>
0C
#32170000000
1!
1*
19
1>
1C
#32180000000
0!
0*
09
0>
0C
#32190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#32200000000
0!
0*
09
0>
0C
#32210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#32220000000
0!
0*
09
0>
0C
#32230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#32240000000
0!
0*
09
0>
0C
#32250000000
1!
1*
b10 6
19
1>
1C
b10 G
#32260000000
0!
0*
09
0>
0C
#32270000000
1!
1*
b11 6
19
1>
1C
b11 G
#32280000000
0!
0*
09
0>
0C
#32290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#32300000000
0!
0*
09
0>
0C
#32310000000
1!
1*
b101 6
19
1>
1C
b101 G
#32320000000
0!
0*
09
0>
0C
#32330000000
1!
1*
b110 6
19
1>
1C
b110 G
#32340000000
0!
0*
09
0>
0C
#32350000000
1!
1*
b111 6
19
1>
1C
b111 G
#32360000000
0!
0*
09
0>
0C
#32370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#32380000000
0!
0*
09
0>
0C
#32390000000
1!
1*
b1 6
19
1>
1C
b1 G
#32400000000
0!
0*
09
0>
0C
#32410000000
1!
1*
b10 6
19
1>
1C
b10 G
#32420000000
0!
0*
09
0>
0C
#32430000000
1!
1*
b11 6
19
1>
1C
b11 G
#32440000000
0!
0*
09
0>
0C
#32450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#32460000000
0!
0*
09
0>
0C
#32470000000
1!
1*
b101 6
19
1>
1C
b101 G
#32480000000
0!
0*
09
0>
0C
#32490000000
1!
1*
b110 6
19
1>
1C
b110 G
#32500000000
0!
0*
09
0>
0C
#32510000000
1!
1*
b111 6
19
1>
1C
b111 G
#32520000000
0!
0*
09
0>
0C
#32530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#32540000000
0!
0*
09
0>
0C
#32550000000
1!
1*
b1 6
19
1>
1C
b1 G
#32560000000
0!
0*
09
0>
0C
#32570000000
1!
1*
b10 6
19
1>
1C
b10 G
#32580000000
0!
0*
09
0>
0C
#32590000000
1!
1*
b11 6
19
1>
1C
b11 G
#32600000000
0!
0*
09
0>
0C
#32610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#32620000000
0!
0*
09
0>
0C
#32630000000
1!
1*
b101 6
19
1>
1C
b101 G
#32640000000
0!
0*
09
0>
0C
#32650000000
1!
1*
b110 6
19
1>
1C
b110 G
#32660000000
0!
0*
09
0>
0C
#32670000000
1!
1*
b111 6
19
1>
1C
b111 G
#32680000000
0!
1"
0*
1+
09
1:
0>
0C
#32690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#32700000000
0!
0*
09
0>
0C
#32710000000
1!
1*
b1 6
19
1>
1C
b1 G
#32720000000
0!
0*
09
0>
0C
#32730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#32740000000
0!
0*
09
0>
0C
#32750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#32760000000
0!
0*
09
0>
0C
#32770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#32780000000
0!
0*
09
0>
0C
#32790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#32800000000
0!
0#
0*
0,
09
0>
0?
0C
#32810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#32820000000
0!
0*
09
0>
0C
#32830000000
1!
1*
19
1>
1C
#32840000000
0!
0*
09
0>
0C
#32850000000
1!
1*
19
1>
1C
#32860000000
0!
0*
09
0>
0C
#32870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#32880000000
0!
0*
09
0>
0C
#32890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#32900000000
0!
0*
09
0>
0C
#32910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#32920000000
0!
0*
09
0>
0C
#32930000000
1!
1*
b10 6
19
1>
1C
b10 G
#32940000000
0!
0*
09
0>
0C
#32950000000
1!
1*
b11 6
19
1>
1C
b11 G
#32960000000
0!
0*
09
0>
0C
#32970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#32980000000
0!
0*
09
0>
0C
#32990000000
1!
1*
b101 6
19
1>
1C
b101 G
#33000000000
0!
0*
09
0>
0C
#33010000000
1!
1*
b110 6
19
1>
1C
b110 G
#33020000000
0!
0*
09
0>
0C
#33030000000
1!
1*
b111 6
19
1>
1C
b111 G
#33040000000
0!
0*
09
0>
0C
#33050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#33060000000
0!
0*
09
0>
0C
#33070000000
1!
1*
b1 6
19
1>
1C
b1 G
#33080000000
0!
0*
09
0>
0C
#33090000000
1!
1*
b10 6
19
1>
1C
b10 G
#33100000000
0!
0*
09
0>
0C
#33110000000
1!
1*
b11 6
19
1>
1C
b11 G
#33120000000
0!
0*
09
0>
0C
#33130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#33140000000
0!
0*
09
0>
0C
#33150000000
1!
1*
b101 6
19
1>
1C
b101 G
#33160000000
0!
0*
09
0>
0C
#33170000000
1!
1*
b110 6
19
1>
1C
b110 G
#33180000000
0!
0*
09
0>
0C
#33190000000
1!
1*
b111 6
19
1>
1C
b111 G
#33200000000
0!
0*
09
0>
0C
#33210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#33220000000
0!
0*
09
0>
0C
#33230000000
1!
1*
b1 6
19
1>
1C
b1 G
#33240000000
0!
0*
09
0>
0C
#33250000000
1!
1*
b10 6
19
1>
1C
b10 G
#33260000000
0!
0*
09
0>
0C
#33270000000
1!
1*
b11 6
19
1>
1C
b11 G
#33280000000
0!
0*
09
0>
0C
#33290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#33300000000
0!
0*
09
0>
0C
#33310000000
1!
1*
b101 6
19
1>
1C
b101 G
#33320000000
0!
0*
09
0>
0C
#33330000000
1!
1*
b110 6
19
1>
1C
b110 G
#33340000000
0!
0*
09
0>
0C
#33350000000
1!
1*
b111 6
19
1>
1C
b111 G
#33360000000
0!
1"
0*
1+
09
1:
0>
0C
#33370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#33380000000
0!
0*
09
0>
0C
#33390000000
1!
1*
b1 6
19
1>
1C
b1 G
#33400000000
0!
0*
09
0>
0C
#33410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#33420000000
0!
0*
09
0>
0C
#33430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#33440000000
0!
0*
09
0>
0C
#33450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#33460000000
0!
0*
09
0>
0C
#33470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#33480000000
0!
0#
0*
0,
09
0>
0?
0C
#33490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#33500000000
0!
0*
09
0>
0C
#33510000000
1!
1*
19
1>
1C
#33520000000
0!
0*
09
0>
0C
#33530000000
1!
1*
19
1>
1C
#33540000000
0!
0*
09
0>
0C
#33550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#33560000000
0!
0*
09
0>
0C
#33570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#33580000000
0!
0*
09
0>
0C
#33590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#33600000000
0!
0*
09
0>
0C
#33610000000
1!
1*
b10 6
19
1>
1C
b10 G
#33620000000
0!
0*
09
0>
0C
#33630000000
1!
1*
b11 6
19
1>
1C
b11 G
#33640000000
0!
0*
09
0>
0C
#33650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#33660000000
0!
0*
09
0>
0C
#33670000000
1!
1*
b101 6
19
1>
1C
b101 G
#33680000000
0!
0*
09
0>
0C
#33690000000
1!
1*
b110 6
19
1>
1C
b110 G
#33700000000
0!
0*
09
0>
0C
#33710000000
1!
1*
b111 6
19
1>
1C
b111 G
#33720000000
0!
0*
09
0>
0C
#33730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#33740000000
0!
0*
09
0>
0C
#33750000000
1!
1*
b1 6
19
1>
1C
b1 G
#33760000000
0!
0*
09
0>
0C
#33770000000
1!
1*
b10 6
19
1>
1C
b10 G
#33780000000
0!
0*
09
0>
0C
#33790000000
1!
1*
b11 6
19
1>
1C
b11 G
#33800000000
0!
0*
09
0>
0C
#33810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#33820000000
0!
0*
09
0>
0C
#33830000000
1!
1*
b101 6
19
1>
1C
b101 G
#33840000000
0!
0*
09
0>
0C
#33850000000
1!
1*
b110 6
19
1>
1C
b110 G
#33860000000
0!
0*
09
0>
0C
#33870000000
1!
1*
b111 6
19
1>
1C
b111 G
#33880000000
0!
0*
09
0>
0C
#33890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#33900000000
0!
0*
09
0>
0C
#33910000000
1!
1*
b1 6
19
1>
1C
b1 G
#33920000000
0!
0*
09
0>
0C
#33930000000
1!
1*
b10 6
19
1>
1C
b10 G
#33940000000
0!
0*
09
0>
0C
#33950000000
1!
1*
b11 6
19
1>
1C
b11 G
#33960000000
0!
0*
09
0>
0C
#33970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#33980000000
0!
0*
09
0>
0C
#33990000000
1!
1*
b101 6
19
1>
1C
b101 G
#34000000000
0!
0*
09
0>
0C
#34010000000
1!
1*
b110 6
19
1>
1C
b110 G
#34020000000
0!
0*
09
0>
0C
#34030000000
1!
1*
b111 6
19
1>
1C
b111 G
#34040000000
0!
1"
0*
1+
09
1:
0>
0C
#34050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#34060000000
0!
0*
09
0>
0C
#34070000000
1!
1*
b1 6
19
1>
1C
b1 G
#34080000000
0!
0*
09
0>
0C
#34090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#34100000000
0!
0*
09
0>
0C
#34110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#34120000000
0!
0*
09
0>
0C
#34130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#34140000000
0!
0*
09
0>
0C
#34150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#34160000000
0!
0#
0*
0,
09
0>
0?
0C
#34170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#34180000000
0!
0*
09
0>
0C
#34190000000
1!
1*
19
1>
1C
#34200000000
0!
0*
09
0>
0C
#34210000000
1!
1*
19
1>
1C
#34220000000
0!
0*
09
0>
0C
#34230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#34240000000
0!
0*
09
0>
0C
#34250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#34260000000
0!
0*
09
0>
0C
#34270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#34280000000
0!
0*
09
0>
0C
#34290000000
1!
1*
b10 6
19
1>
1C
b10 G
#34300000000
0!
0*
09
0>
0C
#34310000000
1!
1*
b11 6
19
1>
1C
b11 G
#34320000000
0!
0*
09
0>
0C
#34330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#34340000000
0!
0*
09
0>
0C
#34350000000
1!
1*
b101 6
19
1>
1C
b101 G
#34360000000
0!
0*
09
0>
0C
#34370000000
1!
1*
b110 6
19
1>
1C
b110 G
#34380000000
0!
0*
09
0>
0C
#34390000000
1!
1*
b111 6
19
1>
1C
b111 G
#34400000000
0!
0*
09
0>
0C
#34410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#34420000000
0!
0*
09
0>
0C
#34430000000
1!
1*
b1 6
19
1>
1C
b1 G
#34440000000
0!
0*
09
0>
0C
#34450000000
1!
1*
b10 6
19
1>
1C
b10 G
#34460000000
0!
0*
09
0>
0C
#34470000000
1!
1*
b11 6
19
1>
1C
b11 G
#34480000000
0!
0*
09
0>
0C
#34490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#34500000000
0!
0*
09
0>
0C
#34510000000
1!
1*
b101 6
19
1>
1C
b101 G
#34520000000
0!
0*
09
0>
0C
#34530000000
1!
1*
b110 6
19
1>
1C
b110 G
#34540000000
0!
0*
09
0>
0C
#34550000000
1!
1*
b111 6
19
1>
1C
b111 G
#34560000000
0!
0*
09
0>
0C
#34570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#34580000000
0!
0*
09
0>
0C
#34590000000
1!
1*
b1 6
19
1>
1C
b1 G
#34600000000
0!
0*
09
0>
0C
#34610000000
1!
1*
b10 6
19
1>
1C
b10 G
#34620000000
0!
0*
09
0>
0C
#34630000000
1!
1*
b11 6
19
1>
1C
b11 G
#34640000000
0!
0*
09
0>
0C
#34650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#34660000000
0!
0*
09
0>
0C
#34670000000
1!
1*
b101 6
19
1>
1C
b101 G
#34680000000
0!
0*
09
0>
0C
#34690000000
1!
1*
b110 6
19
1>
1C
b110 G
#34700000000
0!
0*
09
0>
0C
#34710000000
1!
1*
b111 6
19
1>
1C
b111 G
#34720000000
0!
1"
0*
1+
09
1:
0>
0C
#34730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#34740000000
0!
0*
09
0>
0C
#34750000000
1!
1*
b1 6
19
1>
1C
b1 G
#34760000000
0!
0*
09
0>
0C
#34770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#34780000000
0!
0*
09
0>
0C
#34790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#34800000000
0!
0*
09
0>
0C
#34810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#34820000000
0!
0*
09
0>
0C
#34830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#34840000000
0!
0#
0*
0,
09
0>
0?
0C
#34850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#34860000000
0!
0*
09
0>
0C
#34870000000
1!
1*
19
1>
1C
#34880000000
0!
0*
09
0>
0C
#34890000000
1!
1*
19
1>
1C
#34900000000
0!
0*
09
0>
0C
#34910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#34920000000
0!
0*
09
0>
0C
#34930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#34940000000
0!
0*
09
0>
0C
#34950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#34960000000
0!
0*
09
0>
0C
#34970000000
1!
1*
b10 6
19
1>
1C
b10 G
#34980000000
0!
0*
09
0>
0C
#34990000000
1!
1*
b11 6
19
1>
1C
b11 G
#35000000000
0!
0*
09
0>
0C
#35010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#35020000000
0!
0*
09
0>
0C
#35030000000
1!
1*
b101 6
19
1>
1C
b101 G
#35040000000
0!
0*
09
0>
0C
#35050000000
1!
1*
b110 6
19
1>
1C
b110 G
#35060000000
0!
0*
09
0>
0C
#35070000000
1!
1*
b111 6
19
1>
1C
b111 G
#35080000000
0!
0*
09
0>
0C
#35090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#35100000000
0!
0*
09
0>
0C
#35110000000
1!
1*
b1 6
19
1>
1C
b1 G
#35120000000
0!
0*
09
0>
0C
#35130000000
1!
1*
b10 6
19
1>
1C
b10 G
#35140000000
0!
0*
09
0>
0C
#35150000000
1!
1*
b11 6
19
1>
1C
b11 G
#35160000000
0!
0*
09
0>
0C
#35170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#35180000000
0!
0*
09
0>
0C
#35190000000
1!
1*
b101 6
19
1>
1C
b101 G
#35200000000
0!
0*
09
0>
0C
#35210000000
1!
1*
b110 6
19
1>
1C
b110 G
#35220000000
0!
0*
09
0>
0C
#35230000000
1!
1*
b111 6
19
1>
1C
b111 G
#35240000000
0!
0*
09
0>
0C
#35250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#35260000000
0!
0*
09
0>
0C
#35270000000
1!
1*
b1 6
19
1>
1C
b1 G
#35280000000
0!
0*
09
0>
0C
#35290000000
1!
1*
b10 6
19
1>
1C
b10 G
#35300000000
0!
0*
09
0>
0C
#35310000000
1!
1*
b11 6
19
1>
1C
b11 G
#35320000000
0!
0*
09
0>
0C
#35330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#35340000000
0!
0*
09
0>
0C
#35350000000
1!
1*
b101 6
19
1>
1C
b101 G
#35360000000
0!
0*
09
0>
0C
#35370000000
1!
1*
b110 6
19
1>
1C
b110 G
#35380000000
0!
0*
09
0>
0C
#35390000000
1!
1*
b111 6
19
1>
1C
b111 G
#35400000000
0!
1"
0*
1+
09
1:
0>
0C
#35410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#35420000000
0!
0*
09
0>
0C
#35430000000
1!
1*
b1 6
19
1>
1C
b1 G
#35440000000
0!
0*
09
0>
0C
#35450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#35460000000
0!
0*
09
0>
0C
#35470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#35480000000
0!
0*
09
0>
0C
#35490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#35500000000
0!
0*
09
0>
0C
#35510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#35520000000
0!
0#
0*
0,
09
0>
0?
0C
#35530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#35540000000
0!
0*
09
0>
0C
#35550000000
1!
1*
19
1>
1C
#35560000000
0!
0*
09
0>
0C
#35570000000
1!
1*
19
1>
1C
#35580000000
0!
0*
09
0>
0C
#35590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#35600000000
0!
0*
09
0>
0C
#35610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#35620000000
0!
0*
09
0>
0C
#35630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#35640000000
0!
0*
09
0>
0C
#35650000000
1!
1*
b10 6
19
1>
1C
b10 G
#35660000000
0!
0*
09
0>
0C
#35670000000
1!
1*
b11 6
19
1>
1C
b11 G
#35680000000
0!
0*
09
0>
0C
#35690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#35700000000
0!
0*
09
0>
0C
#35710000000
1!
1*
b101 6
19
1>
1C
b101 G
#35720000000
0!
0*
09
0>
0C
#35730000000
1!
1*
b110 6
19
1>
1C
b110 G
#35740000000
0!
0*
09
0>
0C
#35750000000
1!
1*
b111 6
19
1>
1C
b111 G
#35760000000
0!
0*
09
0>
0C
#35770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#35780000000
0!
0*
09
0>
0C
#35790000000
1!
1*
b1 6
19
1>
1C
b1 G
#35800000000
0!
0*
09
0>
0C
#35810000000
1!
1*
b10 6
19
1>
1C
b10 G
#35820000000
0!
0*
09
0>
0C
#35830000000
1!
1*
b11 6
19
1>
1C
b11 G
#35840000000
0!
0*
09
0>
0C
#35850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#35860000000
0!
0*
09
0>
0C
#35870000000
1!
1*
b101 6
19
1>
1C
b101 G
#35880000000
0!
0*
09
0>
0C
#35890000000
1!
1*
b110 6
19
1>
1C
b110 G
#35900000000
0!
0*
09
0>
0C
#35910000000
1!
1*
b111 6
19
1>
1C
b111 G
#35920000000
0!
0*
09
0>
0C
#35930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#35940000000
0!
0*
09
0>
0C
#35950000000
1!
1*
b1 6
19
1>
1C
b1 G
#35960000000
0!
0*
09
0>
0C
#35970000000
1!
1*
b10 6
19
1>
1C
b10 G
#35980000000
0!
0*
09
0>
0C
#35990000000
1!
1*
b11 6
19
1>
1C
b11 G
#36000000000
0!
0*
09
0>
0C
#36010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#36020000000
0!
0*
09
0>
0C
#36030000000
1!
1*
b101 6
19
1>
1C
b101 G
#36040000000
0!
0*
09
0>
0C
#36050000000
1!
1*
b110 6
19
1>
1C
b110 G
#36060000000
0!
0*
09
0>
0C
#36070000000
1!
1*
b111 6
19
1>
1C
b111 G
#36080000000
0!
1"
0*
1+
09
1:
0>
0C
#36090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#36100000000
0!
0*
09
0>
0C
#36110000000
1!
1*
b1 6
19
1>
1C
b1 G
#36120000000
0!
0*
09
0>
0C
#36130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#36140000000
0!
0*
09
0>
0C
#36150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#36160000000
0!
0*
09
0>
0C
#36170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#36180000000
0!
0*
09
0>
0C
#36190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#36200000000
0!
0#
0*
0,
09
0>
0?
0C
#36210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#36220000000
0!
0*
09
0>
0C
#36230000000
1!
1*
19
1>
1C
#36240000000
0!
0*
09
0>
0C
#36250000000
1!
1*
19
1>
1C
#36260000000
0!
0*
09
0>
0C
#36270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#36280000000
0!
0*
09
0>
0C
#36290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#36300000000
0!
0*
09
0>
0C
#36310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#36320000000
0!
0*
09
0>
0C
#36330000000
1!
1*
b10 6
19
1>
1C
b10 G
#36340000000
0!
0*
09
0>
0C
#36350000000
1!
1*
b11 6
19
1>
1C
b11 G
#36360000000
0!
0*
09
0>
0C
#36370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#36380000000
0!
0*
09
0>
0C
#36390000000
1!
1*
b101 6
19
1>
1C
b101 G
#36400000000
0!
0*
09
0>
0C
#36410000000
1!
1*
b110 6
19
1>
1C
b110 G
#36420000000
0!
0*
09
0>
0C
#36430000000
1!
1*
b111 6
19
1>
1C
b111 G
#36440000000
0!
0*
09
0>
0C
#36450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#36460000000
0!
0*
09
0>
0C
#36470000000
1!
1*
b1 6
19
1>
1C
b1 G
#36480000000
0!
0*
09
0>
0C
#36490000000
1!
1*
b10 6
19
1>
1C
b10 G
#36500000000
0!
0*
09
0>
0C
#36510000000
1!
1*
b11 6
19
1>
1C
b11 G
#36520000000
0!
0*
09
0>
0C
#36530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#36540000000
0!
0*
09
0>
0C
#36550000000
1!
1*
b101 6
19
1>
1C
b101 G
#36560000000
0!
0*
09
0>
0C
#36570000000
1!
1*
b110 6
19
1>
1C
b110 G
#36580000000
0!
0*
09
0>
0C
#36590000000
1!
1*
b111 6
19
1>
1C
b111 G
#36600000000
0!
0*
09
0>
0C
#36610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#36620000000
0!
0*
09
0>
0C
#36630000000
1!
1*
b1 6
19
1>
1C
b1 G
#36640000000
0!
0*
09
0>
0C
#36650000000
1!
1*
b10 6
19
1>
1C
b10 G
#36660000000
0!
0*
09
0>
0C
#36670000000
1!
1*
b11 6
19
1>
1C
b11 G
#36680000000
0!
0*
09
0>
0C
#36690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#36700000000
0!
0*
09
0>
0C
#36710000000
1!
1*
b101 6
19
1>
1C
b101 G
#36720000000
0!
0*
09
0>
0C
#36730000000
1!
1*
b110 6
19
1>
1C
b110 G
#36740000000
0!
0*
09
0>
0C
#36750000000
1!
1*
b111 6
19
1>
1C
b111 G
#36760000000
0!
1"
0*
1+
09
1:
0>
0C
#36770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#36780000000
0!
0*
09
0>
0C
#36790000000
1!
1*
b1 6
19
1>
1C
b1 G
#36800000000
0!
0*
09
0>
0C
#36810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#36820000000
0!
0*
09
0>
0C
#36830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#36840000000
0!
0*
09
0>
0C
#36850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#36860000000
0!
0*
09
0>
0C
#36870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#36880000000
0!
0#
0*
0,
09
0>
0?
0C
#36890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#36900000000
0!
0*
09
0>
0C
#36910000000
1!
1*
19
1>
1C
#36920000000
0!
0*
09
0>
0C
#36930000000
1!
1*
19
1>
1C
#36940000000
0!
0*
09
0>
0C
#36950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#36960000000
0!
0*
09
0>
0C
#36970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#36980000000
0!
0*
09
0>
0C
#36990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#37000000000
0!
0*
09
0>
0C
#37010000000
1!
1*
b10 6
19
1>
1C
b10 G
#37020000000
0!
0*
09
0>
0C
#37030000000
1!
1*
b11 6
19
1>
1C
b11 G
#37040000000
0!
0*
09
0>
0C
#37050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#37060000000
0!
0*
09
0>
0C
#37070000000
1!
1*
b101 6
19
1>
1C
b101 G
#37080000000
0!
0*
09
0>
0C
#37090000000
1!
1*
b110 6
19
1>
1C
b110 G
#37100000000
0!
0*
09
0>
0C
#37110000000
1!
1*
b111 6
19
1>
1C
b111 G
#37120000000
0!
0*
09
0>
0C
#37130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#37140000000
0!
0*
09
0>
0C
#37150000000
1!
1*
b1 6
19
1>
1C
b1 G
#37160000000
0!
0*
09
0>
0C
#37170000000
1!
1*
b10 6
19
1>
1C
b10 G
#37180000000
0!
0*
09
0>
0C
#37190000000
1!
1*
b11 6
19
1>
1C
b11 G
#37200000000
0!
0*
09
0>
0C
#37210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#37220000000
0!
0*
09
0>
0C
#37230000000
1!
1*
b101 6
19
1>
1C
b101 G
#37240000000
0!
0*
09
0>
0C
#37250000000
1!
1*
b110 6
19
1>
1C
b110 G
#37260000000
0!
0*
09
0>
0C
#37270000000
1!
1*
b111 6
19
1>
1C
b111 G
#37280000000
0!
0*
09
0>
0C
#37290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#37300000000
0!
0*
09
0>
0C
#37310000000
1!
1*
b1 6
19
1>
1C
b1 G
#37320000000
0!
0*
09
0>
0C
#37330000000
1!
1*
b10 6
19
1>
1C
b10 G
#37340000000
0!
0*
09
0>
0C
#37350000000
1!
1*
b11 6
19
1>
1C
b11 G
#37360000000
0!
0*
09
0>
0C
#37370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#37380000000
0!
0*
09
0>
0C
#37390000000
1!
1*
b101 6
19
1>
1C
b101 G
#37400000000
0!
0*
09
0>
0C
#37410000000
1!
1*
b110 6
19
1>
1C
b110 G
#37420000000
0!
0*
09
0>
0C
#37430000000
1!
1*
b111 6
19
1>
1C
b111 G
#37440000000
0!
1"
0*
1+
09
1:
0>
0C
#37450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#37460000000
0!
0*
09
0>
0C
#37470000000
1!
1*
b1 6
19
1>
1C
b1 G
#37480000000
0!
0*
09
0>
0C
#37490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#37500000000
0!
0*
09
0>
0C
#37510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#37520000000
0!
0*
09
0>
0C
#37530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#37540000000
0!
0*
09
0>
0C
#37550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#37560000000
0!
0#
0*
0,
09
0>
0?
0C
#37570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#37580000000
0!
0*
09
0>
0C
#37590000000
1!
1*
19
1>
1C
#37600000000
0!
0*
09
0>
0C
#37610000000
1!
1*
19
1>
1C
#37620000000
0!
0*
09
0>
0C
#37630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#37640000000
0!
0*
09
0>
0C
#37650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#37660000000
0!
0*
09
0>
0C
#37670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#37680000000
0!
0*
09
0>
0C
#37690000000
1!
1*
b10 6
19
1>
1C
b10 G
#37700000000
0!
0*
09
0>
0C
#37710000000
1!
1*
b11 6
19
1>
1C
b11 G
#37720000000
0!
0*
09
0>
0C
#37730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#37740000000
0!
0*
09
0>
0C
#37750000000
1!
1*
b101 6
19
1>
1C
b101 G
#37760000000
0!
0*
09
0>
0C
#37770000000
1!
1*
b110 6
19
1>
1C
b110 G
#37780000000
0!
0*
09
0>
0C
#37790000000
1!
1*
b111 6
19
1>
1C
b111 G
#37800000000
0!
0*
09
0>
0C
#37810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#37820000000
0!
0*
09
0>
0C
#37830000000
1!
1*
b1 6
19
1>
1C
b1 G
#37840000000
0!
0*
09
0>
0C
#37850000000
1!
1*
b10 6
19
1>
1C
b10 G
#37860000000
0!
0*
09
0>
0C
#37870000000
1!
1*
b11 6
19
1>
1C
b11 G
#37880000000
0!
0*
09
0>
0C
#37890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#37900000000
0!
0*
09
0>
0C
#37910000000
1!
1*
b101 6
19
1>
1C
b101 G
#37920000000
0!
0*
09
0>
0C
#37930000000
1!
1*
b110 6
19
1>
1C
b110 G
#37940000000
0!
0*
09
0>
0C
#37950000000
1!
1*
b111 6
19
1>
1C
b111 G
#37960000000
0!
0*
09
0>
0C
#37970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#37980000000
0!
0*
09
0>
0C
#37990000000
1!
1*
b1 6
19
1>
1C
b1 G
#38000000000
0!
0*
09
0>
0C
#38010000000
1!
1*
b10 6
19
1>
1C
b10 G
#38020000000
0!
0*
09
0>
0C
#38030000000
1!
1*
b11 6
19
1>
1C
b11 G
#38040000000
0!
0*
09
0>
0C
#38050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#38060000000
0!
0*
09
0>
0C
#38070000000
1!
1*
b101 6
19
1>
1C
b101 G
#38080000000
0!
0*
09
0>
0C
#38090000000
1!
1*
b110 6
19
1>
1C
b110 G
#38100000000
0!
0*
09
0>
0C
#38110000000
1!
1*
b111 6
19
1>
1C
b111 G
#38120000000
0!
1"
0*
1+
09
1:
0>
0C
#38130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#38140000000
0!
0*
09
0>
0C
#38150000000
1!
1*
b1 6
19
1>
1C
b1 G
#38160000000
0!
0*
09
0>
0C
#38170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#38180000000
0!
0*
09
0>
0C
#38190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#38200000000
0!
0*
09
0>
0C
#38210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#38220000000
0!
0*
09
0>
0C
#38230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#38240000000
0!
0#
0*
0,
09
0>
0?
0C
#38250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#38260000000
0!
0*
09
0>
0C
#38270000000
1!
1*
19
1>
1C
#38280000000
0!
0*
09
0>
0C
#38290000000
1!
1*
19
1>
1C
#38300000000
0!
0*
09
0>
0C
#38310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#38320000000
0!
0*
09
0>
0C
#38330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#38340000000
0!
0*
09
0>
0C
#38350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#38360000000
0!
0*
09
0>
0C
#38370000000
1!
1*
b10 6
19
1>
1C
b10 G
#38380000000
0!
0*
09
0>
0C
#38390000000
1!
1*
b11 6
19
1>
1C
b11 G
#38400000000
0!
0*
09
0>
0C
#38410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#38420000000
0!
0*
09
0>
0C
#38430000000
1!
1*
b101 6
19
1>
1C
b101 G
#38440000000
0!
0*
09
0>
0C
#38450000000
1!
1*
b110 6
19
1>
1C
b110 G
#38460000000
0!
0*
09
0>
0C
#38470000000
1!
1*
b111 6
19
1>
1C
b111 G
#38480000000
0!
0*
09
0>
0C
#38490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#38500000000
0!
0*
09
0>
0C
#38510000000
1!
1*
b1 6
19
1>
1C
b1 G
#38520000000
0!
0*
09
0>
0C
#38530000000
1!
1*
b10 6
19
1>
1C
b10 G
#38540000000
0!
0*
09
0>
0C
#38550000000
1!
1*
b11 6
19
1>
1C
b11 G
#38560000000
0!
0*
09
0>
0C
#38570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#38580000000
0!
0*
09
0>
0C
#38590000000
1!
1*
b101 6
19
1>
1C
b101 G
#38600000000
0!
0*
09
0>
0C
#38610000000
1!
1*
b110 6
19
1>
1C
b110 G
#38620000000
0!
0*
09
0>
0C
#38630000000
1!
1*
b111 6
19
1>
1C
b111 G
#38640000000
0!
0*
09
0>
0C
#38650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#38660000000
0!
0*
09
0>
0C
#38670000000
1!
1*
b1 6
19
1>
1C
b1 G
#38680000000
0!
0*
09
0>
0C
#38690000000
1!
1*
b10 6
19
1>
1C
b10 G
#38700000000
0!
0*
09
0>
0C
#38710000000
1!
1*
b11 6
19
1>
1C
b11 G
#38720000000
0!
0*
09
0>
0C
#38730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#38740000000
0!
0*
09
0>
0C
#38750000000
1!
1*
b101 6
19
1>
1C
b101 G
#38760000000
0!
0*
09
0>
0C
#38770000000
1!
1*
b110 6
19
1>
1C
b110 G
#38780000000
0!
0*
09
0>
0C
#38790000000
1!
1*
b111 6
19
1>
1C
b111 G
#38800000000
0!
1"
0*
1+
09
1:
0>
0C
#38810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#38820000000
0!
0*
09
0>
0C
#38830000000
1!
1*
b1 6
19
1>
1C
b1 G
#38840000000
0!
0*
09
0>
0C
#38850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#38860000000
0!
0*
09
0>
0C
#38870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#38880000000
0!
0*
09
0>
0C
#38890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#38900000000
0!
0*
09
0>
0C
#38910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#38920000000
0!
0#
0*
0,
09
0>
0?
0C
#38930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#38940000000
0!
0*
09
0>
0C
#38950000000
1!
1*
19
1>
1C
#38960000000
0!
0*
09
0>
0C
#38970000000
1!
1*
19
1>
1C
#38980000000
0!
0*
09
0>
0C
#38990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#39000000000
0!
0*
09
0>
0C
#39010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#39020000000
0!
0*
09
0>
0C
#39030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#39040000000
0!
0*
09
0>
0C
#39050000000
1!
1*
b10 6
19
1>
1C
b10 G
#39060000000
0!
0*
09
0>
0C
#39070000000
1!
1*
b11 6
19
1>
1C
b11 G
#39080000000
0!
0*
09
0>
0C
#39090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#39100000000
0!
0*
09
0>
0C
#39110000000
1!
1*
b101 6
19
1>
1C
b101 G
#39120000000
0!
0*
09
0>
0C
#39130000000
1!
1*
b110 6
19
1>
1C
b110 G
#39140000000
0!
0*
09
0>
0C
#39150000000
1!
1*
b111 6
19
1>
1C
b111 G
#39160000000
0!
0*
09
0>
0C
#39170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#39180000000
0!
0*
09
0>
0C
#39190000000
1!
1*
b1 6
19
1>
1C
b1 G
#39200000000
0!
0*
09
0>
0C
#39210000000
1!
1*
b10 6
19
1>
1C
b10 G
#39220000000
0!
0*
09
0>
0C
#39230000000
1!
1*
b11 6
19
1>
1C
b11 G
#39240000000
0!
0*
09
0>
0C
#39250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#39260000000
0!
0*
09
0>
0C
#39270000000
1!
1*
b101 6
19
1>
1C
b101 G
#39280000000
0!
0*
09
0>
0C
#39290000000
1!
1*
b110 6
19
1>
1C
b110 G
#39300000000
0!
0*
09
0>
0C
#39310000000
1!
1*
b111 6
19
1>
1C
b111 G
#39320000000
0!
0*
09
0>
0C
#39330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#39340000000
0!
0*
09
0>
0C
#39350000000
1!
1*
b1 6
19
1>
1C
b1 G
#39360000000
0!
0*
09
0>
0C
#39370000000
1!
1*
b10 6
19
1>
1C
b10 G
#39380000000
0!
0*
09
0>
0C
#39390000000
1!
1*
b11 6
19
1>
1C
b11 G
#39400000000
0!
0*
09
0>
0C
#39410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#39420000000
0!
0*
09
0>
0C
#39430000000
1!
1*
b101 6
19
1>
1C
b101 G
#39440000000
0!
0*
09
0>
0C
#39450000000
1!
1*
b110 6
19
1>
1C
b110 G
#39460000000
0!
0*
09
0>
0C
#39470000000
1!
1*
b111 6
19
1>
1C
b111 G
#39480000000
0!
1"
0*
1+
09
1:
0>
0C
#39490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#39500000000
0!
0*
09
0>
0C
#39510000000
1!
1*
b1 6
19
1>
1C
b1 G
#39520000000
0!
0*
09
0>
0C
#39530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#39540000000
0!
0*
09
0>
0C
#39550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#39560000000
0!
0*
09
0>
0C
#39570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#39580000000
0!
0*
09
0>
0C
#39590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#39600000000
0!
0#
0*
0,
09
0>
0?
0C
#39610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#39620000000
0!
0*
09
0>
0C
#39630000000
1!
1*
19
1>
1C
#39640000000
0!
0*
09
0>
0C
#39650000000
1!
1*
19
1>
1C
#39660000000
0!
0*
09
0>
0C
#39670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#39680000000
0!
0*
09
0>
0C
#39690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#39700000000
0!
0*
09
0>
0C
#39710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#39720000000
0!
0*
09
0>
0C
#39730000000
1!
1*
b10 6
19
1>
1C
b10 G
#39740000000
0!
0*
09
0>
0C
#39750000000
1!
1*
b11 6
19
1>
1C
b11 G
#39760000000
0!
0*
09
0>
0C
#39770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#39780000000
0!
0*
09
0>
0C
#39790000000
1!
1*
b101 6
19
1>
1C
b101 G
#39800000000
0!
0*
09
0>
0C
#39810000000
1!
1*
b110 6
19
1>
1C
b110 G
#39820000000
0!
0*
09
0>
0C
#39830000000
1!
1*
b111 6
19
1>
1C
b111 G
#39840000000
0!
0*
09
0>
0C
#39850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#39860000000
0!
0*
09
0>
0C
#39870000000
1!
1*
b1 6
19
1>
1C
b1 G
#39880000000
0!
0*
09
0>
0C
#39890000000
1!
1*
b10 6
19
1>
1C
b10 G
#39900000000
0!
0*
09
0>
0C
#39910000000
1!
1*
b11 6
19
1>
1C
b11 G
#39920000000
0!
0*
09
0>
0C
#39930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#39940000000
0!
0*
09
0>
0C
#39950000000
1!
1*
b101 6
19
1>
1C
b101 G
#39960000000
0!
0*
09
0>
0C
#39970000000
1!
1*
b110 6
19
1>
1C
b110 G
#39980000000
0!
0*
09
0>
0C
#39990000000
1!
1*
b111 6
19
1>
1C
b111 G
#40000000000
0!
0*
09
0>
0C
#40010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#40020000000
0!
0*
09
0>
0C
#40030000000
1!
1*
b1 6
19
1>
1C
b1 G
#40040000000
0!
0*
09
0>
0C
#40050000000
1!
1*
b10 6
19
1>
1C
b10 G
#40060000000
0!
0*
09
0>
0C
#40070000000
1!
1*
b11 6
19
1>
1C
b11 G
#40080000000
0!
0*
09
0>
0C
#40090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#40100000000
0!
0*
09
0>
0C
#40110000000
1!
1*
b101 6
19
1>
1C
b101 G
#40120000000
0!
0*
09
0>
0C
#40130000000
1!
1*
b110 6
19
1>
1C
b110 G
#40140000000
0!
0*
09
0>
0C
#40150000000
1!
1*
b111 6
19
1>
1C
b111 G
#40160000000
0!
1"
0*
1+
09
1:
0>
0C
#40170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#40180000000
0!
0*
09
0>
0C
#40190000000
1!
1*
b1 6
19
1>
1C
b1 G
#40200000000
0!
0*
09
0>
0C
#40210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#40220000000
0!
0*
09
0>
0C
#40230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#40240000000
0!
0*
09
0>
0C
#40250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#40260000000
0!
0*
09
0>
0C
#40270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#40280000000
0!
0#
0*
0,
09
0>
0?
0C
#40290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#40300000000
0!
0*
09
0>
0C
#40310000000
1!
1*
19
1>
1C
#40320000000
0!
0*
09
0>
0C
#40330000000
1!
1*
19
1>
1C
#40340000000
0!
0*
09
0>
0C
#40350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#40360000000
0!
0*
09
0>
0C
#40370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#40380000000
0!
0*
09
0>
0C
#40390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#40400000000
0!
0*
09
0>
0C
#40410000000
1!
1*
b10 6
19
1>
1C
b10 G
#40420000000
0!
0*
09
0>
0C
#40430000000
1!
1*
b11 6
19
1>
1C
b11 G
#40440000000
0!
0*
09
0>
0C
#40450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#40460000000
0!
0*
09
0>
0C
#40470000000
1!
1*
b101 6
19
1>
1C
b101 G
#40480000000
0!
0*
09
0>
0C
#40490000000
1!
1*
b110 6
19
1>
1C
b110 G
#40500000000
0!
0*
09
0>
0C
#40510000000
1!
1*
b111 6
19
1>
1C
b111 G
#40520000000
0!
0*
09
0>
0C
#40530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#40540000000
0!
0*
09
0>
0C
#40550000000
1!
1*
b1 6
19
1>
1C
b1 G
#40560000000
0!
0*
09
0>
0C
#40570000000
1!
1*
b10 6
19
1>
1C
b10 G
#40580000000
0!
0*
09
0>
0C
#40590000000
1!
1*
b11 6
19
1>
1C
b11 G
#40600000000
0!
0*
09
0>
0C
#40610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#40620000000
0!
0*
09
0>
0C
#40630000000
1!
1*
b101 6
19
1>
1C
b101 G
#40640000000
0!
0*
09
0>
0C
#40650000000
1!
1*
b110 6
19
1>
1C
b110 G
#40660000000
0!
0*
09
0>
0C
#40670000000
1!
1*
b111 6
19
1>
1C
b111 G
#40680000000
0!
0*
09
0>
0C
#40690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#40700000000
0!
0*
09
0>
0C
#40710000000
1!
1*
b1 6
19
1>
1C
b1 G
#40720000000
0!
0*
09
0>
0C
#40730000000
1!
1*
b10 6
19
1>
1C
b10 G
#40740000000
0!
0*
09
0>
0C
#40750000000
1!
1*
b11 6
19
1>
1C
b11 G
#40760000000
0!
0*
09
0>
0C
#40770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#40780000000
0!
0*
09
0>
0C
#40790000000
1!
1*
b101 6
19
1>
1C
b101 G
#40800000000
0!
0*
09
0>
0C
#40810000000
1!
1*
b110 6
19
1>
1C
b110 G
#40820000000
0!
0*
09
0>
0C
#40830000000
1!
1*
b111 6
19
1>
1C
b111 G
#40840000000
0!
1"
0*
1+
09
1:
0>
0C
#40850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#40860000000
0!
0*
09
0>
0C
#40870000000
1!
1*
b1 6
19
1>
1C
b1 G
#40880000000
0!
0*
09
0>
0C
#40890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#40900000000
0!
0*
09
0>
0C
#40910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#40920000000
0!
0*
09
0>
0C
#40930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#40940000000
0!
0*
09
0>
0C
#40950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#40960000000
0!
0#
0*
0,
09
0>
0?
0C
#40970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#40980000000
0!
0*
09
0>
0C
#40990000000
1!
1*
19
1>
1C
#41000000000
0!
0*
09
0>
0C
#41010000000
1!
1*
19
1>
1C
#41020000000
0!
0*
09
0>
0C
#41030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#41040000000
0!
0*
09
0>
0C
#41050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#41060000000
0!
0*
09
0>
0C
#41070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#41080000000
0!
0*
09
0>
0C
#41090000000
1!
1*
b10 6
19
1>
1C
b10 G
#41100000000
0!
0*
09
0>
0C
#41110000000
1!
1*
b11 6
19
1>
1C
b11 G
#41120000000
0!
0*
09
0>
0C
#41130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#41140000000
0!
0*
09
0>
0C
#41150000000
1!
1*
b101 6
19
1>
1C
b101 G
#41160000000
0!
0*
09
0>
0C
#41170000000
1!
1*
b110 6
19
1>
1C
b110 G
#41180000000
0!
0*
09
0>
0C
#41190000000
1!
1*
b111 6
19
1>
1C
b111 G
#41200000000
0!
0*
09
0>
0C
#41210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#41220000000
0!
0*
09
0>
0C
#41230000000
1!
1*
b1 6
19
1>
1C
b1 G
#41240000000
0!
0*
09
0>
0C
#41250000000
1!
1*
b10 6
19
1>
1C
b10 G
#41260000000
0!
0*
09
0>
0C
#41270000000
1!
1*
b11 6
19
1>
1C
b11 G
#41280000000
0!
0*
09
0>
0C
#41290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#41300000000
0!
0*
09
0>
0C
#41310000000
1!
1*
b101 6
19
1>
1C
b101 G
#41320000000
0!
0*
09
0>
0C
#41330000000
1!
1*
b110 6
19
1>
1C
b110 G
#41340000000
0!
0*
09
0>
0C
#41350000000
1!
1*
b111 6
19
1>
1C
b111 G
#41360000000
0!
0*
09
0>
0C
#41370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#41380000000
0!
0*
09
0>
0C
#41390000000
1!
1*
b1 6
19
1>
1C
b1 G
#41400000000
0!
0*
09
0>
0C
#41410000000
1!
1*
b10 6
19
1>
1C
b10 G
#41420000000
0!
0*
09
0>
0C
#41430000000
1!
1*
b11 6
19
1>
1C
b11 G
#41440000000
0!
0*
09
0>
0C
#41450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#41460000000
0!
0*
09
0>
0C
#41470000000
1!
1*
b101 6
19
1>
1C
b101 G
#41480000000
0!
0*
09
0>
0C
#41490000000
1!
1*
b110 6
19
1>
1C
b110 G
#41500000000
0!
0*
09
0>
0C
#41510000000
1!
1*
b111 6
19
1>
1C
b111 G
#41520000000
0!
1"
0*
1+
09
1:
0>
0C
#41530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#41540000000
0!
0*
09
0>
0C
#41550000000
1!
1*
b1 6
19
1>
1C
b1 G
#41560000000
0!
0*
09
0>
0C
#41570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#41580000000
0!
0*
09
0>
0C
#41590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#41600000000
0!
0*
09
0>
0C
#41610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#41620000000
0!
0*
09
0>
0C
#41630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#41640000000
0!
0#
0*
0,
09
0>
0?
0C
#41650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#41660000000
0!
0*
09
0>
0C
#41670000000
1!
1*
19
1>
1C
#41680000000
0!
0*
09
0>
0C
#41690000000
1!
1*
19
1>
1C
#41700000000
0!
0*
09
0>
0C
#41710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#41720000000
0!
0*
09
0>
0C
#41730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#41740000000
0!
0*
09
0>
0C
#41750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#41760000000
0!
0*
09
0>
0C
#41770000000
1!
1*
b10 6
19
1>
1C
b10 G
#41780000000
0!
0*
09
0>
0C
#41790000000
1!
1*
b11 6
19
1>
1C
b11 G
#41800000000
0!
0*
09
0>
0C
#41810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#41820000000
0!
0*
09
0>
0C
#41830000000
1!
1*
b101 6
19
1>
1C
b101 G
#41840000000
0!
0*
09
0>
0C
#41850000000
1!
1*
b110 6
19
1>
1C
b110 G
#41860000000
0!
0*
09
0>
0C
#41870000000
1!
1*
b111 6
19
1>
1C
b111 G
#41880000000
0!
0*
09
0>
0C
#41890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#41900000000
0!
0*
09
0>
0C
#41910000000
1!
1*
b1 6
19
1>
1C
b1 G
#41920000000
0!
0*
09
0>
0C
#41930000000
1!
1*
b10 6
19
1>
1C
b10 G
#41940000000
0!
0*
09
0>
0C
#41950000000
1!
1*
b11 6
19
1>
1C
b11 G
#41960000000
0!
0*
09
0>
0C
#41970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#41980000000
0!
0*
09
0>
0C
#41990000000
1!
1*
b101 6
19
1>
1C
b101 G
#42000000000
0!
0*
09
0>
0C
#42010000000
1!
1*
b110 6
19
1>
1C
b110 G
#42020000000
0!
0*
09
0>
0C
#42030000000
1!
1*
b111 6
19
1>
1C
b111 G
#42040000000
0!
0*
09
0>
0C
#42050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#42060000000
0!
0*
09
0>
0C
#42070000000
1!
1*
b1 6
19
1>
1C
b1 G
#42080000000
0!
0*
09
0>
0C
#42090000000
1!
1*
b10 6
19
1>
1C
b10 G
#42100000000
0!
0*
09
0>
0C
#42110000000
1!
1*
b11 6
19
1>
1C
b11 G
#42120000000
0!
0*
09
0>
0C
#42130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#42140000000
0!
0*
09
0>
0C
#42150000000
1!
1*
b101 6
19
1>
1C
b101 G
#42160000000
0!
0*
09
0>
0C
#42170000000
1!
1*
b110 6
19
1>
1C
b110 G
#42180000000
0!
0*
09
0>
0C
#42190000000
1!
1*
b111 6
19
1>
1C
b111 G
#42200000000
0!
1"
0*
1+
09
1:
0>
0C
#42210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#42220000000
0!
0*
09
0>
0C
#42230000000
1!
1*
b1 6
19
1>
1C
b1 G
#42240000000
0!
0*
09
0>
0C
#42250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#42260000000
0!
0*
09
0>
0C
#42270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#42280000000
0!
0*
09
0>
0C
#42290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#42300000000
0!
0*
09
0>
0C
#42310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#42320000000
0!
0#
0*
0,
09
0>
0?
0C
#42330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#42340000000
0!
0*
09
0>
0C
#42350000000
1!
1*
19
1>
1C
#42360000000
0!
0*
09
0>
0C
#42370000000
1!
1*
19
1>
1C
#42380000000
0!
0*
09
0>
0C
#42390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#42400000000
0!
0*
09
0>
0C
#42410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#42420000000
0!
0*
09
0>
0C
#42430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#42440000000
0!
0*
09
0>
0C
#42450000000
1!
1*
b10 6
19
1>
1C
b10 G
#42460000000
0!
0*
09
0>
0C
#42470000000
1!
1*
b11 6
19
1>
1C
b11 G
#42480000000
0!
0*
09
0>
0C
#42490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#42500000000
0!
0*
09
0>
0C
#42510000000
1!
1*
b101 6
19
1>
1C
b101 G
#42520000000
0!
0*
09
0>
0C
#42530000000
1!
1*
b110 6
19
1>
1C
b110 G
#42540000000
0!
0*
09
0>
0C
#42550000000
1!
1*
b111 6
19
1>
1C
b111 G
#42560000000
0!
0*
09
0>
0C
#42570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#42580000000
0!
0*
09
0>
0C
#42590000000
1!
1*
b1 6
19
1>
1C
b1 G
#42600000000
0!
0*
09
0>
0C
#42610000000
1!
1*
b10 6
19
1>
1C
b10 G
#42620000000
0!
0*
09
0>
0C
#42630000000
1!
1*
b11 6
19
1>
1C
b11 G
#42640000000
0!
0*
09
0>
0C
#42650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#42660000000
0!
0*
09
0>
0C
#42670000000
1!
1*
b101 6
19
1>
1C
b101 G
#42680000000
0!
0*
09
0>
0C
#42690000000
1!
1*
b110 6
19
1>
1C
b110 G
#42700000000
0!
0*
09
0>
0C
#42710000000
1!
1*
b111 6
19
1>
1C
b111 G
#42720000000
0!
0*
09
0>
0C
#42730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#42740000000
0!
0*
09
0>
0C
#42750000000
1!
1*
b1 6
19
1>
1C
b1 G
#42760000000
0!
0*
09
0>
0C
#42770000000
1!
1*
b10 6
19
1>
1C
b10 G
#42780000000
0!
0*
09
0>
0C
#42790000000
1!
1*
b11 6
19
1>
1C
b11 G
#42800000000
0!
0*
09
0>
0C
#42810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#42820000000
0!
0*
09
0>
0C
#42830000000
1!
1*
b101 6
19
1>
1C
b101 G
#42840000000
0!
0*
09
0>
0C
#42850000000
1!
1*
b110 6
19
1>
1C
b110 G
#42860000000
0!
0*
09
0>
0C
#42870000000
1!
1*
b111 6
19
1>
1C
b111 G
#42880000000
0!
1"
0*
1+
09
1:
0>
0C
#42890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#42900000000
0!
0*
09
0>
0C
#42910000000
1!
1*
b1 6
19
1>
1C
b1 G
#42920000000
0!
0*
09
0>
0C
#42930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#42940000000
0!
0*
09
0>
0C
#42950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#42960000000
0!
0*
09
0>
0C
#42970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#42980000000
0!
0*
09
0>
0C
#42990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#43000000000
0!
0#
0*
0,
09
0>
0?
0C
#43010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#43020000000
0!
0*
09
0>
0C
#43030000000
1!
1*
19
1>
1C
#43040000000
0!
0*
09
0>
0C
#43050000000
1!
1*
19
1>
1C
#43060000000
0!
0*
09
0>
0C
#43070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#43080000000
0!
0*
09
0>
0C
#43090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#43100000000
0!
0*
09
0>
0C
#43110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#43120000000
0!
0*
09
0>
0C
#43130000000
1!
1*
b10 6
19
1>
1C
b10 G
#43140000000
0!
0*
09
0>
0C
#43150000000
1!
1*
b11 6
19
1>
1C
b11 G
#43160000000
0!
0*
09
0>
0C
#43170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#43180000000
0!
0*
09
0>
0C
#43190000000
1!
1*
b101 6
19
1>
1C
b101 G
#43200000000
0!
0*
09
0>
0C
#43210000000
1!
1*
b110 6
19
1>
1C
b110 G
#43220000000
0!
0*
09
0>
0C
#43230000000
1!
1*
b111 6
19
1>
1C
b111 G
#43240000000
0!
0*
09
0>
0C
#43250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#43260000000
0!
0*
09
0>
0C
#43270000000
1!
1*
b1 6
19
1>
1C
b1 G
#43280000000
0!
0*
09
0>
0C
#43290000000
1!
1*
b10 6
19
1>
1C
b10 G
#43300000000
0!
0*
09
0>
0C
#43310000000
1!
1*
b11 6
19
1>
1C
b11 G
#43320000000
0!
0*
09
0>
0C
#43330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#43340000000
0!
0*
09
0>
0C
#43350000000
1!
1*
b101 6
19
1>
1C
b101 G
#43360000000
0!
0*
09
0>
0C
#43370000000
1!
1*
b110 6
19
1>
1C
b110 G
#43380000000
0!
0*
09
0>
0C
#43390000000
1!
1*
b111 6
19
1>
1C
b111 G
#43400000000
0!
0*
09
0>
0C
#43410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#43420000000
0!
0*
09
0>
0C
#43430000000
1!
1*
b1 6
19
1>
1C
b1 G
#43440000000
0!
0*
09
0>
0C
#43450000000
1!
1*
b10 6
19
1>
1C
b10 G
#43460000000
0!
0*
09
0>
0C
#43470000000
1!
1*
b11 6
19
1>
1C
b11 G
#43480000000
0!
0*
09
0>
0C
#43490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#43500000000
0!
0*
09
0>
0C
#43510000000
1!
1*
b101 6
19
1>
1C
b101 G
#43520000000
0!
0*
09
0>
0C
#43530000000
1!
1*
b110 6
19
1>
1C
b110 G
#43540000000
0!
0*
09
0>
0C
#43550000000
1!
1*
b111 6
19
1>
1C
b111 G
#43560000000
0!
1"
0*
1+
09
1:
0>
0C
#43570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#43580000000
0!
0*
09
0>
0C
#43590000000
1!
1*
b1 6
19
1>
1C
b1 G
#43600000000
0!
0*
09
0>
0C
#43610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#43620000000
0!
0*
09
0>
0C
#43630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#43640000000
0!
0*
09
0>
0C
#43650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#43660000000
0!
0*
09
0>
0C
#43670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#43680000000
0!
0#
0*
0,
09
0>
0?
0C
#43690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#43700000000
0!
0*
09
0>
0C
#43710000000
1!
1*
19
1>
1C
#43720000000
0!
0*
09
0>
0C
#43730000000
1!
1*
19
1>
1C
#43740000000
0!
0*
09
0>
0C
#43750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#43760000000
0!
0*
09
0>
0C
#43770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#43780000000
0!
0*
09
0>
0C
#43790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#43800000000
0!
0*
09
0>
0C
#43810000000
1!
1*
b10 6
19
1>
1C
b10 G
#43820000000
0!
0*
09
0>
0C
#43830000000
1!
1*
b11 6
19
1>
1C
b11 G
#43840000000
0!
0*
09
0>
0C
#43850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#43860000000
0!
0*
09
0>
0C
#43870000000
1!
1*
b101 6
19
1>
1C
b101 G
#43880000000
0!
0*
09
0>
0C
#43890000000
1!
1*
b110 6
19
1>
1C
b110 G
#43900000000
0!
0*
09
0>
0C
#43910000000
1!
1*
b111 6
19
1>
1C
b111 G
#43920000000
0!
0*
09
0>
0C
#43930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#43940000000
0!
0*
09
0>
0C
#43950000000
1!
1*
b1 6
19
1>
1C
b1 G
#43960000000
0!
0*
09
0>
0C
#43970000000
1!
1*
b10 6
19
1>
1C
b10 G
#43980000000
0!
0*
09
0>
0C
#43990000000
1!
1*
b11 6
19
1>
1C
b11 G
#44000000000
0!
0*
09
0>
0C
#44010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#44020000000
0!
0*
09
0>
0C
#44030000000
1!
1*
b101 6
19
1>
1C
b101 G
#44040000000
0!
0*
09
0>
0C
#44050000000
1!
1*
b110 6
19
1>
1C
b110 G
#44060000000
0!
0*
09
0>
0C
#44070000000
1!
1*
b111 6
19
1>
1C
b111 G
#44080000000
0!
0*
09
0>
0C
#44090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#44100000000
0!
0*
09
0>
0C
#44110000000
1!
1*
b1 6
19
1>
1C
b1 G
#44120000000
0!
0*
09
0>
0C
#44130000000
1!
1*
b10 6
19
1>
1C
b10 G
#44140000000
0!
0*
09
0>
0C
#44150000000
1!
1*
b11 6
19
1>
1C
b11 G
#44160000000
0!
0*
09
0>
0C
#44170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#44180000000
0!
0*
09
0>
0C
#44190000000
1!
1*
b101 6
19
1>
1C
b101 G
#44200000000
0!
0*
09
0>
0C
#44210000000
1!
1*
b110 6
19
1>
1C
b110 G
#44220000000
0!
0*
09
0>
0C
#44230000000
1!
1*
b111 6
19
1>
1C
b111 G
#44240000000
0!
1"
0*
1+
09
1:
0>
0C
#44250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#44260000000
0!
0*
09
0>
0C
#44270000000
1!
1*
b1 6
19
1>
1C
b1 G
#44280000000
0!
0*
09
0>
0C
#44290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#44300000000
0!
0*
09
0>
0C
#44310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#44320000000
0!
0*
09
0>
0C
#44330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#44340000000
0!
0*
09
0>
0C
#44350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#44360000000
0!
0#
0*
0,
09
0>
0?
0C
#44370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#44380000000
0!
0*
09
0>
0C
#44390000000
1!
1*
19
1>
1C
#44400000000
0!
0*
09
0>
0C
#44410000000
1!
1*
19
1>
1C
#44420000000
0!
0*
09
0>
0C
#44430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#44440000000
0!
0*
09
0>
0C
#44450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#44460000000
0!
0*
09
0>
0C
#44470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#44480000000
0!
0*
09
0>
0C
#44490000000
1!
1*
b10 6
19
1>
1C
b10 G
#44500000000
0!
0*
09
0>
0C
#44510000000
1!
1*
b11 6
19
1>
1C
b11 G
#44520000000
0!
0*
09
0>
0C
#44530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#44540000000
0!
0*
09
0>
0C
#44550000000
1!
1*
b101 6
19
1>
1C
b101 G
#44560000000
0!
0*
09
0>
0C
#44570000000
1!
1*
b110 6
19
1>
1C
b110 G
#44580000000
0!
0*
09
0>
0C
#44590000000
1!
1*
b111 6
19
1>
1C
b111 G
#44600000000
0!
0*
09
0>
0C
#44610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#44620000000
0!
0*
09
0>
0C
#44630000000
1!
1*
b1 6
19
1>
1C
b1 G
#44640000000
0!
0*
09
0>
0C
#44650000000
1!
1*
b10 6
19
1>
1C
b10 G
#44660000000
0!
0*
09
0>
0C
#44670000000
1!
1*
b11 6
19
1>
1C
b11 G
#44680000000
0!
0*
09
0>
0C
#44690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#44700000000
0!
0*
09
0>
0C
#44710000000
1!
1*
b101 6
19
1>
1C
b101 G
#44720000000
0!
0*
09
0>
0C
#44730000000
1!
1*
b110 6
19
1>
1C
b110 G
#44740000000
0!
0*
09
0>
0C
#44750000000
1!
1*
b111 6
19
1>
1C
b111 G
#44760000000
0!
0*
09
0>
0C
#44770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#44780000000
0!
0*
09
0>
0C
#44790000000
1!
1*
b1 6
19
1>
1C
b1 G
#44800000000
0!
0*
09
0>
0C
#44810000000
1!
1*
b10 6
19
1>
1C
b10 G
#44820000000
0!
0*
09
0>
0C
#44830000000
1!
1*
b11 6
19
1>
1C
b11 G
#44840000000
0!
0*
09
0>
0C
#44850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#44860000000
0!
0*
09
0>
0C
#44870000000
1!
1*
b101 6
19
1>
1C
b101 G
#44880000000
0!
0*
09
0>
0C
#44890000000
1!
1*
b110 6
19
1>
1C
b110 G
#44900000000
0!
0*
09
0>
0C
#44910000000
1!
1*
b111 6
19
1>
1C
b111 G
#44920000000
0!
1"
0*
1+
09
1:
0>
0C
#44930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#44940000000
0!
0*
09
0>
0C
#44950000000
1!
1*
b1 6
19
1>
1C
b1 G
#44960000000
0!
0*
09
0>
0C
#44970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#44980000000
0!
0*
09
0>
0C
#44990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#45000000000
0!
0*
09
0>
0C
#45010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#45020000000
0!
0*
09
0>
0C
#45030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#45040000000
0!
0#
0*
0,
09
0>
0?
0C
#45050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#45060000000
0!
0*
09
0>
0C
#45070000000
1!
1*
19
1>
1C
#45080000000
0!
0*
09
0>
0C
#45090000000
1!
1*
19
1>
1C
#45100000000
0!
0*
09
0>
0C
#45110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#45120000000
0!
0*
09
0>
0C
#45130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#45140000000
0!
0*
09
0>
0C
#45150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#45160000000
0!
0*
09
0>
0C
#45170000000
1!
1*
b10 6
19
1>
1C
b10 G
#45180000000
0!
0*
09
0>
0C
#45190000000
1!
1*
b11 6
19
1>
1C
b11 G
#45200000000
0!
0*
09
0>
0C
#45210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#45220000000
0!
0*
09
0>
0C
#45230000000
1!
1*
b101 6
19
1>
1C
b101 G
#45240000000
0!
0*
09
0>
0C
#45250000000
1!
1*
b110 6
19
1>
1C
b110 G
#45260000000
0!
0*
09
0>
0C
#45270000000
1!
1*
b111 6
19
1>
1C
b111 G
#45280000000
0!
0*
09
0>
0C
#45290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#45300000000
0!
0*
09
0>
0C
#45310000000
1!
1*
b1 6
19
1>
1C
b1 G
#45320000000
0!
0*
09
0>
0C
#45330000000
1!
1*
b10 6
19
1>
1C
b10 G
#45340000000
0!
0*
09
0>
0C
#45350000000
1!
1*
b11 6
19
1>
1C
b11 G
#45360000000
0!
0*
09
0>
0C
#45370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#45380000000
0!
0*
09
0>
0C
#45390000000
1!
1*
b101 6
19
1>
1C
b101 G
#45400000000
0!
0*
09
0>
0C
#45410000000
1!
1*
b110 6
19
1>
1C
b110 G
#45420000000
0!
0*
09
0>
0C
#45430000000
1!
1*
b111 6
19
1>
1C
b111 G
#45440000000
0!
0*
09
0>
0C
#45450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#45460000000
0!
0*
09
0>
0C
#45470000000
1!
1*
b1 6
19
1>
1C
b1 G
#45480000000
0!
0*
09
0>
0C
#45490000000
1!
1*
b10 6
19
1>
1C
b10 G
#45500000000
0!
0*
09
0>
0C
#45510000000
1!
1*
b11 6
19
1>
1C
b11 G
#45520000000
0!
0*
09
0>
0C
#45530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#45540000000
0!
0*
09
0>
0C
#45550000000
1!
1*
b101 6
19
1>
1C
b101 G
#45560000000
0!
0*
09
0>
0C
#45570000000
1!
1*
b110 6
19
1>
1C
b110 G
#45580000000
0!
0*
09
0>
0C
#45590000000
1!
1*
b111 6
19
1>
1C
b111 G
#45600000000
0!
1"
0*
1+
09
1:
0>
0C
#45610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#45620000000
0!
0*
09
0>
0C
#45630000000
1!
1*
b1 6
19
1>
1C
b1 G
#45640000000
0!
0*
09
0>
0C
#45650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#45660000000
0!
0*
09
0>
0C
#45670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#45680000000
0!
0*
09
0>
0C
#45690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#45700000000
0!
0*
09
0>
0C
#45710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#45720000000
0!
0#
0*
0,
09
0>
0?
0C
#45730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#45740000000
0!
0*
09
0>
0C
#45750000000
1!
1*
19
1>
1C
#45760000000
0!
0*
09
0>
0C
#45770000000
1!
1*
19
1>
1C
#45780000000
0!
0*
09
0>
0C
#45790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#45800000000
0!
0*
09
0>
0C
#45810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#45820000000
0!
0*
09
0>
0C
#45830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#45840000000
0!
0*
09
0>
0C
#45850000000
1!
1*
b10 6
19
1>
1C
b10 G
#45860000000
0!
0*
09
0>
0C
#45870000000
1!
1*
b11 6
19
1>
1C
b11 G
#45880000000
0!
0*
09
0>
0C
#45890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#45900000000
0!
0*
09
0>
0C
#45910000000
1!
1*
b101 6
19
1>
1C
b101 G
#45920000000
0!
0*
09
0>
0C
#45930000000
1!
1*
b110 6
19
1>
1C
b110 G
#45940000000
0!
0*
09
0>
0C
#45950000000
1!
1*
b111 6
19
1>
1C
b111 G
#45960000000
0!
0*
09
0>
0C
#45970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#45980000000
0!
0*
09
0>
0C
#45990000000
1!
1*
b1 6
19
1>
1C
b1 G
#46000000000
0!
0*
09
0>
0C
#46010000000
1!
1*
b10 6
19
1>
1C
b10 G
#46020000000
0!
0*
09
0>
0C
#46030000000
1!
1*
b11 6
19
1>
1C
b11 G
#46040000000
0!
0*
09
0>
0C
#46050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#46060000000
0!
0*
09
0>
0C
#46070000000
1!
1*
b101 6
19
1>
1C
b101 G
#46080000000
0!
0*
09
0>
0C
#46090000000
1!
1*
b110 6
19
1>
1C
b110 G
#46100000000
0!
0*
09
0>
0C
#46110000000
1!
1*
b111 6
19
1>
1C
b111 G
#46120000000
0!
0*
09
0>
0C
#46130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#46140000000
0!
0*
09
0>
0C
#46150000000
1!
1*
b1 6
19
1>
1C
b1 G
#46160000000
0!
0*
09
0>
0C
#46170000000
1!
1*
b10 6
19
1>
1C
b10 G
#46180000000
0!
0*
09
0>
0C
#46190000000
1!
1*
b11 6
19
1>
1C
b11 G
#46200000000
0!
0*
09
0>
0C
#46210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#46220000000
0!
0*
09
0>
0C
#46230000000
1!
1*
b101 6
19
1>
1C
b101 G
#46240000000
0!
0*
09
0>
0C
#46250000000
1!
1*
b110 6
19
1>
1C
b110 G
#46260000000
0!
0*
09
0>
0C
#46270000000
1!
1*
b111 6
19
1>
1C
b111 G
#46280000000
0!
1"
0*
1+
09
1:
0>
0C
#46290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#46300000000
0!
0*
09
0>
0C
#46310000000
1!
1*
b1 6
19
1>
1C
b1 G
#46320000000
0!
0*
09
0>
0C
#46330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#46340000000
0!
0*
09
0>
0C
#46350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#46360000000
0!
0*
09
0>
0C
#46370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#46380000000
0!
0*
09
0>
0C
#46390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#46400000000
0!
0#
0*
0,
09
0>
0?
0C
#46410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#46420000000
0!
0*
09
0>
0C
#46430000000
1!
1*
19
1>
1C
#46440000000
0!
0*
09
0>
0C
#46450000000
1!
1*
19
1>
1C
#46460000000
0!
0*
09
0>
0C
#46470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#46480000000
0!
0*
09
0>
0C
#46490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#46500000000
0!
0*
09
0>
0C
#46510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#46520000000
0!
0*
09
0>
0C
#46530000000
1!
1*
b10 6
19
1>
1C
b10 G
#46540000000
0!
0*
09
0>
0C
#46550000000
1!
1*
b11 6
19
1>
1C
b11 G
#46560000000
0!
0*
09
0>
0C
#46570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#46580000000
0!
0*
09
0>
0C
#46590000000
1!
1*
b101 6
19
1>
1C
b101 G
#46600000000
0!
0*
09
0>
0C
#46610000000
1!
1*
b110 6
19
1>
1C
b110 G
#46620000000
0!
0*
09
0>
0C
#46630000000
1!
1*
b111 6
19
1>
1C
b111 G
#46640000000
0!
0*
09
0>
0C
#46650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#46660000000
0!
0*
09
0>
0C
#46670000000
1!
1*
b1 6
19
1>
1C
b1 G
#46680000000
0!
0*
09
0>
0C
#46690000000
1!
1*
b10 6
19
1>
1C
b10 G
#46700000000
0!
0*
09
0>
0C
#46710000000
1!
1*
b11 6
19
1>
1C
b11 G
#46720000000
0!
0*
09
0>
0C
#46730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#46740000000
0!
0*
09
0>
0C
#46750000000
1!
1*
b101 6
19
1>
1C
b101 G
#46760000000
0!
0*
09
0>
0C
#46770000000
1!
1*
b110 6
19
1>
1C
b110 G
#46780000000
0!
0*
09
0>
0C
#46790000000
1!
1*
b111 6
19
1>
1C
b111 G
#46800000000
0!
0*
09
0>
0C
#46810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#46820000000
0!
0*
09
0>
0C
#46830000000
1!
1*
b1 6
19
1>
1C
b1 G
#46840000000
0!
0*
09
0>
0C
#46850000000
1!
1*
b10 6
19
1>
1C
b10 G
#46860000000
0!
0*
09
0>
0C
#46870000000
1!
1*
b11 6
19
1>
1C
b11 G
#46880000000
0!
0*
09
0>
0C
#46890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#46900000000
0!
0*
09
0>
0C
#46910000000
1!
1*
b101 6
19
1>
1C
b101 G
#46920000000
0!
0*
09
0>
0C
#46930000000
1!
1*
b110 6
19
1>
1C
b110 G
#46940000000
0!
0*
09
0>
0C
#46950000000
1!
1*
b111 6
19
1>
1C
b111 G
#46960000000
0!
1"
0*
1+
09
1:
0>
0C
#46970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#46980000000
0!
0*
09
0>
0C
#46990000000
1!
1*
b1 6
19
1>
1C
b1 G
#47000000000
0!
0*
09
0>
0C
#47010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#47020000000
0!
0*
09
0>
0C
#47030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#47040000000
0!
0*
09
0>
0C
#47050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#47060000000
0!
0*
09
0>
0C
#47070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#47080000000
0!
0#
0*
0,
09
0>
0?
0C
#47090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#47100000000
0!
0*
09
0>
0C
#47110000000
1!
1*
19
1>
1C
#47120000000
0!
0*
09
0>
0C
#47130000000
1!
1*
19
1>
1C
#47140000000
0!
0*
09
0>
0C
#47150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#47160000000
0!
0*
09
0>
0C
#47170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#47180000000
0!
0*
09
0>
0C
#47190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#47200000000
0!
0*
09
0>
0C
#47210000000
1!
1*
b10 6
19
1>
1C
b10 G
#47220000000
0!
0*
09
0>
0C
#47230000000
1!
1*
b11 6
19
1>
1C
b11 G
#47240000000
0!
0*
09
0>
0C
#47250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#47260000000
0!
0*
09
0>
0C
#47270000000
1!
1*
b101 6
19
1>
1C
b101 G
#47280000000
0!
0*
09
0>
0C
#47290000000
1!
1*
b110 6
19
1>
1C
b110 G
#47300000000
0!
0*
09
0>
0C
#47310000000
1!
1*
b111 6
19
1>
1C
b111 G
#47320000000
0!
0*
09
0>
0C
#47330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#47340000000
0!
0*
09
0>
0C
#47350000000
1!
1*
b1 6
19
1>
1C
b1 G
#47360000000
0!
0*
09
0>
0C
#47370000000
1!
1*
b10 6
19
1>
1C
b10 G
#47380000000
0!
0*
09
0>
0C
#47390000000
1!
1*
b11 6
19
1>
1C
b11 G
#47400000000
0!
0*
09
0>
0C
#47410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#47420000000
0!
0*
09
0>
0C
#47430000000
1!
1*
b101 6
19
1>
1C
b101 G
#47440000000
0!
0*
09
0>
0C
#47450000000
1!
1*
b110 6
19
1>
1C
b110 G
#47460000000
0!
0*
09
0>
0C
#47470000000
1!
1*
b111 6
19
1>
1C
b111 G
#47480000000
0!
0*
09
0>
0C
#47490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#47500000000
0!
0*
09
0>
0C
#47510000000
1!
1*
b1 6
19
1>
1C
b1 G
#47520000000
0!
0*
09
0>
0C
#47530000000
1!
1*
b10 6
19
1>
1C
b10 G
#47540000000
0!
0*
09
0>
0C
#47550000000
1!
1*
b11 6
19
1>
1C
b11 G
#47560000000
0!
0*
09
0>
0C
#47570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#47580000000
0!
0*
09
0>
0C
#47590000000
1!
1*
b101 6
19
1>
1C
b101 G
#47600000000
0!
0*
09
0>
0C
#47610000000
1!
1*
b110 6
19
1>
1C
b110 G
#47620000000
0!
0*
09
0>
0C
#47630000000
1!
1*
b111 6
19
1>
1C
b111 G
#47640000000
0!
1"
0*
1+
09
1:
0>
0C
#47650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#47660000000
0!
0*
09
0>
0C
#47670000000
1!
1*
b1 6
19
1>
1C
b1 G
#47680000000
0!
0*
09
0>
0C
#47690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#47700000000
0!
0*
09
0>
0C
#47710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#47720000000
0!
0*
09
0>
0C
#47730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#47740000000
0!
0*
09
0>
0C
#47750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#47760000000
0!
0#
0*
0,
09
0>
0?
0C
#47770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#47780000000
0!
0*
09
0>
0C
#47790000000
1!
1*
19
1>
1C
#47800000000
0!
0*
09
0>
0C
#47810000000
1!
1*
19
1>
1C
#47820000000
0!
0*
09
0>
0C
#47830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#47840000000
0!
0*
09
0>
0C
#47850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#47860000000
0!
0*
09
0>
0C
#47870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#47880000000
0!
0*
09
0>
0C
#47890000000
1!
1*
b10 6
19
1>
1C
b10 G
#47900000000
0!
0*
09
0>
0C
#47910000000
1!
1*
b11 6
19
1>
1C
b11 G
#47920000000
0!
0*
09
0>
0C
#47930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#47940000000
0!
0*
09
0>
0C
#47950000000
1!
1*
b101 6
19
1>
1C
b101 G
#47960000000
0!
0*
09
0>
0C
#47970000000
1!
1*
b110 6
19
1>
1C
b110 G
#47980000000
0!
0*
09
0>
0C
#47990000000
1!
1*
b111 6
19
1>
1C
b111 G
#48000000000
0!
0*
09
0>
0C
#48010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#48020000000
0!
0*
09
0>
0C
#48030000000
1!
1*
b1 6
19
1>
1C
b1 G
#48040000000
0!
0*
09
0>
0C
#48050000000
1!
1*
b10 6
19
1>
1C
b10 G
#48060000000
0!
0*
09
0>
0C
#48070000000
1!
1*
b11 6
19
1>
1C
b11 G
#48080000000
0!
0*
09
0>
0C
#48090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#48100000000
0!
0*
09
0>
0C
#48110000000
1!
1*
b101 6
19
1>
1C
b101 G
#48120000000
0!
0*
09
0>
0C
#48130000000
1!
1*
b110 6
19
1>
1C
b110 G
#48140000000
0!
0*
09
0>
0C
#48150000000
1!
1*
b111 6
19
1>
1C
b111 G
#48160000000
0!
0*
09
0>
0C
#48170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#48180000000
0!
0*
09
0>
0C
#48190000000
1!
1*
b1 6
19
1>
1C
b1 G
#48200000000
0!
0*
09
0>
0C
#48210000000
1!
1*
b10 6
19
1>
1C
b10 G
#48220000000
0!
0*
09
0>
0C
#48230000000
1!
1*
b11 6
19
1>
1C
b11 G
#48240000000
0!
0*
09
0>
0C
#48250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#48260000000
0!
0*
09
0>
0C
#48270000000
1!
1*
b101 6
19
1>
1C
b101 G
#48280000000
0!
0*
09
0>
0C
#48290000000
1!
1*
b110 6
19
1>
1C
b110 G
#48300000000
0!
0*
09
0>
0C
#48310000000
1!
1*
b111 6
19
1>
1C
b111 G
#48320000000
0!
1"
0*
1+
09
1:
0>
0C
#48330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#48340000000
0!
0*
09
0>
0C
#48350000000
1!
1*
b1 6
19
1>
1C
b1 G
#48360000000
0!
0*
09
0>
0C
#48370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#48380000000
0!
0*
09
0>
0C
#48390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#48400000000
0!
0*
09
0>
0C
#48410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#48420000000
0!
0*
09
0>
0C
#48430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#48440000000
0!
0#
0*
0,
09
0>
0?
0C
#48450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#48460000000
0!
0*
09
0>
0C
#48470000000
1!
1*
19
1>
1C
#48480000000
0!
0*
09
0>
0C
#48490000000
1!
1*
19
1>
1C
#48500000000
0!
0*
09
0>
0C
#48510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#48520000000
0!
0*
09
0>
0C
#48530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#48540000000
0!
0*
09
0>
0C
#48550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#48560000000
0!
0*
09
0>
0C
#48570000000
1!
1*
b10 6
19
1>
1C
b10 G
#48580000000
0!
0*
09
0>
0C
#48590000000
1!
1*
b11 6
19
1>
1C
b11 G
#48600000000
0!
0*
09
0>
0C
#48610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#48620000000
0!
0*
09
0>
0C
#48630000000
1!
1*
b101 6
19
1>
1C
b101 G
#48640000000
0!
0*
09
0>
0C
#48650000000
1!
1*
b110 6
19
1>
1C
b110 G
#48660000000
0!
0*
09
0>
0C
#48670000000
1!
1*
b111 6
19
1>
1C
b111 G
#48680000000
0!
0*
09
0>
0C
#48690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#48700000000
0!
0*
09
0>
0C
#48710000000
1!
1*
b1 6
19
1>
1C
b1 G
#48720000000
0!
0*
09
0>
0C
#48730000000
1!
1*
b10 6
19
1>
1C
b10 G
#48740000000
0!
0*
09
0>
0C
#48750000000
1!
1*
b11 6
19
1>
1C
b11 G
#48760000000
0!
0*
09
0>
0C
#48770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#48780000000
0!
0*
09
0>
0C
#48790000000
1!
1*
b101 6
19
1>
1C
b101 G
#48800000000
0!
0*
09
0>
0C
#48810000000
1!
1*
b110 6
19
1>
1C
b110 G
#48820000000
0!
0*
09
0>
0C
#48830000000
1!
1*
b111 6
19
1>
1C
b111 G
#48840000000
0!
0*
09
0>
0C
#48850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#48860000000
0!
0*
09
0>
0C
#48870000000
1!
1*
b1 6
19
1>
1C
b1 G
#48880000000
0!
0*
09
0>
0C
#48890000000
1!
1*
b10 6
19
1>
1C
b10 G
#48900000000
0!
0*
09
0>
0C
#48910000000
1!
1*
b11 6
19
1>
1C
b11 G
#48920000000
0!
0*
09
0>
0C
#48930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#48940000000
0!
0*
09
0>
0C
#48950000000
1!
1*
b101 6
19
1>
1C
b101 G
#48960000000
0!
0*
09
0>
0C
#48970000000
1!
1*
b110 6
19
1>
1C
b110 G
#48980000000
0!
0*
09
0>
0C
#48990000000
1!
1*
b111 6
19
1>
1C
b111 G
#49000000000
0!
1"
0*
1+
09
1:
0>
0C
#49010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#49020000000
0!
0*
09
0>
0C
#49030000000
1!
1*
b1 6
19
1>
1C
b1 G
#49040000000
0!
0*
09
0>
0C
#49050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#49060000000
0!
0*
09
0>
0C
#49070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#49080000000
0!
0*
09
0>
0C
#49090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#49100000000
0!
0*
09
0>
0C
#49110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#49120000000
0!
0#
0*
0,
09
0>
0?
0C
#49130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#49140000000
0!
0*
09
0>
0C
#49150000000
1!
1*
19
1>
1C
#49160000000
0!
0*
09
0>
0C
#49170000000
1!
1*
19
1>
1C
#49180000000
0!
0*
09
0>
0C
#49190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#49200000000
0!
0*
09
0>
0C
#49210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#49220000000
0!
0*
09
0>
0C
#49230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#49240000000
0!
0*
09
0>
0C
#49250000000
1!
1*
b10 6
19
1>
1C
b10 G
#49260000000
0!
0*
09
0>
0C
#49270000000
1!
1*
b11 6
19
1>
1C
b11 G
#49280000000
0!
0*
09
0>
0C
#49290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#49300000000
0!
0*
09
0>
0C
#49310000000
1!
1*
b101 6
19
1>
1C
b101 G
#49320000000
0!
0*
09
0>
0C
#49330000000
1!
1*
b110 6
19
1>
1C
b110 G
#49340000000
0!
0*
09
0>
0C
#49350000000
1!
1*
b111 6
19
1>
1C
b111 G
#49360000000
0!
0*
09
0>
0C
#49370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#49380000000
0!
0*
09
0>
0C
#49390000000
1!
1*
b1 6
19
1>
1C
b1 G
#49400000000
0!
0*
09
0>
0C
#49410000000
1!
1*
b10 6
19
1>
1C
b10 G
#49420000000
0!
0*
09
0>
0C
#49430000000
1!
1*
b11 6
19
1>
1C
b11 G
#49440000000
0!
0*
09
0>
0C
#49450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#49460000000
0!
0*
09
0>
0C
#49470000000
1!
1*
b101 6
19
1>
1C
b101 G
#49480000000
0!
0*
09
0>
0C
#49490000000
1!
1*
b110 6
19
1>
1C
b110 G
#49500000000
0!
0*
09
0>
0C
#49510000000
1!
1*
b111 6
19
1>
1C
b111 G
#49520000000
0!
0*
09
0>
0C
#49530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#49540000000
0!
0*
09
0>
0C
#49550000000
1!
1*
b1 6
19
1>
1C
b1 G
#49560000000
0!
0*
09
0>
0C
#49570000000
1!
1*
b10 6
19
1>
1C
b10 G
#49580000000
0!
0*
09
0>
0C
#49590000000
1!
1*
b11 6
19
1>
1C
b11 G
#49600000000
0!
0*
09
0>
0C
#49610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#49620000000
0!
0*
09
0>
0C
#49630000000
1!
1*
b101 6
19
1>
1C
b101 G
#49640000000
0!
0*
09
0>
0C
#49650000000
1!
1*
b110 6
19
1>
1C
b110 G
#49660000000
0!
0*
09
0>
0C
#49670000000
1!
1*
b111 6
19
1>
1C
b111 G
#49680000000
0!
1"
0*
1+
09
1:
0>
0C
#49690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#49700000000
0!
0*
09
0>
0C
#49710000000
1!
1*
b1 6
19
1>
1C
b1 G
#49720000000
0!
0*
09
0>
0C
#49730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#49740000000
0!
0*
09
0>
0C
#49750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#49760000000
0!
0*
09
0>
0C
#49770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#49780000000
0!
0*
09
0>
0C
#49790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#49800000000
0!
0#
0*
0,
09
0>
0?
0C
#49810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#49820000000
0!
0*
09
0>
0C
#49830000000
1!
1*
19
1>
1C
#49840000000
0!
0*
09
0>
0C
#49850000000
1!
1*
19
1>
1C
#49860000000
0!
0*
09
0>
0C
#49870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#49880000000
0!
0*
09
0>
0C
#49890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#49900000000
0!
0*
09
0>
0C
#49910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#49920000000
0!
0*
09
0>
0C
#49930000000
1!
1*
b10 6
19
1>
1C
b10 G
#49940000000
0!
0*
09
0>
0C
#49950000000
1!
1*
b11 6
19
1>
1C
b11 G
#49960000000
0!
0*
09
0>
0C
#49970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#49980000000
0!
0*
09
0>
0C
#49990000000
1!
1*
b101 6
19
1>
1C
b101 G
#50000000000
0!
0*
09
0>
0C
#50010000000
1!
1*
b110 6
19
1>
1C
b110 G
#50020000000
0!
0*
09
0>
0C
#50030000000
1!
1*
b111 6
19
1>
1C
b111 G
#50040000000
0!
0*
09
0>
0C
#50050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#50060000000
0!
0*
09
0>
0C
#50070000000
1!
1*
b1 6
19
1>
1C
b1 G
#50080000000
0!
0*
09
0>
0C
#50090000000
1!
1*
b10 6
19
1>
1C
b10 G
#50100000000
0!
0*
09
0>
0C
#50110000000
1!
1*
b11 6
19
1>
1C
b11 G
#50120000000
0!
0*
09
0>
0C
#50130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#50140000000
0!
0*
09
0>
0C
#50150000000
1!
1*
b101 6
19
1>
1C
b101 G
#50160000000
0!
0*
09
0>
0C
#50170000000
1!
1*
b110 6
19
1>
1C
b110 G
#50180000000
0!
0*
09
0>
0C
#50190000000
1!
1*
b111 6
19
1>
1C
b111 G
#50200000000
0!
0*
09
0>
0C
#50210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#50220000000
0!
0*
09
0>
0C
#50230000000
1!
1*
b1 6
19
1>
1C
b1 G
#50240000000
0!
0*
09
0>
0C
#50250000000
1!
1*
b10 6
19
1>
1C
b10 G
#50260000000
0!
0*
09
0>
0C
#50270000000
1!
1*
b11 6
19
1>
1C
b11 G
#50280000000
0!
0*
09
0>
0C
#50290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#50300000000
0!
0*
09
0>
0C
#50310000000
1!
1*
b101 6
19
1>
1C
b101 G
#50320000000
0!
0*
09
0>
0C
#50330000000
1!
1*
b110 6
19
1>
1C
b110 G
#50340000000
0!
0*
09
0>
0C
#50350000000
1!
1*
b111 6
19
1>
1C
b111 G
#50360000000
0!
1"
0*
1+
09
1:
0>
0C
#50370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#50380000000
0!
0*
09
0>
0C
#50390000000
1!
1*
b1 6
19
1>
1C
b1 G
#50400000000
0!
0*
09
0>
0C
#50410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#50420000000
0!
0*
09
0>
0C
#50430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#50440000000
0!
0*
09
0>
0C
#50450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#50460000000
0!
0*
09
0>
0C
#50470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#50480000000
0!
0#
0*
0,
09
0>
0?
0C
#50490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#50500000000
0!
0*
09
0>
0C
#50510000000
1!
1*
19
1>
1C
#50520000000
0!
0*
09
0>
0C
#50530000000
1!
1*
19
1>
1C
#50540000000
0!
0*
09
0>
0C
#50550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#50560000000
0!
0*
09
0>
0C
#50570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#50580000000
0!
0*
09
0>
0C
#50590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#50600000000
0!
0*
09
0>
0C
#50610000000
1!
1*
b10 6
19
1>
1C
b10 G
#50620000000
0!
0*
09
0>
0C
#50630000000
1!
1*
b11 6
19
1>
1C
b11 G
#50640000000
0!
0*
09
0>
0C
#50650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#50660000000
0!
0*
09
0>
0C
#50670000000
1!
1*
b101 6
19
1>
1C
b101 G
#50680000000
0!
0*
09
0>
0C
#50690000000
1!
1*
b110 6
19
1>
1C
b110 G
#50700000000
0!
0*
09
0>
0C
#50710000000
1!
1*
b111 6
19
1>
1C
b111 G
#50720000000
0!
0*
09
0>
0C
#50730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#50740000000
0!
0*
09
0>
0C
#50750000000
1!
1*
b1 6
19
1>
1C
b1 G
#50760000000
0!
0*
09
0>
0C
#50770000000
1!
1*
b10 6
19
1>
1C
b10 G
#50780000000
0!
0*
09
0>
0C
#50790000000
1!
1*
b11 6
19
1>
1C
b11 G
#50800000000
0!
0*
09
0>
0C
#50810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#50820000000
0!
0*
09
0>
0C
#50830000000
1!
1*
b101 6
19
1>
1C
b101 G
#50840000000
0!
0*
09
0>
0C
#50850000000
1!
1*
b110 6
19
1>
1C
b110 G
#50860000000
0!
0*
09
0>
0C
#50870000000
1!
1*
b111 6
19
1>
1C
b111 G
#50880000000
0!
0*
09
0>
0C
#50890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#50900000000
0!
0*
09
0>
0C
#50910000000
1!
1*
b1 6
19
1>
1C
b1 G
#50920000000
0!
0*
09
0>
0C
#50930000000
1!
1*
b10 6
19
1>
1C
b10 G
#50940000000
0!
0*
09
0>
0C
#50950000000
1!
1*
b11 6
19
1>
1C
b11 G
#50960000000
0!
0*
09
0>
0C
#50970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#50980000000
0!
0*
09
0>
0C
#50990000000
1!
1*
b101 6
19
1>
1C
b101 G
#51000000000
0!
0*
09
0>
0C
#51010000000
1!
1*
b110 6
19
1>
1C
b110 G
#51020000000
0!
0*
09
0>
0C
#51030000000
1!
1*
b111 6
19
1>
1C
b111 G
#51040000000
0!
1"
0*
1+
09
1:
0>
0C
#51050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#51060000000
0!
0*
09
0>
0C
#51070000000
1!
1*
b1 6
19
1>
1C
b1 G
#51080000000
0!
0*
09
0>
0C
#51090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#51100000000
0!
0*
09
0>
0C
#51110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#51120000000
0!
0*
09
0>
0C
#51130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#51140000000
0!
0*
09
0>
0C
#51150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#51160000000
0!
0#
0*
0,
09
0>
0?
0C
#51170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#51180000000
0!
0*
09
0>
0C
#51190000000
1!
1*
19
1>
1C
#51200000000
0!
0*
09
0>
0C
#51210000000
1!
1*
19
1>
1C
#51220000000
0!
0*
09
0>
0C
#51230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#51240000000
0!
0*
09
0>
0C
#51250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#51260000000
0!
0*
09
0>
0C
#51270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#51280000000
0!
0*
09
0>
0C
#51290000000
1!
1*
b10 6
19
1>
1C
b10 G
#51300000000
0!
0*
09
0>
0C
#51310000000
1!
1*
b11 6
19
1>
1C
b11 G
#51320000000
0!
0*
09
0>
0C
#51330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#51340000000
0!
0*
09
0>
0C
#51350000000
1!
1*
b101 6
19
1>
1C
b101 G
#51360000000
0!
0*
09
0>
0C
#51370000000
1!
1*
b110 6
19
1>
1C
b110 G
#51380000000
0!
0*
09
0>
0C
#51390000000
1!
1*
b111 6
19
1>
1C
b111 G
#51400000000
0!
0*
09
0>
0C
#51410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#51420000000
0!
0*
09
0>
0C
#51430000000
1!
1*
b1 6
19
1>
1C
b1 G
#51440000000
0!
0*
09
0>
0C
#51450000000
1!
1*
b10 6
19
1>
1C
b10 G
#51460000000
0!
0*
09
0>
0C
#51470000000
1!
1*
b11 6
19
1>
1C
b11 G
#51480000000
0!
0*
09
0>
0C
#51490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#51500000000
0!
0*
09
0>
0C
#51510000000
1!
1*
b101 6
19
1>
1C
b101 G
#51520000000
0!
0*
09
0>
0C
#51530000000
1!
1*
b110 6
19
1>
1C
b110 G
#51540000000
0!
0*
09
0>
0C
#51550000000
1!
1*
b111 6
19
1>
1C
b111 G
#51560000000
0!
0*
09
0>
0C
#51570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#51580000000
0!
0*
09
0>
0C
#51590000000
1!
1*
b1 6
19
1>
1C
b1 G
#51600000000
0!
0*
09
0>
0C
#51610000000
1!
1*
b10 6
19
1>
1C
b10 G
#51620000000
0!
0*
09
0>
0C
#51630000000
1!
1*
b11 6
19
1>
1C
b11 G
#51640000000
0!
0*
09
0>
0C
#51650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#51660000000
0!
0*
09
0>
0C
#51670000000
1!
1*
b101 6
19
1>
1C
b101 G
#51680000000
0!
0*
09
0>
0C
#51690000000
1!
1*
b110 6
19
1>
1C
b110 G
#51700000000
0!
0*
09
0>
0C
#51710000000
1!
1*
b111 6
19
1>
1C
b111 G
#51720000000
0!
1"
0*
1+
09
1:
0>
0C
#51730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#51740000000
0!
0*
09
0>
0C
#51750000000
1!
1*
b1 6
19
1>
1C
b1 G
#51760000000
0!
0*
09
0>
0C
#51770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#51780000000
0!
0*
09
0>
0C
#51790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#51800000000
0!
0*
09
0>
0C
#51810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#51820000000
0!
0*
09
0>
0C
#51830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#51840000000
0!
0#
0*
0,
09
0>
0?
0C
#51850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#51860000000
0!
0*
09
0>
0C
#51870000000
1!
1*
19
1>
1C
#51880000000
0!
0*
09
0>
0C
#51890000000
1!
1*
19
1>
1C
#51900000000
0!
0*
09
0>
0C
#51910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#51920000000
0!
0*
09
0>
0C
#51930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#51940000000
0!
0*
09
0>
0C
#51950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#51960000000
0!
0*
09
0>
0C
#51970000000
1!
1*
b10 6
19
1>
1C
b10 G
#51980000000
0!
0*
09
0>
0C
#51990000000
1!
1*
b11 6
19
1>
1C
b11 G
#52000000000
0!
0*
09
0>
0C
#52010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#52020000000
0!
0*
09
0>
0C
#52030000000
1!
1*
b101 6
19
1>
1C
b101 G
#52040000000
0!
0*
09
0>
0C
#52050000000
1!
1*
b110 6
19
1>
1C
b110 G
#52060000000
0!
0*
09
0>
0C
#52070000000
1!
1*
b111 6
19
1>
1C
b111 G
#52080000000
0!
0*
09
0>
0C
#52090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#52100000000
0!
0*
09
0>
0C
#52110000000
1!
1*
b1 6
19
1>
1C
b1 G
#52120000000
0!
0*
09
0>
0C
#52130000000
1!
1*
b10 6
19
1>
1C
b10 G
#52140000000
0!
0*
09
0>
0C
#52150000000
1!
1*
b11 6
19
1>
1C
b11 G
#52160000000
0!
0*
09
0>
0C
#52170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#52180000000
0!
0*
09
0>
0C
#52190000000
1!
1*
b101 6
19
1>
1C
b101 G
#52200000000
0!
0*
09
0>
0C
#52210000000
1!
1*
b110 6
19
1>
1C
b110 G
#52220000000
0!
0*
09
0>
0C
#52230000000
1!
1*
b111 6
19
1>
1C
b111 G
#52240000000
0!
0*
09
0>
0C
#52250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#52260000000
0!
0*
09
0>
0C
#52270000000
1!
1*
b1 6
19
1>
1C
b1 G
#52280000000
0!
0*
09
0>
0C
#52290000000
1!
1*
b10 6
19
1>
1C
b10 G
#52300000000
0!
0*
09
0>
0C
#52310000000
1!
1*
b11 6
19
1>
1C
b11 G
#52320000000
0!
0*
09
0>
0C
#52330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#52340000000
0!
0*
09
0>
0C
#52350000000
1!
1*
b101 6
19
1>
1C
b101 G
#52360000000
0!
0*
09
0>
0C
#52370000000
1!
1*
b110 6
19
1>
1C
b110 G
#52380000000
0!
0*
09
0>
0C
#52390000000
1!
1*
b111 6
19
1>
1C
b111 G
#52400000000
0!
1"
0*
1+
09
1:
0>
0C
#52410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#52420000000
0!
0*
09
0>
0C
#52430000000
1!
1*
b1 6
19
1>
1C
b1 G
#52440000000
0!
0*
09
0>
0C
#52450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#52460000000
0!
0*
09
0>
0C
#52470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#52480000000
0!
0*
09
0>
0C
#52490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#52500000000
0!
0*
09
0>
0C
#52510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#52520000000
0!
0#
0*
0,
09
0>
0?
0C
#52530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#52540000000
0!
0*
09
0>
0C
#52550000000
1!
1*
19
1>
1C
#52560000000
0!
0*
09
0>
0C
#52570000000
1!
1*
19
1>
1C
#52580000000
0!
0*
09
0>
0C
#52590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#52600000000
0!
0*
09
0>
0C
#52610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#52620000000
0!
0*
09
0>
0C
#52630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#52640000000
0!
0*
09
0>
0C
#52650000000
1!
1*
b10 6
19
1>
1C
b10 G
#52660000000
0!
0*
09
0>
0C
#52670000000
1!
1*
b11 6
19
1>
1C
b11 G
#52680000000
0!
0*
09
0>
0C
#52690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#52700000000
0!
0*
09
0>
0C
#52710000000
1!
1*
b101 6
19
1>
1C
b101 G
#52720000000
0!
0*
09
0>
0C
#52730000000
1!
1*
b110 6
19
1>
1C
b110 G
#52740000000
0!
0*
09
0>
0C
#52750000000
1!
1*
b111 6
19
1>
1C
b111 G
#52760000000
0!
0*
09
0>
0C
#52770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#52780000000
0!
0*
09
0>
0C
#52790000000
1!
1*
b1 6
19
1>
1C
b1 G
#52800000000
0!
0*
09
0>
0C
#52810000000
1!
1*
b10 6
19
1>
1C
b10 G
#52820000000
0!
0*
09
0>
0C
#52830000000
1!
1*
b11 6
19
1>
1C
b11 G
#52840000000
0!
0*
09
0>
0C
#52850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#52860000000
0!
0*
09
0>
0C
#52870000000
1!
1*
b101 6
19
1>
1C
b101 G
#52880000000
0!
0*
09
0>
0C
#52890000000
1!
1*
b110 6
19
1>
1C
b110 G
#52900000000
0!
0*
09
0>
0C
#52910000000
1!
1*
b111 6
19
1>
1C
b111 G
#52920000000
0!
0*
09
0>
0C
#52930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#52940000000
0!
0*
09
0>
0C
#52950000000
1!
1*
b1 6
19
1>
1C
b1 G
#52960000000
0!
0*
09
0>
0C
#52970000000
1!
1*
b10 6
19
1>
1C
b10 G
#52980000000
0!
0*
09
0>
0C
#52990000000
1!
1*
b11 6
19
1>
1C
b11 G
#53000000000
0!
0*
09
0>
0C
#53010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#53020000000
0!
0*
09
0>
0C
#53030000000
1!
1*
b101 6
19
1>
1C
b101 G
#53040000000
0!
0*
09
0>
0C
#53050000000
1!
1*
b110 6
19
1>
1C
b110 G
#53060000000
0!
0*
09
0>
0C
#53070000000
1!
1*
b111 6
19
1>
1C
b111 G
#53080000000
0!
1"
0*
1+
09
1:
0>
0C
#53090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#53100000000
0!
0*
09
0>
0C
#53110000000
1!
1*
b1 6
19
1>
1C
b1 G
#53120000000
0!
0*
09
0>
0C
#53130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#53140000000
0!
0*
09
0>
0C
#53150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#53160000000
0!
0*
09
0>
0C
#53170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#53180000000
0!
0*
09
0>
0C
#53190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#53200000000
0!
0#
0*
0,
09
0>
0?
0C
#53210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#53220000000
0!
0*
09
0>
0C
#53230000000
1!
1*
19
1>
1C
#53240000000
0!
0*
09
0>
0C
#53250000000
1!
1*
19
1>
1C
#53260000000
0!
0*
09
0>
0C
#53270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#53280000000
0!
0*
09
0>
0C
#53290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#53300000000
0!
0*
09
0>
0C
#53310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#53320000000
0!
0*
09
0>
0C
#53330000000
1!
1*
b10 6
19
1>
1C
b10 G
#53340000000
0!
0*
09
0>
0C
#53350000000
1!
1*
b11 6
19
1>
1C
b11 G
#53360000000
0!
0*
09
0>
0C
#53370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#53380000000
0!
0*
09
0>
0C
#53390000000
1!
1*
b101 6
19
1>
1C
b101 G
#53400000000
0!
0*
09
0>
0C
#53410000000
1!
1*
b110 6
19
1>
1C
b110 G
#53420000000
0!
0*
09
0>
0C
#53430000000
1!
1*
b111 6
19
1>
1C
b111 G
#53440000000
0!
0*
09
0>
0C
#53450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#53460000000
0!
0*
09
0>
0C
#53470000000
1!
1*
b1 6
19
1>
1C
b1 G
#53480000000
0!
0*
09
0>
0C
#53490000000
1!
1*
b10 6
19
1>
1C
b10 G
#53500000000
0!
0*
09
0>
0C
#53510000000
1!
1*
b11 6
19
1>
1C
b11 G
#53520000000
0!
0*
09
0>
0C
#53530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#53540000000
0!
0*
09
0>
0C
#53550000000
1!
1*
b101 6
19
1>
1C
b101 G
#53560000000
0!
0*
09
0>
0C
#53570000000
1!
1*
b110 6
19
1>
1C
b110 G
#53580000000
0!
0*
09
0>
0C
#53590000000
1!
1*
b111 6
19
1>
1C
b111 G
#53600000000
0!
0*
09
0>
0C
#53610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#53620000000
0!
0*
09
0>
0C
#53630000000
1!
1*
b1 6
19
1>
1C
b1 G
#53640000000
0!
0*
09
0>
0C
#53650000000
1!
1*
b10 6
19
1>
1C
b10 G
#53660000000
0!
0*
09
0>
0C
#53670000000
1!
1*
b11 6
19
1>
1C
b11 G
#53680000000
0!
0*
09
0>
0C
#53690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#53700000000
0!
0*
09
0>
0C
#53710000000
1!
1*
b101 6
19
1>
1C
b101 G
#53720000000
0!
0*
09
0>
0C
#53730000000
1!
1*
b110 6
19
1>
1C
b110 G
#53740000000
0!
0*
09
0>
0C
#53750000000
1!
1*
b111 6
19
1>
1C
b111 G
#53760000000
0!
1"
0*
1+
09
1:
0>
0C
#53770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#53780000000
0!
0*
09
0>
0C
#53790000000
1!
1*
b1 6
19
1>
1C
b1 G
#53800000000
0!
0*
09
0>
0C
#53810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#53820000000
0!
0*
09
0>
0C
#53830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#53840000000
0!
0*
09
0>
0C
#53850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#53860000000
0!
0*
09
0>
0C
#53870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#53880000000
0!
0#
0*
0,
09
0>
0?
0C
#53890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#53900000000
0!
0*
09
0>
0C
#53910000000
1!
1*
19
1>
1C
#53920000000
0!
0*
09
0>
0C
#53930000000
1!
1*
19
1>
1C
#53940000000
0!
0*
09
0>
0C
#53950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#53960000000
0!
0*
09
0>
0C
#53970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#53980000000
0!
0*
09
0>
0C
#53990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#54000000000
0!
0*
09
0>
0C
#54010000000
1!
1*
b10 6
19
1>
1C
b10 G
#54020000000
0!
0*
09
0>
0C
#54030000000
1!
1*
b11 6
19
1>
1C
b11 G
#54040000000
0!
0*
09
0>
0C
#54050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#54060000000
0!
0*
09
0>
0C
#54070000000
1!
1*
b101 6
19
1>
1C
b101 G
#54080000000
0!
0*
09
0>
0C
#54090000000
1!
1*
b110 6
19
1>
1C
b110 G
#54100000000
0!
0*
09
0>
0C
#54110000000
1!
1*
b111 6
19
1>
1C
b111 G
#54120000000
0!
0*
09
0>
0C
#54130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#54140000000
0!
0*
09
0>
0C
#54150000000
1!
1*
b1 6
19
1>
1C
b1 G
#54160000000
0!
0*
09
0>
0C
#54170000000
1!
1*
b10 6
19
1>
1C
b10 G
#54180000000
0!
0*
09
0>
0C
#54190000000
1!
1*
b11 6
19
1>
1C
b11 G
#54200000000
0!
0*
09
0>
0C
#54210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#54220000000
0!
0*
09
0>
0C
#54230000000
1!
1*
b101 6
19
1>
1C
b101 G
#54240000000
0!
0*
09
0>
0C
#54250000000
1!
1*
b110 6
19
1>
1C
b110 G
#54260000000
0!
0*
09
0>
0C
#54270000000
1!
1*
b111 6
19
1>
1C
b111 G
#54280000000
0!
0*
09
0>
0C
#54290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#54300000000
0!
0*
09
0>
0C
#54310000000
1!
1*
b1 6
19
1>
1C
b1 G
#54320000000
0!
0*
09
0>
0C
#54330000000
1!
1*
b10 6
19
1>
1C
b10 G
#54340000000
0!
0*
09
0>
0C
#54350000000
1!
1*
b11 6
19
1>
1C
b11 G
#54360000000
0!
0*
09
0>
0C
#54370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#54380000000
0!
0*
09
0>
0C
#54390000000
1!
1*
b101 6
19
1>
1C
b101 G
#54400000000
0!
0*
09
0>
0C
#54410000000
1!
1*
b110 6
19
1>
1C
b110 G
#54420000000
0!
0*
09
0>
0C
#54430000000
1!
1*
b111 6
19
1>
1C
b111 G
#54440000000
0!
1"
0*
1+
09
1:
0>
0C
#54450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#54460000000
0!
0*
09
0>
0C
#54470000000
1!
1*
b1 6
19
1>
1C
b1 G
#54480000000
0!
0*
09
0>
0C
#54490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#54500000000
0!
0*
09
0>
0C
#54510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#54520000000
0!
0*
09
0>
0C
#54530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#54540000000
0!
0*
09
0>
0C
#54550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#54560000000
0!
0#
0*
0,
09
0>
0?
0C
#54570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#54580000000
0!
0*
09
0>
0C
#54590000000
1!
1*
19
1>
1C
#54600000000
0!
0*
09
0>
0C
#54610000000
1!
1*
19
1>
1C
#54620000000
0!
0*
09
0>
0C
#54630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#54640000000
0!
0*
09
0>
0C
#54650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#54660000000
0!
0*
09
0>
0C
#54670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#54680000000
0!
0*
09
0>
0C
#54690000000
1!
1*
b10 6
19
1>
1C
b10 G
#54700000000
0!
0*
09
0>
0C
#54710000000
1!
1*
b11 6
19
1>
1C
b11 G
#54720000000
0!
0*
09
0>
0C
#54730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#54740000000
0!
0*
09
0>
0C
#54750000000
1!
1*
b101 6
19
1>
1C
b101 G
#54760000000
0!
0*
09
0>
0C
#54770000000
1!
1*
b110 6
19
1>
1C
b110 G
#54780000000
0!
0*
09
0>
0C
#54790000000
1!
1*
b111 6
19
1>
1C
b111 G
#54800000000
0!
0*
09
0>
0C
#54810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#54820000000
0!
0*
09
0>
0C
#54830000000
1!
1*
b1 6
19
1>
1C
b1 G
#54840000000
0!
0*
09
0>
0C
#54850000000
1!
1*
b10 6
19
1>
1C
b10 G
#54860000000
0!
0*
09
0>
0C
#54870000000
1!
1*
b11 6
19
1>
1C
b11 G
#54880000000
0!
0*
09
0>
0C
#54890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#54900000000
0!
0*
09
0>
0C
#54910000000
1!
1*
b101 6
19
1>
1C
b101 G
#54920000000
0!
0*
09
0>
0C
#54930000000
1!
1*
b110 6
19
1>
1C
b110 G
#54940000000
0!
0*
09
0>
0C
#54950000000
1!
1*
b111 6
19
1>
1C
b111 G
#54960000000
0!
0*
09
0>
0C
#54970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#54980000000
0!
0*
09
0>
0C
#54990000000
1!
1*
b1 6
19
1>
1C
b1 G
#55000000000
0!
0*
09
0>
0C
#55010000000
1!
1*
b10 6
19
1>
1C
b10 G
#55020000000
0!
0*
09
0>
0C
#55030000000
1!
1*
b11 6
19
1>
1C
b11 G
#55040000000
0!
0*
09
0>
0C
#55050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#55060000000
0!
0*
09
0>
0C
#55070000000
1!
1*
b101 6
19
1>
1C
b101 G
#55080000000
0!
0*
09
0>
0C
#55090000000
1!
1*
b110 6
19
1>
1C
b110 G
#55100000000
0!
0*
09
0>
0C
#55110000000
1!
1*
b111 6
19
1>
1C
b111 G
#55120000000
0!
1"
0*
1+
09
1:
0>
0C
#55130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#55140000000
0!
0*
09
0>
0C
#55150000000
1!
1*
b1 6
19
1>
1C
b1 G
#55160000000
0!
0*
09
0>
0C
#55170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#55180000000
0!
0*
09
0>
0C
#55190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#55200000000
0!
0*
09
0>
0C
#55210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#55220000000
0!
0*
09
0>
0C
#55230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#55240000000
0!
0#
0*
0,
09
0>
0?
0C
#55250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#55260000000
0!
0*
09
0>
0C
#55270000000
1!
1*
19
1>
1C
#55280000000
0!
0*
09
0>
0C
#55290000000
1!
1*
19
1>
1C
#55300000000
0!
0*
09
0>
0C
#55310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#55320000000
0!
0*
09
0>
0C
#55330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#55340000000
0!
0*
09
0>
0C
#55350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#55360000000
0!
0*
09
0>
0C
#55370000000
1!
1*
b10 6
19
1>
1C
b10 G
#55380000000
0!
0*
09
0>
0C
#55390000000
1!
1*
b11 6
19
1>
1C
b11 G
#55400000000
0!
0*
09
0>
0C
#55410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#55420000000
0!
0*
09
0>
0C
#55430000000
1!
1*
b101 6
19
1>
1C
b101 G
#55440000000
0!
0*
09
0>
0C
#55450000000
1!
1*
b110 6
19
1>
1C
b110 G
#55460000000
0!
0*
09
0>
0C
#55470000000
1!
1*
b111 6
19
1>
1C
b111 G
#55480000000
0!
0*
09
0>
0C
#55490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#55500000000
0!
0*
09
0>
0C
#55510000000
1!
1*
b1 6
19
1>
1C
b1 G
#55520000000
0!
0*
09
0>
0C
#55530000000
1!
1*
b10 6
19
1>
1C
b10 G
#55540000000
0!
0*
09
0>
0C
#55550000000
1!
1*
b11 6
19
1>
1C
b11 G
#55560000000
0!
0*
09
0>
0C
#55570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#55580000000
0!
0*
09
0>
0C
#55590000000
1!
1*
b101 6
19
1>
1C
b101 G
#55600000000
0!
0*
09
0>
0C
#55610000000
1!
1*
b110 6
19
1>
1C
b110 G
#55620000000
0!
0*
09
0>
0C
#55630000000
1!
1*
b111 6
19
1>
1C
b111 G
#55640000000
0!
0*
09
0>
0C
#55650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#55660000000
0!
0*
09
0>
0C
#55670000000
1!
1*
b1 6
19
1>
1C
b1 G
#55680000000
0!
0*
09
0>
0C
#55690000000
1!
1*
b10 6
19
1>
1C
b10 G
#55700000000
0!
0*
09
0>
0C
#55710000000
1!
1*
b11 6
19
1>
1C
b11 G
#55720000000
0!
0*
09
0>
0C
#55730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#55740000000
0!
0*
09
0>
0C
#55750000000
1!
1*
b101 6
19
1>
1C
b101 G
#55760000000
0!
0*
09
0>
0C
#55770000000
1!
1*
b110 6
19
1>
1C
b110 G
#55780000000
0!
0*
09
0>
0C
#55790000000
1!
1*
b111 6
19
1>
1C
b111 G
#55800000000
0!
1"
0*
1+
09
1:
0>
0C
#55810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#55820000000
0!
0*
09
0>
0C
#55830000000
1!
1*
b1 6
19
1>
1C
b1 G
#55840000000
0!
0*
09
0>
0C
#55850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#55860000000
0!
0*
09
0>
0C
#55870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#55880000000
0!
0*
09
0>
0C
#55890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#55900000000
0!
0*
09
0>
0C
#55910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#55920000000
0!
0#
0*
0,
09
0>
0?
0C
#55930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#55940000000
0!
0*
09
0>
0C
#55950000000
1!
1*
19
1>
1C
#55960000000
0!
0*
09
0>
0C
#55970000000
1!
1*
19
1>
1C
#55980000000
0!
0*
09
0>
0C
#55990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#56000000000
0!
0*
09
0>
0C
#56010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#56020000000
0!
0*
09
0>
0C
#56030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#56040000000
0!
0*
09
0>
0C
#56050000000
1!
1*
b10 6
19
1>
1C
b10 G
#56060000000
0!
0*
09
0>
0C
#56070000000
1!
1*
b11 6
19
1>
1C
b11 G
#56080000000
0!
0*
09
0>
0C
#56090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#56100000000
0!
0*
09
0>
0C
#56110000000
1!
1*
b101 6
19
1>
1C
b101 G
#56120000000
0!
0*
09
0>
0C
#56130000000
1!
1*
b110 6
19
1>
1C
b110 G
#56140000000
0!
0*
09
0>
0C
#56150000000
1!
1*
b111 6
19
1>
1C
b111 G
#56160000000
0!
0*
09
0>
0C
#56170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#56180000000
0!
0*
09
0>
0C
#56190000000
1!
1*
b1 6
19
1>
1C
b1 G
#56200000000
0!
0*
09
0>
0C
#56210000000
1!
1*
b10 6
19
1>
1C
b10 G
#56220000000
0!
0*
09
0>
0C
#56230000000
1!
1*
b11 6
19
1>
1C
b11 G
#56240000000
0!
0*
09
0>
0C
#56250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#56260000000
0!
0*
09
0>
0C
#56270000000
1!
1*
b101 6
19
1>
1C
b101 G
#56280000000
0!
0*
09
0>
0C
#56290000000
1!
1*
b110 6
19
1>
1C
b110 G
#56300000000
0!
0*
09
0>
0C
#56310000000
1!
1*
b111 6
19
1>
1C
b111 G
#56320000000
0!
0*
09
0>
0C
#56330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#56340000000
0!
0*
09
0>
0C
#56350000000
1!
1*
b1 6
19
1>
1C
b1 G
#56360000000
0!
0*
09
0>
0C
#56370000000
1!
1*
b10 6
19
1>
1C
b10 G
#56380000000
0!
0*
09
0>
0C
#56390000000
1!
1*
b11 6
19
1>
1C
b11 G
#56400000000
0!
0*
09
0>
0C
#56410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#56420000000
0!
0*
09
0>
0C
#56430000000
1!
1*
b101 6
19
1>
1C
b101 G
#56440000000
0!
0*
09
0>
0C
#56450000000
1!
1*
b110 6
19
1>
1C
b110 G
#56460000000
0!
0*
09
0>
0C
#56470000000
1!
1*
b111 6
19
1>
1C
b111 G
#56480000000
0!
1"
0*
1+
09
1:
0>
0C
#56490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#56500000000
0!
0*
09
0>
0C
#56510000000
1!
1*
b1 6
19
1>
1C
b1 G
#56520000000
0!
0*
09
0>
0C
#56530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#56540000000
0!
0*
09
0>
0C
#56550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#56560000000
0!
0*
09
0>
0C
#56570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#56580000000
0!
0*
09
0>
0C
#56590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#56600000000
0!
0#
0*
0,
09
0>
0?
0C
#56610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#56620000000
0!
0*
09
0>
0C
#56630000000
1!
1*
19
1>
1C
#56640000000
0!
0*
09
0>
0C
#56650000000
1!
1*
19
1>
1C
#56660000000
0!
0*
09
0>
0C
#56670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#56680000000
0!
0*
09
0>
0C
#56690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#56700000000
0!
0*
09
0>
0C
#56710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#56720000000
0!
0*
09
0>
0C
#56730000000
1!
1*
b10 6
19
1>
1C
b10 G
#56740000000
0!
0*
09
0>
0C
#56750000000
1!
1*
b11 6
19
1>
1C
b11 G
#56760000000
0!
0*
09
0>
0C
#56770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#56780000000
0!
0*
09
0>
0C
#56790000000
1!
1*
b101 6
19
1>
1C
b101 G
#56800000000
0!
0*
09
0>
0C
#56810000000
1!
1*
b110 6
19
1>
1C
b110 G
#56820000000
0!
0*
09
0>
0C
#56830000000
1!
1*
b111 6
19
1>
1C
b111 G
#56840000000
0!
0*
09
0>
0C
#56850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#56860000000
0!
0*
09
0>
0C
#56870000000
1!
1*
b1 6
19
1>
1C
b1 G
#56880000000
0!
0*
09
0>
0C
#56890000000
1!
1*
b10 6
19
1>
1C
b10 G
#56900000000
0!
0*
09
0>
0C
#56910000000
1!
1*
b11 6
19
1>
1C
b11 G
#56920000000
0!
0*
09
0>
0C
#56930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#56940000000
0!
0*
09
0>
0C
#56950000000
1!
1*
b101 6
19
1>
1C
b101 G
#56960000000
0!
0*
09
0>
0C
#56970000000
1!
1*
b110 6
19
1>
1C
b110 G
#56980000000
0!
0*
09
0>
0C
#56990000000
1!
1*
b111 6
19
1>
1C
b111 G
#57000000000
0!
0*
09
0>
0C
#57010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#57020000000
0!
0*
09
0>
0C
#57030000000
1!
1*
b1 6
19
1>
1C
b1 G
#57040000000
0!
0*
09
0>
0C
#57050000000
1!
1*
b10 6
19
1>
1C
b10 G
#57060000000
0!
0*
09
0>
0C
#57070000000
1!
1*
b11 6
19
1>
1C
b11 G
#57080000000
0!
0*
09
0>
0C
#57090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#57100000000
0!
0*
09
0>
0C
#57110000000
1!
1*
b101 6
19
1>
1C
b101 G
#57120000000
0!
0*
09
0>
0C
#57130000000
1!
1*
b110 6
19
1>
1C
b110 G
#57140000000
0!
0*
09
0>
0C
#57150000000
1!
1*
b111 6
19
1>
1C
b111 G
#57160000000
0!
1"
0*
1+
09
1:
0>
0C
#57170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#57180000000
0!
0*
09
0>
0C
#57190000000
1!
1*
b1 6
19
1>
1C
b1 G
#57200000000
0!
0*
09
0>
0C
#57210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#57220000000
0!
0*
09
0>
0C
#57230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#57240000000
0!
0*
09
0>
0C
#57250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#57260000000
0!
0*
09
0>
0C
#57270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#57280000000
0!
0#
0*
0,
09
0>
0?
0C
#57290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#57300000000
0!
0*
09
0>
0C
#57310000000
1!
1*
19
1>
1C
#57320000000
0!
0*
09
0>
0C
#57330000000
1!
1*
19
1>
1C
#57340000000
0!
0*
09
0>
0C
#57350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#57360000000
0!
0*
09
0>
0C
#57370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#57380000000
0!
0*
09
0>
0C
#57390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#57400000000
0!
0*
09
0>
0C
#57410000000
1!
1*
b10 6
19
1>
1C
b10 G
#57420000000
0!
0*
09
0>
0C
#57430000000
1!
1*
b11 6
19
1>
1C
b11 G
#57440000000
0!
0*
09
0>
0C
#57450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#57460000000
0!
0*
09
0>
0C
#57470000000
1!
1*
b101 6
19
1>
1C
b101 G
#57480000000
0!
0*
09
0>
0C
#57490000000
1!
1*
b110 6
19
1>
1C
b110 G
#57500000000
0!
0*
09
0>
0C
#57510000000
1!
1*
b111 6
19
1>
1C
b111 G
#57520000000
0!
0*
09
0>
0C
#57530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#57540000000
0!
0*
09
0>
0C
#57550000000
1!
1*
b1 6
19
1>
1C
b1 G
#57560000000
0!
0*
09
0>
0C
#57570000000
1!
1*
b10 6
19
1>
1C
b10 G
#57580000000
0!
0*
09
0>
0C
#57590000000
1!
1*
b11 6
19
1>
1C
b11 G
#57600000000
0!
0*
09
0>
0C
#57610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#57620000000
0!
0*
09
0>
0C
#57630000000
1!
1*
b101 6
19
1>
1C
b101 G
#57640000000
0!
0*
09
0>
0C
#57650000000
1!
1*
b110 6
19
1>
1C
b110 G
#57660000000
0!
0*
09
0>
0C
#57670000000
1!
1*
b111 6
19
1>
1C
b111 G
#57680000000
0!
0*
09
0>
0C
#57690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#57700000000
0!
0*
09
0>
0C
#57710000000
1!
1*
b1 6
19
1>
1C
b1 G
#57720000000
0!
0*
09
0>
0C
#57730000000
1!
1*
b10 6
19
1>
1C
b10 G
#57740000000
0!
0*
09
0>
0C
#57750000000
1!
1*
b11 6
19
1>
1C
b11 G
#57760000000
0!
0*
09
0>
0C
#57770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#57780000000
0!
0*
09
0>
0C
#57790000000
1!
1*
b101 6
19
1>
1C
b101 G
#57800000000
0!
0*
09
0>
0C
#57810000000
1!
1*
b110 6
19
1>
1C
b110 G
#57820000000
0!
0*
09
0>
0C
#57830000000
1!
1*
b111 6
19
1>
1C
b111 G
#57840000000
0!
1"
0*
1+
09
1:
0>
0C
#57850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#57860000000
0!
0*
09
0>
0C
#57870000000
1!
1*
b1 6
19
1>
1C
b1 G
#57880000000
0!
0*
09
0>
0C
#57890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#57900000000
0!
0*
09
0>
0C
#57910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#57920000000
0!
0*
09
0>
0C
#57930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#57940000000
0!
0*
09
0>
0C
#57950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#57960000000
0!
0#
0*
0,
09
0>
0?
0C
#57970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#57980000000
0!
0*
09
0>
0C
#57990000000
1!
1*
19
1>
1C
#58000000000
0!
0*
09
0>
0C
#58010000000
1!
1*
19
1>
1C
#58020000000
0!
0*
09
0>
0C
#58030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#58040000000
0!
0*
09
0>
0C
#58050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#58060000000
0!
0*
09
0>
0C
#58070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#58080000000
0!
0*
09
0>
0C
#58090000000
1!
1*
b10 6
19
1>
1C
b10 G
#58100000000
0!
0*
09
0>
0C
#58110000000
1!
1*
b11 6
19
1>
1C
b11 G
#58120000000
0!
0*
09
0>
0C
#58130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#58140000000
0!
0*
09
0>
0C
#58150000000
1!
1*
b101 6
19
1>
1C
b101 G
#58160000000
0!
0*
09
0>
0C
#58170000000
1!
1*
b110 6
19
1>
1C
b110 G
#58180000000
0!
0*
09
0>
0C
#58190000000
1!
1*
b111 6
19
1>
1C
b111 G
#58200000000
0!
0*
09
0>
0C
#58210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#58220000000
0!
0*
09
0>
0C
#58230000000
1!
1*
b1 6
19
1>
1C
b1 G
#58240000000
0!
0*
09
0>
0C
#58250000000
1!
1*
b10 6
19
1>
1C
b10 G
#58260000000
0!
0*
09
0>
0C
#58270000000
1!
1*
b11 6
19
1>
1C
b11 G
#58280000000
0!
0*
09
0>
0C
#58290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#58300000000
0!
0*
09
0>
0C
#58310000000
1!
1*
b101 6
19
1>
1C
b101 G
#58320000000
0!
0*
09
0>
0C
#58330000000
1!
1*
b110 6
19
1>
1C
b110 G
#58340000000
0!
0*
09
0>
0C
#58350000000
1!
1*
b111 6
19
1>
1C
b111 G
#58360000000
0!
0*
09
0>
0C
#58370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#58380000000
0!
0*
09
0>
0C
#58390000000
1!
1*
b1 6
19
1>
1C
b1 G
#58400000000
0!
0*
09
0>
0C
#58410000000
1!
1*
b10 6
19
1>
1C
b10 G
#58420000000
0!
0*
09
0>
0C
#58430000000
1!
1*
b11 6
19
1>
1C
b11 G
#58440000000
0!
0*
09
0>
0C
#58450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#58460000000
0!
0*
09
0>
0C
#58470000000
1!
1*
b101 6
19
1>
1C
b101 G
#58480000000
0!
0*
09
0>
0C
#58490000000
1!
1*
b110 6
19
1>
1C
b110 G
#58500000000
0!
0*
09
0>
0C
#58510000000
1!
1*
b111 6
19
1>
1C
b111 G
#58520000000
0!
1"
0*
1+
09
1:
0>
0C
#58530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#58540000000
0!
0*
09
0>
0C
#58550000000
1!
1*
b1 6
19
1>
1C
b1 G
#58560000000
0!
0*
09
0>
0C
#58570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#58580000000
0!
0*
09
0>
0C
#58590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#58600000000
0!
0*
09
0>
0C
#58610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#58620000000
0!
0*
09
0>
0C
#58630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#58640000000
0!
0#
0*
0,
09
0>
0?
0C
#58650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#58660000000
0!
0*
09
0>
0C
#58670000000
1!
1*
19
1>
1C
#58680000000
0!
0*
09
0>
0C
#58690000000
1!
1*
19
1>
1C
#58700000000
0!
0*
09
0>
0C
#58710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#58720000000
0!
0*
09
0>
0C
#58730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#58740000000
0!
0*
09
0>
0C
#58750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#58760000000
0!
0*
09
0>
0C
#58770000000
1!
1*
b10 6
19
1>
1C
b10 G
#58780000000
0!
0*
09
0>
0C
#58790000000
1!
1*
b11 6
19
1>
1C
b11 G
#58800000000
0!
0*
09
0>
0C
#58810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#58820000000
0!
0*
09
0>
0C
#58830000000
1!
1*
b101 6
19
1>
1C
b101 G
#58840000000
0!
0*
09
0>
0C
#58850000000
1!
1*
b110 6
19
1>
1C
b110 G
#58860000000
0!
0*
09
0>
0C
#58870000000
1!
1*
b111 6
19
1>
1C
b111 G
#58880000000
0!
0*
09
0>
0C
#58890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#58900000000
0!
0*
09
0>
0C
#58910000000
1!
1*
b1 6
19
1>
1C
b1 G
#58920000000
0!
0*
09
0>
0C
#58930000000
1!
1*
b10 6
19
1>
1C
b10 G
#58940000000
0!
0*
09
0>
0C
#58950000000
1!
1*
b11 6
19
1>
1C
b11 G
#58960000000
0!
0*
09
0>
0C
#58970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#58980000000
0!
0*
09
0>
0C
#58990000000
1!
1*
b101 6
19
1>
1C
b101 G
#59000000000
0!
0*
09
0>
0C
#59010000000
1!
1*
b110 6
19
1>
1C
b110 G
#59020000000
0!
0*
09
0>
0C
#59030000000
1!
1*
b111 6
19
1>
1C
b111 G
#59040000000
0!
0*
09
0>
0C
#59050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#59060000000
0!
0*
09
0>
0C
#59070000000
1!
1*
b1 6
19
1>
1C
b1 G
#59080000000
0!
0*
09
0>
0C
#59090000000
1!
1*
b10 6
19
1>
1C
b10 G
#59100000000
0!
0*
09
0>
0C
#59110000000
1!
1*
b11 6
19
1>
1C
b11 G
#59120000000
0!
0*
09
0>
0C
#59130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#59140000000
0!
0*
09
0>
0C
#59150000000
1!
1*
b101 6
19
1>
1C
b101 G
#59160000000
0!
0*
09
0>
0C
#59170000000
1!
1*
b110 6
19
1>
1C
b110 G
#59180000000
0!
0*
09
0>
0C
#59190000000
1!
1*
b111 6
19
1>
1C
b111 G
#59200000000
0!
1"
0*
1+
09
1:
0>
0C
#59210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#59220000000
0!
0*
09
0>
0C
#59230000000
1!
1*
b1 6
19
1>
1C
b1 G
#59240000000
0!
0*
09
0>
0C
#59250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#59260000000
0!
0*
09
0>
0C
#59270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#59280000000
0!
0*
09
0>
0C
#59290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#59300000000
0!
0*
09
0>
0C
#59310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#59320000000
0!
0#
0*
0,
09
0>
0?
0C
#59330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#59340000000
0!
0*
09
0>
0C
#59350000000
1!
1*
19
1>
1C
#59360000000
0!
0*
09
0>
0C
#59370000000
1!
1*
19
1>
1C
#59380000000
0!
0*
09
0>
0C
#59390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#59400000000
0!
0*
09
0>
0C
#59410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#59420000000
0!
0*
09
0>
0C
#59430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#59440000000
0!
0*
09
0>
0C
#59450000000
1!
1*
b10 6
19
1>
1C
b10 G
#59460000000
0!
0*
09
0>
0C
#59470000000
1!
1*
b11 6
19
1>
1C
b11 G
#59480000000
0!
0*
09
0>
0C
#59490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#59500000000
0!
0*
09
0>
0C
#59510000000
1!
1*
b101 6
19
1>
1C
b101 G
#59520000000
0!
0*
09
0>
0C
#59530000000
1!
1*
b110 6
19
1>
1C
b110 G
#59540000000
0!
0*
09
0>
0C
#59550000000
1!
1*
b111 6
19
1>
1C
b111 G
#59560000000
0!
0*
09
0>
0C
#59570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#59580000000
0!
0*
09
0>
0C
#59590000000
1!
1*
b1 6
19
1>
1C
b1 G
#59600000000
0!
0*
09
0>
0C
#59610000000
1!
1*
b10 6
19
1>
1C
b10 G
#59620000000
0!
0*
09
0>
0C
#59630000000
1!
1*
b11 6
19
1>
1C
b11 G
#59640000000
0!
0*
09
0>
0C
#59650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#59660000000
0!
0*
09
0>
0C
#59670000000
1!
1*
b101 6
19
1>
1C
b101 G
#59680000000
0!
0*
09
0>
0C
#59690000000
1!
1*
b110 6
19
1>
1C
b110 G
#59700000000
0!
0*
09
0>
0C
#59710000000
1!
1*
b111 6
19
1>
1C
b111 G
#59720000000
0!
0*
09
0>
0C
#59730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#59740000000
0!
0*
09
0>
0C
#59750000000
1!
1*
b1 6
19
1>
1C
b1 G
#59760000000
0!
0*
09
0>
0C
#59770000000
1!
1*
b10 6
19
1>
1C
b10 G
#59780000000
0!
0*
09
0>
0C
#59790000000
1!
1*
b11 6
19
1>
1C
b11 G
#59800000000
0!
0*
09
0>
0C
#59810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#59820000000
0!
0*
09
0>
0C
#59830000000
1!
1*
b101 6
19
1>
1C
b101 G
#59840000000
0!
0*
09
0>
0C
#59850000000
1!
1*
b110 6
19
1>
1C
b110 G
#59860000000
0!
0*
09
0>
0C
#59870000000
1!
1*
b111 6
19
1>
1C
b111 G
#59880000000
0!
1"
0*
1+
09
1:
0>
0C
#59890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#59900000000
0!
0*
09
0>
0C
#59910000000
1!
1*
b1 6
19
1>
1C
b1 G
#59920000000
0!
0*
09
0>
0C
#59930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#59940000000
0!
0*
09
0>
0C
#59950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#59960000000
0!
0*
09
0>
0C
#59970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#59980000000
0!
0*
09
0>
0C
#59990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#60000000000
0!
0#
0*
0,
09
0>
0?
0C
#60010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#60020000000
0!
0*
09
0>
0C
#60030000000
1!
1*
19
1>
1C
#60040000000
0!
0*
09
0>
0C
#60050000000
1!
1*
19
1>
1C
#60060000000
0!
0*
09
0>
0C
#60070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#60080000000
0!
0*
09
0>
0C
#60090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#60100000000
0!
0*
09
0>
0C
#60110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#60120000000
0!
0*
09
0>
0C
#60130000000
1!
1*
b10 6
19
1>
1C
b10 G
#60140000000
0!
0*
09
0>
0C
#60150000000
1!
1*
b11 6
19
1>
1C
b11 G
#60160000000
0!
0*
09
0>
0C
#60170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#60180000000
0!
0*
09
0>
0C
#60190000000
1!
1*
b101 6
19
1>
1C
b101 G
#60200000000
0!
0*
09
0>
0C
#60210000000
1!
1*
b110 6
19
1>
1C
b110 G
#60220000000
0!
0*
09
0>
0C
#60230000000
1!
1*
b111 6
19
1>
1C
b111 G
#60240000000
0!
0*
09
0>
0C
#60250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#60260000000
0!
0*
09
0>
0C
#60270000000
1!
1*
b1 6
19
1>
1C
b1 G
#60280000000
0!
0*
09
0>
0C
#60290000000
1!
1*
b10 6
19
1>
1C
b10 G
#60300000000
0!
0*
09
0>
0C
#60310000000
1!
1*
b11 6
19
1>
1C
b11 G
#60320000000
0!
0*
09
0>
0C
#60330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#60340000000
0!
0*
09
0>
0C
#60350000000
1!
1*
b101 6
19
1>
1C
b101 G
#60360000000
0!
0*
09
0>
0C
#60370000000
1!
1*
b110 6
19
1>
1C
b110 G
#60380000000
0!
0*
09
0>
0C
#60390000000
1!
1*
b111 6
19
1>
1C
b111 G
#60400000000
0!
0*
09
0>
0C
#60410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#60420000000
0!
0*
09
0>
0C
#60430000000
1!
1*
b1 6
19
1>
1C
b1 G
#60440000000
0!
0*
09
0>
0C
#60450000000
1!
1*
b10 6
19
1>
1C
b10 G
#60460000000
0!
0*
09
0>
0C
#60470000000
1!
1*
b11 6
19
1>
1C
b11 G
#60480000000
0!
0*
09
0>
0C
#60490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#60500000000
0!
0*
09
0>
0C
#60510000000
1!
1*
b101 6
19
1>
1C
b101 G
#60520000000
0!
0*
09
0>
0C
#60530000000
1!
1*
b110 6
19
1>
1C
b110 G
#60540000000
0!
0*
09
0>
0C
#60550000000
1!
1*
b111 6
19
1>
1C
b111 G
#60560000000
0!
1"
0*
1+
09
1:
0>
0C
#60570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#60580000000
0!
0*
09
0>
0C
#60590000000
1!
1*
b1 6
19
1>
1C
b1 G
#60600000000
0!
0*
09
0>
0C
#60610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#60620000000
0!
0*
09
0>
0C
#60630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#60640000000
0!
0*
09
0>
0C
#60650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#60660000000
0!
0*
09
0>
0C
#60670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#60680000000
0!
0#
0*
0,
09
0>
0?
0C
#60690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#60700000000
0!
0*
09
0>
0C
#60710000000
1!
1*
19
1>
1C
#60720000000
0!
0*
09
0>
0C
#60730000000
1!
1*
19
1>
1C
#60740000000
0!
0*
09
0>
0C
#60750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#60760000000
0!
0*
09
0>
0C
#60770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#60780000000
0!
0*
09
0>
0C
#60790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#60800000000
0!
0*
09
0>
0C
#60810000000
1!
1*
b10 6
19
1>
1C
b10 G
#60820000000
0!
0*
09
0>
0C
#60830000000
1!
1*
b11 6
19
1>
1C
b11 G
#60840000000
0!
0*
09
0>
0C
#60850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#60860000000
0!
0*
09
0>
0C
#60870000000
1!
1*
b101 6
19
1>
1C
b101 G
#60880000000
0!
0*
09
0>
0C
#60890000000
1!
1*
b110 6
19
1>
1C
b110 G
#60900000000
0!
0*
09
0>
0C
#60910000000
1!
1*
b111 6
19
1>
1C
b111 G
#60920000000
0!
0*
09
0>
0C
#60930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#60940000000
0!
0*
09
0>
0C
#60950000000
1!
1*
b1 6
19
1>
1C
b1 G
#60960000000
0!
0*
09
0>
0C
#60970000000
1!
1*
b10 6
19
1>
1C
b10 G
#60980000000
0!
0*
09
0>
0C
#60990000000
1!
1*
b11 6
19
1>
1C
b11 G
#61000000000
0!
0*
09
0>
0C
#61010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#61020000000
0!
0*
09
0>
0C
#61030000000
1!
1*
b101 6
19
1>
1C
b101 G
#61040000000
0!
0*
09
0>
0C
#61050000000
1!
1*
b110 6
19
1>
1C
b110 G
#61060000000
0!
0*
09
0>
0C
#61070000000
1!
1*
b111 6
19
1>
1C
b111 G
#61080000000
0!
0*
09
0>
0C
#61090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#61100000000
0!
0*
09
0>
0C
#61110000000
1!
1*
b1 6
19
1>
1C
b1 G
#61120000000
0!
0*
09
0>
0C
#61130000000
1!
1*
b10 6
19
1>
1C
b10 G
#61140000000
0!
0*
09
0>
0C
#61150000000
1!
1*
b11 6
19
1>
1C
b11 G
#61160000000
0!
0*
09
0>
0C
#61170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#61180000000
0!
0*
09
0>
0C
#61190000000
1!
1*
b101 6
19
1>
1C
b101 G
#61200000000
0!
0*
09
0>
0C
#61210000000
1!
1*
b110 6
19
1>
1C
b110 G
#61220000000
0!
0*
09
0>
0C
#61230000000
1!
1*
b111 6
19
1>
1C
b111 G
#61240000000
0!
1"
0*
1+
09
1:
0>
0C
#61250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#61260000000
0!
0*
09
0>
0C
#61270000000
1!
1*
b1 6
19
1>
1C
b1 G
#61280000000
0!
0*
09
0>
0C
#61290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#61300000000
0!
0*
09
0>
0C
#61310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#61320000000
0!
0*
09
0>
0C
#61330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#61340000000
0!
0*
09
0>
0C
#61350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#61360000000
0!
0#
0*
0,
09
0>
0?
0C
#61370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#61380000000
0!
0*
09
0>
0C
#61390000000
1!
1*
19
1>
1C
#61400000000
0!
0*
09
0>
0C
#61410000000
1!
1*
19
1>
1C
#61420000000
0!
0*
09
0>
0C
#61430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#61440000000
0!
0*
09
0>
0C
#61450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#61460000000
0!
0*
09
0>
0C
#61470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#61480000000
0!
0*
09
0>
0C
#61490000000
1!
1*
b10 6
19
1>
1C
b10 G
#61500000000
0!
0*
09
0>
0C
#61510000000
1!
1*
b11 6
19
1>
1C
b11 G
#61520000000
0!
0*
09
0>
0C
#61530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#61540000000
0!
0*
09
0>
0C
#61550000000
1!
1*
b101 6
19
1>
1C
b101 G
#61560000000
0!
0*
09
0>
0C
#61570000000
1!
1*
b110 6
19
1>
1C
b110 G
#61580000000
0!
0*
09
0>
0C
#61590000000
1!
1*
b111 6
19
1>
1C
b111 G
#61600000000
0!
0*
09
0>
0C
#61610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#61620000000
0!
0*
09
0>
0C
#61630000000
1!
1*
b1 6
19
1>
1C
b1 G
#61640000000
0!
0*
09
0>
0C
#61650000000
1!
1*
b10 6
19
1>
1C
b10 G
#61660000000
0!
0*
09
0>
0C
#61670000000
1!
1*
b11 6
19
1>
1C
b11 G
#61680000000
0!
0*
09
0>
0C
#61690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#61700000000
0!
0*
09
0>
0C
#61710000000
1!
1*
b101 6
19
1>
1C
b101 G
#61720000000
0!
0*
09
0>
0C
#61730000000
1!
1*
b110 6
19
1>
1C
b110 G
#61740000000
0!
0*
09
0>
0C
#61750000000
1!
1*
b111 6
19
1>
1C
b111 G
#61760000000
0!
0*
09
0>
0C
#61770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#61780000000
0!
0*
09
0>
0C
#61790000000
1!
1*
b1 6
19
1>
1C
b1 G
#61800000000
0!
0*
09
0>
0C
#61810000000
1!
1*
b10 6
19
1>
1C
b10 G
#61820000000
0!
0*
09
0>
0C
#61830000000
1!
1*
b11 6
19
1>
1C
b11 G
#61840000000
0!
0*
09
0>
0C
#61850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#61860000000
0!
0*
09
0>
0C
#61870000000
1!
1*
b101 6
19
1>
1C
b101 G
#61880000000
0!
0*
09
0>
0C
#61890000000
1!
1*
b110 6
19
1>
1C
b110 G
#61900000000
0!
0*
09
0>
0C
#61910000000
1!
1*
b111 6
19
1>
1C
b111 G
#61920000000
0!
1"
0*
1+
09
1:
0>
0C
#61930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#61940000000
0!
0*
09
0>
0C
#61950000000
1!
1*
b1 6
19
1>
1C
b1 G
#61960000000
0!
0*
09
0>
0C
#61970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#61980000000
0!
0*
09
0>
0C
#61990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#62000000000
0!
0*
09
0>
0C
#62010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#62020000000
0!
0*
09
0>
0C
#62030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#62040000000
0!
0#
0*
0,
09
0>
0?
0C
#62050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#62060000000
0!
0*
09
0>
0C
#62070000000
1!
1*
19
1>
1C
#62080000000
0!
0*
09
0>
0C
#62090000000
1!
1*
19
1>
1C
#62100000000
0!
0*
09
0>
0C
#62110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#62120000000
0!
0*
09
0>
0C
#62130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#62140000000
0!
0*
09
0>
0C
#62150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#62160000000
0!
0*
09
0>
0C
#62170000000
1!
1*
b10 6
19
1>
1C
b10 G
#62180000000
0!
0*
09
0>
0C
#62190000000
1!
1*
b11 6
19
1>
1C
b11 G
#62200000000
0!
0*
09
0>
0C
#62210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#62220000000
0!
0*
09
0>
0C
#62230000000
1!
1*
b101 6
19
1>
1C
b101 G
#62240000000
0!
0*
09
0>
0C
#62250000000
1!
1*
b110 6
19
1>
1C
b110 G
#62260000000
0!
0*
09
0>
0C
#62270000000
1!
1*
b111 6
19
1>
1C
b111 G
#62280000000
0!
0*
09
0>
0C
#62290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#62300000000
0!
0*
09
0>
0C
#62310000000
1!
1*
b1 6
19
1>
1C
b1 G
#62320000000
0!
0*
09
0>
0C
#62330000000
1!
1*
b10 6
19
1>
1C
b10 G
#62340000000
0!
0*
09
0>
0C
#62350000000
1!
1*
b11 6
19
1>
1C
b11 G
#62360000000
0!
0*
09
0>
0C
#62370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#62380000000
0!
0*
09
0>
0C
#62390000000
1!
1*
b101 6
19
1>
1C
b101 G
#62400000000
0!
0*
09
0>
0C
#62410000000
1!
1*
b110 6
19
1>
1C
b110 G
#62420000000
0!
0*
09
0>
0C
#62430000000
1!
1*
b111 6
19
1>
1C
b111 G
#62440000000
0!
0*
09
0>
0C
#62450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#62460000000
0!
0*
09
0>
0C
#62470000000
1!
1*
b1 6
19
1>
1C
b1 G
#62480000000
0!
0*
09
0>
0C
#62490000000
1!
1*
b10 6
19
1>
1C
b10 G
#62500000000
0!
0*
09
0>
0C
#62510000000
1!
1*
b11 6
19
1>
1C
b11 G
#62520000000
0!
0*
09
0>
0C
#62530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#62540000000
0!
0*
09
0>
0C
#62550000000
1!
1*
b101 6
19
1>
1C
b101 G
#62560000000
0!
0*
09
0>
0C
#62570000000
1!
1*
b110 6
19
1>
1C
b110 G
#62580000000
0!
0*
09
0>
0C
#62590000000
1!
1*
b111 6
19
1>
1C
b111 G
#62600000000
0!
1"
0*
1+
09
1:
0>
0C
#62610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#62620000000
0!
0*
09
0>
0C
#62630000000
1!
1*
b1 6
19
1>
1C
b1 G
#62640000000
0!
0*
09
0>
0C
#62650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#62660000000
0!
0*
09
0>
0C
#62670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#62680000000
0!
0*
09
0>
0C
#62690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#62700000000
0!
0*
09
0>
0C
#62710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#62720000000
0!
0#
0*
0,
09
0>
0?
0C
#62730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#62740000000
0!
0*
09
0>
0C
#62750000000
1!
1*
19
1>
1C
#62760000000
0!
0*
09
0>
0C
#62770000000
1!
1*
19
1>
1C
#62780000000
0!
0*
09
0>
0C
#62790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#62800000000
0!
0*
09
0>
0C
#62810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#62820000000
0!
0*
09
0>
0C
#62830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#62840000000
0!
0*
09
0>
0C
#62850000000
1!
1*
b10 6
19
1>
1C
b10 G
#62860000000
0!
0*
09
0>
0C
#62870000000
1!
1*
b11 6
19
1>
1C
b11 G
#62880000000
0!
0*
09
0>
0C
#62890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#62900000000
0!
0*
09
0>
0C
#62910000000
1!
1*
b101 6
19
1>
1C
b101 G
#62920000000
0!
0*
09
0>
0C
#62930000000
1!
1*
b110 6
19
1>
1C
b110 G
#62940000000
0!
0*
09
0>
0C
#62950000000
1!
1*
b111 6
19
1>
1C
b111 G
#62960000000
0!
0*
09
0>
0C
#62970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#62980000000
0!
0*
09
0>
0C
#62990000000
1!
1*
b1 6
19
1>
1C
b1 G
#63000000000
0!
0*
09
0>
0C
#63010000000
1!
1*
b10 6
19
1>
1C
b10 G
#63020000000
0!
0*
09
0>
0C
#63030000000
1!
1*
b11 6
19
1>
1C
b11 G
#63040000000
0!
0*
09
0>
0C
#63050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#63060000000
0!
0*
09
0>
0C
#63070000000
1!
1*
b101 6
19
1>
1C
b101 G
#63080000000
0!
0*
09
0>
0C
#63090000000
1!
1*
b110 6
19
1>
1C
b110 G
#63100000000
0!
0*
09
0>
0C
#63110000000
1!
1*
b111 6
19
1>
1C
b111 G
#63120000000
0!
0*
09
0>
0C
#63130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#63140000000
0!
0*
09
0>
0C
#63150000000
1!
1*
b1 6
19
1>
1C
b1 G
#63160000000
0!
0*
09
0>
0C
#63170000000
1!
1*
b10 6
19
1>
1C
b10 G
#63180000000
0!
0*
09
0>
0C
#63190000000
1!
1*
b11 6
19
1>
1C
b11 G
#63200000000
0!
0*
09
0>
0C
#63210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#63220000000
0!
0*
09
0>
0C
#63230000000
1!
1*
b101 6
19
1>
1C
b101 G
#63240000000
0!
0*
09
0>
0C
#63250000000
1!
1*
b110 6
19
1>
1C
b110 G
#63260000000
0!
0*
09
0>
0C
#63270000000
1!
1*
b111 6
19
1>
1C
b111 G
#63280000000
0!
1"
0*
1+
09
1:
0>
0C
#63290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#63300000000
0!
0*
09
0>
0C
#63310000000
1!
1*
b1 6
19
1>
1C
b1 G
#63320000000
0!
0*
09
0>
0C
#63330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#63340000000
0!
0*
09
0>
0C
#63350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#63360000000
0!
0*
09
0>
0C
#63370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#63380000000
0!
0*
09
0>
0C
#63390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#63400000000
0!
0#
0*
0,
09
0>
0?
0C
#63410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#63420000000
0!
0*
09
0>
0C
#63430000000
1!
1*
19
1>
1C
#63440000000
0!
0*
09
0>
0C
#63450000000
1!
1*
19
1>
1C
#63460000000
0!
0*
09
0>
0C
#63470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#63480000000
0!
0*
09
0>
0C
#63490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#63500000000
0!
0*
09
0>
0C
#63510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#63520000000
0!
0*
09
0>
0C
#63530000000
1!
1*
b10 6
19
1>
1C
b10 G
#63540000000
0!
0*
09
0>
0C
#63550000000
1!
1*
b11 6
19
1>
1C
b11 G
#63560000000
0!
0*
09
0>
0C
#63570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#63580000000
0!
0*
09
0>
0C
#63590000000
1!
1*
b101 6
19
1>
1C
b101 G
#63600000000
0!
0*
09
0>
0C
#63610000000
1!
1*
b110 6
19
1>
1C
b110 G
#63620000000
0!
0*
09
0>
0C
#63630000000
1!
1*
b111 6
19
1>
1C
b111 G
#63640000000
0!
0*
09
0>
0C
#63650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#63660000000
0!
0*
09
0>
0C
#63670000000
1!
1*
b1 6
19
1>
1C
b1 G
#63680000000
0!
0*
09
0>
0C
#63690000000
1!
1*
b10 6
19
1>
1C
b10 G
#63700000000
0!
0*
09
0>
0C
#63710000000
1!
1*
b11 6
19
1>
1C
b11 G
#63720000000
0!
0*
09
0>
0C
#63730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#63740000000
0!
0*
09
0>
0C
#63750000000
1!
1*
b101 6
19
1>
1C
b101 G
#63760000000
0!
0*
09
0>
0C
#63770000000
1!
1*
b110 6
19
1>
1C
b110 G
#63780000000
0!
0*
09
0>
0C
#63790000000
1!
1*
b111 6
19
1>
1C
b111 G
#63800000000
0!
0*
09
0>
0C
#63810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#63820000000
0!
0*
09
0>
0C
#63830000000
1!
1*
b1 6
19
1>
1C
b1 G
#63840000000
0!
0*
09
0>
0C
#63850000000
1!
1*
b10 6
19
1>
1C
b10 G
#63860000000
0!
0*
09
0>
0C
#63870000000
1!
1*
b11 6
19
1>
1C
b11 G
#63880000000
0!
0*
09
0>
0C
#63890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#63900000000
0!
0*
09
0>
0C
#63910000000
1!
1*
b101 6
19
1>
1C
b101 G
#63920000000
0!
0*
09
0>
0C
#63930000000
1!
1*
b110 6
19
1>
1C
b110 G
#63940000000
0!
0*
09
0>
0C
#63950000000
1!
1*
b111 6
19
1>
1C
b111 G
#63960000000
0!
1"
0*
1+
09
1:
0>
0C
#63970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#63980000000
0!
0*
09
0>
0C
#63990000000
1!
1*
b1 6
19
1>
1C
b1 G
#64000000000
0!
0*
09
0>
0C
#64010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#64020000000
0!
0*
09
0>
0C
#64030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#64040000000
0!
0*
09
0>
0C
#64050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#64060000000
0!
0*
09
0>
0C
#64070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#64080000000
0!
0#
0*
0,
09
0>
0?
0C
#64090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#64100000000
0!
0*
09
0>
0C
#64110000000
1!
1*
19
1>
1C
#64120000000
0!
0*
09
0>
0C
#64130000000
1!
1*
19
1>
1C
#64140000000
0!
0*
09
0>
0C
#64150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#64160000000
0!
0*
09
0>
0C
#64170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#64180000000
0!
0*
09
0>
0C
#64190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#64200000000
0!
0*
09
0>
0C
#64210000000
1!
1*
b10 6
19
1>
1C
b10 G
#64220000000
0!
0*
09
0>
0C
#64230000000
1!
1*
b11 6
19
1>
1C
b11 G
#64240000000
0!
0*
09
0>
0C
#64250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#64260000000
0!
0*
09
0>
0C
#64270000000
1!
1*
b101 6
19
1>
1C
b101 G
#64280000000
0!
0*
09
0>
0C
#64290000000
1!
1*
b110 6
19
1>
1C
b110 G
#64300000000
0!
0*
09
0>
0C
#64310000000
1!
1*
b111 6
19
1>
1C
b111 G
#64320000000
0!
0*
09
0>
0C
#64330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#64340000000
0!
0*
09
0>
0C
#64350000000
1!
1*
b1 6
19
1>
1C
b1 G
#64360000000
0!
0*
09
0>
0C
#64370000000
1!
1*
b10 6
19
1>
1C
b10 G
#64380000000
0!
0*
09
0>
0C
#64390000000
1!
1*
b11 6
19
1>
1C
b11 G
#64400000000
0!
0*
09
0>
0C
#64410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#64420000000
0!
0*
09
0>
0C
#64430000000
1!
1*
b101 6
19
1>
1C
b101 G
#64440000000
0!
0*
09
0>
0C
#64450000000
1!
1*
b110 6
19
1>
1C
b110 G
#64460000000
0!
0*
09
0>
0C
#64470000000
1!
1*
b111 6
19
1>
1C
b111 G
#64480000000
0!
0*
09
0>
0C
#64490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#64500000000
0!
0*
09
0>
0C
#64510000000
1!
1*
b1 6
19
1>
1C
b1 G
#64520000000
0!
0*
09
0>
0C
#64530000000
1!
1*
b10 6
19
1>
1C
b10 G
#64540000000
0!
0*
09
0>
0C
#64550000000
1!
1*
b11 6
19
1>
1C
b11 G
#64560000000
0!
0*
09
0>
0C
#64570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#64580000000
0!
0*
09
0>
0C
#64590000000
1!
1*
b101 6
19
1>
1C
b101 G
#64600000000
0!
0*
09
0>
0C
#64610000000
1!
1*
b110 6
19
1>
1C
b110 G
#64620000000
0!
0*
09
0>
0C
#64630000000
1!
1*
b111 6
19
1>
1C
b111 G
#64640000000
0!
1"
0*
1+
09
1:
0>
0C
#64650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#64660000000
0!
0*
09
0>
0C
#64670000000
1!
1*
b1 6
19
1>
1C
b1 G
#64680000000
0!
0*
09
0>
0C
#64690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#64700000000
0!
0*
09
0>
0C
#64710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#64720000000
0!
0*
09
0>
0C
#64730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#64740000000
0!
0*
09
0>
0C
#64750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#64760000000
0!
0#
0*
0,
09
0>
0?
0C
#64770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#64780000000
0!
0*
09
0>
0C
#64790000000
1!
1*
19
1>
1C
#64800000000
0!
0*
09
0>
0C
#64810000000
1!
1*
19
1>
1C
#64820000000
0!
0*
09
0>
0C
#64830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#64840000000
0!
0*
09
0>
0C
#64850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#64860000000
0!
0*
09
0>
0C
#64870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#64880000000
0!
0*
09
0>
0C
#64890000000
1!
1*
b10 6
19
1>
1C
b10 G
#64900000000
0!
0*
09
0>
0C
#64910000000
1!
1*
b11 6
19
1>
1C
b11 G
#64920000000
0!
0*
09
0>
0C
#64930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#64940000000
0!
0*
09
0>
0C
#64950000000
1!
1*
b101 6
19
1>
1C
b101 G
#64960000000
0!
0*
09
0>
0C
#64970000000
1!
1*
b110 6
19
1>
1C
b110 G
#64980000000
0!
0*
09
0>
0C
#64990000000
1!
1*
b111 6
19
1>
1C
b111 G
#65000000000
0!
0*
09
0>
0C
#65010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#65020000000
0!
0*
09
0>
0C
#65030000000
1!
1*
b1 6
19
1>
1C
b1 G
#65040000000
0!
0*
09
0>
0C
#65050000000
1!
1*
b10 6
19
1>
1C
b10 G
#65060000000
0!
0*
09
0>
0C
#65070000000
1!
1*
b11 6
19
1>
1C
b11 G
#65080000000
0!
0*
09
0>
0C
#65090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#65100000000
0!
0*
09
0>
0C
#65110000000
1!
1*
b101 6
19
1>
1C
b101 G
#65120000000
0!
0*
09
0>
0C
#65130000000
1!
1*
b110 6
19
1>
1C
b110 G
#65140000000
0!
0*
09
0>
0C
#65150000000
1!
1*
b111 6
19
1>
1C
b111 G
#65160000000
0!
0*
09
0>
0C
#65170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#65180000000
0!
0*
09
0>
0C
#65190000000
1!
1*
b1 6
19
1>
1C
b1 G
#65200000000
0!
0*
09
0>
0C
#65210000000
1!
1*
b10 6
19
1>
1C
b10 G
#65220000000
0!
0*
09
0>
0C
#65230000000
1!
1*
b11 6
19
1>
1C
b11 G
#65240000000
0!
0*
09
0>
0C
#65250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#65260000000
0!
0*
09
0>
0C
#65270000000
1!
1*
b101 6
19
1>
1C
b101 G
#65280000000
0!
0*
09
0>
0C
#65290000000
1!
1*
b110 6
19
1>
1C
b110 G
#65300000000
0!
0*
09
0>
0C
#65310000000
1!
1*
b111 6
19
1>
1C
b111 G
#65320000000
0!
1"
0*
1+
09
1:
0>
0C
#65330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#65340000000
0!
0*
09
0>
0C
#65350000000
1!
1*
b1 6
19
1>
1C
b1 G
#65360000000
0!
0*
09
0>
0C
#65370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#65380000000
0!
0*
09
0>
0C
#65390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#65400000000
0!
0*
09
0>
0C
#65410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#65420000000
0!
0*
09
0>
0C
#65430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#65440000000
0!
0#
0*
0,
09
0>
0?
0C
#65450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#65460000000
0!
0*
09
0>
0C
#65470000000
1!
1*
19
1>
1C
#65480000000
0!
0*
09
0>
0C
#65490000000
1!
1*
19
1>
1C
#65500000000
0!
0*
09
0>
0C
#65510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#65520000000
0!
0*
09
0>
0C
#65530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#65540000000
0!
0*
09
0>
0C
#65550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#65560000000
0!
0*
09
0>
0C
#65570000000
1!
1*
b10 6
19
1>
1C
b10 G
#65580000000
0!
0*
09
0>
0C
#65590000000
1!
1*
b11 6
19
1>
1C
b11 G
#65600000000
0!
0*
09
0>
0C
#65610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#65620000000
0!
0*
09
0>
0C
#65630000000
1!
1*
b101 6
19
1>
1C
b101 G
#65640000000
0!
0*
09
0>
0C
#65650000000
1!
1*
b110 6
19
1>
1C
b110 G
#65660000000
0!
0*
09
0>
0C
#65670000000
1!
1*
b111 6
19
1>
1C
b111 G
#65680000000
0!
0*
09
0>
0C
#65690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#65700000000
0!
0*
09
0>
0C
#65710000000
1!
1*
b1 6
19
1>
1C
b1 G
#65720000000
0!
0*
09
0>
0C
#65730000000
1!
1*
b10 6
19
1>
1C
b10 G
#65740000000
0!
0*
09
0>
0C
#65750000000
1!
1*
b11 6
19
1>
1C
b11 G
#65760000000
0!
0*
09
0>
0C
#65770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#65780000000
0!
0*
09
0>
0C
#65790000000
1!
1*
b101 6
19
1>
1C
b101 G
#65800000000
0!
0*
09
0>
0C
#65810000000
1!
1*
b110 6
19
1>
1C
b110 G
#65820000000
0!
0*
09
0>
0C
#65830000000
1!
1*
b111 6
19
1>
1C
b111 G
#65840000000
0!
0*
09
0>
0C
#65850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#65860000000
0!
0*
09
0>
0C
#65870000000
1!
1*
b1 6
19
1>
1C
b1 G
#65880000000
0!
0*
09
0>
0C
#65890000000
1!
1*
b10 6
19
1>
1C
b10 G
#65900000000
0!
0*
09
0>
0C
#65910000000
1!
1*
b11 6
19
1>
1C
b11 G
#65920000000
0!
0*
09
0>
0C
#65930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#65940000000
0!
0*
09
0>
0C
#65950000000
1!
1*
b101 6
19
1>
1C
b101 G
#65960000000
0!
0*
09
0>
0C
#65970000000
1!
1*
b110 6
19
1>
1C
b110 G
#65980000000
0!
0*
09
0>
0C
#65990000000
1!
1*
b111 6
19
1>
1C
b111 G
#66000000000
0!
1"
0*
1+
09
1:
0>
0C
#66010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#66020000000
0!
0*
09
0>
0C
#66030000000
1!
1*
b1 6
19
1>
1C
b1 G
#66040000000
0!
0*
09
0>
0C
#66050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#66060000000
0!
0*
09
0>
0C
#66070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#66080000000
0!
0*
09
0>
0C
#66090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#66100000000
0!
0*
09
0>
0C
#66110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#66120000000
0!
0#
0*
0,
09
0>
0?
0C
#66130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#66140000000
0!
0*
09
0>
0C
#66150000000
1!
1*
19
1>
1C
#66160000000
0!
0*
09
0>
0C
#66170000000
1!
1*
19
1>
1C
#66180000000
0!
0*
09
0>
0C
#66190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#66200000000
0!
0*
09
0>
0C
#66210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#66220000000
0!
0*
09
0>
0C
#66230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#66240000000
0!
0*
09
0>
0C
#66250000000
1!
1*
b10 6
19
1>
1C
b10 G
#66260000000
0!
0*
09
0>
0C
#66270000000
1!
1*
b11 6
19
1>
1C
b11 G
#66280000000
0!
0*
09
0>
0C
#66290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#66300000000
0!
0*
09
0>
0C
#66310000000
1!
1*
b101 6
19
1>
1C
b101 G
#66320000000
0!
0*
09
0>
0C
#66330000000
1!
1*
b110 6
19
1>
1C
b110 G
#66340000000
0!
0*
09
0>
0C
#66350000000
1!
1*
b111 6
19
1>
1C
b111 G
#66360000000
0!
0*
09
0>
0C
#66370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#66380000000
0!
0*
09
0>
0C
#66390000000
1!
1*
b1 6
19
1>
1C
b1 G
#66400000000
0!
0*
09
0>
0C
#66410000000
1!
1*
b10 6
19
1>
1C
b10 G
#66420000000
0!
0*
09
0>
0C
#66430000000
1!
1*
b11 6
19
1>
1C
b11 G
#66440000000
0!
0*
09
0>
0C
#66450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#66460000000
0!
0*
09
0>
0C
#66470000000
1!
1*
b101 6
19
1>
1C
b101 G
#66480000000
0!
0*
09
0>
0C
#66490000000
1!
1*
b110 6
19
1>
1C
b110 G
#66500000000
0!
0*
09
0>
0C
#66510000000
1!
1*
b111 6
19
1>
1C
b111 G
#66520000000
0!
0*
09
0>
0C
#66530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#66540000000
0!
0*
09
0>
0C
#66550000000
1!
1*
b1 6
19
1>
1C
b1 G
#66560000000
0!
0*
09
0>
0C
#66570000000
1!
1*
b10 6
19
1>
1C
b10 G
#66580000000
0!
0*
09
0>
0C
#66590000000
1!
1*
b11 6
19
1>
1C
b11 G
#66600000000
0!
0*
09
0>
0C
#66610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#66620000000
0!
0*
09
0>
0C
#66630000000
1!
1*
b101 6
19
1>
1C
b101 G
#66640000000
0!
0*
09
0>
0C
#66650000000
1!
1*
b110 6
19
1>
1C
b110 G
#66660000000
0!
0*
09
0>
0C
#66670000000
1!
1*
b111 6
19
1>
1C
b111 G
#66680000000
0!
1"
0*
1+
09
1:
0>
0C
#66690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#66700000000
0!
0*
09
0>
0C
#66710000000
1!
1*
b1 6
19
1>
1C
b1 G
#66720000000
0!
0*
09
0>
0C
#66730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#66740000000
0!
0*
09
0>
0C
#66750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#66760000000
0!
0*
09
0>
0C
#66770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#66780000000
0!
0*
09
0>
0C
#66790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#66800000000
0!
0#
0*
0,
09
0>
0?
0C
#66810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#66820000000
0!
0*
09
0>
0C
#66830000000
1!
1*
19
1>
1C
#66840000000
0!
0*
09
0>
0C
#66850000000
1!
1*
19
1>
1C
#66860000000
0!
0*
09
0>
0C
#66870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#66880000000
0!
0*
09
0>
0C
#66890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#66900000000
0!
0*
09
0>
0C
#66910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#66920000000
0!
0*
09
0>
0C
#66930000000
1!
1*
b10 6
19
1>
1C
b10 G
#66940000000
0!
0*
09
0>
0C
#66950000000
1!
1*
b11 6
19
1>
1C
b11 G
#66960000000
0!
0*
09
0>
0C
#66970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#66980000000
0!
0*
09
0>
0C
#66990000000
1!
1*
b101 6
19
1>
1C
b101 G
#67000000000
0!
0*
09
0>
0C
#67010000000
1!
1*
b110 6
19
1>
1C
b110 G
#67020000000
0!
0*
09
0>
0C
#67030000000
1!
1*
b111 6
19
1>
1C
b111 G
#67040000000
0!
0*
09
0>
0C
#67050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#67060000000
0!
0*
09
0>
0C
#67070000000
1!
1*
b1 6
19
1>
1C
b1 G
#67080000000
0!
0*
09
0>
0C
#67090000000
1!
1*
b10 6
19
1>
1C
b10 G
#67100000000
0!
0*
09
0>
0C
#67110000000
1!
1*
b11 6
19
1>
1C
b11 G
#67120000000
0!
0*
09
0>
0C
#67130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#67140000000
0!
0*
09
0>
0C
#67150000000
1!
1*
b101 6
19
1>
1C
b101 G
#67160000000
0!
0*
09
0>
0C
#67170000000
1!
1*
b110 6
19
1>
1C
b110 G
#67180000000
0!
0*
09
0>
0C
#67190000000
1!
1*
b111 6
19
1>
1C
b111 G
#67200000000
0!
0*
09
0>
0C
#67210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#67220000000
0!
0*
09
0>
0C
#67230000000
1!
1*
b1 6
19
1>
1C
b1 G
#67240000000
0!
0*
09
0>
0C
#67250000000
1!
1*
b10 6
19
1>
1C
b10 G
#67260000000
0!
0*
09
0>
0C
#67270000000
1!
1*
b11 6
19
1>
1C
b11 G
#67280000000
0!
0*
09
0>
0C
#67290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#67300000000
0!
0*
09
0>
0C
#67310000000
1!
1*
b101 6
19
1>
1C
b101 G
#67320000000
0!
0*
09
0>
0C
#67330000000
1!
1*
b110 6
19
1>
1C
b110 G
#67340000000
0!
0*
09
0>
0C
#67350000000
1!
1*
b111 6
19
1>
1C
b111 G
#67360000000
0!
1"
0*
1+
09
1:
0>
0C
#67370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#67380000000
0!
0*
09
0>
0C
#67390000000
1!
1*
b1 6
19
1>
1C
b1 G
#67400000000
0!
0*
09
0>
0C
#67410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#67420000000
0!
0*
09
0>
0C
#67430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#67440000000
0!
0*
09
0>
0C
#67450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#67460000000
0!
0*
09
0>
0C
#67470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#67480000000
0!
0#
0*
0,
09
0>
0?
0C
#67490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#67500000000
0!
0*
09
0>
0C
#67510000000
1!
1*
19
1>
1C
#67520000000
0!
0*
09
0>
0C
#67530000000
1!
1*
19
1>
1C
#67540000000
0!
0*
09
0>
0C
#67550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#67560000000
0!
0*
09
0>
0C
#67570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#67580000000
0!
0*
09
0>
0C
#67590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#67600000000
0!
0*
09
0>
0C
#67610000000
1!
1*
b10 6
19
1>
1C
b10 G
#67620000000
0!
0*
09
0>
0C
#67630000000
1!
1*
b11 6
19
1>
1C
b11 G
#67640000000
0!
0*
09
0>
0C
#67650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#67660000000
0!
0*
09
0>
0C
#67670000000
1!
1*
b101 6
19
1>
1C
b101 G
#67680000000
0!
0*
09
0>
0C
#67690000000
1!
1*
b110 6
19
1>
1C
b110 G
#67700000000
0!
0*
09
0>
0C
#67710000000
1!
1*
b111 6
19
1>
1C
b111 G
#67720000000
0!
0*
09
0>
0C
#67730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#67740000000
0!
0*
09
0>
0C
#67750000000
1!
1*
b1 6
19
1>
1C
b1 G
#67760000000
0!
0*
09
0>
0C
#67770000000
1!
1*
b10 6
19
1>
1C
b10 G
#67780000000
0!
0*
09
0>
0C
#67790000000
1!
1*
b11 6
19
1>
1C
b11 G
#67800000000
0!
0*
09
0>
0C
#67810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#67820000000
0!
0*
09
0>
0C
#67830000000
1!
1*
b101 6
19
1>
1C
b101 G
#67840000000
0!
0*
09
0>
0C
#67850000000
1!
1*
b110 6
19
1>
1C
b110 G
#67860000000
0!
0*
09
0>
0C
#67870000000
1!
1*
b111 6
19
1>
1C
b111 G
#67880000000
0!
0*
09
0>
0C
#67890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#67900000000
0!
0*
09
0>
0C
#67910000000
1!
1*
b1 6
19
1>
1C
b1 G
#67920000000
0!
0*
09
0>
0C
#67930000000
1!
1*
b10 6
19
1>
1C
b10 G
#67940000000
0!
0*
09
0>
0C
#67950000000
1!
1*
b11 6
19
1>
1C
b11 G
#67960000000
0!
0*
09
0>
0C
#67970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#67980000000
0!
0*
09
0>
0C
#67990000000
1!
1*
b101 6
19
1>
1C
b101 G
#68000000000
0!
0*
09
0>
0C
#68010000000
1!
1*
b110 6
19
1>
1C
b110 G
#68020000000
0!
0*
09
0>
0C
#68030000000
1!
1*
b111 6
19
1>
1C
b111 G
#68040000000
0!
1"
0*
1+
09
1:
0>
0C
#68050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#68060000000
0!
0*
09
0>
0C
#68070000000
1!
1*
b1 6
19
1>
1C
b1 G
#68080000000
0!
0*
09
0>
0C
#68090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#68100000000
0!
0*
09
0>
0C
#68110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#68120000000
0!
0*
09
0>
0C
#68130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#68140000000
0!
0*
09
0>
0C
#68150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#68160000000
0!
0#
0*
0,
09
0>
0?
0C
#68170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#68180000000
0!
0*
09
0>
0C
#68190000000
1!
1*
19
1>
1C
#68200000000
0!
0*
09
0>
0C
#68210000000
1!
1*
19
1>
1C
#68220000000
0!
0*
09
0>
0C
#68230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#68240000000
0!
0*
09
0>
0C
#68250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#68260000000
0!
0*
09
0>
0C
#68270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#68280000000
0!
0*
09
0>
0C
#68290000000
1!
1*
b10 6
19
1>
1C
b10 G
#68300000000
0!
0*
09
0>
0C
#68310000000
1!
1*
b11 6
19
1>
1C
b11 G
#68320000000
0!
0*
09
0>
0C
#68330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#68340000000
0!
0*
09
0>
0C
#68350000000
1!
1*
b101 6
19
1>
1C
b101 G
#68360000000
0!
0*
09
0>
0C
#68370000000
1!
1*
b110 6
19
1>
1C
b110 G
#68380000000
0!
0*
09
0>
0C
#68390000000
1!
1*
b111 6
19
1>
1C
b111 G
#68400000000
0!
0*
09
0>
0C
#68410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#68420000000
0!
0*
09
0>
0C
#68430000000
1!
1*
b1 6
19
1>
1C
b1 G
#68440000000
0!
0*
09
0>
0C
#68450000000
1!
1*
b10 6
19
1>
1C
b10 G
#68460000000
0!
0*
09
0>
0C
#68470000000
1!
1*
b11 6
19
1>
1C
b11 G
#68480000000
0!
0*
09
0>
0C
#68490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#68500000000
0!
0*
09
0>
0C
#68510000000
1!
1*
b101 6
19
1>
1C
b101 G
#68520000000
0!
0*
09
0>
0C
#68530000000
1!
1*
b110 6
19
1>
1C
b110 G
#68540000000
0!
0*
09
0>
0C
#68550000000
1!
1*
b111 6
19
1>
1C
b111 G
#68560000000
0!
0*
09
0>
0C
#68570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#68580000000
0!
0*
09
0>
0C
#68590000000
1!
1*
b1 6
19
1>
1C
b1 G
#68600000000
0!
0*
09
0>
0C
#68610000000
1!
1*
b10 6
19
1>
1C
b10 G
#68620000000
0!
0*
09
0>
0C
#68630000000
1!
1*
b11 6
19
1>
1C
b11 G
#68640000000
0!
0*
09
0>
0C
#68650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#68660000000
0!
0*
09
0>
0C
#68670000000
1!
1*
b101 6
19
1>
1C
b101 G
#68680000000
0!
0*
09
0>
0C
#68690000000
1!
1*
b110 6
19
1>
1C
b110 G
#68700000000
0!
0*
09
0>
0C
#68710000000
1!
1*
b111 6
19
1>
1C
b111 G
#68720000000
0!
1"
0*
1+
09
1:
0>
0C
#68730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#68740000000
0!
0*
09
0>
0C
#68750000000
1!
1*
b1 6
19
1>
1C
b1 G
#68760000000
0!
0*
09
0>
0C
#68770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#68780000000
0!
0*
09
0>
0C
#68790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#68800000000
0!
0*
09
0>
0C
#68810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#68820000000
0!
0*
09
0>
0C
#68830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#68840000000
0!
0#
0*
0,
09
0>
0?
0C
#68850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#68860000000
0!
0*
09
0>
0C
#68870000000
1!
1*
19
1>
1C
#68880000000
0!
0*
09
0>
0C
#68890000000
1!
1*
19
1>
1C
#68900000000
0!
0*
09
0>
0C
#68910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#68920000000
0!
0*
09
0>
0C
#68930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#68940000000
0!
0*
09
0>
0C
#68950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#68960000000
0!
0*
09
0>
0C
#68970000000
1!
1*
b10 6
19
1>
1C
b10 G
#68980000000
0!
0*
09
0>
0C
#68990000000
1!
1*
b11 6
19
1>
1C
b11 G
#69000000000
0!
0*
09
0>
0C
#69010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#69020000000
0!
0*
09
0>
0C
#69030000000
1!
1*
b101 6
19
1>
1C
b101 G
#69040000000
0!
0*
09
0>
0C
#69050000000
1!
1*
b110 6
19
1>
1C
b110 G
#69060000000
0!
0*
09
0>
0C
#69070000000
1!
1*
b111 6
19
1>
1C
b111 G
#69080000000
0!
0*
09
0>
0C
#69090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#69100000000
0!
0*
09
0>
0C
#69110000000
1!
1*
b1 6
19
1>
1C
b1 G
#69120000000
0!
0*
09
0>
0C
#69130000000
1!
1*
b10 6
19
1>
1C
b10 G
#69140000000
0!
0*
09
0>
0C
#69150000000
1!
1*
b11 6
19
1>
1C
b11 G
#69160000000
0!
0*
09
0>
0C
#69170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#69180000000
0!
0*
09
0>
0C
#69190000000
1!
1*
b101 6
19
1>
1C
b101 G
#69200000000
0!
0*
09
0>
0C
#69210000000
1!
1*
b110 6
19
1>
1C
b110 G
#69220000000
0!
0*
09
0>
0C
#69230000000
1!
1*
b111 6
19
1>
1C
b111 G
#69240000000
0!
0*
09
0>
0C
#69250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#69260000000
0!
0*
09
0>
0C
#69270000000
1!
1*
b1 6
19
1>
1C
b1 G
#69280000000
0!
0*
09
0>
0C
#69290000000
1!
1*
b10 6
19
1>
1C
b10 G
#69300000000
0!
0*
09
0>
0C
#69310000000
1!
1*
b11 6
19
1>
1C
b11 G
#69320000000
0!
0*
09
0>
0C
#69330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#69340000000
0!
0*
09
0>
0C
#69350000000
1!
1*
b101 6
19
1>
1C
b101 G
#69360000000
0!
0*
09
0>
0C
#69370000000
1!
1*
b110 6
19
1>
1C
b110 G
#69380000000
0!
0*
09
0>
0C
#69390000000
1!
1*
b111 6
19
1>
1C
b111 G
#69400000000
0!
1"
0*
1+
09
1:
0>
0C
#69410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#69420000000
0!
0*
09
0>
0C
#69430000000
1!
1*
b1 6
19
1>
1C
b1 G
#69440000000
0!
0*
09
0>
0C
#69450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#69460000000
0!
0*
09
0>
0C
#69470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#69480000000
0!
0*
09
0>
0C
#69490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#69500000000
0!
0*
09
0>
0C
#69510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#69520000000
0!
0#
0*
0,
09
0>
0?
0C
#69530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#69540000000
0!
0*
09
0>
0C
#69550000000
1!
1*
19
1>
1C
#69560000000
0!
0*
09
0>
0C
#69570000000
1!
1*
19
1>
1C
#69580000000
0!
0*
09
0>
0C
#69590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#69600000000
0!
0*
09
0>
0C
#69610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#69620000000
0!
0*
09
0>
0C
#69630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#69640000000
0!
0*
09
0>
0C
#69650000000
1!
1*
b10 6
19
1>
1C
b10 G
#69660000000
0!
0*
09
0>
0C
#69670000000
1!
1*
b11 6
19
1>
1C
b11 G
#69680000000
0!
0*
09
0>
0C
#69690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#69700000000
0!
0*
09
0>
0C
#69710000000
1!
1*
b101 6
19
1>
1C
b101 G
#69720000000
0!
0*
09
0>
0C
#69730000000
1!
1*
b110 6
19
1>
1C
b110 G
#69740000000
0!
0*
09
0>
0C
#69750000000
1!
1*
b111 6
19
1>
1C
b111 G
#69760000000
0!
0*
09
0>
0C
#69770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#69780000000
0!
0*
09
0>
0C
#69790000000
1!
1*
b1 6
19
1>
1C
b1 G
#69800000000
0!
0*
09
0>
0C
#69810000000
1!
1*
b10 6
19
1>
1C
b10 G
#69820000000
0!
0*
09
0>
0C
#69830000000
1!
1*
b11 6
19
1>
1C
b11 G
#69840000000
0!
0*
09
0>
0C
#69850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#69860000000
0!
0*
09
0>
0C
#69870000000
1!
1*
b101 6
19
1>
1C
b101 G
#69880000000
0!
0*
09
0>
0C
#69890000000
1!
1*
b110 6
19
1>
1C
b110 G
#69900000000
0!
0*
09
0>
0C
#69910000000
1!
1*
b111 6
19
1>
1C
b111 G
#69920000000
0!
0*
09
0>
0C
#69930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#69940000000
0!
0*
09
0>
0C
#69950000000
1!
1*
b1 6
19
1>
1C
b1 G
#69960000000
0!
0*
09
0>
0C
#69970000000
1!
1*
b10 6
19
1>
1C
b10 G
#69980000000
0!
0*
09
0>
0C
#69990000000
1!
1*
b11 6
19
1>
1C
b11 G
#70000000000
0!
0*
09
0>
0C
#70010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#70020000000
0!
0*
09
0>
0C
#70030000000
1!
1*
b101 6
19
1>
1C
b101 G
#70040000000
0!
0*
09
0>
0C
#70050000000
1!
1*
b110 6
19
1>
1C
b110 G
#70060000000
0!
0*
09
0>
0C
#70070000000
1!
1*
b111 6
19
1>
1C
b111 G
#70080000000
0!
1"
0*
1+
09
1:
0>
0C
#70090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#70100000000
0!
0*
09
0>
0C
#70110000000
1!
1*
b1 6
19
1>
1C
b1 G
#70120000000
0!
0*
09
0>
0C
#70130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#70140000000
0!
0*
09
0>
0C
#70150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#70160000000
0!
0*
09
0>
0C
#70170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#70180000000
0!
0*
09
0>
0C
#70190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#70200000000
0!
0#
0*
0,
09
0>
0?
0C
#70210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#70220000000
0!
0*
09
0>
0C
#70230000000
1!
1*
19
1>
1C
#70240000000
0!
0*
09
0>
0C
#70250000000
1!
1*
19
1>
1C
#70260000000
0!
0*
09
0>
0C
#70270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#70280000000
0!
0*
09
0>
0C
#70290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#70300000000
0!
0*
09
0>
0C
#70310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#70320000000
0!
0*
09
0>
0C
#70330000000
1!
1*
b10 6
19
1>
1C
b10 G
#70340000000
0!
0*
09
0>
0C
#70350000000
1!
1*
b11 6
19
1>
1C
b11 G
#70360000000
0!
0*
09
0>
0C
#70370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#70380000000
0!
0*
09
0>
0C
#70390000000
1!
1*
b101 6
19
1>
1C
b101 G
#70400000000
0!
0*
09
0>
0C
#70410000000
1!
1*
b110 6
19
1>
1C
b110 G
#70420000000
0!
0*
09
0>
0C
#70430000000
1!
1*
b111 6
19
1>
1C
b111 G
#70440000000
0!
0*
09
0>
0C
#70450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#70460000000
0!
0*
09
0>
0C
#70470000000
1!
1*
b1 6
19
1>
1C
b1 G
#70480000000
0!
0*
09
0>
0C
#70490000000
1!
1*
b10 6
19
1>
1C
b10 G
#70500000000
0!
0*
09
0>
0C
#70510000000
1!
1*
b11 6
19
1>
1C
b11 G
#70520000000
0!
0*
09
0>
0C
#70530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#70540000000
0!
0*
09
0>
0C
#70550000000
1!
1*
b101 6
19
1>
1C
b101 G
#70560000000
0!
0*
09
0>
0C
#70570000000
1!
1*
b110 6
19
1>
1C
b110 G
#70580000000
0!
0*
09
0>
0C
#70590000000
1!
1*
b111 6
19
1>
1C
b111 G
#70600000000
0!
0*
09
0>
0C
#70610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#70620000000
0!
0*
09
0>
0C
#70630000000
1!
1*
b1 6
19
1>
1C
b1 G
#70640000000
0!
0*
09
0>
0C
#70650000000
1!
1*
b10 6
19
1>
1C
b10 G
#70660000000
0!
0*
09
0>
0C
#70670000000
1!
1*
b11 6
19
1>
1C
b11 G
#70680000000
0!
0*
09
0>
0C
#70690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#70700000000
0!
0*
09
0>
0C
#70710000000
1!
1*
b101 6
19
1>
1C
b101 G
#70720000000
0!
0*
09
0>
0C
#70730000000
1!
1*
b110 6
19
1>
1C
b110 G
#70740000000
0!
0*
09
0>
0C
#70750000000
1!
1*
b111 6
19
1>
1C
b111 G
#70760000000
0!
1"
0*
1+
09
1:
0>
0C
#70770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#70780000000
0!
0*
09
0>
0C
#70790000000
1!
1*
b1 6
19
1>
1C
b1 G
#70800000000
0!
0*
09
0>
0C
#70810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#70820000000
0!
0*
09
0>
0C
#70830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#70840000000
0!
0*
09
0>
0C
#70850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#70860000000
0!
0*
09
0>
0C
#70870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#70880000000
0!
0#
0*
0,
09
0>
0?
0C
#70890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#70900000000
0!
0*
09
0>
0C
#70910000000
1!
1*
19
1>
1C
#70920000000
0!
0*
09
0>
0C
#70930000000
1!
1*
19
1>
1C
#70940000000
0!
0*
09
0>
0C
#70950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#70960000000
0!
0*
09
0>
0C
#70970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#70980000000
0!
0*
09
0>
0C
#70990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#71000000000
0!
0*
09
0>
0C
#71010000000
1!
1*
b10 6
19
1>
1C
b10 G
#71020000000
0!
0*
09
0>
0C
#71030000000
1!
1*
b11 6
19
1>
1C
b11 G
#71040000000
0!
0*
09
0>
0C
#71050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#71060000000
0!
0*
09
0>
0C
#71070000000
1!
1*
b101 6
19
1>
1C
b101 G
#71080000000
0!
0*
09
0>
0C
#71090000000
1!
1*
b110 6
19
1>
1C
b110 G
#71100000000
0!
0*
09
0>
0C
#71110000000
1!
1*
b111 6
19
1>
1C
b111 G
#71120000000
0!
0*
09
0>
0C
#71130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#71140000000
0!
0*
09
0>
0C
#71150000000
1!
1*
b1 6
19
1>
1C
b1 G
#71160000000
0!
0*
09
0>
0C
#71170000000
1!
1*
b10 6
19
1>
1C
b10 G
#71180000000
0!
0*
09
0>
0C
#71190000000
1!
1*
b11 6
19
1>
1C
b11 G
#71200000000
0!
0*
09
0>
0C
#71210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#71220000000
0!
0*
09
0>
0C
#71230000000
1!
1*
b101 6
19
1>
1C
b101 G
#71240000000
0!
0*
09
0>
0C
#71250000000
1!
1*
b110 6
19
1>
1C
b110 G
#71260000000
0!
0*
09
0>
0C
#71270000000
1!
1*
b111 6
19
1>
1C
b111 G
#71280000000
0!
0*
09
0>
0C
#71290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#71300000000
0!
0*
09
0>
0C
#71310000000
1!
1*
b1 6
19
1>
1C
b1 G
#71320000000
0!
0*
09
0>
0C
#71330000000
1!
1*
b10 6
19
1>
1C
b10 G
#71340000000
0!
0*
09
0>
0C
#71350000000
1!
1*
b11 6
19
1>
1C
b11 G
#71360000000
0!
0*
09
0>
0C
#71370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#71380000000
0!
0*
09
0>
0C
#71390000000
1!
1*
b101 6
19
1>
1C
b101 G
#71400000000
0!
0*
09
0>
0C
#71410000000
1!
1*
b110 6
19
1>
1C
b110 G
#71420000000
0!
0*
09
0>
0C
#71430000000
1!
1*
b111 6
19
1>
1C
b111 G
#71440000000
0!
1"
0*
1+
09
1:
0>
0C
#71450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#71460000000
0!
0*
09
0>
0C
#71470000000
1!
1*
b1 6
19
1>
1C
b1 G
#71480000000
0!
0*
09
0>
0C
#71490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#71500000000
0!
0*
09
0>
0C
#71510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#71520000000
0!
0*
09
0>
0C
#71530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#71540000000
0!
0*
09
0>
0C
#71550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#71560000000
0!
0#
0*
0,
09
0>
0?
0C
#71570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#71580000000
0!
0*
09
0>
0C
#71590000000
1!
1*
19
1>
1C
#71600000000
0!
0*
09
0>
0C
#71610000000
1!
1*
19
1>
1C
#71620000000
0!
0*
09
0>
0C
#71630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#71640000000
0!
0*
09
0>
0C
#71650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#71660000000
0!
0*
09
0>
0C
#71670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#71680000000
0!
0*
09
0>
0C
#71690000000
1!
1*
b10 6
19
1>
1C
b10 G
#71700000000
0!
0*
09
0>
0C
#71710000000
1!
1*
b11 6
19
1>
1C
b11 G
#71720000000
0!
0*
09
0>
0C
#71730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#71740000000
0!
0*
09
0>
0C
#71750000000
1!
1*
b101 6
19
1>
1C
b101 G
#71760000000
0!
0*
09
0>
0C
#71770000000
1!
1*
b110 6
19
1>
1C
b110 G
#71780000000
0!
0*
09
0>
0C
#71790000000
1!
1*
b111 6
19
1>
1C
b111 G
#71800000000
0!
0*
09
0>
0C
#71810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#71820000000
0!
0*
09
0>
0C
#71830000000
1!
1*
b1 6
19
1>
1C
b1 G
#71840000000
0!
0*
09
0>
0C
#71850000000
1!
1*
b10 6
19
1>
1C
b10 G
#71860000000
0!
0*
09
0>
0C
#71870000000
1!
1*
b11 6
19
1>
1C
b11 G
#71880000000
0!
0*
09
0>
0C
#71890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#71900000000
0!
0*
09
0>
0C
#71910000000
1!
1*
b101 6
19
1>
1C
b101 G
#71920000000
0!
0*
09
0>
0C
#71930000000
1!
1*
b110 6
19
1>
1C
b110 G
#71940000000
0!
0*
09
0>
0C
#71950000000
1!
1*
b111 6
19
1>
1C
b111 G
#71960000000
0!
0*
09
0>
0C
#71970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#71980000000
0!
0*
09
0>
0C
#71990000000
1!
1*
b1 6
19
1>
1C
b1 G
#72000000000
0!
0*
09
0>
0C
#72010000000
1!
1*
b10 6
19
1>
1C
b10 G
#72020000000
0!
0*
09
0>
0C
#72030000000
1!
1*
b11 6
19
1>
1C
b11 G
#72040000000
0!
0*
09
0>
0C
#72050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#72060000000
0!
0*
09
0>
0C
#72070000000
1!
1*
b101 6
19
1>
1C
b101 G
#72080000000
0!
0*
09
0>
0C
#72090000000
1!
1*
b110 6
19
1>
1C
b110 G
#72100000000
0!
0*
09
0>
0C
#72110000000
1!
1*
b111 6
19
1>
1C
b111 G
#72120000000
0!
1"
0*
1+
09
1:
0>
0C
#72130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#72140000000
0!
0*
09
0>
0C
#72150000000
1!
1*
b1 6
19
1>
1C
b1 G
#72160000000
0!
0*
09
0>
0C
#72170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#72180000000
0!
0*
09
0>
0C
#72190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#72200000000
0!
0*
09
0>
0C
#72210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#72220000000
0!
0*
09
0>
0C
#72230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#72240000000
0!
0#
0*
0,
09
0>
0?
0C
#72250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#72260000000
0!
0*
09
0>
0C
#72270000000
1!
1*
19
1>
1C
#72280000000
0!
0*
09
0>
0C
#72290000000
1!
1*
19
1>
1C
#72300000000
0!
0*
09
0>
0C
#72310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#72320000000
0!
0*
09
0>
0C
#72330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#72340000000
0!
0*
09
0>
0C
#72350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#72360000000
0!
0*
09
0>
0C
#72370000000
1!
1*
b10 6
19
1>
1C
b10 G
#72380000000
0!
0*
09
0>
0C
#72390000000
1!
1*
b11 6
19
1>
1C
b11 G
#72400000000
0!
0*
09
0>
0C
#72410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#72420000000
0!
0*
09
0>
0C
#72430000000
1!
1*
b101 6
19
1>
1C
b101 G
#72440000000
0!
0*
09
0>
0C
#72450000000
1!
1*
b110 6
19
1>
1C
b110 G
#72460000000
0!
0*
09
0>
0C
#72470000000
1!
1*
b111 6
19
1>
1C
b111 G
#72480000000
0!
0*
09
0>
0C
#72490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#72500000000
0!
0*
09
0>
0C
#72510000000
1!
1*
b1 6
19
1>
1C
b1 G
#72520000000
0!
0*
09
0>
0C
#72530000000
1!
1*
b10 6
19
1>
1C
b10 G
#72540000000
0!
0*
09
0>
0C
#72550000000
1!
1*
b11 6
19
1>
1C
b11 G
#72560000000
0!
0*
09
0>
0C
#72570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#72580000000
0!
0*
09
0>
0C
#72590000000
1!
1*
b101 6
19
1>
1C
b101 G
#72600000000
0!
0*
09
0>
0C
#72610000000
1!
1*
b110 6
19
1>
1C
b110 G
#72620000000
0!
0*
09
0>
0C
#72630000000
1!
1*
b111 6
19
1>
1C
b111 G
#72640000000
0!
0*
09
0>
0C
#72650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#72660000000
0!
0*
09
0>
0C
#72670000000
1!
1*
b1 6
19
1>
1C
b1 G
#72680000000
0!
0*
09
0>
0C
#72690000000
1!
1*
b10 6
19
1>
1C
b10 G
#72700000000
0!
0*
09
0>
0C
#72710000000
1!
1*
b11 6
19
1>
1C
b11 G
#72720000000
0!
0*
09
0>
0C
#72730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#72740000000
0!
0*
09
0>
0C
#72750000000
1!
1*
b101 6
19
1>
1C
b101 G
#72760000000
0!
0*
09
0>
0C
#72770000000
1!
1*
b110 6
19
1>
1C
b110 G
#72780000000
0!
0*
09
0>
0C
#72790000000
1!
1*
b111 6
19
1>
1C
b111 G
#72800000000
0!
1"
0*
1+
09
1:
0>
0C
#72810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#72820000000
0!
0*
09
0>
0C
#72830000000
1!
1*
b1 6
19
1>
1C
b1 G
#72840000000
0!
0*
09
0>
0C
#72850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#72860000000
0!
0*
09
0>
0C
#72870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#72880000000
0!
0*
09
0>
0C
#72890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#72900000000
0!
0*
09
0>
0C
#72910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#72920000000
0!
0#
0*
0,
09
0>
0?
0C
#72930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#72940000000
0!
0*
09
0>
0C
#72950000000
1!
1*
19
1>
1C
#72960000000
0!
0*
09
0>
0C
#72970000000
1!
1*
19
1>
1C
#72980000000
0!
0*
09
0>
0C
#72990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#73000000000
0!
0*
09
0>
0C
#73010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#73020000000
0!
0*
09
0>
0C
#73030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#73040000000
0!
0*
09
0>
0C
#73050000000
1!
1*
b10 6
19
1>
1C
b10 G
#73060000000
0!
0*
09
0>
0C
#73070000000
1!
1*
b11 6
19
1>
1C
b11 G
#73080000000
0!
0*
09
0>
0C
#73090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#73100000000
0!
0*
09
0>
0C
#73110000000
1!
1*
b101 6
19
1>
1C
b101 G
#73120000000
0!
0*
09
0>
0C
#73130000000
1!
1*
b110 6
19
1>
1C
b110 G
#73140000000
0!
0*
09
0>
0C
#73150000000
1!
1*
b111 6
19
1>
1C
b111 G
#73160000000
0!
0*
09
0>
0C
#73170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#73180000000
0!
0*
09
0>
0C
#73190000000
1!
1*
b1 6
19
1>
1C
b1 G
#73200000000
0!
0*
09
0>
0C
#73210000000
1!
1*
b10 6
19
1>
1C
b10 G
#73220000000
0!
0*
09
0>
0C
#73230000000
1!
1*
b11 6
19
1>
1C
b11 G
#73240000000
0!
0*
09
0>
0C
#73250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#73260000000
0!
0*
09
0>
0C
#73270000000
1!
1*
b101 6
19
1>
1C
b101 G
#73280000000
0!
0*
09
0>
0C
#73290000000
1!
1*
b110 6
19
1>
1C
b110 G
#73300000000
0!
0*
09
0>
0C
#73310000000
1!
1*
b111 6
19
1>
1C
b111 G
#73320000000
0!
0*
09
0>
0C
#73330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#73340000000
0!
0*
09
0>
0C
#73350000000
1!
1*
b1 6
19
1>
1C
b1 G
#73360000000
0!
0*
09
0>
0C
#73370000000
1!
1*
b10 6
19
1>
1C
b10 G
#73380000000
0!
0*
09
0>
0C
#73390000000
1!
1*
b11 6
19
1>
1C
b11 G
#73400000000
0!
0*
09
0>
0C
#73410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#73420000000
0!
0*
09
0>
0C
#73430000000
1!
1*
b101 6
19
1>
1C
b101 G
#73440000000
0!
0*
09
0>
0C
#73450000000
1!
1*
b110 6
19
1>
1C
b110 G
#73460000000
0!
0*
09
0>
0C
#73470000000
1!
1*
b111 6
19
1>
1C
b111 G
#73480000000
0!
1"
0*
1+
09
1:
0>
0C
#73490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#73500000000
0!
0*
09
0>
0C
#73510000000
1!
1*
b1 6
19
1>
1C
b1 G
#73520000000
0!
0*
09
0>
0C
#73530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#73540000000
0!
0*
09
0>
0C
#73550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#73560000000
0!
0*
09
0>
0C
#73570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#73580000000
0!
0*
09
0>
0C
#73590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#73600000000
0!
0#
0*
0,
09
0>
0?
0C
#73610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#73620000000
0!
0*
09
0>
0C
#73630000000
1!
1*
19
1>
1C
#73640000000
0!
0*
09
0>
0C
#73650000000
1!
1*
19
1>
1C
#73660000000
0!
0*
09
0>
0C
#73670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#73680000000
0!
0*
09
0>
0C
#73690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#73700000000
0!
0*
09
0>
0C
#73710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#73720000000
0!
0*
09
0>
0C
#73730000000
1!
1*
b10 6
19
1>
1C
b10 G
#73740000000
0!
0*
09
0>
0C
#73750000000
1!
1*
b11 6
19
1>
1C
b11 G
#73760000000
0!
0*
09
0>
0C
#73770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#73780000000
0!
0*
09
0>
0C
#73790000000
1!
1*
b101 6
19
1>
1C
b101 G
#73800000000
0!
0*
09
0>
0C
#73810000000
1!
1*
b110 6
19
1>
1C
b110 G
#73820000000
0!
0*
09
0>
0C
#73830000000
1!
1*
b111 6
19
1>
1C
b111 G
#73840000000
0!
0*
09
0>
0C
#73850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#73860000000
0!
0*
09
0>
0C
#73870000000
1!
1*
b1 6
19
1>
1C
b1 G
#73880000000
0!
0*
09
0>
0C
#73890000000
1!
1*
b10 6
19
1>
1C
b10 G
#73900000000
0!
0*
09
0>
0C
#73910000000
1!
1*
b11 6
19
1>
1C
b11 G
#73920000000
0!
0*
09
0>
0C
#73930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#73940000000
0!
0*
09
0>
0C
#73950000000
1!
1*
b101 6
19
1>
1C
b101 G
#73960000000
0!
0*
09
0>
0C
#73970000000
1!
1*
b110 6
19
1>
1C
b110 G
#73980000000
0!
0*
09
0>
0C
#73990000000
1!
1*
b111 6
19
1>
1C
b111 G
#74000000000
0!
0*
09
0>
0C
#74010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#74020000000
0!
0*
09
0>
0C
#74030000000
1!
1*
b1 6
19
1>
1C
b1 G
#74040000000
0!
0*
09
0>
0C
#74050000000
1!
1*
b10 6
19
1>
1C
b10 G
#74060000000
0!
0*
09
0>
0C
#74070000000
1!
1*
b11 6
19
1>
1C
b11 G
#74080000000
0!
0*
09
0>
0C
#74090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#74100000000
0!
0*
09
0>
0C
#74110000000
1!
1*
b101 6
19
1>
1C
b101 G
#74120000000
0!
0*
09
0>
0C
#74130000000
1!
1*
b110 6
19
1>
1C
b110 G
#74140000000
0!
0*
09
0>
0C
#74150000000
1!
1*
b111 6
19
1>
1C
b111 G
#74160000000
0!
1"
0*
1+
09
1:
0>
0C
#74170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#74180000000
0!
0*
09
0>
0C
#74190000000
1!
1*
b1 6
19
1>
1C
b1 G
#74200000000
0!
0*
09
0>
0C
#74210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#74220000000
0!
0*
09
0>
0C
#74230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#74240000000
0!
0*
09
0>
0C
#74250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#74260000000
0!
0*
09
0>
0C
#74270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#74280000000
0!
0#
0*
0,
09
0>
0?
0C
#74290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#74300000000
0!
0*
09
0>
0C
#74310000000
1!
1*
19
1>
1C
#74320000000
0!
0*
09
0>
0C
#74330000000
1!
1*
19
1>
1C
#74340000000
0!
0*
09
0>
0C
#74350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#74360000000
0!
0*
09
0>
0C
#74370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#74380000000
0!
0*
09
0>
0C
#74390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#74400000000
0!
0*
09
0>
0C
#74410000000
1!
1*
b10 6
19
1>
1C
b10 G
#74420000000
0!
0*
09
0>
0C
#74430000000
1!
1*
b11 6
19
1>
1C
b11 G
#74440000000
0!
0*
09
0>
0C
#74450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#74460000000
0!
0*
09
0>
0C
#74470000000
1!
1*
b101 6
19
1>
1C
b101 G
#74480000000
0!
0*
09
0>
0C
#74490000000
1!
1*
b110 6
19
1>
1C
b110 G
#74500000000
0!
0*
09
0>
0C
#74510000000
1!
1*
b111 6
19
1>
1C
b111 G
#74520000000
0!
0*
09
0>
0C
#74530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#74540000000
0!
0*
09
0>
0C
#74550000000
1!
1*
b1 6
19
1>
1C
b1 G
#74560000000
0!
0*
09
0>
0C
#74570000000
1!
1*
b10 6
19
1>
1C
b10 G
#74580000000
0!
0*
09
0>
0C
#74590000000
1!
1*
b11 6
19
1>
1C
b11 G
#74600000000
0!
0*
09
0>
0C
#74610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#74620000000
0!
0*
09
0>
0C
#74630000000
1!
1*
b101 6
19
1>
1C
b101 G
#74640000000
0!
0*
09
0>
0C
#74650000000
1!
1*
b110 6
19
1>
1C
b110 G
#74660000000
0!
0*
09
0>
0C
#74670000000
1!
1*
b111 6
19
1>
1C
b111 G
#74680000000
0!
0*
09
0>
0C
#74690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#74700000000
0!
0*
09
0>
0C
#74710000000
1!
1*
b1 6
19
1>
1C
b1 G
#74720000000
0!
0*
09
0>
0C
#74730000000
1!
1*
b10 6
19
1>
1C
b10 G
#74740000000
0!
0*
09
0>
0C
#74750000000
1!
1*
b11 6
19
1>
1C
b11 G
#74760000000
0!
0*
09
0>
0C
#74770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#74780000000
0!
0*
09
0>
0C
#74790000000
1!
1*
b101 6
19
1>
1C
b101 G
#74800000000
0!
0*
09
0>
0C
#74810000000
1!
1*
b110 6
19
1>
1C
b110 G
#74820000000
0!
0*
09
0>
0C
#74830000000
1!
1*
b111 6
19
1>
1C
b111 G
#74840000000
0!
1"
0*
1+
09
1:
0>
0C
#74850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#74860000000
0!
0*
09
0>
0C
#74870000000
1!
1*
b1 6
19
1>
1C
b1 G
#74880000000
0!
0*
09
0>
0C
#74890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#74900000000
0!
0*
09
0>
0C
#74910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#74920000000
0!
0*
09
0>
0C
#74930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#74940000000
0!
0*
09
0>
0C
#74950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#74960000000
0!
0#
0*
0,
09
0>
0?
0C
#74970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#74980000000
0!
0*
09
0>
0C
#74990000000
1!
1*
19
1>
1C
#75000000000
0!
0*
09
0>
0C
#75010000000
1!
1*
19
1>
1C
#75020000000
0!
0*
09
0>
0C
#75030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#75040000000
0!
0*
09
0>
0C
#75050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#75060000000
0!
0*
09
0>
0C
#75070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#75080000000
0!
0*
09
0>
0C
#75090000000
1!
1*
b10 6
19
1>
1C
b10 G
#75100000000
0!
0*
09
0>
0C
#75110000000
1!
1*
b11 6
19
1>
1C
b11 G
#75120000000
0!
0*
09
0>
0C
#75130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#75140000000
0!
0*
09
0>
0C
#75150000000
1!
1*
b101 6
19
1>
1C
b101 G
#75160000000
0!
0*
09
0>
0C
#75170000000
1!
1*
b110 6
19
1>
1C
b110 G
#75180000000
0!
0*
09
0>
0C
#75190000000
1!
1*
b111 6
19
1>
1C
b111 G
#75200000000
0!
0*
09
0>
0C
#75210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#75220000000
0!
0*
09
0>
0C
#75230000000
1!
1*
b1 6
19
1>
1C
b1 G
#75240000000
0!
0*
09
0>
0C
#75250000000
1!
1*
b10 6
19
1>
1C
b10 G
#75260000000
0!
0*
09
0>
0C
#75270000000
1!
1*
b11 6
19
1>
1C
b11 G
#75280000000
0!
0*
09
0>
0C
#75290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#75300000000
0!
0*
09
0>
0C
#75310000000
1!
1*
b101 6
19
1>
1C
b101 G
#75320000000
0!
0*
09
0>
0C
#75330000000
1!
1*
b110 6
19
1>
1C
b110 G
#75340000000
0!
0*
09
0>
0C
#75350000000
1!
1*
b111 6
19
1>
1C
b111 G
#75360000000
0!
0*
09
0>
0C
#75370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#75380000000
0!
0*
09
0>
0C
#75390000000
1!
1*
b1 6
19
1>
1C
b1 G
#75400000000
0!
0*
09
0>
0C
#75410000000
1!
1*
b10 6
19
1>
1C
b10 G
#75420000000
0!
0*
09
0>
0C
#75430000000
1!
1*
b11 6
19
1>
1C
b11 G
#75440000000
0!
0*
09
0>
0C
#75450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#75460000000
0!
0*
09
0>
0C
#75470000000
1!
1*
b101 6
19
1>
1C
b101 G
#75480000000
0!
0*
09
0>
0C
#75490000000
1!
1*
b110 6
19
1>
1C
b110 G
#75500000000
0!
0*
09
0>
0C
#75510000000
1!
1*
b111 6
19
1>
1C
b111 G
#75520000000
0!
1"
0*
1+
09
1:
0>
0C
#75530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#75540000000
0!
0*
09
0>
0C
#75550000000
1!
1*
b1 6
19
1>
1C
b1 G
#75560000000
0!
0*
09
0>
0C
#75570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#75580000000
0!
0*
09
0>
0C
#75590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#75600000000
0!
0*
09
0>
0C
#75610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#75620000000
0!
0*
09
0>
0C
#75630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#75640000000
0!
0#
0*
0,
09
0>
0?
0C
#75650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#75660000000
0!
0*
09
0>
0C
#75670000000
1!
1*
19
1>
1C
#75680000000
0!
0*
09
0>
0C
#75690000000
1!
1*
19
1>
1C
#75700000000
0!
0*
09
0>
0C
#75710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#75720000000
0!
0*
09
0>
0C
#75730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#75740000000
0!
0*
09
0>
0C
#75750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#75760000000
0!
0*
09
0>
0C
#75770000000
1!
1*
b10 6
19
1>
1C
b10 G
#75780000000
0!
0*
09
0>
0C
#75790000000
1!
1*
b11 6
19
1>
1C
b11 G
#75800000000
0!
0*
09
0>
0C
#75810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#75820000000
0!
0*
09
0>
0C
#75830000000
1!
1*
b101 6
19
1>
1C
b101 G
#75840000000
0!
0*
09
0>
0C
#75850000000
1!
1*
b110 6
19
1>
1C
b110 G
#75860000000
0!
0*
09
0>
0C
#75870000000
1!
1*
b111 6
19
1>
1C
b111 G
#75880000000
0!
0*
09
0>
0C
#75890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#75900000000
0!
0*
09
0>
0C
#75910000000
1!
1*
b1 6
19
1>
1C
b1 G
#75920000000
0!
0*
09
0>
0C
#75930000000
1!
1*
b10 6
19
1>
1C
b10 G
#75940000000
0!
0*
09
0>
0C
#75950000000
1!
1*
b11 6
19
1>
1C
b11 G
#75960000000
0!
0*
09
0>
0C
#75970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#75980000000
0!
0*
09
0>
0C
#75990000000
1!
1*
b101 6
19
1>
1C
b101 G
#76000000000
0!
0*
09
0>
0C
#76010000000
1!
1*
b110 6
19
1>
1C
b110 G
#76020000000
0!
0*
09
0>
0C
#76030000000
1!
1*
b111 6
19
1>
1C
b111 G
#76040000000
0!
0*
09
0>
0C
#76050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#76060000000
0!
0*
09
0>
0C
#76070000000
1!
1*
b1 6
19
1>
1C
b1 G
#76080000000
0!
0*
09
0>
0C
#76090000000
1!
1*
b10 6
19
1>
1C
b10 G
#76100000000
0!
0*
09
0>
0C
#76110000000
1!
1*
b11 6
19
1>
1C
b11 G
#76120000000
0!
0*
09
0>
0C
#76130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#76140000000
0!
0*
09
0>
0C
#76150000000
1!
1*
b101 6
19
1>
1C
b101 G
#76160000000
0!
0*
09
0>
0C
#76170000000
1!
1*
b110 6
19
1>
1C
b110 G
#76180000000
0!
0*
09
0>
0C
#76190000000
1!
1*
b111 6
19
1>
1C
b111 G
#76200000000
0!
1"
0*
1+
09
1:
0>
0C
#76210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#76220000000
0!
0*
09
0>
0C
#76230000000
1!
1*
b1 6
19
1>
1C
b1 G
#76240000000
0!
0*
09
0>
0C
#76250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#76260000000
0!
0*
09
0>
0C
#76270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#76280000000
0!
0*
09
0>
0C
#76290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#76300000000
0!
0*
09
0>
0C
#76310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#76320000000
0!
0#
0*
0,
09
0>
0?
0C
#76330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#76340000000
0!
0*
09
0>
0C
#76350000000
1!
1*
19
1>
1C
#76360000000
0!
0*
09
0>
0C
#76370000000
1!
1*
19
1>
1C
#76380000000
0!
0*
09
0>
0C
#76390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#76400000000
0!
0*
09
0>
0C
#76410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#76420000000
0!
0*
09
0>
0C
#76430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#76440000000
0!
0*
09
0>
0C
#76450000000
1!
1*
b10 6
19
1>
1C
b10 G
#76460000000
0!
0*
09
0>
0C
#76470000000
1!
1*
b11 6
19
1>
1C
b11 G
#76480000000
0!
0*
09
0>
0C
#76490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#76500000000
0!
0*
09
0>
0C
#76510000000
1!
1*
b101 6
19
1>
1C
b101 G
#76520000000
0!
0*
09
0>
0C
#76530000000
1!
1*
b110 6
19
1>
1C
b110 G
#76540000000
0!
0*
09
0>
0C
#76550000000
1!
1*
b111 6
19
1>
1C
b111 G
#76560000000
0!
0*
09
0>
0C
#76570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#76580000000
0!
0*
09
0>
0C
#76590000000
1!
1*
b1 6
19
1>
1C
b1 G
#76600000000
0!
0*
09
0>
0C
#76610000000
1!
1*
b10 6
19
1>
1C
b10 G
#76620000000
0!
0*
09
0>
0C
#76630000000
1!
1*
b11 6
19
1>
1C
b11 G
#76640000000
0!
0*
09
0>
0C
#76650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#76660000000
0!
0*
09
0>
0C
#76670000000
1!
1*
b101 6
19
1>
1C
b101 G
#76680000000
0!
0*
09
0>
0C
#76690000000
1!
1*
b110 6
19
1>
1C
b110 G
#76700000000
0!
0*
09
0>
0C
#76710000000
1!
1*
b111 6
19
1>
1C
b111 G
#76720000000
0!
0*
09
0>
0C
#76730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#76740000000
0!
0*
09
0>
0C
#76750000000
1!
1*
b1 6
19
1>
1C
b1 G
#76760000000
0!
0*
09
0>
0C
#76770000000
1!
1*
b10 6
19
1>
1C
b10 G
#76780000000
0!
0*
09
0>
0C
#76790000000
1!
1*
b11 6
19
1>
1C
b11 G
#76800000000
0!
0*
09
0>
0C
#76810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#76820000000
0!
0*
09
0>
0C
#76830000000
1!
1*
b101 6
19
1>
1C
b101 G
#76840000000
0!
0*
09
0>
0C
#76850000000
1!
1*
b110 6
19
1>
1C
b110 G
#76860000000
0!
0*
09
0>
0C
#76870000000
1!
1*
b111 6
19
1>
1C
b111 G
#76880000000
0!
1"
0*
1+
09
1:
0>
0C
#76890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#76900000000
0!
0*
09
0>
0C
#76910000000
1!
1*
b1 6
19
1>
1C
b1 G
#76920000000
0!
0*
09
0>
0C
#76930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#76940000000
0!
0*
09
0>
0C
#76950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#76960000000
0!
0*
09
0>
0C
#76970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#76980000000
0!
0*
09
0>
0C
#76990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#77000000000
0!
0#
0*
0,
09
0>
0?
0C
#77010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#77020000000
0!
0*
09
0>
0C
#77030000000
1!
1*
19
1>
1C
#77040000000
0!
0*
09
0>
0C
#77050000000
1!
1*
19
1>
1C
#77060000000
0!
0*
09
0>
0C
#77070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#77080000000
0!
0*
09
0>
0C
#77090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#77100000000
0!
0*
09
0>
0C
#77110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#77120000000
0!
0*
09
0>
0C
#77130000000
1!
1*
b10 6
19
1>
1C
b10 G
#77140000000
0!
0*
09
0>
0C
#77150000000
1!
1*
b11 6
19
1>
1C
b11 G
#77160000000
0!
0*
09
0>
0C
#77170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#77180000000
0!
0*
09
0>
0C
#77190000000
1!
1*
b101 6
19
1>
1C
b101 G
#77200000000
0!
0*
09
0>
0C
#77210000000
1!
1*
b110 6
19
1>
1C
b110 G
#77220000000
0!
0*
09
0>
0C
#77230000000
1!
1*
b111 6
19
1>
1C
b111 G
#77240000000
0!
0*
09
0>
0C
#77250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#77260000000
0!
0*
09
0>
0C
#77270000000
1!
1*
b1 6
19
1>
1C
b1 G
#77280000000
0!
0*
09
0>
0C
#77290000000
1!
1*
b10 6
19
1>
1C
b10 G
#77300000000
0!
0*
09
0>
0C
#77310000000
1!
1*
b11 6
19
1>
1C
b11 G
#77320000000
0!
0*
09
0>
0C
#77330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#77340000000
0!
0*
09
0>
0C
#77350000000
1!
1*
b101 6
19
1>
1C
b101 G
#77360000000
0!
0*
09
0>
0C
#77370000000
1!
1*
b110 6
19
1>
1C
b110 G
#77380000000
0!
0*
09
0>
0C
#77390000000
1!
1*
b111 6
19
1>
1C
b111 G
#77400000000
0!
0*
09
0>
0C
#77410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#77420000000
0!
0*
09
0>
0C
#77430000000
1!
1*
b1 6
19
1>
1C
b1 G
#77440000000
0!
0*
09
0>
0C
#77450000000
1!
1*
b10 6
19
1>
1C
b10 G
#77460000000
0!
0*
09
0>
0C
#77470000000
1!
1*
b11 6
19
1>
1C
b11 G
#77480000000
0!
0*
09
0>
0C
#77490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#77500000000
0!
0*
09
0>
0C
#77510000000
1!
1*
b101 6
19
1>
1C
b101 G
#77520000000
0!
0*
09
0>
0C
#77530000000
1!
1*
b110 6
19
1>
1C
b110 G
#77540000000
0!
0*
09
0>
0C
#77550000000
1!
1*
b111 6
19
1>
1C
b111 G
#77560000000
0!
1"
0*
1+
09
1:
0>
0C
#77570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#77580000000
0!
0*
09
0>
0C
#77590000000
1!
1*
b1 6
19
1>
1C
b1 G
#77600000000
0!
0*
09
0>
0C
#77610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#77620000000
0!
0*
09
0>
0C
#77630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#77640000000
0!
0*
09
0>
0C
#77650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#77660000000
0!
0*
09
0>
0C
#77670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#77680000000
0!
0#
0*
0,
09
0>
0?
0C
#77690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#77700000000
0!
0*
09
0>
0C
#77710000000
1!
1*
19
1>
1C
#77720000000
0!
0*
09
0>
0C
#77730000000
1!
1*
19
1>
1C
#77740000000
0!
0*
09
0>
0C
#77750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#77760000000
0!
0*
09
0>
0C
#77770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#77780000000
0!
0*
09
0>
0C
#77790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#77800000000
0!
0*
09
0>
0C
#77810000000
1!
1*
b10 6
19
1>
1C
b10 G
#77820000000
0!
0*
09
0>
0C
#77830000000
1!
1*
b11 6
19
1>
1C
b11 G
#77840000000
0!
0*
09
0>
0C
#77850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#77860000000
0!
0*
09
0>
0C
#77870000000
1!
1*
b101 6
19
1>
1C
b101 G
#77880000000
0!
0*
09
0>
0C
#77890000000
1!
1*
b110 6
19
1>
1C
b110 G
#77900000000
0!
0*
09
0>
0C
#77910000000
1!
1*
b111 6
19
1>
1C
b111 G
#77920000000
0!
0*
09
0>
0C
#77930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#77940000000
0!
0*
09
0>
0C
#77950000000
1!
1*
b1 6
19
1>
1C
b1 G
#77960000000
0!
0*
09
0>
0C
#77970000000
1!
1*
b10 6
19
1>
1C
b10 G
#77980000000
0!
0*
09
0>
0C
#77990000000
1!
1*
b11 6
19
1>
1C
b11 G
#78000000000
0!
0*
09
0>
0C
#78010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#78020000000
0!
0*
09
0>
0C
#78030000000
1!
1*
b101 6
19
1>
1C
b101 G
#78040000000
0!
0*
09
0>
0C
#78050000000
1!
1*
b110 6
19
1>
1C
b110 G
#78060000000
0!
0*
09
0>
0C
#78070000000
1!
1*
b111 6
19
1>
1C
b111 G
#78080000000
0!
0*
09
0>
0C
#78090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#78100000000
0!
0*
09
0>
0C
#78110000000
1!
1*
b1 6
19
1>
1C
b1 G
#78120000000
0!
0*
09
0>
0C
#78130000000
1!
1*
b10 6
19
1>
1C
b10 G
#78140000000
0!
0*
09
0>
0C
#78150000000
1!
1*
b11 6
19
1>
1C
b11 G
#78160000000
0!
0*
09
0>
0C
#78170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#78180000000
0!
0*
09
0>
0C
#78190000000
1!
1*
b101 6
19
1>
1C
b101 G
#78200000000
0!
0*
09
0>
0C
#78210000000
1!
1*
b110 6
19
1>
1C
b110 G
#78220000000
0!
0*
09
0>
0C
#78230000000
1!
1*
b111 6
19
1>
1C
b111 G
#78240000000
0!
1"
0*
1+
09
1:
0>
0C
#78250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#78260000000
0!
0*
09
0>
0C
#78270000000
1!
1*
b1 6
19
1>
1C
b1 G
#78280000000
0!
0*
09
0>
0C
#78290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#78300000000
0!
0*
09
0>
0C
#78310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#78320000000
0!
0*
09
0>
0C
#78330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#78340000000
0!
0*
09
0>
0C
#78350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#78360000000
0!
0#
0*
0,
09
0>
0?
0C
#78370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#78380000000
0!
0*
09
0>
0C
#78390000000
1!
1*
19
1>
1C
#78400000000
0!
0*
09
0>
0C
#78410000000
1!
1*
19
1>
1C
#78420000000
0!
0*
09
0>
0C
#78430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#78440000000
0!
0*
09
0>
0C
#78450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#78460000000
0!
0*
09
0>
0C
#78470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#78480000000
0!
0*
09
0>
0C
#78490000000
1!
1*
b10 6
19
1>
1C
b10 G
#78500000000
0!
0*
09
0>
0C
#78510000000
1!
1*
b11 6
19
1>
1C
b11 G
#78520000000
0!
0*
09
0>
0C
#78530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#78540000000
0!
0*
09
0>
0C
#78550000000
1!
1*
b101 6
19
1>
1C
b101 G
#78560000000
0!
0*
09
0>
0C
#78570000000
1!
1*
b110 6
19
1>
1C
b110 G
#78580000000
0!
0*
09
0>
0C
#78590000000
1!
1*
b111 6
19
1>
1C
b111 G
#78600000000
0!
0*
09
0>
0C
#78610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#78620000000
0!
0*
09
0>
0C
#78630000000
1!
1*
b1 6
19
1>
1C
b1 G
#78640000000
0!
0*
09
0>
0C
#78650000000
1!
1*
b10 6
19
1>
1C
b10 G
#78660000000
0!
0*
09
0>
0C
#78670000000
1!
1*
b11 6
19
1>
1C
b11 G
#78680000000
0!
0*
09
0>
0C
#78690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#78700000000
0!
0*
09
0>
0C
#78710000000
1!
1*
b101 6
19
1>
1C
b101 G
#78720000000
0!
0*
09
0>
0C
#78730000000
1!
1*
b110 6
19
1>
1C
b110 G
#78740000000
0!
0*
09
0>
0C
#78750000000
1!
1*
b111 6
19
1>
1C
b111 G
#78760000000
0!
0*
09
0>
0C
#78770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#78780000000
0!
0*
09
0>
0C
#78790000000
1!
1*
b1 6
19
1>
1C
b1 G
#78800000000
0!
0*
09
0>
0C
#78810000000
1!
1*
b10 6
19
1>
1C
b10 G
#78820000000
0!
0*
09
0>
0C
#78830000000
1!
1*
b11 6
19
1>
1C
b11 G
#78840000000
0!
0*
09
0>
0C
#78850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#78860000000
0!
0*
09
0>
0C
#78870000000
1!
1*
b101 6
19
1>
1C
b101 G
#78880000000
0!
0*
09
0>
0C
#78890000000
1!
1*
b110 6
19
1>
1C
b110 G
#78900000000
0!
0*
09
0>
0C
#78910000000
1!
1*
b111 6
19
1>
1C
b111 G
#78920000000
0!
1"
0*
1+
09
1:
0>
0C
#78930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#78940000000
0!
0*
09
0>
0C
#78950000000
1!
1*
b1 6
19
1>
1C
b1 G
#78960000000
0!
0*
09
0>
0C
#78970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#78980000000
0!
0*
09
0>
0C
#78990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#79000000000
0!
0*
09
0>
0C
#79010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#79020000000
0!
0*
09
0>
0C
#79030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#79040000000
0!
0#
0*
0,
09
0>
0?
0C
#79050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#79060000000
0!
0*
09
0>
0C
#79070000000
1!
1*
19
1>
1C
#79080000000
0!
0*
09
0>
0C
#79090000000
1!
1*
19
1>
1C
#79100000000
0!
0*
09
0>
0C
#79110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#79120000000
0!
0*
09
0>
0C
#79130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#79140000000
0!
0*
09
0>
0C
#79150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#79160000000
0!
0*
09
0>
0C
#79170000000
1!
1*
b10 6
19
1>
1C
b10 G
#79180000000
0!
0*
09
0>
0C
#79190000000
1!
1*
b11 6
19
1>
1C
b11 G
#79200000000
0!
0*
09
0>
0C
#79210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#79220000000
0!
0*
09
0>
0C
#79230000000
1!
1*
b101 6
19
1>
1C
b101 G
#79240000000
0!
0*
09
0>
0C
#79250000000
1!
1*
b110 6
19
1>
1C
b110 G
#79260000000
0!
0*
09
0>
0C
#79270000000
1!
1*
b111 6
19
1>
1C
b111 G
#79280000000
0!
0*
09
0>
0C
#79290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#79300000000
0!
0*
09
0>
0C
#79310000000
1!
1*
b1 6
19
1>
1C
b1 G
#79320000000
0!
0*
09
0>
0C
#79330000000
1!
1*
b10 6
19
1>
1C
b10 G
#79340000000
0!
0*
09
0>
0C
#79350000000
1!
1*
b11 6
19
1>
1C
b11 G
#79360000000
0!
0*
09
0>
0C
#79370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#79380000000
0!
0*
09
0>
0C
#79390000000
1!
1*
b101 6
19
1>
1C
b101 G
#79400000000
0!
0*
09
0>
0C
#79410000000
1!
1*
b110 6
19
1>
1C
b110 G
#79420000000
0!
0*
09
0>
0C
#79430000000
1!
1*
b111 6
19
1>
1C
b111 G
#79440000000
0!
0*
09
0>
0C
#79450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#79460000000
0!
0*
09
0>
0C
#79470000000
1!
1*
b1 6
19
1>
1C
b1 G
#79480000000
0!
0*
09
0>
0C
#79490000000
1!
1*
b10 6
19
1>
1C
b10 G
#79500000000
0!
0*
09
0>
0C
#79510000000
1!
1*
b11 6
19
1>
1C
b11 G
#79520000000
0!
0*
09
0>
0C
#79530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#79540000000
0!
0*
09
0>
0C
#79550000000
1!
1*
b101 6
19
1>
1C
b101 G
#79560000000
0!
0*
09
0>
0C
#79570000000
1!
1*
b110 6
19
1>
1C
b110 G
#79580000000
0!
0*
09
0>
0C
#79590000000
1!
1*
b111 6
19
1>
1C
b111 G
#79600000000
0!
1"
0*
1+
09
1:
0>
0C
#79610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#79620000000
0!
0*
09
0>
0C
#79630000000
1!
1*
b1 6
19
1>
1C
b1 G
#79640000000
0!
0*
09
0>
0C
#79650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#79660000000
0!
0*
09
0>
0C
#79670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#79680000000
0!
0*
09
0>
0C
#79690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#79700000000
0!
0*
09
0>
0C
#79710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#79720000000
0!
0#
0*
0,
09
0>
0?
0C
#79730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#79740000000
0!
0*
09
0>
0C
#79750000000
1!
1*
19
1>
1C
#79760000000
0!
0*
09
0>
0C
#79770000000
1!
1*
19
1>
1C
#79780000000
0!
0*
09
0>
0C
#79790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#79800000000
0!
0*
09
0>
0C
#79810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#79820000000
0!
0*
09
0>
0C
#79830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#79840000000
0!
0*
09
0>
0C
#79850000000
1!
1*
b10 6
19
1>
1C
b10 G
#79860000000
0!
0*
09
0>
0C
#79870000000
1!
1*
b11 6
19
1>
1C
b11 G
#79880000000
0!
0*
09
0>
0C
#79890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#79900000000
0!
0*
09
0>
0C
#79910000000
1!
1*
b101 6
19
1>
1C
b101 G
#79920000000
0!
0*
09
0>
0C
#79930000000
1!
1*
b110 6
19
1>
1C
b110 G
#79940000000
0!
0*
09
0>
0C
#79950000000
1!
1*
b111 6
19
1>
1C
b111 G
#79960000000
0!
0*
09
0>
0C
#79970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#79980000000
0!
0*
09
0>
0C
#79990000000
1!
1*
b1 6
19
1>
1C
b1 G
#80000000000
0!
0*
09
0>
0C
#80010000000
1!
1*
b10 6
19
1>
1C
b10 G
#80020000000
0!
0*
09
0>
0C
#80030000000
1!
1*
b11 6
19
1>
1C
b11 G
#80040000000
0!
0*
09
0>
0C
#80050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#80060000000
0!
0*
09
0>
0C
#80070000000
1!
1*
b101 6
19
1>
1C
b101 G
#80080000000
0!
0*
09
0>
0C
#80090000000
1!
1*
b110 6
19
1>
1C
b110 G
#80100000000
0!
0*
09
0>
0C
#80110000000
1!
1*
b111 6
19
1>
1C
b111 G
#80120000000
0!
0*
09
0>
0C
#80130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#80140000000
0!
0*
09
0>
0C
#80150000000
1!
1*
b1 6
19
1>
1C
b1 G
#80160000000
0!
0*
09
0>
0C
#80170000000
1!
1*
b10 6
19
1>
1C
b10 G
#80180000000
0!
0*
09
0>
0C
#80190000000
1!
1*
b11 6
19
1>
1C
b11 G
#80200000000
0!
0*
09
0>
0C
#80210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#80220000000
0!
0*
09
0>
0C
#80230000000
1!
1*
b101 6
19
1>
1C
b101 G
#80240000000
0!
0*
09
0>
0C
#80250000000
1!
1*
b110 6
19
1>
1C
b110 G
#80260000000
0!
0*
09
0>
0C
#80270000000
1!
1*
b111 6
19
1>
1C
b111 G
#80280000000
0!
1"
0*
1+
09
1:
0>
0C
#80290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#80300000000
0!
0*
09
0>
0C
#80310000000
1!
1*
b1 6
19
1>
1C
b1 G
#80320000000
0!
0*
09
0>
0C
#80330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#80340000000
0!
0*
09
0>
0C
#80350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#80360000000
0!
0*
09
0>
0C
#80370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#80380000000
0!
0*
09
0>
0C
#80390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#80400000000
0!
0#
0*
0,
09
0>
0?
0C
#80410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#80420000000
0!
0*
09
0>
0C
#80430000000
1!
1*
19
1>
1C
#80440000000
0!
0*
09
0>
0C
#80450000000
1!
1*
19
1>
1C
#80460000000
0!
0*
09
0>
0C
#80470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#80480000000
0!
0*
09
0>
0C
#80490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#80500000000
0!
0*
09
0>
0C
#80510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#80520000000
0!
0*
09
0>
0C
#80530000000
1!
1*
b10 6
19
1>
1C
b10 G
#80540000000
0!
0*
09
0>
0C
#80550000000
1!
1*
b11 6
19
1>
1C
b11 G
#80560000000
0!
0*
09
0>
0C
#80570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#80580000000
0!
0*
09
0>
0C
#80590000000
1!
1*
b101 6
19
1>
1C
b101 G
#80600000000
0!
0*
09
0>
0C
#80610000000
1!
1*
b110 6
19
1>
1C
b110 G
#80620000000
0!
0*
09
0>
0C
#80630000000
1!
1*
b111 6
19
1>
1C
b111 G
#80640000000
0!
0*
09
0>
0C
#80650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#80660000000
0!
0*
09
0>
0C
#80670000000
1!
1*
b1 6
19
1>
1C
b1 G
#80680000000
0!
0*
09
0>
0C
#80690000000
1!
1*
b10 6
19
1>
1C
b10 G
#80700000000
0!
0*
09
0>
0C
#80710000000
1!
1*
b11 6
19
1>
1C
b11 G
#80720000000
0!
0*
09
0>
0C
#80730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#80740000000
0!
0*
09
0>
0C
#80750000000
1!
1*
b101 6
19
1>
1C
b101 G
#80760000000
0!
0*
09
0>
0C
#80770000000
1!
1*
b110 6
19
1>
1C
b110 G
#80780000000
0!
0*
09
0>
0C
#80790000000
1!
1*
b111 6
19
1>
1C
b111 G
#80800000000
0!
0*
09
0>
0C
#80810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#80820000000
0!
0*
09
0>
0C
#80830000000
1!
1*
b1 6
19
1>
1C
b1 G
#80840000000
0!
0*
09
0>
0C
#80850000000
1!
1*
b10 6
19
1>
1C
b10 G
#80860000000
0!
0*
09
0>
0C
#80870000000
1!
1*
b11 6
19
1>
1C
b11 G
#80880000000
0!
0*
09
0>
0C
#80890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#80900000000
0!
0*
09
0>
0C
#80910000000
1!
1*
b101 6
19
1>
1C
b101 G
#80920000000
0!
0*
09
0>
0C
#80930000000
1!
1*
b110 6
19
1>
1C
b110 G
#80940000000
0!
0*
09
0>
0C
#80950000000
1!
1*
b111 6
19
1>
1C
b111 G
#80960000000
0!
1"
0*
1+
09
1:
0>
0C
#80970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#80980000000
0!
0*
09
0>
0C
#80990000000
1!
1*
b1 6
19
1>
1C
b1 G
#81000000000
0!
0*
09
0>
0C
#81010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#81020000000
0!
0*
09
0>
0C
#81030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#81040000000
0!
0*
09
0>
0C
#81050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#81060000000
0!
0*
09
0>
0C
#81070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#81080000000
0!
0#
0*
0,
09
0>
0?
0C
#81090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#81100000000
0!
0*
09
0>
0C
#81110000000
1!
1*
19
1>
1C
#81120000000
0!
0*
09
0>
0C
#81130000000
1!
1*
19
1>
1C
#81140000000
0!
0*
09
0>
0C
#81150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#81160000000
0!
0*
09
0>
0C
#81170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#81180000000
0!
0*
09
0>
0C
#81190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#81200000000
0!
0*
09
0>
0C
#81210000000
1!
1*
b10 6
19
1>
1C
b10 G
#81220000000
0!
0*
09
0>
0C
#81230000000
1!
1*
b11 6
19
1>
1C
b11 G
#81240000000
0!
0*
09
0>
0C
#81250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#81260000000
0!
0*
09
0>
0C
#81270000000
1!
1*
b101 6
19
1>
1C
b101 G
#81280000000
0!
0*
09
0>
0C
#81290000000
1!
1*
b110 6
19
1>
1C
b110 G
#81300000000
0!
0*
09
0>
0C
#81310000000
1!
1*
b111 6
19
1>
1C
b111 G
#81320000000
0!
0*
09
0>
0C
#81330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#81340000000
0!
0*
09
0>
0C
#81350000000
1!
1*
b1 6
19
1>
1C
b1 G
#81360000000
0!
0*
09
0>
0C
#81370000000
1!
1*
b10 6
19
1>
1C
b10 G
#81380000000
0!
0*
09
0>
0C
#81390000000
1!
1*
b11 6
19
1>
1C
b11 G
#81400000000
0!
0*
09
0>
0C
#81410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#81420000000
0!
0*
09
0>
0C
#81430000000
1!
1*
b101 6
19
1>
1C
b101 G
#81440000000
0!
0*
09
0>
0C
#81450000000
1!
1*
b110 6
19
1>
1C
b110 G
#81460000000
0!
0*
09
0>
0C
#81470000000
1!
1*
b111 6
19
1>
1C
b111 G
#81480000000
0!
0*
09
0>
0C
#81490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#81500000000
0!
0*
09
0>
0C
#81510000000
1!
1*
b1 6
19
1>
1C
b1 G
#81520000000
0!
0*
09
0>
0C
#81530000000
1!
1*
b10 6
19
1>
1C
b10 G
#81540000000
0!
0*
09
0>
0C
#81550000000
1!
1*
b11 6
19
1>
1C
b11 G
#81560000000
0!
0*
09
0>
0C
#81570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#81580000000
0!
0*
09
0>
0C
#81590000000
1!
1*
b101 6
19
1>
1C
b101 G
#81600000000
0!
0*
09
0>
0C
#81610000000
1!
1*
b110 6
19
1>
1C
b110 G
#81620000000
0!
0*
09
0>
0C
#81630000000
1!
1*
b111 6
19
1>
1C
b111 G
#81640000000
0!
1"
0*
1+
09
1:
0>
0C
#81650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#81660000000
0!
0*
09
0>
0C
#81670000000
1!
1*
b1 6
19
1>
1C
b1 G
#81680000000
0!
0*
09
0>
0C
#81690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#81700000000
0!
0*
09
0>
0C
#81710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#81720000000
0!
0*
09
0>
0C
#81730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#81740000000
0!
0*
09
0>
0C
#81750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#81760000000
0!
0#
0*
0,
09
0>
0?
0C
#81770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#81780000000
0!
0*
09
0>
0C
#81790000000
1!
1*
19
1>
1C
#81800000000
0!
0*
09
0>
0C
#81810000000
1!
1*
19
1>
1C
#81820000000
0!
0*
09
0>
0C
#81830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#81840000000
0!
0*
09
0>
0C
#81850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#81860000000
0!
0*
09
0>
0C
#81870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#81880000000
0!
0*
09
0>
0C
#81890000000
1!
1*
b10 6
19
1>
1C
b10 G
#81900000000
0!
0*
09
0>
0C
#81910000000
1!
1*
b11 6
19
1>
1C
b11 G
#81920000000
0!
0*
09
0>
0C
#81930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#81940000000
0!
0*
09
0>
0C
#81950000000
1!
1*
b101 6
19
1>
1C
b101 G
#81960000000
0!
0*
09
0>
0C
#81970000000
1!
1*
b110 6
19
1>
1C
b110 G
#81980000000
0!
0*
09
0>
0C
#81990000000
1!
1*
b111 6
19
1>
1C
b111 G
#82000000000
0!
0*
09
0>
0C
#82010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#82020000000
0!
0*
09
0>
0C
#82030000000
1!
1*
b1 6
19
1>
1C
b1 G
#82040000000
0!
0*
09
0>
0C
#82050000000
1!
1*
b10 6
19
1>
1C
b10 G
#82060000000
0!
0*
09
0>
0C
#82070000000
1!
1*
b11 6
19
1>
1C
b11 G
#82080000000
0!
0*
09
0>
0C
#82090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#82100000000
0!
0*
09
0>
0C
#82110000000
1!
1*
b101 6
19
1>
1C
b101 G
#82120000000
0!
0*
09
0>
0C
#82130000000
1!
1*
b110 6
19
1>
1C
b110 G
#82140000000
0!
0*
09
0>
0C
#82150000000
1!
1*
b111 6
19
1>
1C
b111 G
#82160000000
0!
0*
09
0>
0C
#82170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#82180000000
0!
0*
09
0>
0C
#82190000000
1!
1*
b1 6
19
1>
1C
b1 G
#82200000000
0!
0*
09
0>
0C
#82210000000
1!
1*
b10 6
19
1>
1C
b10 G
#82220000000
0!
0*
09
0>
0C
#82230000000
1!
1*
b11 6
19
1>
1C
b11 G
#82240000000
0!
0*
09
0>
0C
#82250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#82260000000
0!
0*
09
0>
0C
#82270000000
1!
1*
b101 6
19
1>
1C
b101 G
#82280000000
0!
0*
09
0>
0C
#82290000000
1!
1*
b110 6
19
1>
1C
b110 G
#82300000000
0!
0*
09
0>
0C
#82310000000
1!
1*
b111 6
19
1>
1C
b111 G
#82320000000
0!
1"
0*
1+
09
1:
0>
0C
#82330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#82340000000
0!
0*
09
0>
0C
#82350000000
1!
1*
b1 6
19
1>
1C
b1 G
#82360000000
0!
0*
09
0>
0C
#82370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#82380000000
0!
0*
09
0>
0C
#82390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#82400000000
0!
0*
09
0>
0C
#82410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#82420000000
0!
0*
09
0>
0C
#82430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#82440000000
0!
0#
0*
0,
09
0>
0?
0C
#82450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#82460000000
0!
0*
09
0>
0C
#82470000000
1!
1*
19
1>
1C
#82480000000
0!
0*
09
0>
0C
#82490000000
1!
1*
19
1>
1C
#82500000000
0!
0*
09
0>
0C
#82510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#82520000000
0!
0*
09
0>
0C
#82530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#82540000000
0!
0*
09
0>
0C
#82550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#82560000000
0!
0*
09
0>
0C
#82570000000
1!
1*
b10 6
19
1>
1C
b10 G
#82580000000
0!
0*
09
0>
0C
#82590000000
1!
1*
b11 6
19
1>
1C
b11 G
#82600000000
0!
0*
09
0>
0C
#82610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#82620000000
0!
0*
09
0>
0C
#82630000000
1!
1*
b101 6
19
1>
1C
b101 G
#82640000000
0!
0*
09
0>
0C
#82650000000
1!
1*
b110 6
19
1>
1C
b110 G
#82660000000
0!
0*
09
0>
0C
#82670000000
1!
1*
b111 6
19
1>
1C
b111 G
#82680000000
0!
0*
09
0>
0C
#82690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#82700000000
0!
0*
09
0>
0C
#82710000000
1!
1*
b1 6
19
1>
1C
b1 G
#82720000000
0!
0*
09
0>
0C
#82730000000
1!
1*
b10 6
19
1>
1C
b10 G
#82740000000
0!
0*
09
0>
0C
#82750000000
1!
1*
b11 6
19
1>
1C
b11 G
#82760000000
0!
0*
09
0>
0C
#82770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#82780000000
0!
0*
09
0>
0C
#82790000000
1!
1*
b101 6
19
1>
1C
b101 G
#82800000000
0!
0*
09
0>
0C
#82810000000
1!
1*
b110 6
19
1>
1C
b110 G
#82820000000
0!
0*
09
0>
0C
#82830000000
1!
1*
b111 6
19
1>
1C
b111 G
#82840000000
0!
0*
09
0>
0C
#82850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#82860000000
0!
0*
09
0>
0C
#82870000000
1!
1*
b1 6
19
1>
1C
b1 G
#82880000000
0!
0*
09
0>
0C
#82890000000
1!
1*
b10 6
19
1>
1C
b10 G
#82900000000
0!
0*
09
0>
0C
#82910000000
1!
1*
b11 6
19
1>
1C
b11 G
#82920000000
0!
0*
09
0>
0C
#82930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#82940000000
0!
0*
09
0>
0C
#82950000000
1!
1*
b101 6
19
1>
1C
b101 G
#82960000000
0!
0*
09
0>
0C
#82970000000
1!
1*
b110 6
19
1>
1C
b110 G
#82980000000
0!
0*
09
0>
0C
#82990000000
1!
1*
b111 6
19
1>
1C
b111 G
#83000000000
0!
1"
0*
1+
09
1:
0>
0C
#83010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#83020000000
0!
0*
09
0>
0C
#83030000000
1!
1*
b1 6
19
1>
1C
b1 G
#83040000000
0!
0*
09
0>
0C
#83050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#83060000000
0!
0*
09
0>
0C
#83070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#83080000000
0!
0*
09
0>
0C
#83090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#83100000000
0!
0*
09
0>
0C
#83110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#83120000000
0!
0#
0*
0,
09
0>
0?
0C
#83130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#83140000000
0!
0*
09
0>
0C
#83150000000
1!
1*
19
1>
1C
#83160000000
0!
0*
09
0>
0C
#83170000000
1!
1*
19
1>
1C
#83180000000
0!
0*
09
0>
0C
#83190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#83200000000
0!
0*
09
0>
0C
#83210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#83220000000
0!
0*
09
0>
0C
#83230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#83240000000
0!
0*
09
0>
0C
#83250000000
1!
1*
b10 6
19
1>
1C
b10 G
#83260000000
0!
0*
09
0>
0C
#83270000000
1!
1*
b11 6
19
1>
1C
b11 G
#83280000000
0!
0*
09
0>
0C
#83290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#83300000000
0!
0*
09
0>
0C
#83310000000
1!
1*
b101 6
19
1>
1C
b101 G
#83320000000
0!
0*
09
0>
0C
#83330000000
1!
1*
b110 6
19
1>
1C
b110 G
#83340000000
0!
0*
09
0>
0C
#83350000000
1!
1*
b111 6
19
1>
1C
b111 G
#83360000000
0!
0*
09
0>
0C
#83370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#83380000000
0!
0*
09
0>
0C
#83390000000
1!
1*
b1 6
19
1>
1C
b1 G
#83400000000
0!
0*
09
0>
0C
#83410000000
1!
1*
b10 6
19
1>
1C
b10 G
#83420000000
0!
0*
09
0>
0C
#83430000000
1!
1*
b11 6
19
1>
1C
b11 G
#83440000000
0!
0*
09
0>
0C
#83450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#83460000000
0!
0*
09
0>
0C
#83470000000
1!
1*
b101 6
19
1>
1C
b101 G
#83480000000
0!
0*
09
0>
0C
#83490000000
1!
1*
b110 6
19
1>
1C
b110 G
#83500000000
0!
0*
09
0>
0C
#83510000000
1!
1*
b111 6
19
1>
1C
b111 G
#83520000000
0!
0*
09
0>
0C
#83530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#83540000000
0!
0*
09
0>
0C
#83550000000
1!
1*
b1 6
19
1>
1C
b1 G
#83560000000
0!
0*
09
0>
0C
#83570000000
1!
1*
b10 6
19
1>
1C
b10 G
#83580000000
0!
0*
09
0>
0C
#83590000000
1!
1*
b11 6
19
1>
1C
b11 G
#83600000000
0!
0*
09
0>
0C
#83610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#83620000000
0!
0*
09
0>
0C
#83630000000
1!
1*
b101 6
19
1>
1C
b101 G
#83640000000
0!
0*
09
0>
0C
#83650000000
1!
1*
b110 6
19
1>
1C
b110 G
#83660000000
0!
0*
09
0>
0C
#83670000000
1!
1*
b111 6
19
1>
1C
b111 G
#83680000000
0!
1"
0*
1+
09
1:
0>
0C
#83690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#83700000000
0!
0*
09
0>
0C
#83710000000
1!
1*
b1 6
19
1>
1C
b1 G
#83720000000
0!
0*
09
0>
0C
#83730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#83740000000
0!
0*
09
0>
0C
#83750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#83760000000
0!
0*
09
0>
0C
#83770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#83780000000
0!
0*
09
0>
0C
#83790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#83800000000
0!
0#
0*
0,
09
0>
0?
0C
#83810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#83820000000
0!
0*
09
0>
0C
#83830000000
1!
1*
19
1>
1C
#83840000000
0!
0*
09
0>
0C
#83850000000
1!
1*
19
1>
1C
#83860000000
0!
0*
09
0>
0C
#83870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#83880000000
0!
0*
09
0>
0C
#83890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#83900000000
0!
0*
09
0>
0C
#83910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#83920000000
0!
0*
09
0>
0C
#83930000000
1!
1*
b10 6
19
1>
1C
b10 G
#83940000000
0!
0*
09
0>
0C
#83950000000
1!
1*
b11 6
19
1>
1C
b11 G
#83960000000
0!
0*
09
0>
0C
#83970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#83980000000
0!
0*
09
0>
0C
#83990000000
1!
1*
b101 6
19
1>
1C
b101 G
#84000000000
0!
0*
09
0>
0C
#84010000000
1!
1*
b110 6
19
1>
1C
b110 G
#84020000000
0!
0*
09
0>
0C
#84030000000
1!
1*
b111 6
19
1>
1C
b111 G
#84040000000
0!
0*
09
0>
0C
#84050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#84060000000
0!
0*
09
0>
0C
#84070000000
1!
1*
b1 6
19
1>
1C
b1 G
#84080000000
0!
0*
09
0>
0C
#84090000000
1!
1*
b10 6
19
1>
1C
b10 G
#84100000000
0!
0*
09
0>
0C
#84110000000
1!
1*
b11 6
19
1>
1C
b11 G
#84120000000
0!
0*
09
0>
0C
#84130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#84140000000
0!
0*
09
0>
0C
#84150000000
1!
1*
b101 6
19
1>
1C
b101 G
#84160000000
0!
0*
09
0>
0C
#84170000000
1!
1*
b110 6
19
1>
1C
b110 G
#84180000000
0!
0*
09
0>
0C
#84190000000
1!
1*
b111 6
19
1>
1C
b111 G
#84200000000
0!
0*
09
0>
0C
#84210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#84220000000
0!
0*
09
0>
0C
#84230000000
1!
1*
b1 6
19
1>
1C
b1 G
#84240000000
0!
0*
09
0>
0C
#84250000000
1!
1*
b10 6
19
1>
1C
b10 G
#84260000000
0!
0*
09
0>
0C
#84270000000
1!
1*
b11 6
19
1>
1C
b11 G
#84280000000
0!
0*
09
0>
0C
#84290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#84300000000
0!
0*
09
0>
0C
#84310000000
1!
1*
b101 6
19
1>
1C
b101 G
#84320000000
0!
0*
09
0>
0C
#84330000000
1!
1*
b110 6
19
1>
1C
b110 G
#84340000000
0!
0*
09
0>
0C
#84350000000
1!
1*
b111 6
19
1>
1C
b111 G
#84360000000
0!
1"
0*
1+
09
1:
0>
0C
#84370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#84380000000
0!
0*
09
0>
0C
#84390000000
1!
1*
b1 6
19
1>
1C
b1 G
#84400000000
0!
0*
09
0>
0C
#84410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#84420000000
0!
0*
09
0>
0C
#84430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#84440000000
0!
0*
09
0>
0C
#84450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#84460000000
0!
0*
09
0>
0C
#84470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#84480000000
0!
0#
0*
0,
09
0>
0?
0C
#84490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#84500000000
0!
0*
09
0>
0C
#84510000000
1!
1*
19
1>
1C
#84520000000
0!
0*
09
0>
0C
#84530000000
1!
1*
19
1>
1C
#84540000000
0!
0*
09
0>
0C
#84550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#84560000000
0!
0*
09
0>
0C
#84570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#84580000000
0!
0*
09
0>
0C
#84590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#84600000000
0!
0*
09
0>
0C
#84610000000
1!
1*
b10 6
19
1>
1C
b10 G
#84620000000
0!
0*
09
0>
0C
#84630000000
1!
1*
b11 6
19
1>
1C
b11 G
#84640000000
0!
0*
09
0>
0C
#84650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#84660000000
0!
0*
09
0>
0C
#84670000000
1!
1*
b101 6
19
1>
1C
b101 G
#84680000000
0!
0*
09
0>
0C
#84690000000
1!
1*
b110 6
19
1>
1C
b110 G
#84700000000
0!
0*
09
0>
0C
#84710000000
1!
1*
b111 6
19
1>
1C
b111 G
#84720000000
0!
0*
09
0>
0C
#84730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#84740000000
0!
0*
09
0>
0C
#84750000000
1!
1*
b1 6
19
1>
1C
b1 G
#84760000000
0!
0*
09
0>
0C
#84770000000
1!
1*
b10 6
19
1>
1C
b10 G
#84780000000
0!
0*
09
0>
0C
#84790000000
1!
1*
b11 6
19
1>
1C
b11 G
#84800000000
0!
0*
09
0>
0C
#84810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#84820000000
0!
0*
09
0>
0C
#84830000000
1!
1*
b101 6
19
1>
1C
b101 G
#84840000000
0!
0*
09
0>
0C
#84850000000
1!
1*
b110 6
19
1>
1C
b110 G
#84860000000
0!
0*
09
0>
0C
#84870000000
1!
1*
b111 6
19
1>
1C
b111 G
#84880000000
0!
0*
09
0>
0C
#84890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#84900000000
0!
0*
09
0>
0C
#84910000000
1!
1*
b1 6
19
1>
1C
b1 G
#84920000000
0!
0*
09
0>
0C
#84930000000
1!
1*
b10 6
19
1>
1C
b10 G
#84940000000
0!
0*
09
0>
0C
#84950000000
1!
1*
b11 6
19
1>
1C
b11 G
#84960000000
0!
0*
09
0>
0C
#84970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#84980000000
0!
0*
09
0>
0C
#84990000000
1!
1*
b101 6
19
1>
1C
b101 G
#85000000000
0!
0*
09
0>
0C
#85010000000
1!
1*
b110 6
19
1>
1C
b110 G
#85020000000
0!
0*
09
0>
0C
#85030000000
1!
1*
b111 6
19
1>
1C
b111 G
#85040000000
0!
1"
0*
1+
09
1:
0>
0C
#85050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#85060000000
0!
0*
09
0>
0C
#85070000000
1!
1*
b1 6
19
1>
1C
b1 G
#85080000000
0!
0*
09
0>
0C
#85090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#85100000000
0!
0*
09
0>
0C
#85110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#85120000000
0!
0*
09
0>
0C
#85130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#85140000000
0!
0*
09
0>
0C
#85150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#85160000000
0!
0#
0*
0,
09
0>
0?
0C
#85170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#85180000000
0!
0*
09
0>
0C
#85190000000
1!
1*
19
1>
1C
#85200000000
0!
0*
09
0>
0C
#85210000000
1!
1*
19
1>
1C
#85220000000
0!
0*
09
0>
0C
#85230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#85240000000
0!
0*
09
0>
0C
#85250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#85260000000
0!
0*
09
0>
0C
#85270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#85280000000
0!
0*
09
0>
0C
#85290000000
1!
1*
b10 6
19
1>
1C
b10 G
#85300000000
0!
0*
09
0>
0C
#85310000000
1!
1*
b11 6
19
1>
1C
b11 G
#85320000000
0!
0*
09
0>
0C
#85330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#85340000000
0!
0*
09
0>
0C
#85350000000
1!
1*
b101 6
19
1>
1C
b101 G
#85360000000
0!
0*
09
0>
0C
#85370000000
1!
1*
b110 6
19
1>
1C
b110 G
#85380000000
0!
0*
09
0>
0C
#85390000000
1!
1*
b111 6
19
1>
1C
b111 G
#85400000000
0!
0*
09
0>
0C
#85410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#85420000000
0!
0*
09
0>
0C
#85430000000
1!
1*
b1 6
19
1>
1C
b1 G
#85440000000
0!
0*
09
0>
0C
#85450000000
1!
1*
b10 6
19
1>
1C
b10 G
#85460000000
0!
0*
09
0>
0C
#85470000000
1!
1*
b11 6
19
1>
1C
b11 G
#85480000000
0!
0*
09
0>
0C
#85490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#85500000000
0!
0*
09
0>
0C
#85510000000
1!
1*
b101 6
19
1>
1C
b101 G
#85520000000
0!
0*
09
0>
0C
#85530000000
1!
1*
b110 6
19
1>
1C
b110 G
#85540000000
0!
0*
09
0>
0C
#85550000000
1!
1*
b111 6
19
1>
1C
b111 G
#85560000000
0!
0*
09
0>
0C
#85570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#85580000000
0!
0*
09
0>
0C
#85590000000
1!
1*
b1 6
19
1>
1C
b1 G
#85600000000
0!
0*
09
0>
0C
#85610000000
1!
1*
b10 6
19
1>
1C
b10 G
#85620000000
0!
0*
09
0>
0C
#85630000000
1!
1*
b11 6
19
1>
1C
b11 G
#85640000000
0!
0*
09
0>
0C
#85650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#85660000000
0!
0*
09
0>
0C
#85670000000
1!
1*
b101 6
19
1>
1C
b101 G
#85680000000
0!
0*
09
0>
0C
#85690000000
1!
1*
b110 6
19
1>
1C
b110 G
#85700000000
0!
0*
09
0>
0C
#85710000000
1!
1*
b111 6
19
1>
1C
b111 G
#85720000000
0!
1"
0*
1+
09
1:
0>
0C
#85730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#85740000000
0!
0*
09
0>
0C
#85750000000
1!
1*
b1 6
19
1>
1C
b1 G
#85760000000
0!
0*
09
0>
0C
#85770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#85780000000
0!
0*
09
0>
0C
#85790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#85800000000
0!
0*
09
0>
0C
#85810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#85820000000
0!
0*
09
0>
0C
#85830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#85840000000
0!
0#
0*
0,
09
0>
0?
0C
#85850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#85860000000
0!
0*
09
0>
0C
#85870000000
1!
1*
19
1>
1C
#85880000000
0!
0*
09
0>
0C
#85890000000
1!
1*
19
1>
1C
#85900000000
0!
0*
09
0>
0C
#85910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#85920000000
0!
0*
09
0>
0C
#85930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#85940000000
0!
0*
09
0>
0C
#85950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#85960000000
0!
0*
09
0>
0C
#85970000000
1!
1*
b10 6
19
1>
1C
b10 G
#85980000000
0!
0*
09
0>
0C
#85990000000
1!
1*
b11 6
19
1>
1C
b11 G
#86000000000
0!
0*
09
0>
0C
#86010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#86020000000
0!
0*
09
0>
0C
#86030000000
1!
1*
b101 6
19
1>
1C
b101 G
#86040000000
0!
0*
09
0>
0C
#86050000000
1!
1*
b110 6
19
1>
1C
b110 G
#86060000000
0!
0*
09
0>
0C
#86070000000
1!
1*
b111 6
19
1>
1C
b111 G
#86080000000
0!
0*
09
0>
0C
#86090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#86100000000
0!
0*
09
0>
0C
#86110000000
1!
1*
b1 6
19
1>
1C
b1 G
#86120000000
0!
0*
09
0>
0C
#86130000000
1!
1*
b10 6
19
1>
1C
b10 G
#86140000000
0!
0*
09
0>
0C
#86150000000
1!
1*
b11 6
19
1>
1C
b11 G
#86160000000
0!
0*
09
0>
0C
#86170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#86180000000
0!
0*
09
0>
0C
#86190000000
1!
1*
b101 6
19
1>
1C
b101 G
#86200000000
0!
0*
09
0>
0C
#86210000000
1!
1*
b110 6
19
1>
1C
b110 G
#86220000000
0!
0*
09
0>
0C
#86230000000
1!
1*
b111 6
19
1>
1C
b111 G
#86240000000
0!
0*
09
0>
0C
#86250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#86260000000
0!
0*
09
0>
0C
#86270000000
1!
1*
b1 6
19
1>
1C
b1 G
#86280000000
0!
0*
09
0>
0C
#86290000000
1!
1*
b10 6
19
1>
1C
b10 G
#86300000000
0!
0*
09
0>
0C
#86310000000
1!
1*
b11 6
19
1>
1C
b11 G
#86320000000
0!
0*
09
0>
0C
#86330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#86340000000
0!
0*
09
0>
0C
#86350000000
1!
1*
b101 6
19
1>
1C
b101 G
#86360000000
0!
0*
09
0>
0C
#86370000000
1!
1*
b110 6
19
1>
1C
b110 G
#86380000000
0!
0*
09
0>
0C
#86390000000
1!
1*
b111 6
19
1>
1C
b111 G
#86400000000
0!
1"
0*
1+
09
1:
0>
0C
#86410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#86420000000
0!
0*
09
0>
0C
#86430000000
1!
1*
b1 6
19
1>
1C
b1 G
#86440000000
0!
0*
09
0>
0C
#86450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#86460000000
0!
0*
09
0>
0C
#86470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#86480000000
0!
0*
09
0>
0C
#86490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#86500000000
0!
0*
09
0>
0C
#86510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#86520000000
0!
0#
0*
0,
09
0>
0?
0C
#86530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#86540000000
0!
0*
09
0>
0C
#86550000000
1!
1*
19
1>
1C
#86560000000
0!
0*
09
0>
0C
#86570000000
1!
1*
19
1>
1C
#86580000000
0!
0*
09
0>
0C
#86590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#86600000000
0!
0*
09
0>
0C
#86610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#86620000000
0!
0*
09
0>
0C
#86630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#86640000000
0!
0*
09
0>
0C
#86650000000
1!
1*
b10 6
19
1>
1C
b10 G
#86660000000
0!
0*
09
0>
0C
#86670000000
1!
1*
b11 6
19
1>
1C
b11 G
#86680000000
0!
0*
09
0>
0C
#86690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#86700000000
0!
0*
09
0>
0C
#86710000000
1!
1*
b101 6
19
1>
1C
b101 G
#86720000000
0!
0*
09
0>
0C
#86730000000
1!
1*
b110 6
19
1>
1C
b110 G
#86740000000
0!
0*
09
0>
0C
#86750000000
1!
1*
b111 6
19
1>
1C
b111 G
#86760000000
0!
0*
09
0>
0C
#86770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#86780000000
0!
0*
09
0>
0C
#86790000000
1!
1*
b1 6
19
1>
1C
b1 G
#86800000000
0!
0*
09
0>
0C
#86810000000
1!
1*
b10 6
19
1>
1C
b10 G
#86820000000
0!
0*
09
0>
0C
#86830000000
1!
1*
b11 6
19
1>
1C
b11 G
#86840000000
0!
0*
09
0>
0C
#86850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#86860000000
0!
0*
09
0>
0C
#86870000000
1!
1*
b101 6
19
1>
1C
b101 G
#86880000000
0!
0*
09
0>
0C
#86890000000
1!
1*
b110 6
19
1>
1C
b110 G
#86900000000
0!
0*
09
0>
0C
#86910000000
1!
1*
b111 6
19
1>
1C
b111 G
#86920000000
0!
0*
09
0>
0C
#86930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#86940000000
0!
0*
09
0>
0C
#86950000000
1!
1*
b1 6
19
1>
1C
b1 G
#86960000000
0!
0*
09
0>
0C
#86970000000
1!
1*
b10 6
19
1>
1C
b10 G
#86980000000
0!
0*
09
0>
0C
#86990000000
1!
1*
b11 6
19
1>
1C
b11 G
#87000000000
0!
0*
09
0>
0C
#87010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#87020000000
0!
0*
09
0>
0C
#87030000000
1!
1*
b101 6
19
1>
1C
b101 G
#87040000000
0!
0*
09
0>
0C
#87050000000
1!
1*
b110 6
19
1>
1C
b110 G
#87060000000
0!
0*
09
0>
0C
#87070000000
1!
1*
b111 6
19
1>
1C
b111 G
#87080000000
0!
1"
0*
1+
09
1:
0>
0C
#87090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#87100000000
0!
0*
09
0>
0C
#87110000000
1!
1*
b1 6
19
1>
1C
b1 G
#87120000000
0!
0*
09
0>
0C
#87130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#87140000000
0!
0*
09
0>
0C
#87150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#87160000000
0!
0*
09
0>
0C
#87170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#87180000000
0!
0*
09
0>
0C
#87190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#87200000000
0!
0#
0*
0,
09
0>
0?
0C
#87210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#87220000000
0!
0*
09
0>
0C
#87230000000
1!
1*
19
1>
1C
#87240000000
0!
0*
09
0>
0C
#87250000000
1!
1*
19
1>
1C
#87260000000
0!
0*
09
0>
0C
#87270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#87280000000
0!
0*
09
0>
0C
#87290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#87300000000
0!
0*
09
0>
0C
#87310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#87320000000
0!
0*
09
0>
0C
#87330000000
1!
1*
b10 6
19
1>
1C
b10 G
#87340000000
0!
0*
09
0>
0C
#87350000000
1!
1*
b11 6
19
1>
1C
b11 G
#87360000000
0!
0*
09
0>
0C
#87370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#87380000000
0!
0*
09
0>
0C
#87390000000
1!
1*
b101 6
19
1>
1C
b101 G
#87400000000
0!
0*
09
0>
0C
#87410000000
1!
1*
b110 6
19
1>
1C
b110 G
#87420000000
0!
0*
09
0>
0C
#87430000000
1!
1*
b111 6
19
1>
1C
b111 G
#87440000000
0!
0*
09
0>
0C
#87450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#87460000000
0!
0*
09
0>
0C
#87470000000
1!
1*
b1 6
19
1>
1C
b1 G
#87480000000
0!
0*
09
0>
0C
#87490000000
1!
1*
b10 6
19
1>
1C
b10 G
#87500000000
0!
0*
09
0>
0C
#87510000000
1!
1*
b11 6
19
1>
1C
b11 G
#87520000000
0!
0*
09
0>
0C
#87530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#87540000000
0!
0*
09
0>
0C
#87550000000
1!
1*
b101 6
19
1>
1C
b101 G
#87560000000
0!
0*
09
0>
0C
#87570000000
1!
1*
b110 6
19
1>
1C
b110 G
#87580000000
0!
0*
09
0>
0C
#87590000000
1!
1*
b111 6
19
1>
1C
b111 G
#87600000000
0!
0*
09
0>
0C
#87610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#87620000000
0!
0*
09
0>
0C
#87630000000
1!
1*
b1 6
19
1>
1C
b1 G
#87640000000
0!
0*
09
0>
0C
#87650000000
1!
1*
b10 6
19
1>
1C
b10 G
#87660000000
0!
0*
09
0>
0C
#87670000000
1!
1*
b11 6
19
1>
1C
b11 G
#87680000000
0!
0*
09
0>
0C
#87690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#87700000000
0!
0*
09
0>
0C
#87710000000
1!
1*
b101 6
19
1>
1C
b101 G
#87720000000
0!
0*
09
0>
0C
#87730000000
1!
1*
b110 6
19
1>
1C
b110 G
#87740000000
0!
0*
09
0>
0C
#87750000000
1!
1*
b111 6
19
1>
1C
b111 G
#87760000000
0!
1"
0*
1+
09
1:
0>
0C
#87770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#87780000000
0!
0*
09
0>
0C
#87790000000
1!
1*
b1 6
19
1>
1C
b1 G
#87800000000
0!
0*
09
0>
0C
#87810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#87820000000
0!
0*
09
0>
0C
#87830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#87840000000
0!
0*
09
0>
0C
#87850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#87860000000
0!
0*
09
0>
0C
#87870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#87880000000
0!
0#
0*
0,
09
0>
0?
0C
#87890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#87900000000
0!
0*
09
0>
0C
#87910000000
1!
1*
19
1>
1C
#87920000000
0!
0*
09
0>
0C
#87930000000
1!
1*
19
1>
1C
#87940000000
0!
0*
09
0>
0C
#87950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#87960000000
0!
0*
09
0>
0C
#87970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#87980000000
0!
0*
09
0>
0C
#87990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#88000000000
0!
0*
09
0>
0C
#88010000000
1!
1*
b10 6
19
1>
1C
b10 G
#88020000000
0!
0*
09
0>
0C
#88030000000
1!
1*
b11 6
19
1>
1C
b11 G
#88040000000
0!
0*
09
0>
0C
#88050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#88060000000
0!
0*
09
0>
0C
#88070000000
1!
1*
b101 6
19
1>
1C
b101 G
#88080000000
0!
0*
09
0>
0C
#88090000000
1!
1*
b110 6
19
1>
1C
b110 G
#88100000000
0!
0*
09
0>
0C
#88110000000
1!
1*
b111 6
19
1>
1C
b111 G
#88120000000
0!
0*
09
0>
0C
#88130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#88140000000
0!
0*
09
0>
0C
#88150000000
1!
1*
b1 6
19
1>
1C
b1 G
#88160000000
0!
0*
09
0>
0C
#88170000000
1!
1*
b10 6
19
1>
1C
b10 G
#88180000000
0!
0*
09
0>
0C
#88190000000
1!
1*
b11 6
19
1>
1C
b11 G
#88200000000
0!
0*
09
0>
0C
#88210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#88220000000
0!
0*
09
0>
0C
#88230000000
1!
1*
b101 6
19
1>
1C
b101 G
#88240000000
0!
0*
09
0>
0C
#88250000000
1!
1*
b110 6
19
1>
1C
b110 G
#88260000000
0!
0*
09
0>
0C
#88270000000
1!
1*
b111 6
19
1>
1C
b111 G
#88280000000
0!
0*
09
0>
0C
#88290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#88300000000
0!
0*
09
0>
0C
#88310000000
1!
1*
b1 6
19
1>
1C
b1 G
#88320000000
0!
0*
09
0>
0C
#88330000000
1!
1*
b10 6
19
1>
1C
b10 G
#88340000000
0!
0*
09
0>
0C
#88350000000
1!
1*
b11 6
19
1>
1C
b11 G
#88360000000
0!
0*
09
0>
0C
#88370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#88380000000
0!
0*
09
0>
0C
#88390000000
1!
1*
b101 6
19
1>
1C
b101 G
#88400000000
0!
0*
09
0>
0C
#88410000000
1!
1*
b110 6
19
1>
1C
b110 G
#88420000000
0!
0*
09
0>
0C
#88430000000
1!
1*
b111 6
19
1>
1C
b111 G
#88440000000
0!
1"
0*
1+
09
1:
0>
0C
#88450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#88460000000
0!
0*
09
0>
0C
#88470000000
1!
1*
b1 6
19
1>
1C
b1 G
#88480000000
0!
0*
09
0>
0C
#88490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#88500000000
0!
0*
09
0>
0C
#88510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#88520000000
0!
0*
09
0>
0C
#88530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#88540000000
0!
0*
09
0>
0C
#88550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#88560000000
0!
0#
0*
0,
09
0>
0?
0C
#88570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#88580000000
0!
0*
09
0>
0C
#88590000000
1!
1*
19
1>
1C
#88600000000
0!
0*
09
0>
0C
#88610000000
1!
1*
19
1>
1C
#88620000000
0!
0*
09
0>
0C
#88630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#88640000000
0!
0*
09
0>
0C
#88650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#88660000000
0!
0*
09
0>
0C
#88670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#88680000000
0!
0*
09
0>
0C
#88690000000
1!
1*
b10 6
19
1>
1C
b10 G
#88700000000
0!
0*
09
0>
0C
#88710000000
1!
1*
b11 6
19
1>
1C
b11 G
#88720000000
0!
0*
09
0>
0C
#88730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#88740000000
0!
0*
09
0>
0C
#88750000000
1!
1*
b101 6
19
1>
1C
b101 G
#88760000000
0!
0*
09
0>
0C
#88770000000
1!
1*
b110 6
19
1>
1C
b110 G
#88780000000
0!
0*
09
0>
0C
#88790000000
1!
1*
b111 6
19
1>
1C
b111 G
#88800000000
0!
0*
09
0>
0C
#88810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#88820000000
0!
0*
09
0>
0C
#88830000000
1!
1*
b1 6
19
1>
1C
b1 G
#88840000000
0!
0*
09
0>
0C
#88850000000
1!
1*
b10 6
19
1>
1C
b10 G
#88860000000
0!
0*
09
0>
0C
#88870000000
1!
1*
b11 6
19
1>
1C
b11 G
#88880000000
0!
0*
09
0>
0C
#88890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#88900000000
0!
0*
09
0>
0C
#88910000000
1!
1*
b101 6
19
1>
1C
b101 G
#88920000000
0!
0*
09
0>
0C
#88930000000
1!
1*
b110 6
19
1>
1C
b110 G
#88940000000
0!
0*
09
0>
0C
#88950000000
1!
1*
b111 6
19
1>
1C
b111 G
#88960000000
0!
0*
09
0>
0C
#88970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#88980000000
0!
0*
09
0>
0C
#88990000000
1!
1*
b1 6
19
1>
1C
b1 G
#89000000000
0!
0*
09
0>
0C
#89010000000
1!
1*
b10 6
19
1>
1C
b10 G
#89020000000
0!
0*
09
0>
0C
#89030000000
1!
1*
b11 6
19
1>
1C
b11 G
#89040000000
0!
0*
09
0>
0C
#89050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#89060000000
0!
0*
09
0>
0C
#89070000000
1!
1*
b101 6
19
1>
1C
b101 G
#89080000000
0!
0*
09
0>
0C
#89090000000
1!
1*
b110 6
19
1>
1C
b110 G
#89100000000
0!
0*
09
0>
0C
#89110000000
1!
1*
b111 6
19
1>
1C
b111 G
#89120000000
0!
1"
0*
1+
09
1:
0>
0C
#89130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#89140000000
0!
0*
09
0>
0C
#89150000000
1!
1*
b1 6
19
1>
1C
b1 G
#89160000000
0!
0*
09
0>
0C
#89170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#89180000000
0!
0*
09
0>
0C
#89190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#89200000000
0!
0*
09
0>
0C
#89210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#89220000000
0!
0*
09
0>
0C
#89230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#89240000000
0!
0#
0*
0,
09
0>
0?
0C
#89250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#89260000000
0!
0*
09
0>
0C
#89270000000
1!
1*
19
1>
1C
#89280000000
0!
0*
09
0>
0C
#89290000000
1!
1*
19
1>
1C
#89300000000
0!
0*
09
0>
0C
#89310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#89320000000
0!
0*
09
0>
0C
#89330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#89340000000
0!
0*
09
0>
0C
#89350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#89360000000
0!
0*
09
0>
0C
#89370000000
1!
1*
b10 6
19
1>
1C
b10 G
#89380000000
0!
0*
09
0>
0C
#89390000000
1!
1*
b11 6
19
1>
1C
b11 G
#89400000000
0!
0*
09
0>
0C
#89410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#89420000000
0!
0*
09
0>
0C
#89430000000
1!
1*
b101 6
19
1>
1C
b101 G
#89440000000
0!
0*
09
0>
0C
#89450000000
1!
1*
b110 6
19
1>
1C
b110 G
#89460000000
0!
0*
09
0>
0C
#89470000000
1!
1*
b111 6
19
1>
1C
b111 G
#89480000000
0!
0*
09
0>
0C
#89490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#89500000000
0!
0*
09
0>
0C
#89510000000
1!
1*
b1 6
19
1>
1C
b1 G
#89520000000
0!
0*
09
0>
0C
#89530000000
1!
1*
b10 6
19
1>
1C
b10 G
#89540000000
0!
0*
09
0>
0C
#89550000000
1!
1*
b11 6
19
1>
1C
b11 G
#89560000000
0!
0*
09
0>
0C
#89570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#89580000000
0!
0*
09
0>
0C
#89590000000
1!
1*
b101 6
19
1>
1C
b101 G
#89600000000
0!
0*
09
0>
0C
#89610000000
1!
1*
b110 6
19
1>
1C
b110 G
#89620000000
0!
0*
09
0>
0C
#89630000000
1!
1*
b111 6
19
1>
1C
b111 G
#89640000000
0!
0*
09
0>
0C
#89650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#89660000000
0!
0*
09
0>
0C
#89670000000
1!
1*
b1 6
19
1>
1C
b1 G
#89680000000
0!
0*
09
0>
0C
#89690000000
1!
1*
b10 6
19
1>
1C
b10 G
#89700000000
0!
0*
09
0>
0C
#89710000000
1!
1*
b11 6
19
1>
1C
b11 G
#89720000000
0!
0*
09
0>
0C
#89730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#89740000000
0!
0*
09
0>
0C
#89750000000
1!
1*
b101 6
19
1>
1C
b101 G
#89760000000
0!
0*
09
0>
0C
#89770000000
1!
1*
b110 6
19
1>
1C
b110 G
#89780000000
0!
0*
09
0>
0C
#89790000000
1!
1*
b111 6
19
1>
1C
b111 G
#89800000000
0!
1"
0*
1+
09
1:
0>
0C
#89810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#89820000000
0!
0*
09
0>
0C
#89830000000
1!
1*
b1 6
19
1>
1C
b1 G
#89840000000
0!
0*
09
0>
0C
#89850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#89860000000
0!
0*
09
0>
0C
#89870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#89880000000
0!
0*
09
0>
0C
#89890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#89900000000
0!
0*
09
0>
0C
#89910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#89920000000
0!
0#
0*
0,
09
0>
0?
0C
#89930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#89940000000
0!
0*
09
0>
0C
#89950000000
1!
1*
19
1>
1C
#89960000000
0!
0*
09
0>
0C
#89970000000
1!
1*
19
1>
1C
#89980000000
0!
0*
09
0>
0C
#89990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#90000000000
0!
0*
09
0>
0C
#90010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#90020000000
0!
0*
09
0>
0C
#90030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#90040000000
0!
0*
09
0>
0C
#90050000000
1!
1*
b10 6
19
1>
1C
b10 G
#90060000000
0!
0*
09
0>
0C
#90070000000
1!
1*
b11 6
19
1>
1C
b11 G
#90080000000
0!
0*
09
0>
0C
#90090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#90100000000
0!
0*
09
0>
0C
#90110000000
1!
1*
b101 6
19
1>
1C
b101 G
#90120000000
0!
0*
09
0>
0C
#90130000000
1!
1*
b110 6
19
1>
1C
b110 G
#90140000000
0!
0*
09
0>
0C
#90150000000
1!
1*
b111 6
19
1>
1C
b111 G
#90160000000
0!
0*
09
0>
0C
#90170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#90180000000
0!
0*
09
0>
0C
#90190000000
1!
1*
b1 6
19
1>
1C
b1 G
#90200000000
0!
0*
09
0>
0C
#90210000000
1!
1*
b10 6
19
1>
1C
b10 G
#90220000000
0!
0*
09
0>
0C
#90230000000
1!
1*
b11 6
19
1>
1C
b11 G
#90240000000
0!
0*
09
0>
0C
#90250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#90260000000
0!
0*
09
0>
0C
#90270000000
1!
1*
b101 6
19
1>
1C
b101 G
#90280000000
0!
0*
09
0>
0C
#90290000000
1!
1*
b110 6
19
1>
1C
b110 G
#90300000000
0!
0*
09
0>
0C
#90310000000
1!
1*
b111 6
19
1>
1C
b111 G
#90320000000
0!
0*
09
0>
0C
#90330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#90340000000
0!
0*
09
0>
0C
#90350000000
1!
1*
b1 6
19
1>
1C
b1 G
#90360000000
0!
0*
09
0>
0C
#90370000000
1!
1*
b10 6
19
1>
1C
b10 G
#90380000000
0!
0*
09
0>
0C
#90390000000
1!
1*
b11 6
19
1>
1C
b11 G
#90400000000
0!
0*
09
0>
0C
#90410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#90420000000
0!
0*
09
0>
0C
#90430000000
1!
1*
b101 6
19
1>
1C
b101 G
#90440000000
0!
0*
09
0>
0C
#90450000000
1!
1*
b110 6
19
1>
1C
b110 G
#90460000000
0!
0*
09
0>
0C
#90470000000
1!
1*
b111 6
19
1>
1C
b111 G
#90480000000
0!
1"
0*
1+
09
1:
0>
0C
#90490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#90500000000
0!
0*
09
0>
0C
#90510000000
1!
1*
b1 6
19
1>
1C
b1 G
#90520000000
0!
0*
09
0>
0C
#90530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#90540000000
0!
0*
09
0>
0C
#90550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#90560000000
0!
0*
09
0>
0C
#90570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#90580000000
0!
0*
09
0>
0C
#90590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#90600000000
0!
0#
0*
0,
09
0>
0?
0C
#90610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#90620000000
0!
0*
09
0>
0C
#90630000000
1!
1*
19
1>
1C
#90640000000
0!
0*
09
0>
0C
#90650000000
1!
1*
19
1>
1C
#90660000000
0!
0*
09
0>
0C
#90670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#90680000000
0!
0*
09
0>
0C
#90690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#90700000000
0!
0*
09
0>
0C
#90710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#90720000000
0!
0*
09
0>
0C
#90730000000
1!
1*
b10 6
19
1>
1C
b10 G
#90740000000
0!
0*
09
0>
0C
#90750000000
1!
1*
b11 6
19
1>
1C
b11 G
#90760000000
0!
0*
09
0>
0C
#90770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#90780000000
0!
0*
09
0>
0C
#90790000000
1!
1*
b101 6
19
1>
1C
b101 G
#90800000000
0!
0*
09
0>
0C
#90810000000
1!
1*
b110 6
19
1>
1C
b110 G
#90820000000
0!
0*
09
0>
0C
#90830000000
1!
1*
b111 6
19
1>
1C
b111 G
#90840000000
0!
0*
09
0>
0C
#90850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#90860000000
0!
0*
09
0>
0C
#90870000000
1!
1*
b1 6
19
1>
1C
b1 G
#90880000000
0!
0*
09
0>
0C
#90890000000
1!
1*
b10 6
19
1>
1C
b10 G
#90900000000
0!
0*
09
0>
0C
#90910000000
1!
1*
b11 6
19
1>
1C
b11 G
#90920000000
0!
0*
09
0>
0C
#90930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#90940000000
0!
0*
09
0>
0C
#90950000000
1!
1*
b101 6
19
1>
1C
b101 G
#90960000000
0!
0*
09
0>
0C
#90970000000
1!
1*
b110 6
19
1>
1C
b110 G
#90980000000
0!
0*
09
0>
0C
#90990000000
1!
1*
b111 6
19
1>
1C
b111 G
#91000000000
0!
0*
09
0>
0C
#91010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#91020000000
0!
0*
09
0>
0C
#91030000000
1!
1*
b1 6
19
1>
1C
b1 G
#91040000000
0!
0*
09
0>
0C
#91050000000
1!
1*
b10 6
19
1>
1C
b10 G
#91060000000
0!
0*
09
0>
0C
#91070000000
1!
1*
b11 6
19
1>
1C
b11 G
#91080000000
0!
0*
09
0>
0C
#91090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#91100000000
0!
0*
09
0>
0C
#91110000000
1!
1*
b101 6
19
1>
1C
b101 G
#91120000000
0!
0*
09
0>
0C
#91130000000
1!
1*
b110 6
19
1>
1C
b110 G
#91140000000
0!
0*
09
0>
0C
#91150000000
1!
1*
b111 6
19
1>
1C
b111 G
#91160000000
0!
1"
0*
1+
09
1:
0>
0C
#91170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#91180000000
0!
0*
09
0>
0C
#91190000000
1!
1*
b1 6
19
1>
1C
b1 G
#91200000000
0!
0*
09
0>
0C
#91210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#91220000000
0!
0*
09
0>
0C
#91230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#91240000000
0!
0*
09
0>
0C
#91250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#91260000000
0!
0*
09
0>
0C
#91270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#91280000000
0!
0#
0*
0,
09
0>
0?
0C
#91290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#91300000000
0!
0*
09
0>
0C
#91310000000
1!
1*
19
1>
1C
#91320000000
0!
0*
09
0>
0C
#91330000000
1!
1*
19
1>
1C
#91340000000
0!
0*
09
0>
0C
#91350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#91360000000
0!
0*
09
0>
0C
#91370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#91380000000
0!
0*
09
0>
0C
#91390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#91400000000
0!
0*
09
0>
0C
#91410000000
1!
1*
b10 6
19
1>
1C
b10 G
#91420000000
0!
0*
09
0>
0C
#91430000000
1!
1*
b11 6
19
1>
1C
b11 G
#91440000000
0!
0*
09
0>
0C
#91450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#91460000000
0!
0*
09
0>
0C
#91470000000
1!
1*
b101 6
19
1>
1C
b101 G
#91480000000
0!
0*
09
0>
0C
#91490000000
1!
1*
b110 6
19
1>
1C
b110 G
#91500000000
0!
0*
09
0>
0C
#91510000000
1!
1*
b111 6
19
1>
1C
b111 G
#91520000000
0!
0*
09
0>
0C
#91530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#91540000000
0!
0*
09
0>
0C
#91550000000
1!
1*
b1 6
19
1>
1C
b1 G
#91560000000
0!
0*
09
0>
0C
#91570000000
1!
1*
b10 6
19
1>
1C
b10 G
#91580000000
0!
0*
09
0>
0C
#91590000000
1!
1*
b11 6
19
1>
1C
b11 G
#91600000000
0!
0*
09
0>
0C
#91610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#91620000000
0!
0*
09
0>
0C
#91630000000
1!
1*
b101 6
19
1>
1C
b101 G
#91640000000
0!
0*
09
0>
0C
#91650000000
1!
1*
b110 6
19
1>
1C
b110 G
#91660000000
0!
0*
09
0>
0C
#91670000000
1!
1*
b111 6
19
1>
1C
b111 G
#91680000000
0!
0*
09
0>
0C
#91690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#91700000000
0!
0*
09
0>
0C
#91710000000
1!
1*
b1 6
19
1>
1C
b1 G
#91720000000
0!
0*
09
0>
0C
#91730000000
1!
1*
b10 6
19
1>
1C
b10 G
#91740000000
0!
0*
09
0>
0C
#91750000000
1!
1*
b11 6
19
1>
1C
b11 G
#91760000000
0!
0*
09
0>
0C
#91770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#91780000000
0!
0*
09
0>
0C
#91790000000
1!
1*
b101 6
19
1>
1C
b101 G
#91800000000
0!
0*
09
0>
0C
#91810000000
1!
1*
b110 6
19
1>
1C
b110 G
#91820000000
0!
0*
09
0>
0C
#91830000000
1!
1*
b111 6
19
1>
1C
b111 G
#91840000000
0!
1"
0*
1+
09
1:
0>
0C
#91850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#91860000000
0!
0*
09
0>
0C
#91870000000
1!
1*
b1 6
19
1>
1C
b1 G
#91880000000
0!
0*
09
0>
0C
#91890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#91900000000
0!
0*
09
0>
0C
#91910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#91920000000
0!
0*
09
0>
0C
#91930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#91940000000
0!
0*
09
0>
0C
#91950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#91960000000
0!
0#
0*
0,
09
0>
0?
0C
#91970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#91980000000
0!
0*
09
0>
0C
#91990000000
1!
1*
19
1>
1C
#92000000000
0!
0*
09
0>
0C
#92010000000
1!
1*
19
1>
1C
#92020000000
0!
0*
09
0>
0C
#92030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#92040000000
0!
0*
09
0>
0C
#92050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#92060000000
0!
0*
09
0>
0C
#92070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#92080000000
0!
0*
09
0>
0C
#92090000000
1!
1*
b10 6
19
1>
1C
b10 G
#92100000000
0!
0*
09
0>
0C
#92110000000
1!
1*
b11 6
19
1>
1C
b11 G
#92120000000
0!
0*
09
0>
0C
#92130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#92140000000
0!
0*
09
0>
0C
#92150000000
1!
1*
b101 6
19
1>
1C
b101 G
#92160000000
0!
0*
09
0>
0C
#92170000000
1!
1*
b110 6
19
1>
1C
b110 G
#92180000000
0!
0*
09
0>
0C
#92190000000
1!
1*
b111 6
19
1>
1C
b111 G
#92200000000
0!
0*
09
0>
0C
#92210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#92220000000
0!
0*
09
0>
0C
#92230000000
1!
1*
b1 6
19
1>
1C
b1 G
#92240000000
0!
0*
09
0>
0C
#92250000000
1!
1*
b10 6
19
1>
1C
b10 G
#92260000000
0!
0*
09
0>
0C
#92270000000
1!
1*
b11 6
19
1>
1C
b11 G
#92280000000
0!
0*
09
0>
0C
#92290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#92300000000
0!
0*
09
0>
0C
#92310000000
1!
1*
b101 6
19
1>
1C
b101 G
#92320000000
0!
0*
09
0>
0C
#92330000000
1!
1*
b110 6
19
1>
1C
b110 G
#92340000000
0!
0*
09
0>
0C
#92350000000
1!
1*
b111 6
19
1>
1C
b111 G
#92360000000
0!
0*
09
0>
0C
#92370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#92380000000
0!
0*
09
0>
0C
#92390000000
1!
1*
b1 6
19
1>
1C
b1 G
#92400000000
0!
0*
09
0>
0C
#92410000000
1!
1*
b10 6
19
1>
1C
b10 G
#92420000000
0!
0*
09
0>
0C
#92430000000
1!
1*
b11 6
19
1>
1C
b11 G
#92440000000
0!
0*
09
0>
0C
#92450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#92460000000
0!
0*
09
0>
0C
#92470000000
1!
1*
b101 6
19
1>
1C
b101 G
#92480000000
0!
0*
09
0>
0C
#92490000000
1!
1*
b110 6
19
1>
1C
b110 G
#92500000000
0!
0*
09
0>
0C
#92510000000
1!
1*
b111 6
19
1>
1C
b111 G
#92520000000
0!
1"
0*
1+
09
1:
0>
0C
#92530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#92540000000
0!
0*
09
0>
0C
#92550000000
1!
1*
b1 6
19
1>
1C
b1 G
#92560000000
0!
0*
09
0>
0C
#92570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#92580000000
0!
0*
09
0>
0C
#92590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#92600000000
0!
0*
09
0>
0C
#92610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#92620000000
0!
0*
09
0>
0C
#92630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#92640000000
0!
0#
0*
0,
09
0>
0?
0C
#92650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#92660000000
0!
0*
09
0>
0C
#92670000000
1!
1*
19
1>
1C
#92680000000
0!
0*
09
0>
0C
#92690000000
1!
1*
19
1>
1C
#92700000000
0!
0*
09
0>
0C
#92710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#92720000000
0!
0*
09
0>
0C
#92730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#92740000000
0!
0*
09
0>
0C
#92750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#92760000000
0!
0*
09
0>
0C
#92770000000
1!
1*
b10 6
19
1>
1C
b10 G
#92780000000
0!
0*
09
0>
0C
#92790000000
1!
1*
b11 6
19
1>
1C
b11 G
#92800000000
0!
0*
09
0>
0C
#92810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#92820000000
0!
0*
09
0>
0C
#92830000000
1!
1*
b101 6
19
1>
1C
b101 G
#92840000000
0!
0*
09
0>
0C
#92850000000
1!
1*
b110 6
19
1>
1C
b110 G
#92860000000
0!
0*
09
0>
0C
#92870000000
1!
1*
b111 6
19
1>
1C
b111 G
#92880000000
0!
0*
09
0>
0C
#92890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#92900000000
0!
0*
09
0>
0C
#92910000000
1!
1*
b1 6
19
1>
1C
b1 G
#92920000000
0!
0*
09
0>
0C
#92930000000
1!
1*
b10 6
19
1>
1C
b10 G
#92940000000
0!
0*
09
0>
0C
#92950000000
1!
1*
b11 6
19
1>
1C
b11 G
#92960000000
0!
0*
09
0>
0C
#92970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#92980000000
0!
0*
09
0>
0C
#92990000000
1!
1*
b101 6
19
1>
1C
b101 G
#93000000000
0!
0*
09
0>
0C
#93010000000
1!
1*
b110 6
19
1>
1C
b110 G
#93020000000
0!
0*
09
0>
0C
#93030000000
1!
1*
b111 6
19
1>
1C
b111 G
#93040000000
0!
0*
09
0>
0C
#93050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#93060000000
0!
0*
09
0>
0C
#93070000000
1!
1*
b1 6
19
1>
1C
b1 G
#93080000000
0!
0*
09
0>
0C
#93090000000
1!
1*
b10 6
19
1>
1C
b10 G
#93100000000
0!
0*
09
0>
0C
#93110000000
1!
1*
b11 6
19
1>
1C
b11 G
#93120000000
0!
0*
09
0>
0C
#93130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#93140000000
0!
0*
09
0>
0C
#93150000000
1!
1*
b101 6
19
1>
1C
b101 G
#93160000000
0!
0*
09
0>
0C
#93170000000
1!
1*
b110 6
19
1>
1C
b110 G
#93180000000
0!
0*
09
0>
0C
#93190000000
1!
1*
b111 6
19
1>
1C
b111 G
#93200000000
0!
1"
0*
1+
09
1:
0>
0C
#93210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#93220000000
0!
0*
09
0>
0C
#93230000000
1!
1*
b1 6
19
1>
1C
b1 G
#93240000000
0!
0*
09
0>
0C
#93250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#93260000000
0!
0*
09
0>
0C
#93270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#93280000000
0!
0*
09
0>
0C
#93290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#93300000000
0!
0*
09
0>
0C
#93310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#93320000000
0!
0#
0*
0,
09
0>
0?
0C
#93330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#93340000000
0!
0*
09
0>
0C
#93350000000
1!
1*
19
1>
1C
#93360000000
0!
0*
09
0>
0C
#93370000000
1!
1*
19
1>
1C
#93380000000
0!
0*
09
0>
0C
#93390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#93400000000
0!
0*
09
0>
0C
#93410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#93420000000
0!
0*
09
0>
0C
#93430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#93440000000
0!
0*
09
0>
0C
#93450000000
1!
1*
b10 6
19
1>
1C
b10 G
#93460000000
0!
0*
09
0>
0C
#93470000000
1!
1*
b11 6
19
1>
1C
b11 G
#93480000000
0!
0*
09
0>
0C
#93490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#93500000000
0!
0*
09
0>
0C
#93510000000
1!
1*
b101 6
19
1>
1C
b101 G
#93520000000
0!
0*
09
0>
0C
#93530000000
1!
1*
b110 6
19
1>
1C
b110 G
#93540000000
0!
0*
09
0>
0C
#93550000000
1!
1*
b111 6
19
1>
1C
b111 G
#93560000000
0!
0*
09
0>
0C
#93570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#93580000000
0!
0*
09
0>
0C
#93590000000
1!
1*
b1 6
19
1>
1C
b1 G
#93600000000
0!
0*
09
0>
0C
#93610000000
1!
1*
b10 6
19
1>
1C
b10 G
#93620000000
0!
0*
09
0>
0C
#93630000000
1!
1*
b11 6
19
1>
1C
b11 G
#93640000000
0!
0*
09
0>
0C
#93650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#93660000000
0!
0*
09
0>
0C
#93670000000
1!
1*
b101 6
19
1>
1C
b101 G
#93680000000
0!
0*
09
0>
0C
#93690000000
1!
1*
b110 6
19
1>
1C
b110 G
#93700000000
0!
0*
09
0>
0C
#93710000000
1!
1*
b111 6
19
1>
1C
b111 G
#93720000000
0!
0*
09
0>
0C
#93730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#93740000000
0!
0*
09
0>
0C
#93750000000
1!
1*
b1 6
19
1>
1C
b1 G
#93760000000
0!
0*
09
0>
0C
#93770000000
1!
1*
b10 6
19
1>
1C
b10 G
#93780000000
0!
0*
09
0>
0C
#93790000000
1!
1*
b11 6
19
1>
1C
b11 G
#93800000000
0!
0*
09
0>
0C
#93810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#93820000000
0!
0*
09
0>
0C
#93830000000
1!
1*
b101 6
19
1>
1C
b101 G
#93840000000
0!
0*
09
0>
0C
#93850000000
1!
1*
b110 6
19
1>
1C
b110 G
#93860000000
0!
0*
09
0>
0C
#93870000000
1!
1*
b111 6
19
1>
1C
b111 G
#93880000000
0!
1"
0*
1+
09
1:
0>
0C
#93890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#93900000000
0!
0*
09
0>
0C
#93910000000
1!
1*
b1 6
19
1>
1C
b1 G
#93920000000
0!
0*
09
0>
0C
#93930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#93940000000
0!
0*
09
0>
0C
#93950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#93960000000
0!
0*
09
0>
0C
#93970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#93980000000
0!
0*
09
0>
0C
#93990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#94000000000
0!
0#
0*
0,
09
0>
0?
0C
#94010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#94020000000
0!
0*
09
0>
0C
#94030000000
1!
1*
19
1>
1C
#94040000000
0!
0*
09
0>
0C
#94050000000
1!
1*
19
1>
1C
#94060000000
0!
0*
09
0>
0C
#94070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#94080000000
0!
0*
09
0>
0C
#94090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#94100000000
0!
0*
09
0>
0C
#94110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#94120000000
0!
0*
09
0>
0C
#94130000000
1!
1*
b10 6
19
1>
1C
b10 G
#94140000000
0!
0*
09
0>
0C
#94150000000
1!
1*
b11 6
19
1>
1C
b11 G
#94160000000
0!
0*
09
0>
0C
#94170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#94180000000
0!
0*
09
0>
0C
#94190000000
1!
1*
b101 6
19
1>
1C
b101 G
#94200000000
0!
0*
09
0>
0C
#94210000000
1!
1*
b110 6
19
1>
1C
b110 G
#94220000000
0!
0*
09
0>
0C
#94230000000
1!
1*
b111 6
19
1>
1C
b111 G
#94240000000
0!
0*
09
0>
0C
#94250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#94260000000
0!
0*
09
0>
0C
#94270000000
1!
1*
b1 6
19
1>
1C
b1 G
#94280000000
0!
0*
09
0>
0C
#94290000000
1!
1*
b10 6
19
1>
1C
b10 G
#94300000000
0!
0*
09
0>
0C
#94310000000
1!
1*
b11 6
19
1>
1C
b11 G
#94320000000
0!
0*
09
0>
0C
#94330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#94340000000
0!
0*
09
0>
0C
#94350000000
1!
1*
b101 6
19
1>
1C
b101 G
#94360000000
0!
0*
09
0>
0C
#94370000000
1!
1*
b110 6
19
1>
1C
b110 G
#94380000000
0!
0*
09
0>
0C
#94390000000
1!
1*
b111 6
19
1>
1C
b111 G
#94400000000
0!
0*
09
0>
0C
#94410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#94420000000
0!
0*
09
0>
0C
#94430000000
1!
1*
b1 6
19
1>
1C
b1 G
#94440000000
0!
0*
09
0>
0C
#94450000000
1!
1*
b10 6
19
1>
1C
b10 G
#94460000000
0!
0*
09
0>
0C
#94470000000
1!
1*
b11 6
19
1>
1C
b11 G
#94480000000
0!
0*
09
0>
0C
#94490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#94500000000
0!
0*
09
0>
0C
#94510000000
1!
1*
b101 6
19
1>
1C
b101 G
#94520000000
0!
0*
09
0>
0C
#94530000000
1!
1*
b110 6
19
1>
1C
b110 G
#94540000000
0!
0*
09
0>
0C
#94550000000
1!
1*
b111 6
19
1>
1C
b111 G
#94560000000
0!
1"
0*
1+
09
1:
0>
0C
#94570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#94580000000
0!
0*
09
0>
0C
#94590000000
1!
1*
b1 6
19
1>
1C
b1 G
#94600000000
0!
0*
09
0>
0C
#94610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#94620000000
0!
0*
09
0>
0C
#94630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#94640000000
0!
0*
09
0>
0C
#94650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#94660000000
0!
0*
09
0>
0C
#94670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#94680000000
0!
0#
0*
0,
09
0>
0?
0C
#94690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#94700000000
0!
0*
09
0>
0C
#94710000000
1!
1*
19
1>
1C
#94720000000
0!
0*
09
0>
0C
#94730000000
1!
1*
19
1>
1C
#94740000000
0!
0*
09
0>
0C
#94750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#94760000000
0!
0*
09
0>
0C
#94770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#94780000000
0!
0*
09
0>
0C
#94790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#94800000000
0!
0*
09
0>
0C
#94810000000
1!
1*
b10 6
19
1>
1C
b10 G
#94820000000
0!
0*
09
0>
0C
#94830000000
1!
1*
b11 6
19
1>
1C
b11 G
#94840000000
0!
0*
09
0>
0C
#94850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#94860000000
0!
0*
09
0>
0C
#94870000000
1!
1*
b101 6
19
1>
1C
b101 G
#94880000000
0!
0*
09
0>
0C
#94890000000
1!
1*
b110 6
19
1>
1C
b110 G
#94900000000
0!
0*
09
0>
0C
#94910000000
1!
1*
b111 6
19
1>
1C
b111 G
#94920000000
0!
0*
09
0>
0C
#94930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#94940000000
0!
0*
09
0>
0C
#94950000000
1!
1*
b1 6
19
1>
1C
b1 G
#94960000000
0!
0*
09
0>
0C
#94970000000
1!
1*
b10 6
19
1>
1C
b10 G
#94980000000
0!
0*
09
0>
0C
#94990000000
1!
1*
b11 6
19
1>
1C
b11 G
#95000000000
0!
0*
09
0>
0C
#95010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#95020000000
0!
0*
09
0>
0C
#95030000000
1!
1*
b101 6
19
1>
1C
b101 G
#95040000000
0!
0*
09
0>
0C
#95050000000
1!
1*
b110 6
19
1>
1C
b110 G
#95060000000
0!
0*
09
0>
0C
#95070000000
1!
1*
b111 6
19
1>
1C
b111 G
#95080000000
0!
0*
09
0>
0C
#95090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#95100000000
0!
0*
09
0>
0C
#95110000000
1!
1*
b1 6
19
1>
1C
b1 G
#95120000000
0!
0*
09
0>
0C
#95130000000
1!
1*
b10 6
19
1>
1C
b10 G
#95140000000
0!
0*
09
0>
0C
#95150000000
1!
1*
b11 6
19
1>
1C
b11 G
#95160000000
0!
0*
09
0>
0C
#95170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#95180000000
0!
0*
09
0>
0C
#95190000000
1!
1*
b101 6
19
1>
1C
b101 G
#95200000000
0!
0*
09
0>
0C
#95210000000
1!
1*
b110 6
19
1>
1C
b110 G
#95220000000
0!
0*
09
0>
0C
#95230000000
1!
1*
b111 6
19
1>
1C
b111 G
#95240000000
0!
1"
0*
1+
09
1:
0>
0C
#95250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#95260000000
0!
0*
09
0>
0C
#95270000000
1!
1*
b1 6
19
1>
1C
b1 G
#95280000000
0!
0*
09
0>
0C
#95290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#95300000000
0!
0*
09
0>
0C
#95310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#95320000000
0!
0*
09
0>
0C
#95330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#95340000000
0!
0*
09
0>
0C
#95350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#95360000000
0!
0#
0*
0,
09
0>
0?
0C
#95370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#95380000000
0!
0*
09
0>
0C
#95390000000
1!
1*
19
1>
1C
#95400000000
0!
0*
09
0>
0C
#95410000000
1!
1*
19
1>
1C
#95420000000
0!
0*
09
0>
0C
#95430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#95440000000
0!
0*
09
0>
0C
#95450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#95460000000
0!
0*
09
0>
0C
#95470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#95480000000
0!
0*
09
0>
0C
#95490000000
1!
1*
b10 6
19
1>
1C
b10 G
#95500000000
0!
0*
09
0>
0C
#95510000000
1!
1*
b11 6
19
1>
1C
b11 G
#95520000000
0!
0*
09
0>
0C
#95530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#95540000000
0!
0*
09
0>
0C
#95550000000
1!
1*
b101 6
19
1>
1C
b101 G
#95560000000
0!
0*
09
0>
0C
#95570000000
1!
1*
b110 6
19
1>
1C
b110 G
#95580000000
0!
0*
09
0>
0C
#95590000000
1!
1*
b111 6
19
1>
1C
b111 G
#95600000000
0!
0*
09
0>
0C
#95610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#95620000000
0!
0*
09
0>
0C
#95630000000
1!
1*
b1 6
19
1>
1C
b1 G
#95640000000
0!
0*
09
0>
0C
#95650000000
1!
1*
b10 6
19
1>
1C
b10 G
#95660000000
0!
0*
09
0>
0C
#95670000000
1!
1*
b11 6
19
1>
1C
b11 G
#95680000000
0!
0*
09
0>
0C
#95690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#95700000000
0!
0*
09
0>
0C
#95710000000
1!
1*
b101 6
19
1>
1C
b101 G
#95720000000
0!
0*
09
0>
0C
#95730000000
1!
1*
b110 6
19
1>
1C
b110 G
#95740000000
0!
0*
09
0>
0C
#95750000000
1!
1*
b111 6
19
1>
1C
b111 G
#95760000000
0!
0*
09
0>
0C
#95770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#95780000000
0!
0*
09
0>
0C
#95790000000
1!
1*
b1 6
19
1>
1C
b1 G
#95800000000
0!
0*
09
0>
0C
#95810000000
1!
1*
b10 6
19
1>
1C
b10 G
#95820000000
0!
0*
09
0>
0C
#95830000000
1!
1*
b11 6
19
1>
1C
b11 G
#95840000000
0!
0*
09
0>
0C
#95850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#95860000000
0!
0*
09
0>
0C
#95870000000
1!
1*
b101 6
19
1>
1C
b101 G
#95880000000
0!
0*
09
0>
0C
#95890000000
1!
1*
b110 6
19
1>
1C
b110 G
#95900000000
0!
0*
09
0>
0C
#95910000000
1!
1*
b111 6
19
1>
1C
b111 G
#95920000000
0!
1"
0*
1+
09
1:
0>
0C
#95930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#95940000000
0!
0*
09
0>
0C
#95950000000
1!
1*
b1 6
19
1>
1C
b1 G
#95960000000
0!
0*
09
0>
0C
#95970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#95980000000
0!
0*
09
0>
0C
#95990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#96000000000
0!
0*
09
0>
0C
#96010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#96020000000
0!
0*
09
0>
0C
#96030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#96040000000
0!
0#
0*
0,
09
0>
0?
0C
#96050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#96060000000
0!
0*
09
0>
0C
#96070000000
1!
1*
19
1>
1C
#96080000000
0!
0*
09
0>
0C
#96090000000
1!
1*
19
1>
1C
#96100000000
0!
0*
09
0>
0C
#96110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#96120000000
0!
0*
09
0>
0C
#96130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#96140000000
0!
0*
09
0>
0C
#96150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#96160000000
0!
0*
09
0>
0C
#96170000000
1!
1*
b10 6
19
1>
1C
b10 G
#96180000000
0!
0*
09
0>
0C
#96190000000
1!
1*
b11 6
19
1>
1C
b11 G
#96200000000
0!
0*
09
0>
0C
#96210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#96220000000
0!
0*
09
0>
0C
#96230000000
1!
1*
b101 6
19
1>
1C
b101 G
#96240000000
0!
0*
09
0>
0C
#96250000000
1!
1*
b110 6
19
1>
1C
b110 G
#96260000000
0!
0*
09
0>
0C
#96270000000
1!
1*
b111 6
19
1>
1C
b111 G
#96280000000
0!
0*
09
0>
0C
#96290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#96300000000
0!
0*
09
0>
0C
#96310000000
1!
1*
b1 6
19
1>
1C
b1 G
#96320000000
0!
0*
09
0>
0C
#96330000000
1!
1*
b10 6
19
1>
1C
b10 G
#96340000000
0!
0*
09
0>
0C
#96350000000
1!
1*
b11 6
19
1>
1C
b11 G
#96360000000
0!
0*
09
0>
0C
#96370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#96380000000
0!
0*
09
0>
0C
#96390000000
1!
1*
b101 6
19
1>
1C
b101 G
#96400000000
0!
0*
09
0>
0C
#96410000000
1!
1*
b110 6
19
1>
1C
b110 G
#96420000000
0!
0*
09
0>
0C
#96430000000
1!
1*
b111 6
19
1>
1C
b111 G
#96440000000
0!
0*
09
0>
0C
#96450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#96460000000
0!
0*
09
0>
0C
#96470000000
1!
1*
b1 6
19
1>
1C
b1 G
#96480000000
0!
0*
09
0>
0C
#96490000000
1!
1*
b10 6
19
1>
1C
b10 G
#96500000000
0!
0*
09
0>
0C
#96510000000
1!
1*
b11 6
19
1>
1C
b11 G
#96520000000
0!
0*
09
0>
0C
#96530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#96540000000
0!
0*
09
0>
0C
#96550000000
1!
1*
b101 6
19
1>
1C
b101 G
#96560000000
0!
0*
09
0>
0C
#96570000000
1!
1*
b110 6
19
1>
1C
b110 G
#96580000000
0!
0*
09
0>
0C
#96590000000
1!
1*
b111 6
19
1>
1C
b111 G
#96600000000
0!
1"
0*
1+
09
1:
0>
0C
#96610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#96620000000
0!
0*
09
0>
0C
#96630000000
1!
1*
b1 6
19
1>
1C
b1 G
#96640000000
0!
0*
09
0>
0C
#96650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#96660000000
0!
0*
09
0>
0C
#96670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#96680000000
0!
0*
09
0>
0C
#96690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#96700000000
0!
0*
09
0>
0C
#96710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#96720000000
0!
0#
0*
0,
09
0>
0?
0C
#96730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#96740000000
0!
0*
09
0>
0C
#96750000000
1!
1*
19
1>
1C
#96760000000
0!
0*
09
0>
0C
#96770000000
1!
1*
19
1>
1C
#96780000000
0!
0*
09
0>
0C
#96790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#96800000000
0!
0*
09
0>
0C
#96810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#96820000000
0!
0*
09
0>
0C
#96830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#96840000000
0!
0*
09
0>
0C
#96850000000
1!
1*
b10 6
19
1>
1C
b10 G
#96860000000
0!
0*
09
0>
0C
#96870000000
1!
1*
b11 6
19
1>
1C
b11 G
#96880000000
0!
0*
09
0>
0C
#96890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#96900000000
0!
0*
09
0>
0C
#96910000000
1!
1*
b101 6
19
1>
1C
b101 G
#96920000000
0!
0*
09
0>
0C
#96930000000
1!
1*
b110 6
19
1>
1C
b110 G
#96940000000
0!
0*
09
0>
0C
#96950000000
1!
1*
b111 6
19
1>
1C
b111 G
#96960000000
0!
0*
09
0>
0C
#96970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#96980000000
0!
0*
09
0>
0C
#96990000000
1!
1*
b1 6
19
1>
1C
b1 G
#97000000000
0!
0*
09
0>
0C
#97010000000
1!
1*
b10 6
19
1>
1C
b10 G
#97020000000
0!
0*
09
0>
0C
#97030000000
1!
1*
b11 6
19
1>
1C
b11 G
#97040000000
0!
0*
09
0>
0C
#97050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#97060000000
0!
0*
09
0>
0C
#97070000000
1!
1*
b101 6
19
1>
1C
b101 G
#97080000000
0!
0*
09
0>
0C
#97090000000
1!
1*
b110 6
19
1>
1C
b110 G
#97100000000
0!
0*
09
0>
0C
#97110000000
1!
1*
b111 6
19
1>
1C
b111 G
#97120000000
0!
0*
09
0>
0C
#97130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#97140000000
0!
0*
09
0>
0C
#97150000000
1!
1*
b1 6
19
1>
1C
b1 G
#97160000000
0!
0*
09
0>
0C
#97170000000
1!
1*
b10 6
19
1>
1C
b10 G
#97180000000
0!
0*
09
0>
0C
#97190000000
1!
1*
b11 6
19
1>
1C
b11 G
#97200000000
0!
0*
09
0>
0C
#97210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#97220000000
0!
0*
09
0>
0C
#97230000000
1!
1*
b101 6
19
1>
1C
b101 G
#97240000000
0!
0*
09
0>
0C
#97250000000
1!
1*
b110 6
19
1>
1C
b110 G
#97260000000
0!
0*
09
0>
0C
#97270000000
1!
1*
b111 6
19
1>
1C
b111 G
#97280000000
0!
1"
0*
1+
09
1:
0>
0C
#97290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#97300000000
0!
0*
09
0>
0C
#97310000000
1!
1*
b1 6
19
1>
1C
b1 G
#97320000000
0!
0*
09
0>
0C
#97330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#97340000000
0!
0*
09
0>
0C
#97350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#97360000000
0!
0*
09
0>
0C
#97370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#97380000000
0!
0*
09
0>
0C
#97390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#97400000000
0!
0#
0*
0,
09
0>
0?
0C
#97410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#97420000000
0!
0*
09
0>
0C
#97430000000
1!
1*
19
1>
1C
#97440000000
0!
0*
09
0>
0C
#97450000000
1!
1*
19
1>
1C
#97460000000
0!
0*
09
0>
0C
#97470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#97480000000
0!
0*
09
0>
0C
#97490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#97500000000
0!
0*
09
0>
0C
#97510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#97520000000
0!
0*
09
0>
0C
#97530000000
1!
1*
b10 6
19
1>
1C
b10 G
#97540000000
0!
0*
09
0>
0C
#97550000000
1!
1*
b11 6
19
1>
1C
b11 G
#97560000000
0!
0*
09
0>
0C
#97570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#97580000000
0!
0*
09
0>
0C
#97590000000
1!
1*
b101 6
19
1>
1C
b101 G
#97600000000
0!
0*
09
0>
0C
#97610000000
1!
1*
b110 6
19
1>
1C
b110 G
#97620000000
0!
0*
09
0>
0C
#97630000000
1!
1*
b111 6
19
1>
1C
b111 G
#97640000000
0!
0*
09
0>
0C
#97650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#97660000000
0!
0*
09
0>
0C
#97670000000
1!
1*
b1 6
19
1>
1C
b1 G
#97680000000
0!
0*
09
0>
0C
#97690000000
1!
1*
b10 6
19
1>
1C
b10 G
#97700000000
0!
0*
09
0>
0C
#97710000000
1!
1*
b11 6
19
1>
1C
b11 G
#97720000000
0!
0*
09
0>
0C
#97730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#97740000000
0!
0*
09
0>
0C
#97750000000
1!
1*
b101 6
19
1>
1C
b101 G
#97760000000
0!
0*
09
0>
0C
#97770000000
1!
1*
b110 6
19
1>
1C
b110 G
#97780000000
0!
0*
09
0>
0C
#97790000000
1!
1*
b111 6
19
1>
1C
b111 G
#97800000000
0!
0*
09
0>
0C
#97810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#97820000000
0!
0*
09
0>
0C
#97830000000
1!
1*
b1 6
19
1>
1C
b1 G
#97840000000
0!
0*
09
0>
0C
#97850000000
1!
1*
b10 6
19
1>
1C
b10 G
#97860000000
0!
0*
09
0>
0C
#97870000000
1!
1*
b11 6
19
1>
1C
b11 G
#97880000000
0!
0*
09
0>
0C
#97890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#97900000000
0!
0*
09
0>
0C
#97910000000
1!
1*
b101 6
19
1>
1C
b101 G
#97920000000
0!
0*
09
0>
0C
#97930000000
1!
1*
b110 6
19
1>
1C
b110 G
#97940000000
0!
0*
09
0>
0C
#97950000000
1!
1*
b111 6
19
1>
1C
b111 G
#97960000000
0!
1"
0*
1+
09
1:
0>
0C
#97970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#97980000000
0!
0*
09
0>
0C
#97990000000
1!
1*
b1 6
19
1>
1C
b1 G
#98000000000
0!
0*
09
0>
0C
#98010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#98020000000
0!
0*
09
0>
0C
#98030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#98040000000
0!
0*
09
0>
0C
#98050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#98060000000
0!
0*
09
0>
0C
#98070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#98080000000
0!
0#
0*
0,
09
0>
0?
0C
#98090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#98100000000
0!
0*
09
0>
0C
#98110000000
1!
1*
19
1>
1C
#98120000000
0!
0*
09
0>
0C
#98130000000
1!
1*
19
1>
1C
#98140000000
0!
0*
09
0>
0C
#98150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#98160000000
0!
0*
09
0>
0C
#98170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#98180000000
0!
0*
09
0>
0C
#98190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#98200000000
0!
0*
09
0>
0C
#98210000000
1!
1*
b10 6
19
1>
1C
b10 G
#98220000000
0!
0*
09
0>
0C
#98230000000
1!
1*
b11 6
19
1>
1C
b11 G
#98240000000
0!
0*
09
0>
0C
#98250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#98260000000
0!
0*
09
0>
0C
#98270000000
1!
1*
b101 6
19
1>
1C
b101 G
#98280000000
0!
0*
09
0>
0C
#98290000000
1!
1*
b110 6
19
1>
1C
b110 G
#98300000000
0!
0*
09
0>
0C
#98310000000
1!
1*
b111 6
19
1>
1C
b111 G
#98320000000
0!
0*
09
0>
0C
#98330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#98340000000
0!
0*
09
0>
0C
#98350000000
1!
1*
b1 6
19
1>
1C
b1 G
#98360000000
0!
0*
09
0>
0C
#98370000000
1!
1*
b10 6
19
1>
1C
b10 G
#98380000000
0!
0*
09
0>
0C
#98390000000
1!
1*
b11 6
19
1>
1C
b11 G
#98400000000
0!
0*
09
0>
0C
#98410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#98420000000
0!
0*
09
0>
0C
#98430000000
1!
1*
b101 6
19
1>
1C
b101 G
#98440000000
0!
0*
09
0>
0C
#98450000000
1!
1*
b110 6
19
1>
1C
b110 G
#98460000000
0!
0*
09
0>
0C
#98470000000
1!
1*
b111 6
19
1>
1C
b111 G
#98480000000
0!
0*
09
0>
0C
#98490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#98500000000
0!
0*
09
0>
0C
#98510000000
1!
1*
b1 6
19
1>
1C
b1 G
#98520000000
0!
0*
09
0>
0C
#98530000000
1!
1*
b10 6
19
1>
1C
b10 G
#98540000000
0!
0*
09
0>
0C
#98550000000
1!
1*
b11 6
19
1>
1C
b11 G
#98560000000
0!
0*
09
0>
0C
#98570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#98580000000
0!
0*
09
0>
0C
#98590000000
1!
1*
b101 6
19
1>
1C
b101 G
#98600000000
0!
0*
09
0>
0C
#98610000000
1!
1*
b110 6
19
1>
1C
b110 G
#98620000000
0!
0*
09
0>
0C
#98630000000
1!
1*
b111 6
19
1>
1C
b111 G
#98640000000
0!
1"
0*
1+
09
1:
0>
0C
#98650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#98660000000
0!
0*
09
0>
0C
#98670000000
1!
1*
b1 6
19
1>
1C
b1 G
#98680000000
0!
0*
09
0>
0C
#98690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#98700000000
0!
0*
09
0>
0C
#98710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#98720000000
0!
0*
09
0>
0C
#98730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#98740000000
0!
0*
09
0>
0C
#98750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#98760000000
0!
0#
0*
0,
09
0>
0?
0C
#98770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#98780000000
0!
0*
09
0>
0C
#98790000000
1!
1*
19
1>
1C
#98800000000
0!
0*
09
0>
0C
#98810000000
1!
1*
19
1>
1C
#98820000000
0!
0*
09
0>
0C
#98830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#98840000000
0!
0*
09
0>
0C
#98850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#98860000000
0!
0*
09
0>
0C
#98870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#98880000000
0!
0*
09
0>
0C
#98890000000
1!
1*
b10 6
19
1>
1C
b10 G
#98900000000
0!
0*
09
0>
0C
#98910000000
1!
1*
b11 6
19
1>
1C
b11 G
#98920000000
0!
0*
09
0>
0C
#98930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#98940000000
0!
0*
09
0>
0C
#98950000000
1!
1*
b101 6
19
1>
1C
b101 G
#98960000000
0!
0*
09
0>
0C
#98970000000
1!
1*
b110 6
19
1>
1C
b110 G
#98980000000
0!
0*
09
0>
0C
#98990000000
1!
1*
b111 6
19
1>
1C
b111 G
#99000000000
0!
0*
09
0>
0C
#99010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#99020000000
0!
0*
09
0>
0C
#99030000000
1!
1*
b1 6
19
1>
1C
b1 G
#99040000000
0!
0*
09
0>
0C
#99050000000
1!
1*
b10 6
19
1>
1C
b10 G
#99060000000
0!
0*
09
0>
0C
#99070000000
1!
1*
b11 6
19
1>
1C
b11 G
#99080000000
0!
0*
09
0>
0C
#99090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#99100000000
0!
0*
09
0>
0C
#99110000000
1!
1*
b101 6
19
1>
1C
b101 G
#99120000000
0!
0*
09
0>
0C
#99130000000
1!
1*
b110 6
19
1>
1C
b110 G
#99140000000
0!
0*
09
0>
0C
#99150000000
1!
1*
b111 6
19
1>
1C
b111 G
#99160000000
0!
0*
09
0>
0C
#99170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#99180000000
0!
0*
09
0>
0C
#99190000000
1!
1*
b1 6
19
1>
1C
b1 G
#99200000000
0!
0*
09
0>
0C
#99210000000
1!
1*
b10 6
19
1>
1C
b10 G
#99220000000
0!
0*
09
0>
0C
#99230000000
1!
1*
b11 6
19
1>
1C
b11 G
#99240000000
0!
0*
09
0>
0C
#99250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#99260000000
0!
0*
09
0>
0C
#99270000000
1!
1*
b101 6
19
1>
1C
b101 G
#99280000000
0!
0*
09
0>
0C
#99290000000
1!
1*
b110 6
19
1>
1C
b110 G
#99300000000
0!
0*
09
0>
0C
#99310000000
1!
1*
b111 6
19
1>
1C
b111 G
#99320000000
0!
1"
0*
1+
09
1:
0>
0C
#99330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#99340000000
0!
0*
09
0>
0C
#99350000000
1!
1*
b1 6
19
1>
1C
b1 G
#99360000000
0!
0*
09
0>
0C
#99370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#99380000000
0!
0*
09
0>
0C
#99390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#99400000000
0!
0*
09
0>
0C
#99410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#99420000000
0!
0*
09
0>
0C
#99430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#99440000000
0!
0#
0*
0,
09
0>
0?
0C
#99450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#99460000000
0!
0*
09
0>
0C
#99470000000
1!
1*
19
1>
1C
#99480000000
0!
0*
09
0>
0C
#99490000000
1!
1*
19
1>
1C
#99500000000
0!
0*
09
0>
0C
#99510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#99520000000
0!
0*
09
0>
0C
#99530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#99540000000
0!
0*
09
0>
0C
#99550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#99560000000
0!
0*
09
0>
0C
#99570000000
1!
1*
b10 6
19
1>
1C
b10 G
#99580000000
0!
0*
09
0>
0C
#99590000000
1!
1*
b11 6
19
1>
1C
b11 G
#99600000000
0!
0*
09
0>
0C
#99610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#99620000000
0!
0*
09
0>
0C
#99630000000
1!
1*
b101 6
19
1>
1C
b101 G
#99640000000
0!
0*
09
0>
0C
#99650000000
1!
1*
b110 6
19
1>
1C
b110 G
#99660000000
0!
0*
09
0>
0C
#99670000000
1!
1*
b111 6
19
1>
1C
b111 G
#99680000000
0!
0*
09
0>
0C
#99690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#99700000000
0!
0*
09
0>
0C
#99710000000
1!
1*
b1 6
19
1>
1C
b1 G
#99720000000
0!
0*
09
0>
0C
#99730000000
1!
1*
b10 6
19
1>
1C
b10 G
#99740000000
0!
0*
09
0>
0C
#99750000000
1!
1*
b11 6
19
1>
1C
b11 G
#99760000000
0!
0*
09
0>
0C
#99770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#99780000000
0!
0*
09
0>
0C
#99790000000
1!
1*
b101 6
19
1>
1C
b101 G
#99800000000
0!
0*
09
0>
0C
#99810000000
1!
1*
b110 6
19
1>
1C
b110 G
#99820000000
0!
0*
09
0>
0C
#99830000000
1!
1*
b111 6
19
1>
1C
b111 G
#99840000000
0!
0*
09
0>
0C
#99850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#99860000000
0!
0*
09
0>
0C
#99870000000
1!
1*
b1 6
19
1>
1C
b1 G
#99880000000
0!
0*
09
0>
0C
#99890000000
1!
1*
b10 6
19
1>
1C
b10 G
#99900000000
0!
0*
09
0>
0C
#99910000000
1!
1*
b11 6
19
1>
1C
b11 G
#99920000000
0!
0*
09
0>
0C
#99930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#99940000000
0!
0*
09
0>
0C
#99950000000
1!
1*
b101 6
19
1>
1C
b101 G
#99960000000
0!
0*
09
0>
0C
#99970000000
1!
1*
b110 6
19
1>
1C
b110 G
#99980000000
0!
0*
09
0>
0C
#99990000000
1!
1*
b111 6
19
1>
1C
b111 G
#100000000000
0!
1"
0*
1+
09
1:
0>
0C
#100010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#100020000000
0!
0*
09
0>
0C
#100030000000
1!
1*
b1 6
19
1>
1C
b1 G
#100040000000
0!
0*
09
0>
0C
#100050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#100060000000
0!
0*
09
0>
0C
#100070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#100080000000
0!
0*
09
0>
0C
#100090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#100100000000
0!
0*
09
0>
0C
#100110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#100120000000
0!
0#
0*
0,
09
0>
0?
0C
#100130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#100140000000
0!
0*
09
0>
0C
#100150000000
1!
1*
19
1>
1C
#100160000000
0!
0*
09
0>
0C
#100170000000
1!
1*
19
1>
1C
#100180000000
0!
0*
09
0>
0C
#100190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#100200000000
0!
0*
09
0>
0C
#100210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#100220000000
0!
0*
09
0>
0C
#100230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#100240000000
0!
0*
09
0>
0C
#100250000000
1!
1*
b10 6
19
1>
1C
b10 G
#100260000000
0!
0*
09
0>
0C
#100270000000
1!
1*
b11 6
19
1>
1C
b11 G
#100280000000
0!
0*
09
0>
0C
#100290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#100300000000
0!
0*
09
0>
0C
#100310000000
1!
1*
b101 6
19
1>
1C
b101 G
#100320000000
0!
0*
09
0>
0C
#100330000000
1!
1*
b110 6
19
1>
1C
b110 G
#100340000000
0!
0*
09
0>
0C
#100350000000
1!
1*
b111 6
19
1>
1C
b111 G
#100360000000
0!
0*
09
0>
0C
#100370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#100380000000
0!
0*
09
0>
0C
#100390000000
1!
1*
b1 6
19
1>
1C
b1 G
#100400000000
0!
0*
09
0>
0C
#100410000000
1!
1*
b10 6
19
1>
1C
b10 G
#100420000000
0!
0*
09
0>
0C
#100430000000
1!
1*
b11 6
19
1>
1C
b11 G
#100440000000
0!
0*
09
0>
0C
#100450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#100460000000
0!
0*
09
0>
0C
#100470000000
1!
1*
b101 6
19
1>
1C
b101 G
#100480000000
0!
0*
09
0>
0C
#100490000000
1!
1*
b110 6
19
1>
1C
b110 G
#100500000000
0!
0*
09
0>
0C
#100510000000
1!
1*
b111 6
19
1>
1C
b111 G
#100520000000
0!
0*
09
0>
0C
#100530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#100540000000
0!
0*
09
0>
0C
#100550000000
1!
1*
b1 6
19
1>
1C
b1 G
#100560000000
0!
0*
09
0>
0C
#100570000000
1!
1*
b10 6
19
1>
1C
b10 G
#100580000000
0!
0*
09
0>
0C
#100590000000
1!
1*
b11 6
19
1>
1C
b11 G
#100600000000
0!
0*
09
0>
0C
#100610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#100620000000
0!
0*
09
0>
0C
#100630000000
1!
1*
b101 6
19
1>
1C
b101 G
#100640000000
0!
0*
09
0>
0C
#100650000000
1!
1*
b110 6
19
1>
1C
b110 G
#100660000000
0!
0*
09
0>
0C
#100670000000
1!
1*
b111 6
19
1>
1C
b111 G
#100680000000
0!
1"
0*
1+
09
1:
0>
0C
#100690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#100700000000
0!
0*
09
0>
0C
#100710000000
1!
1*
b1 6
19
1>
1C
b1 G
#100720000000
0!
0*
09
0>
0C
#100730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#100740000000
0!
0*
09
0>
0C
#100750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#100760000000
0!
0*
09
0>
0C
#100770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#100780000000
0!
0*
09
0>
0C
#100790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#100800000000
0!
0#
0*
0,
09
0>
0?
0C
#100810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#100820000000
0!
0*
09
0>
0C
#100830000000
1!
1*
19
1>
1C
#100840000000
0!
0*
09
0>
0C
#100850000000
1!
1*
19
1>
1C
#100860000000
0!
0*
09
0>
0C
#100870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#100880000000
0!
0*
09
0>
0C
#100890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#100900000000
0!
0*
09
0>
0C
#100910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#100920000000
0!
0*
09
0>
0C
#100930000000
1!
1*
b10 6
19
1>
1C
b10 G
#100940000000
0!
0*
09
0>
0C
#100950000000
1!
1*
b11 6
19
1>
1C
b11 G
#100960000000
0!
0*
09
0>
0C
#100970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#100980000000
0!
0*
09
0>
0C
#100990000000
1!
1*
b101 6
19
1>
1C
b101 G
#101000000000
0!
0*
09
0>
0C
#101010000000
1!
1*
b110 6
19
1>
1C
b110 G
#101020000000
0!
0*
09
0>
0C
#101030000000
1!
1*
b111 6
19
1>
1C
b111 G
#101040000000
0!
0*
09
0>
0C
#101050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#101060000000
0!
0*
09
0>
0C
#101070000000
1!
1*
b1 6
19
1>
1C
b1 G
#101080000000
0!
0*
09
0>
0C
#101090000000
1!
1*
b10 6
19
1>
1C
b10 G
#101100000000
0!
0*
09
0>
0C
#101110000000
1!
1*
b11 6
19
1>
1C
b11 G
#101120000000
0!
0*
09
0>
0C
#101130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#101140000000
0!
0*
09
0>
0C
#101150000000
1!
1*
b101 6
19
1>
1C
b101 G
#101160000000
0!
0*
09
0>
0C
#101170000000
1!
1*
b110 6
19
1>
1C
b110 G
#101180000000
0!
0*
09
0>
0C
#101190000000
1!
1*
b111 6
19
1>
1C
b111 G
#101200000000
0!
0*
09
0>
0C
#101210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#101220000000
0!
0*
09
0>
0C
#101230000000
1!
1*
b1 6
19
1>
1C
b1 G
#101240000000
0!
0*
09
0>
0C
#101250000000
1!
1*
b10 6
19
1>
1C
b10 G
#101260000000
0!
0*
09
0>
0C
#101270000000
1!
1*
b11 6
19
1>
1C
b11 G
#101280000000
0!
0*
09
0>
0C
#101290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#101300000000
0!
0*
09
0>
0C
#101310000000
1!
1*
b101 6
19
1>
1C
b101 G
#101320000000
0!
0*
09
0>
0C
#101330000000
1!
1*
b110 6
19
1>
1C
b110 G
#101340000000
0!
0*
09
0>
0C
#101350000000
1!
1*
b111 6
19
1>
1C
b111 G
#101360000000
0!
1"
0*
1+
09
1:
0>
0C
#101370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#101380000000
0!
0*
09
0>
0C
#101390000000
1!
1*
b1 6
19
1>
1C
b1 G
#101400000000
0!
0*
09
0>
0C
#101410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#101420000000
0!
0*
09
0>
0C
#101430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#101440000000
0!
0*
09
0>
0C
#101450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#101460000000
0!
0*
09
0>
0C
#101470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#101480000000
0!
0#
0*
0,
09
0>
0?
0C
#101490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#101500000000
0!
0*
09
0>
0C
#101510000000
1!
1*
19
1>
1C
#101520000000
0!
0*
09
0>
0C
#101530000000
1!
1*
19
1>
1C
#101540000000
0!
0*
09
0>
0C
#101550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#101560000000
0!
0*
09
0>
0C
#101570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#101580000000
0!
0*
09
0>
0C
#101590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#101600000000
0!
0*
09
0>
0C
#101610000000
1!
1*
b10 6
19
1>
1C
b10 G
#101620000000
0!
0*
09
0>
0C
#101630000000
1!
1*
b11 6
19
1>
1C
b11 G
#101640000000
0!
0*
09
0>
0C
#101650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#101660000000
0!
0*
09
0>
0C
#101670000000
1!
1*
b101 6
19
1>
1C
b101 G
#101680000000
0!
0*
09
0>
0C
#101690000000
1!
1*
b110 6
19
1>
1C
b110 G
#101700000000
0!
0*
09
0>
0C
#101710000000
1!
1*
b111 6
19
1>
1C
b111 G
#101720000000
0!
0*
09
0>
0C
#101730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#101740000000
0!
0*
09
0>
0C
#101750000000
1!
1*
b1 6
19
1>
1C
b1 G
#101760000000
0!
0*
09
0>
0C
#101770000000
1!
1*
b10 6
19
1>
1C
b10 G
#101780000000
0!
0*
09
0>
0C
#101790000000
1!
1*
b11 6
19
1>
1C
b11 G
#101800000000
0!
0*
09
0>
0C
#101810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#101820000000
0!
0*
09
0>
0C
#101830000000
1!
1*
b101 6
19
1>
1C
b101 G
#101840000000
0!
0*
09
0>
0C
#101850000000
1!
1*
b110 6
19
1>
1C
b110 G
#101860000000
0!
0*
09
0>
0C
#101870000000
1!
1*
b111 6
19
1>
1C
b111 G
#101880000000
0!
0*
09
0>
0C
#101890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#101900000000
0!
0*
09
0>
0C
#101910000000
1!
1*
b1 6
19
1>
1C
b1 G
#101920000000
0!
0*
09
0>
0C
#101930000000
1!
1*
b10 6
19
1>
1C
b10 G
#101940000000
0!
0*
09
0>
0C
#101950000000
1!
1*
b11 6
19
1>
1C
b11 G
#101960000000
0!
0*
09
0>
0C
#101970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#101980000000
0!
0*
09
0>
0C
#101990000000
1!
1*
b101 6
19
1>
1C
b101 G
#102000000000
0!
0*
09
0>
0C
#102010000000
1!
1*
b110 6
19
1>
1C
b110 G
#102020000000
0!
0*
09
0>
0C
#102030000000
1!
1*
b111 6
19
1>
1C
b111 G
#102040000000
0!
1"
0*
1+
09
1:
0>
0C
#102050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#102060000000
0!
0*
09
0>
0C
#102070000000
1!
1*
b1 6
19
1>
1C
b1 G
#102080000000
0!
0*
09
0>
0C
#102090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#102100000000
0!
0*
09
0>
0C
#102110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#102120000000
0!
0*
09
0>
0C
#102130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#102140000000
0!
0*
09
0>
0C
#102150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#102160000000
0!
0#
0*
0,
09
0>
0?
0C
#102170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#102180000000
0!
0*
09
0>
0C
#102190000000
1!
1*
19
1>
1C
#102200000000
0!
0*
09
0>
0C
#102210000000
1!
1*
19
1>
1C
#102220000000
0!
0*
09
0>
0C
#102230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#102240000000
0!
0*
09
0>
0C
#102250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#102260000000
0!
0*
09
0>
0C
#102270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#102280000000
0!
0*
09
0>
0C
#102290000000
1!
1*
b10 6
19
1>
1C
b10 G
#102300000000
0!
0*
09
0>
0C
#102310000000
1!
1*
b11 6
19
1>
1C
b11 G
#102320000000
0!
0*
09
0>
0C
#102330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#102340000000
0!
0*
09
0>
0C
#102350000000
1!
1*
b101 6
19
1>
1C
b101 G
#102360000000
0!
0*
09
0>
0C
#102370000000
1!
1*
b110 6
19
1>
1C
b110 G
#102380000000
0!
0*
09
0>
0C
#102390000000
1!
1*
b111 6
19
1>
1C
b111 G
#102400000000
0!
0*
09
0>
0C
#102410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#102420000000
0!
0*
09
0>
0C
#102430000000
1!
1*
b1 6
19
1>
1C
b1 G
#102440000000
0!
0*
09
0>
0C
#102450000000
1!
1*
b10 6
19
1>
1C
b10 G
#102460000000
0!
0*
09
0>
0C
#102470000000
1!
1*
b11 6
19
1>
1C
b11 G
#102480000000
0!
0*
09
0>
0C
#102490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#102500000000
0!
0*
09
0>
0C
#102510000000
1!
1*
b101 6
19
1>
1C
b101 G
#102520000000
0!
0*
09
0>
0C
#102530000000
1!
1*
b110 6
19
1>
1C
b110 G
#102540000000
0!
0*
09
0>
0C
#102550000000
1!
1*
b111 6
19
1>
1C
b111 G
#102560000000
0!
0*
09
0>
0C
#102570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#102580000000
0!
0*
09
0>
0C
#102590000000
1!
1*
b1 6
19
1>
1C
b1 G
#102600000000
0!
0*
09
0>
0C
#102610000000
1!
1*
b10 6
19
1>
1C
b10 G
#102620000000
0!
0*
09
0>
0C
#102630000000
1!
1*
b11 6
19
1>
1C
b11 G
#102640000000
0!
0*
09
0>
0C
#102650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#102660000000
0!
0*
09
0>
0C
#102670000000
1!
1*
b101 6
19
1>
1C
b101 G
#102680000000
0!
0*
09
0>
0C
#102690000000
1!
1*
b110 6
19
1>
1C
b110 G
#102700000000
0!
0*
09
0>
0C
#102710000000
1!
1*
b111 6
19
1>
1C
b111 G
#102720000000
0!
1"
0*
1+
09
1:
0>
0C
#102730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#102740000000
0!
0*
09
0>
0C
#102750000000
1!
1*
b1 6
19
1>
1C
b1 G
#102760000000
0!
0*
09
0>
0C
#102770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#102780000000
0!
0*
09
0>
0C
#102790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#102800000000
0!
0*
09
0>
0C
#102810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#102820000000
0!
0*
09
0>
0C
#102830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#102840000000
0!
0#
0*
0,
09
0>
0?
0C
#102850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#102860000000
0!
0*
09
0>
0C
#102870000000
1!
1*
19
1>
1C
#102880000000
0!
0*
09
0>
0C
#102890000000
1!
1*
19
1>
1C
#102900000000
0!
0*
09
0>
0C
#102910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#102920000000
0!
0*
09
0>
0C
#102930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#102940000000
0!
0*
09
0>
0C
#102950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#102960000000
0!
0*
09
0>
0C
#102970000000
1!
1*
b10 6
19
1>
1C
b10 G
#102980000000
0!
0*
09
0>
0C
#102990000000
1!
1*
b11 6
19
1>
1C
b11 G
#103000000000
0!
0*
09
0>
0C
#103010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#103020000000
0!
0*
09
0>
0C
#103030000000
1!
1*
b101 6
19
1>
1C
b101 G
#103040000000
0!
0*
09
0>
0C
#103050000000
1!
1*
b110 6
19
1>
1C
b110 G
#103060000000
0!
0*
09
0>
0C
#103070000000
1!
1*
b111 6
19
1>
1C
b111 G
#103080000000
0!
0*
09
0>
0C
#103090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#103100000000
0!
0*
09
0>
0C
#103110000000
1!
1*
b1 6
19
1>
1C
b1 G
#103120000000
0!
0*
09
0>
0C
#103130000000
1!
1*
b10 6
19
1>
1C
b10 G
#103140000000
0!
0*
09
0>
0C
#103150000000
1!
1*
b11 6
19
1>
1C
b11 G
#103160000000
0!
0*
09
0>
0C
#103170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#103180000000
0!
0*
09
0>
0C
#103190000000
1!
1*
b101 6
19
1>
1C
b101 G
#103200000000
0!
0*
09
0>
0C
#103210000000
1!
1*
b110 6
19
1>
1C
b110 G
#103220000000
0!
0*
09
0>
0C
#103230000000
1!
1*
b111 6
19
1>
1C
b111 G
#103240000000
0!
0*
09
0>
0C
#103250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#103260000000
0!
0*
09
0>
0C
#103270000000
1!
1*
b1 6
19
1>
1C
b1 G
#103280000000
0!
0*
09
0>
0C
#103290000000
1!
1*
b10 6
19
1>
1C
b10 G
#103300000000
0!
0*
09
0>
0C
#103310000000
1!
1*
b11 6
19
1>
1C
b11 G
#103320000000
0!
0*
09
0>
0C
#103330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#103340000000
0!
0*
09
0>
0C
#103350000000
1!
1*
b101 6
19
1>
1C
b101 G
#103360000000
0!
0*
09
0>
0C
#103370000000
1!
1*
b110 6
19
1>
1C
b110 G
#103380000000
0!
0*
09
0>
0C
#103390000000
1!
1*
b111 6
19
1>
1C
b111 G
#103400000000
0!
1"
0*
1+
09
1:
0>
0C
#103410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#103420000000
0!
0*
09
0>
0C
#103430000000
1!
1*
b1 6
19
1>
1C
b1 G
#103440000000
0!
0*
09
0>
0C
#103450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#103460000000
0!
0*
09
0>
0C
#103470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#103480000000
0!
0*
09
0>
0C
#103490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#103500000000
0!
0*
09
0>
0C
#103510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#103520000000
0!
0#
0*
0,
09
0>
0?
0C
#103530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#103540000000
0!
0*
09
0>
0C
#103550000000
1!
1*
19
1>
1C
#103560000000
0!
0*
09
0>
0C
#103570000000
1!
1*
19
1>
1C
#103580000000
0!
0*
09
0>
0C
#103590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#103600000000
0!
0*
09
0>
0C
#103610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#103620000000
0!
0*
09
0>
0C
#103630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#103640000000
0!
0*
09
0>
0C
#103650000000
1!
1*
b10 6
19
1>
1C
b10 G
#103660000000
0!
0*
09
0>
0C
#103670000000
1!
1*
b11 6
19
1>
1C
b11 G
#103680000000
0!
0*
09
0>
0C
#103690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#103700000000
0!
0*
09
0>
0C
#103710000000
1!
1*
b101 6
19
1>
1C
b101 G
#103720000000
0!
0*
09
0>
0C
#103730000000
1!
1*
b110 6
19
1>
1C
b110 G
#103740000000
0!
0*
09
0>
0C
#103750000000
1!
1*
b111 6
19
1>
1C
b111 G
#103760000000
0!
0*
09
0>
0C
#103770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#103780000000
0!
0*
09
0>
0C
#103790000000
1!
1*
b1 6
19
1>
1C
b1 G
#103800000000
0!
0*
09
0>
0C
#103810000000
1!
1*
b10 6
19
1>
1C
b10 G
#103820000000
0!
0*
09
0>
0C
#103830000000
1!
1*
b11 6
19
1>
1C
b11 G
#103840000000
0!
0*
09
0>
0C
#103850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#103860000000
0!
0*
09
0>
0C
#103870000000
1!
1*
b101 6
19
1>
1C
b101 G
#103880000000
0!
0*
09
0>
0C
#103890000000
1!
1*
b110 6
19
1>
1C
b110 G
#103900000000
0!
0*
09
0>
0C
#103910000000
1!
1*
b111 6
19
1>
1C
b111 G
#103920000000
0!
0*
09
0>
0C
#103930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#103940000000
0!
0*
09
0>
0C
#103950000000
1!
1*
b1 6
19
1>
1C
b1 G
#103960000000
0!
0*
09
0>
0C
#103970000000
1!
1*
b10 6
19
1>
1C
b10 G
#103980000000
0!
0*
09
0>
0C
#103990000000
1!
1*
b11 6
19
1>
1C
b11 G
#104000000000
0!
0*
09
0>
0C
#104010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#104020000000
0!
0*
09
0>
0C
#104030000000
1!
1*
b101 6
19
1>
1C
b101 G
#104040000000
0!
0*
09
0>
0C
#104050000000
1!
1*
b110 6
19
1>
1C
b110 G
#104060000000
0!
0*
09
0>
0C
#104070000000
1!
1*
b111 6
19
1>
1C
b111 G
#104080000000
0!
1"
0*
1+
09
1:
0>
0C
#104090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#104100000000
0!
0*
09
0>
0C
#104110000000
1!
1*
b1 6
19
1>
1C
b1 G
#104120000000
0!
0*
09
0>
0C
#104130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#104140000000
0!
0*
09
0>
0C
#104150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#104160000000
0!
0*
09
0>
0C
#104170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#104180000000
0!
0*
09
0>
0C
#104190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#104200000000
0!
0#
0*
0,
09
0>
0?
0C
#104210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#104220000000
0!
0*
09
0>
0C
#104230000000
1!
1*
19
1>
1C
#104240000000
0!
0*
09
0>
0C
#104250000000
1!
1*
19
1>
1C
#104260000000
0!
0*
09
0>
0C
#104270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#104280000000
0!
0*
09
0>
0C
#104290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#104300000000
0!
0*
09
0>
0C
#104310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#104320000000
0!
0*
09
0>
0C
#104330000000
1!
1*
b10 6
19
1>
1C
b10 G
#104340000000
0!
0*
09
0>
0C
#104350000000
1!
1*
b11 6
19
1>
1C
b11 G
#104360000000
0!
0*
09
0>
0C
#104370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#104380000000
0!
0*
09
0>
0C
#104390000000
1!
1*
b101 6
19
1>
1C
b101 G
#104400000000
0!
0*
09
0>
0C
#104410000000
1!
1*
b110 6
19
1>
1C
b110 G
#104420000000
0!
0*
09
0>
0C
#104430000000
1!
1*
b111 6
19
1>
1C
b111 G
#104440000000
0!
0*
09
0>
0C
#104450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#104460000000
0!
0*
09
0>
0C
#104470000000
1!
1*
b1 6
19
1>
1C
b1 G
#104480000000
0!
0*
09
0>
0C
#104490000000
1!
1*
b10 6
19
1>
1C
b10 G
#104500000000
0!
0*
09
0>
0C
#104510000000
1!
1*
b11 6
19
1>
1C
b11 G
#104520000000
0!
0*
09
0>
0C
#104530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#104540000000
0!
0*
09
0>
0C
#104550000000
1!
1*
b101 6
19
1>
1C
b101 G
#104560000000
0!
0*
09
0>
0C
#104570000000
1!
1*
b110 6
19
1>
1C
b110 G
#104580000000
0!
0*
09
0>
0C
#104590000000
1!
1*
b111 6
19
1>
1C
b111 G
#104600000000
0!
0*
09
0>
0C
#104610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#104620000000
0!
0*
09
0>
0C
#104630000000
1!
1*
b1 6
19
1>
1C
b1 G
#104640000000
0!
0*
09
0>
0C
#104650000000
1!
1*
b10 6
19
1>
1C
b10 G
#104660000000
0!
0*
09
0>
0C
#104670000000
1!
1*
b11 6
19
1>
1C
b11 G
#104680000000
0!
0*
09
0>
0C
#104690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#104700000000
0!
0*
09
0>
0C
#104710000000
1!
1*
b101 6
19
1>
1C
b101 G
#104720000000
0!
0*
09
0>
0C
#104730000000
1!
1*
b110 6
19
1>
1C
b110 G
#104740000000
0!
0*
09
0>
0C
#104750000000
1!
1*
b111 6
19
1>
1C
b111 G
#104760000000
0!
1"
0*
1+
09
1:
0>
0C
#104770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#104780000000
0!
0*
09
0>
0C
#104790000000
1!
1*
b1 6
19
1>
1C
b1 G
#104800000000
0!
0*
09
0>
0C
#104810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#104820000000
0!
0*
09
0>
0C
#104830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#104840000000
0!
0*
09
0>
0C
#104850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#104860000000
0!
0*
09
0>
0C
#104870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#104880000000
0!
0#
0*
0,
09
0>
0?
0C
#104890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#104900000000
0!
0*
09
0>
0C
#104910000000
1!
1*
19
1>
1C
#104920000000
0!
0*
09
0>
0C
#104930000000
1!
1*
19
1>
1C
#104940000000
0!
0*
09
0>
0C
#104950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#104960000000
0!
0*
09
0>
0C
#104970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#104980000000
0!
0*
09
0>
0C
#104990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#105000000000
0!
0*
09
0>
0C
#105010000000
1!
1*
b10 6
19
1>
1C
b10 G
#105020000000
0!
0*
09
0>
0C
#105030000000
1!
1*
b11 6
19
1>
1C
b11 G
#105040000000
0!
0*
09
0>
0C
#105050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#105060000000
0!
0*
09
0>
0C
#105070000000
1!
1*
b101 6
19
1>
1C
b101 G
#105080000000
0!
0*
09
0>
0C
#105090000000
1!
1*
b110 6
19
1>
1C
b110 G
#105100000000
0!
0*
09
0>
0C
#105110000000
1!
1*
b111 6
19
1>
1C
b111 G
#105120000000
0!
0*
09
0>
0C
#105130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#105140000000
0!
0*
09
0>
0C
#105150000000
1!
1*
b1 6
19
1>
1C
b1 G
#105160000000
0!
0*
09
0>
0C
#105170000000
1!
1*
b10 6
19
1>
1C
b10 G
#105180000000
0!
0*
09
0>
0C
#105190000000
1!
1*
b11 6
19
1>
1C
b11 G
#105200000000
0!
0*
09
0>
0C
#105210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#105220000000
0!
0*
09
0>
0C
#105230000000
1!
1*
b101 6
19
1>
1C
b101 G
#105240000000
0!
0*
09
0>
0C
#105250000000
1!
1*
b110 6
19
1>
1C
b110 G
#105260000000
0!
0*
09
0>
0C
#105270000000
1!
1*
b111 6
19
1>
1C
b111 G
#105280000000
0!
0*
09
0>
0C
#105290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#105300000000
0!
0*
09
0>
0C
#105310000000
1!
1*
b1 6
19
1>
1C
b1 G
#105320000000
0!
0*
09
0>
0C
#105330000000
1!
1*
b10 6
19
1>
1C
b10 G
#105340000000
0!
0*
09
0>
0C
#105350000000
1!
1*
b11 6
19
1>
1C
b11 G
#105360000000
0!
0*
09
0>
0C
#105370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#105380000000
0!
0*
09
0>
0C
#105390000000
1!
1*
b101 6
19
1>
1C
b101 G
#105400000000
0!
0*
09
0>
0C
#105410000000
1!
1*
b110 6
19
1>
1C
b110 G
#105420000000
0!
0*
09
0>
0C
#105430000000
1!
1*
b111 6
19
1>
1C
b111 G
#105440000000
0!
1"
0*
1+
09
1:
0>
0C
#105450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#105460000000
0!
0*
09
0>
0C
#105470000000
1!
1*
b1 6
19
1>
1C
b1 G
#105480000000
0!
0*
09
0>
0C
#105490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#105500000000
0!
0*
09
0>
0C
#105510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#105520000000
0!
0*
09
0>
0C
#105530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#105540000000
0!
0*
09
0>
0C
#105550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#105560000000
0!
0#
0*
0,
09
0>
0?
0C
#105570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#105580000000
0!
0*
09
0>
0C
#105590000000
1!
1*
19
1>
1C
#105600000000
0!
0*
09
0>
0C
#105610000000
1!
1*
19
1>
1C
#105620000000
0!
0*
09
0>
0C
#105630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#105640000000
0!
0*
09
0>
0C
#105650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#105660000000
0!
0*
09
0>
0C
#105670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#105680000000
0!
0*
09
0>
0C
#105690000000
1!
1*
b10 6
19
1>
1C
b10 G
#105700000000
0!
0*
09
0>
0C
#105710000000
1!
1*
b11 6
19
1>
1C
b11 G
#105720000000
0!
0*
09
0>
0C
#105730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#105740000000
0!
0*
09
0>
0C
#105750000000
1!
1*
b101 6
19
1>
1C
b101 G
#105760000000
0!
0*
09
0>
0C
#105770000000
1!
1*
b110 6
19
1>
1C
b110 G
#105780000000
0!
0*
09
0>
0C
#105790000000
1!
1*
b111 6
19
1>
1C
b111 G
#105800000000
0!
0*
09
0>
0C
#105810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#105820000000
0!
0*
09
0>
0C
#105830000000
1!
1*
b1 6
19
1>
1C
b1 G
#105840000000
0!
0*
09
0>
0C
#105850000000
1!
1*
b10 6
19
1>
1C
b10 G
#105860000000
0!
0*
09
0>
0C
#105870000000
1!
1*
b11 6
19
1>
1C
b11 G
#105880000000
0!
0*
09
0>
0C
#105890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#105900000000
0!
0*
09
0>
0C
#105910000000
1!
1*
b101 6
19
1>
1C
b101 G
#105920000000
0!
0*
09
0>
0C
#105930000000
1!
1*
b110 6
19
1>
1C
b110 G
#105940000000
0!
0*
09
0>
0C
#105950000000
1!
1*
b111 6
19
1>
1C
b111 G
#105960000000
0!
0*
09
0>
0C
#105970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#105980000000
0!
0*
09
0>
0C
#105990000000
1!
1*
b1 6
19
1>
1C
b1 G
#106000000000
0!
0*
09
0>
0C
#106010000000
1!
1*
b10 6
19
1>
1C
b10 G
#106020000000
0!
0*
09
0>
0C
#106030000000
1!
1*
b11 6
19
1>
1C
b11 G
#106040000000
0!
0*
09
0>
0C
#106050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#106060000000
0!
0*
09
0>
0C
#106070000000
1!
1*
b101 6
19
1>
1C
b101 G
#106080000000
0!
0*
09
0>
0C
#106090000000
1!
1*
b110 6
19
1>
1C
b110 G
#106100000000
0!
0*
09
0>
0C
#106110000000
1!
1*
b111 6
19
1>
1C
b111 G
#106120000000
0!
1"
0*
1+
09
1:
0>
0C
#106130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#106140000000
0!
0*
09
0>
0C
#106150000000
1!
1*
b1 6
19
1>
1C
b1 G
#106160000000
0!
0*
09
0>
0C
#106170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#106180000000
0!
0*
09
0>
0C
#106190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#106200000000
0!
0*
09
0>
0C
#106210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#106220000000
0!
0*
09
0>
0C
#106230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#106240000000
0!
0#
0*
0,
09
0>
0?
0C
#106250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#106260000000
0!
0*
09
0>
0C
#106270000000
1!
1*
19
1>
1C
#106280000000
0!
0*
09
0>
0C
#106290000000
1!
1*
19
1>
1C
#106300000000
0!
0*
09
0>
0C
#106310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#106320000000
0!
0*
09
0>
0C
#106330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#106340000000
0!
0*
09
0>
0C
#106350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#106360000000
0!
0*
09
0>
0C
#106370000000
1!
1*
b10 6
19
1>
1C
b10 G
#106380000000
0!
0*
09
0>
0C
#106390000000
1!
1*
b11 6
19
1>
1C
b11 G
#106400000000
0!
0*
09
0>
0C
#106410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#106420000000
0!
0*
09
0>
0C
#106430000000
1!
1*
b101 6
19
1>
1C
b101 G
#106440000000
0!
0*
09
0>
0C
#106450000000
1!
1*
b110 6
19
1>
1C
b110 G
#106460000000
0!
0*
09
0>
0C
#106470000000
1!
1*
b111 6
19
1>
1C
b111 G
#106480000000
0!
0*
09
0>
0C
#106490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#106500000000
0!
0*
09
0>
0C
#106510000000
1!
1*
b1 6
19
1>
1C
b1 G
#106520000000
0!
0*
09
0>
0C
#106530000000
1!
1*
b10 6
19
1>
1C
b10 G
#106540000000
0!
0*
09
0>
0C
#106550000000
1!
1*
b11 6
19
1>
1C
b11 G
#106560000000
0!
0*
09
0>
0C
#106570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#106580000000
0!
0*
09
0>
0C
#106590000000
1!
1*
b101 6
19
1>
1C
b101 G
#106600000000
0!
0*
09
0>
0C
#106610000000
1!
1*
b110 6
19
1>
1C
b110 G
#106620000000
0!
0*
09
0>
0C
#106630000000
1!
1*
b111 6
19
1>
1C
b111 G
#106640000000
0!
0*
09
0>
0C
#106650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#106660000000
0!
0*
09
0>
0C
#106670000000
1!
1*
b1 6
19
1>
1C
b1 G
#106680000000
0!
0*
09
0>
0C
#106690000000
1!
1*
b10 6
19
1>
1C
b10 G
#106700000000
0!
0*
09
0>
0C
#106710000000
1!
1*
b11 6
19
1>
1C
b11 G
#106720000000
0!
0*
09
0>
0C
#106730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#106740000000
0!
0*
09
0>
0C
#106750000000
1!
1*
b101 6
19
1>
1C
b101 G
#106760000000
0!
0*
09
0>
0C
#106770000000
1!
1*
b110 6
19
1>
1C
b110 G
#106780000000
0!
0*
09
0>
0C
#106790000000
1!
1*
b111 6
19
1>
1C
b111 G
#106800000000
0!
1"
0*
1+
09
1:
0>
0C
#106810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#106820000000
0!
0*
09
0>
0C
#106830000000
1!
1*
b1 6
19
1>
1C
b1 G
#106840000000
0!
0*
09
0>
0C
#106850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#106860000000
0!
0*
09
0>
0C
#106870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#106880000000
0!
0*
09
0>
0C
#106890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#106900000000
0!
0*
09
0>
0C
#106910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#106920000000
0!
0#
0*
0,
09
0>
0?
0C
#106930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#106940000000
0!
0*
09
0>
0C
#106950000000
1!
1*
19
1>
1C
#106960000000
0!
0*
09
0>
0C
#106970000000
1!
1*
19
1>
1C
#106980000000
0!
0*
09
0>
0C
#106990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#107000000000
0!
0*
09
0>
0C
#107010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#107020000000
0!
0*
09
0>
0C
#107030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#107040000000
0!
0*
09
0>
0C
#107050000000
1!
1*
b10 6
19
1>
1C
b10 G
#107060000000
0!
0*
09
0>
0C
#107070000000
1!
1*
b11 6
19
1>
1C
b11 G
#107080000000
0!
0*
09
0>
0C
#107090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#107100000000
0!
0*
09
0>
0C
#107110000000
1!
1*
b101 6
19
1>
1C
b101 G
#107120000000
0!
0*
09
0>
0C
#107130000000
1!
1*
b110 6
19
1>
1C
b110 G
#107140000000
0!
0*
09
0>
0C
#107150000000
1!
1*
b111 6
19
1>
1C
b111 G
#107160000000
0!
0*
09
0>
0C
#107170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#107180000000
0!
0*
09
0>
0C
#107190000000
1!
1*
b1 6
19
1>
1C
b1 G
#107200000000
0!
0*
09
0>
0C
#107210000000
1!
1*
b10 6
19
1>
1C
b10 G
#107220000000
0!
0*
09
0>
0C
#107230000000
1!
1*
b11 6
19
1>
1C
b11 G
#107240000000
0!
0*
09
0>
0C
#107250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#107260000000
0!
0*
09
0>
0C
#107270000000
1!
1*
b101 6
19
1>
1C
b101 G
#107280000000
0!
0*
09
0>
0C
#107290000000
1!
1*
b110 6
19
1>
1C
b110 G
#107300000000
0!
0*
09
0>
0C
#107310000000
1!
1*
b111 6
19
1>
1C
b111 G
#107320000000
0!
0*
09
0>
0C
#107330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#107340000000
0!
0*
09
0>
0C
#107350000000
1!
1*
b1 6
19
1>
1C
b1 G
#107360000000
0!
0*
09
0>
0C
#107370000000
1!
1*
b10 6
19
1>
1C
b10 G
#107380000000
0!
0*
09
0>
0C
#107390000000
1!
1*
b11 6
19
1>
1C
b11 G
#107400000000
0!
0*
09
0>
0C
#107410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#107420000000
0!
0*
09
0>
0C
#107430000000
1!
1*
b101 6
19
1>
1C
b101 G
#107440000000
0!
0*
09
0>
0C
#107450000000
1!
1*
b110 6
19
1>
1C
b110 G
#107460000000
0!
0*
09
0>
0C
#107470000000
1!
1*
b111 6
19
1>
1C
b111 G
#107480000000
0!
1"
0*
1+
09
1:
0>
0C
#107490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#107500000000
0!
0*
09
0>
0C
#107510000000
1!
1*
b1 6
19
1>
1C
b1 G
#107520000000
0!
0*
09
0>
0C
#107530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#107540000000
0!
0*
09
0>
0C
#107550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#107560000000
0!
0*
09
0>
0C
#107570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#107580000000
0!
0*
09
0>
0C
#107590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#107600000000
0!
0#
0*
0,
09
0>
0?
0C
#107610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#107620000000
0!
0*
09
0>
0C
#107630000000
1!
1*
19
1>
1C
#107640000000
0!
0*
09
0>
0C
#107650000000
1!
1*
19
1>
1C
#107660000000
0!
0*
09
0>
0C
#107670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#107680000000
0!
0*
09
0>
0C
#107690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#107700000000
0!
0*
09
0>
0C
#107710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#107720000000
0!
0*
09
0>
0C
#107730000000
1!
1*
b10 6
19
1>
1C
b10 G
#107740000000
0!
0*
09
0>
0C
#107750000000
1!
1*
b11 6
19
1>
1C
b11 G
#107760000000
0!
0*
09
0>
0C
#107770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#107780000000
0!
0*
09
0>
0C
#107790000000
1!
1*
b101 6
19
1>
1C
b101 G
#107800000000
0!
0*
09
0>
0C
#107810000000
1!
1*
b110 6
19
1>
1C
b110 G
#107820000000
0!
0*
09
0>
0C
#107830000000
1!
1*
b111 6
19
1>
1C
b111 G
#107840000000
0!
0*
09
0>
0C
#107850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#107860000000
0!
0*
09
0>
0C
#107870000000
1!
1*
b1 6
19
1>
1C
b1 G
#107880000000
0!
0*
09
0>
0C
#107890000000
1!
1*
b10 6
19
1>
1C
b10 G
#107900000000
0!
0*
09
0>
0C
#107910000000
1!
1*
b11 6
19
1>
1C
b11 G
#107920000000
0!
0*
09
0>
0C
#107930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#107940000000
0!
0*
09
0>
0C
#107950000000
1!
1*
b101 6
19
1>
1C
b101 G
#107960000000
0!
0*
09
0>
0C
#107970000000
1!
1*
b110 6
19
1>
1C
b110 G
#107980000000
0!
0*
09
0>
0C
#107990000000
1!
1*
b111 6
19
1>
1C
b111 G
#108000000000
0!
0*
09
0>
0C
#108010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#108020000000
0!
0*
09
0>
0C
#108030000000
1!
1*
b1 6
19
1>
1C
b1 G
#108040000000
0!
0*
09
0>
0C
#108050000000
1!
1*
b10 6
19
1>
1C
b10 G
#108060000000
0!
0*
09
0>
0C
#108070000000
1!
1*
b11 6
19
1>
1C
b11 G
#108080000000
0!
0*
09
0>
0C
#108090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#108100000000
0!
0*
09
0>
0C
#108110000000
1!
1*
b101 6
19
1>
1C
b101 G
#108120000000
0!
0*
09
0>
0C
#108130000000
1!
1*
b110 6
19
1>
1C
b110 G
#108140000000
0!
0*
09
0>
0C
#108150000000
1!
1*
b111 6
19
1>
1C
b111 G
#108160000000
0!
1"
0*
1+
09
1:
0>
0C
#108170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#108180000000
0!
0*
09
0>
0C
#108190000000
1!
1*
b1 6
19
1>
1C
b1 G
#108200000000
0!
0*
09
0>
0C
#108210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#108220000000
0!
0*
09
0>
0C
#108230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#108240000000
0!
0*
09
0>
0C
#108250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#108260000000
0!
0*
09
0>
0C
#108270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#108280000000
0!
0#
0*
0,
09
0>
0?
0C
#108290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#108300000000
0!
0*
09
0>
0C
#108310000000
1!
1*
19
1>
1C
#108320000000
0!
0*
09
0>
0C
#108330000000
1!
1*
19
1>
1C
#108340000000
0!
0*
09
0>
0C
#108350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#108360000000
0!
0*
09
0>
0C
#108370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#108380000000
0!
0*
09
0>
0C
#108390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#108400000000
0!
0*
09
0>
0C
#108410000000
1!
1*
b10 6
19
1>
1C
b10 G
#108420000000
0!
0*
09
0>
0C
#108430000000
1!
1*
b11 6
19
1>
1C
b11 G
#108440000000
0!
0*
09
0>
0C
#108450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#108460000000
0!
0*
09
0>
0C
#108470000000
1!
1*
b101 6
19
1>
1C
b101 G
#108480000000
0!
0*
09
0>
0C
#108490000000
1!
1*
b110 6
19
1>
1C
b110 G
#108500000000
0!
0*
09
0>
0C
#108510000000
1!
1*
b111 6
19
1>
1C
b111 G
#108520000000
0!
0*
09
0>
0C
#108530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#108540000000
0!
0*
09
0>
0C
#108550000000
1!
1*
b1 6
19
1>
1C
b1 G
#108560000000
0!
0*
09
0>
0C
#108570000000
1!
1*
b10 6
19
1>
1C
b10 G
#108580000000
0!
0*
09
0>
0C
#108590000000
1!
1*
b11 6
19
1>
1C
b11 G
#108600000000
0!
0*
09
0>
0C
#108610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#108620000000
0!
0*
09
0>
0C
#108630000000
1!
1*
b101 6
19
1>
1C
b101 G
#108640000000
0!
0*
09
0>
0C
#108650000000
1!
1*
b110 6
19
1>
1C
b110 G
#108660000000
0!
0*
09
0>
0C
#108670000000
1!
1*
b111 6
19
1>
1C
b111 G
#108680000000
0!
0*
09
0>
0C
#108690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#108700000000
0!
0*
09
0>
0C
#108710000000
1!
1*
b1 6
19
1>
1C
b1 G
#108720000000
0!
0*
09
0>
0C
#108730000000
1!
1*
b10 6
19
1>
1C
b10 G
#108740000000
0!
0*
09
0>
0C
#108750000000
1!
1*
b11 6
19
1>
1C
b11 G
#108760000000
0!
0*
09
0>
0C
#108770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#108780000000
0!
0*
09
0>
0C
#108790000000
1!
1*
b101 6
19
1>
1C
b101 G
#108800000000
0!
0*
09
0>
0C
#108810000000
1!
1*
b110 6
19
1>
1C
b110 G
#108820000000
0!
0*
09
0>
0C
#108830000000
1!
1*
b111 6
19
1>
1C
b111 G
#108840000000
0!
1"
0*
1+
09
1:
0>
0C
#108850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#108860000000
0!
0*
09
0>
0C
#108870000000
1!
1*
b1 6
19
1>
1C
b1 G
#108880000000
0!
0*
09
0>
0C
#108890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#108900000000
0!
0*
09
0>
0C
#108910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#108920000000
0!
0*
09
0>
0C
#108930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#108940000000
0!
0*
09
0>
0C
#108950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#108960000000
0!
0#
0*
0,
09
0>
0?
0C
#108970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#108980000000
0!
0*
09
0>
0C
#108990000000
1!
1*
19
1>
1C
#109000000000
0!
0*
09
0>
0C
#109010000000
1!
1*
19
1>
1C
#109020000000
0!
0*
09
0>
0C
#109030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#109040000000
0!
0*
09
0>
0C
#109050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#109060000000
0!
0*
09
0>
0C
#109070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#109080000000
0!
0*
09
0>
0C
#109090000000
1!
1*
b10 6
19
1>
1C
b10 G
#109100000000
0!
0*
09
0>
0C
#109110000000
1!
1*
b11 6
19
1>
1C
b11 G
#109120000000
0!
0*
09
0>
0C
#109130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#109140000000
0!
0*
09
0>
0C
#109150000000
1!
1*
b101 6
19
1>
1C
b101 G
#109160000000
0!
0*
09
0>
0C
#109170000000
1!
1*
b110 6
19
1>
1C
b110 G
#109180000000
0!
0*
09
0>
0C
#109190000000
1!
1*
b111 6
19
1>
1C
b111 G
#109200000000
0!
0*
09
0>
0C
#109210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#109220000000
0!
0*
09
0>
0C
#109230000000
1!
1*
b1 6
19
1>
1C
b1 G
#109240000000
0!
0*
09
0>
0C
#109250000000
1!
1*
b10 6
19
1>
1C
b10 G
#109260000000
0!
0*
09
0>
0C
#109270000000
1!
1*
b11 6
19
1>
1C
b11 G
#109280000000
0!
0*
09
0>
0C
#109290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#109300000000
0!
0*
09
0>
0C
#109310000000
1!
1*
b101 6
19
1>
1C
b101 G
#109320000000
0!
0*
09
0>
0C
#109330000000
1!
1*
b110 6
19
1>
1C
b110 G
#109340000000
0!
0*
09
0>
0C
#109350000000
1!
1*
b111 6
19
1>
1C
b111 G
#109360000000
0!
0*
09
0>
0C
#109370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#109380000000
0!
0*
09
0>
0C
#109390000000
1!
1*
b1 6
19
1>
1C
b1 G
#109400000000
0!
0*
09
0>
0C
#109410000000
1!
1*
b10 6
19
1>
1C
b10 G
#109420000000
0!
0*
09
0>
0C
#109430000000
1!
1*
b11 6
19
1>
1C
b11 G
#109440000000
0!
0*
09
0>
0C
#109450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#109460000000
0!
0*
09
0>
0C
#109470000000
1!
1*
b101 6
19
1>
1C
b101 G
#109480000000
0!
0*
09
0>
0C
#109490000000
1!
1*
b110 6
19
1>
1C
b110 G
#109500000000
0!
0*
09
0>
0C
#109510000000
1!
1*
b111 6
19
1>
1C
b111 G
#109520000000
0!
1"
0*
1+
09
1:
0>
0C
#109530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#109540000000
0!
0*
09
0>
0C
#109550000000
1!
1*
b1 6
19
1>
1C
b1 G
#109560000000
0!
0*
09
0>
0C
#109570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#109580000000
0!
0*
09
0>
0C
#109590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#109600000000
0!
0*
09
0>
0C
#109610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#109620000000
0!
0*
09
0>
0C
#109630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#109640000000
0!
0#
0*
0,
09
0>
0?
0C
#109650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#109660000000
0!
0*
09
0>
0C
#109670000000
1!
1*
19
1>
1C
#109680000000
0!
0*
09
0>
0C
#109690000000
1!
1*
19
1>
1C
#109700000000
0!
0*
09
0>
0C
#109710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#109720000000
0!
0*
09
0>
0C
#109730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#109740000000
0!
0*
09
0>
0C
#109750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#109760000000
0!
0*
09
0>
0C
#109770000000
1!
1*
b10 6
19
1>
1C
b10 G
#109780000000
0!
0*
09
0>
0C
#109790000000
1!
1*
b11 6
19
1>
1C
b11 G
#109800000000
0!
0*
09
0>
0C
#109810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#109820000000
0!
0*
09
0>
0C
#109830000000
1!
1*
b101 6
19
1>
1C
b101 G
#109840000000
0!
0*
09
0>
0C
#109850000000
1!
1*
b110 6
19
1>
1C
b110 G
#109860000000
0!
0*
09
0>
0C
#109870000000
1!
1*
b111 6
19
1>
1C
b111 G
#109880000000
0!
0*
09
0>
0C
#109890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#109900000000
0!
0*
09
0>
0C
#109910000000
1!
1*
b1 6
19
1>
1C
b1 G
#109920000000
0!
0*
09
0>
0C
#109930000000
1!
1*
b10 6
19
1>
1C
b10 G
#109940000000
0!
0*
09
0>
0C
#109950000000
1!
1*
b11 6
19
1>
1C
b11 G
#109960000000
0!
0*
09
0>
0C
#109970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#109980000000
0!
0*
09
0>
0C
#109990000000
1!
1*
b101 6
19
1>
1C
b101 G
#110000000000
0!
0*
09
0>
0C
#110010000000
1!
1*
b110 6
19
1>
1C
b110 G
#110020000000
0!
0*
09
0>
0C
#110030000000
1!
1*
b111 6
19
1>
1C
b111 G
#110040000000
0!
0*
09
0>
0C
#110050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#110060000000
0!
0*
09
0>
0C
#110070000000
1!
1*
b1 6
19
1>
1C
b1 G
#110080000000
0!
0*
09
0>
0C
#110090000000
1!
1*
b10 6
19
1>
1C
b10 G
#110100000000
0!
0*
09
0>
0C
#110110000000
1!
1*
b11 6
19
1>
1C
b11 G
#110120000000
0!
0*
09
0>
0C
#110130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#110140000000
0!
0*
09
0>
0C
#110150000000
1!
1*
b101 6
19
1>
1C
b101 G
#110160000000
0!
0*
09
0>
0C
#110170000000
1!
1*
b110 6
19
1>
1C
b110 G
#110180000000
0!
0*
09
0>
0C
#110190000000
1!
1*
b111 6
19
1>
1C
b111 G
#110200000000
0!
1"
0*
1+
09
1:
0>
0C
#110210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#110220000000
0!
0*
09
0>
0C
#110230000000
1!
1*
b1 6
19
1>
1C
b1 G
#110240000000
0!
0*
09
0>
0C
#110250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#110260000000
0!
0*
09
0>
0C
#110270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#110280000000
0!
0*
09
0>
0C
#110290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#110300000000
0!
0*
09
0>
0C
#110310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#110320000000
0!
0#
0*
0,
09
0>
0?
0C
#110330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#110340000000
0!
0*
09
0>
0C
#110350000000
1!
1*
19
1>
1C
#110360000000
0!
0*
09
0>
0C
#110370000000
1!
1*
19
1>
1C
#110380000000
0!
0*
09
0>
0C
#110390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#110400000000
0!
0*
09
0>
0C
#110410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#110420000000
0!
0*
09
0>
0C
#110430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#110440000000
0!
0*
09
0>
0C
#110450000000
1!
1*
b10 6
19
1>
1C
b10 G
#110460000000
0!
0*
09
0>
0C
#110470000000
1!
1*
b11 6
19
1>
1C
b11 G
#110480000000
0!
0*
09
0>
0C
#110490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#110500000000
0!
0*
09
0>
0C
#110510000000
1!
1*
b101 6
19
1>
1C
b101 G
#110520000000
0!
0*
09
0>
0C
#110530000000
1!
1*
b110 6
19
1>
1C
b110 G
#110540000000
0!
0*
09
0>
0C
#110550000000
1!
1*
b111 6
19
1>
1C
b111 G
#110560000000
0!
0*
09
0>
0C
#110570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#110580000000
0!
0*
09
0>
0C
#110590000000
1!
1*
b1 6
19
1>
1C
b1 G
#110600000000
0!
0*
09
0>
0C
#110610000000
1!
1*
b10 6
19
1>
1C
b10 G
#110620000000
0!
0*
09
0>
0C
#110630000000
1!
1*
b11 6
19
1>
1C
b11 G
#110640000000
0!
0*
09
0>
0C
#110650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#110660000000
0!
0*
09
0>
0C
#110670000000
1!
1*
b101 6
19
1>
1C
b101 G
#110680000000
0!
0*
09
0>
0C
#110690000000
1!
1*
b110 6
19
1>
1C
b110 G
#110700000000
0!
0*
09
0>
0C
#110710000000
1!
1*
b111 6
19
1>
1C
b111 G
#110720000000
0!
0*
09
0>
0C
#110730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#110740000000
0!
0*
09
0>
0C
#110750000000
1!
1*
b1 6
19
1>
1C
b1 G
#110760000000
0!
0*
09
0>
0C
#110770000000
1!
1*
b10 6
19
1>
1C
b10 G
#110780000000
0!
0*
09
0>
0C
#110790000000
1!
1*
b11 6
19
1>
1C
b11 G
#110800000000
0!
0*
09
0>
0C
#110810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#110820000000
0!
0*
09
0>
0C
#110830000000
1!
1*
b101 6
19
1>
1C
b101 G
#110840000000
0!
0*
09
0>
0C
#110850000000
1!
1*
b110 6
19
1>
1C
b110 G
#110860000000
0!
0*
09
0>
0C
#110870000000
1!
1*
b111 6
19
1>
1C
b111 G
#110880000000
0!
1"
0*
1+
09
1:
0>
0C
#110890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#110900000000
0!
0*
09
0>
0C
#110910000000
1!
1*
b1 6
19
1>
1C
b1 G
#110920000000
0!
0*
09
0>
0C
#110930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#110940000000
0!
0*
09
0>
0C
#110950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#110960000000
0!
0*
09
0>
0C
#110970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#110980000000
0!
0*
09
0>
0C
#110990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#111000000000
0!
0#
0*
0,
09
0>
0?
0C
#111010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#111020000000
0!
0*
09
0>
0C
#111030000000
1!
1*
19
1>
1C
#111040000000
0!
0*
09
0>
0C
#111050000000
1!
1*
19
1>
1C
#111060000000
0!
0*
09
0>
0C
#111070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#111080000000
0!
0*
09
0>
0C
#111090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#111100000000
0!
0*
09
0>
0C
#111110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#111120000000
0!
0*
09
0>
0C
#111130000000
1!
1*
b10 6
19
1>
1C
b10 G
#111140000000
0!
0*
09
0>
0C
#111150000000
1!
1*
b11 6
19
1>
1C
b11 G
#111160000000
0!
0*
09
0>
0C
#111170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#111180000000
0!
0*
09
0>
0C
#111190000000
1!
1*
b101 6
19
1>
1C
b101 G
#111200000000
0!
0*
09
0>
0C
#111210000000
1!
1*
b110 6
19
1>
1C
b110 G
#111220000000
0!
0*
09
0>
0C
#111230000000
1!
1*
b111 6
19
1>
1C
b111 G
#111240000000
0!
0*
09
0>
0C
#111250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#111260000000
0!
0*
09
0>
0C
#111270000000
1!
1*
b1 6
19
1>
1C
b1 G
#111280000000
0!
0*
09
0>
0C
#111290000000
1!
1*
b10 6
19
1>
1C
b10 G
#111300000000
0!
0*
09
0>
0C
#111310000000
1!
1*
b11 6
19
1>
1C
b11 G
#111320000000
0!
0*
09
0>
0C
#111330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#111340000000
0!
0*
09
0>
0C
#111350000000
1!
1*
b101 6
19
1>
1C
b101 G
#111360000000
0!
0*
09
0>
0C
#111370000000
1!
1*
b110 6
19
1>
1C
b110 G
#111380000000
0!
0*
09
0>
0C
#111390000000
1!
1*
b111 6
19
1>
1C
b111 G
#111400000000
0!
0*
09
0>
0C
#111410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#111420000000
0!
0*
09
0>
0C
#111430000000
1!
1*
b1 6
19
1>
1C
b1 G
#111440000000
0!
0*
09
0>
0C
#111450000000
1!
1*
b10 6
19
1>
1C
b10 G
#111460000000
0!
0*
09
0>
0C
#111470000000
1!
1*
b11 6
19
1>
1C
b11 G
#111480000000
0!
0*
09
0>
0C
#111490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#111500000000
0!
0*
09
0>
0C
#111510000000
1!
1*
b101 6
19
1>
1C
b101 G
#111520000000
0!
0*
09
0>
0C
#111530000000
1!
1*
b110 6
19
1>
1C
b110 G
#111540000000
0!
0*
09
0>
0C
#111550000000
1!
1*
b111 6
19
1>
1C
b111 G
#111560000000
0!
1"
0*
1+
09
1:
0>
0C
#111570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#111580000000
0!
0*
09
0>
0C
#111590000000
1!
1*
b1 6
19
1>
1C
b1 G
#111600000000
0!
0*
09
0>
0C
#111610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#111620000000
0!
0*
09
0>
0C
#111630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#111640000000
0!
0*
09
0>
0C
#111650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#111660000000
0!
0*
09
0>
0C
#111670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#111680000000
0!
0#
0*
0,
09
0>
0?
0C
#111690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#111700000000
0!
0*
09
0>
0C
#111710000000
1!
1*
19
1>
1C
#111720000000
0!
0*
09
0>
0C
#111730000000
1!
1*
19
1>
1C
#111740000000
0!
0*
09
0>
0C
#111750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#111760000000
0!
0*
09
0>
0C
#111770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#111780000000
0!
0*
09
0>
0C
#111790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#111800000000
0!
0*
09
0>
0C
#111810000000
1!
1*
b10 6
19
1>
1C
b10 G
#111820000000
0!
0*
09
0>
0C
#111830000000
1!
1*
b11 6
19
1>
1C
b11 G
#111840000000
0!
0*
09
0>
0C
#111850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#111860000000
0!
0*
09
0>
0C
#111870000000
1!
1*
b101 6
19
1>
1C
b101 G
#111880000000
0!
0*
09
0>
0C
#111890000000
1!
1*
b110 6
19
1>
1C
b110 G
#111900000000
0!
0*
09
0>
0C
#111910000000
1!
1*
b111 6
19
1>
1C
b111 G
#111920000000
0!
0*
09
0>
0C
#111930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#111940000000
0!
0*
09
0>
0C
#111950000000
1!
1*
b1 6
19
1>
1C
b1 G
#111960000000
0!
0*
09
0>
0C
#111970000000
1!
1*
b10 6
19
1>
1C
b10 G
#111980000000
0!
0*
09
0>
0C
#111990000000
1!
1*
b11 6
19
1>
1C
b11 G
#112000000000
0!
0*
09
0>
0C
#112010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#112020000000
0!
0*
09
0>
0C
#112030000000
1!
1*
b101 6
19
1>
1C
b101 G
#112040000000
0!
0*
09
0>
0C
#112050000000
1!
1*
b110 6
19
1>
1C
b110 G
#112060000000
0!
0*
09
0>
0C
#112070000000
1!
1*
b111 6
19
1>
1C
b111 G
#112080000000
0!
0*
09
0>
0C
#112090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#112100000000
0!
0*
09
0>
0C
#112110000000
1!
1*
b1 6
19
1>
1C
b1 G
#112120000000
0!
0*
09
0>
0C
#112130000000
1!
1*
b10 6
19
1>
1C
b10 G
#112140000000
0!
0*
09
0>
0C
#112150000000
1!
1*
b11 6
19
1>
1C
b11 G
#112160000000
0!
0*
09
0>
0C
#112170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#112180000000
0!
0*
09
0>
0C
#112190000000
1!
1*
b101 6
19
1>
1C
b101 G
#112200000000
0!
0*
09
0>
0C
#112210000000
1!
1*
b110 6
19
1>
1C
b110 G
#112220000000
0!
0*
09
0>
0C
#112230000000
1!
1*
b111 6
19
1>
1C
b111 G
#112240000000
0!
1"
0*
1+
09
1:
0>
0C
#112250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#112260000000
0!
0*
09
0>
0C
#112270000000
1!
1*
b1 6
19
1>
1C
b1 G
#112280000000
0!
0*
09
0>
0C
#112290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#112300000000
0!
0*
09
0>
0C
#112310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#112320000000
0!
0*
09
0>
0C
#112330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#112340000000
0!
0*
09
0>
0C
#112350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#112360000000
0!
0#
0*
0,
09
0>
0?
0C
#112370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#112380000000
0!
0*
09
0>
0C
#112390000000
1!
1*
19
1>
1C
#112400000000
0!
0*
09
0>
0C
#112410000000
1!
1*
19
1>
1C
#112420000000
0!
0*
09
0>
0C
#112430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#112440000000
0!
0*
09
0>
0C
#112450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#112460000000
0!
0*
09
0>
0C
#112470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#112480000000
0!
0*
09
0>
0C
#112490000000
1!
1*
b10 6
19
1>
1C
b10 G
#112500000000
0!
0*
09
0>
0C
#112510000000
1!
1*
b11 6
19
1>
1C
b11 G
#112520000000
0!
0*
09
0>
0C
#112530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#112540000000
0!
0*
09
0>
0C
#112550000000
1!
1*
b101 6
19
1>
1C
b101 G
#112560000000
0!
0*
09
0>
0C
#112570000000
1!
1*
b110 6
19
1>
1C
b110 G
#112580000000
0!
0*
09
0>
0C
#112590000000
1!
1*
b111 6
19
1>
1C
b111 G
#112600000000
0!
0*
09
0>
0C
#112610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#112620000000
0!
0*
09
0>
0C
#112630000000
1!
1*
b1 6
19
1>
1C
b1 G
#112640000000
0!
0*
09
0>
0C
#112650000000
1!
1*
b10 6
19
1>
1C
b10 G
#112660000000
0!
0*
09
0>
0C
#112670000000
1!
1*
b11 6
19
1>
1C
b11 G
#112680000000
0!
0*
09
0>
0C
#112690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#112700000000
0!
0*
09
0>
0C
#112710000000
1!
1*
b101 6
19
1>
1C
b101 G
#112720000000
0!
0*
09
0>
0C
#112730000000
1!
1*
b110 6
19
1>
1C
b110 G
#112740000000
0!
0*
09
0>
0C
#112750000000
1!
1*
b111 6
19
1>
1C
b111 G
#112760000000
0!
0*
09
0>
0C
#112770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#112780000000
0!
0*
09
0>
0C
#112790000000
1!
1*
b1 6
19
1>
1C
b1 G
#112800000000
0!
0*
09
0>
0C
#112810000000
1!
1*
b10 6
19
1>
1C
b10 G
#112820000000
0!
0*
09
0>
0C
#112830000000
1!
1*
b11 6
19
1>
1C
b11 G
#112840000000
0!
0*
09
0>
0C
#112850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#112860000000
0!
0*
09
0>
0C
#112870000000
1!
1*
b101 6
19
1>
1C
b101 G
#112880000000
0!
0*
09
0>
0C
#112890000000
1!
1*
b110 6
19
1>
1C
b110 G
#112900000000
0!
0*
09
0>
0C
#112910000000
1!
1*
b111 6
19
1>
1C
b111 G
#112920000000
0!
1"
0*
1+
09
1:
0>
0C
#112930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#112940000000
0!
0*
09
0>
0C
#112950000000
1!
1*
b1 6
19
1>
1C
b1 G
#112960000000
0!
0*
09
0>
0C
#112970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#112980000000
0!
0*
09
0>
0C
#112990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#113000000000
0!
0*
09
0>
0C
#113010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#113020000000
0!
0*
09
0>
0C
#113030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#113040000000
0!
0#
0*
0,
09
0>
0?
0C
#113050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#113060000000
0!
0*
09
0>
0C
#113070000000
1!
1*
19
1>
1C
#113080000000
0!
0*
09
0>
0C
#113090000000
1!
1*
19
1>
1C
#113100000000
0!
0*
09
0>
0C
#113110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#113120000000
0!
0*
09
0>
0C
#113130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#113140000000
0!
0*
09
0>
0C
#113150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#113160000000
0!
0*
09
0>
0C
#113170000000
1!
1*
b10 6
19
1>
1C
b10 G
#113180000000
0!
0*
09
0>
0C
#113190000000
1!
1*
b11 6
19
1>
1C
b11 G
#113200000000
0!
0*
09
0>
0C
#113210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#113220000000
0!
0*
09
0>
0C
#113230000000
1!
1*
b101 6
19
1>
1C
b101 G
#113240000000
0!
0*
09
0>
0C
#113250000000
1!
1*
b110 6
19
1>
1C
b110 G
#113260000000
0!
0*
09
0>
0C
#113270000000
1!
1*
b111 6
19
1>
1C
b111 G
#113280000000
0!
0*
09
0>
0C
#113290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#113300000000
0!
0*
09
0>
0C
#113310000000
1!
1*
b1 6
19
1>
1C
b1 G
#113320000000
0!
0*
09
0>
0C
#113330000000
1!
1*
b10 6
19
1>
1C
b10 G
#113340000000
0!
0*
09
0>
0C
#113350000000
1!
1*
b11 6
19
1>
1C
b11 G
#113360000000
0!
0*
09
0>
0C
#113370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#113380000000
0!
0*
09
0>
0C
#113390000000
1!
1*
b101 6
19
1>
1C
b101 G
#113400000000
0!
0*
09
0>
0C
#113410000000
1!
1*
b110 6
19
1>
1C
b110 G
#113420000000
0!
0*
09
0>
0C
#113430000000
1!
1*
b111 6
19
1>
1C
b111 G
#113440000000
0!
0*
09
0>
0C
#113450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#113460000000
0!
0*
09
0>
0C
#113470000000
1!
1*
b1 6
19
1>
1C
b1 G
#113480000000
0!
0*
09
0>
0C
#113490000000
1!
1*
b10 6
19
1>
1C
b10 G
#113500000000
0!
0*
09
0>
0C
#113510000000
1!
1*
b11 6
19
1>
1C
b11 G
#113520000000
0!
0*
09
0>
0C
#113530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#113540000000
0!
0*
09
0>
0C
#113550000000
1!
1*
b101 6
19
1>
1C
b101 G
#113560000000
0!
0*
09
0>
0C
#113570000000
1!
1*
b110 6
19
1>
1C
b110 G
#113580000000
0!
0*
09
0>
0C
#113590000000
1!
1*
b111 6
19
1>
1C
b111 G
#113600000000
0!
1"
0*
1+
09
1:
0>
0C
#113610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#113620000000
0!
0*
09
0>
0C
#113630000000
1!
1*
b1 6
19
1>
1C
b1 G
#113640000000
0!
0*
09
0>
0C
#113650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#113660000000
0!
0*
09
0>
0C
#113670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#113680000000
0!
0*
09
0>
0C
#113690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#113700000000
0!
0*
09
0>
0C
#113710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#113720000000
0!
0#
0*
0,
09
0>
0?
0C
#113730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#113740000000
0!
0*
09
0>
0C
#113750000000
1!
1*
19
1>
1C
#113760000000
0!
0*
09
0>
0C
#113770000000
1!
1*
19
1>
1C
#113780000000
0!
0*
09
0>
0C
#113790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#113800000000
0!
0*
09
0>
0C
#113810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#113820000000
0!
0*
09
0>
0C
#113830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#113840000000
0!
0*
09
0>
0C
#113850000000
1!
1*
b10 6
19
1>
1C
b10 G
#113860000000
0!
0*
09
0>
0C
#113870000000
1!
1*
b11 6
19
1>
1C
b11 G
#113880000000
0!
0*
09
0>
0C
#113890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#113900000000
0!
0*
09
0>
0C
#113910000000
1!
1*
b101 6
19
1>
1C
b101 G
#113920000000
0!
0*
09
0>
0C
#113930000000
1!
1*
b110 6
19
1>
1C
b110 G
#113940000000
0!
0*
09
0>
0C
#113950000000
1!
1*
b111 6
19
1>
1C
b111 G
#113960000000
0!
0*
09
0>
0C
#113970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#113980000000
0!
0*
09
0>
0C
#113990000000
1!
1*
b1 6
19
1>
1C
b1 G
#114000000000
0!
0*
09
0>
0C
#114010000000
1!
1*
b10 6
19
1>
1C
b10 G
#114020000000
0!
0*
09
0>
0C
#114030000000
1!
1*
b11 6
19
1>
1C
b11 G
#114040000000
0!
0*
09
0>
0C
#114050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#114060000000
0!
0*
09
0>
0C
#114070000000
1!
1*
b101 6
19
1>
1C
b101 G
#114080000000
0!
0*
09
0>
0C
#114090000000
1!
1*
b110 6
19
1>
1C
b110 G
#114100000000
0!
0*
09
0>
0C
#114110000000
1!
1*
b111 6
19
1>
1C
b111 G
#114120000000
0!
0*
09
0>
0C
#114130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#114140000000
0!
0*
09
0>
0C
#114150000000
1!
1*
b1 6
19
1>
1C
b1 G
#114160000000
0!
0*
09
0>
0C
#114170000000
1!
1*
b10 6
19
1>
1C
b10 G
#114180000000
0!
0*
09
0>
0C
#114190000000
1!
1*
b11 6
19
1>
1C
b11 G
#114200000000
0!
0*
09
0>
0C
#114210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#114220000000
0!
0*
09
0>
0C
#114230000000
1!
1*
b101 6
19
1>
1C
b101 G
#114240000000
0!
0*
09
0>
0C
#114250000000
1!
1*
b110 6
19
1>
1C
b110 G
#114260000000
0!
0*
09
0>
0C
#114270000000
1!
1*
b111 6
19
1>
1C
b111 G
#114280000000
0!
1"
0*
1+
09
1:
0>
0C
#114290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#114300000000
0!
0*
09
0>
0C
#114310000000
1!
1*
b1 6
19
1>
1C
b1 G
#114320000000
0!
0*
09
0>
0C
#114330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#114340000000
0!
0*
09
0>
0C
#114350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#114360000000
0!
0*
09
0>
0C
#114370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#114380000000
0!
0*
09
0>
0C
#114390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#114400000000
0!
0#
0*
0,
09
0>
0?
0C
#114410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#114420000000
0!
0*
09
0>
0C
#114430000000
1!
1*
19
1>
1C
#114440000000
0!
0*
09
0>
0C
#114450000000
1!
1*
19
1>
1C
#114460000000
0!
0*
09
0>
0C
#114470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#114480000000
0!
0*
09
0>
0C
#114490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#114500000000
0!
0*
09
0>
0C
#114510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#114520000000
0!
0*
09
0>
0C
#114530000000
1!
1*
b10 6
19
1>
1C
b10 G
#114540000000
0!
0*
09
0>
0C
#114550000000
1!
1*
b11 6
19
1>
1C
b11 G
#114560000000
0!
0*
09
0>
0C
#114570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#114580000000
0!
0*
09
0>
0C
#114590000000
1!
1*
b101 6
19
1>
1C
b101 G
#114600000000
0!
0*
09
0>
0C
#114610000000
1!
1*
b110 6
19
1>
1C
b110 G
#114620000000
0!
0*
09
0>
0C
#114630000000
1!
1*
b111 6
19
1>
1C
b111 G
#114640000000
0!
0*
09
0>
0C
#114650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#114660000000
0!
0*
09
0>
0C
#114670000000
1!
1*
b1 6
19
1>
1C
b1 G
#114680000000
0!
0*
09
0>
0C
#114690000000
1!
1*
b10 6
19
1>
1C
b10 G
#114700000000
0!
0*
09
0>
0C
#114710000000
1!
1*
b11 6
19
1>
1C
b11 G
#114720000000
0!
0*
09
0>
0C
#114730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#114740000000
0!
0*
09
0>
0C
#114750000000
1!
1*
b101 6
19
1>
1C
b101 G
#114760000000
0!
0*
09
0>
0C
#114770000000
1!
1*
b110 6
19
1>
1C
b110 G
#114780000000
0!
0*
09
0>
0C
#114790000000
1!
1*
b111 6
19
1>
1C
b111 G
#114800000000
0!
0*
09
0>
0C
#114810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#114820000000
0!
0*
09
0>
0C
#114830000000
1!
1*
b1 6
19
1>
1C
b1 G
#114840000000
0!
0*
09
0>
0C
#114850000000
1!
1*
b10 6
19
1>
1C
b10 G
#114860000000
0!
0*
09
0>
0C
#114870000000
1!
1*
b11 6
19
1>
1C
b11 G
#114880000000
0!
0*
09
0>
0C
#114890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#114900000000
0!
0*
09
0>
0C
#114910000000
1!
1*
b101 6
19
1>
1C
b101 G
#114920000000
0!
0*
09
0>
0C
#114930000000
1!
1*
b110 6
19
1>
1C
b110 G
#114940000000
0!
0*
09
0>
0C
#114950000000
1!
1*
b111 6
19
1>
1C
b111 G
#114960000000
0!
1"
0*
1+
09
1:
0>
0C
#114970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#114980000000
0!
0*
09
0>
0C
#114990000000
1!
1*
b1 6
19
1>
1C
b1 G
#115000000000
0!
0*
09
0>
0C
#115010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#115020000000
0!
0*
09
0>
0C
#115030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#115040000000
0!
0*
09
0>
0C
#115050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#115060000000
0!
0*
09
0>
0C
#115070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#115080000000
0!
0#
0*
0,
09
0>
0?
0C
#115090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#115100000000
0!
0*
09
0>
0C
#115110000000
1!
1*
19
1>
1C
#115120000000
0!
0*
09
0>
0C
#115130000000
1!
1*
19
1>
1C
#115140000000
0!
0*
09
0>
0C
#115150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#115160000000
0!
0*
09
0>
0C
#115170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#115180000000
0!
0*
09
0>
0C
#115190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#115200000000
0!
0*
09
0>
0C
#115210000000
1!
1*
b10 6
19
1>
1C
b10 G
#115220000000
0!
0*
09
0>
0C
#115230000000
1!
1*
b11 6
19
1>
1C
b11 G
#115240000000
0!
0*
09
0>
0C
#115250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#115260000000
0!
0*
09
0>
0C
#115270000000
1!
1*
b101 6
19
1>
1C
b101 G
#115280000000
0!
0*
09
0>
0C
#115290000000
1!
1*
b110 6
19
1>
1C
b110 G
#115300000000
0!
0*
09
0>
0C
#115310000000
1!
1*
b111 6
19
1>
1C
b111 G
#115320000000
0!
0*
09
0>
0C
#115330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#115340000000
0!
0*
09
0>
0C
#115350000000
1!
1*
b1 6
19
1>
1C
b1 G
#115360000000
0!
0*
09
0>
0C
#115370000000
1!
1*
b10 6
19
1>
1C
b10 G
#115380000000
0!
0*
09
0>
0C
#115390000000
1!
1*
b11 6
19
1>
1C
b11 G
#115400000000
0!
0*
09
0>
0C
#115410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#115420000000
0!
0*
09
0>
0C
#115430000000
1!
1*
b101 6
19
1>
1C
b101 G
#115440000000
0!
0*
09
0>
0C
#115450000000
1!
1*
b110 6
19
1>
1C
b110 G
#115460000000
0!
0*
09
0>
0C
#115470000000
1!
1*
b111 6
19
1>
1C
b111 G
#115480000000
0!
0*
09
0>
0C
#115490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#115500000000
0!
0*
09
0>
0C
#115510000000
1!
1*
b1 6
19
1>
1C
b1 G
#115520000000
0!
0*
09
0>
0C
#115530000000
1!
1*
b10 6
19
1>
1C
b10 G
#115540000000
0!
0*
09
0>
0C
#115550000000
1!
1*
b11 6
19
1>
1C
b11 G
#115560000000
0!
0*
09
0>
0C
#115570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#115580000000
0!
0*
09
0>
0C
#115590000000
1!
1*
b101 6
19
1>
1C
b101 G
#115600000000
0!
0*
09
0>
0C
#115610000000
1!
1*
b110 6
19
1>
1C
b110 G
#115620000000
0!
0*
09
0>
0C
#115630000000
1!
1*
b111 6
19
1>
1C
b111 G
#115640000000
0!
1"
0*
1+
09
1:
0>
0C
#115650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#115660000000
0!
0*
09
0>
0C
#115670000000
1!
1*
b1 6
19
1>
1C
b1 G
#115680000000
0!
0*
09
0>
0C
#115690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#115700000000
0!
0*
09
0>
0C
#115710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#115720000000
0!
0*
09
0>
0C
#115730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#115740000000
0!
0*
09
0>
0C
#115750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#115760000000
0!
0#
0*
0,
09
0>
0?
0C
#115770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#115780000000
0!
0*
09
0>
0C
#115790000000
1!
1*
19
1>
1C
#115800000000
0!
0*
09
0>
0C
#115810000000
1!
1*
19
1>
1C
#115820000000
0!
0*
09
0>
0C
#115830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#115840000000
0!
0*
09
0>
0C
#115850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#115860000000
0!
0*
09
0>
0C
#115870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#115880000000
0!
0*
09
0>
0C
#115890000000
1!
1*
b10 6
19
1>
1C
b10 G
#115900000000
0!
0*
09
0>
0C
#115910000000
1!
1*
b11 6
19
1>
1C
b11 G
#115920000000
0!
0*
09
0>
0C
#115930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#115940000000
0!
0*
09
0>
0C
#115950000000
1!
1*
b101 6
19
1>
1C
b101 G
#115960000000
0!
0*
09
0>
0C
#115970000000
1!
1*
b110 6
19
1>
1C
b110 G
#115980000000
0!
0*
09
0>
0C
#115990000000
1!
1*
b111 6
19
1>
1C
b111 G
#116000000000
0!
0*
09
0>
0C
#116010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#116020000000
0!
0*
09
0>
0C
#116030000000
1!
1*
b1 6
19
1>
1C
b1 G
#116040000000
0!
0*
09
0>
0C
#116050000000
1!
1*
b10 6
19
1>
1C
b10 G
#116060000000
0!
0*
09
0>
0C
#116070000000
1!
1*
b11 6
19
1>
1C
b11 G
#116080000000
0!
0*
09
0>
0C
#116090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#116100000000
0!
0*
09
0>
0C
#116110000000
1!
1*
b101 6
19
1>
1C
b101 G
#116120000000
0!
0*
09
0>
0C
#116130000000
1!
1*
b110 6
19
1>
1C
b110 G
#116140000000
0!
0*
09
0>
0C
#116150000000
1!
1*
b111 6
19
1>
1C
b111 G
#116160000000
0!
0*
09
0>
0C
#116170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#116180000000
0!
0*
09
0>
0C
#116190000000
1!
1*
b1 6
19
1>
1C
b1 G
#116200000000
0!
0*
09
0>
0C
#116210000000
1!
1*
b10 6
19
1>
1C
b10 G
#116220000000
0!
0*
09
0>
0C
#116230000000
1!
1*
b11 6
19
1>
1C
b11 G
#116240000000
0!
0*
09
0>
0C
#116250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#116260000000
0!
0*
09
0>
0C
#116270000000
1!
1*
b101 6
19
1>
1C
b101 G
#116280000000
0!
0*
09
0>
0C
#116290000000
1!
1*
b110 6
19
1>
1C
b110 G
#116300000000
0!
0*
09
0>
0C
#116310000000
1!
1*
b111 6
19
1>
1C
b111 G
#116320000000
0!
1"
0*
1+
09
1:
0>
0C
#116330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#116340000000
0!
0*
09
0>
0C
#116350000000
1!
1*
b1 6
19
1>
1C
b1 G
#116360000000
0!
0*
09
0>
0C
#116370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#116380000000
0!
0*
09
0>
0C
#116390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#116400000000
0!
0*
09
0>
0C
#116410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#116420000000
0!
0*
09
0>
0C
#116430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#116440000000
0!
0#
0*
0,
09
0>
0?
0C
#116450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#116460000000
0!
0*
09
0>
0C
#116470000000
1!
1*
19
1>
1C
#116480000000
0!
0*
09
0>
0C
#116490000000
1!
1*
19
1>
1C
#116500000000
0!
0*
09
0>
0C
#116510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#116520000000
0!
0*
09
0>
0C
#116530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#116540000000
0!
0*
09
0>
0C
#116550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#116560000000
0!
0*
09
0>
0C
#116570000000
1!
1*
b10 6
19
1>
1C
b10 G
#116580000000
0!
0*
09
0>
0C
#116590000000
1!
1*
b11 6
19
1>
1C
b11 G
#116600000000
0!
0*
09
0>
0C
#116610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#116620000000
0!
0*
09
0>
0C
#116630000000
1!
1*
b101 6
19
1>
1C
b101 G
#116640000000
0!
0*
09
0>
0C
#116650000000
1!
1*
b110 6
19
1>
1C
b110 G
#116660000000
0!
0*
09
0>
0C
#116670000000
1!
1*
b111 6
19
1>
1C
b111 G
#116680000000
0!
0*
09
0>
0C
#116690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#116700000000
0!
0*
09
0>
0C
#116710000000
1!
1*
b1 6
19
1>
1C
b1 G
#116720000000
0!
0*
09
0>
0C
#116730000000
1!
1*
b10 6
19
1>
1C
b10 G
#116740000000
0!
0*
09
0>
0C
#116750000000
1!
1*
b11 6
19
1>
1C
b11 G
#116760000000
0!
0*
09
0>
0C
#116770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#116780000000
0!
0*
09
0>
0C
#116790000000
1!
1*
b101 6
19
1>
1C
b101 G
#116800000000
0!
0*
09
0>
0C
#116810000000
1!
1*
b110 6
19
1>
1C
b110 G
#116820000000
0!
0*
09
0>
0C
#116830000000
1!
1*
b111 6
19
1>
1C
b111 G
#116840000000
0!
0*
09
0>
0C
#116850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#116860000000
0!
0*
09
0>
0C
#116870000000
1!
1*
b1 6
19
1>
1C
b1 G
#116880000000
0!
0*
09
0>
0C
#116890000000
1!
1*
b10 6
19
1>
1C
b10 G
#116900000000
0!
0*
09
0>
0C
#116910000000
1!
1*
b11 6
19
1>
1C
b11 G
#116920000000
0!
0*
09
0>
0C
#116930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#116940000000
0!
0*
09
0>
0C
#116950000000
1!
1*
b101 6
19
1>
1C
b101 G
#116960000000
0!
0*
09
0>
0C
#116970000000
1!
1*
b110 6
19
1>
1C
b110 G
#116980000000
0!
0*
09
0>
0C
#116990000000
1!
1*
b111 6
19
1>
1C
b111 G
#117000000000
0!
1"
0*
1+
09
1:
0>
0C
#117010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#117020000000
0!
0*
09
0>
0C
#117030000000
1!
1*
b1 6
19
1>
1C
b1 G
#117040000000
0!
0*
09
0>
0C
#117050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#117060000000
0!
0*
09
0>
0C
#117070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#117080000000
0!
0*
09
0>
0C
#117090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#117100000000
0!
0*
09
0>
0C
#117110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#117120000000
0!
0#
0*
0,
09
0>
0?
0C
#117130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#117140000000
0!
0*
09
0>
0C
#117150000000
1!
1*
19
1>
1C
#117160000000
0!
0*
09
0>
0C
#117170000000
1!
1*
19
1>
1C
#117180000000
0!
0*
09
0>
0C
#117190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#117200000000
0!
0*
09
0>
0C
#117210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#117220000000
0!
0*
09
0>
0C
#117230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#117240000000
0!
0*
09
0>
0C
#117250000000
1!
1*
b10 6
19
1>
1C
b10 G
#117260000000
0!
0*
09
0>
0C
#117270000000
1!
1*
b11 6
19
1>
1C
b11 G
#117280000000
0!
0*
09
0>
0C
#117290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#117300000000
0!
0*
09
0>
0C
#117310000000
1!
1*
b101 6
19
1>
1C
b101 G
#117320000000
0!
0*
09
0>
0C
#117330000000
1!
1*
b110 6
19
1>
1C
b110 G
#117340000000
0!
0*
09
0>
0C
#117350000000
1!
1*
b111 6
19
1>
1C
b111 G
#117360000000
0!
0*
09
0>
0C
#117370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#117380000000
0!
0*
09
0>
0C
#117390000000
1!
1*
b1 6
19
1>
1C
b1 G
#117400000000
0!
0*
09
0>
0C
#117410000000
1!
1*
b10 6
19
1>
1C
b10 G
#117420000000
0!
0*
09
0>
0C
#117430000000
1!
1*
b11 6
19
1>
1C
b11 G
#117440000000
0!
0*
09
0>
0C
#117450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#117460000000
0!
0*
09
0>
0C
#117470000000
1!
1*
b101 6
19
1>
1C
b101 G
#117480000000
0!
0*
09
0>
0C
#117490000000
1!
1*
b110 6
19
1>
1C
b110 G
#117500000000
0!
0*
09
0>
0C
#117510000000
1!
1*
b111 6
19
1>
1C
b111 G
#117520000000
0!
0*
09
0>
0C
#117530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#117540000000
0!
0*
09
0>
0C
#117550000000
1!
1*
b1 6
19
1>
1C
b1 G
#117560000000
0!
0*
09
0>
0C
#117570000000
1!
1*
b10 6
19
1>
1C
b10 G
#117580000000
0!
0*
09
0>
0C
#117590000000
1!
1*
b11 6
19
1>
1C
b11 G
#117600000000
0!
0*
09
0>
0C
#117610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#117620000000
0!
0*
09
0>
0C
#117630000000
1!
1*
b101 6
19
1>
1C
b101 G
#117640000000
0!
0*
09
0>
0C
#117650000000
1!
1*
b110 6
19
1>
1C
b110 G
#117660000000
0!
0*
09
0>
0C
#117670000000
1!
1*
b111 6
19
1>
1C
b111 G
#117680000000
0!
1"
0*
1+
09
1:
0>
0C
#117690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#117700000000
0!
0*
09
0>
0C
#117710000000
1!
1*
b1 6
19
1>
1C
b1 G
#117720000000
0!
0*
09
0>
0C
#117730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#117740000000
0!
0*
09
0>
0C
#117750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#117760000000
0!
0*
09
0>
0C
#117770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#117780000000
0!
0*
09
0>
0C
#117790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#117800000000
0!
0#
0*
0,
09
0>
0?
0C
#117810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#117820000000
0!
0*
09
0>
0C
#117830000000
1!
1*
19
1>
1C
#117840000000
0!
0*
09
0>
0C
#117850000000
1!
1*
19
1>
1C
#117860000000
0!
0*
09
0>
0C
#117870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#117880000000
0!
0*
09
0>
0C
#117890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#117900000000
0!
0*
09
0>
0C
#117910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#117920000000
0!
0*
09
0>
0C
#117930000000
1!
1*
b10 6
19
1>
1C
b10 G
#117940000000
0!
0*
09
0>
0C
#117950000000
1!
1*
b11 6
19
1>
1C
b11 G
#117960000000
0!
0*
09
0>
0C
#117970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#117980000000
0!
0*
09
0>
0C
#117990000000
1!
1*
b101 6
19
1>
1C
b101 G
#118000000000
0!
0*
09
0>
0C
#118010000000
1!
1*
b110 6
19
1>
1C
b110 G
#118020000000
0!
0*
09
0>
0C
#118030000000
1!
1*
b111 6
19
1>
1C
b111 G
#118040000000
0!
0*
09
0>
0C
#118050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#118060000000
0!
0*
09
0>
0C
#118070000000
1!
1*
b1 6
19
1>
1C
b1 G
#118080000000
0!
0*
09
0>
0C
#118090000000
1!
1*
b10 6
19
1>
1C
b10 G
#118100000000
0!
0*
09
0>
0C
#118110000000
1!
1*
b11 6
19
1>
1C
b11 G
#118120000000
0!
0*
09
0>
0C
#118130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#118140000000
0!
0*
09
0>
0C
#118150000000
1!
1*
b101 6
19
1>
1C
b101 G
#118160000000
0!
0*
09
0>
0C
#118170000000
1!
1*
b110 6
19
1>
1C
b110 G
#118180000000
0!
0*
09
0>
0C
#118190000000
1!
1*
b111 6
19
1>
1C
b111 G
#118200000000
0!
0*
09
0>
0C
#118210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#118220000000
0!
0*
09
0>
0C
#118230000000
1!
1*
b1 6
19
1>
1C
b1 G
#118240000000
0!
0*
09
0>
0C
#118250000000
1!
1*
b10 6
19
1>
1C
b10 G
#118260000000
0!
0*
09
0>
0C
#118270000000
1!
1*
b11 6
19
1>
1C
b11 G
#118280000000
0!
0*
09
0>
0C
#118290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#118300000000
0!
0*
09
0>
0C
#118310000000
1!
1*
b101 6
19
1>
1C
b101 G
#118320000000
0!
0*
09
0>
0C
#118330000000
1!
1*
b110 6
19
1>
1C
b110 G
#118340000000
0!
0*
09
0>
0C
#118350000000
1!
1*
b111 6
19
1>
1C
b111 G
#118360000000
0!
1"
0*
1+
09
1:
0>
0C
#118370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#118380000000
0!
0*
09
0>
0C
#118390000000
1!
1*
b1 6
19
1>
1C
b1 G
#118400000000
0!
0*
09
0>
0C
#118410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#118420000000
0!
0*
09
0>
0C
#118430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#118440000000
0!
0*
09
0>
0C
#118450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#118460000000
0!
0*
09
0>
0C
#118470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#118480000000
0!
0#
0*
0,
09
0>
0?
0C
#118490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#118500000000
0!
0*
09
0>
0C
#118510000000
1!
1*
19
1>
1C
#118520000000
0!
0*
09
0>
0C
#118530000000
1!
1*
19
1>
1C
#118540000000
0!
0*
09
0>
0C
#118550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#118560000000
0!
0*
09
0>
0C
#118570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#118580000000
0!
0*
09
0>
0C
#118590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#118600000000
0!
0*
09
0>
0C
#118610000000
1!
1*
b10 6
19
1>
1C
b10 G
#118620000000
0!
0*
09
0>
0C
#118630000000
1!
1*
b11 6
19
1>
1C
b11 G
#118640000000
0!
0*
09
0>
0C
#118650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#118660000000
0!
0*
09
0>
0C
#118670000000
1!
1*
b101 6
19
1>
1C
b101 G
#118680000000
0!
0*
09
0>
0C
#118690000000
1!
1*
b110 6
19
1>
1C
b110 G
#118700000000
0!
0*
09
0>
0C
#118710000000
1!
1*
b111 6
19
1>
1C
b111 G
#118720000000
0!
0*
09
0>
0C
#118730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#118740000000
0!
0*
09
0>
0C
#118750000000
1!
1*
b1 6
19
1>
1C
b1 G
#118760000000
0!
0*
09
0>
0C
#118770000000
1!
1*
b10 6
19
1>
1C
b10 G
#118780000000
0!
0*
09
0>
0C
#118790000000
1!
1*
b11 6
19
1>
1C
b11 G
#118800000000
0!
0*
09
0>
0C
#118810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#118820000000
0!
0*
09
0>
0C
#118830000000
1!
1*
b101 6
19
1>
1C
b101 G
#118840000000
0!
0*
09
0>
0C
#118850000000
1!
1*
b110 6
19
1>
1C
b110 G
#118860000000
0!
0*
09
0>
0C
#118870000000
1!
1*
b111 6
19
1>
1C
b111 G
#118880000000
0!
0*
09
0>
0C
#118890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#118900000000
0!
0*
09
0>
0C
#118910000000
1!
1*
b1 6
19
1>
1C
b1 G
#118920000000
0!
0*
09
0>
0C
#118930000000
1!
1*
b10 6
19
1>
1C
b10 G
#118940000000
0!
0*
09
0>
0C
#118950000000
1!
1*
b11 6
19
1>
1C
b11 G
#118960000000
0!
0*
09
0>
0C
#118970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#118980000000
0!
0*
09
0>
0C
#118990000000
1!
1*
b101 6
19
1>
1C
b101 G
#119000000000
0!
0*
09
0>
0C
#119010000000
1!
1*
b110 6
19
1>
1C
b110 G
#119020000000
0!
0*
09
0>
0C
#119030000000
1!
1*
b111 6
19
1>
1C
b111 G
#119040000000
0!
1"
0*
1+
09
1:
0>
0C
#119050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#119060000000
0!
0*
09
0>
0C
#119070000000
1!
1*
b1 6
19
1>
1C
b1 G
#119080000000
0!
0*
09
0>
0C
#119090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#119100000000
0!
0*
09
0>
0C
#119110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#119120000000
0!
0*
09
0>
0C
#119130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#119140000000
0!
0*
09
0>
0C
#119150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#119160000000
0!
0#
0*
0,
09
0>
0?
0C
#119170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#119180000000
0!
0*
09
0>
0C
#119190000000
1!
1*
19
1>
1C
#119200000000
0!
0*
09
0>
0C
#119210000000
1!
1*
19
1>
1C
#119220000000
0!
0*
09
0>
0C
#119230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#119240000000
0!
0*
09
0>
0C
#119250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#119260000000
0!
0*
09
0>
0C
#119270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#119280000000
0!
0*
09
0>
0C
#119290000000
1!
1*
b10 6
19
1>
1C
b10 G
#119300000000
0!
0*
09
0>
0C
#119310000000
1!
1*
b11 6
19
1>
1C
b11 G
#119320000000
0!
0*
09
0>
0C
#119330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#119340000000
0!
0*
09
0>
0C
#119350000000
1!
1*
b101 6
19
1>
1C
b101 G
#119360000000
0!
0*
09
0>
0C
#119370000000
1!
1*
b110 6
19
1>
1C
b110 G
#119380000000
0!
0*
09
0>
0C
#119390000000
1!
1*
b111 6
19
1>
1C
b111 G
#119400000000
0!
0*
09
0>
0C
#119410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#119420000000
0!
0*
09
0>
0C
#119430000000
1!
1*
b1 6
19
1>
1C
b1 G
#119440000000
0!
0*
09
0>
0C
#119450000000
1!
1*
b10 6
19
1>
1C
b10 G
#119460000000
0!
0*
09
0>
0C
#119470000000
1!
1*
b11 6
19
1>
1C
b11 G
#119480000000
0!
0*
09
0>
0C
#119490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#119500000000
0!
0*
09
0>
0C
#119510000000
1!
1*
b101 6
19
1>
1C
b101 G
#119520000000
0!
0*
09
0>
0C
#119530000000
1!
1*
b110 6
19
1>
1C
b110 G
#119540000000
0!
0*
09
0>
0C
#119550000000
1!
1*
b111 6
19
1>
1C
b111 G
#119560000000
0!
0*
09
0>
0C
#119570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#119580000000
0!
0*
09
0>
0C
#119590000000
1!
1*
b1 6
19
1>
1C
b1 G
#119600000000
0!
0*
09
0>
0C
#119610000000
1!
1*
b10 6
19
1>
1C
b10 G
#119620000000
0!
0*
09
0>
0C
#119630000000
1!
1*
b11 6
19
1>
1C
b11 G
#119640000000
0!
0*
09
0>
0C
#119650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#119660000000
0!
0*
09
0>
0C
#119670000000
1!
1*
b101 6
19
1>
1C
b101 G
#119680000000
0!
0*
09
0>
0C
#119690000000
1!
1*
b110 6
19
1>
1C
b110 G
#119700000000
0!
0*
09
0>
0C
#119710000000
1!
1*
b111 6
19
1>
1C
b111 G
#119720000000
0!
1"
0*
1+
09
1:
0>
0C
#119730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#119740000000
0!
0*
09
0>
0C
#119750000000
1!
1*
b1 6
19
1>
1C
b1 G
#119760000000
0!
0*
09
0>
0C
#119770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#119780000000
0!
0*
09
0>
0C
#119790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#119800000000
0!
0*
09
0>
0C
#119810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#119820000000
0!
0*
09
0>
0C
#119830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#119840000000
0!
0#
0*
0,
09
0>
0?
0C
#119850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#119860000000
0!
0*
09
0>
0C
#119870000000
1!
1*
19
1>
1C
#119880000000
0!
0*
09
0>
0C
#119890000000
1!
1*
19
1>
1C
#119900000000
0!
0*
09
0>
0C
#119910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#119920000000
0!
0*
09
0>
0C
#119930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#119940000000
0!
0*
09
0>
0C
#119950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#119960000000
0!
0*
09
0>
0C
#119970000000
1!
1*
b10 6
19
1>
1C
b10 G
#119980000000
0!
0*
09
0>
0C
#119990000000
1!
1*
b11 6
19
1>
1C
b11 G
#120000000000
0!
0*
09
0>
0C
#120010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#120020000000
0!
0*
09
0>
0C
#120030000000
1!
1*
b101 6
19
1>
1C
b101 G
#120040000000
0!
0*
09
0>
0C
#120050000000
1!
1*
b110 6
19
1>
1C
b110 G
#120060000000
0!
0*
09
0>
0C
#120070000000
1!
1*
b111 6
19
1>
1C
b111 G
#120080000000
0!
0*
09
0>
0C
#120090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#120100000000
0!
0*
09
0>
0C
#120110000000
1!
1*
b1 6
19
1>
1C
b1 G
#120120000000
0!
0*
09
0>
0C
#120130000000
1!
1*
b10 6
19
1>
1C
b10 G
#120140000000
0!
0*
09
0>
0C
#120150000000
1!
1*
b11 6
19
1>
1C
b11 G
#120160000000
0!
0*
09
0>
0C
#120170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#120180000000
0!
0*
09
0>
0C
#120190000000
1!
1*
b101 6
19
1>
1C
b101 G
#120200000000
0!
0*
09
0>
0C
#120210000000
1!
1*
b110 6
19
1>
1C
b110 G
#120220000000
0!
0*
09
0>
0C
#120230000000
1!
1*
b111 6
19
1>
1C
b111 G
#120240000000
0!
0*
09
0>
0C
#120250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#120260000000
0!
0*
09
0>
0C
#120270000000
1!
1*
b1 6
19
1>
1C
b1 G
#120280000000
0!
0*
09
0>
0C
#120290000000
1!
1*
b10 6
19
1>
1C
b10 G
#120300000000
0!
0*
09
0>
0C
#120310000000
1!
1*
b11 6
19
1>
1C
b11 G
#120320000000
0!
0*
09
0>
0C
#120330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#120340000000
0!
0*
09
0>
0C
#120350000000
1!
1*
b101 6
19
1>
1C
b101 G
#120360000000
0!
0*
09
0>
0C
#120370000000
1!
1*
b110 6
19
1>
1C
b110 G
#120380000000
0!
0*
09
0>
0C
#120390000000
1!
1*
b111 6
19
1>
1C
b111 G
#120400000000
0!
1"
0*
1+
09
1:
0>
0C
#120410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#120420000000
0!
0*
09
0>
0C
#120430000000
1!
1*
b1 6
19
1>
1C
b1 G
#120440000000
0!
0*
09
0>
0C
#120450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#120460000000
0!
0*
09
0>
0C
#120470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#120480000000
0!
0*
09
0>
0C
#120490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#120500000000
0!
0*
09
0>
0C
#120510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#120520000000
0!
0#
0*
0,
09
0>
0?
0C
#120530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#120540000000
0!
0*
09
0>
0C
#120550000000
1!
1*
19
1>
1C
#120560000000
0!
0*
09
0>
0C
#120570000000
1!
1*
19
1>
1C
#120580000000
0!
0*
09
0>
0C
#120590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#120600000000
0!
0*
09
0>
0C
#120610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#120620000000
0!
0*
09
0>
0C
#120630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#120640000000
0!
0*
09
0>
0C
#120650000000
1!
1*
b10 6
19
1>
1C
b10 G
#120660000000
0!
0*
09
0>
0C
#120670000000
1!
1*
b11 6
19
1>
1C
b11 G
#120680000000
0!
0*
09
0>
0C
#120690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#120700000000
0!
0*
09
0>
0C
#120710000000
1!
1*
b101 6
19
1>
1C
b101 G
#120720000000
0!
0*
09
0>
0C
#120730000000
1!
1*
b110 6
19
1>
1C
b110 G
#120740000000
0!
0*
09
0>
0C
#120750000000
1!
1*
b111 6
19
1>
1C
b111 G
#120760000000
0!
0*
09
0>
0C
#120770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#120780000000
0!
0*
09
0>
0C
#120790000000
1!
1*
b1 6
19
1>
1C
b1 G
#120800000000
0!
0*
09
0>
0C
#120810000000
1!
1*
b10 6
19
1>
1C
b10 G
#120820000000
0!
0*
09
0>
0C
#120830000000
1!
1*
b11 6
19
1>
1C
b11 G
#120840000000
0!
0*
09
0>
0C
#120850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#120860000000
0!
0*
09
0>
0C
#120870000000
1!
1*
b101 6
19
1>
1C
b101 G
#120880000000
0!
0*
09
0>
0C
#120890000000
1!
1*
b110 6
19
1>
1C
b110 G
#120900000000
0!
0*
09
0>
0C
#120910000000
1!
1*
b111 6
19
1>
1C
b111 G
#120920000000
0!
0*
09
0>
0C
#120930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#120940000000
0!
0*
09
0>
0C
#120950000000
1!
1*
b1 6
19
1>
1C
b1 G
#120960000000
0!
0*
09
0>
0C
#120970000000
1!
1*
b10 6
19
1>
1C
b10 G
#120980000000
0!
0*
09
0>
0C
#120990000000
1!
1*
b11 6
19
1>
1C
b11 G
#121000000000
0!
0*
09
0>
0C
#121010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#121020000000
0!
0*
09
0>
0C
#121030000000
1!
1*
b101 6
19
1>
1C
b101 G
#121040000000
0!
0*
09
0>
0C
#121050000000
1!
1*
b110 6
19
1>
1C
b110 G
#121060000000
0!
0*
09
0>
0C
#121070000000
1!
1*
b111 6
19
1>
1C
b111 G
#121080000000
0!
1"
0*
1+
09
1:
0>
0C
#121090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#121100000000
0!
0*
09
0>
0C
#121110000000
1!
1*
b1 6
19
1>
1C
b1 G
#121120000000
0!
0*
09
0>
0C
#121130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#121140000000
0!
0*
09
0>
0C
#121150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#121160000000
0!
0*
09
0>
0C
#121170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#121180000000
0!
0*
09
0>
0C
#121190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#121200000000
0!
0#
0*
0,
09
0>
0?
0C
#121210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#121220000000
0!
0*
09
0>
0C
#121230000000
1!
1*
19
1>
1C
#121240000000
0!
0*
09
0>
0C
#121250000000
1!
1*
19
1>
1C
#121260000000
0!
0*
09
0>
0C
#121270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#121280000000
0!
0*
09
0>
0C
#121290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#121300000000
0!
0*
09
0>
0C
#121310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#121320000000
0!
0*
09
0>
0C
#121330000000
1!
1*
b10 6
19
1>
1C
b10 G
#121340000000
0!
0*
09
0>
0C
#121350000000
1!
1*
b11 6
19
1>
1C
b11 G
#121360000000
0!
0*
09
0>
0C
#121370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#121380000000
0!
0*
09
0>
0C
#121390000000
1!
1*
b101 6
19
1>
1C
b101 G
#121400000000
0!
0*
09
0>
0C
#121410000000
1!
1*
b110 6
19
1>
1C
b110 G
#121420000000
0!
0*
09
0>
0C
#121430000000
1!
1*
b111 6
19
1>
1C
b111 G
#121440000000
0!
0*
09
0>
0C
#121450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#121460000000
0!
0*
09
0>
0C
#121470000000
1!
1*
b1 6
19
1>
1C
b1 G
#121480000000
0!
0*
09
0>
0C
#121490000000
1!
1*
b10 6
19
1>
1C
b10 G
#121500000000
0!
0*
09
0>
0C
#121510000000
1!
1*
b11 6
19
1>
1C
b11 G
#121520000000
0!
0*
09
0>
0C
#121530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#121540000000
0!
0*
09
0>
0C
#121550000000
1!
1*
b101 6
19
1>
1C
b101 G
#121560000000
0!
0*
09
0>
0C
#121570000000
1!
1*
b110 6
19
1>
1C
b110 G
#121580000000
0!
0*
09
0>
0C
#121590000000
1!
1*
b111 6
19
1>
1C
b111 G
#121600000000
0!
0*
09
0>
0C
#121610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#121620000000
0!
0*
09
0>
0C
#121630000000
1!
1*
b1 6
19
1>
1C
b1 G
#121640000000
0!
0*
09
0>
0C
#121650000000
1!
1*
b10 6
19
1>
1C
b10 G
#121660000000
0!
0*
09
0>
0C
#121670000000
1!
1*
b11 6
19
1>
1C
b11 G
#121680000000
0!
0*
09
0>
0C
#121690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#121700000000
0!
0*
09
0>
0C
#121710000000
1!
1*
b101 6
19
1>
1C
b101 G
#121720000000
0!
0*
09
0>
0C
#121730000000
1!
1*
b110 6
19
1>
1C
b110 G
#121740000000
0!
0*
09
0>
0C
#121750000000
1!
1*
b111 6
19
1>
1C
b111 G
#121760000000
0!
1"
0*
1+
09
1:
0>
0C
#121770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#121780000000
0!
0*
09
0>
0C
#121790000000
1!
1*
b1 6
19
1>
1C
b1 G
#121800000000
0!
0*
09
0>
0C
#121810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#121820000000
0!
0*
09
0>
0C
#121830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#121840000000
0!
0*
09
0>
0C
#121850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#121860000000
0!
0*
09
0>
0C
#121870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#121880000000
0!
0#
0*
0,
09
0>
0?
0C
#121890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#121900000000
0!
0*
09
0>
0C
#121910000000
1!
1*
19
1>
1C
#121920000000
0!
0*
09
0>
0C
#121930000000
1!
1*
19
1>
1C
#121940000000
0!
0*
09
0>
0C
#121950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#121960000000
0!
0*
09
0>
0C
#121970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#121980000000
0!
0*
09
0>
0C
#121990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#122000000000
0!
0*
09
0>
0C
#122010000000
1!
1*
b10 6
19
1>
1C
b10 G
#122020000000
0!
0*
09
0>
0C
#122030000000
1!
1*
b11 6
19
1>
1C
b11 G
#122040000000
0!
0*
09
0>
0C
#122050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#122060000000
0!
0*
09
0>
0C
#122070000000
1!
1*
b101 6
19
1>
1C
b101 G
#122080000000
0!
0*
09
0>
0C
#122090000000
1!
1*
b110 6
19
1>
1C
b110 G
#122100000000
0!
0*
09
0>
0C
#122110000000
1!
1*
b111 6
19
1>
1C
b111 G
#122120000000
0!
0*
09
0>
0C
#122130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#122140000000
0!
0*
09
0>
0C
#122150000000
1!
1*
b1 6
19
1>
1C
b1 G
#122160000000
0!
0*
09
0>
0C
#122170000000
1!
1*
b10 6
19
1>
1C
b10 G
#122180000000
0!
0*
09
0>
0C
#122190000000
1!
1*
b11 6
19
1>
1C
b11 G
#122200000000
0!
0*
09
0>
0C
#122210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#122220000000
0!
0*
09
0>
0C
#122230000000
1!
1*
b101 6
19
1>
1C
b101 G
#122240000000
0!
0*
09
0>
0C
#122250000000
1!
1*
b110 6
19
1>
1C
b110 G
#122260000000
0!
0*
09
0>
0C
#122270000000
1!
1*
b111 6
19
1>
1C
b111 G
#122280000000
0!
0*
09
0>
0C
#122290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#122300000000
0!
0*
09
0>
0C
#122310000000
1!
1*
b1 6
19
1>
1C
b1 G
#122320000000
0!
0*
09
0>
0C
#122330000000
1!
1*
b10 6
19
1>
1C
b10 G
#122340000000
0!
0*
09
0>
0C
#122350000000
1!
1*
b11 6
19
1>
1C
b11 G
#122360000000
0!
0*
09
0>
0C
#122370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#122380000000
0!
0*
09
0>
0C
#122390000000
1!
1*
b101 6
19
1>
1C
b101 G
#122400000000
0!
0*
09
0>
0C
#122410000000
1!
1*
b110 6
19
1>
1C
b110 G
#122420000000
0!
0*
09
0>
0C
#122430000000
1!
1*
b111 6
19
1>
1C
b111 G
#122440000000
0!
1"
0*
1+
09
1:
0>
0C
#122450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#122460000000
0!
0*
09
0>
0C
#122470000000
1!
1*
b1 6
19
1>
1C
b1 G
#122480000000
0!
0*
09
0>
0C
#122490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#122500000000
0!
0*
09
0>
0C
#122510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#122520000000
0!
0*
09
0>
0C
#122530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#122540000000
0!
0*
09
0>
0C
#122550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#122560000000
0!
0#
0*
0,
09
0>
0?
0C
#122570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#122580000000
0!
0*
09
0>
0C
#122590000000
1!
1*
19
1>
1C
#122600000000
0!
0*
09
0>
0C
#122610000000
1!
1*
19
1>
1C
#122620000000
0!
0*
09
0>
0C
#122630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#122640000000
0!
0*
09
0>
0C
#122650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#122660000000
0!
0*
09
0>
0C
#122670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#122680000000
0!
0*
09
0>
0C
#122690000000
1!
1*
b10 6
19
1>
1C
b10 G
#122700000000
0!
0*
09
0>
0C
#122710000000
1!
1*
b11 6
19
1>
1C
b11 G
#122720000000
0!
0*
09
0>
0C
#122730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#122740000000
0!
0*
09
0>
0C
#122750000000
1!
1*
b101 6
19
1>
1C
b101 G
#122760000000
0!
0*
09
0>
0C
#122770000000
1!
1*
b110 6
19
1>
1C
b110 G
#122780000000
0!
0*
09
0>
0C
#122790000000
1!
1*
b111 6
19
1>
1C
b111 G
#122800000000
0!
0*
09
0>
0C
#122810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#122820000000
0!
0*
09
0>
0C
#122830000000
1!
1*
b1 6
19
1>
1C
b1 G
#122840000000
0!
0*
09
0>
0C
#122850000000
1!
1*
b10 6
19
1>
1C
b10 G
#122860000000
0!
0*
09
0>
0C
#122870000000
1!
1*
b11 6
19
1>
1C
b11 G
#122880000000
0!
0*
09
0>
0C
#122890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#122900000000
0!
0*
09
0>
0C
#122910000000
1!
1*
b101 6
19
1>
1C
b101 G
#122920000000
0!
0*
09
0>
0C
#122930000000
1!
1*
b110 6
19
1>
1C
b110 G
#122940000000
0!
0*
09
0>
0C
#122950000000
1!
1*
b111 6
19
1>
1C
b111 G
#122960000000
0!
0*
09
0>
0C
#122970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#122980000000
0!
0*
09
0>
0C
#122990000000
1!
1*
b1 6
19
1>
1C
b1 G
#123000000000
0!
0*
09
0>
0C
#123010000000
1!
1*
b10 6
19
1>
1C
b10 G
#123020000000
0!
0*
09
0>
0C
#123030000000
1!
1*
b11 6
19
1>
1C
b11 G
#123040000000
0!
0*
09
0>
0C
#123050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#123060000000
0!
0*
09
0>
0C
#123070000000
1!
1*
b101 6
19
1>
1C
b101 G
#123080000000
0!
0*
09
0>
0C
#123090000000
1!
1*
b110 6
19
1>
1C
b110 G
#123100000000
0!
0*
09
0>
0C
#123110000000
1!
1*
b111 6
19
1>
1C
b111 G
#123120000000
0!
1"
0*
1+
09
1:
0>
0C
#123130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#123140000000
0!
0*
09
0>
0C
#123150000000
1!
1*
b1 6
19
1>
1C
b1 G
#123160000000
0!
0*
09
0>
0C
#123170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#123180000000
0!
0*
09
0>
0C
#123190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#123200000000
0!
0*
09
0>
0C
#123210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#123220000000
0!
0*
09
0>
0C
#123230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#123240000000
0!
0#
0*
0,
09
0>
0?
0C
#123250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#123260000000
0!
0*
09
0>
0C
#123270000000
1!
1*
19
1>
1C
#123280000000
0!
0*
09
0>
0C
#123290000000
1!
1*
19
1>
1C
#123300000000
0!
0*
09
0>
0C
#123310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#123320000000
0!
0*
09
0>
0C
#123330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#123340000000
0!
0*
09
0>
0C
#123350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#123360000000
0!
0*
09
0>
0C
#123370000000
1!
1*
b10 6
19
1>
1C
b10 G
#123380000000
0!
0*
09
0>
0C
#123390000000
1!
1*
b11 6
19
1>
1C
b11 G
#123400000000
0!
0*
09
0>
0C
#123410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#123420000000
0!
0*
09
0>
0C
#123430000000
1!
1*
b101 6
19
1>
1C
b101 G
#123440000000
0!
0*
09
0>
0C
#123450000000
1!
1*
b110 6
19
1>
1C
b110 G
#123460000000
0!
0*
09
0>
0C
#123470000000
1!
1*
b111 6
19
1>
1C
b111 G
#123480000000
0!
0*
09
0>
0C
#123490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#123500000000
0!
0*
09
0>
0C
#123510000000
1!
1*
b1 6
19
1>
1C
b1 G
#123520000000
0!
0*
09
0>
0C
#123530000000
1!
1*
b10 6
19
1>
1C
b10 G
#123540000000
0!
0*
09
0>
0C
#123550000000
1!
1*
b11 6
19
1>
1C
b11 G
#123560000000
0!
0*
09
0>
0C
#123570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#123580000000
0!
0*
09
0>
0C
#123590000000
1!
1*
b101 6
19
1>
1C
b101 G
#123600000000
0!
0*
09
0>
0C
#123610000000
1!
1*
b110 6
19
1>
1C
b110 G
#123620000000
0!
0*
09
0>
0C
#123630000000
1!
1*
b111 6
19
1>
1C
b111 G
#123640000000
0!
0*
09
0>
0C
#123650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#123660000000
0!
0*
09
0>
0C
#123670000000
1!
1*
b1 6
19
1>
1C
b1 G
#123680000000
0!
0*
09
0>
0C
#123690000000
1!
1*
b10 6
19
1>
1C
b10 G
#123700000000
0!
0*
09
0>
0C
#123710000000
1!
1*
b11 6
19
1>
1C
b11 G
#123720000000
0!
0*
09
0>
0C
#123730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#123740000000
0!
0*
09
0>
0C
#123750000000
1!
1*
b101 6
19
1>
1C
b101 G
#123760000000
0!
0*
09
0>
0C
#123770000000
1!
1*
b110 6
19
1>
1C
b110 G
#123780000000
0!
0*
09
0>
0C
#123790000000
1!
1*
b111 6
19
1>
1C
b111 G
#123800000000
0!
1"
0*
1+
09
1:
0>
0C
#123810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#123820000000
0!
0*
09
0>
0C
#123830000000
1!
1*
b1 6
19
1>
1C
b1 G
#123840000000
0!
0*
09
0>
0C
#123850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#123860000000
0!
0*
09
0>
0C
#123870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#123880000000
0!
0*
09
0>
0C
#123890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#123900000000
0!
0*
09
0>
0C
#123910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#123920000000
0!
0#
0*
0,
09
0>
0?
0C
#123930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#123940000000
0!
0*
09
0>
0C
#123950000000
1!
1*
19
1>
1C
#123960000000
0!
0*
09
0>
0C
#123970000000
1!
1*
19
1>
1C
#123980000000
0!
0*
09
0>
0C
#123990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#124000000000
0!
0*
09
0>
0C
#124010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#124020000000
0!
0*
09
0>
0C
#124030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#124040000000
0!
0*
09
0>
0C
#124050000000
1!
1*
b10 6
19
1>
1C
b10 G
#124060000000
0!
0*
09
0>
0C
#124070000000
1!
1*
b11 6
19
1>
1C
b11 G
#124080000000
0!
0*
09
0>
0C
#124090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#124100000000
0!
0*
09
0>
0C
#124110000000
1!
1*
b101 6
19
1>
1C
b101 G
#124120000000
0!
0*
09
0>
0C
#124130000000
1!
1*
b110 6
19
1>
1C
b110 G
#124140000000
0!
0*
09
0>
0C
#124150000000
1!
1*
b111 6
19
1>
1C
b111 G
#124160000000
0!
0*
09
0>
0C
#124170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#124180000000
0!
0*
09
0>
0C
#124190000000
1!
1*
b1 6
19
1>
1C
b1 G
#124200000000
0!
0*
09
0>
0C
#124210000000
1!
1*
b10 6
19
1>
1C
b10 G
#124220000000
0!
0*
09
0>
0C
#124230000000
1!
1*
b11 6
19
1>
1C
b11 G
#124240000000
0!
0*
09
0>
0C
#124250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#124260000000
0!
0*
09
0>
0C
#124270000000
1!
1*
b101 6
19
1>
1C
b101 G
#124280000000
0!
0*
09
0>
0C
#124290000000
1!
1*
b110 6
19
1>
1C
b110 G
#124300000000
0!
0*
09
0>
0C
#124310000000
1!
1*
b111 6
19
1>
1C
b111 G
#124320000000
0!
0*
09
0>
0C
#124330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#124340000000
0!
0*
09
0>
0C
#124350000000
1!
1*
b1 6
19
1>
1C
b1 G
#124360000000
0!
0*
09
0>
0C
#124370000000
1!
1*
b10 6
19
1>
1C
b10 G
#124380000000
0!
0*
09
0>
0C
#124390000000
1!
1*
b11 6
19
1>
1C
b11 G
#124400000000
0!
0*
09
0>
0C
#124410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#124420000000
0!
0*
09
0>
0C
#124430000000
1!
1*
b101 6
19
1>
1C
b101 G
#124440000000
0!
0*
09
0>
0C
#124450000000
1!
1*
b110 6
19
1>
1C
b110 G
#124460000000
0!
0*
09
0>
0C
#124470000000
1!
1*
b111 6
19
1>
1C
b111 G
#124480000000
0!
1"
0*
1+
09
1:
0>
0C
#124490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#124500000000
0!
0*
09
0>
0C
#124510000000
1!
1*
b1 6
19
1>
1C
b1 G
#124520000000
0!
0*
09
0>
0C
#124530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#124540000000
0!
0*
09
0>
0C
#124550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#124560000000
0!
0*
09
0>
0C
#124570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#124580000000
0!
0*
09
0>
0C
#124590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#124600000000
0!
0#
0*
0,
09
0>
0?
0C
#124610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#124620000000
0!
0*
09
0>
0C
#124630000000
1!
1*
19
1>
1C
#124640000000
0!
0*
09
0>
0C
#124650000000
1!
1*
19
1>
1C
#124660000000
0!
0*
09
0>
0C
#124670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#124680000000
0!
0*
09
0>
0C
#124690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#124700000000
0!
0*
09
0>
0C
#124710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#124720000000
0!
0*
09
0>
0C
#124730000000
1!
1*
b10 6
19
1>
1C
b10 G
#124740000000
0!
0*
09
0>
0C
#124750000000
1!
1*
b11 6
19
1>
1C
b11 G
#124760000000
0!
0*
09
0>
0C
#124770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#124780000000
0!
0*
09
0>
0C
#124790000000
1!
1*
b101 6
19
1>
1C
b101 G
#124800000000
0!
0*
09
0>
0C
#124810000000
1!
1*
b110 6
19
1>
1C
b110 G
#124820000000
0!
0*
09
0>
0C
#124830000000
1!
1*
b111 6
19
1>
1C
b111 G
#124840000000
0!
0*
09
0>
0C
#124850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#124860000000
0!
0*
09
0>
0C
#124870000000
1!
1*
b1 6
19
1>
1C
b1 G
#124880000000
0!
0*
09
0>
0C
#124890000000
1!
1*
b10 6
19
1>
1C
b10 G
#124900000000
0!
0*
09
0>
0C
#124910000000
1!
1*
b11 6
19
1>
1C
b11 G
#124920000000
0!
0*
09
0>
0C
#124930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#124940000000
0!
0*
09
0>
0C
#124950000000
1!
1*
b101 6
19
1>
1C
b101 G
#124960000000
0!
0*
09
0>
0C
#124970000000
1!
1*
b110 6
19
1>
1C
b110 G
#124980000000
0!
0*
09
0>
0C
#124990000000
1!
1*
b111 6
19
1>
1C
b111 G
#125000000000
0!
0*
09
0>
0C
#125010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#125020000000
0!
0*
09
0>
0C
#125030000000
1!
1*
b1 6
19
1>
1C
b1 G
#125040000000
0!
0*
09
0>
0C
#125050000000
1!
1*
b10 6
19
1>
1C
b10 G
#125060000000
0!
0*
09
0>
0C
#125070000000
1!
1*
b11 6
19
1>
1C
b11 G
#125080000000
0!
0*
09
0>
0C
#125090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#125100000000
0!
0*
09
0>
0C
#125110000000
1!
1*
b101 6
19
1>
1C
b101 G
#125120000000
0!
0*
09
0>
0C
#125130000000
1!
1*
b110 6
19
1>
1C
b110 G
#125140000000
0!
0*
09
0>
0C
#125150000000
1!
1*
b111 6
19
1>
1C
b111 G
#125160000000
0!
1"
0*
1+
09
1:
0>
0C
#125170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#125180000000
0!
0*
09
0>
0C
#125190000000
1!
1*
b1 6
19
1>
1C
b1 G
#125200000000
0!
0*
09
0>
0C
#125210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#125220000000
0!
0*
09
0>
0C
#125230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#125240000000
0!
0*
09
0>
0C
#125250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#125260000000
0!
0*
09
0>
0C
#125270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#125280000000
0!
0#
0*
0,
09
0>
0?
0C
#125290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#125300000000
0!
0*
09
0>
0C
#125310000000
1!
1*
19
1>
1C
#125320000000
0!
0*
09
0>
0C
#125330000000
1!
1*
19
1>
1C
#125340000000
0!
0*
09
0>
0C
#125350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#125360000000
0!
0*
09
0>
0C
#125370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#125380000000
0!
0*
09
0>
0C
#125390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#125400000000
0!
0*
09
0>
0C
#125410000000
1!
1*
b10 6
19
1>
1C
b10 G
#125420000000
0!
0*
09
0>
0C
#125430000000
1!
1*
b11 6
19
1>
1C
b11 G
#125440000000
0!
0*
09
0>
0C
#125450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#125460000000
0!
0*
09
0>
0C
#125470000000
1!
1*
b101 6
19
1>
1C
b101 G
#125480000000
0!
0*
09
0>
0C
#125490000000
1!
1*
b110 6
19
1>
1C
b110 G
#125500000000
0!
0*
09
0>
0C
#125510000000
1!
1*
b111 6
19
1>
1C
b111 G
#125520000000
0!
0*
09
0>
0C
#125530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#125540000000
0!
0*
09
0>
0C
#125550000000
1!
1*
b1 6
19
1>
1C
b1 G
#125560000000
0!
0*
09
0>
0C
#125570000000
1!
1*
b10 6
19
1>
1C
b10 G
#125580000000
0!
0*
09
0>
0C
#125590000000
1!
1*
b11 6
19
1>
1C
b11 G
#125600000000
0!
0*
09
0>
0C
#125610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#125620000000
0!
0*
09
0>
0C
#125630000000
1!
1*
b101 6
19
1>
1C
b101 G
#125640000000
0!
0*
09
0>
0C
#125650000000
1!
1*
b110 6
19
1>
1C
b110 G
#125660000000
0!
0*
09
0>
0C
#125670000000
1!
1*
b111 6
19
1>
1C
b111 G
#125680000000
0!
0*
09
0>
0C
#125690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#125700000000
0!
0*
09
0>
0C
#125710000000
1!
1*
b1 6
19
1>
1C
b1 G
#125720000000
0!
0*
09
0>
0C
#125730000000
1!
1*
b10 6
19
1>
1C
b10 G
#125740000000
0!
0*
09
0>
0C
#125750000000
1!
1*
b11 6
19
1>
1C
b11 G
#125760000000
0!
0*
09
0>
0C
#125770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#125780000000
0!
0*
09
0>
0C
#125790000000
1!
1*
b101 6
19
1>
1C
b101 G
#125800000000
0!
0*
09
0>
0C
#125810000000
1!
1*
b110 6
19
1>
1C
b110 G
#125820000000
0!
0*
09
0>
0C
#125830000000
1!
1*
b111 6
19
1>
1C
b111 G
#125840000000
0!
1"
0*
1+
09
1:
0>
0C
#125850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#125860000000
0!
0*
09
0>
0C
#125870000000
1!
1*
b1 6
19
1>
1C
b1 G
#125880000000
0!
0*
09
0>
0C
#125890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#125900000000
0!
0*
09
0>
0C
#125910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#125920000000
0!
0*
09
0>
0C
#125930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#125940000000
0!
0*
09
0>
0C
#125950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#125960000000
0!
0#
0*
0,
09
0>
0?
0C
#125970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#125980000000
0!
0*
09
0>
0C
#125990000000
1!
1*
19
1>
1C
#126000000000
0!
0*
09
0>
0C
#126010000000
1!
1*
19
1>
1C
#126020000000
0!
0*
09
0>
0C
#126030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#126040000000
0!
0*
09
0>
0C
#126050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#126060000000
0!
0*
09
0>
0C
#126070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#126080000000
0!
0*
09
0>
0C
#126090000000
1!
1*
b10 6
19
1>
1C
b10 G
#126100000000
0!
0*
09
0>
0C
#126110000000
1!
1*
b11 6
19
1>
1C
b11 G
#126120000000
0!
0*
09
0>
0C
#126130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#126140000000
0!
0*
09
0>
0C
#126150000000
1!
1*
b101 6
19
1>
1C
b101 G
#126160000000
0!
0*
09
0>
0C
#126170000000
1!
1*
b110 6
19
1>
1C
b110 G
#126180000000
0!
0*
09
0>
0C
#126190000000
1!
1*
b111 6
19
1>
1C
b111 G
#126200000000
0!
0*
09
0>
0C
#126210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#126220000000
0!
0*
09
0>
0C
#126230000000
1!
1*
b1 6
19
1>
1C
b1 G
#126240000000
0!
0*
09
0>
0C
#126250000000
1!
1*
b10 6
19
1>
1C
b10 G
#126260000000
0!
0*
09
0>
0C
#126270000000
1!
1*
b11 6
19
1>
1C
b11 G
#126280000000
0!
0*
09
0>
0C
#126290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#126300000000
0!
0*
09
0>
0C
#126310000000
1!
1*
b101 6
19
1>
1C
b101 G
#126320000000
0!
0*
09
0>
0C
#126330000000
1!
1*
b110 6
19
1>
1C
b110 G
#126340000000
0!
0*
09
0>
0C
#126350000000
1!
1*
b111 6
19
1>
1C
b111 G
#126360000000
0!
0*
09
0>
0C
#126370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#126380000000
0!
0*
09
0>
0C
#126390000000
1!
1*
b1 6
19
1>
1C
b1 G
#126400000000
0!
0*
09
0>
0C
#126410000000
1!
1*
b10 6
19
1>
1C
b10 G
#126420000000
0!
0*
09
0>
0C
#126430000000
1!
1*
b11 6
19
1>
1C
b11 G
#126440000000
0!
0*
09
0>
0C
#126450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#126460000000
0!
0*
09
0>
0C
#126470000000
1!
1*
b101 6
19
1>
1C
b101 G
#126480000000
0!
0*
09
0>
0C
#126490000000
1!
1*
b110 6
19
1>
1C
b110 G
#126500000000
0!
0*
09
0>
0C
#126510000000
1!
1*
b111 6
19
1>
1C
b111 G
#126520000000
0!
1"
0*
1+
09
1:
0>
0C
#126530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#126540000000
0!
0*
09
0>
0C
#126550000000
1!
1*
b1 6
19
1>
1C
b1 G
#126560000000
0!
0*
09
0>
0C
#126570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#126580000000
0!
0*
09
0>
0C
#126590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#126600000000
0!
0*
09
0>
0C
#126610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#126620000000
0!
0*
09
0>
0C
#126630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#126640000000
0!
0#
0*
0,
09
0>
0?
0C
#126650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#126660000000
0!
0*
09
0>
0C
#126670000000
1!
1*
19
1>
1C
#126680000000
0!
0*
09
0>
0C
#126690000000
1!
1*
19
1>
1C
#126700000000
0!
0*
09
0>
0C
#126710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#126720000000
0!
0*
09
0>
0C
#126730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#126740000000
0!
0*
09
0>
0C
#126750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#126760000000
0!
0*
09
0>
0C
#126770000000
1!
1*
b10 6
19
1>
1C
b10 G
#126780000000
0!
0*
09
0>
0C
#126790000000
1!
1*
b11 6
19
1>
1C
b11 G
#126800000000
0!
0*
09
0>
0C
#126810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#126820000000
0!
0*
09
0>
0C
#126830000000
1!
1*
b101 6
19
1>
1C
b101 G
#126840000000
0!
0*
09
0>
0C
#126850000000
1!
1*
b110 6
19
1>
1C
b110 G
#126860000000
0!
0*
09
0>
0C
#126870000000
1!
1*
b111 6
19
1>
1C
b111 G
#126880000000
0!
0*
09
0>
0C
#126890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#126900000000
0!
0*
09
0>
0C
#126910000000
1!
1*
b1 6
19
1>
1C
b1 G
#126920000000
0!
0*
09
0>
0C
#126930000000
1!
1*
b10 6
19
1>
1C
b10 G
#126940000000
0!
0*
09
0>
0C
#126950000000
1!
1*
b11 6
19
1>
1C
b11 G
#126960000000
0!
0*
09
0>
0C
#126970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#126980000000
0!
0*
09
0>
0C
#126990000000
1!
1*
b101 6
19
1>
1C
b101 G
#127000000000
0!
0*
09
0>
0C
#127010000000
1!
1*
b110 6
19
1>
1C
b110 G
#127020000000
0!
0*
09
0>
0C
#127030000000
1!
1*
b111 6
19
1>
1C
b111 G
#127040000000
0!
0*
09
0>
0C
#127050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#127060000000
0!
0*
09
0>
0C
#127070000000
1!
1*
b1 6
19
1>
1C
b1 G
#127080000000
0!
0*
09
0>
0C
#127090000000
1!
1*
b10 6
19
1>
1C
b10 G
#127100000000
0!
0*
09
0>
0C
#127110000000
1!
1*
b11 6
19
1>
1C
b11 G
#127120000000
0!
0*
09
0>
0C
#127130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#127140000000
0!
0*
09
0>
0C
#127150000000
1!
1*
b101 6
19
1>
1C
b101 G
#127160000000
0!
0*
09
0>
0C
#127170000000
1!
1*
b110 6
19
1>
1C
b110 G
#127180000000
0!
0*
09
0>
0C
#127190000000
1!
1*
b111 6
19
1>
1C
b111 G
#127200000000
0!
1"
0*
1+
09
1:
0>
0C
#127210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#127220000000
0!
0*
09
0>
0C
#127230000000
1!
1*
b1 6
19
1>
1C
b1 G
#127240000000
0!
0*
09
0>
0C
#127250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#127260000000
0!
0*
09
0>
0C
#127270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#127280000000
0!
0*
09
0>
0C
#127290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#127300000000
0!
0*
09
0>
0C
#127310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#127320000000
0!
0#
0*
0,
09
0>
0?
0C
#127330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#127340000000
0!
0*
09
0>
0C
#127350000000
1!
1*
19
1>
1C
#127360000000
0!
0*
09
0>
0C
#127370000000
1!
1*
19
1>
1C
#127380000000
0!
0*
09
0>
0C
#127390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#127400000000
0!
0*
09
0>
0C
#127410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#127420000000
0!
0*
09
0>
0C
#127430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#127440000000
0!
0*
09
0>
0C
#127450000000
1!
1*
b10 6
19
1>
1C
b10 G
#127460000000
0!
0*
09
0>
0C
#127470000000
1!
1*
b11 6
19
1>
1C
b11 G
#127480000000
0!
0*
09
0>
0C
#127490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#127500000000
0!
0*
09
0>
0C
#127510000000
1!
1*
b101 6
19
1>
1C
b101 G
#127520000000
0!
0*
09
0>
0C
#127530000000
1!
1*
b110 6
19
1>
1C
b110 G
#127540000000
0!
0*
09
0>
0C
#127550000000
1!
1*
b111 6
19
1>
1C
b111 G
#127560000000
0!
0*
09
0>
0C
#127570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#127580000000
0!
0*
09
0>
0C
#127590000000
1!
1*
b1 6
19
1>
1C
b1 G
#127600000000
0!
0*
09
0>
0C
#127610000000
1!
1*
b10 6
19
1>
1C
b10 G
#127620000000
0!
0*
09
0>
0C
#127630000000
1!
1*
b11 6
19
1>
1C
b11 G
#127640000000
0!
0*
09
0>
0C
#127650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#127660000000
0!
0*
09
0>
0C
#127670000000
1!
1*
b101 6
19
1>
1C
b101 G
#127680000000
0!
0*
09
0>
0C
#127690000000
1!
1*
b110 6
19
1>
1C
b110 G
#127700000000
0!
0*
09
0>
0C
#127710000000
1!
1*
b111 6
19
1>
1C
b111 G
#127720000000
0!
0*
09
0>
0C
#127730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#127740000000
0!
0*
09
0>
0C
#127750000000
1!
1*
b1 6
19
1>
1C
b1 G
#127760000000
0!
0*
09
0>
0C
#127770000000
1!
1*
b10 6
19
1>
1C
b10 G
#127780000000
0!
0*
09
0>
0C
#127790000000
1!
1*
b11 6
19
1>
1C
b11 G
#127800000000
0!
0*
09
0>
0C
#127810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#127820000000
0!
0*
09
0>
0C
#127830000000
1!
1*
b101 6
19
1>
1C
b101 G
#127840000000
0!
0*
09
0>
0C
#127850000000
1!
1*
b110 6
19
1>
1C
b110 G
#127860000000
0!
0*
09
0>
0C
#127870000000
1!
1*
b111 6
19
1>
1C
b111 G
#127880000000
0!
1"
0*
1+
09
1:
0>
0C
#127890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#127900000000
0!
0*
09
0>
0C
#127910000000
1!
1*
b1 6
19
1>
1C
b1 G
#127920000000
0!
0*
09
0>
0C
#127930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#127940000000
0!
0*
09
0>
0C
#127950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#127960000000
0!
0*
09
0>
0C
#127970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#127980000000
0!
0*
09
0>
0C
#127990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#128000000000
0!
0#
0*
0,
09
0>
0?
0C
#128010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#128020000000
0!
0*
09
0>
0C
#128030000000
1!
1*
19
1>
1C
#128040000000
0!
0*
09
0>
0C
#128050000000
1!
1*
19
1>
1C
#128060000000
0!
0*
09
0>
0C
#128070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#128080000000
0!
0*
09
0>
0C
#128090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#128100000000
0!
0*
09
0>
0C
#128110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#128120000000
0!
0*
09
0>
0C
#128130000000
1!
1*
b10 6
19
1>
1C
b10 G
#128140000000
0!
0*
09
0>
0C
#128150000000
1!
1*
b11 6
19
1>
1C
b11 G
#128160000000
0!
0*
09
0>
0C
#128170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#128180000000
0!
0*
09
0>
0C
#128190000000
1!
1*
b101 6
19
1>
1C
b101 G
#128200000000
0!
0*
09
0>
0C
#128210000000
1!
1*
b110 6
19
1>
1C
b110 G
#128220000000
0!
0*
09
0>
0C
#128230000000
1!
1*
b111 6
19
1>
1C
b111 G
#128240000000
0!
0*
09
0>
0C
#128250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#128260000000
0!
0*
09
0>
0C
#128270000000
1!
1*
b1 6
19
1>
1C
b1 G
#128280000000
0!
0*
09
0>
0C
#128290000000
1!
1*
b10 6
19
1>
1C
b10 G
#128300000000
0!
0*
09
0>
0C
#128310000000
1!
1*
b11 6
19
1>
1C
b11 G
#128320000000
0!
0*
09
0>
0C
#128330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#128340000000
0!
0*
09
0>
0C
#128350000000
1!
1*
b101 6
19
1>
1C
b101 G
#128360000000
0!
0*
09
0>
0C
#128370000000
1!
1*
b110 6
19
1>
1C
b110 G
#128380000000
0!
0*
09
0>
0C
#128390000000
1!
1*
b111 6
19
1>
1C
b111 G
#128400000000
0!
0*
09
0>
0C
#128410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#128420000000
0!
0*
09
0>
0C
#128430000000
1!
1*
b1 6
19
1>
1C
b1 G
#128440000000
0!
0*
09
0>
0C
#128450000000
1!
1*
b10 6
19
1>
1C
b10 G
#128460000000
0!
0*
09
0>
0C
#128470000000
1!
1*
b11 6
19
1>
1C
b11 G
#128480000000
0!
0*
09
0>
0C
#128490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#128500000000
0!
0*
09
0>
0C
#128510000000
1!
1*
b101 6
19
1>
1C
b101 G
#128520000000
0!
0*
09
0>
0C
#128530000000
1!
1*
b110 6
19
1>
1C
b110 G
#128540000000
0!
0*
09
0>
0C
#128550000000
1!
1*
b111 6
19
1>
1C
b111 G
#128560000000
0!
1"
0*
1+
09
1:
0>
0C
#128570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#128580000000
0!
0*
09
0>
0C
#128590000000
1!
1*
b1 6
19
1>
1C
b1 G
#128600000000
0!
0*
09
0>
0C
#128610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#128620000000
0!
0*
09
0>
0C
#128630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#128640000000
0!
0*
09
0>
0C
#128650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#128660000000
0!
0*
09
0>
0C
#128670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#128680000000
0!
0#
0*
0,
09
0>
0?
0C
#128690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#128700000000
0!
0*
09
0>
0C
#128710000000
1!
1*
19
1>
1C
#128720000000
0!
0*
09
0>
0C
#128730000000
1!
1*
19
1>
1C
#128740000000
0!
0*
09
0>
0C
#128750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#128760000000
0!
0*
09
0>
0C
#128770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#128780000000
0!
0*
09
0>
0C
#128790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#128800000000
0!
0*
09
0>
0C
#128810000000
1!
1*
b10 6
19
1>
1C
b10 G
#128820000000
0!
0*
09
0>
0C
#128830000000
1!
1*
b11 6
19
1>
1C
b11 G
#128840000000
0!
0*
09
0>
0C
#128850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#128860000000
0!
0*
09
0>
0C
#128870000000
1!
1*
b101 6
19
1>
1C
b101 G
#128880000000
0!
0*
09
0>
0C
#128890000000
1!
1*
b110 6
19
1>
1C
b110 G
#128900000000
0!
0*
09
0>
0C
#128910000000
1!
1*
b111 6
19
1>
1C
b111 G
#128920000000
0!
0*
09
0>
0C
#128930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#128940000000
0!
0*
09
0>
0C
#128950000000
1!
1*
b1 6
19
1>
1C
b1 G
#128960000000
0!
0*
09
0>
0C
#128970000000
1!
1*
b10 6
19
1>
1C
b10 G
#128980000000
0!
0*
09
0>
0C
#128990000000
1!
1*
b11 6
19
1>
1C
b11 G
#129000000000
0!
0*
09
0>
0C
#129010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#129020000000
0!
0*
09
0>
0C
#129030000000
1!
1*
b101 6
19
1>
1C
b101 G
#129040000000
0!
0*
09
0>
0C
#129050000000
1!
1*
b110 6
19
1>
1C
b110 G
#129060000000
0!
0*
09
0>
0C
#129070000000
1!
1*
b111 6
19
1>
1C
b111 G
#129080000000
0!
0*
09
0>
0C
#129090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#129100000000
0!
0*
09
0>
0C
#129110000000
1!
1*
b1 6
19
1>
1C
b1 G
#129120000000
0!
0*
09
0>
0C
#129130000000
1!
1*
b10 6
19
1>
1C
b10 G
#129140000000
0!
0*
09
0>
0C
#129150000000
1!
1*
b11 6
19
1>
1C
b11 G
#129160000000
0!
0*
09
0>
0C
#129170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#129180000000
0!
0*
09
0>
0C
#129190000000
1!
1*
b101 6
19
1>
1C
b101 G
#129200000000
0!
0*
09
0>
0C
#129210000000
1!
1*
b110 6
19
1>
1C
b110 G
#129220000000
0!
0*
09
0>
0C
#129230000000
1!
1*
b111 6
19
1>
1C
b111 G
#129240000000
0!
1"
0*
1+
09
1:
0>
0C
#129250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#129260000000
0!
0*
09
0>
0C
#129270000000
1!
1*
b1 6
19
1>
1C
b1 G
#129280000000
0!
0*
09
0>
0C
#129290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#129300000000
0!
0*
09
0>
0C
#129310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#129320000000
0!
0*
09
0>
0C
#129330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#129340000000
0!
0*
09
0>
0C
#129350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#129360000000
0!
0#
0*
0,
09
0>
0?
0C
#129370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#129380000000
0!
0*
09
0>
0C
#129390000000
1!
1*
19
1>
1C
#129400000000
0!
0*
09
0>
0C
#129410000000
1!
1*
19
1>
1C
#129420000000
0!
0*
09
0>
0C
#129430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#129440000000
0!
0*
09
0>
0C
#129450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#129460000000
0!
0*
09
0>
0C
#129470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#129480000000
0!
0*
09
0>
0C
#129490000000
1!
1*
b10 6
19
1>
1C
b10 G
#129500000000
0!
0*
09
0>
0C
#129510000000
1!
1*
b11 6
19
1>
1C
b11 G
#129520000000
0!
0*
09
0>
0C
#129530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#129540000000
0!
0*
09
0>
0C
#129550000000
1!
1*
b101 6
19
1>
1C
b101 G
#129560000000
0!
0*
09
0>
0C
#129570000000
1!
1*
b110 6
19
1>
1C
b110 G
#129580000000
0!
0*
09
0>
0C
#129590000000
1!
1*
b111 6
19
1>
1C
b111 G
#129600000000
0!
0*
09
0>
0C
#129610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#129620000000
0!
0*
09
0>
0C
#129630000000
1!
1*
b1 6
19
1>
1C
b1 G
#129640000000
0!
0*
09
0>
0C
#129650000000
1!
1*
b10 6
19
1>
1C
b10 G
#129660000000
0!
0*
09
0>
0C
#129670000000
1!
1*
b11 6
19
1>
1C
b11 G
#129680000000
0!
0*
09
0>
0C
#129690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#129700000000
0!
0*
09
0>
0C
#129710000000
1!
1*
b101 6
19
1>
1C
b101 G
#129720000000
0!
0*
09
0>
0C
#129730000000
1!
1*
b110 6
19
1>
1C
b110 G
#129740000000
0!
0*
09
0>
0C
#129750000000
1!
1*
b111 6
19
1>
1C
b111 G
#129760000000
0!
0*
09
0>
0C
#129770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#129780000000
0!
0*
09
0>
0C
#129790000000
1!
1*
b1 6
19
1>
1C
b1 G
#129800000000
0!
0*
09
0>
0C
#129810000000
1!
1*
b10 6
19
1>
1C
b10 G
#129820000000
0!
0*
09
0>
0C
#129830000000
1!
1*
b11 6
19
1>
1C
b11 G
#129840000000
0!
0*
09
0>
0C
#129850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#129860000000
0!
0*
09
0>
0C
#129870000000
1!
1*
b101 6
19
1>
1C
b101 G
#129880000000
0!
0*
09
0>
0C
#129890000000
1!
1*
b110 6
19
1>
1C
b110 G
#129900000000
0!
0*
09
0>
0C
#129910000000
1!
1*
b111 6
19
1>
1C
b111 G
#129920000000
0!
1"
0*
1+
09
1:
0>
0C
#129930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#129940000000
0!
0*
09
0>
0C
#129950000000
1!
1*
b1 6
19
1>
1C
b1 G
#129960000000
0!
0*
09
0>
0C
#129970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#129980000000
0!
0*
09
0>
0C
#129990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#130000000000
0!
0*
09
0>
0C
#130010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#130020000000
0!
0*
09
0>
0C
#130030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#130040000000
0!
0#
0*
0,
09
0>
0?
0C
#130050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#130060000000
0!
0*
09
0>
0C
#130070000000
1!
1*
19
1>
1C
#130080000000
0!
0*
09
0>
0C
#130090000000
1!
1*
19
1>
1C
#130100000000
0!
0*
09
0>
0C
#130110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#130120000000
0!
0*
09
0>
0C
#130130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#130140000000
0!
0*
09
0>
0C
#130150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#130160000000
0!
0*
09
0>
0C
#130170000000
1!
1*
b10 6
19
1>
1C
b10 G
#130180000000
0!
0*
09
0>
0C
#130190000000
1!
1*
b11 6
19
1>
1C
b11 G
#130200000000
0!
0*
09
0>
0C
#130210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#130220000000
0!
0*
09
0>
0C
#130230000000
1!
1*
b101 6
19
1>
1C
b101 G
#130240000000
0!
0*
09
0>
0C
#130250000000
1!
1*
b110 6
19
1>
1C
b110 G
#130260000000
0!
0*
09
0>
0C
#130270000000
1!
1*
b111 6
19
1>
1C
b111 G
#130280000000
0!
0*
09
0>
0C
#130290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#130300000000
0!
0*
09
0>
0C
#130310000000
1!
1*
b1 6
19
1>
1C
b1 G
#130320000000
0!
0*
09
0>
0C
#130330000000
1!
1*
b10 6
19
1>
1C
b10 G
#130340000000
0!
0*
09
0>
0C
#130350000000
1!
1*
b11 6
19
1>
1C
b11 G
#130360000000
0!
0*
09
0>
0C
#130370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#130380000000
0!
0*
09
0>
0C
#130390000000
1!
1*
b101 6
19
1>
1C
b101 G
#130400000000
0!
0*
09
0>
0C
#130410000000
1!
1*
b110 6
19
1>
1C
b110 G
#130420000000
0!
0*
09
0>
0C
#130430000000
1!
1*
b111 6
19
1>
1C
b111 G
#130440000000
0!
0*
09
0>
0C
#130450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#130460000000
0!
0*
09
0>
0C
#130470000000
1!
1*
b1 6
19
1>
1C
b1 G
#130480000000
0!
0*
09
0>
0C
#130490000000
1!
1*
b10 6
19
1>
1C
b10 G
#130500000000
0!
0*
09
0>
0C
#130510000000
1!
1*
b11 6
19
1>
1C
b11 G
#130520000000
0!
0*
09
0>
0C
#130530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#130540000000
0!
0*
09
0>
0C
#130550000000
1!
1*
b101 6
19
1>
1C
b101 G
#130560000000
0!
0*
09
0>
0C
#130570000000
1!
1*
b110 6
19
1>
1C
b110 G
#130580000000
0!
0*
09
0>
0C
#130590000000
1!
1*
b111 6
19
1>
1C
b111 G
#130600000000
0!
1"
0*
1+
09
1:
0>
0C
#130610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#130620000000
0!
0*
09
0>
0C
#130630000000
1!
1*
b1 6
19
1>
1C
b1 G
#130640000000
0!
0*
09
0>
0C
#130650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#130660000000
0!
0*
09
0>
0C
#130670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#130680000000
0!
0*
09
0>
0C
#130690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#130700000000
0!
0*
09
0>
0C
#130710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#130720000000
0!
0#
0*
0,
09
0>
0?
0C
#130730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#130740000000
0!
0*
09
0>
0C
#130750000000
1!
1*
19
1>
1C
#130760000000
0!
0*
09
0>
0C
#130770000000
1!
1*
19
1>
1C
#130780000000
0!
0*
09
0>
0C
#130790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#130800000000
0!
0*
09
0>
0C
#130810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#130820000000
0!
0*
09
0>
0C
#130830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#130840000000
0!
0*
09
0>
0C
#130850000000
1!
1*
b10 6
19
1>
1C
b10 G
#130860000000
0!
0*
09
0>
0C
#130870000000
1!
1*
b11 6
19
1>
1C
b11 G
#130880000000
0!
0*
09
0>
0C
#130890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#130900000000
0!
0*
09
0>
0C
#130910000000
1!
1*
b101 6
19
1>
1C
b101 G
#130920000000
0!
0*
09
0>
0C
#130930000000
1!
1*
b110 6
19
1>
1C
b110 G
#130940000000
0!
0*
09
0>
0C
#130950000000
1!
1*
b111 6
19
1>
1C
b111 G
#130960000000
0!
0*
09
0>
0C
#130970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#130980000000
0!
0*
09
0>
0C
#130990000000
1!
1*
b1 6
19
1>
1C
b1 G
#131000000000
0!
0*
09
0>
0C
#131010000000
1!
1*
b10 6
19
1>
1C
b10 G
#131020000000
0!
0*
09
0>
0C
#131030000000
1!
1*
b11 6
19
1>
1C
b11 G
#131040000000
0!
0*
09
0>
0C
#131050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#131060000000
0!
0*
09
0>
0C
#131070000000
1!
1*
b101 6
19
1>
1C
b101 G
#131080000000
0!
0*
09
0>
0C
#131090000000
1!
1*
b110 6
19
1>
1C
b110 G
#131100000000
0!
0*
09
0>
0C
#131110000000
1!
1*
b111 6
19
1>
1C
b111 G
#131120000000
0!
0*
09
0>
0C
#131130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#131140000000
0!
0*
09
0>
0C
#131150000000
1!
1*
b1 6
19
1>
1C
b1 G
#131160000000
0!
0*
09
0>
0C
#131170000000
1!
1*
b10 6
19
1>
1C
b10 G
#131180000000
0!
0*
09
0>
0C
#131190000000
1!
1*
b11 6
19
1>
1C
b11 G
#131200000000
0!
0*
09
0>
0C
#131210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#131220000000
0!
0*
09
0>
0C
#131230000000
1!
1*
b101 6
19
1>
1C
b101 G
#131240000000
0!
0*
09
0>
0C
#131250000000
1!
1*
b110 6
19
1>
1C
b110 G
#131260000000
0!
0*
09
0>
0C
#131270000000
1!
1*
b111 6
19
1>
1C
b111 G
#131280000000
0!
1"
0*
1+
09
1:
0>
0C
#131290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#131300000000
0!
0*
09
0>
0C
#131310000000
1!
1*
b1 6
19
1>
1C
b1 G
#131320000000
0!
0*
09
0>
0C
#131330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#131340000000
0!
0*
09
0>
0C
#131350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#131360000000
0!
0*
09
0>
0C
#131370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#131380000000
0!
0*
09
0>
0C
#131390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#131400000000
0!
0#
0*
0,
09
0>
0?
0C
#131410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#131420000000
0!
0*
09
0>
0C
#131430000000
1!
1*
19
1>
1C
#131440000000
0!
0*
09
0>
0C
#131450000000
1!
1*
19
1>
1C
#131460000000
0!
0*
09
0>
0C
#131470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#131480000000
0!
0*
09
0>
0C
#131490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#131500000000
0!
0*
09
0>
0C
#131510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#131520000000
0!
0*
09
0>
0C
#131530000000
1!
1*
b10 6
19
1>
1C
b10 G
#131540000000
0!
0*
09
0>
0C
#131550000000
1!
1*
b11 6
19
1>
1C
b11 G
#131560000000
0!
0*
09
0>
0C
#131570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#131580000000
0!
0*
09
0>
0C
#131590000000
1!
1*
b101 6
19
1>
1C
b101 G
#131600000000
0!
0*
09
0>
0C
#131610000000
1!
1*
b110 6
19
1>
1C
b110 G
#131620000000
0!
0*
09
0>
0C
#131630000000
1!
1*
b111 6
19
1>
1C
b111 G
#131640000000
0!
0*
09
0>
0C
#131650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#131660000000
0!
0*
09
0>
0C
#131670000000
1!
1*
b1 6
19
1>
1C
b1 G
#131680000000
0!
0*
09
0>
0C
#131690000000
1!
1*
b10 6
19
1>
1C
b10 G
#131700000000
0!
0*
09
0>
0C
#131710000000
1!
1*
b11 6
19
1>
1C
b11 G
#131720000000
0!
0*
09
0>
0C
#131730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#131740000000
0!
0*
09
0>
0C
#131750000000
1!
1*
b101 6
19
1>
1C
b101 G
#131760000000
0!
0*
09
0>
0C
#131770000000
1!
1*
b110 6
19
1>
1C
b110 G
#131780000000
0!
0*
09
0>
0C
#131790000000
1!
1*
b111 6
19
1>
1C
b111 G
#131800000000
0!
0*
09
0>
0C
#131810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#131820000000
0!
0*
09
0>
0C
#131830000000
1!
1*
b1 6
19
1>
1C
b1 G
#131840000000
0!
0*
09
0>
0C
#131850000000
1!
1*
b10 6
19
1>
1C
b10 G
#131860000000
0!
0*
09
0>
0C
#131870000000
1!
1*
b11 6
19
1>
1C
b11 G
#131880000000
0!
0*
09
0>
0C
#131890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#131900000000
0!
0*
09
0>
0C
#131910000000
1!
1*
b101 6
19
1>
1C
b101 G
#131920000000
0!
0*
09
0>
0C
#131930000000
1!
1*
b110 6
19
1>
1C
b110 G
#131940000000
0!
0*
09
0>
0C
#131950000000
1!
1*
b111 6
19
1>
1C
b111 G
#131960000000
0!
1"
0*
1+
09
1:
0>
0C
#131970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#131980000000
0!
0*
09
0>
0C
#131990000000
1!
1*
b1 6
19
1>
1C
b1 G
#132000000000
0!
0*
09
0>
0C
#132010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#132020000000
0!
0*
09
0>
0C
#132030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#132040000000
0!
0*
09
0>
0C
#132050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#132060000000
0!
0*
09
0>
0C
#132070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#132080000000
0!
0#
0*
0,
09
0>
0?
0C
#132090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#132100000000
0!
0*
09
0>
0C
#132110000000
1!
1*
19
1>
1C
#132120000000
0!
0*
09
0>
0C
#132130000000
1!
1*
19
1>
1C
#132140000000
0!
0*
09
0>
0C
#132150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#132160000000
0!
0*
09
0>
0C
#132170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#132180000000
0!
0*
09
0>
0C
#132190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#132200000000
0!
0*
09
0>
0C
#132210000000
1!
1*
b10 6
19
1>
1C
b10 G
#132220000000
0!
0*
09
0>
0C
#132230000000
1!
1*
b11 6
19
1>
1C
b11 G
#132240000000
0!
0*
09
0>
0C
#132250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#132260000000
0!
0*
09
0>
0C
#132270000000
1!
1*
b101 6
19
1>
1C
b101 G
#132280000000
0!
0*
09
0>
0C
#132290000000
1!
1*
b110 6
19
1>
1C
b110 G
#132300000000
0!
0*
09
0>
0C
#132310000000
1!
1*
b111 6
19
1>
1C
b111 G
#132320000000
0!
0*
09
0>
0C
#132330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#132340000000
0!
0*
09
0>
0C
#132350000000
1!
1*
b1 6
19
1>
1C
b1 G
#132360000000
0!
0*
09
0>
0C
#132370000000
1!
1*
b10 6
19
1>
1C
b10 G
#132380000000
0!
0*
09
0>
0C
#132390000000
1!
1*
b11 6
19
1>
1C
b11 G
#132400000000
0!
0*
09
0>
0C
#132410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#132420000000
0!
0*
09
0>
0C
#132430000000
1!
1*
b101 6
19
1>
1C
b101 G
#132440000000
0!
0*
09
0>
0C
#132450000000
1!
1*
b110 6
19
1>
1C
b110 G
#132460000000
0!
0*
09
0>
0C
#132470000000
1!
1*
b111 6
19
1>
1C
b111 G
#132480000000
0!
0*
09
0>
0C
#132490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#132500000000
0!
0*
09
0>
0C
#132510000000
1!
1*
b1 6
19
1>
1C
b1 G
#132520000000
0!
0*
09
0>
0C
#132530000000
1!
1*
b10 6
19
1>
1C
b10 G
#132540000000
0!
0*
09
0>
0C
#132550000000
1!
1*
b11 6
19
1>
1C
b11 G
#132560000000
0!
0*
09
0>
0C
#132570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#132580000000
0!
0*
09
0>
0C
#132590000000
1!
1*
b101 6
19
1>
1C
b101 G
#132600000000
0!
0*
09
0>
0C
#132610000000
1!
1*
b110 6
19
1>
1C
b110 G
#132620000000
0!
0*
09
0>
0C
#132630000000
1!
1*
b111 6
19
1>
1C
b111 G
#132640000000
0!
1"
0*
1+
09
1:
0>
0C
#132650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#132660000000
0!
0*
09
0>
0C
#132670000000
1!
1*
b1 6
19
1>
1C
b1 G
#132680000000
0!
0*
09
0>
0C
#132690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#132700000000
0!
0*
09
0>
0C
#132710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#132720000000
0!
0*
09
0>
0C
#132730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#132740000000
0!
0*
09
0>
0C
#132750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#132760000000
0!
0#
0*
0,
09
0>
0?
0C
#132770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#132780000000
0!
0*
09
0>
0C
#132790000000
1!
1*
19
1>
1C
#132800000000
0!
0*
09
0>
0C
#132810000000
1!
1*
19
1>
1C
#132820000000
0!
0*
09
0>
0C
#132830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#132840000000
0!
0*
09
0>
0C
#132850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#132860000000
0!
0*
09
0>
0C
#132870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#132880000000
0!
0*
09
0>
0C
#132890000000
1!
1*
b10 6
19
1>
1C
b10 G
#132900000000
0!
0*
09
0>
0C
#132910000000
1!
1*
b11 6
19
1>
1C
b11 G
#132920000000
0!
0*
09
0>
0C
#132930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#132940000000
0!
0*
09
0>
0C
#132950000000
1!
1*
b101 6
19
1>
1C
b101 G
#132960000000
0!
0*
09
0>
0C
#132970000000
1!
1*
b110 6
19
1>
1C
b110 G
#132980000000
0!
0*
09
0>
0C
#132990000000
1!
1*
b111 6
19
1>
1C
b111 G
#133000000000
0!
0*
09
0>
0C
#133010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#133020000000
0!
0*
09
0>
0C
#133030000000
1!
1*
b1 6
19
1>
1C
b1 G
#133040000000
0!
0*
09
0>
0C
#133050000000
1!
1*
b10 6
19
1>
1C
b10 G
#133060000000
0!
0*
09
0>
0C
#133070000000
1!
1*
b11 6
19
1>
1C
b11 G
#133080000000
0!
0*
09
0>
0C
#133090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#133100000000
0!
0*
09
0>
0C
#133110000000
1!
1*
b101 6
19
1>
1C
b101 G
#133120000000
0!
0*
09
0>
0C
#133130000000
1!
1*
b110 6
19
1>
1C
b110 G
#133140000000
0!
0*
09
0>
0C
#133150000000
1!
1*
b111 6
19
1>
1C
b111 G
#133160000000
0!
0*
09
0>
0C
#133170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#133180000000
0!
0*
09
0>
0C
#133190000000
1!
1*
b1 6
19
1>
1C
b1 G
#133200000000
0!
0*
09
0>
0C
#133210000000
1!
1*
b10 6
19
1>
1C
b10 G
#133220000000
0!
0*
09
0>
0C
#133230000000
1!
1*
b11 6
19
1>
1C
b11 G
#133240000000
0!
0*
09
0>
0C
#133250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#133260000000
0!
0*
09
0>
0C
#133270000000
1!
1*
b101 6
19
1>
1C
b101 G
#133280000000
0!
0*
09
0>
0C
#133290000000
1!
1*
b110 6
19
1>
1C
b110 G
#133300000000
0!
0*
09
0>
0C
#133310000000
1!
1*
b111 6
19
1>
1C
b111 G
#133320000000
0!
1"
0*
1+
09
1:
0>
0C
#133330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#133340000000
0!
0*
09
0>
0C
#133350000000
1!
1*
b1 6
19
1>
1C
b1 G
#133360000000
0!
0*
09
0>
0C
#133370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#133380000000
0!
0*
09
0>
0C
#133390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#133400000000
0!
0*
09
0>
0C
#133410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#133420000000
0!
0*
09
0>
0C
#133430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#133440000000
0!
0#
0*
0,
09
0>
0?
0C
#133450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#133460000000
0!
0*
09
0>
0C
#133470000000
1!
1*
19
1>
1C
#133480000000
0!
0*
09
0>
0C
#133490000000
1!
1*
19
1>
1C
#133500000000
0!
0*
09
0>
0C
#133510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#133520000000
0!
0*
09
0>
0C
#133530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#133540000000
0!
0*
09
0>
0C
#133550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#133560000000
0!
0*
09
0>
0C
#133570000000
1!
1*
b10 6
19
1>
1C
b10 G
#133580000000
0!
0*
09
0>
0C
#133590000000
1!
1*
b11 6
19
1>
1C
b11 G
#133600000000
0!
0*
09
0>
0C
#133610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#133620000000
0!
0*
09
0>
0C
#133630000000
1!
1*
b101 6
19
1>
1C
b101 G
#133640000000
0!
0*
09
0>
0C
#133650000000
1!
1*
b110 6
19
1>
1C
b110 G
#133660000000
0!
0*
09
0>
0C
#133670000000
1!
1*
b111 6
19
1>
1C
b111 G
#133680000000
0!
0*
09
0>
0C
#133690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#133700000000
0!
0*
09
0>
0C
#133710000000
1!
1*
b1 6
19
1>
1C
b1 G
#133720000000
0!
0*
09
0>
0C
#133730000000
1!
1*
b10 6
19
1>
1C
b10 G
#133740000000
0!
0*
09
0>
0C
#133750000000
1!
1*
b11 6
19
1>
1C
b11 G
#133760000000
0!
0*
09
0>
0C
#133770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#133780000000
0!
0*
09
0>
0C
#133790000000
1!
1*
b101 6
19
1>
1C
b101 G
#133800000000
0!
0*
09
0>
0C
#133810000000
1!
1*
b110 6
19
1>
1C
b110 G
#133820000000
0!
0*
09
0>
0C
#133830000000
1!
1*
b111 6
19
1>
1C
b111 G
#133840000000
0!
0*
09
0>
0C
#133850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#133860000000
0!
0*
09
0>
0C
#133870000000
1!
1*
b1 6
19
1>
1C
b1 G
#133880000000
0!
0*
09
0>
0C
#133890000000
1!
1*
b10 6
19
1>
1C
b10 G
#133900000000
0!
0*
09
0>
0C
#133910000000
1!
1*
b11 6
19
1>
1C
b11 G
#133920000000
0!
0*
09
0>
0C
#133930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#133940000000
0!
0*
09
0>
0C
#133950000000
1!
1*
b101 6
19
1>
1C
b101 G
#133960000000
0!
0*
09
0>
0C
#133970000000
1!
1*
b110 6
19
1>
1C
b110 G
#133980000000
0!
0*
09
0>
0C
#133990000000
1!
1*
b111 6
19
1>
1C
b111 G
#134000000000
0!
1"
0*
1+
09
1:
0>
0C
#134010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#134020000000
0!
0*
09
0>
0C
#134030000000
1!
1*
b1 6
19
1>
1C
b1 G
#134040000000
0!
0*
09
0>
0C
#134050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#134060000000
0!
0*
09
0>
0C
#134070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#134080000000
0!
0*
09
0>
0C
#134090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#134100000000
0!
0*
09
0>
0C
#134110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#134120000000
0!
0#
0*
0,
09
0>
0?
0C
#134130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#134140000000
0!
0*
09
0>
0C
#134150000000
1!
1*
19
1>
1C
#134160000000
0!
0*
09
0>
0C
#134170000000
1!
1*
19
1>
1C
#134180000000
0!
0*
09
0>
0C
#134190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#134200000000
0!
0*
09
0>
0C
#134210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#134220000000
0!
0*
09
0>
0C
#134230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#134240000000
0!
0*
09
0>
0C
#134250000000
1!
1*
b10 6
19
1>
1C
b10 G
#134260000000
0!
0*
09
0>
0C
#134270000000
1!
1*
b11 6
19
1>
1C
b11 G
#134280000000
0!
0*
09
0>
0C
#134290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#134300000000
0!
0*
09
0>
0C
#134310000000
1!
1*
b101 6
19
1>
1C
b101 G
#134320000000
0!
0*
09
0>
0C
#134330000000
1!
1*
b110 6
19
1>
1C
b110 G
#134340000000
0!
0*
09
0>
0C
#134350000000
1!
1*
b111 6
19
1>
1C
b111 G
#134360000000
0!
0*
09
0>
0C
#134370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#134380000000
0!
0*
09
0>
0C
#134390000000
1!
1*
b1 6
19
1>
1C
b1 G
#134400000000
0!
0*
09
0>
0C
#134410000000
1!
1*
b10 6
19
1>
1C
b10 G
#134420000000
0!
0*
09
0>
0C
#134430000000
1!
1*
b11 6
19
1>
1C
b11 G
#134440000000
0!
0*
09
0>
0C
#134450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#134460000000
0!
0*
09
0>
0C
#134470000000
1!
1*
b101 6
19
1>
1C
b101 G
#134480000000
0!
0*
09
0>
0C
#134490000000
1!
1*
b110 6
19
1>
1C
b110 G
#134500000000
0!
0*
09
0>
0C
#134510000000
1!
1*
b111 6
19
1>
1C
b111 G
#134520000000
0!
0*
09
0>
0C
#134530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#134540000000
0!
0*
09
0>
0C
#134550000000
1!
1*
b1 6
19
1>
1C
b1 G
#134560000000
0!
0*
09
0>
0C
#134570000000
1!
1*
b10 6
19
1>
1C
b10 G
#134580000000
0!
0*
09
0>
0C
#134590000000
1!
1*
b11 6
19
1>
1C
b11 G
#134600000000
0!
0*
09
0>
0C
#134610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#134620000000
0!
0*
09
0>
0C
#134630000000
1!
1*
b101 6
19
1>
1C
b101 G
#134640000000
0!
0*
09
0>
0C
#134650000000
1!
1*
b110 6
19
1>
1C
b110 G
#134660000000
0!
0*
09
0>
0C
#134670000000
1!
1*
b111 6
19
1>
1C
b111 G
#134680000000
0!
1"
0*
1+
09
1:
0>
0C
#134690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#134700000000
0!
0*
09
0>
0C
#134710000000
1!
1*
b1 6
19
1>
1C
b1 G
#134720000000
0!
0*
09
0>
0C
#134730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#134740000000
0!
0*
09
0>
0C
#134750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#134760000000
0!
0*
09
0>
0C
#134770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#134780000000
0!
0*
09
0>
0C
#134790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#134800000000
0!
0#
0*
0,
09
0>
0?
0C
#134810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#134820000000
0!
0*
09
0>
0C
#134830000000
1!
1*
19
1>
1C
#134840000000
0!
0*
09
0>
0C
#134850000000
1!
1*
19
1>
1C
#134860000000
0!
0*
09
0>
0C
#134870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#134880000000
0!
0*
09
0>
0C
#134890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#134900000000
0!
0*
09
0>
0C
#134910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#134920000000
0!
0*
09
0>
0C
#134930000000
1!
1*
b10 6
19
1>
1C
b10 G
#134940000000
0!
0*
09
0>
0C
#134950000000
1!
1*
b11 6
19
1>
1C
b11 G
#134960000000
0!
0*
09
0>
0C
#134970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#134980000000
0!
0*
09
0>
0C
#134990000000
1!
1*
b101 6
19
1>
1C
b101 G
#135000000000
0!
0*
09
0>
0C
#135010000000
1!
1*
b110 6
19
1>
1C
b110 G
#135020000000
0!
0*
09
0>
0C
#135030000000
1!
1*
b111 6
19
1>
1C
b111 G
#135040000000
0!
0*
09
0>
0C
#135050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#135060000000
0!
0*
09
0>
0C
#135070000000
1!
1*
b1 6
19
1>
1C
b1 G
#135080000000
0!
0*
09
0>
0C
#135090000000
1!
1*
b10 6
19
1>
1C
b10 G
#135100000000
0!
0*
09
0>
0C
#135110000000
1!
1*
b11 6
19
1>
1C
b11 G
#135120000000
0!
0*
09
0>
0C
#135130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#135140000000
0!
0*
09
0>
0C
#135150000000
1!
1*
b101 6
19
1>
1C
b101 G
#135160000000
0!
0*
09
0>
0C
#135170000000
1!
1*
b110 6
19
1>
1C
b110 G
#135180000000
0!
0*
09
0>
0C
#135190000000
1!
1*
b111 6
19
1>
1C
b111 G
#135200000000
0!
0*
09
0>
0C
#135210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#135220000000
0!
0*
09
0>
0C
#135230000000
1!
1*
b1 6
19
1>
1C
b1 G
#135240000000
0!
0*
09
0>
0C
#135250000000
1!
1*
b10 6
19
1>
1C
b10 G
#135260000000
0!
0*
09
0>
0C
#135270000000
1!
1*
b11 6
19
1>
1C
b11 G
#135280000000
0!
0*
09
0>
0C
#135290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#135300000000
0!
0*
09
0>
0C
#135310000000
1!
1*
b101 6
19
1>
1C
b101 G
#135320000000
0!
0*
09
0>
0C
#135330000000
1!
1*
b110 6
19
1>
1C
b110 G
#135340000000
0!
0*
09
0>
0C
#135350000000
1!
1*
b111 6
19
1>
1C
b111 G
#135360000000
0!
1"
0*
1+
09
1:
0>
0C
#135370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#135380000000
0!
0*
09
0>
0C
#135390000000
1!
1*
b1 6
19
1>
1C
b1 G
#135400000000
0!
0*
09
0>
0C
#135410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#135420000000
0!
0*
09
0>
0C
#135430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#135440000000
0!
0*
09
0>
0C
#135450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#135460000000
0!
0*
09
0>
0C
#135470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#135480000000
0!
0#
0*
0,
09
0>
0?
0C
#135490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#135500000000
0!
0*
09
0>
0C
#135510000000
1!
1*
19
1>
1C
#135520000000
0!
0*
09
0>
0C
#135530000000
1!
1*
19
1>
1C
#135540000000
0!
0*
09
0>
0C
#135550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#135560000000
0!
0*
09
0>
0C
#135570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#135580000000
0!
0*
09
0>
0C
#135590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#135600000000
0!
0*
09
0>
0C
#135610000000
1!
1*
b10 6
19
1>
1C
b10 G
#135620000000
0!
0*
09
0>
0C
#135630000000
1!
1*
b11 6
19
1>
1C
b11 G
#135640000000
0!
0*
09
0>
0C
#135650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#135660000000
0!
0*
09
0>
0C
#135670000000
1!
1*
b101 6
19
1>
1C
b101 G
#135680000000
0!
0*
09
0>
0C
#135690000000
1!
1*
b110 6
19
1>
1C
b110 G
#135700000000
0!
0*
09
0>
0C
#135710000000
1!
1*
b111 6
19
1>
1C
b111 G
#135720000000
0!
0*
09
0>
0C
#135730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#135740000000
0!
0*
09
0>
0C
#135750000000
1!
1*
b1 6
19
1>
1C
b1 G
#135760000000
0!
0*
09
0>
0C
#135770000000
1!
1*
b10 6
19
1>
1C
b10 G
#135780000000
0!
0*
09
0>
0C
#135790000000
1!
1*
b11 6
19
1>
1C
b11 G
#135800000000
0!
0*
09
0>
0C
#135810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#135820000000
0!
0*
09
0>
0C
#135830000000
1!
1*
b101 6
19
1>
1C
b101 G
#135840000000
0!
0*
09
0>
0C
#135850000000
1!
1*
b110 6
19
1>
1C
b110 G
#135860000000
0!
0*
09
0>
0C
#135870000000
1!
1*
b111 6
19
1>
1C
b111 G
#135880000000
0!
0*
09
0>
0C
#135890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#135900000000
0!
0*
09
0>
0C
#135910000000
1!
1*
b1 6
19
1>
1C
b1 G
#135920000000
0!
0*
09
0>
0C
#135930000000
1!
1*
b10 6
19
1>
1C
b10 G
#135940000000
0!
0*
09
0>
0C
#135950000000
1!
1*
b11 6
19
1>
1C
b11 G
#135960000000
0!
0*
09
0>
0C
#135970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#135980000000
0!
0*
09
0>
0C
#135990000000
1!
1*
b101 6
19
1>
1C
b101 G
#136000000000
0!
0*
09
0>
0C
#136010000000
1!
1*
b110 6
19
1>
1C
b110 G
#136020000000
0!
0*
09
0>
0C
#136030000000
1!
1*
b111 6
19
1>
1C
b111 G
#136040000000
0!
1"
0*
1+
09
1:
0>
0C
#136050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#136060000000
0!
0*
09
0>
0C
#136070000000
1!
1*
b1 6
19
1>
1C
b1 G
#136080000000
0!
0*
09
0>
0C
#136090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#136100000000
0!
0*
09
0>
0C
#136110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#136120000000
0!
0*
09
0>
0C
#136130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#136140000000
0!
0*
09
0>
0C
#136150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#136160000000
0!
0#
0*
0,
09
0>
0?
0C
#136170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#136180000000
0!
0*
09
0>
0C
#136190000000
1!
1*
19
1>
1C
#136200000000
0!
0*
09
0>
0C
#136210000000
1!
1*
19
1>
1C
#136220000000
0!
0*
09
0>
0C
#136230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#136240000000
0!
0*
09
0>
0C
#136250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#136260000000
0!
0*
09
0>
0C
#136270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#136280000000
0!
0*
09
0>
0C
#136290000000
1!
1*
b10 6
19
1>
1C
b10 G
#136300000000
0!
0*
09
0>
0C
#136310000000
1!
1*
b11 6
19
1>
1C
b11 G
#136320000000
0!
0*
09
0>
0C
#136330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#136340000000
0!
0*
09
0>
0C
#136350000000
1!
1*
b101 6
19
1>
1C
b101 G
#136360000000
0!
0*
09
0>
0C
#136370000000
1!
1*
b110 6
19
1>
1C
b110 G
#136380000000
0!
0*
09
0>
0C
#136390000000
1!
1*
b111 6
19
1>
1C
b111 G
#136400000000
0!
0*
09
0>
0C
#136410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#136420000000
0!
0*
09
0>
0C
#136430000000
1!
1*
b1 6
19
1>
1C
b1 G
#136440000000
0!
0*
09
0>
0C
#136450000000
1!
1*
b10 6
19
1>
1C
b10 G
#136460000000
0!
0*
09
0>
0C
#136470000000
1!
1*
b11 6
19
1>
1C
b11 G
#136480000000
0!
0*
09
0>
0C
#136490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#136500000000
0!
0*
09
0>
0C
#136510000000
1!
1*
b101 6
19
1>
1C
b101 G
#136520000000
0!
0*
09
0>
0C
#136530000000
1!
1*
b110 6
19
1>
1C
b110 G
#136540000000
0!
0*
09
0>
0C
#136550000000
1!
1*
b111 6
19
1>
1C
b111 G
#136560000000
0!
0*
09
0>
0C
#136570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#136580000000
0!
0*
09
0>
0C
#136590000000
1!
1*
b1 6
19
1>
1C
b1 G
#136600000000
0!
0*
09
0>
0C
#136610000000
1!
1*
b10 6
19
1>
1C
b10 G
#136620000000
0!
0*
09
0>
0C
#136630000000
1!
1*
b11 6
19
1>
1C
b11 G
#136640000000
0!
0*
09
0>
0C
#136650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#136660000000
0!
0*
09
0>
0C
#136670000000
1!
1*
b101 6
19
1>
1C
b101 G
#136680000000
0!
0*
09
0>
0C
#136690000000
1!
1*
b110 6
19
1>
1C
b110 G
#136700000000
0!
0*
09
0>
0C
#136710000000
1!
1*
b111 6
19
1>
1C
b111 G
#136720000000
0!
1"
0*
1+
09
1:
0>
0C
#136730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#136740000000
0!
0*
09
0>
0C
#136750000000
1!
1*
b1 6
19
1>
1C
b1 G
#136760000000
0!
0*
09
0>
0C
#136770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#136780000000
0!
0*
09
0>
0C
#136790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#136800000000
0!
0*
09
0>
0C
#136810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#136820000000
0!
0*
09
0>
0C
#136830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#136840000000
0!
0#
0*
0,
09
0>
0?
0C
#136850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#136860000000
0!
0*
09
0>
0C
#136870000000
1!
1*
19
1>
1C
#136880000000
0!
0*
09
0>
0C
#136890000000
1!
1*
19
1>
1C
#136900000000
0!
0*
09
0>
0C
#136910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#136920000000
0!
0*
09
0>
0C
#136930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#136940000000
0!
0*
09
0>
0C
#136950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#136960000000
0!
0*
09
0>
0C
#136970000000
1!
1*
b10 6
19
1>
1C
b10 G
#136980000000
0!
0*
09
0>
0C
#136990000000
1!
1*
b11 6
19
1>
1C
b11 G
#137000000000
0!
0*
09
0>
0C
#137010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#137020000000
0!
0*
09
0>
0C
#137030000000
1!
1*
b101 6
19
1>
1C
b101 G
#137040000000
0!
0*
09
0>
0C
#137050000000
1!
1*
b110 6
19
1>
1C
b110 G
#137060000000
0!
0*
09
0>
0C
#137070000000
1!
1*
b111 6
19
1>
1C
b111 G
#137080000000
0!
0*
09
0>
0C
#137090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#137100000000
0!
0*
09
0>
0C
#137110000000
1!
1*
b1 6
19
1>
1C
b1 G
#137120000000
0!
0*
09
0>
0C
#137130000000
1!
1*
b10 6
19
1>
1C
b10 G
#137140000000
0!
0*
09
0>
0C
#137150000000
1!
1*
b11 6
19
1>
1C
b11 G
#137160000000
0!
0*
09
0>
0C
#137170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#137180000000
0!
0*
09
0>
0C
#137190000000
1!
1*
b101 6
19
1>
1C
b101 G
#137200000000
0!
0*
09
0>
0C
#137210000000
1!
1*
b110 6
19
1>
1C
b110 G
#137220000000
0!
0*
09
0>
0C
#137230000000
1!
1*
b111 6
19
1>
1C
b111 G
#137240000000
0!
0*
09
0>
0C
#137250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#137260000000
0!
0*
09
0>
0C
#137270000000
1!
1*
b1 6
19
1>
1C
b1 G
#137280000000
0!
0*
09
0>
0C
#137290000000
1!
1*
b10 6
19
1>
1C
b10 G
#137300000000
0!
0*
09
0>
0C
#137310000000
1!
1*
b11 6
19
1>
1C
b11 G
#137320000000
0!
0*
09
0>
0C
#137330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#137340000000
0!
0*
09
0>
0C
#137350000000
1!
1*
b101 6
19
1>
1C
b101 G
#137360000000
0!
0*
09
0>
0C
#137370000000
1!
1*
b110 6
19
1>
1C
b110 G
#137380000000
0!
0*
09
0>
0C
#137390000000
1!
1*
b111 6
19
1>
1C
b111 G
#137400000000
0!
1"
0*
1+
09
1:
0>
0C
#137410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#137420000000
0!
0*
09
0>
0C
#137430000000
1!
1*
b1 6
19
1>
1C
b1 G
#137440000000
0!
0*
09
0>
0C
#137450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#137460000000
0!
0*
09
0>
0C
#137470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#137480000000
0!
0*
09
0>
0C
#137490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#137500000000
0!
0*
09
0>
0C
#137510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#137520000000
0!
0#
0*
0,
09
0>
0?
0C
#137530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#137540000000
0!
0*
09
0>
0C
#137550000000
1!
1*
19
1>
1C
#137560000000
0!
0*
09
0>
0C
#137570000000
1!
1*
19
1>
1C
#137580000000
0!
0*
09
0>
0C
#137590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#137600000000
0!
0*
09
0>
0C
#137610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#137620000000
0!
0*
09
0>
0C
#137630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#137640000000
0!
0*
09
0>
0C
#137650000000
1!
1*
b10 6
19
1>
1C
b10 G
#137660000000
0!
0*
09
0>
0C
#137670000000
1!
1*
b11 6
19
1>
1C
b11 G
#137680000000
0!
0*
09
0>
0C
#137690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#137700000000
0!
0*
09
0>
0C
#137710000000
1!
1*
b101 6
19
1>
1C
b101 G
#137720000000
0!
0*
09
0>
0C
#137730000000
1!
1*
b110 6
19
1>
1C
b110 G
#137740000000
0!
0*
09
0>
0C
#137750000000
1!
1*
b111 6
19
1>
1C
b111 G
#137760000000
0!
0*
09
0>
0C
#137770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#137780000000
0!
0*
09
0>
0C
#137790000000
1!
1*
b1 6
19
1>
1C
b1 G
#137800000000
0!
0*
09
0>
0C
#137810000000
1!
1*
b10 6
19
1>
1C
b10 G
#137820000000
0!
0*
09
0>
0C
#137830000000
1!
1*
b11 6
19
1>
1C
b11 G
#137840000000
0!
0*
09
0>
0C
#137850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#137860000000
0!
0*
09
0>
0C
#137870000000
1!
1*
b101 6
19
1>
1C
b101 G
#137880000000
0!
0*
09
0>
0C
#137890000000
1!
1*
b110 6
19
1>
1C
b110 G
#137900000000
0!
0*
09
0>
0C
#137910000000
1!
1*
b111 6
19
1>
1C
b111 G
#137920000000
0!
0*
09
0>
0C
#137930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#137940000000
0!
0*
09
0>
0C
#137950000000
1!
1*
b1 6
19
1>
1C
b1 G
#137960000000
0!
0*
09
0>
0C
#137970000000
1!
1*
b10 6
19
1>
1C
b10 G
#137980000000
0!
0*
09
0>
0C
#137990000000
1!
1*
b11 6
19
1>
1C
b11 G
#138000000000
0!
0*
09
0>
0C
#138010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#138020000000
0!
0*
09
0>
0C
#138030000000
1!
1*
b101 6
19
1>
1C
b101 G
#138040000000
0!
0*
09
0>
0C
#138050000000
1!
1*
b110 6
19
1>
1C
b110 G
#138060000000
0!
0*
09
0>
0C
#138070000000
1!
1*
b111 6
19
1>
1C
b111 G
#138080000000
0!
1"
0*
1+
09
1:
0>
0C
#138090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#138100000000
0!
0*
09
0>
0C
#138110000000
1!
1*
b1 6
19
1>
1C
b1 G
#138120000000
0!
0*
09
0>
0C
#138130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#138140000000
0!
0*
09
0>
0C
#138150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#138160000000
0!
0*
09
0>
0C
#138170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#138180000000
0!
0*
09
0>
0C
#138190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#138200000000
0!
0#
0*
0,
09
0>
0?
0C
#138210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#138220000000
0!
0*
09
0>
0C
#138230000000
1!
1*
19
1>
1C
#138240000000
0!
0*
09
0>
0C
#138250000000
1!
1*
19
1>
1C
#138260000000
0!
0*
09
0>
0C
#138270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#138280000000
0!
0*
09
0>
0C
#138290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#138300000000
0!
0*
09
0>
0C
#138310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#138320000000
0!
0*
09
0>
0C
#138330000000
1!
1*
b10 6
19
1>
1C
b10 G
#138340000000
0!
0*
09
0>
0C
#138350000000
1!
1*
b11 6
19
1>
1C
b11 G
#138360000000
0!
0*
09
0>
0C
#138370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#138380000000
0!
0*
09
0>
0C
#138390000000
1!
1*
b101 6
19
1>
1C
b101 G
#138400000000
0!
0*
09
0>
0C
#138410000000
1!
1*
b110 6
19
1>
1C
b110 G
#138420000000
0!
0*
09
0>
0C
#138430000000
1!
1*
b111 6
19
1>
1C
b111 G
#138440000000
0!
0*
09
0>
0C
#138450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#138460000000
0!
0*
09
0>
0C
#138470000000
1!
1*
b1 6
19
1>
1C
b1 G
#138480000000
0!
0*
09
0>
0C
#138490000000
1!
1*
b10 6
19
1>
1C
b10 G
#138500000000
0!
0*
09
0>
0C
#138510000000
1!
1*
b11 6
19
1>
1C
b11 G
#138520000000
0!
0*
09
0>
0C
#138530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#138540000000
0!
0*
09
0>
0C
#138550000000
1!
1*
b101 6
19
1>
1C
b101 G
#138560000000
0!
0*
09
0>
0C
#138570000000
1!
1*
b110 6
19
1>
1C
b110 G
#138580000000
0!
0*
09
0>
0C
#138590000000
1!
1*
b111 6
19
1>
1C
b111 G
#138600000000
0!
0*
09
0>
0C
#138610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#138620000000
0!
0*
09
0>
0C
#138630000000
1!
1*
b1 6
19
1>
1C
b1 G
#138640000000
0!
0*
09
0>
0C
#138650000000
1!
1*
b10 6
19
1>
1C
b10 G
#138660000000
0!
0*
09
0>
0C
#138670000000
1!
1*
b11 6
19
1>
1C
b11 G
#138680000000
0!
0*
09
0>
0C
#138690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#138700000000
0!
0*
09
0>
0C
#138710000000
1!
1*
b101 6
19
1>
1C
b101 G
#138720000000
0!
0*
09
0>
0C
#138730000000
1!
1*
b110 6
19
1>
1C
b110 G
#138740000000
0!
0*
09
0>
0C
#138750000000
1!
1*
b111 6
19
1>
1C
b111 G
#138760000000
0!
1"
0*
1+
09
1:
0>
0C
#138770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#138780000000
0!
0*
09
0>
0C
#138790000000
1!
1*
b1 6
19
1>
1C
b1 G
#138800000000
0!
0*
09
0>
0C
#138810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#138820000000
0!
0*
09
0>
0C
#138830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#138840000000
0!
0*
09
0>
0C
#138850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#138860000000
0!
0*
09
0>
0C
#138870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#138880000000
0!
0#
0*
0,
09
0>
0?
0C
#138890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#138900000000
0!
0*
09
0>
0C
#138910000000
1!
1*
19
1>
1C
#138920000000
0!
0*
09
0>
0C
#138930000000
1!
1*
19
1>
1C
#138940000000
0!
0*
09
0>
0C
#138950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#138960000000
0!
0*
09
0>
0C
#138970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#138980000000
0!
0*
09
0>
0C
#138990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#139000000000
0!
0*
09
0>
0C
#139010000000
1!
1*
b10 6
19
1>
1C
b10 G
#139020000000
0!
0*
09
0>
0C
#139030000000
1!
1*
b11 6
19
1>
1C
b11 G
#139040000000
0!
0*
09
0>
0C
#139050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#139060000000
0!
0*
09
0>
0C
#139070000000
1!
1*
b101 6
19
1>
1C
b101 G
#139080000000
0!
0*
09
0>
0C
#139090000000
1!
1*
b110 6
19
1>
1C
b110 G
#139100000000
0!
0*
09
0>
0C
#139110000000
1!
1*
b111 6
19
1>
1C
b111 G
#139120000000
0!
0*
09
0>
0C
#139130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#139140000000
0!
0*
09
0>
0C
#139150000000
1!
1*
b1 6
19
1>
1C
b1 G
#139160000000
0!
0*
09
0>
0C
#139170000000
1!
1*
b10 6
19
1>
1C
b10 G
#139180000000
0!
0*
09
0>
0C
#139190000000
1!
1*
b11 6
19
1>
1C
b11 G
#139200000000
0!
0*
09
0>
0C
#139210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#139220000000
0!
0*
09
0>
0C
#139230000000
1!
1*
b101 6
19
1>
1C
b101 G
#139240000000
0!
0*
09
0>
0C
#139250000000
1!
1*
b110 6
19
1>
1C
b110 G
#139260000000
0!
0*
09
0>
0C
#139270000000
1!
1*
b111 6
19
1>
1C
b111 G
#139280000000
0!
0*
09
0>
0C
#139290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#139300000000
0!
0*
09
0>
0C
#139310000000
1!
1*
b1 6
19
1>
1C
b1 G
#139320000000
0!
0*
09
0>
0C
#139330000000
1!
1*
b10 6
19
1>
1C
b10 G
#139340000000
0!
0*
09
0>
0C
#139350000000
1!
1*
b11 6
19
1>
1C
b11 G
#139360000000
0!
0*
09
0>
0C
#139370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#139380000000
0!
0*
09
0>
0C
#139390000000
1!
1*
b101 6
19
1>
1C
b101 G
#139400000000
0!
0*
09
0>
0C
#139410000000
1!
1*
b110 6
19
1>
1C
b110 G
#139420000000
0!
0*
09
0>
0C
#139430000000
1!
1*
b111 6
19
1>
1C
b111 G
#139440000000
0!
1"
0*
1+
09
1:
0>
0C
#139450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#139460000000
0!
0*
09
0>
0C
#139470000000
1!
1*
b1 6
19
1>
1C
b1 G
#139480000000
0!
0*
09
0>
0C
#139490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#139500000000
0!
0*
09
0>
0C
#139510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#139520000000
0!
0*
09
0>
0C
#139530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#139540000000
0!
0*
09
0>
0C
#139550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#139560000000
0!
0#
0*
0,
09
0>
0?
0C
#139570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#139580000000
0!
0*
09
0>
0C
#139590000000
1!
1*
19
1>
1C
#139600000000
0!
0*
09
0>
0C
#139610000000
1!
1*
19
1>
1C
#139620000000
0!
0*
09
0>
0C
#139630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#139640000000
0!
0*
09
0>
0C
#139650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#139660000000
0!
0*
09
0>
0C
#139670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#139680000000
0!
0*
09
0>
0C
#139690000000
1!
1*
b10 6
19
1>
1C
b10 G
#139700000000
0!
0*
09
0>
0C
#139710000000
1!
1*
b11 6
19
1>
1C
b11 G
#139720000000
0!
0*
09
0>
0C
#139730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#139740000000
0!
0*
09
0>
0C
#139750000000
1!
1*
b101 6
19
1>
1C
b101 G
#139760000000
0!
0*
09
0>
0C
#139770000000
1!
1*
b110 6
19
1>
1C
b110 G
#139780000000
0!
0*
09
0>
0C
#139790000000
1!
1*
b111 6
19
1>
1C
b111 G
#139800000000
0!
0*
09
0>
0C
#139810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#139820000000
0!
0*
09
0>
0C
#139830000000
1!
1*
b1 6
19
1>
1C
b1 G
#139840000000
0!
0*
09
0>
0C
#139850000000
1!
1*
b10 6
19
1>
1C
b10 G
#139860000000
0!
0*
09
0>
0C
#139870000000
1!
1*
b11 6
19
1>
1C
b11 G
#139880000000
0!
0*
09
0>
0C
#139890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#139900000000
0!
0*
09
0>
0C
#139910000000
1!
1*
b101 6
19
1>
1C
b101 G
#139920000000
0!
0*
09
0>
0C
#139930000000
1!
1*
b110 6
19
1>
1C
b110 G
#139940000000
0!
0*
09
0>
0C
#139950000000
1!
1*
b111 6
19
1>
1C
b111 G
#139960000000
0!
0*
09
0>
0C
#139970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#139980000000
0!
0*
09
0>
0C
#139990000000
1!
1*
b1 6
19
1>
1C
b1 G
#140000000000
0!
0*
09
0>
0C
#140010000000
1!
1*
b10 6
19
1>
1C
b10 G
#140020000000
0!
0*
09
0>
0C
#140030000000
1!
1*
b11 6
19
1>
1C
b11 G
#140040000000
0!
0*
09
0>
0C
#140050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#140060000000
0!
0*
09
0>
0C
#140070000000
1!
1*
b101 6
19
1>
1C
b101 G
#140080000000
0!
0*
09
0>
0C
#140090000000
1!
1*
b110 6
19
1>
1C
b110 G
#140100000000
0!
0*
09
0>
0C
#140110000000
1!
1*
b111 6
19
1>
1C
b111 G
#140120000000
0!
1"
0*
1+
09
1:
0>
0C
#140130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#140140000000
0!
0*
09
0>
0C
#140150000000
1!
1*
b1 6
19
1>
1C
b1 G
#140160000000
0!
0*
09
0>
0C
#140170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#140180000000
0!
0*
09
0>
0C
#140190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#140200000000
0!
0*
09
0>
0C
#140210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#140220000000
0!
0*
09
0>
0C
#140230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#140240000000
0!
0#
0*
0,
09
0>
0?
0C
#140250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#140260000000
0!
0*
09
0>
0C
#140270000000
1!
1*
19
1>
1C
#140280000000
0!
0*
09
0>
0C
#140290000000
1!
1*
19
1>
1C
#140300000000
0!
0*
09
0>
0C
#140310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#140320000000
0!
0*
09
0>
0C
#140330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#140340000000
0!
0*
09
0>
0C
#140350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#140360000000
0!
0*
09
0>
0C
#140370000000
1!
1*
b10 6
19
1>
1C
b10 G
#140380000000
0!
0*
09
0>
0C
#140390000000
1!
1*
b11 6
19
1>
1C
b11 G
#140400000000
0!
0*
09
0>
0C
#140410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#140420000000
0!
0*
09
0>
0C
#140430000000
1!
1*
b101 6
19
1>
1C
b101 G
#140440000000
0!
0*
09
0>
0C
#140450000000
1!
1*
b110 6
19
1>
1C
b110 G
#140460000000
0!
0*
09
0>
0C
#140470000000
1!
1*
b111 6
19
1>
1C
b111 G
#140480000000
0!
0*
09
0>
0C
#140490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#140500000000
0!
0*
09
0>
0C
#140510000000
1!
1*
b1 6
19
1>
1C
b1 G
#140520000000
0!
0*
09
0>
0C
#140530000000
1!
1*
b10 6
19
1>
1C
b10 G
#140540000000
0!
0*
09
0>
0C
#140550000000
1!
1*
b11 6
19
1>
1C
b11 G
#140560000000
0!
0*
09
0>
0C
#140570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#140580000000
0!
0*
09
0>
0C
#140590000000
1!
1*
b101 6
19
1>
1C
b101 G
#140600000000
0!
0*
09
0>
0C
#140610000000
1!
1*
b110 6
19
1>
1C
b110 G
#140620000000
0!
0*
09
0>
0C
#140630000000
1!
1*
b111 6
19
1>
1C
b111 G
#140640000000
0!
0*
09
0>
0C
#140650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#140660000000
0!
0*
09
0>
0C
#140670000000
1!
1*
b1 6
19
1>
1C
b1 G
#140680000000
0!
0*
09
0>
0C
#140690000000
1!
1*
b10 6
19
1>
1C
b10 G
#140700000000
0!
0*
09
0>
0C
#140710000000
1!
1*
b11 6
19
1>
1C
b11 G
#140720000000
0!
0*
09
0>
0C
#140730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#140740000000
0!
0*
09
0>
0C
#140750000000
1!
1*
b101 6
19
1>
1C
b101 G
#140760000000
0!
0*
09
0>
0C
#140770000000
1!
1*
b110 6
19
1>
1C
b110 G
#140780000000
0!
0*
09
0>
0C
#140790000000
1!
1*
b111 6
19
1>
1C
b111 G
#140800000000
0!
1"
0*
1+
09
1:
0>
0C
#140810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#140820000000
0!
0*
09
0>
0C
#140830000000
1!
1*
b1 6
19
1>
1C
b1 G
#140840000000
0!
0*
09
0>
0C
#140850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#140860000000
0!
0*
09
0>
0C
#140870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#140880000000
0!
0*
09
0>
0C
#140890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#140900000000
0!
0*
09
0>
0C
#140910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#140920000000
0!
0#
0*
0,
09
0>
0?
0C
#140930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#140940000000
0!
0*
09
0>
0C
#140950000000
1!
1*
19
1>
1C
#140960000000
0!
0*
09
0>
0C
#140970000000
1!
1*
19
1>
1C
#140980000000
0!
0*
09
0>
0C
#140990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#141000000000
0!
0*
09
0>
0C
#141010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#141020000000
0!
0*
09
0>
0C
#141030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#141040000000
0!
0*
09
0>
0C
#141050000000
1!
1*
b10 6
19
1>
1C
b10 G
#141060000000
0!
0*
09
0>
0C
#141070000000
1!
1*
b11 6
19
1>
1C
b11 G
#141080000000
0!
0*
09
0>
0C
#141090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#141100000000
0!
0*
09
0>
0C
#141110000000
1!
1*
b101 6
19
1>
1C
b101 G
#141120000000
0!
0*
09
0>
0C
#141130000000
1!
1*
b110 6
19
1>
1C
b110 G
#141140000000
0!
0*
09
0>
0C
#141150000000
1!
1*
b111 6
19
1>
1C
b111 G
#141160000000
0!
0*
09
0>
0C
#141170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#141180000000
0!
0*
09
0>
0C
#141190000000
1!
1*
b1 6
19
1>
1C
b1 G
#141200000000
0!
0*
09
0>
0C
#141210000000
1!
1*
b10 6
19
1>
1C
b10 G
#141220000000
0!
0*
09
0>
0C
#141230000000
1!
1*
b11 6
19
1>
1C
b11 G
#141240000000
0!
0*
09
0>
0C
#141250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#141260000000
0!
0*
09
0>
0C
#141270000000
1!
1*
b101 6
19
1>
1C
b101 G
#141280000000
0!
0*
09
0>
0C
#141290000000
1!
1*
b110 6
19
1>
1C
b110 G
#141300000000
0!
0*
09
0>
0C
#141310000000
1!
1*
b111 6
19
1>
1C
b111 G
#141320000000
0!
0*
09
0>
0C
#141330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#141340000000
0!
0*
09
0>
0C
#141350000000
1!
1*
b1 6
19
1>
1C
b1 G
#141360000000
0!
0*
09
0>
0C
#141370000000
1!
1*
b10 6
19
1>
1C
b10 G
#141380000000
0!
0*
09
0>
0C
#141390000000
1!
1*
b11 6
19
1>
1C
b11 G
#141400000000
0!
0*
09
0>
0C
#141410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#141420000000
0!
0*
09
0>
0C
#141430000000
1!
1*
b101 6
19
1>
1C
b101 G
#141440000000
0!
0*
09
0>
0C
#141450000000
1!
1*
b110 6
19
1>
1C
b110 G
#141460000000
0!
0*
09
0>
0C
#141470000000
1!
1*
b111 6
19
1>
1C
b111 G
#141480000000
0!
1"
0*
1+
09
1:
0>
0C
#141490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#141500000000
0!
0*
09
0>
0C
#141510000000
1!
1*
b1 6
19
1>
1C
b1 G
#141520000000
0!
0*
09
0>
0C
#141530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#141540000000
0!
0*
09
0>
0C
#141550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#141560000000
0!
0*
09
0>
0C
#141570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#141580000000
0!
0*
09
0>
0C
#141590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#141600000000
0!
0#
0*
0,
09
0>
0?
0C
#141610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#141620000000
0!
0*
09
0>
0C
#141630000000
1!
1*
19
1>
1C
#141640000000
0!
0*
09
0>
0C
#141650000000
1!
1*
19
1>
1C
#141660000000
0!
0*
09
0>
0C
#141670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#141680000000
0!
0*
09
0>
0C
#141690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#141700000000
0!
0*
09
0>
0C
#141710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#141720000000
0!
0*
09
0>
0C
#141730000000
1!
1*
b10 6
19
1>
1C
b10 G
#141740000000
0!
0*
09
0>
0C
#141750000000
1!
1*
b11 6
19
1>
1C
b11 G
#141760000000
0!
0*
09
0>
0C
#141770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#141780000000
0!
0*
09
0>
0C
#141790000000
1!
1*
b101 6
19
1>
1C
b101 G
#141800000000
0!
0*
09
0>
0C
#141810000000
1!
1*
b110 6
19
1>
1C
b110 G
#141820000000
0!
0*
09
0>
0C
#141830000000
1!
1*
b111 6
19
1>
1C
b111 G
#141840000000
0!
0*
09
0>
0C
#141850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#141860000000
0!
0*
09
0>
0C
#141870000000
1!
1*
b1 6
19
1>
1C
b1 G
#141880000000
0!
0*
09
0>
0C
#141890000000
1!
1*
b10 6
19
1>
1C
b10 G
#141900000000
0!
0*
09
0>
0C
#141910000000
1!
1*
b11 6
19
1>
1C
b11 G
#141920000000
0!
0*
09
0>
0C
#141930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#141940000000
0!
0*
09
0>
0C
#141950000000
1!
1*
b101 6
19
1>
1C
b101 G
#141960000000
0!
0*
09
0>
0C
#141970000000
1!
1*
b110 6
19
1>
1C
b110 G
#141980000000
0!
0*
09
0>
0C
#141990000000
1!
1*
b111 6
19
1>
1C
b111 G
#142000000000
0!
0*
09
0>
0C
#142010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#142020000000
0!
0*
09
0>
0C
#142030000000
1!
1*
b1 6
19
1>
1C
b1 G
#142040000000
0!
0*
09
0>
0C
#142050000000
1!
1*
b10 6
19
1>
1C
b10 G
#142060000000
0!
0*
09
0>
0C
#142070000000
1!
1*
b11 6
19
1>
1C
b11 G
#142080000000
0!
0*
09
0>
0C
#142090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#142100000000
0!
0*
09
0>
0C
#142110000000
1!
1*
b101 6
19
1>
1C
b101 G
#142120000000
0!
0*
09
0>
0C
#142130000000
1!
1*
b110 6
19
1>
1C
b110 G
#142140000000
0!
0*
09
0>
0C
#142150000000
1!
1*
b111 6
19
1>
1C
b111 G
#142160000000
0!
1"
0*
1+
09
1:
0>
0C
#142170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#142180000000
0!
0*
09
0>
0C
#142190000000
1!
1*
b1 6
19
1>
1C
b1 G
#142200000000
0!
0*
09
0>
0C
#142210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#142220000000
0!
0*
09
0>
0C
#142230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#142240000000
0!
0*
09
0>
0C
#142250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#142260000000
0!
0*
09
0>
0C
#142270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#142280000000
0!
0#
0*
0,
09
0>
0?
0C
#142290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#142300000000
0!
0*
09
0>
0C
#142310000000
1!
1*
19
1>
1C
#142320000000
0!
0*
09
0>
0C
#142330000000
1!
1*
19
1>
1C
#142340000000
0!
0*
09
0>
0C
#142350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#142360000000
0!
0*
09
0>
0C
#142370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#142380000000
0!
0*
09
0>
0C
#142390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#142400000000
0!
0*
09
0>
0C
#142410000000
1!
1*
b10 6
19
1>
1C
b10 G
#142420000000
0!
0*
09
0>
0C
#142430000000
1!
1*
b11 6
19
1>
1C
b11 G
#142440000000
0!
0*
09
0>
0C
#142450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#142460000000
0!
0*
09
0>
0C
#142470000000
1!
1*
b101 6
19
1>
1C
b101 G
#142480000000
0!
0*
09
0>
0C
#142490000000
1!
1*
b110 6
19
1>
1C
b110 G
#142500000000
0!
0*
09
0>
0C
#142510000000
1!
1*
b111 6
19
1>
1C
b111 G
#142520000000
0!
0*
09
0>
0C
#142530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#142540000000
0!
0*
09
0>
0C
#142550000000
1!
1*
b1 6
19
1>
1C
b1 G
#142560000000
0!
0*
09
0>
0C
#142570000000
1!
1*
b10 6
19
1>
1C
b10 G
#142580000000
0!
0*
09
0>
0C
#142590000000
1!
1*
b11 6
19
1>
1C
b11 G
#142600000000
0!
0*
09
0>
0C
#142610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#142620000000
0!
0*
09
0>
0C
#142630000000
1!
1*
b101 6
19
1>
1C
b101 G
#142640000000
0!
0*
09
0>
0C
#142650000000
1!
1*
b110 6
19
1>
1C
b110 G
#142660000000
0!
0*
09
0>
0C
#142670000000
1!
1*
b111 6
19
1>
1C
b111 G
#142680000000
0!
0*
09
0>
0C
#142690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#142700000000
0!
0*
09
0>
0C
#142710000000
1!
1*
b1 6
19
1>
1C
b1 G
#142720000000
0!
0*
09
0>
0C
#142730000000
1!
1*
b10 6
19
1>
1C
b10 G
#142740000000
0!
0*
09
0>
0C
#142750000000
1!
1*
b11 6
19
1>
1C
b11 G
#142760000000
0!
0*
09
0>
0C
#142770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#142780000000
0!
0*
09
0>
0C
#142790000000
1!
1*
b101 6
19
1>
1C
b101 G
#142800000000
0!
0*
09
0>
0C
#142810000000
1!
1*
b110 6
19
1>
1C
b110 G
#142820000000
0!
0*
09
0>
0C
#142830000000
1!
1*
b111 6
19
1>
1C
b111 G
#142840000000
0!
1"
0*
1+
09
1:
0>
0C
#142850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#142860000000
0!
0*
09
0>
0C
#142870000000
1!
1*
b1 6
19
1>
1C
b1 G
#142880000000
0!
0*
09
0>
0C
#142890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#142900000000
0!
0*
09
0>
0C
#142910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#142920000000
0!
0*
09
0>
0C
#142930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#142940000000
0!
0*
09
0>
0C
#142950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#142960000000
0!
0#
0*
0,
09
0>
0?
0C
#142970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#142980000000
0!
0*
09
0>
0C
#142990000000
1!
1*
19
1>
1C
#143000000000
0!
0*
09
0>
0C
#143010000000
1!
1*
19
1>
1C
#143020000000
0!
0*
09
0>
0C
#143030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#143040000000
0!
0*
09
0>
0C
#143050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#143060000000
0!
0*
09
0>
0C
#143070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#143080000000
0!
0*
09
0>
0C
#143090000000
1!
1*
b10 6
19
1>
1C
b10 G
#143100000000
0!
0*
09
0>
0C
#143110000000
1!
1*
b11 6
19
1>
1C
b11 G
#143120000000
0!
0*
09
0>
0C
#143130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#143140000000
0!
0*
09
0>
0C
#143150000000
1!
1*
b101 6
19
1>
1C
b101 G
#143160000000
0!
0*
09
0>
0C
#143170000000
1!
1*
b110 6
19
1>
1C
b110 G
#143180000000
0!
0*
09
0>
0C
#143190000000
1!
1*
b111 6
19
1>
1C
b111 G
#143200000000
0!
0*
09
0>
0C
#143210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#143220000000
0!
0*
09
0>
0C
#143230000000
1!
1*
b1 6
19
1>
1C
b1 G
#143240000000
0!
0*
09
0>
0C
#143250000000
1!
1*
b10 6
19
1>
1C
b10 G
#143260000000
0!
0*
09
0>
0C
#143270000000
1!
1*
b11 6
19
1>
1C
b11 G
#143280000000
0!
0*
09
0>
0C
#143290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#143300000000
0!
0*
09
0>
0C
#143310000000
1!
1*
b101 6
19
1>
1C
b101 G
#143320000000
0!
0*
09
0>
0C
#143330000000
1!
1*
b110 6
19
1>
1C
b110 G
#143340000000
0!
0*
09
0>
0C
#143350000000
1!
1*
b111 6
19
1>
1C
b111 G
#143360000000
0!
0*
09
0>
0C
#143370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#143380000000
0!
0*
09
0>
0C
#143390000000
1!
1*
b1 6
19
1>
1C
b1 G
#143400000000
0!
0*
09
0>
0C
#143410000000
1!
1*
b10 6
19
1>
1C
b10 G
#143420000000
0!
0*
09
0>
0C
#143430000000
1!
1*
b11 6
19
1>
1C
b11 G
#143440000000
0!
0*
09
0>
0C
#143450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#143460000000
0!
0*
09
0>
0C
#143470000000
1!
1*
b101 6
19
1>
1C
b101 G
#143480000000
0!
0*
09
0>
0C
#143490000000
1!
1*
b110 6
19
1>
1C
b110 G
#143500000000
0!
0*
09
0>
0C
#143510000000
1!
1*
b111 6
19
1>
1C
b111 G
#143520000000
0!
1"
0*
1+
09
1:
0>
0C
#143530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#143540000000
0!
0*
09
0>
0C
#143550000000
1!
1*
b1 6
19
1>
1C
b1 G
#143560000000
0!
0*
09
0>
0C
#143570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#143580000000
0!
0*
09
0>
0C
#143590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#143600000000
0!
0*
09
0>
0C
#143610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#143620000000
0!
0*
09
0>
0C
#143630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#143640000000
0!
0#
0*
0,
09
0>
0?
0C
#143650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#143660000000
0!
0*
09
0>
0C
#143670000000
1!
1*
19
1>
1C
#143680000000
0!
0*
09
0>
0C
#143690000000
1!
1*
19
1>
1C
#143700000000
0!
0*
09
0>
0C
#143710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#143720000000
0!
0*
09
0>
0C
#143730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#143740000000
0!
0*
09
0>
0C
#143750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#143760000000
0!
0*
09
0>
0C
#143770000000
1!
1*
b10 6
19
1>
1C
b10 G
#143780000000
0!
0*
09
0>
0C
#143790000000
1!
1*
b11 6
19
1>
1C
b11 G
#143800000000
0!
0*
09
0>
0C
#143810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#143820000000
0!
0*
09
0>
0C
#143830000000
1!
1*
b101 6
19
1>
1C
b101 G
#143840000000
0!
0*
09
0>
0C
#143850000000
1!
1*
b110 6
19
1>
1C
b110 G
#143860000000
0!
0*
09
0>
0C
#143870000000
1!
1*
b111 6
19
1>
1C
b111 G
#143880000000
0!
0*
09
0>
0C
#143890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#143900000000
0!
0*
09
0>
0C
#143910000000
1!
1*
b1 6
19
1>
1C
b1 G
#143920000000
0!
0*
09
0>
0C
#143930000000
1!
1*
b10 6
19
1>
1C
b10 G
#143940000000
0!
0*
09
0>
0C
#143950000000
1!
1*
b11 6
19
1>
1C
b11 G
#143960000000
0!
0*
09
0>
0C
#143970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#143980000000
0!
0*
09
0>
0C
#143990000000
1!
1*
b101 6
19
1>
1C
b101 G
#144000000000
0!
0*
09
0>
0C
#144010000000
1!
1*
b110 6
19
1>
1C
b110 G
#144020000000
0!
0*
09
0>
0C
#144030000000
1!
1*
b111 6
19
1>
1C
b111 G
#144040000000
0!
0*
09
0>
0C
#144050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#144060000000
0!
0*
09
0>
0C
#144070000000
1!
1*
b1 6
19
1>
1C
b1 G
#144080000000
0!
0*
09
0>
0C
#144090000000
1!
1*
b10 6
19
1>
1C
b10 G
#144100000000
0!
0*
09
0>
0C
#144110000000
1!
1*
b11 6
19
1>
1C
b11 G
#144120000000
0!
0*
09
0>
0C
#144130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#144140000000
0!
0*
09
0>
0C
#144150000000
1!
1*
b101 6
19
1>
1C
b101 G
#144160000000
0!
0*
09
0>
0C
#144170000000
1!
1*
b110 6
19
1>
1C
b110 G
#144180000000
0!
0*
09
0>
0C
#144190000000
1!
1*
b111 6
19
1>
1C
b111 G
#144200000000
0!
1"
0*
1+
09
1:
0>
0C
#144210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#144220000000
0!
0*
09
0>
0C
#144230000000
1!
1*
b1 6
19
1>
1C
b1 G
#144240000000
0!
0*
09
0>
0C
#144250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#144260000000
0!
0*
09
0>
0C
#144270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#144280000000
0!
0*
09
0>
0C
#144290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#144300000000
0!
0*
09
0>
0C
#144310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#144320000000
0!
0#
0*
0,
09
0>
0?
0C
#144330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#144340000000
0!
0*
09
0>
0C
#144350000000
1!
1*
19
1>
1C
#144360000000
0!
0*
09
0>
0C
#144370000000
1!
1*
19
1>
1C
#144380000000
0!
0*
09
0>
0C
#144390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#144400000000
0!
0*
09
0>
0C
#144410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#144420000000
0!
0*
09
0>
0C
#144430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#144440000000
0!
0*
09
0>
0C
#144450000000
1!
1*
b10 6
19
1>
1C
b10 G
#144460000000
0!
0*
09
0>
0C
#144470000000
1!
1*
b11 6
19
1>
1C
b11 G
#144480000000
0!
0*
09
0>
0C
#144490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#144500000000
0!
0*
09
0>
0C
#144510000000
1!
1*
b101 6
19
1>
1C
b101 G
#144520000000
0!
0*
09
0>
0C
#144530000000
1!
1*
b110 6
19
1>
1C
b110 G
#144540000000
0!
0*
09
0>
0C
#144550000000
1!
1*
b111 6
19
1>
1C
b111 G
#144560000000
0!
0*
09
0>
0C
#144570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#144580000000
0!
0*
09
0>
0C
#144590000000
1!
1*
b1 6
19
1>
1C
b1 G
#144600000000
0!
0*
09
0>
0C
#144610000000
1!
1*
b10 6
19
1>
1C
b10 G
#144620000000
0!
0*
09
0>
0C
#144630000000
1!
1*
b11 6
19
1>
1C
b11 G
#144640000000
0!
0*
09
0>
0C
#144650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#144660000000
0!
0*
09
0>
0C
#144670000000
1!
1*
b101 6
19
1>
1C
b101 G
#144680000000
0!
0*
09
0>
0C
#144690000000
1!
1*
b110 6
19
1>
1C
b110 G
#144700000000
0!
0*
09
0>
0C
#144710000000
1!
1*
b111 6
19
1>
1C
b111 G
#144720000000
0!
0*
09
0>
0C
#144730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#144740000000
0!
0*
09
0>
0C
#144750000000
1!
1*
b1 6
19
1>
1C
b1 G
#144760000000
0!
0*
09
0>
0C
#144770000000
1!
1*
b10 6
19
1>
1C
b10 G
#144780000000
0!
0*
09
0>
0C
#144790000000
1!
1*
b11 6
19
1>
1C
b11 G
#144800000000
0!
0*
09
0>
0C
#144810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#144820000000
0!
0*
09
0>
0C
#144830000000
1!
1*
b101 6
19
1>
1C
b101 G
#144840000000
0!
0*
09
0>
0C
#144850000000
1!
1*
b110 6
19
1>
1C
b110 G
#144860000000
0!
0*
09
0>
0C
#144870000000
1!
1*
b111 6
19
1>
1C
b111 G
#144880000000
0!
1"
0*
1+
09
1:
0>
0C
#144890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#144900000000
0!
0*
09
0>
0C
#144910000000
1!
1*
b1 6
19
1>
1C
b1 G
#144920000000
0!
0*
09
0>
0C
#144930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#144940000000
0!
0*
09
0>
0C
#144950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#144960000000
0!
0*
09
0>
0C
#144970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#144980000000
0!
0*
09
0>
0C
#144990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#145000000000
0!
0#
0*
0,
09
0>
0?
0C
#145010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#145020000000
0!
0*
09
0>
0C
#145030000000
1!
1*
19
1>
1C
#145040000000
0!
0*
09
0>
0C
#145050000000
1!
1*
19
1>
1C
#145060000000
0!
0*
09
0>
0C
#145070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#145080000000
0!
0*
09
0>
0C
#145090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#145100000000
0!
0*
09
0>
0C
#145110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#145120000000
0!
0*
09
0>
0C
#145130000000
1!
1*
b10 6
19
1>
1C
b10 G
#145140000000
0!
0*
09
0>
0C
#145150000000
1!
1*
b11 6
19
1>
1C
b11 G
#145160000000
0!
0*
09
0>
0C
#145170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#145180000000
0!
0*
09
0>
0C
#145190000000
1!
1*
b101 6
19
1>
1C
b101 G
#145200000000
0!
0*
09
0>
0C
#145210000000
1!
1*
b110 6
19
1>
1C
b110 G
#145220000000
0!
0*
09
0>
0C
#145230000000
1!
1*
b111 6
19
1>
1C
b111 G
#145240000000
0!
0*
09
0>
0C
#145250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#145260000000
0!
0*
09
0>
0C
#145270000000
1!
1*
b1 6
19
1>
1C
b1 G
#145280000000
0!
0*
09
0>
0C
#145290000000
1!
1*
b10 6
19
1>
1C
b10 G
#145300000000
0!
0*
09
0>
0C
#145310000000
1!
1*
b11 6
19
1>
1C
b11 G
#145320000000
0!
0*
09
0>
0C
#145330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#145340000000
0!
0*
09
0>
0C
#145350000000
1!
1*
b101 6
19
1>
1C
b101 G
#145360000000
0!
0*
09
0>
0C
#145370000000
1!
1*
b110 6
19
1>
1C
b110 G
#145380000000
0!
0*
09
0>
0C
#145390000000
1!
1*
b111 6
19
1>
1C
b111 G
#145400000000
0!
0*
09
0>
0C
#145410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#145420000000
0!
0*
09
0>
0C
#145430000000
1!
1*
b1 6
19
1>
1C
b1 G
#145440000000
0!
0*
09
0>
0C
#145450000000
1!
1*
b10 6
19
1>
1C
b10 G
#145460000000
0!
0*
09
0>
0C
#145470000000
1!
1*
b11 6
19
1>
1C
b11 G
#145480000000
0!
0*
09
0>
0C
#145490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#145500000000
0!
0*
09
0>
0C
#145510000000
1!
1*
b101 6
19
1>
1C
b101 G
#145520000000
0!
0*
09
0>
0C
#145530000000
1!
1*
b110 6
19
1>
1C
b110 G
#145540000000
0!
0*
09
0>
0C
#145550000000
1!
1*
b111 6
19
1>
1C
b111 G
#145560000000
0!
1"
0*
1+
09
1:
0>
0C
#145570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#145580000000
0!
0*
09
0>
0C
#145590000000
1!
1*
b1 6
19
1>
1C
b1 G
#145600000000
0!
0*
09
0>
0C
#145610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#145620000000
0!
0*
09
0>
0C
#145630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#145640000000
0!
0*
09
0>
0C
#145650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#145660000000
0!
0*
09
0>
0C
#145670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#145680000000
0!
0#
0*
0,
09
0>
0?
0C
#145690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#145700000000
0!
0*
09
0>
0C
#145710000000
1!
1*
19
1>
1C
#145720000000
0!
0*
09
0>
0C
#145730000000
1!
1*
19
1>
1C
#145740000000
0!
0*
09
0>
0C
#145750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#145760000000
0!
0*
09
0>
0C
#145770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#145780000000
0!
0*
09
0>
0C
#145790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#145800000000
0!
0*
09
0>
0C
#145810000000
1!
1*
b10 6
19
1>
1C
b10 G
#145820000000
0!
0*
09
0>
0C
#145830000000
1!
1*
b11 6
19
1>
1C
b11 G
#145840000000
0!
0*
09
0>
0C
#145850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#145860000000
0!
0*
09
0>
0C
#145870000000
1!
1*
b101 6
19
1>
1C
b101 G
#145880000000
0!
0*
09
0>
0C
#145890000000
1!
1*
b110 6
19
1>
1C
b110 G
#145900000000
0!
0*
09
0>
0C
#145910000000
1!
1*
b111 6
19
1>
1C
b111 G
#145920000000
0!
0*
09
0>
0C
#145930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#145940000000
0!
0*
09
0>
0C
#145950000000
1!
1*
b1 6
19
1>
1C
b1 G
#145960000000
0!
0*
09
0>
0C
#145970000000
1!
1*
b10 6
19
1>
1C
b10 G
#145980000000
0!
0*
09
0>
0C
#145990000000
1!
1*
b11 6
19
1>
1C
b11 G
#146000000000
0!
0*
09
0>
0C
#146010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#146020000000
0!
0*
09
0>
0C
#146030000000
1!
1*
b101 6
19
1>
1C
b101 G
#146040000000
0!
0*
09
0>
0C
#146050000000
1!
1*
b110 6
19
1>
1C
b110 G
#146060000000
0!
0*
09
0>
0C
#146070000000
1!
1*
b111 6
19
1>
1C
b111 G
#146080000000
0!
0*
09
0>
0C
#146090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#146100000000
0!
0*
09
0>
0C
#146110000000
1!
1*
b1 6
19
1>
1C
b1 G
#146120000000
0!
0*
09
0>
0C
#146130000000
1!
1*
b10 6
19
1>
1C
b10 G
#146140000000
0!
0*
09
0>
0C
#146150000000
1!
1*
b11 6
19
1>
1C
b11 G
#146160000000
0!
0*
09
0>
0C
#146170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#146180000000
0!
0*
09
0>
0C
#146190000000
1!
1*
b101 6
19
1>
1C
b101 G
#146200000000
0!
0*
09
0>
0C
#146210000000
1!
1*
b110 6
19
1>
1C
b110 G
#146220000000
0!
0*
09
0>
0C
#146230000000
1!
1*
b111 6
19
1>
1C
b111 G
#146240000000
0!
1"
0*
1+
09
1:
0>
0C
#146250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#146260000000
0!
0*
09
0>
0C
#146270000000
1!
1*
b1 6
19
1>
1C
b1 G
#146280000000
0!
0*
09
0>
0C
#146290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#146300000000
0!
0*
09
0>
0C
#146310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#146320000000
0!
0*
09
0>
0C
#146330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#146340000000
0!
0*
09
0>
0C
#146350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#146360000000
0!
0#
0*
0,
09
0>
0?
0C
#146370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#146380000000
0!
0*
09
0>
0C
#146390000000
1!
1*
19
1>
1C
#146400000000
0!
0*
09
0>
0C
#146410000000
1!
1*
19
1>
1C
#146420000000
0!
0*
09
0>
0C
#146430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#146440000000
0!
0*
09
0>
0C
#146450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#146460000000
0!
0*
09
0>
0C
#146470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#146480000000
0!
0*
09
0>
0C
#146490000000
1!
1*
b10 6
19
1>
1C
b10 G
#146500000000
0!
0*
09
0>
0C
#146510000000
1!
1*
b11 6
19
1>
1C
b11 G
#146520000000
0!
0*
09
0>
0C
#146530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#146540000000
0!
0*
09
0>
0C
#146550000000
1!
1*
b101 6
19
1>
1C
b101 G
#146560000000
0!
0*
09
0>
0C
#146570000000
1!
1*
b110 6
19
1>
1C
b110 G
#146580000000
0!
0*
09
0>
0C
#146590000000
1!
1*
b111 6
19
1>
1C
b111 G
#146600000000
0!
0*
09
0>
0C
#146610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#146620000000
0!
0*
09
0>
0C
#146630000000
1!
1*
b1 6
19
1>
1C
b1 G
#146640000000
0!
0*
09
0>
0C
#146650000000
1!
1*
b10 6
19
1>
1C
b10 G
#146660000000
0!
0*
09
0>
0C
#146670000000
1!
1*
b11 6
19
1>
1C
b11 G
#146680000000
0!
0*
09
0>
0C
#146690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#146700000000
0!
0*
09
0>
0C
#146710000000
1!
1*
b101 6
19
1>
1C
b101 G
#146720000000
0!
0*
09
0>
0C
#146730000000
1!
1*
b110 6
19
1>
1C
b110 G
#146740000000
0!
0*
09
0>
0C
#146750000000
1!
1*
b111 6
19
1>
1C
b111 G
#146760000000
0!
0*
09
0>
0C
#146770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#146780000000
0!
0*
09
0>
0C
#146790000000
1!
1*
b1 6
19
1>
1C
b1 G
#146800000000
0!
0*
09
0>
0C
#146810000000
1!
1*
b10 6
19
1>
1C
b10 G
#146820000000
0!
0*
09
0>
0C
#146830000000
1!
1*
b11 6
19
1>
1C
b11 G
#146840000000
0!
0*
09
0>
0C
#146850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#146860000000
0!
0*
09
0>
0C
#146870000000
1!
1*
b101 6
19
1>
1C
b101 G
#146880000000
0!
0*
09
0>
0C
#146890000000
1!
1*
b110 6
19
1>
1C
b110 G
#146900000000
0!
0*
09
0>
0C
#146910000000
1!
1*
b111 6
19
1>
1C
b111 G
#146920000000
0!
1"
0*
1+
09
1:
0>
0C
#146930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#146940000000
0!
0*
09
0>
0C
#146950000000
1!
1*
b1 6
19
1>
1C
b1 G
#146960000000
0!
0*
09
0>
0C
#146970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#146980000000
0!
0*
09
0>
0C
#146990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#147000000000
0!
0*
09
0>
0C
#147010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#147020000000
0!
0*
09
0>
0C
#147030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#147040000000
0!
0#
0*
0,
09
0>
0?
0C
#147050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#147060000000
0!
0*
09
0>
0C
#147070000000
1!
1*
19
1>
1C
#147080000000
0!
0*
09
0>
0C
#147090000000
1!
1*
19
1>
1C
#147100000000
0!
0*
09
0>
0C
#147110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#147120000000
0!
0*
09
0>
0C
#147130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#147140000000
0!
0*
09
0>
0C
#147150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#147160000000
0!
0*
09
0>
0C
#147170000000
1!
1*
b10 6
19
1>
1C
b10 G
#147180000000
0!
0*
09
0>
0C
#147190000000
1!
1*
b11 6
19
1>
1C
b11 G
#147200000000
0!
0*
09
0>
0C
#147210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#147220000000
0!
0*
09
0>
0C
#147230000000
1!
1*
b101 6
19
1>
1C
b101 G
#147240000000
0!
0*
09
0>
0C
#147250000000
1!
1*
b110 6
19
1>
1C
b110 G
#147260000000
0!
0*
09
0>
0C
#147270000000
1!
1*
b111 6
19
1>
1C
b111 G
#147280000000
0!
0*
09
0>
0C
#147290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#147300000000
0!
0*
09
0>
0C
#147310000000
1!
1*
b1 6
19
1>
1C
b1 G
#147320000000
0!
0*
09
0>
0C
#147330000000
1!
1*
b10 6
19
1>
1C
b10 G
#147340000000
0!
0*
09
0>
0C
#147350000000
1!
1*
b11 6
19
1>
1C
b11 G
#147360000000
0!
0*
09
0>
0C
#147370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#147380000000
0!
0*
09
0>
0C
#147390000000
1!
1*
b101 6
19
1>
1C
b101 G
#147400000000
0!
0*
09
0>
0C
#147410000000
1!
1*
b110 6
19
1>
1C
b110 G
#147420000000
0!
0*
09
0>
0C
#147430000000
1!
1*
b111 6
19
1>
1C
b111 G
#147440000000
0!
0*
09
0>
0C
#147450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#147460000000
0!
0*
09
0>
0C
#147470000000
1!
1*
b1 6
19
1>
1C
b1 G
#147480000000
0!
0*
09
0>
0C
#147490000000
1!
1*
b10 6
19
1>
1C
b10 G
#147500000000
0!
0*
09
0>
0C
#147510000000
1!
1*
b11 6
19
1>
1C
b11 G
#147520000000
0!
0*
09
0>
0C
#147530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#147540000000
0!
0*
09
0>
0C
#147550000000
1!
1*
b101 6
19
1>
1C
b101 G
#147560000000
0!
0*
09
0>
0C
#147570000000
1!
1*
b110 6
19
1>
1C
b110 G
#147580000000
0!
0*
09
0>
0C
#147590000000
1!
1*
b111 6
19
1>
1C
b111 G
#147600000000
0!
1"
0*
1+
09
1:
0>
0C
#147610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#147620000000
0!
0*
09
0>
0C
#147630000000
1!
1*
b1 6
19
1>
1C
b1 G
#147640000000
0!
0*
09
0>
0C
#147650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#147660000000
0!
0*
09
0>
0C
#147670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#147680000000
0!
0*
09
0>
0C
#147690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#147700000000
0!
0*
09
0>
0C
#147710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#147720000000
0!
0#
0*
0,
09
0>
0?
0C
#147730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#147740000000
0!
0*
09
0>
0C
#147750000000
1!
1*
19
1>
1C
#147760000000
0!
0*
09
0>
0C
#147770000000
1!
1*
19
1>
1C
#147780000000
0!
0*
09
0>
0C
#147790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#147800000000
0!
0*
09
0>
0C
#147810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#147820000000
0!
0*
09
0>
0C
#147830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#147840000000
0!
0*
09
0>
0C
#147850000000
1!
1*
b10 6
19
1>
1C
b10 G
#147860000000
0!
0*
09
0>
0C
#147870000000
1!
1*
b11 6
19
1>
1C
b11 G
#147880000000
0!
0*
09
0>
0C
#147890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#147900000000
0!
0*
09
0>
0C
#147910000000
1!
1*
b101 6
19
1>
1C
b101 G
#147920000000
0!
0*
09
0>
0C
#147930000000
1!
1*
b110 6
19
1>
1C
b110 G
#147940000000
0!
0*
09
0>
0C
#147950000000
1!
1*
b111 6
19
1>
1C
b111 G
#147960000000
0!
0*
09
0>
0C
#147970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#147980000000
0!
0*
09
0>
0C
#147990000000
1!
1*
b1 6
19
1>
1C
b1 G
#148000000000
0!
0*
09
0>
0C
#148010000000
1!
1*
b10 6
19
1>
1C
b10 G
#148020000000
0!
0*
09
0>
0C
#148030000000
1!
1*
b11 6
19
1>
1C
b11 G
#148040000000
0!
0*
09
0>
0C
#148050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#148060000000
0!
0*
09
0>
0C
#148070000000
1!
1*
b101 6
19
1>
1C
b101 G
#148080000000
0!
0*
09
0>
0C
#148090000000
1!
1*
b110 6
19
1>
1C
b110 G
#148100000000
0!
0*
09
0>
0C
#148110000000
1!
1*
b111 6
19
1>
1C
b111 G
#148120000000
0!
0*
09
0>
0C
#148130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#148140000000
0!
0*
09
0>
0C
#148150000000
1!
1*
b1 6
19
1>
1C
b1 G
#148160000000
0!
0*
09
0>
0C
#148170000000
1!
1*
b10 6
19
1>
1C
b10 G
#148180000000
0!
0*
09
0>
0C
#148190000000
1!
1*
b11 6
19
1>
1C
b11 G
#148200000000
0!
0*
09
0>
0C
#148210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#148220000000
0!
0*
09
0>
0C
#148230000000
1!
1*
b101 6
19
1>
1C
b101 G
#148240000000
0!
0*
09
0>
0C
#148250000000
1!
1*
b110 6
19
1>
1C
b110 G
#148260000000
0!
0*
09
0>
0C
#148270000000
1!
1*
b111 6
19
1>
1C
b111 G
#148280000000
0!
1"
0*
1+
09
1:
0>
0C
#148290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#148300000000
0!
0*
09
0>
0C
#148310000000
1!
1*
b1 6
19
1>
1C
b1 G
#148320000000
0!
0*
09
0>
0C
#148330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#148340000000
0!
0*
09
0>
0C
#148350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#148360000000
0!
0*
09
0>
0C
#148370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#148380000000
0!
0*
09
0>
0C
#148390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#148400000000
0!
0#
0*
0,
09
0>
0?
0C
#148410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#148420000000
0!
0*
09
0>
0C
#148430000000
1!
1*
19
1>
1C
#148440000000
0!
0*
09
0>
0C
#148450000000
1!
1*
19
1>
1C
#148460000000
0!
0*
09
0>
0C
#148470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#148480000000
0!
0*
09
0>
0C
#148490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#148500000000
0!
0*
09
0>
0C
#148510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#148520000000
0!
0*
09
0>
0C
#148530000000
1!
1*
b10 6
19
1>
1C
b10 G
#148540000000
0!
0*
09
0>
0C
#148550000000
1!
1*
b11 6
19
1>
1C
b11 G
#148560000000
0!
0*
09
0>
0C
#148570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#148580000000
0!
0*
09
0>
0C
#148590000000
1!
1*
b101 6
19
1>
1C
b101 G
#148600000000
0!
0*
09
0>
0C
#148610000000
1!
1*
b110 6
19
1>
1C
b110 G
#148620000000
0!
0*
09
0>
0C
#148630000000
1!
1*
b111 6
19
1>
1C
b111 G
#148640000000
0!
0*
09
0>
0C
#148650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#148660000000
0!
0*
09
0>
0C
#148670000000
1!
1*
b1 6
19
1>
1C
b1 G
#148680000000
0!
0*
09
0>
0C
#148690000000
1!
1*
b10 6
19
1>
1C
b10 G
#148700000000
0!
0*
09
0>
0C
#148710000000
1!
1*
b11 6
19
1>
1C
b11 G
#148720000000
0!
0*
09
0>
0C
#148730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#148740000000
0!
0*
09
0>
0C
#148750000000
1!
1*
b101 6
19
1>
1C
b101 G
#148760000000
0!
0*
09
0>
0C
#148770000000
1!
1*
b110 6
19
1>
1C
b110 G
#148780000000
0!
0*
09
0>
0C
#148790000000
1!
1*
b111 6
19
1>
1C
b111 G
#148800000000
0!
0*
09
0>
0C
#148810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#148820000000
0!
0*
09
0>
0C
#148830000000
1!
1*
b1 6
19
1>
1C
b1 G
#148840000000
0!
0*
09
0>
0C
#148850000000
1!
1*
b10 6
19
1>
1C
b10 G
#148860000000
0!
0*
09
0>
0C
#148870000000
1!
1*
b11 6
19
1>
1C
b11 G
#148880000000
0!
0*
09
0>
0C
#148890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#148900000000
0!
0*
09
0>
0C
#148910000000
1!
1*
b101 6
19
1>
1C
b101 G
#148920000000
0!
0*
09
0>
0C
#148930000000
1!
1*
b110 6
19
1>
1C
b110 G
#148940000000
0!
0*
09
0>
0C
#148950000000
1!
1*
b111 6
19
1>
1C
b111 G
#148960000000
0!
1"
0*
1+
09
1:
0>
0C
#148970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#148980000000
0!
0*
09
0>
0C
#148990000000
1!
1*
b1 6
19
1>
1C
b1 G
#149000000000
0!
0*
09
0>
0C
#149010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#149020000000
0!
0*
09
0>
0C
#149030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#149040000000
0!
0*
09
0>
0C
#149050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#149060000000
0!
0*
09
0>
0C
#149070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#149080000000
0!
0#
0*
0,
09
0>
0?
0C
#149090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#149100000000
0!
0*
09
0>
0C
#149110000000
1!
1*
19
1>
1C
#149120000000
0!
0*
09
0>
0C
#149130000000
1!
1*
19
1>
1C
#149140000000
0!
0*
09
0>
0C
#149150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#149160000000
0!
0*
09
0>
0C
#149170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#149180000000
0!
0*
09
0>
0C
#149190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#149200000000
0!
0*
09
0>
0C
#149210000000
1!
1*
b10 6
19
1>
1C
b10 G
#149220000000
0!
0*
09
0>
0C
#149230000000
1!
1*
b11 6
19
1>
1C
b11 G
#149240000000
0!
0*
09
0>
0C
#149250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#149260000000
0!
0*
09
0>
0C
#149270000000
1!
1*
b101 6
19
1>
1C
b101 G
#149280000000
0!
0*
09
0>
0C
#149290000000
1!
1*
b110 6
19
1>
1C
b110 G
#149300000000
0!
0*
09
0>
0C
#149310000000
1!
1*
b111 6
19
1>
1C
b111 G
#149320000000
0!
0*
09
0>
0C
#149330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#149340000000
0!
0*
09
0>
0C
#149350000000
1!
1*
b1 6
19
1>
1C
b1 G
#149360000000
0!
0*
09
0>
0C
#149370000000
1!
1*
b10 6
19
1>
1C
b10 G
#149380000000
0!
0*
09
0>
0C
#149390000000
1!
1*
b11 6
19
1>
1C
b11 G
#149400000000
0!
0*
09
0>
0C
#149410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#149420000000
0!
0*
09
0>
0C
#149430000000
1!
1*
b101 6
19
1>
1C
b101 G
#149440000000
0!
0*
09
0>
0C
#149450000000
1!
1*
b110 6
19
1>
1C
b110 G
#149460000000
0!
0*
09
0>
0C
#149470000000
1!
1*
b111 6
19
1>
1C
b111 G
#149480000000
0!
0*
09
0>
0C
#149490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#149500000000
0!
0*
09
0>
0C
#149510000000
1!
1*
b1 6
19
1>
1C
b1 G
#149520000000
0!
0*
09
0>
0C
#149530000000
1!
1*
b10 6
19
1>
1C
b10 G
#149540000000
0!
0*
09
0>
0C
#149550000000
1!
1*
b11 6
19
1>
1C
b11 G
#149560000000
0!
0*
09
0>
0C
#149570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#149580000000
0!
0*
09
0>
0C
#149590000000
1!
1*
b101 6
19
1>
1C
b101 G
#149600000000
0!
0*
09
0>
0C
#149610000000
1!
1*
b110 6
19
1>
1C
b110 G
#149620000000
0!
0*
09
0>
0C
#149630000000
1!
1*
b111 6
19
1>
1C
b111 G
#149640000000
0!
1"
0*
1+
09
1:
0>
0C
#149650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#149660000000
0!
0*
09
0>
0C
#149670000000
1!
1*
b1 6
19
1>
1C
b1 G
#149680000000
0!
0*
09
0>
0C
#149690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#149700000000
0!
0*
09
0>
0C
#149710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#149720000000
0!
0*
09
0>
0C
#149730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#149740000000
0!
0*
09
0>
0C
#149750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#149760000000
0!
0#
0*
0,
09
0>
0?
0C
#149770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#149780000000
0!
0*
09
0>
0C
#149790000000
1!
1*
19
1>
1C
#149800000000
0!
0*
09
0>
0C
#149810000000
1!
1*
19
1>
1C
#149820000000
0!
0*
09
0>
0C
#149830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#149840000000
0!
0*
09
0>
0C
#149850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#149860000000
0!
0*
09
0>
0C
#149870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#149880000000
0!
0*
09
0>
0C
#149890000000
1!
1*
b10 6
19
1>
1C
b10 G
#149900000000
0!
0*
09
0>
0C
#149910000000
1!
1*
b11 6
19
1>
1C
b11 G
#149920000000
0!
0*
09
0>
0C
#149930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#149940000000
0!
0*
09
0>
0C
#149950000000
1!
1*
b101 6
19
1>
1C
b101 G
#149960000000
0!
0*
09
0>
0C
#149970000000
1!
1*
b110 6
19
1>
1C
b110 G
#149980000000
0!
0*
09
0>
0C
#149990000000
1!
1*
b111 6
19
1>
1C
b111 G
#150000000000
0!
0*
09
0>
0C
#150010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#150020000000
0!
0*
09
0>
0C
#150030000000
1!
1*
b1 6
19
1>
1C
b1 G
#150040000000
0!
0*
09
0>
0C
#150050000000
1!
1*
b10 6
19
1>
1C
b10 G
#150060000000
0!
0*
09
0>
0C
#150070000000
1!
1*
b11 6
19
1>
1C
b11 G
#150080000000
0!
0*
09
0>
0C
#150090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#150100000000
0!
0*
09
0>
0C
#150110000000
1!
1*
b101 6
19
1>
1C
b101 G
#150120000000
0!
0*
09
0>
0C
#150130000000
1!
1*
b110 6
19
1>
1C
b110 G
#150140000000
0!
0*
09
0>
0C
#150150000000
1!
1*
b111 6
19
1>
1C
b111 G
#150160000000
0!
0*
09
0>
0C
#150170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#150180000000
0!
0*
09
0>
0C
#150190000000
1!
1*
b1 6
19
1>
1C
b1 G
#150200000000
0!
0*
09
0>
0C
#150210000000
1!
1*
b10 6
19
1>
1C
b10 G
#150220000000
0!
0*
09
0>
0C
#150230000000
1!
1*
b11 6
19
1>
1C
b11 G
#150240000000
0!
0*
09
0>
0C
#150250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#150260000000
0!
0*
09
0>
0C
#150270000000
1!
1*
b101 6
19
1>
1C
b101 G
#150280000000
0!
0*
09
0>
0C
#150290000000
1!
1*
b110 6
19
1>
1C
b110 G
#150300000000
0!
0*
09
0>
0C
#150310000000
1!
1*
b111 6
19
1>
1C
b111 G
#150320000000
0!
1"
0*
1+
09
1:
0>
0C
#150330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#150340000000
0!
0*
09
0>
0C
#150350000000
1!
1*
b1 6
19
1>
1C
b1 G
#150360000000
0!
0*
09
0>
0C
#150370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#150380000000
0!
0*
09
0>
0C
#150390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#150400000000
0!
0*
09
0>
0C
#150410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#150420000000
0!
0*
09
0>
0C
#150430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#150440000000
0!
0#
0*
0,
09
0>
0?
0C
#150450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#150460000000
0!
0*
09
0>
0C
#150470000000
1!
1*
19
1>
1C
#150480000000
0!
0*
09
0>
0C
#150490000000
1!
1*
19
1>
1C
#150500000000
0!
0*
09
0>
0C
#150510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#150520000000
0!
0*
09
0>
0C
#150530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#150540000000
0!
0*
09
0>
0C
#150550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#150560000000
0!
0*
09
0>
0C
#150570000000
1!
1*
b10 6
19
1>
1C
b10 G
#150580000000
0!
0*
09
0>
0C
#150590000000
1!
1*
b11 6
19
1>
1C
b11 G
#150600000000
0!
0*
09
0>
0C
#150610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#150620000000
0!
0*
09
0>
0C
#150630000000
1!
1*
b101 6
19
1>
1C
b101 G
#150640000000
0!
0*
09
0>
0C
#150650000000
1!
1*
b110 6
19
1>
1C
b110 G
#150660000000
0!
0*
09
0>
0C
#150670000000
1!
1*
b111 6
19
1>
1C
b111 G
#150680000000
0!
0*
09
0>
0C
#150690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#150700000000
0!
0*
09
0>
0C
#150710000000
1!
1*
b1 6
19
1>
1C
b1 G
#150720000000
0!
0*
09
0>
0C
#150730000000
1!
1*
b10 6
19
1>
1C
b10 G
#150740000000
0!
0*
09
0>
0C
#150750000000
1!
1*
b11 6
19
1>
1C
b11 G
#150760000000
0!
0*
09
0>
0C
#150770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#150780000000
0!
0*
09
0>
0C
#150790000000
1!
1*
b101 6
19
1>
1C
b101 G
#150800000000
0!
0*
09
0>
0C
#150810000000
1!
1*
b110 6
19
1>
1C
b110 G
#150820000000
0!
0*
09
0>
0C
#150830000000
1!
1*
b111 6
19
1>
1C
b111 G
#150840000000
0!
0*
09
0>
0C
#150850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#150860000000
0!
0*
09
0>
0C
#150870000000
1!
1*
b1 6
19
1>
1C
b1 G
#150880000000
0!
0*
09
0>
0C
#150890000000
1!
1*
b10 6
19
1>
1C
b10 G
#150900000000
0!
0*
09
0>
0C
#150910000000
1!
1*
b11 6
19
1>
1C
b11 G
#150920000000
0!
0*
09
0>
0C
#150930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#150940000000
0!
0*
09
0>
0C
#150950000000
1!
1*
b101 6
19
1>
1C
b101 G
#150960000000
0!
0*
09
0>
0C
#150970000000
1!
1*
b110 6
19
1>
1C
b110 G
#150980000000
0!
0*
09
0>
0C
#150990000000
1!
1*
b111 6
19
1>
1C
b111 G
#151000000000
0!
1"
0*
1+
09
1:
0>
0C
#151010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#151020000000
0!
0*
09
0>
0C
#151030000000
1!
1*
b1 6
19
1>
1C
b1 G
#151040000000
0!
0*
09
0>
0C
#151050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#151060000000
0!
0*
09
0>
0C
#151070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#151080000000
0!
0*
09
0>
0C
#151090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#151100000000
0!
0*
09
0>
0C
#151110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#151120000000
0!
0#
0*
0,
09
0>
0?
0C
#151130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#151140000000
0!
0*
09
0>
0C
#151150000000
1!
1*
19
1>
1C
#151160000000
0!
0*
09
0>
0C
#151170000000
1!
1*
19
1>
1C
#151180000000
0!
0*
09
0>
0C
#151190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#151200000000
0!
0*
09
0>
0C
#151210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#151220000000
0!
0*
09
0>
0C
#151230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#151240000000
0!
0*
09
0>
0C
#151250000000
1!
1*
b10 6
19
1>
1C
b10 G
#151260000000
0!
0*
09
0>
0C
#151270000000
1!
1*
b11 6
19
1>
1C
b11 G
#151280000000
0!
0*
09
0>
0C
#151290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#151300000000
0!
0*
09
0>
0C
#151310000000
1!
1*
b101 6
19
1>
1C
b101 G
#151320000000
0!
0*
09
0>
0C
#151330000000
1!
1*
b110 6
19
1>
1C
b110 G
#151340000000
0!
0*
09
0>
0C
#151350000000
1!
1*
b111 6
19
1>
1C
b111 G
#151360000000
0!
0*
09
0>
0C
#151370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#151380000000
0!
0*
09
0>
0C
#151390000000
1!
1*
b1 6
19
1>
1C
b1 G
#151400000000
0!
0*
09
0>
0C
#151410000000
1!
1*
b10 6
19
1>
1C
b10 G
#151420000000
0!
0*
09
0>
0C
#151430000000
1!
1*
b11 6
19
1>
1C
b11 G
#151440000000
0!
0*
09
0>
0C
#151450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#151460000000
0!
0*
09
0>
0C
#151470000000
1!
1*
b101 6
19
1>
1C
b101 G
#151480000000
0!
0*
09
0>
0C
#151490000000
1!
1*
b110 6
19
1>
1C
b110 G
#151500000000
0!
0*
09
0>
0C
#151510000000
1!
1*
b111 6
19
1>
1C
b111 G
#151520000000
0!
0*
09
0>
0C
#151530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#151540000000
0!
0*
09
0>
0C
#151550000000
1!
1*
b1 6
19
1>
1C
b1 G
#151560000000
0!
0*
09
0>
0C
#151570000000
1!
1*
b10 6
19
1>
1C
b10 G
#151580000000
0!
0*
09
0>
0C
#151590000000
1!
1*
b11 6
19
1>
1C
b11 G
#151600000000
0!
0*
09
0>
0C
#151610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#151620000000
0!
0*
09
0>
0C
#151630000000
1!
1*
b101 6
19
1>
1C
b101 G
#151640000000
0!
0*
09
0>
0C
#151650000000
1!
1*
b110 6
19
1>
1C
b110 G
#151660000000
0!
0*
09
0>
0C
#151670000000
1!
1*
b111 6
19
1>
1C
b111 G
#151680000000
0!
1"
0*
1+
09
1:
0>
0C
#151690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#151700000000
0!
0*
09
0>
0C
#151710000000
1!
1*
b1 6
19
1>
1C
b1 G
#151720000000
0!
0*
09
0>
0C
#151730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#151740000000
0!
0*
09
0>
0C
#151750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#151760000000
0!
0*
09
0>
0C
#151770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#151780000000
0!
0*
09
0>
0C
#151790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#151800000000
0!
0#
0*
0,
09
0>
0?
0C
#151810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#151820000000
0!
0*
09
0>
0C
#151830000000
1!
1*
19
1>
1C
#151840000000
0!
0*
09
0>
0C
#151850000000
1!
1*
19
1>
1C
#151860000000
0!
0*
09
0>
0C
#151870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#151880000000
0!
0*
09
0>
0C
#151890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#151900000000
0!
0*
09
0>
0C
#151910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#151920000000
0!
0*
09
0>
0C
#151930000000
1!
1*
b10 6
19
1>
1C
b10 G
#151940000000
0!
0*
09
0>
0C
#151950000000
1!
1*
b11 6
19
1>
1C
b11 G
#151960000000
0!
0*
09
0>
0C
#151970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#151980000000
0!
0*
09
0>
0C
#151990000000
1!
1*
b101 6
19
1>
1C
b101 G
#152000000000
0!
0*
09
0>
0C
#152010000000
1!
1*
b110 6
19
1>
1C
b110 G
#152020000000
0!
0*
09
0>
0C
#152030000000
1!
1*
b111 6
19
1>
1C
b111 G
#152040000000
0!
0*
09
0>
0C
#152050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#152060000000
0!
0*
09
0>
0C
#152070000000
1!
1*
b1 6
19
1>
1C
b1 G
#152080000000
0!
0*
09
0>
0C
#152090000000
1!
1*
b10 6
19
1>
1C
b10 G
#152100000000
0!
0*
09
0>
0C
#152110000000
1!
1*
b11 6
19
1>
1C
b11 G
#152120000000
0!
0*
09
0>
0C
#152130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#152140000000
0!
0*
09
0>
0C
#152150000000
1!
1*
b101 6
19
1>
1C
b101 G
#152160000000
0!
0*
09
0>
0C
#152170000000
1!
1*
b110 6
19
1>
1C
b110 G
#152180000000
0!
0*
09
0>
0C
#152190000000
1!
1*
b111 6
19
1>
1C
b111 G
#152200000000
0!
0*
09
0>
0C
#152210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#152220000000
0!
0*
09
0>
0C
#152230000000
1!
1*
b1 6
19
1>
1C
b1 G
#152240000000
0!
0*
09
0>
0C
#152250000000
1!
1*
b10 6
19
1>
1C
b10 G
#152260000000
0!
0*
09
0>
0C
#152270000000
1!
1*
b11 6
19
1>
1C
b11 G
#152280000000
0!
0*
09
0>
0C
#152290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#152300000000
0!
0*
09
0>
0C
#152310000000
1!
1*
b101 6
19
1>
1C
b101 G
#152320000000
0!
0*
09
0>
0C
#152330000000
1!
1*
b110 6
19
1>
1C
b110 G
#152340000000
0!
0*
09
0>
0C
#152350000000
1!
1*
b111 6
19
1>
1C
b111 G
#152360000000
0!
1"
0*
1+
09
1:
0>
0C
#152370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#152380000000
0!
0*
09
0>
0C
#152390000000
1!
1*
b1 6
19
1>
1C
b1 G
#152400000000
0!
0*
09
0>
0C
#152410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#152420000000
0!
0*
09
0>
0C
#152430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#152440000000
0!
0*
09
0>
0C
#152450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#152460000000
0!
0*
09
0>
0C
#152470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#152480000000
0!
0#
0*
0,
09
0>
0?
0C
#152490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#152500000000
0!
0*
09
0>
0C
#152510000000
1!
1*
19
1>
1C
#152520000000
0!
0*
09
0>
0C
#152530000000
1!
1*
19
1>
1C
#152540000000
0!
0*
09
0>
0C
#152550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#152560000000
0!
0*
09
0>
0C
#152570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#152580000000
0!
0*
09
0>
0C
#152590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#152600000000
0!
0*
09
0>
0C
#152610000000
1!
1*
b10 6
19
1>
1C
b10 G
#152620000000
0!
0*
09
0>
0C
#152630000000
1!
1*
b11 6
19
1>
1C
b11 G
#152640000000
0!
0*
09
0>
0C
#152650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#152660000000
0!
0*
09
0>
0C
#152670000000
1!
1*
b101 6
19
1>
1C
b101 G
#152680000000
0!
0*
09
0>
0C
#152690000000
1!
1*
b110 6
19
1>
1C
b110 G
#152700000000
0!
0*
09
0>
0C
#152710000000
1!
1*
b111 6
19
1>
1C
b111 G
#152720000000
0!
0*
09
0>
0C
#152730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#152740000000
0!
0*
09
0>
0C
#152750000000
1!
1*
b1 6
19
1>
1C
b1 G
#152760000000
0!
0*
09
0>
0C
#152770000000
1!
1*
b10 6
19
1>
1C
b10 G
#152780000000
0!
0*
09
0>
0C
#152790000000
1!
1*
b11 6
19
1>
1C
b11 G
#152800000000
0!
0*
09
0>
0C
#152810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#152820000000
0!
0*
09
0>
0C
#152830000000
1!
1*
b101 6
19
1>
1C
b101 G
#152840000000
0!
0*
09
0>
0C
#152850000000
1!
1*
b110 6
19
1>
1C
b110 G
#152860000000
0!
0*
09
0>
0C
#152870000000
1!
1*
b111 6
19
1>
1C
b111 G
#152880000000
0!
0*
09
0>
0C
#152890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#152900000000
0!
0*
09
0>
0C
#152910000000
1!
1*
b1 6
19
1>
1C
b1 G
#152920000000
0!
0*
09
0>
0C
#152930000000
1!
1*
b10 6
19
1>
1C
b10 G
#152940000000
0!
0*
09
0>
0C
#152950000000
1!
1*
b11 6
19
1>
1C
b11 G
#152960000000
0!
0*
09
0>
0C
#152970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#152980000000
0!
0*
09
0>
0C
#152990000000
1!
1*
b101 6
19
1>
1C
b101 G
#153000000000
0!
0*
09
0>
0C
#153010000000
1!
1*
b110 6
19
1>
1C
b110 G
#153020000000
0!
0*
09
0>
0C
#153030000000
1!
1*
b111 6
19
1>
1C
b111 G
#153040000000
0!
1"
0*
1+
09
1:
0>
0C
#153050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#153060000000
0!
0*
09
0>
0C
#153070000000
1!
1*
b1 6
19
1>
1C
b1 G
#153080000000
0!
0*
09
0>
0C
#153090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#153100000000
0!
0*
09
0>
0C
#153110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#153120000000
0!
0*
09
0>
0C
#153130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#153140000000
0!
0*
09
0>
0C
#153150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#153160000000
0!
0#
0*
0,
09
0>
0?
0C
#153170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#153180000000
0!
0*
09
0>
0C
#153190000000
1!
1*
19
1>
1C
#153200000000
0!
0*
09
0>
0C
#153210000000
1!
1*
19
1>
1C
#153220000000
0!
0*
09
0>
0C
#153230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#153240000000
0!
0*
09
0>
0C
#153250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#153260000000
0!
0*
09
0>
0C
#153270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#153280000000
0!
0*
09
0>
0C
#153290000000
1!
1*
b10 6
19
1>
1C
b10 G
#153300000000
0!
0*
09
0>
0C
#153310000000
1!
1*
b11 6
19
1>
1C
b11 G
#153320000000
0!
0*
09
0>
0C
#153330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#153340000000
0!
0*
09
0>
0C
#153350000000
1!
1*
b101 6
19
1>
1C
b101 G
#153360000000
0!
0*
09
0>
0C
#153370000000
1!
1*
b110 6
19
1>
1C
b110 G
#153380000000
0!
0*
09
0>
0C
#153390000000
1!
1*
b111 6
19
1>
1C
b111 G
#153400000000
0!
0*
09
0>
0C
#153410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#153420000000
0!
0*
09
0>
0C
#153430000000
1!
1*
b1 6
19
1>
1C
b1 G
#153440000000
0!
0*
09
0>
0C
#153450000000
1!
1*
b10 6
19
1>
1C
b10 G
#153460000000
0!
0*
09
0>
0C
#153470000000
1!
1*
b11 6
19
1>
1C
b11 G
#153480000000
0!
0*
09
0>
0C
#153490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#153500000000
0!
0*
09
0>
0C
#153510000000
1!
1*
b101 6
19
1>
1C
b101 G
#153520000000
0!
0*
09
0>
0C
#153530000000
1!
1*
b110 6
19
1>
1C
b110 G
#153540000000
0!
0*
09
0>
0C
#153550000000
1!
1*
b111 6
19
1>
1C
b111 G
#153560000000
0!
0*
09
0>
0C
#153570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#153580000000
0!
0*
09
0>
0C
#153590000000
1!
1*
b1 6
19
1>
1C
b1 G
#153600000000
0!
0*
09
0>
0C
#153610000000
1!
1*
b10 6
19
1>
1C
b10 G
#153620000000
0!
0*
09
0>
0C
#153630000000
1!
1*
b11 6
19
1>
1C
b11 G
#153640000000
0!
0*
09
0>
0C
#153650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#153660000000
0!
0*
09
0>
0C
#153670000000
1!
1*
b101 6
19
1>
1C
b101 G
#153680000000
0!
0*
09
0>
0C
#153690000000
1!
1*
b110 6
19
1>
1C
b110 G
#153700000000
0!
0*
09
0>
0C
#153710000000
1!
1*
b111 6
19
1>
1C
b111 G
#153720000000
0!
1"
0*
1+
09
1:
0>
0C
#153730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#153740000000
0!
0*
09
0>
0C
#153750000000
1!
1*
b1 6
19
1>
1C
b1 G
#153760000000
0!
0*
09
0>
0C
#153770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#153780000000
0!
0*
09
0>
0C
#153790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#153800000000
0!
0*
09
0>
0C
#153810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#153820000000
0!
0*
09
0>
0C
#153830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#153840000000
0!
0#
0*
0,
09
0>
0?
0C
#153850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#153860000000
0!
0*
09
0>
0C
#153870000000
1!
1*
19
1>
1C
#153880000000
0!
0*
09
0>
0C
#153890000000
1!
1*
19
1>
1C
#153900000000
0!
0*
09
0>
0C
#153910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#153920000000
0!
0*
09
0>
0C
#153930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#153940000000
0!
0*
09
0>
0C
#153950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#153960000000
0!
0*
09
0>
0C
#153970000000
1!
1*
b10 6
19
1>
1C
b10 G
#153980000000
0!
0*
09
0>
0C
#153990000000
1!
1*
b11 6
19
1>
1C
b11 G
#154000000000
0!
0*
09
0>
0C
#154010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#154020000000
0!
0*
09
0>
0C
#154030000000
1!
1*
b101 6
19
1>
1C
b101 G
#154040000000
0!
0*
09
0>
0C
#154050000000
1!
1*
b110 6
19
1>
1C
b110 G
#154060000000
0!
0*
09
0>
0C
#154070000000
1!
1*
b111 6
19
1>
1C
b111 G
#154080000000
0!
0*
09
0>
0C
#154090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#154100000000
0!
0*
09
0>
0C
#154110000000
1!
1*
b1 6
19
1>
1C
b1 G
#154120000000
0!
0*
09
0>
0C
#154130000000
1!
1*
b10 6
19
1>
1C
b10 G
#154140000000
0!
0*
09
0>
0C
#154150000000
1!
1*
b11 6
19
1>
1C
b11 G
#154160000000
0!
0*
09
0>
0C
#154170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#154180000000
0!
0*
09
0>
0C
#154190000000
1!
1*
b101 6
19
1>
1C
b101 G
#154200000000
0!
0*
09
0>
0C
#154210000000
1!
1*
b110 6
19
1>
1C
b110 G
#154220000000
0!
0*
09
0>
0C
#154230000000
1!
1*
b111 6
19
1>
1C
b111 G
#154240000000
0!
0*
09
0>
0C
#154250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#154260000000
0!
0*
09
0>
0C
#154270000000
1!
1*
b1 6
19
1>
1C
b1 G
#154280000000
0!
0*
09
0>
0C
#154290000000
1!
1*
b10 6
19
1>
1C
b10 G
#154300000000
0!
0*
09
0>
0C
#154310000000
1!
1*
b11 6
19
1>
1C
b11 G
#154320000000
0!
0*
09
0>
0C
#154330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#154340000000
0!
0*
09
0>
0C
#154350000000
1!
1*
b101 6
19
1>
1C
b101 G
#154360000000
0!
0*
09
0>
0C
#154370000000
1!
1*
b110 6
19
1>
1C
b110 G
#154380000000
0!
0*
09
0>
0C
#154390000000
1!
1*
b111 6
19
1>
1C
b111 G
#154400000000
0!
1"
0*
1+
09
1:
0>
0C
#154410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#154420000000
0!
0*
09
0>
0C
#154430000000
1!
1*
b1 6
19
1>
1C
b1 G
#154440000000
0!
0*
09
0>
0C
#154450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#154460000000
0!
0*
09
0>
0C
#154470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#154480000000
0!
0*
09
0>
0C
#154490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#154500000000
0!
0*
09
0>
0C
#154510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#154520000000
0!
0#
0*
0,
09
0>
0?
0C
#154530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#154540000000
0!
0*
09
0>
0C
#154550000000
1!
1*
19
1>
1C
#154560000000
0!
0*
09
0>
0C
#154570000000
1!
1*
19
1>
1C
#154580000000
0!
0*
09
0>
0C
#154590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#154600000000
0!
0*
09
0>
0C
#154610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#154620000000
0!
0*
09
0>
0C
#154630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#154640000000
0!
0*
09
0>
0C
#154650000000
1!
1*
b10 6
19
1>
1C
b10 G
#154660000000
0!
0*
09
0>
0C
#154670000000
1!
1*
b11 6
19
1>
1C
b11 G
#154680000000
0!
0*
09
0>
0C
#154690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#154700000000
0!
0*
09
0>
0C
#154710000000
1!
1*
b101 6
19
1>
1C
b101 G
#154720000000
0!
0*
09
0>
0C
#154730000000
1!
1*
b110 6
19
1>
1C
b110 G
#154740000000
0!
0*
09
0>
0C
#154750000000
1!
1*
b111 6
19
1>
1C
b111 G
#154760000000
0!
0*
09
0>
0C
#154770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#154780000000
0!
0*
09
0>
0C
#154790000000
1!
1*
b1 6
19
1>
1C
b1 G
#154800000000
0!
0*
09
0>
0C
#154810000000
1!
1*
b10 6
19
1>
1C
b10 G
#154820000000
0!
0*
09
0>
0C
#154830000000
1!
1*
b11 6
19
1>
1C
b11 G
#154840000000
0!
0*
09
0>
0C
#154850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#154860000000
0!
0*
09
0>
0C
#154870000000
1!
1*
b101 6
19
1>
1C
b101 G
#154880000000
0!
0*
09
0>
0C
#154890000000
1!
1*
b110 6
19
1>
1C
b110 G
#154900000000
0!
0*
09
0>
0C
#154910000000
1!
1*
b111 6
19
1>
1C
b111 G
#154920000000
0!
0*
09
0>
0C
#154930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#154940000000
0!
0*
09
0>
0C
#154950000000
1!
1*
b1 6
19
1>
1C
b1 G
#154960000000
0!
0*
09
0>
0C
#154970000000
1!
1*
b10 6
19
1>
1C
b10 G
#154980000000
0!
0*
09
0>
0C
#154990000000
1!
1*
b11 6
19
1>
1C
b11 G
#155000000000
0!
0*
09
0>
0C
#155010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#155020000000
0!
0*
09
0>
0C
#155030000000
1!
1*
b101 6
19
1>
1C
b101 G
#155040000000
0!
0*
09
0>
0C
#155050000000
1!
1*
b110 6
19
1>
1C
b110 G
#155060000000
0!
0*
09
0>
0C
#155070000000
1!
1*
b111 6
19
1>
1C
b111 G
#155080000000
0!
1"
0*
1+
09
1:
0>
0C
#155090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#155100000000
0!
0*
09
0>
0C
#155110000000
1!
1*
b1 6
19
1>
1C
b1 G
#155120000000
0!
0*
09
0>
0C
#155130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#155140000000
0!
0*
09
0>
0C
#155150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#155160000000
0!
0*
09
0>
0C
#155170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#155180000000
0!
0*
09
0>
0C
#155190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#155200000000
0!
0#
0*
0,
09
0>
0?
0C
#155210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#155220000000
0!
0*
09
0>
0C
#155230000000
1!
1*
19
1>
1C
#155240000000
0!
0*
09
0>
0C
#155250000000
1!
1*
19
1>
1C
#155260000000
0!
0*
09
0>
0C
#155270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#155280000000
0!
0*
09
0>
0C
#155290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#155300000000
0!
0*
09
0>
0C
#155310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#155320000000
0!
0*
09
0>
0C
#155330000000
1!
1*
b10 6
19
1>
1C
b10 G
#155340000000
0!
0*
09
0>
0C
#155350000000
1!
1*
b11 6
19
1>
1C
b11 G
#155360000000
0!
0*
09
0>
0C
#155370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#155380000000
0!
0*
09
0>
0C
#155390000000
1!
1*
b101 6
19
1>
1C
b101 G
#155400000000
0!
0*
09
0>
0C
#155410000000
1!
1*
b110 6
19
1>
1C
b110 G
#155420000000
0!
0*
09
0>
0C
#155430000000
1!
1*
b111 6
19
1>
1C
b111 G
#155440000000
0!
0*
09
0>
0C
#155450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#155460000000
0!
0*
09
0>
0C
#155470000000
1!
1*
b1 6
19
1>
1C
b1 G
#155480000000
0!
0*
09
0>
0C
#155490000000
1!
1*
b10 6
19
1>
1C
b10 G
#155500000000
0!
0*
09
0>
0C
#155510000000
1!
1*
b11 6
19
1>
1C
b11 G
#155520000000
0!
0*
09
0>
0C
#155530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#155540000000
0!
0*
09
0>
0C
#155550000000
1!
1*
b101 6
19
1>
1C
b101 G
#155560000000
0!
0*
09
0>
0C
#155570000000
1!
1*
b110 6
19
1>
1C
b110 G
#155580000000
0!
0*
09
0>
0C
#155590000000
1!
1*
b111 6
19
1>
1C
b111 G
#155600000000
0!
0*
09
0>
0C
#155610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#155620000000
0!
0*
09
0>
0C
#155630000000
1!
1*
b1 6
19
1>
1C
b1 G
#155640000000
0!
0*
09
0>
0C
#155650000000
1!
1*
b10 6
19
1>
1C
b10 G
#155660000000
0!
0*
09
0>
0C
#155670000000
1!
1*
b11 6
19
1>
1C
b11 G
#155680000000
0!
0*
09
0>
0C
#155690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#155700000000
0!
0*
09
0>
0C
#155710000000
1!
1*
b101 6
19
1>
1C
b101 G
#155720000000
0!
0*
09
0>
0C
#155730000000
1!
1*
b110 6
19
1>
1C
b110 G
#155740000000
0!
0*
09
0>
0C
#155750000000
1!
1*
b111 6
19
1>
1C
b111 G
#155760000000
0!
1"
0*
1+
09
1:
0>
0C
#155770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#155780000000
0!
0*
09
0>
0C
#155790000000
1!
1*
b1 6
19
1>
1C
b1 G
#155800000000
0!
0*
09
0>
0C
#155810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#155820000000
0!
0*
09
0>
0C
#155830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#155840000000
0!
0*
09
0>
0C
#155850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#155860000000
0!
0*
09
0>
0C
#155870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#155880000000
0!
0#
0*
0,
09
0>
0?
0C
#155890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#155900000000
0!
0*
09
0>
0C
#155910000000
1!
1*
19
1>
1C
#155920000000
0!
0*
09
0>
0C
#155930000000
1!
1*
19
1>
1C
#155940000000
0!
0*
09
0>
0C
#155950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#155960000000
0!
0*
09
0>
0C
#155970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#155980000000
0!
0*
09
0>
0C
#155990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#156000000000
0!
0*
09
0>
0C
#156010000000
1!
1*
b10 6
19
1>
1C
b10 G
#156020000000
0!
0*
09
0>
0C
#156030000000
1!
1*
b11 6
19
1>
1C
b11 G
#156040000000
0!
0*
09
0>
0C
#156050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#156060000000
0!
0*
09
0>
0C
#156070000000
1!
1*
b101 6
19
1>
1C
b101 G
#156080000000
0!
0*
09
0>
0C
#156090000000
1!
1*
b110 6
19
1>
1C
b110 G
#156100000000
0!
0*
09
0>
0C
#156110000000
1!
1*
b111 6
19
1>
1C
b111 G
#156120000000
0!
0*
09
0>
0C
#156130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#156140000000
0!
0*
09
0>
0C
#156150000000
1!
1*
b1 6
19
1>
1C
b1 G
#156160000000
0!
0*
09
0>
0C
#156170000000
1!
1*
b10 6
19
1>
1C
b10 G
#156180000000
0!
0*
09
0>
0C
#156190000000
1!
1*
b11 6
19
1>
1C
b11 G
#156200000000
0!
0*
09
0>
0C
#156210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#156220000000
0!
0*
09
0>
0C
#156230000000
1!
1*
b101 6
19
1>
1C
b101 G
#156240000000
0!
0*
09
0>
0C
#156250000000
1!
1*
b110 6
19
1>
1C
b110 G
#156260000000
0!
0*
09
0>
0C
#156270000000
1!
1*
b111 6
19
1>
1C
b111 G
#156280000000
0!
0*
09
0>
0C
#156290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#156300000000
0!
0*
09
0>
0C
#156310000000
1!
1*
b1 6
19
1>
1C
b1 G
#156320000000
0!
0*
09
0>
0C
#156330000000
1!
1*
b10 6
19
1>
1C
b10 G
#156340000000
0!
0*
09
0>
0C
#156350000000
1!
1*
b11 6
19
1>
1C
b11 G
#156360000000
0!
0*
09
0>
0C
#156370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#156380000000
0!
0*
09
0>
0C
#156390000000
1!
1*
b101 6
19
1>
1C
b101 G
#156400000000
0!
0*
09
0>
0C
#156410000000
1!
1*
b110 6
19
1>
1C
b110 G
#156420000000
0!
0*
09
0>
0C
#156430000000
1!
1*
b111 6
19
1>
1C
b111 G
#156440000000
0!
1"
0*
1+
09
1:
0>
0C
#156450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#156460000000
0!
0*
09
0>
0C
#156470000000
1!
1*
b1 6
19
1>
1C
b1 G
#156480000000
0!
0*
09
0>
0C
#156490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#156500000000
0!
0*
09
0>
0C
#156510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#156520000000
0!
0*
09
0>
0C
#156530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#156540000000
0!
0*
09
0>
0C
#156550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#156560000000
0!
0#
0*
0,
09
0>
0?
0C
#156570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#156580000000
0!
0*
09
0>
0C
#156590000000
1!
1*
19
1>
1C
#156600000000
0!
0*
09
0>
0C
#156610000000
1!
1*
19
1>
1C
#156620000000
0!
0*
09
0>
0C
#156630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#156640000000
0!
0*
09
0>
0C
#156650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#156660000000
0!
0*
09
0>
0C
#156670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#156680000000
0!
0*
09
0>
0C
#156690000000
1!
1*
b10 6
19
1>
1C
b10 G
#156700000000
0!
0*
09
0>
0C
#156710000000
1!
1*
b11 6
19
1>
1C
b11 G
#156720000000
0!
0*
09
0>
0C
#156730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#156740000000
0!
0*
09
0>
0C
#156750000000
1!
1*
b101 6
19
1>
1C
b101 G
#156760000000
0!
0*
09
0>
0C
#156770000000
1!
1*
b110 6
19
1>
1C
b110 G
#156780000000
0!
0*
09
0>
0C
#156790000000
1!
1*
b111 6
19
1>
1C
b111 G
#156800000000
0!
0*
09
0>
0C
#156810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#156820000000
0!
0*
09
0>
0C
#156830000000
1!
1*
b1 6
19
1>
1C
b1 G
#156840000000
0!
0*
09
0>
0C
#156850000000
1!
1*
b10 6
19
1>
1C
b10 G
#156860000000
0!
0*
09
0>
0C
#156870000000
1!
1*
b11 6
19
1>
1C
b11 G
#156880000000
0!
0*
09
0>
0C
#156890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#156900000000
0!
0*
09
0>
0C
#156910000000
1!
1*
b101 6
19
1>
1C
b101 G
#156920000000
0!
0*
09
0>
0C
#156930000000
1!
1*
b110 6
19
1>
1C
b110 G
#156940000000
0!
0*
09
0>
0C
#156950000000
1!
1*
b111 6
19
1>
1C
b111 G
#156960000000
0!
0*
09
0>
0C
#156970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#156980000000
0!
0*
09
0>
0C
#156990000000
1!
1*
b1 6
19
1>
1C
b1 G
#157000000000
0!
0*
09
0>
0C
#157010000000
1!
1*
b10 6
19
1>
1C
b10 G
#157020000000
0!
0*
09
0>
0C
#157030000000
1!
1*
b11 6
19
1>
1C
b11 G
#157040000000
0!
0*
09
0>
0C
#157050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#157060000000
0!
0*
09
0>
0C
#157070000000
1!
1*
b101 6
19
1>
1C
b101 G
#157080000000
0!
0*
09
0>
0C
#157090000000
1!
1*
b110 6
19
1>
1C
b110 G
#157100000000
0!
0*
09
0>
0C
#157110000000
1!
1*
b111 6
19
1>
1C
b111 G
#157120000000
0!
1"
0*
1+
09
1:
0>
0C
#157130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#157140000000
0!
0*
09
0>
0C
#157150000000
1!
1*
b1 6
19
1>
1C
b1 G
#157160000000
0!
0*
09
0>
0C
#157170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#157180000000
0!
0*
09
0>
0C
#157190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#157200000000
0!
0*
09
0>
0C
#157210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#157220000000
0!
0*
09
0>
0C
#157230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#157240000000
0!
0#
0*
0,
09
0>
0?
0C
#157250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#157260000000
0!
0*
09
0>
0C
#157270000000
1!
1*
19
1>
1C
#157280000000
0!
0*
09
0>
0C
#157290000000
1!
1*
19
1>
1C
#157300000000
0!
0*
09
0>
0C
#157310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#157320000000
0!
0*
09
0>
0C
#157330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#157340000000
0!
0*
09
0>
0C
#157350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#157360000000
0!
0*
09
0>
0C
#157370000000
1!
1*
b10 6
19
1>
1C
b10 G
#157380000000
0!
0*
09
0>
0C
#157390000000
1!
1*
b11 6
19
1>
1C
b11 G
#157400000000
0!
0*
09
0>
0C
#157410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#157420000000
0!
0*
09
0>
0C
#157430000000
1!
1*
b101 6
19
1>
1C
b101 G
#157440000000
0!
0*
09
0>
0C
#157450000000
1!
1*
b110 6
19
1>
1C
b110 G
#157460000000
0!
0*
09
0>
0C
#157470000000
1!
1*
b111 6
19
1>
1C
b111 G
#157480000000
0!
0*
09
0>
0C
#157490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#157500000000
0!
0*
09
0>
0C
#157510000000
1!
1*
b1 6
19
1>
1C
b1 G
#157520000000
0!
0*
09
0>
0C
#157530000000
1!
1*
b10 6
19
1>
1C
b10 G
#157540000000
0!
0*
09
0>
0C
#157550000000
1!
1*
b11 6
19
1>
1C
b11 G
#157560000000
0!
0*
09
0>
0C
#157570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#157580000000
0!
0*
09
0>
0C
#157590000000
1!
1*
b101 6
19
1>
1C
b101 G
#157600000000
0!
0*
09
0>
0C
#157610000000
1!
1*
b110 6
19
1>
1C
b110 G
#157620000000
0!
0*
09
0>
0C
#157630000000
1!
1*
b111 6
19
1>
1C
b111 G
#157640000000
0!
0*
09
0>
0C
#157650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#157660000000
0!
0*
09
0>
0C
#157670000000
1!
1*
b1 6
19
1>
1C
b1 G
#157680000000
0!
0*
09
0>
0C
#157690000000
1!
1*
b10 6
19
1>
1C
b10 G
#157700000000
0!
0*
09
0>
0C
#157710000000
1!
1*
b11 6
19
1>
1C
b11 G
#157720000000
0!
0*
09
0>
0C
#157730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#157740000000
0!
0*
09
0>
0C
#157750000000
1!
1*
b101 6
19
1>
1C
b101 G
#157760000000
0!
0*
09
0>
0C
#157770000000
1!
1*
b110 6
19
1>
1C
b110 G
#157780000000
0!
0*
09
0>
0C
#157790000000
1!
1*
b111 6
19
1>
1C
b111 G
#157800000000
0!
1"
0*
1+
09
1:
0>
0C
#157810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#157820000000
0!
0*
09
0>
0C
#157830000000
1!
1*
b1 6
19
1>
1C
b1 G
#157840000000
0!
0*
09
0>
0C
#157850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#157860000000
0!
0*
09
0>
0C
#157870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#157880000000
0!
0*
09
0>
0C
#157890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#157900000000
0!
0*
09
0>
0C
#157910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#157920000000
0!
0#
0*
0,
09
0>
0?
0C
#157930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#157940000000
0!
0*
09
0>
0C
#157950000000
1!
1*
19
1>
1C
#157960000000
0!
0*
09
0>
0C
#157970000000
1!
1*
19
1>
1C
#157980000000
0!
0*
09
0>
0C
#157990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#158000000000
0!
0*
09
0>
0C
#158010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#158020000000
0!
0*
09
0>
0C
#158030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#158040000000
0!
0*
09
0>
0C
#158050000000
1!
1*
b10 6
19
1>
1C
b10 G
#158060000000
0!
0*
09
0>
0C
#158070000000
1!
1*
b11 6
19
1>
1C
b11 G
#158080000000
0!
0*
09
0>
0C
#158090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#158100000000
0!
0*
09
0>
0C
#158110000000
1!
1*
b101 6
19
1>
1C
b101 G
#158120000000
0!
0*
09
0>
0C
#158130000000
1!
1*
b110 6
19
1>
1C
b110 G
#158140000000
0!
0*
09
0>
0C
#158150000000
1!
1*
b111 6
19
1>
1C
b111 G
#158160000000
0!
0*
09
0>
0C
#158170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#158180000000
0!
0*
09
0>
0C
#158190000000
1!
1*
b1 6
19
1>
1C
b1 G
#158200000000
0!
0*
09
0>
0C
#158210000000
1!
1*
b10 6
19
1>
1C
b10 G
#158220000000
0!
0*
09
0>
0C
#158230000000
1!
1*
b11 6
19
1>
1C
b11 G
#158240000000
0!
0*
09
0>
0C
#158250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#158260000000
0!
0*
09
0>
0C
#158270000000
1!
1*
b101 6
19
1>
1C
b101 G
#158280000000
0!
0*
09
0>
0C
#158290000000
1!
1*
b110 6
19
1>
1C
b110 G
#158300000000
0!
0*
09
0>
0C
#158310000000
1!
1*
b111 6
19
1>
1C
b111 G
#158320000000
0!
0*
09
0>
0C
#158330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#158340000000
0!
0*
09
0>
0C
#158350000000
1!
1*
b1 6
19
1>
1C
b1 G
#158360000000
0!
0*
09
0>
0C
#158370000000
1!
1*
b10 6
19
1>
1C
b10 G
#158380000000
0!
0*
09
0>
0C
#158390000000
1!
1*
b11 6
19
1>
1C
b11 G
#158400000000
0!
0*
09
0>
0C
#158410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#158420000000
0!
0*
09
0>
0C
#158430000000
1!
1*
b101 6
19
1>
1C
b101 G
#158440000000
0!
0*
09
0>
0C
#158450000000
1!
1*
b110 6
19
1>
1C
b110 G
#158460000000
0!
0*
09
0>
0C
#158470000000
1!
1*
b111 6
19
1>
1C
b111 G
#158480000000
0!
1"
0*
1+
09
1:
0>
0C
#158490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#158500000000
0!
0*
09
0>
0C
#158510000000
1!
1*
b1 6
19
1>
1C
b1 G
#158520000000
0!
0*
09
0>
0C
#158530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#158540000000
0!
0*
09
0>
0C
#158550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#158560000000
0!
0*
09
0>
0C
#158570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#158580000000
0!
0*
09
0>
0C
#158590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#158600000000
0!
0#
0*
0,
09
0>
0?
0C
#158610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#158620000000
0!
0*
09
0>
0C
#158630000000
1!
1*
19
1>
1C
#158640000000
0!
0*
09
0>
0C
#158650000000
1!
1*
19
1>
1C
#158660000000
0!
0*
09
0>
0C
#158670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#158680000000
0!
0*
09
0>
0C
#158690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#158700000000
0!
0*
09
0>
0C
#158710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#158720000000
0!
0*
09
0>
0C
#158730000000
1!
1*
b10 6
19
1>
1C
b10 G
#158740000000
0!
0*
09
0>
0C
#158750000000
1!
1*
b11 6
19
1>
1C
b11 G
#158760000000
0!
0*
09
0>
0C
#158770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#158780000000
0!
0*
09
0>
0C
#158790000000
1!
1*
b101 6
19
1>
1C
b101 G
#158800000000
0!
0*
09
0>
0C
#158810000000
1!
1*
b110 6
19
1>
1C
b110 G
#158820000000
0!
0*
09
0>
0C
#158830000000
1!
1*
b111 6
19
1>
1C
b111 G
#158840000000
0!
0*
09
0>
0C
#158850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#158860000000
0!
0*
09
0>
0C
#158870000000
1!
1*
b1 6
19
1>
1C
b1 G
#158880000000
0!
0*
09
0>
0C
#158890000000
1!
1*
b10 6
19
1>
1C
b10 G
#158900000000
0!
0*
09
0>
0C
#158910000000
1!
1*
b11 6
19
1>
1C
b11 G
#158920000000
0!
0*
09
0>
0C
#158930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#158940000000
0!
0*
09
0>
0C
#158950000000
1!
1*
b101 6
19
1>
1C
b101 G
#158960000000
0!
0*
09
0>
0C
#158970000000
1!
1*
b110 6
19
1>
1C
b110 G
#158980000000
0!
0*
09
0>
0C
#158990000000
1!
1*
b111 6
19
1>
1C
b111 G
#159000000000
0!
0*
09
0>
0C
#159010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#159020000000
0!
0*
09
0>
0C
#159030000000
1!
1*
b1 6
19
1>
1C
b1 G
#159040000000
0!
0*
09
0>
0C
#159050000000
1!
1*
b10 6
19
1>
1C
b10 G
#159060000000
0!
0*
09
0>
0C
#159070000000
1!
1*
b11 6
19
1>
1C
b11 G
#159080000000
0!
0*
09
0>
0C
#159090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#159100000000
0!
0*
09
0>
0C
#159110000000
1!
1*
b101 6
19
1>
1C
b101 G
#159120000000
0!
0*
09
0>
0C
#159130000000
1!
1*
b110 6
19
1>
1C
b110 G
#159140000000
0!
0*
09
0>
0C
#159150000000
1!
1*
b111 6
19
1>
1C
b111 G
#159160000000
0!
1"
0*
1+
09
1:
0>
0C
#159170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#159180000000
0!
0*
09
0>
0C
#159190000000
1!
1*
b1 6
19
1>
1C
b1 G
#159200000000
0!
0*
09
0>
0C
#159210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#159220000000
0!
0*
09
0>
0C
#159230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#159240000000
0!
0*
09
0>
0C
#159250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#159260000000
0!
0*
09
0>
0C
#159270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#159280000000
0!
0#
0*
0,
09
0>
0?
0C
#159290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#159300000000
0!
0*
09
0>
0C
#159310000000
1!
1*
19
1>
1C
#159320000000
0!
0*
09
0>
0C
#159330000000
1!
1*
19
1>
1C
#159340000000
0!
0*
09
0>
0C
#159350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#159360000000
0!
0*
09
0>
0C
#159370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#159380000000
0!
0*
09
0>
0C
#159390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#159400000000
0!
0*
09
0>
0C
#159410000000
1!
1*
b10 6
19
1>
1C
b10 G
#159420000000
0!
0*
09
0>
0C
#159430000000
1!
1*
b11 6
19
1>
1C
b11 G
#159440000000
0!
0*
09
0>
0C
#159450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#159460000000
0!
0*
09
0>
0C
#159470000000
1!
1*
b101 6
19
1>
1C
b101 G
#159480000000
0!
0*
09
0>
0C
#159490000000
1!
1*
b110 6
19
1>
1C
b110 G
#159500000000
0!
0*
09
0>
0C
#159510000000
1!
1*
b111 6
19
1>
1C
b111 G
#159520000000
0!
0*
09
0>
0C
#159530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#159540000000
0!
0*
09
0>
0C
#159550000000
1!
1*
b1 6
19
1>
1C
b1 G
#159560000000
0!
0*
09
0>
0C
#159570000000
1!
1*
b10 6
19
1>
1C
b10 G
#159580000000
0!
0*
09
0>
0C
#159590000000
1!
1*
b11 6
19
1>
1C
b11 G
#159600000000
0!
0*
09
0>
0C
#159610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#159620000000
0!
0*
09
0>
0C
#159630000000
1!
1*
b101 6
19
1>
1C
b101 G
#159640000000
0!
0*
09
0>
0C
#159650000000
1!
1*
b110 6
19
1>
1C
b110 G
#159660000000
0!
0*
09
0>
0C
#159670000000
1!
1*
b111 6
19
1>
1C
b111 G
#159680000000
0!
0*
09
0>
0C
#159690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#159700000000
0!
0*
09
0>
0C
#159710000000
1!
1*
b1 6
19
1>
1C
b1 G
#159720000000
0!
0*
09
0>
0C
#159730000000
1!
1*
b10 6
19
1>
1C
b10 G
#159740000000
0!
0*
09
0>
0C
#159750000000
1!
1*
b11 6
19
1>
1C
b11 G
#159760000000
0!
0*
09
0>
0C
#159770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#159780000000
0!
0*
09
0>
0C
#159790000000
1!
1*
b101 6
19
1>
1C
b101 G
#159800000000
0!
0*
09
0>
0C
#159810000000
1!
1*
b110 6
19
1>
1C
b110 G
#159820000000
0!
0*
09
0>
0C
#159830000000
1!
1*
b111 6
19
1>
1C
b111 G
#159840000000
0!
1"
0*
1+
09
1:
0>
0C
#159850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#159860000000
0!
0*
09
0>
0C
#159870000000
1!
1*
b1 6
19
1>
1C
b1 G
#159880000000
0!
0*
09
0>
0C
#159890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#159900000000
0!
0*
09
0>
0C
#159910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#159920000000
0!
0*
09
0>
0C
#159930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#159940000000
0!
0*
09
0>
0C
#159950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#159960000000
0!
0#
0*
0,
09
0>
0?
0C
#159970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#159980000000
0!
0*
09
0>
0C
#159990000000
1!
1*
19
1>
1C
#160000000000
0!
0*
09
0>
0C
#160010000000
1!
1*
19
1>
1C
#160020000000
0!
0*
09
0>
0C
#160030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#160040000000
0!
0*
09
0>
0C
#160050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#160060000000
0!
0*
09
0>
0C
#160070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#160080000000
0!
0*
09
0>
0C
#160090000000
1!
1*
b10 6
19
1>
1C
b10 G
#160100000000
0!
0*
09
0>
0C
#160110000000
1!
1*
b11 6
19
1>
1C
b11 G
#160120000000
0!
0*
09
0>
0C
#160130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#160140000000
0!
0*
09
0>
0C
#160150000000
1!
1*
b101 6
19
1>
1C
b101 G
#160160000000
0!
0*
09
0>
0C
#160170000000
1!
1*
b110 6
19
1>
1C
b110 G
#160180000000
0!
0*
09
0>
0C
#160190000000
1!
1*
b111 6
19
1>
1C
b111 G
#160200000000
0!
0*
09
0>
0C
#160210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#160220000000
0!
0*
09
0>
0C
#160230000000
1!
1*
b1 6
19
1>
1C
b1 G
#160240000000
0!
0*
09
0>
0C
#160250000000
1!
1*
b10 6
19
1>
1C
b10 G
#160260000000
0!
0*
09
0>
0C
#160270000000
1!
1*
b11 6
19
1>
1C
b11 G
#160280000000
0!
0*
09
0>
0C
#160290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#160300000000
0!
0*
09
0>
0C
#160310000000
1!
1*
b101 6
19
1>
1C
b101 G
#160320000000
0!
0*
09
0>
0C
#160330000000
1!
1*
b110 6
19
1>
1C
b110 G
#160340000000
0!
0*
09
0>
0C
#160350000000
1!
1*
b111 6
19
1>
1C
b111 G
#160360000000
0!
0*
09
0>
0C
#160370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#160380000000
0!
0*
09
0>
0C
#160390000000
1!
1*
b1 6
19
1>
1C
b1 G
#160400000000
0!
0*
09
0>
0C
#160410000000
1!
1*
b10 6
19
1>
1C
b10 G
#160420000000
0!
0*
09
0>
0C
#160430000000
1!
1*
b11 6
19
1>
1C
b11 G
#160440000000
0!
0*
09
0>
0C
#160450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#160460000000
0!
0*
09
0>
0C
#160470000000
1!
1*
b101 6
19
1>
1C
b101 G
#160480000000
0!
0*
09
0>
0C
#160490000000
1!
1*
b110 6
19
1>
1C
b110 G
#160500000000
0!
0*
09
0>
0C
#160510000000
1!
1*
b111 6
19
1>
1C
b111 G
#160520000000
0!
1"
0*
1+
09
1:
0>
0C
#160530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#160540000000
0!
0*
09
0>
0C
#160550000000
1!
1*
b1 6
19
1>
1C
b1 G
#160560000000
0!
0*
09
0>
0C
#160570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#160580000000
0!
0*
09
0>
0C
#160590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#160600000000
0!
0*
09
0>
0C
#160610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#160620000000
0!
0*
09
0>
0C
#160630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#160640000000
0!
0#
0*
0,
09
0>
0?
0C
#160650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#160660000000
0!
0*
09
0>
0C
#160670000000
1!
1*
19
1>
1C
#160680000000
0!
0*
09
0>
0C
#160690000000
1!
1*
19
1>
1C
#160700000000
0!
0*
09
0>
0C
#160710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#160720000000
0!
0*
09
0>
0C
#160730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#160740000000
0!
0*
09
0>
0C
#160750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#160760000000
0!
0*
09
0>
0C
#160770000000
1!
1*
b10 6
19
1>
1C
b10 G
#160780000000
0!
0*
09
0>
0C
#160790000000
1!
1*
b11 6
19
1>
1C
b11 G
#160800000000
0!
0*
09
0>
0C
#160810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#160820000000
0!
0*
09
0>
0C
#160830000000
1!
1*
b101 6
19
1>
1C
b101 G
#160840000000
0!
0*
09
0>
0C
#160850000000
1!
1*
b110 6
19
1>
1C
b110 G
#160860000000
0!
0*
09
0>
0C
#160870000000
1!
1*
b111 6
19
1>
1C
b111 G
#160880000000
0!
0*
09
0>
0C
#160890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#160900000000
0!
0*
09
0>
0C
#160910000000
1!
1*
b1 6
19
1>
1C
b1 G
#160920000000
0!
0*
09
0>
0C
#160930000000
1!
1*
b10 6
19
1>
1C
b10 G
#160940000000
0!
0*
09
0>
0C
#160950000000
1!
1*
b11 6
19
1>
1C
b11 G
#160960000000
0!
0*
09
0>
0C
#160970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#160980000000
0!
0*
09
0>
0C
#160990000000
1!
1*
b101 6
19
1>
1C
b101 G
#161000000000
0!
0*
09
0>
0C
#161010000000
1!
1*
b110 6
19
1>
1C
b110 G
#161020000000
0!
0*
09
0>
0C
#161030000000
1!
1*
b111 6
19
1>
1C
b111 G
#161040000000
0!
0*
09
0>
0C
#161050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#161060000000
0!
0*
09
0>
0C
#161070000000
1!
1*
b1 6
19
1>
1C
b1 G
#161080000000
0!
0*
09
0>
0C
#161090000000
1!
1*
b10 6
19
1>
1C
b10 G
#161100000000
0!
0*
09
0>
0C
#161110000000
1!
1*
b11 6
19
1>
1C
b11 G
#161120000000
0!
0*
09
0>
0C
#161130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#161140000000
0!
0*
09
0>
0C
#161150000000
1!
1*
b101 6
19
1>
1C
b101 G
#161160000000
0!
0*
09
0>
0C
#161170000000
1!
1*
b110 6
19
1>
1C
b110 G
#161180000000
0!
0*
09
0>
0C
#161190000000
1!
1*
b111 6
19
1>
1C
b111 G
#161200000000
0!
1"
0*
1+
09
1:
0>
0C
#161210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#161220000000
0!
0*
09
0>
0C
#161230000000
1!
1*
b1 6
19
1>
1C
b1 G
#161240000000
0!
0*
09
0>
0C
#161250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#161260000000
0!
0*
09
0>
0C
#161270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#161280000000
0!
0*
09
0>
0C
#161290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#161300000000
0!
0*
09
0>
0C
#161310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#161320000000
0!
0#
0*
0,
09
0>
0?
0C
#161330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#161340000000
0!
0*
09
0>
0C
#161350000000
1!
1*
19
1>
1C
#161360000000
0!
0*
09
0>
0C
#161370000000
1!
1*
19
1>
1C
#161380000000
0!
0*
09
0>
0C
#161390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#161400000000
0!
0*
09
0>
0C
#161410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#161420000000
0!
0*
09
0>
0C
#161430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#161440000000
0!
0*
09
0>
0C
#161450000000
1!
1*
b10 6
19
1>
1C
b10 G
#161460000000
0!
0*
09
0>
0C
#161470000000
1!
1*
b11 6
19
1>
1C
b11 G
#161480000000
0!
0*
09
0>
0C
#161490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#161500000000
0!
0*
09
0>
0C
#161510000000
1!
1*
b101 6
19
1>
1C
b101 G
#161520000000
0!
0*
09
0>
0C
#161530000000
1!
1*
b110 6
19
1>
1C
b110 G
#161540000000
0!
0*
09
0>
0C
#161550000000
1!
1*
b111 6
19
1>
1C
b111 G
#161560000000
0!
0*
09
0>
0C
#161570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#161580000000
0!
0*
09
0>
0C
#161590000000
1!
1*
b1 6
19
1>
1C
b1 G
#161600000000
0!
0*
09
0>
0C
#161610000000
1!
1*
b10 6
19
1>
1C
b10 G
#161620000000
0!
0*
09
0>
0C
#161630000000
1!
1*
b11 6
19
1>
1C
b11 G
#161640000000
0!
0*
09
0>
0C
#161650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#161660000000
0!
0*
09
0>
0C
#161670000000
1!
1*
b101 6
19
1>
1C
b101 G
#161680000000
0!
0*
09
0>
0C
#161690000000
1!
1*
b110 6
19
1>
1C
b110 G
#161700000000
0!
0*
09
0>
0C
#161710000000
1!
1*
b111 6
19
1>
1C
b111 G
#161720000000
0!
0*
09
0>
0C
#161730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#161740000000
0!
0*
09
0>
0C
#161750000000
1!
1*
b1 6
19
1>
1C
b1 G
#161760000000
0!
0*
09
0>
0C
#161770000000
1!
1*
b10 6
19
1>
1C
b10 G
#161780000000
0!
0*
09
0>
0C
#161790000000
1!
1*
b11 6
19
1>
1C
b11 G
#161800000000
0!
0*
09
0>
0C
#161810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#161820000000
0!
0*
09
0>
0C
#161830000000
1!
1*
b101 6
19
1>
1C
b101 G
#161840000000
0!
0*
09
0>
0C
#161850000000
1!
1*
b110 6
19
1>
1C
b110 G
#161860000000
0!
0*
09
0>
0C
#161870000000
1!
1*
b111 6
19
1>
1C
b111 G
#161880000000
0!
1"
0*
1+
09
1:
0>
0C
#161890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#161900000000
0!
0*
09
0>
0C
#161910000000
1!
1*
b1 6
19
1>
1C
b1 G
#161920000000
0!
0*
09
0>
0C
#161930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#161940000000
0!
0*
09
0>
0C
#161950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#161960000000
0!
0*
09
0>
0C
#161970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#161980000000
0!
0*
09
0>
0C
#161990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#162000000000
0!
0#
0*
0,
09
0>
0?
0C
#162010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#162020000000
0!
0*
09
0>
0C
#162030000000
1!
1*
19
1>
1C
#162040000000
0!
0*
09
0>
0C
#162050000000
1!
1*
19
1>
1C
#162060000000
0!
0*
09
0>
0C
#162070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#162080000000
0!
0*
09
0>
0C
#162090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#162100000000
0!
0*
09
0>
0C
#162110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#162120000000
0!
0*
09
0>
0C
#162130000000
1!
1*
b10 6
19
1>
1C
b10 G
#162140000000
0!
0*
09
0>
0C
#162150000000
1!
1*
b11 6
19
1>
1C
b11 G
#162160000000
0!
0*
09
0>
0C
#162170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#162180000000
0!
0*
09
0>
0C
#162190000000
1!
1*
b101 6
19
1>
1C
b101 G
#162200000000
0!
0*
09
0>
0C
#162210000000
1!
1*
b110 6
19
1>
1C
b110 G
#162220000000
0!
0*
09
0>
0C
#162230000000
1!
1*
b111 6
19
1>
1C
b111 G
#162240000000
0!
0*
09
0>
0C
#162250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#162260000000
0!
0*
09
0>
0C
#162270000000
1!
1*
b1 6
19
1>
1C
b1 G
#162280000000
0!
0*
09
0>
0C
#162290000000
1!
1*
b10 6
19
1>
1C
b10 G
#162300000000
0!
0*
09
0>
0C
#162310000000
1!
1*
b11 6
19
1>
1C
b11 G
#162320000000
0!
0*
09
0>
0C
#162330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#162340000000
0!
0*
09
0>
0C
#162350000000
1!
1*
b101 6
19
1>
1C
b101 G
#162360000000
0!
0*
09
0>
0C
#162370000000
1!
1*
b110 6
19
1>
1C
b110 G
#162380000000
0!
0*
09
0>
0C
#162390000000
1!
1*
b111 6
19
1>
1C
b111 G
#162400000000
0!
0*
09
0>
0C
#162410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#162420000000
0!
0*
09
0>
0C
#162430000000
1!
1*
b1 6
19
1>
1C
b1 G
#162440000000
0!
0*
09
0>
0C
#162450000000
1!
1*
b10 6
19
1>
1C
b10 G
#162460000000
0!
0*
09
0>
0C
#162470000000
1!
1*
b11 6
19
1>
1C
b11 G
#162480000000
0!
0*
09
0>
0C
#162490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#162500000000
0!
0*
09
0>
0C
#162510000000
1!
1*
b101 6
19
1>
1C
b101 G
#162520000000
0!
0*
09
0>
0C
#162530000000
1!
1*
b110 6
19
1>
1C
b110 G
#162540000000
0!
0*
09
0>
0C
#162550000000
1!
1*
b111 6
19
1>
1C
b111 G
#162560000000
0!
1"
0*
1+
09
1:
0>
0C
#162570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#162580000000
0!
0*
09
0>
0C
#162590000000
1!
1*
b1 6
19
1>
1C
b1 G
#162600000000
0!
0*
09
0>
0C
#162610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#162620000000
0!
0*
09
0>
0C
#162630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#162640000000
0!
0*
09
0>
0C
#162650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#162660000000
0!
0*
09
0>
0C
#162670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#162680000000
0!
0#
0*
0,
09
0>
0?
0C
#162690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#162700000000
0!
0*
09
0>
0C
#162710000000
1!
1*
19
1>
1C
#162720000000
0!
0*
09
0>
0C
#162730000000
1!
1*
19
1>
1C
#162740000000
0!
0*
09
0>
0C
#162750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#162760000000
0!
0*
09
0>
0C
#162770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#162780000000
0!
0*
09
0>
0C
#162790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#162800000000
0!
0*
09
0>
0C
#162810000000
1!
1*
b10 6
19
1>
1C
b10 G
#162820000000
0!
0*
09
0>
0C
#162830000000
1!
1*
b11 6
19
1>
1C
b11 G
#162840000000
0!
0*
09
0>
0C
#162850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#162860000000
0!
0*
09
0>
0C
#162870000000
1!
1*
b101 6
19
1>
1C
b101 G
#162880000000
0!
0*
09
0>
0C
#162890000000
1!
1*
b110 6
19
1>
1C
b110 G
#162900000000
0!
0*
09
0>
0C
#162910000000
1!
1*
b111 6
19
1>
1C
b111 G
#162920000000
0!
0*
09
0>
0C
#162930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#162940000000
0!
0*
09
0>
0C
#162950000000
1!
1*
b1 6
19
1>
1C
b1 G
#162960000000
0!
0*
09
0>
0C
#162970000000
1!
1*
b10 6
19
1>
1C
b10 G
#162980000000
0!
0*
09
0>
0C
#162990000000
1!
1*
b11 6
19
1>
1C
b11 G
#163000000000
0!
0*
09
0>
0C
#163010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#163020000000
0!
0*
09
0>
0C
#163030000000
1!
1*
b101 6
19
1>
1C
b101 G
#163040000000
0!
0*
09
0>
0C
#163050000000
1!
1*
b110 6
19
1>
1C
b110 G
#163060000000
0!
0*
09
0>
0C
#163070000000
1!
1*
b111 6
19
1>
1C
b111 G
#163080000000
0!
0*
09
0>
0C
#163090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#163100000000
0!
0*
09
0>
0C
#163110000000
1!
1*
b1 6
19
1>
1C
b1 G
#163120000000
0!
0*
09
0>
0C
#163130000000
1!
1*
b10 6
19
1>
1C
b10 G
#163140000000
0!
0*
09
0>
0C
#163150000000
1!
1*
b11 6
19
1>
1C
b11 G
#163160000000
0!
0*
09
0>
0C
#163170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#163180000000
0!
0*
09
0>
0C
#163190000000
1!
1*
b101 6
19
1>
1C
b101 G
#163200000000
0!
0*
09
0>
0C
#163210000000
1!
1*
b110 6
19
1>
1C
b110 G
#163220000000
0!
0*
09
0>
0C
#163230000000
1!
1*
b111 6
19
1>
1C
b111 G
#163240000000
0!
1"
0*
1+
09
1:
0>
0C
#163250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#163260000000
0!
0*
09
0>
0C
#163270000000
1!
1*
b1 6
19
1>
1C
b1 G
#163280000000
0!
0*
09
0>
0C
#163290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#163300000000
0!
0*
09
0>
0C
#163310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#163320000000
0!
0*
09
0>
0C
#163330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#163340000000
0!
0*
09
0>
0C
#163350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#163360000000
0!
0#
0*
0,
09
0>
0?
0C
#163370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#163380000000
0!
0*
09
0>
0C
#163390000000
1!
1*
19
1>
1C
#163400000000
0!
0*
09
0>
0C
#163410000000
1!
1*
19
1>
1C
#163420000000
0!
0*
09
0>
0C
#163430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#163440000000
0!
0*
09
0>
0C
#163450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#163460000000
0!
0*
09
0>
0C
#163470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#163480000000
0!
0*
09
0>
0C
#163490000000
1!
1*
b10 6
19
1>
1C
b10 G
#163500000000
0!
0*
09
0>
0C
#163510000000
1!
1*
b11 6
19
1>
1C
b11 G
#163520000000
0!
0*
09
0>
0C
#163530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#163540000000
0!
0*
09
0>
0C
#163550000000
1!
1*
b101 6
19
1>
1C
b101 G
#163560000000
0!
0*
09
0>
0C
#163570000000
1!
1*
b110 6
19
1>
1C
b110 G
#163580000000
0!
0*
09
0>
0C
#163590000000
1!
1*
b111 6
19
1>
1C
b111 G
#163600000000
0!
0*
09
0>
0C
#163610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#163620000000
0!
0*
09
0>
0C
#163630000000
1!
1*
b1 6
19
1>
1C
b1 G
#163640000000
0!
0*
09
0>
0C
#163650000000
1!
1*
b10 6
19
1>
1C
b10 G
#163660000000
0!
0*
09
0>
0C
#163670000000
1!
1*
b11 6
19
1>
1C
b11 G
#163680000000
0!
0*
09
0>
0C
#163690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#163700000000
0!
0*
09
0>
0C
#163710000000
1!
1*
b101 6
19
1>
1C
b101 G
#163720000000
0!
0*
09
0>
0C
#163730000000
1!
1*
b110 6
19
1>
1C
b110 G
#163740000000
0!
0*
09
0>
0C
#163750000000
1!
1*
b111 6
19
1>
1C
b111 G
#163760000000
0!
0*
09
0>
0C
#163770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#163780000000
0!
0*
09
0>
0C
#163790000000
1!
1*
b1 6
19
1>
1C
b1 G
#163800000000
0!
0*
09
0>
0C
#163810000000
1!
1*
b10 6
19
1>
1C
b10 G
#163820000000
0!
0*
09
0>
0C
#163830000000
1!
1*
b11 6
19
1>
1C
b11 G
#163840000000
0!
0*
09
0>
0C
#163850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#163860000000
0!
0*
09
0>
0C
#163870000000
1!
1*
b101 6
19
1>
1C
b101 G
#163880000000
0!
0*
09
0>
0C
#163890000000
1!
1*
b110 6
19
1>
1C
b110 G
#163900000000
0!
0*
09
0>
0C
#163910000000
1!
1*
b111 6
19
1>
1C
b111 G
#163920000000
0!
1"
0*
1+
09
1:
0>
0C
#163930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#163940000000
0!
0*
09
0>
0C
#163950000000
1!
1*
b1 6
19
1>
1C
b1 G
#163960000000
0!
0*
09
0>
0C
#163970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#163980000000
0!
0*
09
0>
0C
#163990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#164000000000
0!
0*
09
0>
0C
#164010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#164020000000
0!
0*
09
0>
0C
#164030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#164040000000
0!
0#
0*
0,
09
0>
0?
0C
#164050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#164060000000
0!
0*
09
0>
0C
#164070000000
1!
1*
19
1>
1C
#164080000000
0!
0*
09
0>
0C
#164090000000
1!
1*
19
1>
1C
#164100000000
0!
0*
09
0>
0C
#164110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#164120000000
0!
0*
09
0>
0C
#164130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#164140000000
0!
0*
09
0>
0C
#164150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#164160000000
0!
0*
09
0>
0C
#164170000000
1!
1*
b10 6
19
1>
1C
b10 G
#164180000000
0!
0*
09
0>
0C
#164190000000
1!
1*
b11 6
19
1>
1C
b11 G
#164200000000
0!
0*
09
0>
0C
#164210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#164220000000
0!
0*
09
0>
0C
#164230000000
1!
1*
b101 6
19
1>
1C
b101 G
#164240000000
0!
0*
09
0>
0C
#164250000000
1!
1*
b110 6
19
1>
1C
b110 G
#164260000000
0!
0*
09
0>
0C
#164270000000
1!
1*
b111 6
19
1>
1C
b111 G
#164280000000
0!
0*
09
0>
0C
#164290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#164300000000
0!
0*
09
0>
0C
#164310000000
1!
1*
b1 6
19
1>
1C
b1 G
#164320000000
0!
0*
09
0>
0C
#164330000000
1!
1*
b10 6
19
1>
1C
b10 G
#164340000000
0!
0*
09
0>
0C
#164350000000
1!
1*
b11 6
19
1>
1C
b11 G
#164360000000
0!
0*
09
0>
0C
#164370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#164380000000
0!
0*
09
0>
0C
#164390000000
1!
1*
b101 6
19
1>
1C
b101 G
#164400000000
0!
0*
09
0>
0C
#164410000000
1!
1*
b110 6
19
1>
1C
b110 G
#164420000000
0!
0*
09
0>
0C
#164430000000
1!
1*
b111 6
19
1>
1C
b111 G
#164440000000
0!
0*
09
0>
0C
#164450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#164460000000
0!
0*
09
0>
0C
#164470000000
1!
1*
b1 6
19
1>
1C
b1 G
#164480000000
0!
0*
09
0>
0C
#164490000000
1!
1*
b10 6
19
1>
1C
b10 G
#164500000000
0!
0*
09
0>
0C
#164510000000
1!
1*
b11 6
19
1>
1C
b11 G
#164520000000
0!
0*
09
0>
0C
#164530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#164540000000
0!
0*
09
0>
0C
#164550000000
1!
1*
b101 6
19
1>
1C
b101 G
#164560000000
0!
0*
09
0>
0C
#164570000000
1!
1*
b110 6
19
1>
1C
b110 G
#164580000000
0!
0*
09
0>
0C
#164590000000
1!
1*
b111 6
19
1>
1C
b111 G
#164600000000
0!
1"
0*
1+
09
1:
0>
0C
#164610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#164620000000
0!
0*
09
0>
0C
#164630000000
1!
1*
b1 6
19
1>
1C
b1 G
#164640000000
0!
0*
09
0>
0C
#164650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#164660000000
0!
0*
09
0>
0C
#164670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#164680000000
0!
0*
09
0>
0C
#164690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#164700000000
0!
0*
09
0>
0C
#164710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#164720000000
0!
0#
0*
0,
09
0>
0?
0C
#164730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#164740000000
0!
0*
09
0>
0C
#164750000000
1!
1*
19
1>
1C
#164760000000
0!
0*
09
0>
0C
#164770000000
1!
1*
19
1>
1C
#164780000000
0!
0*
09
0>
0C
#164790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#164800000000
0!
0*
09
0>
0C
#164810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#164820000000
0!
0*
09
0>
0C
#164830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#164840000000
0!
0*
09
0>
0C
#164850000000
1!
1*
b10 6
19
1>
1C
b10 G
#164860000000
0!
0*
09
0>
0C
#164870000000
1!
1*
b11 6
19
1>
1C
b11 G
#164880000000
0!
0*
09
0>
0C
#164890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#164900000000
0!
0*
09
0>
0C
#164910000000
1!
1*
b101 6
19
1>
1C
b101 G
#164920000000
0!
0*
09
0>
0C
#164930000000
1!
1*
b110 6
19
1>
1C
b110 G
#164940000000
0!
0*
09
0>
0C
#164950000000
1!
1*
b111 6
19
1>
1C
b111 G
#164960000000
0!
0*
09
0>
0C
#164970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#164980000000
0!
0*
09
0>
0C
#164990000000
1!
1*
b1 6
19
1>
1C
b1 G
#165000000000
0!
0*
09
0>
0C
#165010000000
1!
1*
b10 6
19
1>
1C
b10 G
#165020000000
0!
0*
09
0>
0C
#165030000000
1!
1*
b11 6
19
1>
1C
b11 G
#165040000000
0!
0*
09
0>
0C
#165050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#165060000000
0!
0*
09
0>
0C
#165070000000
1!
1*
b101 6
19
1>
1C
b101 G
#165080000000
0!
0*
09
0>
0C
#165090000000
1!
1*
b110 6
19
1>
1C
b110 G
#165100000000
0!
0*
09
0>
0C
#165110000000
1!
1*
b111 6
19
1>
1C
b111 G
#165120000000
0!
0*
09
0>
0C
#165130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#165140000000
0!
0*
09
0>
0C
#165150000000
1!
1*
b1 6
19
1>
1C
b1 G
#165160000000
0!
0*
09
0>
0C
#165170000000
1!
1*
b10 6
19
1>
1C
b10 G
#165180000000
0!
0*
09
0>
0C
#165190000000
1!
1*
b11 6
19
1>
1C
b11 G
#165200000000
0!
0*
09
0>
0C
#165210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#165220000000
0!
0*
09
0>
0C
#165230000000
1!
1*
b101 6
19
1>
1C
b101 G
#165240000000
0!
0*
09
0>
0C
#165250000000
1!
1*
b110 6
19
1>
1C
b110 G
#165260000000
0!
0*
09
0>
0C
#165270000000
1!
1*
b111 6
19
1>
1C
b111 G
#165280000000
0!
1"
0*
1+
09
1:
0>
0C
#165290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#165300000000
0!
0*
09
0>
0C
#165310000000
1!
1*
b1 6
19
1>
1C
b1 G
#165320000000
0!
0*
09
0>
0C
#165330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#165340000000
0!
0*
09
0>
0C
#165350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#165360000000
0!
0*
09
0>
0C
#165370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#165380000000
0!
0*
09
0>
0C
#165390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#165400000000
0!
0#
0*
0,
09
0>
0?
0C
#165410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#165420000000
0!
0*
09
0>
0C
#165430000000
1!
1*
19
1>
1C
#165440000000
0!
0*
09
0>
0C
#165450000000
1!
1*
19
1>
1C
#165460000000
0!
0*
09
0>
0C
#165470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#165480000000
0!
0*
09
0>
0C
#165490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#165500000000
0!
0*
09
0>
0C
#165510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#165520000000
0!
0*
09
0>
0C
#165530000000
1!
1*
b10 6
19
1>
1C
b10 G
#165540000000
0!
0*
09
0>
0C
#165550000000
1!
1*
b11 6
19
1>
1C
b11 G
#165560000000
0!
0*
09
0>
0C
#165570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#165580000000
0!
0*
09
0>
0C
#165590000000
1!
1*
b101 6
19
1>
1C
b101 G
#165600000000
0!
0*
09
0>
0C
#165610000000
1!
1*
b110 6
19
1>
1C
b110 G
#165620000000
0!
0*
09
0>
0C
#165630000000
1!
1*
b111 6
19
1>
1C
b111 G
#165640000000
0!
0*
09
0>
0C
#165650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#165660000000
0!
0*
09
0>
0C
#165670000000
1!
1*
b1 6
19
1>
1C
b1 G
#165680000000
0!
0*
09
0>
0C
#165690000000
1!
1*
b10 6
19
1>
1C
b10 G
#165700000000
0!
0*
09
0>
0C
#165710000000
1!
1*
b11 6
19
1>
1C
b11 G
#165720000000
0!
0*
09
0>
0C
#165730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#165740000000
0!
0*
09
0>
0C
#165750000000
1!
1*
b101 6
19
1>
1C
b101 G
#165760000000
0!
0*
09
0>
0C
#165770000000
1!
1*
b110 6
19
1>
1C
b110 G
#165780000000
0!
0*
09
0>
0C
#165790000000
1!
1*
b111 6
19
1>
1C
b111 G
#165800000000
0!
0*
09
0>
0C
#165810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#165820000000
0!
0*
09
0>
0C
#165830000000
1!
1*
b1 6
19
1>
1C
b1 G
#165840000000
0!
0*
09
0>
0C
#165850000000
1!
1*
b10 6
19
1>
1C
b10 G
#165860000000
0!
0*
09
0>
0C
#165870000000
1!
1*
b11 6
19
1>
1C
b11 G
#165880000000
0!
0*
09
0>
0C
#165890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#165900000000
0!
0*
09
0>
0C
#165910000000
1!
1*
b101 6
19
1>
1C
b101 G
#165920000000
0!
0*
09
0>
0C
#165930000000
1!
1*
b110 6
19
1>
1C
b110 G
#165940000000
0!
0*
09
0>
0C
#165950000000
1!
1*
b111 6
19
1>
1C
b111 G
#165960000000
0!
1"
0*
1+
09
1:
0>
0C
#165970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#165980000000
0!
0*
09
0>
0C
#165990000000
1!
1*
b1 6
19
1>
1C
b1 G
#166000000000
0!
0*
09
0>
0C
#166010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#166020000000
0!
0*
09
0>
0C
#166030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#166040000000
0!
0*
09
0>
0C
#166050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#166060000000
0!
0*
09
0>
0C
#166070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#166080000000
0!
0#
0*
0,
09
0>
0?
0C
#166090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#166100000000
0!
0*
09
0>
0C
#166110000000
1!
1*
19
1>
1C
#166120000000
0!
0*
09
0>
0C
#166130000000
1!
1*
19
1>
1C
#166140000000
0!
0*
09
0>
0C
#166150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#166160000000
0!
0*
09
0>
0C
#166170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#166180000000
0!
0*
09
0>
0C
#166190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#166200000000
0!
0*
09
0>
0C
#166210000000
1!
1*
b10 6
19
1>
1C
b10 G
#166220000000
0!
0*
09
0>
0C
#166230000000
1!
1*
b11 6
19
1>
1C
b11 G
#166240000000
0!
0*
09
0>
0C
#166250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#166260000000
0!
0*
09
0>
0C
#166270000000
1!
1*
b101 6
19
1>
1C
b101 G
#166280000000
0!
0*
09
0>
0C
#166290000000
1!
1*
b110 6
19
1>
1C
b110 G
#166300000000
0!
0*
09
0>
0C
#166310000000
1!
1*
b111 6
19
1>
1C
b111 G
#166320000000
0!
0*
09
0>
0C
#166330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#166340000000
0!
0*
09
0>
0C
#166350000000
1!
1*
b1 6
19
1>
1C
b1 G
#166360000000
0!
0*
09
0>
0C
#166370000000
1!
1*
b10 6
19
1>
1C
b10 G
#166380000000
0!
0*
09
0>
0C
#166390000000
1!
1*
b11 6
19
1>
1C
b11 G
#166400000000
0!
0*
09
0>
0C
#166410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#166420000000
0!
0*
09
0>
0C
#166430000000
1!
1*
b101 6
19
1>
1C
b101 G
#166440000000
0!
0*
09
0>
0C
#166450000000
1!
1*
b110 6
19
1>
1C
b110 G
#166460000000
0!
0*
09
0>
0C
#166470000000
1!
1*
b111 6
19
1>
1C
b111 G
#166480000000
0!
0*
09
0>
0C
#166490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#166500000000
0!
0*
09
0>
0C
#166510000000
1!
1*
b1 6
19
1>
1C
b1 G
#166520000000
0!
0*
09
0>
0C
#166530000000
1!
1*
b10 6
19
1>
1C
b10 G
#166540000000
0!
0*
09
0>
0C
#166550000000
1!
1*
b11 6
19
1>
1C
b11 G
#166560000000
0!
0*
09
0>
0C
#166570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#166580000000
0!
0*
09
0>
0C
#166590000000
1!
1*
b101 6
19
1>
1C
b101 G
#166600000000
0!
0*
09
0>
0C
#166610000000
1!
1*
b110 6
19
1>
1C
b110 G
#166620000000
0!
0*
09
0>
0C
#166630000000
1!
1*
b111 6
19
1>
1C
b111 G
#166640000000
0!
1"
0*
1+
09
1:
0>
0C
#166650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#166660000000
0!
0*
09
0>
0C
#166670000000
1!
1*
b1 6
19
1>
1C
b1 G
#166680000000
0!
0*
09
0>
0C
#166690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#166700000000
0!
0*
09
0>
0C
#166710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#166720000000
0!
0*
09
0>
0C
#166730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#166740000000
0!
0*
09
0>
0C
#166750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#166760000000
0!
0#
0*
0,
09
0>
0?
0C
#166770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#166780000000
0!
0*
09
0>
0C
#166790000000
1!
1*
19
1>
1C
#166800000000
0!
0*
09
0>
0C
#166810000000
1!
1*
19
1>
1C
#166820000000
0!
0*
09
0>
0C
#166830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#166840000000
0!
0*
09
0>
0C
#166850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#166860000000
0!
0*
09
0>
0C
#166870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#166880000000
0!
0*
09
0>
0C
#166890000000
1!
1*
b10 6
19
1>
1C
b10 G
#166900000000
0!
0*
09
0>
0C
#166910000000
1!
1*
b11 6
19
1>
1C
b11 G
#166920000000
0!
0*
09
0>
0C
#166930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#166940000000
0!
0*
09
0>
0C
#166950000000
1!
1*
b101 6
19
1>
1C
b101 G
#166960000000
0!
0*
09
0>
0C
#166970000000
1!
1*
b110 6
19
1>
1C
b110 G
#166980000000
0!
0*
09
0>
0C
#166990000000
1!
1*
b111 6
19
1>
1C
b111 G
#167000000000
0!
0*
09
0>
0C
#167010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#167020000000
0!
0*
09
0>
0C
#167030000000
1!
1*
b1 6
19
1>
1C
b1 G
#167040000000
0!
0*
09
0>
0C
#167050000000
1!
1*
b10 6
19
1>
1C
b10 G
#167060000000
0!
0*
09
0>
0C
#167070000000
1!
1*
b11 6
19
1>
1C
b11 G
#167080000000
0!
0*
09
0>
0C
#167090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#167100000000
0!
0*
09
0>
0C
#167110000000
1!
1*
b101 6
19
1>
1C
b101 G
#167120000000
0!
0*
09
0>
0C
#167130000000
1!
1*
b110 6
19
1>
1C
b110 G
#167140000000
0!
0*
09
0>
0C
#167150000000
1!
1*
b111 6
19
1>
1C
b111 G
#167160000000
0!
0*
09
0>
0C
#167170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#167180000000
0!
0*
09
0>
0C
#167190000000
1!
1*
b1 6
19
1>
1C
b1 G
#167200000000
0!
0*
09
0>
0C
#167210000000
1!
1*
b10 6
19
1>
1C
b10 G
#167220000000
0!
0*
09
0>
0C
#167230000000
1!
1*
b11 6
19
1>
1C
b11 G
#167240000000
0!
0*
09
0>
0C
#167250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#167260000000
0!
0*
09
0>
0C
#167270000000
1!
1*
b101 6
19
1>
1C
b101 G
#167280000000
0!
0*
09
0>
0C
#167290000000
1!
1*
b110 6
19
1>
1C
b110 G
#167300000000
0!
0*
09
0>
0C
#167310000000
1!
1*
b111 6
19
1>
1C
b111 G
#167320000000
0!
1"
0*
1+
09
1:
0>
0C
#167330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#167340000000
0!
0*
09
0>
0C
#167350000000
1!
1*
b1 6
19
1>
1C
b1 G
#167360000000
0!
0*
09
0>
0C
#167370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#167380000000
0!
0*
09
0>
0C
#167390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#167400000000
0!
0*
09
0>
0C
#167410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#167420000000
0!
0*
09
0>
0C
#167430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#167440000000
0!
0#
0*
0,
09
0>
0?
0C
#167450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#167460000000
0!
0*
09
0>
0C
#167470000000
1!
1*
19
1>
1C
#167480000000
0!
0*
09
0>
0C
#167490000000
1!
1*
19
1>
1C
#167500000000
0!
0*
09
0>
0C
#167510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#167520000000
0!
0*
09
0>
0C
#167530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#167540000000
0!
0*
09
0>
0C
#167550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#167560000000
0!
0*
09
0>
0C
#167570000000
1!
1*
b10 6
19
1>
1C
b10 G
#167580000000
0!
0*
09
0>
0C
#167590000000
1!
1*
b11 6
19
1>
1C
b11 G
#167600000000
0!
0*
09
0>
0C
#167610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#167620000000
0!
0*
09
0>
0C
#167630000000
1!
1*
b101 6
19
1>
1C
b101 G
#167640000000
0!
0*
09
0>
0C
#167650000000
1!
1*
b110 6
19
1>
1C
b110 G
#167660000000
0!
0*
09
0>
0C
#167670000000
1!
1*
b111 6
19
1>
1C
b111 G
#167680000000
0!
0*
09
0>
0C
#167690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#167700000000
0!
0*
09
0>
0C
#167710000000
1!
1*
b1 6
19
1>
1C
b1 G
#167720000000
0!
0*
09
0>
0C
#167730000000
1!
1*
b10 6
19
1>
1C
b10 G
#167740000000
0!
0*
09
0>
0C
#167750000000
1!
1*
b11 6
19
1>
1C
b11 G
#167760000000
0!
0*
09
0>
0C
#167770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#167780000000
0!
0*
09
0>
0C
#167790000000
1!
1*
b101 6
19
1>
1C
b101 G
#167800000000
0!
0*
09
0>
0C
#167810000000
1!
1*
b110 6
19
1>
1C
b110 G
#167820000000
0!
0*
09
0>
0C
#167830000000
1!
1*
b111 6
19
1>
1C
b111 G
#167840000000
0!
0*
09
0>
0C
#167850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#167860000000
0!
0*
09
0>
0C
#167870000000
1!
1*
b1 6
19
1>
1C
b1 G
#167880000000
0!
0*
09
0>
0C
#167890000000
1!
1*
b10 6
19
1>
1C
b10 G
#167900000000
0!
0*
09
0>
0C
#167910000000
1!
1*
b11 6
19
1>
1C
b11 G
#167920000000
0!
0*
09
0>
0C
#167930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#167940000000
0!
0*
09
0>
0C
#167950000000
1!
1*
b101 6
19
1>
1C
b101 G
#167960000000
0!
0*
09
0>
0C
#167970000000
1!
1*
b110 6
19
1>
1C
b110 G
#167980000000
0!
0*
09
0>
0C
#167990000000
1!
1*
b111 6
19
1>
1C
b111 G
#168000000000
0!
1"
0*
1+
09
1:
0>
0C
#168010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#168020000000
0!
0*
09
0>
0C
#168030000000
1!
1*
b1 6
19
1>
1C
b1 G
#168040000000
0!
0*
09
0>
0C
#168050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#168060000000
0!
0*
09
0>
0C
#168070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#168080000000
0!
0*
09
0>
0C
#168090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#168100000000
0!
0*
09
0>
0C
#168110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#168120000000
0!
0#
0*
0,
09
0>
0?
0C
#168130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#168140000000
0!
0*
09
0>
0C
#168150000000
1!
1*
19
1>
1C
#168160000000
0!
0*
09
0>
0C
#168170000000
1!
1*
19
1>
1C
#168180000000
0!
0*
09
0>
0C
#168190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#168200000000
0!
0*
09
0>
0C
#168210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#168220000000
0!
0*
09
0>
0C
#168230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#168240000000
0!
0*
09
0>
0C
#168250000000
1!
1*
b10 6
19
1>
1C
b10 G
#168260000000
0!
0*
09
0>
0C
#168270000000
1!
1*
b11 6
19
1>
1C
b11 G
#168280000000
0!
0*
09
0>
0C
#168290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#168300000000
0!
0*
09
0>
0C
#168310000000
1!
1*
b101 6
19
1>
1C
b101 G
#168320000000
0!
0*
09
0>
0C
#168330000000
1!
1*
b110 6
19
1>
1C
b110 G
#168340000000
0!
0*
09
0>
0C
#168350000000
1!
1*
b111 6
19
1>
1C
b111 G
#168360000000
0!
0*
09
0>
0C
#168370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#168380000000
0!
0*
09
0>
0C
#168390000000
1!
1*
b1 6
19
1>
1C
b1 G
#168400000000
0!
0*
09
0>
0C
#168410000000
1!
1*
b10 6
19
1>
1C
b10 G
#168420000000
0!
0*
09
0>
0C
#168430000000
1!
1*
b11 6
19
1>
1C
b11 G
#168440000000
0!
0*
09
0>
0C
#168450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#168460000000
0!
0*
09
0>
0C
#168470000000
1!
1*
b101 6
19
1>
1C
b101 G
#168480000000
0!
0*
09
0>
0C
#168490000000
1!
1*
b110 6
19
1>
1C
b110 G
#168500000000
0!
0*
09
0>
0C
#168510000000
1!
1*
b111 6
19
1>
1C
b111 G
#168520000000
0!
0*
09
0>
0C
#168530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#168540000000
0!
0*
09
0>
0C
#168550000000
1!
1*
b1 6
19
1>
1C
b1 G
#168560000000
0!
0*
09
0>
0C
#168570000000
1!
1*
b10 6
19
1>
1C
b10 G
#168580000000
0!
0*
09
0>
0C
#168590000000
1!
1*
b11 6
19
1>
1C
b11 G
#168600000000
0!
0*
09
0>
0C
#168610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#168620000000
0!
0*
09
0>
0C
#168630000000
1!
1*
b101 6
19
1>
1C
b101 G
#168640000000
0!
0*
09
0>
0C
#168650000000
1!
1*
b110 6
19
1>
1C
b110 G
#168660000000
0!
0*
09
0>
0C
#168670000000
1!
1*
b111 6
19
1>
1C
b111 G
#168680000000
0!
1"
0*
1+
09
1:
0>
0C
#168690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#168700000000
0!
0*
09
0>
0C
#168710000000
1!
1*
b1 6
19
1>
1C
b1 G
#168720000000
0!
0*
09
0>
0C
#168730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#168740000000
0!
0*
09
0>
0C
#168750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#168760000000
0!
0*
09
0>
0C
#168770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#168780000000
0!
0*
09
0>
0C
#168790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#168800000000
0!
0#
0*
0,
09
0>
0?
0C
#168810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#168820000000
0!
0*
09
0>
0C
#168830000000
1!
1*
19
1>
1C
#168840000000
0!
0*
09
0>
0C
#168850000000
1!
1*
19
1>
1C
#168860000000
0!
0*
09
0>
0C
#168870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#168880000000
0!
0*
09
0>
0C
#168890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#168900000000
0!
0*
09
0>
0C
#168910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#168920000000
0!
0*
09
0>
0C
#168930000000
1!
1*
b10 6
19
1>
1C
b10 G
#168940000000
0!
0*
09
0>
0C
#168950000000
1!
1*
b11 6
19
1>
1C
b11 G
#168960000000
0!
0*
09
0>
0C
#168970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#168980000000
0!
0*
09
0>
0C
#168990000000
1!
1*
b101 6
19
1>
1C
b101 G
#169000000000
0!
0*
09
0>
0C
#169010000000
1!
1*
b110 6
19
1>
1C
b110 G
#169020000000
0!
0*
09
0>
0C
#169030000000
1!
1*
b111 6
19
1>
1C
b111 G
#169040000000
0!
0*
09
0>
0C
#169050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#169060000000
0!
0*
09
0>
0C
#169070000000
1!
1*
b1 6
19
1>
1C
b1 G
#169080000000
0!
0*
09
0>
0C
#169090000000
1!
1*
b10 6
19
1>
1C
b10 G
#169100000000
0!
0*
09
0>
0C
#169110000000
1!
1*
b11 6
19
1>
1C
b11 G
#169120000000
0!
0*
09
0>
0C
#169130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#169140000000
0!
0*
09
0>
0C
#169150000000
1!
1*
b101 6
19
1>
1C
b101 G
#169160000000
0!
0*
09
0>
0C
#169170000000
1!
1*
b110 6
19
1>
1C
b110 G
#169180000000
0!
0*
09
0>
0C
#169190000000
1!
1*
b111 6
19
1>
1C
b111 G
#169200000000
0!
0*
09
0>
0C
#169210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#169220000000
0!
0*
09
0>
0C
#169230000000
1!
1*
b1 6
19
1>
1C
b1 G
#169240000000
0!
0*
09
0>
0C
#169250000000
1!
1*
b10 6
19
1>
1C
b10 G
#169260000000
0!
0*
09
0>
0C
#169270000000
1!
1*
b11 6
19
1>
1C
b11 G
#169280000000
0!
0*
09
0>
0C
#169290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#169300000000
0!
0*
09
0>
0C
#169310000000
1!
1*
b101 6
19
1>
1C
b101 G
#169320000000
0!
0*
09
0>
0C
#169330000000
1!
1*
b110 6
19
1>
1C
b110 G
#169340000000
0!
0*
09
0>
0C
#169350000000
1!
1*
b111 6
19
1>
1C
b111 G
#169360000000
0!
1"
0*
1+
09
1:
0>
0C
#169370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#169380000000
0!
0*
09
0>
0C
#169390000000
1!
1*
b1 6
19
1>
1C
b1 G
#169400000000
0!
0*
09
0>
0C
#169410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#169420000000
0!
0*
09
0>
0C
#169430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#169440000000
0!
0*
09
0>
0C
#169450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#169460000000
0!
0*
09
0>
0C
#169470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#169480000000
0!
0#
0*
0,
09
0>
0?
0C
#169490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#169500000000
0!
0*
09
0>
0C
#169510000000
1!
1*
19
1>
1C
#169520000000
0!
0*
09
0>
0C
#169530000000
1!
1*
19
1>
1C
#169540000000
0!
0*
09
0>
0C
#169550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#169560000000
0!
0*
09
0>
0C
#169570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#169580000000
0!
0*
09
0>
0C
#169590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#169600000000
0!
0*
09
0>
0C
#169610000000
1!
1*
b10 6
19
1>
1C
b10 G
#169620000000
0!
0*
09
0>
0C
#169630000000
1!
1*
b11 6
19
1>
1C
b11 G
#169640000000
0!
0*
09
0>
0C
#169650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#169660000000
0!
0*
09
0>
0C
#169670000000
1!
1*
b101 6
19
1>
1C
b101 G
#169680000000
0!
0*
09
0>
0C
#169690000000
1!
1*
b110 6
19
1>
1C
b110 G
#169700000000
0!
0*
09
0>
0C
#169710000000
1!
1*
b111 6
19
1>
1C
b111 G
#169720000000
0!
0*
09
0>
0C
#169730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#169740000000
0!
0*
09
0>
0C
#169750000000
1!
1*
b1 6
19
1>
1C
b1 G
#169760000000
0!
0*
09
0>
0C
#169770000000
1!
1*
b10 6
19
1>
1C
b10 G
#169780000000
0!
0*
09
0>
0C
#169790000000
1!
1*
b11 6
19
1>
1C
b11 G
#169800000000
0!
0*
09
0>
0C
#169810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#169820000000
0!
0*
09
0>
0C
#169830000000
1!
1*
b101 6
19
1>
1C
b101 G
#169840000000
0!
0*
09
0>
0C
#169850000000
1!
1*
b110 6
19
1>
1C
b110 G
#169860000000
0!
0*
09
0>
0C
#169870000000
1!
1*
b111 6
19
1>
1C
b111 G
#169880000000
0!
0*
09
0>
0C
#169890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#169900000000
0!
0*
09
0>
0C
#169910000000
1!
1*
b1 6
19
1>
1C
b1 G
#169920000000
0!
0*
09
0>
0C
#169930000000
1!
1*
b10 6
19
1>
1C
b10 G
#169940000000
0!
0*
09
0>
0C
#169950000000
1!
1*
b11 6
19
1>
1C
b11 G
#169960000000
0!
0*
09
0>
0C
#169970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#169980000000
0!
0*
09
0>
0C
#169990000000
1!
1*
b101 6
19
1>
1C
b101 G
#170000000000
0!
0*
09
0>
0C
#170010000000
1!
1*
b110 6
19
1>
1C
b110 G
#170020000000
0!
0*
09
0>
0C
#170030000000
1!
1*
b111 6
19
1>
1C
b111 G
#170040000000
0!
1"
0*
1+
09
1:
0>
0C
#170050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#170060000000
0!
0*
09
0>
0C
#170070000000
1!
1*
b1 6
19
1>
1C
b1 G
#170080000000
0!
0*
09
0>
0C
#170090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#170100000000
0!
0*
09
0>
0C
#170110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#170120000000
0!
0*
09
0>
0C
#170130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#170140000000
0!
0*
09
0>
0C
#170150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#170160000000
0!
0#
0*
0,
09
0>
0?
0C
#170170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#170180000000
0!
0*
09
0>
0C
#170190000000
1!
1*
19
1>
1C
#170200000000
0!
0*
09
0>
0C
#170210000000
1!
1*
19
1>
1C
#170220000000
0!
0*
09
0>
0C
#170230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#170240000000
0!
0*
09
0>
0C
#170250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#170260000000
0!
0*
09
0>
0C
#170270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#170280000000
0!
0*
09
0>
0C
#170290000000
1!
1*
b10 6
19
1>
1C
b10 G
#170300000000
0!
0*
09
0>
0C
#170310000000
1!
1*
b11 6
19
1>
1C
b11 G
#170320000000
0!
0*
09
0>
0C
#170330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#170340000000
0!
0*
09
0>
0C
#170350000000
1!
1*
b101 6
19
1>
1C
b101 G
#170360000000
0!
0*
09
0>
0C
#170370000000
1!
1*
b110 6
19
1>
1C
b110 G
#170380000000
0!
0*
09
0>
0C
#170390000000
1!
1*
b111 6
19
1>
1C
b111 G
#170400000000
0!
0*
09
0>
0C
#170410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#170420000000
0!
0*
09
0>
0C
#170430000000
1!
1*
b1 6
19
1>
1C
b1 G
#170440000000
0!
0*
09
0>
0C
#170450000000
1!
1*
b10 6
19
1>
1C
b10 G
#170460000000
0!
0*
09
0>
0C
#170470000000
1!
1*
b11 6
19
1>
1C
b11 G
#170480000000
0!
0*
09
0>
0C
#170490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#170500000000
0!
0*
09
0>
0C
#170510000000
1!
1*
b101 6
19
1>
1C
b101 G
#170520000000
0!
0*
09
0>
0C
#170530000000
1!
1*
b110 6
19
1>
1C
b110 G
#170540000000
0!
0*
09
0>
0C
#170550000000
1!
1*
b111 6
19
1>
1C
b111 G
#170560000000
0!
0*
09
0>
0C
#170570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#170580000000
0!
0*
09
0>
0C
#170590000000
1!
1*
b1 6
19
1>
1C
b1 G
#170600000000
0!
0*
09
0>
0C
#170610000000
1!
1*
b10 6
19
1>
1C
b10 G
#170620000000
0!
0*
09
0>
0C
#170630000000
1!
1*
b11 6
19
1>
1C
b11 G
#170640000000
0!
0*
09
0>
0C
#170650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#170660000000
0!
0*
09
0>
0C
#170670000000
1!
1*
b101 6
19
1>
1C
b101 G
#170680000000
0!
0*
09
0>
0C
#170690000000
1!
1*
b110 6
19
1>
1C
b110 G
#170700000000
0!
0*
09
0>
0C
#170710000000
1!
1*
b111 6
19
1>
1C
b111 G
#170720000000
0!
1"
0*
1+
09
1:
0>
0C
#170730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#170740000000
0!
0*
09
0>
0C
#170750000000
1!
1*
b1 6
19
1>
1C
b1 G
#170760000000
0!
0*
09
0>
0C
#170770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#170780000000
0!
0*
09
0>
0C
#170790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#170800000000
0!
0*
09
0>
0C
#170810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#170820000000
0!
0*
09
0>
0C
#170830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#170840000000
0!
0#
0*
0,
09
0>
0?
0C
#170850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#170860000000
0!
0*
09
0>
0C
#170870000000
1!
1*
19
1>
1C
#170880000000
0!
0*
09
0>
0C
#170890000000
1!
1*
19
1>
1C
#170900000000
0!
0*
09
0>
0C
#170910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#170920000000
0!
0*
09
0>
0C
#170930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#170940000000
0!
0*
09
0>
0C
#170950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#170960000000
0!
0*
09
0>
0C
#170970000000
1!
1*
b10 6
19
1>
1C
b10 G
#170980000000
0!
0*
09
0>
0C
#170990000000
1!
1*
b11 6
19
1>
1C
b11 G
#171000000000
0!
0*
09
0>
0C
#171010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#171020000000
0!
0*
09
0>
0C
#171030000000
1!
1*
b101 6
19
1>
1C
b101 G
#171040000000
0!
0*
09
0>
0C
#171050000000
1!
1*
b110 6
19
1>
1C
b110 G
#171060000000
0!
0*
09
0>
0C
#171070000000
1!
1*
b111 6
19
1>
1C
b111 G
#171080000000
0!
0*
09
0>
0C
#171090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#171100000000
0!
0*
09
0>
0C
#171110000000
1!
1*
b1 6
19
1>
1C
b1 G
#171120000000
0!
0*
09
0>
0C
#171130000000
1!
1*
b10 6
19
1>
1C
b10 G
#171140000000
0!
0*
09
0>
0C
#171150000000
1!
1*
b11 6
19
1>
1C
b11 G
#171160000000
0!
0*
09
0>
0C
#171170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#171180000000
0!
0*
09
0>
0C
#171190000000
1!
1*
b101 6
19
1>
1C
b101 G
#171200000000
0!
0*
09
0>
0C
#171210000000
1!
1*
b110 6
19
1>
1C
b110 G
#171220000000
0!
0*
09
0>
0C
#171230000000
1!
1*
b111 6
19
1>
1C
b111 G
#171240000000
0!
0*
09
0>
0C
#171250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#171260000000
0!
0*
09
0>
0C
#171270000000
1!
1*
b1 6
19
1>
1C
b1 G
#171280000000
0!
0*
09
0>
0C
#171290000000
1!
1*
b10 6
19
1>
1C
b10 G
#171300000000
0!
0*
09
0>
0C
#171310000000
1!
1*
b11 6
19
1>
1C
b11 G
#171320000000
0!
0*
09
0>
0C
#171330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#171340000000
0!
0*
09
0>
0C
#171350000000
1!
1*
b101 6
19
1>
1C
b101 G
#171360000000
0!
0*
09
0>
0C
#171370000000
1!
1*
b110 6
19
1>
1C
b110 G
#171380000000
0!
0*
09
0>
0C
#171390000000
1!
1*
b111 6
19
1>
1C
b111 G
#171400000000
0!
1"
0*
1+
09
1:
0>
0C
#171410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#171420000000
0!
0*
09
0>
0C
#171430000000
1!
1*
b1 6
19
1>
1C
b1 G
#171440000000
0!
0*
09
0>
0C
#171450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#171460000000
0!
0*
09
0>
0C
#171470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#171480000000
0!
0*
09
0>
0C
#171490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#171500000000
0!
0*
09
0>
0C
#171510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#171520000000
0!
0#
0*
0,
09
0>
0?
0C
#171530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#171540000000
0!
0*
09
0>
0C
#171550000000
1!
1*
19
1>
1C
#171560000000
0!
0*
09
0>
0C
#171570000000
1!
1*
19
1>
1C
#171580000000
0!
0*
09
0>
0C
#171590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#171600000000
0!
0*
09
0>
0C
#171610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#171620000000
0!
0*
09
0>
0C
#171630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#171640000000
0!
0*
09
0>
0C
#171650000000
1!
1*
b10 6
19
1>
1C
b10 G
#171660000000
0!
0*
09
0>
0C
#171670000000
1!
1*
b11 6
19
1>
1C
b11 G
#171680000000
0!
0*
09
0>
0C
#171690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#171700000000
0!
0*
09
0>
0C
#171710000000
1!
1*
b101 6
19
1>
1C
b101 G
#171720000000
0!
0*
09
0>
0C
#171730000000
1!
1*
b110 6
19
1>
1C
b110 G
#171740000000
0!
0*
09
0>
0C
#171750000000
1!
1*
b111 6
19
1>
1C
b111 G
#171760000000
0!
0*
09
0>
0C
#171770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#171780000000
0!
0*
09
0>
0C
#171790000000
1!
1*
b1 6
19
1>
1C
b1 G
#171800000000
0!
0*
09
0>
0C
#171810000000
1!
1*
b10 6
19
1>
1C
b10 G
#171820000000
0!
0*
09
0>
0C
#171830000000
1!
1*
b11 6
19
1>
1C
b11 G
#171840000000
0!
0*
09
0>
0C
#171850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#171860000000
0!
0*
09
0>
0C
#171870000000
1!
1*
b101 6
19
1>
1C
b101 G
#171880000000
0!
0*
09
0>
0C
#171890000000
1!
1*
b110 6
19
1>
1C
b110 G
#171900000000
0!
0*
09
0>
0C
#171910000000
1!
1*
b111 6
19
1>
1C
b111 G
#171920000000
0!
0*
09
0>
0C
#171930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#171940000000
0!
0*
09
0>
0C
#171950000000
1!
1*
b1 6
19
1>
1C
b1 G
#171960000000
0!
0*
09
0>
0C
#171970000000
1!
1*
b10 6
19
1>
1C
b10 G
#171980000000
0!
0*
09
0>
0C
#171990000000
1!
1*
b11 6
19
1>
1C
b11 G
#172000000000
0!
0*
09
0>
0C
#172010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#172020000000
0!
0*
09
0>
0C
#172030000000
1!
1*
b101 6
19
1>
1C
b101 G
#172040000000
0!
0*
09
0>
0C
#172050000000
1!
1*
b110 6
19
1>
1C
b110 G
#172060000000
0!
0*
09
0>
0C
#172070000000
1!
1*
b111 6
19
1>
1C
b111 G
#172080000000
0!
1"
0*
1+
09
1:
0>
0C
#172090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#172100000000
0!
0*
09
0>
0C
#172110000000
1!
1*
b1 6
19
1>
1C
b1 G
#172120000000
0!
0*
09
0>
0C
#172130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#172140000000
0!
0*
09
0>
0C
#172150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#172160000000
0!
0*
09
0>
0C
#172170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#172180000000
0!
0*
09
0>
0C
#172190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#172200000000
0!
0#
0*
0,
09
0>
0?
0C
#172210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#172220000000
0!
0*
09
0>
0C
#172230000000
1!
1*
19
1>
1C
#172240000000
0!
0*
09
0>
0C
#172250000000
1!
1*
19
1>
1C
#172260000000
0!
0*
09
0>
0C
#172270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#172280000000
0!
0*
09
0>
0C
#172290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#172300000000
0!
0*
09
0>
0C
#172310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#172320000000
0!
0*
09
0>
0C
#172330000000
1!
1*
b10 6
19
1>
1C
b10 G
#172340000000
0!
0*
09
0>
0C
#172350000000
1!
1*
b11 6
19
1>
1C
b11 G
#172360000000
0!
0*
09
0>
0C
#172370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#172380000000
0!
0*
09
0>
0C
#172390000000
1!
1*
b101 6
19
1>
1C
b101 G
#172400000000
0!
0*
09
0>
0C
#172410000000
1!
1*
b110 6
19
1>
1C
b110 G
#172420000000
0!
0*
09
0>
0C
#172430000000
1!
1*
b111 6
19
1>
1C
b111 G
#172440000000
0!
0*
09
0>
0C
#172450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#172460000000
0!
0*
09
0>
0C
#172470000000
1!
1*
b1 6
19
1>
1C
b1 G
#172480000000
0!
0*
09
0>
0C
#172490000000
1!
1*
b10 6
19
1>
1C
b10 G
#172500000000
0!
0*
09
0>
0C
#172510000000
1!
1*
b11 6
19
1>
1C
b11 G
#172520000000
0!
0*
09
0>
0C
#172530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#172540000000
0!
0*
09
0>
0C
#172550000000
1!
1*
b101 6
19
1>
1C
b101 G
#172560000000
0!
0*
09
0>
0C
#172570000000
1!
1*
b110 6
19
1>
1C
b110 G
#172580000000
0!
0*
09
0>
0C
#172590000000
1!
1*
b111 6
19
1>
1C
b111 G
#172600000000
0!
0*
09
0>
0C
#172610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#172620000000
0!
0*
09
0>
0C
#172630000000
1!
1*
b1 6
19
1>
1C
b1 G
#172640000000
0!
0*
09
0>
0C
#172650000000
1!
1*
b10 6
19
1>
1C
b10 G
#172660000000
0!
0*
09
0>
0C
#172670000000
1!
1*
b11 6
19
1>
1C
b11 G
#172680000000
0!
0*
09
0>
0C
#172690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#172700000000
0!
0*
09
0>
0C
#172710000000
1!
1*
b101 6
19
1>
1C
b101 G
#172720000000
0!
0*
09
0>
0C
#172730000000
1!
1*
b110 6
19
1>
1C
b110 G
#172740000000
0!
0*
09
0>
0C
#172750000000
1!
1*
b111 6
19
1>
1C
b111 G
#172760000000
0!
1"
0*
1+
09
1:
0>
0C
#172770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#172780000000
0!
0*
09
0>
0C
#172790000000
1!
1*
b1 6
19
1>
1C
b1 G
#172800000000
0!
0*
09
0>
0C
#172810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#172820000000
0!
0*
09
0>
0C
#172830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#172840000000
0!
0*
09
0>
0C
#172850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#172860000000
0!
0*
09
0>
0C
#172870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#172880000000
0!
0#
0*
0,
09
0>
0?
0C
#172890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#172900000000
0!
0*
09
0>
0C
#172910000000
1!
1*
19
1>
1C
#172920000000
0!
0*
09
0>
0C
#172930000000
1!
1*
19
1>
1C
#172940000000
0!
0*
09
0>
0C
#172950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#172960000000
0!
0*
09
0>
0C
#172970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#172980000000
0!
0*
09
0>
0C
#172990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#173000000000
0!
0*
09
0>
0C
#173010000000
1!
1*
b10 6
19
1>
1C
b10 G
#173020000000
0!
0*
09
0>
0C
#173030000000
1!
1*
b11 6
19
1>
1C
b11 G
#173040000000
0!
0*
09
0>
0C
#173050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#173060000000
0!
0*
09
0>
0C
#173070000000
1!
1*
b101 6
19
1>
1C
b101 G
#173080000000
0!
0*
09
0>
0C
#173090000000
1!
1*
b110 6
19
1>
1C
b110 G
#173100000000
0!
0*
09
0>
0C
#173110000000
1!
1*
b111 6
19
1>
1C
b111 G
#173120000000
0!
0*
09
0>
0C
#173130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#173140000000
0!
0*
09
0>
0C
#173150000000
1!
1*
b1 6
19
1>
1C
b1 G
#173160000000
0!
0*
09
0>
0C
#173170000000
1!
1*
b10 6
19
1>
1C
b10 G
#173180000000
0!
0*
09
0>
0C
#173190000000
1!
1*
b11 6
19
1>
1C
b11 G
#173200000000
0!
0*
09
0>
0C
#173210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#173220000000
0!
0*
09
0>
0C
#173230000000
1!
1*
b101 6
19
1>
1C
b101 G
#173240000000
0!
0*
09
0>
0C
#173250000000
1!
1*
b110 6
19
1>
1C
b110 G
#173260000000
0!
0*
09
0>
0C
#173270000000
1!
1*
b111 6
19
1>
1C
b111 G
#173280000000
0!
0*
09
0>
0C
#173290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#173300000000
0!
0*
09
0>
0C
#173310000000
1!
1*
b1 6
19
1>
1C
b1 G
#173320000000
0!
0*
09
0>
0C
#173330000000
1!
1*
b10 6
19
1>
1C
b10 G
#173340000000
0!
0*
09
0>
0C
#173350000000
1!
1*
b11 6
19
1>
1C
b11 G
#173360000000
0!
0*
09
0>
0C
#173370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#173380000000
0!
0*
09
0>
0C
#173390000000
1!
1*
b101 6
19
1>
1C
b101 G
#173400000000
0!
0*
09
0>
0C
#173410000000
1!
1*
b110 6
19
1>
1C
b110 G
#173420000000
0!
0*
09
0>
0C
#173430000000
1!
1*
b111 6
19
1>
1C
b111 G
#173440000000
0!
1"
0*
1+
09
1:
0>
0C
#173450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#173460000000
0!
0*
09
0>
0C
#173470000000
1!
1*
b1 6
19
1>
1C
b1 G
#173480000000
0!
0*
09
0>
0C
#173490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#173500000000
0!
0*
09
0>
0C
#173510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#173520000000
0!
0*
09
0>
0C
#173530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#173540000000
0!
0*
09
0>
0C
#173550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#173560000000
0!
0#
0*
0,
09
0>
0?
0C
#173570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#173580000000
0!
0*
09
0>
0C
#173590000000
1!
1*
19
1>
1C
#173600000000
0!
0*
09
0>
0C
#173610000000
1!
1*
19
1>
1C
#173620000000
0!
0*
09
0>
0C
#173630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#173640000000
0!
0*
09
0>
0C
#173650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#173660000000
0!
0*
09
0>
0C
#173670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#173680000000
0!
0*
09
0>
0C
#173690000000
1!
1*
b10 6
19
1>
1C
b10 G
#173700000000
0!
0*
09
0>
0C
#173710000000
1!
1*
b11 6
19
1>
1C
b11 G
#173720000000
0!
0*
09
0>
0C
#173730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#173740000000
0!
0*
09
0>
0C
#173750000000
1!
1*
b101 6
19
1>
1C
b101 G
#173760000000
0!
0*
09
0>
0C
#173770000000
1!
1*
b110 6
19
1>
1C
b110 G
#173780000000
0!
0*
09
0>
0C
#173790000000
1!
1*
b111 6
19
1>
1C
b111 G
#173800000000
0!
0*
09
0>
0C
#173810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#173820000000
0!
0*
09
0>
0C
#173830000000
1!
1*
b1 6
19
1>
1C
b1 G
#173840000000
0!
0*
09
0>
0C
#173850000000
1!
1*
b10 6
19
1>
1C
b10 G
#173860000000
0!
0*
09
0>
0C
#173870000000
1!
1*
b11 6
19
1>
1C
b11 G
#173880000000
0!
0*
09
0>
0C
#173890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#173900000000
0!
0*
09
0>
0C
#173910000000
1!
1*
b101 6
19
1>
1C
b101 G
#173920000000
0!
0*
09
0>
0C
#173930000000
1!
1*
b110 6
19
1>
1C
b110 G
#173940000000
0!
0*
09
0>
0C
#173950000000
1!
1*
b111 6
19
1>
1C
b111 G
#173960000000
0!
0*
09
0>
0C
#173970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#173980000000
0!
0*
09
0>
0C
#173990000000
1!
1*
b1 6
19
1>
1C
b1 G
#174000000000
0!
0*
09
0>
0C
#174010000000
1!
1*
b10 6
19
1>
1C
b10 G
#174020000000
0!
0*
09
0>
0C
#174030000000
1!
1*
b11 6
19
1>
1C
b11 G
#174040000000
0!
0*
09
0>
0C
#174050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#174060000000
0!
0*
09
0>
0C
#174070000000
1!
1*
b101 6
19
1>
1C
b101 G
#174080000000
0!
0*
09
0>
0C
#174090000000
1!
1*
b110 6
19
1>
1C
b110 G
#174100000000
0!
0*
09
0>
0C
#174110000000
1!
1*
b111 6
19
1>
1C
b111 G
#174120000000
0!
1"
0*
1+
09
1:
0>
0C
#174130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#174140000000
0!
0*
09
0>
0C
#174150000000
1!
1*
b1 6
19
1>
1C
b1 G
#174160000000
0!
0*
09
0>
0C
#174170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#174180000000
0!
0*
09
0>
0C
#174190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#174200000000
0!
0*
09
0>
0C
#174210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#174220000000
0!
0*
09
0>
0C
#174230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#174240000000
0!
0#
0*
0,
09
0>
0?
0C
#174250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#174260000000
0!
0*
09
0>
0C
#174270000000
1!
1*
19
1>
1C
#174280000000
0!
0*
09
0>
0C
#174290000000
1!
1*
19
1>
1C
#174300000000
0!
0*
09
0>
0C
#174310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#174320000000
0!
0*
09
0>
0C
#174330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#174340000000
0!
0*
09
0>
0C
#174350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#174360000000
0!
0*
09
0>
0C
#174370000000
1!
1*
b10 6
19
1>
1C
b10 G
#174380000000
0!
0*
09
0>
0C
#174390000000
1!
1*
b11 6
19
1>
1C
b11 G
#174400000000
0!
0*
09
0>
0C
#174410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#174420000000
0!
0*
09
0>
0C
#174430000000
1!
1*
b101 6
19
1>
1C
b101 G
#174440000000
0!
0*
09
0>
0C
#174450000000
1!
1*
b110 6
19
1>
1C
b110 G
#174460000000
0!
0*
09
0>
0C
#174470000000
1!
1*
b111 6
19
1>
1C
b111 G
#174480000000
0!
0*
09
0>
0C
#174490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#174500000000
0!
0*
09
0>
0C
#174510000000
1!
1*
b1 6
19
1>
1C
b1 G
#174520000000
0!
0*
09
0>
0C
#174530000000
1!
1*
b10 6
19
1>
1C
b10 G
#174540000000
0!
0*
09
0>
0C
#174550000000
1!
1*
b11 6
19
1>
1C
b11 G
#174560000000
0!
0*
09
0>
0C
#174570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#174580000000
0!
0*
09
0>
0C
#174590000000
1!
1*
b101 6
19
1>
1C
b101 G
#174600000000
0!
0*
09
0>
0C
#174610000000
1!
1*
b110 6
19
1>
1C
b110 G
#174620000000
0!
0*
09
0>
0C
#174630000000
1!
1*
b111 6
19
1>
1C
b111 G
#174640000000
0!
0*
09
0>
0C
#174650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#174660000000
0!
0*
09
0>
0C
#174670000000
1!
1*
b1 6
19
1>
1C
b1 G
#174680000000
0!
0*
09
0>
0C
#174690000000
1!
1*
b10 6
19
1>
1C
b10 G
#174700000000
0!
0*
09
0>
0C
#174710000000
1!
1*
b11 6
19
1>
1C
b11 G
#174720000000
0!
0*
09
0>
0C
#174730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#174740000000
0!
0*
09
0>
0C
#174750000000
1!
1*
b101 6
19
1>
1C
b101 G
#174760000000
0!
0*
09
0>
0C
#174770000000
1!
1*
b110 6
19
1>
1C
b110 G
#174780000000
0!
0*
09
0>
0C
#174790000000
1!
1*
b111 6
19
1>
1C
b111 G
#174800000000
0!
1"
0*
1+
09
1:
0>
0C
#174810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#174820000000
0!
0*
09
0>
0C
#174830000000
1!
1*
b1 6
19
1>
1C
b1 G
#174840000000
0!
0*
09
0>
0C
#174850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#174860000000
0!
0*
09
0>
0C
#174870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#174880000000
0!
0*
09
0>
0C
#174890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#174900000000
0!
0*
09
0>
0C
#174910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#174920000000
0!
0#
0*
0,
09
0>
0?
0C
#174930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#174940000000
0!
0*
09
0>
0C
#174950000000
1!
1*
19
1>
1C
#174960000000
0!
0*
09
0>
0C
#174970000000
1!
1*
19
1>
1C
#174980000000
0!
0*
09
0>
0C
#174990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#175000000000
0!
0*
09
0>
0C
#175010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#175020000000
0!
0*
09
0>
0C
#175030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#175040000000
0!
0*
09
0>
0C
#175050000000
1!
1*
b10 6
19
1>
1C
b10 G
#175060000000
0!
0*
09
0>
0C
#175070000000
1!
1*
b11 6
19
1>
1C
b11 G
#175080000000
0!
0*
09
0>
0C
#175090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#175100000000
0!
0*
09
0>
0C
#175110000000
1!
1*
b101 6
19
1>
1C
b101 G
#175120000000
0!
0*
09
0>
0C
#175130000000
1!
1*
b110 6
19
1>
1C
b110 G
#175140000000
0!
0*
09
0>
0C
#175150000000
1!
1*
b111 6
19
1>
1C
b111 G
#175160000000
0!
0*
09
0>
0C
#175170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#175180000000
0!
0*
09
0>
0C
#175190000000
1!
1*
b1 6
19
1>
1C
b1 G
#175200000000
0!
0*
09
0>
0C
#175210000000
1!
1*
b10 6
19
1>
1C
b10 G
#175220000000
0!
0*
09
0>
0C
#175230000000
1!
1*
b11 6
19
1>
1C
b11 G
#175240000000
0!
0*
09
0>
0C
#175250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#175260000000
0!
0*
09
0>
0C
#175270000000
1!
1*
b101 6
19
1>
1C
b101 G
#175280000000
0!
0*
09
0>
0C
#175290000000
1!
1*
b110 6
19
1>
1C
b110 G
#175300000000
0!
0*
09
0>
0C
#175310000000
1!
1*
b111 6
19
1>
1C
b111 G
#175320000000
0!
0*
09
0>
0C
#175330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#175340000000
0!
0*
09
0>
0C
#175350000000
1!
1*
b1 6
19
1>
1C
b1 G
#175360000000
0!
0*
09
0>
0C
#175370000000
1!
1*
b10 6
19
1>
1C
b10 G
#175380000000
0!
0*
09
0>
0C
#175390000000
1!
1*
b11 6
19
1>
1C
b11 G
#175400000000
0!
0*
09
0>
0C
#175410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#175420000000
0!
0*
09
0>
0C
#175430000000
1!
1*
b101 6
19
1>
1C
b101 G
#175440000000
0!
0*
09
0>
0C
#175450000000
1!
1*
b110 6
19
1>
1C
b110 G
#175460000000
0!
0*
09
0>
0C
#175470000000
1!
1*
b111 6
19
1>
1C
b111 G
#175480000000
0!
1"
0*
1+
09
1:
0>
0C
#175490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#175500000000
0!
0*
09
0>
0C
#175510000000
1!
1*
b1 6
19
1>
1C
b1 G
#175520000000
0!
0*
09
0>
0C
#175530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#175540000000
0!
0*
09
0>
0C
#175550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#175560000000
0!
0*
09
0>
0C
#175570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#175580000000
0!
0*
09
0>
0C
#175590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#175600000000
0!
0#
0*
0,
09
0>
0?
0C
#175610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#175620000000
0!
0*
09
0>
0C
#175630000000
1!
1*
19
1>
1C
#175640000000
0!
0*
09
0>
0C
#175650000000
1!
1*
19
1>
1C
#175660000000
0!
0*
09
0>
0C
#175670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#175680000000
0!
0*
09
0>
0C
#175690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#175700000000
0!
0*
09
0>
0C
#175710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#175720000000
0!
0*
09
0>
0C
#175730000000
1!
1*
b10 6
19
1>
1C
b10 G
#175740000000
0!
0*
09
0>
0C
#175750000000
1!
1*
b11 6
19
1>
1C
b11 G
#175760000000
0!
0*
09
0>
0C
#175770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#175780000000
0!
0*
09
0>
0C
#175790000000
1!
1*
b101 6
19
1>
1C
b101 G
#175800000000
0!
0*
09
0>
0C
#175810000000
1!
1*
b110 6
19
1>
1C
b110 G
#175820000000
0!
0*
09
0>
0C
#175830000000
1!
1*
b111 6
19
1>
1C
b111 G
#175840000000
0!
0*
09
0>
0C
#175850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#175860000000
0!
0*
09
0>
0C
#175870000000
1!
1*
b1 6
19
1>
1C
b1 G
#175880000000
0!
0*
09
0>
0C
#175890000000
1!
1*
b10 6
19
1>
1C
b10 G
#175900000000
0!
0*
09
0>
0C
#175910000000
1!
1*
b11 6
19
1>
1C
b11 G
#175920000000
0!
0*
09
0>
0C
#175930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#175940000000
0!
0*
09
0>
0C
#175950000000
1!
1*
b101 6
19
1>
1C
b101 G
#175960000000
0!
0*
09
0>
0C
#175970000000
1!
1*
b110 6
19
1>
1C
b110 G
#175980000000
0!
0*
09
0>
0C
#175990000000
1!
1*
b111 6
19
1>
1C
b111 G
#176000000000
0!
0*
09
0>
0C
#176010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#176020000000
0!
0*
09
0>
0C
#176030000000
1!
1*
b1 6
19
1>
1C
b1 G
#176040000000
0!
0*
09
0>
0C
#176050000000
1!
1*
b10 6
19
1>
1C
b10 G
#176060000000
0!
0*
09
0>
0C
#176070000000
1!
1*
b11 6
19
1>
1C
b11 G
#176080000000
0!
0*
09
0>
0C
#176090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#176100000000
0!
0*
09
0>
0C
#176110000000
1!
1*
b101 6
19
1>
1C
b101 G
#176120000000
0!
0*
09
0>
0C
#176130000000
1!
1*
b110 6
19
1>
1C
b110 G
#176140000000
0!
0*
09
0>
0C
#176150000000
1!
1*
b111 6
19
1>
1C
b111 G
#176160000000
0!
1"
0*
1+
09
1:
0>
0C
#176170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#176180000000
0!
0*
09
0>
0C
#176190000000
1!
1*
b1 6
19
1>
1C
b1 G
#176200000000
0!
0*
09
0>
0C
#176210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#176220000000
0!
0*
09
0>
0C
#176230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#176240000000
0!
0*
09
0>
0C
#176250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#176260000000
0!
0*
09
0>
0C
#176270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#176280000000
0!
0#
0*
0,
09
0>
0?
0C
#176290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#176300000000
0!
0*
09
0>
0C
#176310000000
1!
1*
19
1>
1C
#176320000000
0!
0*
09
0>
0C
#176330000000
1!
1*
19
1>
1C
#176340000000
0!
0*
09
0>
0C
#176350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#176360000000
0!
0*
09
0>
0C
#176370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#176380000000
0!
0*
09
0>
0C
#176390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#176400000000
0!
0*
09
0>
0C
#176410000000
1!
1*
b10 6
19
1>
1C
b10 G
#176420000000
0!
0*
09
0>
0C
#176430000000
1!
1*
b11 6
19
1>
1C
b11 G
#176440000000
0!
0*
09
0>
0C
#176450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#176460000000
0!
0*
09
0>
0C
#176470000000
1!
1*
b101 6
19
1>
1C
b101 G
#176480000000
0!
0*
09
0>
0C
#176490000000
1!
1*
b110 6
19
1>
1C
b110 G
#176500000000
0!
0*
09
0>
0C
#176510000000
1!
1*
b111 6
19
1>
1C
b111 G
#176520000000
0!
0*
09
0>
0C
#176530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#176540000000
0!
0*
09
0>
0C
#176550000000
1!
1*
b1 6
19
1>
1C
b1 G
#176560000000
0!
0*
09
0>
0C
#176570000000
1!
1*
b10 6
19
1>
1C
b10 G
#176580000000
0!
0*
09
0>
0C
#176590000000
1!
1*
b11 6
19
1>
1C
b11 G
#176600000000
0!
0*
09
0>
0C
#176610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#176620000000
0!
0*
09
0>
0C
#176630000000
1!
1*
b101 6
19
1>
1C
b101 G
#176640000000
0!
0*
09
0>
0C
#176650000000
1!
1*
b110 6
19
1>
1C
b110 G
#176660000000
0!
0*
09
0>
0C
#176670000000
1!
1*
b111 6
19
1>
1C
b111 G
#176680000000
0!
0*
09
0>
0C
#176690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#176700000000
0!
0*
09
0>
0C
#176710000000
1!
1*
b1 6
19
1>
1C
b1 G
#176720000000
0!
0*
09
0>
0C
#176730000000
1!
1*
b10 6
19
1>
1C
b10 G
#176740000000
0!
0*
09
0>
0C
#176750000000
1!
1*
b11 6
19
1>
1C
b11 G
#176760000000
0!
0*
09
0>
0C
#176770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#176780000000
0!
0*
09
0>
0C
#176790000000
1!
1*
b101 6
19
1>
1C
b101 G
#176800000000
0!
0*
09
0>
0C
#176810000000
1!
1*
b110 6
19
1>
1C
b110 G
#176820000000
0!
0*
09
0>
0C
#176830000000
1!
1*
b111 6
19
1>
1C
b111 G
#176840000000
0!
1"
0*
1+
09
1:
0>
0C
#176850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#176860000000
0!
0*
09
0>
0C
#176870000000
1!
1*
b1 6
19
1>
1C
b1 G
#176880000000
0!
0*
09
0>
0C
#176890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#176900000000
0!
0*
09
0>
0C
#176910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#176920000000
0!
0*
09
0>
0C
#176930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#176940000000
0!
0*
09
0>
0C
#176950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#176960000000
0!
0#
0*
0,
09
0>
0?
0C
#176970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#176980000000
0!
0*
09
0>
0C
#176990000000
1!
1*
19
1>
1C
#177000000000
0!
0*
09
0>
0C
#177010000000
1!
1*
19
1>
1C
#177020000000
0!
0*
09
0>
0C
#177030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#177040000000
0!
0*
09
0>
0C
#177050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#177060000000
0!
0*
09
0>
0C
#177070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#177080000000
0!
0*
09
0>
0C
#177090000000
1!
1*
b10 6
19
1>
1C
b10 G
#177100000000
0!
0*
09
0>
0C
#177110000000
1!
1*
b11 6
19
1>
1C
b11 G
#177120000000
0!
0*
09
0>
0C
#177130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#177140000000
0!
0*
09
0>
0C
#177150000000
1!
1*
b101 6
19
1>
1C
b101 G
#177160000000
0!
0*
09
0>
0C
#177170000000
1!
1*
b110 6
19
1>
1C
b110 G
#177180000000
0!
0*
09
0>
0C
#177190000000
1!
1*
b111 6
19
1>
1C
b111 G
#177200000000
0!
0*
09
0>
0C
#177210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#177220000000
0!
0*
09
0>
0C
#177230000000
1!
1*
b1 6
19
1>
1C
b1 G
#177240000000
0!
0*
09
0>
0C
#177250000000
1!
1*
b10 6
19
1>
1C
b10 G
#177260000000
0!
0*
09
0>
0C
#177270000000
1!
1*
b11 6
19
1>
1C
b11 G
#177280000000
0!
0*
09
0>
0C
#177290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#177300000000
0!
0*
09
0>
0C
#177310000000
1!
1*
b101 6
19
1>
1C
b101 G
#177320000000
0!
0*
09
0>
0C
#177330000000
1!
1*
b110 6
19
1>
1C
b110 G
#177340000000
0!
0*
09
0>
0C
#177350000000
1!
1*
b111 6
19
1>
1C
b111 G
#177360000000
0!
0*
09
0>
0C
#177370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#177380000000
0!
0*
09
0>
0C
#177390000000
1!
1*
b1 6
19
1>
1C
b1 G
#177400000000
0!
0*
09
0>
0C
#177410000000
1!
1*
b10 6
19
1>
1C
b10 G
#177420000000
0!
0*
09
0>
0C
#177430000000
1!
1*
b11 6
19
1>
1C
b11 G
#177440000000
0!
0*
09
0>
0C
#177450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#177460000000
0!
0*
09
0>
0C
#177470000000
1!
1*
b101 6
19
1>
1C
b101 G
#177480000000
0!
0*
09
0>
0C
#177490000000
1!
1*
b110 6
19
1>
1C
b110 G
#177500000000
0!
0*
09
0>
0C
#177510000000
1!
1*
b111 6
19
1>
1C
b111 G
#177520000000
0!
1"
0*
1+
09
1:
0>
0C
#177530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#177540000000
0!
0*
09
0>
0C
#177550000000
1!
1*
b1 6
19
1>
1C
b1 G
#177560000000
0!
0*
09
0>
0C
#177570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#177580000000
0!
0*
09
0>
0C
#177590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#177600000000
0!
0*
09
0>
0C
#177610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#177620000000
0!
0*
09
0>
0C
#177630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#177640000000
0!
0#
0*
0,
09
0>
0?
0C
#177650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#177660000000
0!
0*
09
0>
0C
#177670000000
1!
1*
19
1>
1C
#177680000000
0!
0*
09
0>
0C
#177690000000
1!
1*
19
1>
1C
#177700000000
0!
0*
09
0>
0C
#177710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#177720000000
0!
0*
09
0>
0C
#177730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#177740000000
0!
0*
09
0>
0C
#177750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#177760000000
0!
0*
09
0>
0C
#177770000000
1!
1*
b10 6
19
1>
1C
b10 G
#177780000000
0!
0*
09
0>
0C
#177790000000
1!
1*
b11 6
19
1>
1C
b11 G
#177800000000
0!
0*
09
0>
0C
#177810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#177820000000
0!
0*
09
0>
0C
#177830000000
1!
1*
b101 6
19
1>
1C
b101 G
#177840000000
0!
0*
09
0>
0C
#177850000000
1!
1*
b110 6
19
1>
1C
b110 G
#177860000000
0!
0*
09
0>
0C
#177870000000
1!
1*
b111 6
19
1>
1C
b111 G
#177880000000
0!
0*
09
0>
0C
#177890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#177900000000
0!
0*
09
0>
0C
#177910000000
1!
1*
b1 6
19
1>
1C
b1 G
#177920000000
0!
0*
09
0>
0C
#177930000000
1!
1*
b10 6
19
1>
1C
b10 G
#177940000000
0!
0*
09
0>
0C
#177950000000
1!
1*
b11 6
19
1>
1C
b11 G
#177960000000
0!
0*
09
0>
0C
#177970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#177980000000
0!
0*
09
0>
0C
#177990000000
1!
1*
b101 6
19
1>
1C
b101 G
#178000000000
0!
0*
09
0>
0C
#178010000000
1!
1*
b110 6
19
1>
1C
b110 G
#178020000000
0!
0*
09
0>
0C
#178030000000
1!
1*
b111 6
19
1>
1C
b111 G
#178040000000
0!
0*
09
0>
0C
#178050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#178060000000
0!
0*
09
0>
0C
#178070000000
1!
1*
b1 6
19
1>
1C
b1 G
#178080000000
0!
0*
09
0>
0C
#178090000000
1!
1*
b10 6
19
1>
1C
b10 G
#178100000000
0!
0*
09
0>
0C
#178110000000
1!
1*
b11 6
19
1>
1C
b11 G
#178120000000
0!
0*
09
0>
0C
#178130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#178140000000
0!
0*
09
0>
0C
#178150000000
1!
1*
b101 6
19
1>
1C
b101 G
#178160000000
0!
0*
09
0>
0C
#178170000000
1!
1*
b110 6
19
1>
1C
b110 G
#178180000000
0!
0*
09
0>
0C
#178190000000
1!
1*
b111 6
19
1>
1C
b111 G
#178200000000
0!
1"
0*
1+
09
1:
0>
0C
#178210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#178220000000
0!
0*
09
0>
0C
#178230000000
1!
1*
b1 6
19
1>
1C
b1 G
#178240000000
0!
0*
09
0>
0C
#178250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#178260000000
0!
0*
09
0>
0C
#178270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#178280000000
0!
0*
09
0>
0C
#178290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#178300000000
0!
0*
09
0>
0C
#178310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#178320000000
0!
0#
0*
0,
09
0>
0?
0C
#178330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#178340000000
0!
0*
09
0>
0C
#178350000000
1!
1*
19
1>
1C
#178360000000
0!
0*
09
0>
0C
#178370000000
1!
1*
19
1>
1C
#178380000000
0!
0*
09
0>
0C
#178390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#178400000000
0!
0*
09
0>
0C
#178410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#178420000000
0!
0*
09
0>
0C
#178430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#178440000000
0!
0*
09
0>
0C
#178450000000
1!
1*
b10 6
19
1>
1C
b10 G
#178460000000
0!
0*
09
0>
0C
#178470000000
1!
1*
b11 6
19
1>
1C
b11 G
#178480000000
0!
0*
09
0>
0C
#178490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#178500000000
0!
0*
09
0>
0C
#178510000000
1!
1*
b101 6
19
1>
1C
b101 G
#178520000000
0!
0*
09
0>
0C
#178530000000
1!
1*
b110 6
19
1>
1C
b110 G
#178540000000
0!
0*
09
0>
0C
#178550000000
1!
1*
b111 6
19
1>
1C
b111 G
#178560000000
0!
0*
09
0>
0C
#178570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#178580000000
0!
0*
09
0>
0C
#178590000000
1!
1*
b1 6
19
1>
1C
b1 G
#178600000000
0!
0*
09
0>
0C
#178610000000
1!
1*
b10 6
19
1>
1C
b10 G
#178620000000
0!
0*
09
0>
0C
#178630000000
1!
1*
b11 6
19
1>
1C
b11 G
#178640000000
0!
0*
09
0>
0C
#178650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#178660000000
0!
0*
09
0>
0C
#178670000000
1!
1*
b101 6
19
1>
1C
b101 G
#178680000000
0!
0*
09
0>
0C
#178690000000
1!
1*
b110 6
19
1>
1C
b110 G
#178700000000
0!
0*
09
0>
0C
#178710000000
1!
1*
b111 6
19
1>
1C
b111 G
#178720000000
0!
0*
09
0>
0C
#178730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#178740000000
0!
0*
09
0>
0C
#178750000000
1!
1*
b1 6
19
1>
1C
b1 G
#178760000000
0!
0*
09
0>
0C
#178770000000
1!
1*
b10 6
19
1>
1C
b10 G
#178780000000
0!
0*
09
0>
0C
#178790000000
1!
1*
b11 6
19
1>
1C
b11 G
#178800000000
0!
0*
09
0>
0C
#178810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#178820000000
0!
0*
09
0>
0C
#178830000000
1!
1*
b101 6
19
1>
1C
b101 G
#178840000000
0!
0*
09
0>
0C
#178850000000
1!
1*
b110 6
19
1>
1C
b110 G
#178860000000
0!
0*
09
0>
0C
#178870000000
1!
1*
b111 6
19
1>
1C
b111 G
#178880000000
0!
1"
0*
1+
09
1:
0>
0C
#178890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#178900000000
0!
0*
09
0>
0C
#178910000000
1!
1*
b1 6
19
1>
1C
b1 G
#178920000000
0!
0*
09
0>
0C
#178930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#178940000000
0!
0*
09
0>
0C
#178950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#178960000000
0!
0*
09
0>
0C
#178970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#178980000000
0!
0*
09
0>
0C
#178990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#179000000000
0!
0#
0*
0,
09
0>
0?
0C
#179010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#179020000000
0!
0*
09
0>
0C
#179030000000
1!
1*
19
1>
1C
#179040000000
0!
0*
09
0>
0C
#179050000000
1!
1*
19
1>
1C
#179060000000
0!
0*
09
0>
0C
#179070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#179080000000
0!
0*
09
0>
0C
#179090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#179100000000
0!
0*
09
0>
0C
#179110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#179120000000
0!
0*
09
0>
0C
#179130000000
1!
1*
b10 6
19
1>
1C
b10 G
#179140000000
0!
0*
09
0>
0C
#179150000000
1!
1*
b11 6
19
1>
1C
b11 G
#179160000000
0!
0*
09
0>
0C
#179170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#179180000000
0!
0*
09
0>
0C
#179190000000
1!
1*
b101 6
19
1>
1C
b101 G
#179200000000
0!
0*
09
0>
0C
#179210000000
1!
1*
b110 6
19
1>
1C
b110 G
#179220000000
0!
0*
09
0>
0C
#179230000000
1!
1*
b111 6
19
1>
1C
b111 G
#179240000000
0!
0*
09
0>
0C
#179250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#179260000000
0!
0*
09
0>
0C
#179270000000
1!
1*
b1 6
19
1>
1C
b1 G
#179280000000
0!
0*
09
0>
0C
#179290000000
1!
1*
b10 6
19
1>
1C
b10 G
#179300000000
0!
0*
09
0>
0C
#179310000000
1!
1*
b11 6
19
1>
1C
b11 G
#179320000000
0!
0*
09
0>
0C
#179330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#179340000000
0!
0*
09
0>
0C
#179350000000
1!
1*
b101 6
19
1>
1C
b101 G
#179360000000
0!
0*
09
0>
0C
#179370000000
1!
1*
b110 6
19
1>
1C
b110 G
#179380000000
0!
0*
09
0>
0C
#179390000000
1!
1*
b111 6
19
1>
1C
b111 G
#179400000000
0!
0*
09
0>
0C
#179410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#179420000000
0!
0*
09
0>
0C
#179430000000
1!
1*
b1 6
19
1>
1C
b1 G
#179440000000
0!
0*
09
0>
0C
#179450000000
1!
1*
b10 6
19
1>
1C
b10 G
#179460000000
0!
0*
09
0>
0C
#179470000000
1!
1*
b11 6
19
1>
1C
b11 G
#179480000000
0!
0*
09
0>
0C
#179490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#179500000000
0!
0*
09
0>
0C
#179510000000
1!
1*
b101 6
19
1>
1C
b101 G
#179520000000
0!
0*
09
0>
0C
#179530000000
1!
1*
b110 6
19
1>
1C
b110 G
#179540000000
0!
0*
09
0>
0C
#179550000000
1!
1*
b111 6
19
1>
1C
b111 G
#179560000000
0!
1"
0*
1+
09
1:
0>
0C
#179570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#179580000000
0!
0*
09
0>
0C
#179590000000
1!
1*
b1 6
19
1>
1C
b1 G
#179600000000
0!
0*
09
0>
0C
#179610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#179620000000
0!
0*
09
0>
0C
#179630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#179640000000
0!
0*
09
0>
0C
#179650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#179660000000
0!
0*
09
0>
0C
#179670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#179680000000
0!
0#
0*
0,
09
0>
0?
0C
#179690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#179700000000
0!
0*
09
0>
0C
#179710000000
1!
1*
19
1>
1C
#179720000000
0!
0*
09
0>
0C
#179730000000
1!
1*
19
1>
1C
#179740000000
0!
0*
09
0>
0C
#179750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#179760000000
0!
0*
09
0>
0C
#179770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#179780000000
0!
0*
09
0>
0C
#179790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#179800000000
0!
0*
09
0>
0C
#179810000000
1!
1*
b10 6
19
1>
1C
b10 G
#179820000000
0!
0*
09
0>
0C
#179830000000
1!
1*
b11 6
19
1>
1C
b11 G
#179840000000
0!
0*
09
0>
0C
#179850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#179860000000
0!
0*
09
0>
0C
#179870000000
1!
1*
b101 6
19
1>
1C
b101 G
#179880000000
0!
0*
09
0>
0C
#179890000000
1!
1*
b110 6
19
1>
1C
b110 G
#179900000000
0!
0*
09
0>
0C
#179910000000
1!
1*
b111 6
19
1>
1C
b111 G
#179920000000
0!
0*
09
0>
0C
#179930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#179940000000
0!
0*
09
0>
0C
#179950000000
1!
1*
b1 6
19
1>
1C
b1 G
#179960000000
0!
0*
09
0>
0C
#179970000000
1!
1*
b10 6
19
1>
1C
b10 G
#179980000000
0!
0*
09
0>
0C
#179990000000
1!
1*
b11 6
19
1>
1C
b11 G
#180000000000
0!
0*
09
0>
0C
#180010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#180020000000
0!
0*
09
0>
0C
#180030000000
1!
1*
b101 6
19
1>
1C
b101 G
#180040000000
0!
0*
09
0>
0C
#180050000000
1!
1*
b110 6
19
1>
1C
b110 G
#180060000000
0!
0*
09
0>
0C
#180070000000
1!
1*
b111 6
19
1>
1C
b111 G
#180080000000
0!
0*
09
0>
0C
#180090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#180100000000
0!
0*
09
0>
0C
#180110000000
1!
1*
b1 6
19
1>
1C
b1 G
#180120000000
0!
0*
09
0>
0C
#180130000000
1!
1*
b10 6
19
1>
1C
b10 G
#180140000000
0!
0*
09
0>
0C
#180150000000
1!
1*
b11 6
19
1>
1C
b11 G
#180160000000
0!
0*
09
0>
0C
#180170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#180180000000
0!
0*
09
0>
0C
#180190000000
1!
1*
b101 6
19
1>
1C
b101 G
#180200000000
0!
0*
09
0>
0C
#180210000000
1!
1*
b110 6
19
1>
1C
b110 G
#180220000000
0!
0*
09
0>
0C
#180230000000
1!
1*
b111 6
19
1>
1C
b111 G
#180240000000
0!
1"
0*
1+
09
1:
0>
0C
#180250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#180260000000
0!
0*
09
0>
0C
#180270000000
1!
1*
b1 6
19
1>
1C
b1 G
#180280000000
0!
0*
09
0>
0C
#180290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#180300000000
0!
0*
09
0>
0C
#180310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#180320000000
0!
0*
09
0>
0C
#180330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#180340000000
0!
0*
09
0>
0C
#180350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#180360000000
0!
0#
0*
0,
09
0>
0?
0C
#180370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#180380000000
0!
0*
09
0>
0C
#180390000000
1!
1*
19
1>
1C
#180400000000
0!
0*
09
0>
0C
#180410000000
1!
1*
19
1>
1C
#180420000000
0!
0*
09
0>
0C
#180430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#180440000000
0!
0*
09
0>
0C
#180450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#180460000000
0!
0*
09
0>
0C
#180470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#180480000000
0!
0*
09
0>
0C
#180490000000
1!
1*
b10 6
19
1>
1C
b10 G
#180500000000
0!
0*
09
0>
0C
#180510000000
1!
1*
b11 6
19
1>
1C
b11 G
#180520000000
0!
0*
09
0>
0C
#180530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#180540000000
0!
0*
09
0>
0C
#180550000000
1!
1*
b101 6
19
1>
1C
b101 G
#180560000000
0!
0*
09
0>
0C
#180570000000
1!
1*
b110 6
19
1>
1C
b110 G
#180580000000
0!
0*
09
0>
0C
#180590000000
1!
1*
b111 6
19
1>
1C
b111 G
#180600000000
0!
0*
09
0>
0C
#180610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#180620000000
0!
0*
09
0>
0C
#180630000000
1!
1*
b1 6
19
1>
1C
b1 G
#180640000000
0!
0*
09
0>
0C
#180650000000
1!
1*
b10 6
19
1>
1C
b10 G
#180660000000
0!
0*
09
0>
0C
#180670000000
1!
1*
b11 6
19
1>
1C
b11 G
#180680000000
0!
0*
09
0>
0C
#180690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#180700000000
0!
0*
09
0>
0C
#180710000000
1!
1*
b101 6
19
1>
1C
b101 G
#180720000000
0!
0*
09
0>
0C
#180730000000
1!
1*
b110 6
19
1>
1C
b110 G
#180740000000
0!
0*
09
0>
0C
#180750000000
1!
1*
b111 6
19
1>
1C
b111 G
#180760000000
0!
0*
09
0>
0C
#180770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#180780000000
0!
0*
09
0>
0C
#180790000000
1!
1*
b1 6
19
1>
1C
b1 G
#180800000000
0!
0*
09
0>
0C
#180810000000
1!
1*
b10 6
19
1>
1C
b10 G
#180820000000
0!
0*
09
0>
0C
#180830000000
1!
1*
b11 6
19
1>
1C
b11 G
#180840000000
0!
0*
09
0>
0C
#180850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#180860000000
0!
0*
09
0>
0C
#180870000000
1!
1*
b101 6
19
1>
1C
b101 G
#180880000000
0!
0*
09
0>
0C
#180890000000
1!
1*
b110 6
19
1>
1C
b110 G
#180900000000
0!
0*
09
0>
0C
#180910000000
1!
1*
b111 6
19
1>
1C
b111 G
#180920000000
0!
1"
0*
1+
09
1:
0>
0C
#180930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#180940000000
0!
0*
09
0>
0C
#180950000000
1!
1*
b1 6
19
1>
1C
b1 G
#180960000000
0!
0*
09
0>
0C
#180970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#180980000000
0!
0*
09
0>
0C
#180990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#181000000000
0!
0*
09
0>
0C
#181010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#181020000000
0!
0*
09
0>
0C
#181030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#181040000000
0!
0#
0*
0,
09
0>
0?
0C
#181050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#181060000000
0!
0*
09
0>
0C
#181070000000
1!
1*
19
1>
1C
#181080000000
0!
0*
09
0>
0C
#181090000000
1!
1*
19
1>
1C
#181100000000
0!
0*
09
0>
0C
#181110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#181120000000
0!
0*
09
0>
0C
#181130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#181140000000
0!
0*
09
0>
0C
#181150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#181160000000
0!
0*
09
0>
0C
#181170000000
1!
1*
b10 6
19
1>
1C
b10 G
#181180000000
0!
0*
09
0>
0C
#181190000000
1!
1*
b11 6
19
1>
1C
b11 G
#181200000000
0!
0*
09
0>
0C
#181210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#181220000000
0!
0*
09
0>
0C
#181230000000
1!
1*
b101 6
19
1>
1C
b101 G
#181240000000
0!
0*
09
0>
0C
#181250000000
1!
1*
b110 6
19
1>
1C
b110 G
#181260000000
0!
0*
09
0>
0C
#181270000000
1!
1*
b111 6
19
1>
1C
b111 G
#181280000000
0!
0*
09
0>
0C
#181290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#181300000000
0!
0*
09
0>
0C
#181310000000
1!
1*
b1 6
19
1>
1C
b1 G
#181320000000
0!
0*
09
0>
0C
#181330000000
1!
1*
b10 6
19
1>
1C
b10 G
#181340000000
0!
0*
09
0>
0C
#181350000000
1!
1*
b11 6
19
1>
1C
b11 G
#181360000000
0!
0*
09
0>
0C
#181370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#181380000000
0!
0*
09
0>
0C
#181390000000
1!
1*
b101 6
19
1>
1C
b101 G
#181400000000
0!
0*
09
0>
0C
#181410000000
1!
1*
b110 6
19
1>
1C
b110 G
#181420000000
0!
0*
09
0>
0C
#181430000000
1!
1*
b111 6
19
1>
1C
b111 G
#181440000000
0!
0*
09
0>
0C
#181450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#181460000000
0!
0*
09
0>
0C
#181470000000
1!
1*
b1 6
19
1>
1C
b1 G
#181480000000
0!
0*
09
0>
0C
#181490000000
1!
1*
b10 6
19
1>
1C
b10 G
#181500000000
0!
0*
09
0>
0C
#181510000000
1!
1*
b11 6
19
1>
1C
b11 G
#181520000000
0!
0*
09
0>
0C
#181530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#181540000000
0!
0*
09
0>
0C
#181550000000
1!
1*
b101 6
19
1>
1C
b101 G
#181560000000
0!
0*
09
0>
0C
#181570000000
1!
1*
b110 6
19
1>
1C
b110 G
#181580000000
0!
0*
09
0>
0C
#181590000000
1!
1*
b111 6
19
1>
1C
b111 G
#181600000000
0!
1"
0*
1+
09
1:
0>
0C
#181610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#181620000000
0!
0*
09
0>
0C
#181630000000
1!
1*
b1 6
19
1>
1C
b1 G
#181640000000
0!
0*
09
0>
0C
#181650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#181660000000
0!
0*
09
0>
0C
#181670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#181680000000
0!
0*
09
0>
0C
#181690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#181700000000
0!
0*
09
0>
0C
#181710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#181720000000
0!
0#
0*
0,
09
0>
0?
0C
#181730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#181740000000
0!
0*
09
0>
0C
#181750000000
1!
1*
19
1>
1C
#181760000000
0!
0*
09
0>
0C
#181770000000
1!
1*
19
1>
1C
#181780000000
0!
0*
09
0>
0C
#181790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#181800000000
0!
0*
09
0>
0C
#181810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#181820000000
0!
0*
09
0>
0C
#181830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#181840000000
0!
0*
09
0>
0C
#181850000000
1!
1*
b10 6
19
1>
1C
b10 G
#181860000000
0!
0*
09
0>
0C
#181870000000
1!
1*
b11 6
19
1>
1C
b11 G
#181880000000
0!
0*
09
0>
0C
#181890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#181900000000
0!
0*
09
0>
0C
#181910000000
1!
1*
b101 6
19
1>
1C
b101 G
#181920000000
0!
0*
09
0>
0C
#181930000000
1!
1*
b110 6
19
1>
1C
b110 G
#181940000000
0!
0*
09
0>
0C
#181950000000
1!
1*
b111 6
19
1>
1C
b111 G
#181960000000
0!
0*
09
0>
0C
#181970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#181980000000
0!
0*
09
0>
0C
#181990000000
1!
1*
b1 6
19
1>
1C
b1 G
#182000000000
0!
0*
09
0>
0C
#182010000000
1!
1*
b10 6
19
1>
1C
b10 G
#182020000000
0!
0*
09
0>
0C
#182030000000
1!
1*
b11 6
19
1>
1C
b11 G
#182040000000
0!
0*
09
0>
0C
#182050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#182060000000
0!
0*
09
0>
0C
#182070000000
1!
1*
b101 6
19
1>
1C
b101 G
#182080000000
0!
0*
09
0>
0C
#182090000000
1!
1*
b110 6
19
1>
1C
b110 G
#182100000000
0!
0*
09
0>
0C
#182110000000
1!
1*
b111 6
19
1>
1C
b111 G
#182120000000
0!
0*
09
0>
0C
#182130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#182140000000
0!
0*
09
0>
0C
#182150000000
1!
1*
b1 6
19
1>
1C
b1 G
#182160000000
0!
0*
09
0>
0C
#182170000000
1!
1*
b10 6
19
1>
1C
b10 G
#182180000000
0!
0*
09
0>
0C
#182190000000
1!
1*
b11 6
19
1>
1C
b11 G
#182200000000
0!
0*
09
0>
0C
#182210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#182220000000
0!
0*
09
0>
0C
#182230000000
1!
1*
b101 6
19
1>
1C
b101 G
#182240000000
0!
0*
09
0>
0C
#182250000000
1!
1*
b110 6
19
1>
1C
b110 G
#182260000000
0!
0*
09
0>
0C
#182270000000
1!
1*
b111 6
19
1>
1C
b111 G
#182280000000
0!
1"
0*
1+
09
1:
0>
0C
#182290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#182300000000
0!
0*
09
0>
0C
#182310000000
1!
1*
b1 6
19
1>
1C
b1 G
#182320000000
0!
0*
09
0>
0C
#182330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#182340000000
0!
0*
09
0>
0C
#182350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#182360000000
0!
0*
09
0>
0C
#182370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#182380000000
0!
0*
09
0>
0C
#182390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#182400000000
0!
0#
0*
0,
09
0>
0?
0C
#182410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#182420000000
0!
0*
09
0>
0C
#182430000000
1!
1*
19
1>
1C
#182440000000
0!
0*
09
0>
0C
#182450000000
1!
1*
19
1>
1C
#182460000000
0!
0*
09
0>
0C
#182470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#182480000000
0!
0*
09
0>
0C
#182490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#182500000000
0!
0*
09
0>
0C
#182510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#182520000000
0!
0*
09
0>
0C
#182530000000
1!
1*
b10 6
19
1>
1C
b10 G
#182540000000
0!
0*
09
0>
0C
#182550000000
1!
1*
b11 6
19
1>
1C
b11 G
#182560000000
0!
0*
09
0>
0C
#182570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#182580000000
0!
0*
09
0>
0C
#182590000000
1!
1*
b101 6
19
1>
1C
b101 G
#182600000000
0!
0*
09
0>
0C
#182610000000
1!
1*
b110 6
19
1>
1C
b110 G
#182620000000
0!
0*
09
0>
0C
#182630000000
1!
1*
b111 6
19
1>
1C
b111 G
#182640000000
0!
0*
09
0>
0C
#182650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#182660000000
0!
0*
09
0>
0C
#182670000000
1!
1*
b1 6
19
1>
1C
b1 G
#182680000000
0!
0*
09
0>
0C
#182690000000
1!
1*
b10 6
19
1>
1C
b10 G
#182700000000
0!
0*
09
0>
0C
#182710000000
1!
1*
b11 6
19
1>
1C
b11 G
#182720000000
0!
0*
09
0>
0C
#182730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#182740000000
0!
0*
09
0>
0C
#182750000000
1!
1*
b101 6
19
1>
1C
b101 G
#182760000000
0!
0*
09
0>
0C
#182770000000
1!
1*
b110 6
19
1>
1C
b110 G
#182780000000
0!
0*
09
0>
0C
#182790000000
1!
1*
b111 6
19
1>
1C
b111 G
#182800000000
0!
0*
09
0>
0C
#182810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#182820000000
0!
0*
09
0>
0C
#182830000000
1!
1*
b1 6
19
1>
1C
b1 G
#182840000000
0!
0*
09
0>
0C
#182850000000
1!
1*
b10 6
19
1>
1C
b10 G
#182860000000
0!
0*
09
0>
0C
#182870000000
1!
1*
b11 6
19
1>
1C
b11 G
#182880000000
0!
0*
09
0>
0C
#182890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#182900000000
0!
0*
09
0>
0C
#182910000000
1!
1*
b101 6
19
1>
1C
b101 G
#182920000000
0!
0*
09
0>
0C
#182930000000
1!
1*
b110 6
19
1>
1C
b110 G
#182940000000
0!
0*
09
0>
0C
#182950000000
1!
1*
b111 6
19
1>
1C
b111 G
#182960000000
0!
1"
0*
1+
09
1:
0>
0C
#182970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#182980000000
0!
0*
09
0>
0C
#182990000000
1!
1*
b1 6
19
1>
1C
b1 G
#183000000000
0!
0*
09
0>
0C
#183010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#183020000000
0!
0*
09
0>
0C
#183030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#183040000000
0!
0*
09
0>
0C
#183050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#183060000000
0!
0*
09
0>
0C
#183070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#183080000000
0!
0#
0*
0,
09
0>
0?
0C
#183090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#183100000000
0!
0*
09
0>
0C
#183110000000
1!
1*
19
1>
1C
#183120000000
0!
0*
09
0>
0C
#183130000000
1!
1*
19
1>
1C
#183140000000
0!
0*
09
0>
0C
#183150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#183160000000
0!
0*
09
0>
0C
#183170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#183180000000
0!
0*
09
0>
0C
#183190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#183200000000
0!
0*
09
0>
0C
#183210000000
1!
1*
b10 6
19
1>
1C
b10 G
#183220000000
0!
0*
09
0>
0C
#183230000000
1!
1*
b11 6
19
1>
1C
b11 G
#183240000000
0!
0*
09
0>
0C
#183250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#183260000000
0!
0*
09
0>
0C
#183270000000
1!
1*
b101 6
19
1>
1C
b101 G
#183280000000
0!
0*
09
0>
0C
#183290000000
1!
1*
b110 6
19
1>
1C
b110 G
#183300000000
0!
0*
09
0>
0C
#183310000000
1!
1*
b111 6
19
1>
1C
b111 G
#183320000000
0!
0*
09
0>
0C
#183330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#183340000000
0!
0*
09
0>
0C
#183350000000
1!
1*
b1 6
19
1>
1C
b1 G
#183360000000
0!
0*
09
0>
0C
#183370000000
1!
1*
b10 6
19
1>
1C
b10 G
#183380000000
0!
0*
09
0>
0C
#183390000000
1!
1*
b11 6
19
1>
1C
b11 G
#183400000000
0!
0*
09
0>
0C
#183410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#183420000000
0!
0*
09
0>
0C
#183430000000
1!
1*
b101 6
19
1>
1C
b101 G
#183440000000
0!
0*
09
0>
0C
#183450000000
1!
1*
b110 6
19
1>
1C
b110 G
#183460000000
0!
0*
09
0>
0C
#183470000000
1!
1*
b111 6
19
1>
1C
b111 G
#183480000000
0!
0*
09
0>
0C
#183490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#183500000000
0!
0*
09
0>
0C
#183510000000
1!
1*
b1 6
19
1>
1C
b1 G
#183520000000
0!
0*
09
0>
0C
#183530000000
1!
1*
b10 6
19
1>
1C
b10 G
#183540000000
0!
0*
09
0>
0C
#183550000000
1!
1*
b11 6
19
1>
1C
b11 G
#183560000000
0!
0*
09
0>
0C
#183570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#183580000000
0!
0*
09
0>
0C
#183590000000
1!
1*
b101 6
19
1>
1C
b101 G
#183600000000
0!
0*
09
0>
0C
#183610000000
1!
1*
b110 6
19
1>
1C
b110 G
#183620000000
0!
0*
09
0>
0C
#183630000000
1!
1*
b111 6
19
1>
1C
b111 G
#183640000000
0!
1"
0*
1+
09
1:
0>
0C
#183650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#183660000000
0!
0*
09
0>
0C
#183670000000
1!
1*
b1 6
19
1>
1C
b1 G
#183680000000
0!
0*
09
0>
0C
#183690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#183700000000
0!
0*
09
0>
0C
#183710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#183720000000
0!
0*
09
0>
0C
#183730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#183740000000
0!
0*
09
0>
0C
#183750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#183760000000
0!
0#
0*
0,
09
0>
0?
0C
#183770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#183780000000
0!
0*
09
0>
0C
#183790000000
1!
1*
19
1>
1C
#183800000000
0!
0*
09
0>
0C
#183810000000
1!
1*
19
1>
1C
#183820000000
0!
0*
09
0>
0C
#183830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#183840000000
0!
0*
09
0>
0C
#183850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#183860000000
0!
0*
09
0>
0C
#183870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#183880000000
0!
0*
09
0>
0C
#183890000000
1!
1*
b10 6
19
1>
1C
b10 G
#183900000000
0!
0*
09
0>
0C
#183910000000
1!
1*
b11 6
19
1>
1C
b11 G
#183920000000
0!
0*
09
0>
0C
#183930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#183940000000
0!
0*
09
0>
0C
#183950000000
1!
1*
b101 6
19
1>
1C
b101 G
#183960000000
0!
0*
09
0>
0C
#183970000000
1!
1*
b110 6
19
1>
1C
b110 G
#183980000000
0!
0*
09
0>
0C
#183990000000
1!
1*
b111 6
19
1>
1C
b111 G
#184000000000
0!
0*
09
0>
0C
#184010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#184020000000
0!
0*
09
0>
0C
#184030000000
1!
1*
b1 6
19
1>
1C
b1 G
#184040000000
0!
0*
09
0>
0C
#184050000000
1!
1*
b10 6
19
1>
1C
b10 G
#184060000000
0!
0*
09
0>
0C
#184070000000
1!
1*
b11 6
19
1>
1C
b11 G
#184080000000
0!
0*
09
0>
0C
#184090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#184100000000
0!
0*
09
0>
0C
#184110000000
1!
1*
b101 6
19
1>
1C
b101 G
#184120000000
0!
0*
09
0>
0C
#184130000000
1!
1*
b110 6
19
1>
1C
b110 G
#184140000000
0!
0*
09
0>
0C
#184150000000
1!
1*
b111 6
19
1>
1C
b111 G
#184160000000
0!
0*
09
0>
0C
#184170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#184180000000
0!
0*
09
0>
0C
#184190000000
1!
1*
b1 6
19
1>
1C
b1 G
#184200000000
0!
0*
09
0>
0C
#184210000000
1!
1*
b10 6
19
1>
1C
b10 G
#184220000000
0!
0*
09
0>
0C
#184230000000
1!
1*
b11 6
19
1>
1C
b11 G
#184240000000
0!
0*
09
0>
0C
#184250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#184260000000
0!
0*
09
0>
0C
#184270000000
1!
1*
b101 6
19
1>
1C
b101 G
#184280000000
0!
0*
09
0>
0C
#184290000000
1!
1*
b110 6
19
1>
1C
b110 G
#184300000000
0!
0*
09
0>
0C
#184310000000
1!
1*
b111 6
19
1>
1C
b111 G
#184320000000
0!
1"
0*
1+
09
1:
0>
0C
#184330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#184340000000
0!
0*
09
0>
0C
#184350000000
1!
1*
b1 6
19
1>
1C
b1 G
#184360000000
0!
0*
09
0>
0C
#184370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#184380000000
0!
0*
09
0>
0C
#184390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#184400000000
0!
0*
09
0>
0C
#184410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#184420000000
0!
0*
09
0>
0C
#184430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#184440000000
0!
0#
0*
0,
09
0>
0?
0C
#184450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#184460000000
0!
0*
09
0>
0C
#184470000000
1!
1*
19
1>
1C
#184480000000
0!
0*
09
0>
0C
#184490000000
1!
1*
19
1>
1C
#184500000000
0!
0*
09
0>
0C
#184510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#184520000000
0!
0*
09
0>
0C
#184530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#184540000000
0!
0*
09
0>
0C
#184550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#184560000000
0!
0*
09
0>
0C
#184570000000
1!
1*
b10 6
19
1>
1C
b10 G
#184580000000
0!
0*
09
0>
0C
#184590000000
1!
1*
b11 6
19
1>
1C
b11 G
#184600000000
0!
0*
09
0>
0C
#184610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#184620000000
0!
0*
09
0>
0C
#184630000000
1!
1*
b101 6
19
1>
1C
b101 G
#184640000000
0!
0*
09
0>
0C
#184650000000
1!
1*
b110 6
19
1>
1C
b110 G
#184660000000
0!
0*
09
0>
0C
#184670000000
1!
1*
b111 6
19
1>
1C
b111 G
#184680000000
0!
0*
09
0>
0C
#184690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#184700000000
0!
0*
09
0>
0C
#184710000000
1!
1*
b1 6
19
1>
1C
b1 G
#184720000000
0!
0*
09
0>
0C
#184730000000
1!
1*
b10 6
19
1>
1C
b10 G
#184740000000
0!
0*
09
0>
0C
#184750000000
1!
1*
b11 6
19
1>
1C
b11 G
#184760000000
0!
0*
09
0>
0C
#184770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#184780000000
0!
0*
09
0>
0C
#184790000000
1!
1*
b101 6
19
1>
1C
b101 G
#184800000000
0!
0*
09
0>
0C
#184810000000
1!
1*
b110 6
19
1>
1C
b110 G
#184820000000
0!
0*
09
0>
0C
#184830000000
1!
1*
b111 6
19
1>
1C
b111 G
#184840000000
0!
0*
09
0>
0C
#184850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#184860000000
0!
0*
09
0>
0C
#184870000000
1!
1*
b1 6
19
1>
1C
b1 G
#184880000000
0!
0*
09
0>
0C
#184890000000
1!
1*
b10 6
19
1>
1C
b10 G
#184900000000
0!
0*
09
0>
0C
#184910000000
1!
1*
b11 6
19
1>
1C
b11 G
#184920000000
0!
0*
09
0>
0C
#184930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#184940000000
0!
0*
09
0>
0C
#184950000000
1!
1*
b101 6
19
1>
1C
b101 G
#184960000000
0!
0*
09
0>
0C
#184970000000
1!
1*
b110 6
19
1>
1C
b110 G
#184980000000
0!
0*
09
0>
0C
#184990000000
1!
1*
b111 6
19
1>
1C
b111 G
#185000000000
0!
1"
0*
1+
09
1:
0>
0C
#185010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#185020000000
0!
0*
09
0>
0C
#185030000000
1!
1*
b1 6
19
1>
1C
b1 G
#185040000000
0!
0*
09
0>
0C
#185050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#185060000000
0!
0*
09
0>
0C
#185070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#185080000000
0!
0*
09
0>
0C
#185090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#185100000000
0!
0*
09
0>
0C
#185110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#185120000000
0!
0#
0*
0,
09
0>
0?
0C
#185130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#185140000000
0!
0*
09
0>
0C
#185150000000
1!
1*
19
1>
1C
#185160000000
0!
0*
09
0>
0C
#185170000000
1!
1*
19
1>
1C
#185180000000
0!
0*
09
0>
0C
#185190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#185200000000
0!
0*
09
0>
0C
#185210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#185220000000
0!
0*
09
0>
0C
#185230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#185240000000
0!
0*
09
0>
0C
#185250000000
1!
1*
b10 6
19
1>
1C
b10 G
#185260000000
0!
0*
09
0>
0C
#185270000000
1!
1*
b11 6
19
1>
1C
b11 G
#185280000000
0!
0*
09
0>
0C
#185290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#185300000000
0!
0*
09
0>
0C
#185310000000
1!
1*
b101 6
19
1>
1C
b101 G
#185320000000
0!
0*
09
0>
0C
#185330000000
1!
1*
b110 6
19
1>
1C
b110 G
#185340000000
0!
0*
09
0>
0C
#185350000000
1!
1*
b111 6
19
1>
1C
b111 G
#185360000000
0!
0*
09
0>
0C
#185370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#185380000000
0!
0*
09
0>
0C
#185390000000
1!
1*
b1 6
19
1>
1C
b1 G
#185400000000
0!
0*
09
0>
0C
#185410000000
1!
1*
b10 6
19
1>
1C
b10 G
#185420000000
0!
0*
09
0>
0C
#185430000000
1!
1*
b11 6
19
1>
1C
b11 G
#185440000000
0!
0*
09
0>
0C
#185450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#185460000000
0!
0*
09
0>
0C
#185470000000
1!
1*
b101 6
19
1>
1C
b101 G
#185480000000
0!
0*
09
0>
0C
#185490000000
1!
1*
b110 6
19
1>
1C
b110 G
#185500000000
0!
0*
09
0>
0C
#185510000000
1!
1*
b111 6
19
1>
1C
b111 G
#185520000000
0!
0*
09
0>
0C
#185530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#185540000000
0!
0*
09
0>
0C
#185550000000
1!
1*
b1 6
19
1>
1C
b1 G
#185560000000
0!
0*
09
0>
0C
#185570000000
1!
1*
b10 6
19
1>
1C
b10 G
#185580000000
0!
0*
09
0>
0C
#185590000000
1!
1*
b11 6
19
1>
1C
b11 G
#185600000000
0!
0*
09
0>
0C
#185610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#185620000000
0!
0*
09
0>
0C
#185630000000
1!
1*
b101 6
19
1>
1C
b101 G
#185640000000
0!
0*
09
0>
0C
#185650000000
1!
1*
b110 6
19
1>
1C
b110 G
#185660000000
0!
0*
09
0>
0C
#185670000000
1!
1*
b111 6
19
1>
1C
b111 G
#185680000000
0!
1"
0*
1+
09
1:
0>
0C
#185690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#185700000000
0!
0*
09
0>
0C
#185710000000
1!
1*
b1 6
19
1>
1C
b1 G
#185720000000
0!
0*
09
0>
0C
#185730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#185740000000
0!
0*
09
0>
0C
#185750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#185760000000
0!
0*
09
0>
0C
#185770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#185780000000
0!
0*
09
0>
0C
#185790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#185800000000
0!
0#
0*
0,
09
0>
0?
0C
#185810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#185820000000
0!
0*
09
0>
0C
#185830000000
1!
1*
19
1>
1C
#185840000000
0!
0*
09
0>
0C
#185850000000
1!
1*
19
1>
1C
#185860000000
0!
0*
09
0>
0C
#185870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#185880000000
0!
0*
09
0>
0C
#185890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#185900000000
0!
0*
09
0>
0C
#185910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#185920000000
0!
0*
09
0>
0C
#185930000000
1!
1*
b10 6
19
1>
1C
b10 G
#185940000000
0!
0*
09
0>
0C
#185950000000
1!
1*
b11 6
19
1>
1C
b11 G
#185960000000
0!
0*
09
0>
0C
#185970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#185980000000
0!
0*
09
0>
0C
#185990000000
1!
1*
b101 6
19
1>
1C
b101 G
#186000000000
0!
0*
09
0>
0C
#186010000000
1!
1*
b110 6
19
1>
1C
b110 G
#186020000000
0!
0*
09
0>
0C
#186030000000
1!
1*
b111 6
19
1>
1C
b111 G
#186040000000
0!
0*
09
0>
0C
#186050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#186060000000
0!
0*
09
0>
0C
#186070000000
1!
1*
b1 6
19
1>
1C
b1 G
#186080000000
0!
0*
09
0>
0C
#186090000000
1!
1*
b10 6
19
1>
1C
b10 G
#186100000000
0!
0*
09
0>
0C
#186110000000
1!
1*
b11 6
19
1>
1C
b11 G
#186120000000
0!
0*
09
0>
0C
#186130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#186140000000
0!
0*
09
0>
0C
#186150000000
1!
1*
b101 6
19
1>
1C
b101 G
#186160000000
0!
0*
09
0>
0C
#186170000000
1!
1*
b110 6
19
1>
1C
b110 G
#186180000000
0!
0*
09
0>
0C
#186190000000
1!
1*
b111 6
19
1>
1C
b111 G
#186200000000
0!
0*
09
0>
0C
#186210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#186220000000
0!
0*
09
0>
0C
#186230000000
1!
1*
b1 6
19
1>
1C
b1 G
#186240000000
0!
0*
09
0>
0C
#186250000000
1!
1*
b10 6
19
1>
1C
b10 G
#186260000000
0!
0*
09
0>
0C
#186270000000
1!
1*
b11 6
19
1>
1C
b11 G
#186280000000
0!
0*
09
0>
0C
#186290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#186300000000
0!
0*
09
0>
0C
#186310000000
1!
1*
b101 6
19
1>
1C
b101 G
#186320000000
0!
0*
09
0>
0C
#186330000000
1!
1*
b110 6
19
1>
1C
b110 G
#186340000000
0!
0*
09
0>
0C
#186350000000
1!
1*
b111 6
19
1>
1C
b111 G
#186360000000
0!
1"
0*
1+
09
1:
0>
0C
#186370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#186380000000
0!
0*
09
0>
0C
#186390000000
1!
1*
b1 6
19
1>
1C
b1 G
#186400000000
0!
0*
09
0>
0C
#186410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#186420000000
0!
0*
09
0>
0C
#186430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#186440000000
0!
0*
09
0>
0C
#186450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#186460000000
0!
0*
09
0>
0C
#186470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#186480000000
0!
0#
0*
0,
09
0>
0?
0C
#186490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#186500000000
0!
0*
09
0>
0C
#186510000000
1!
1*
19
1>
1C
#186520000000
0!
0*
09
0>
0C
#186530000000
1!
1*
19
1>
1C
#186540000000
0!
0*
09
0>
0C
#186550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#186560000000
0!
0*
09
0>
0C
#186570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#186580000000
0!
0*
09
0>
0C
#186590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#186600000000
0!
0*
09
0>
0C
#186610000000
1!
1*
b10 6
19
1>
1C
b10 G
#186620000000
0!
0*
09
0>
0C
#186630000000
1!
1*
b11 6
19
1>
1C
b11 G
#186640000000
0!
0*
09
0>
0C
#186650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#186660000000
0!
0*
09
0>
0C
#186670000000
1!
1*
b101 6
19
1>
1C
b101 G
#186680000000
0!
0*
09
0>
0C
#186690000000
1!
1*
b110 6
19
1>
1C
b110 G
#186700000000
0!
0*
09
0>
0C
#186710000000
1!
1*
b111 6
19
1>
1C
b111 G
#186720000000
0!
0*
09
0>
0C
#186730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#186740000000
0!
0*
09
0>
0C
#186750000000
1!
1*
b1 6
19
1>
1C
b1 G
#186760000000
0!
0*
09
0>
0C
#186770000000
1!
1*
b10 6
19
1>
1C
b10 G
#186780000000
0!
0*
09
0>
0C
#186790000000
1!
1*
b11 6
19
1>
1C
b11 G
#186800000000
0!
0*
09
0>
0C
#186810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#186820000000
0!
0*
09
0>
0C
#186830000000
1!
1*
b101 6
19
1>
1C
b101 G
#186840000000
0!
0*
09
0>
0C
#186850000000
1!
1*
b110 6
19
1>
1C
b110 G
#186860000000
0!
0*
09
0>
0C
#186870000000
1!
1*
b111 6
19
1>
1C
b111 G
#186880000000
0!
0*
09
0>
0C
#186890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#186900000000
0!
0*
09
0>
0C
#186910000000
1!
1*
b1 6
19
1>
1C
b1 G
#186920000000
0!
0*
09
0>
0C
#186930000000
1!
1*
b10 6
19
1>
1C
b10 G
#186940000000
0!
0*
09
0>
0C
#186950000000
1!
1*
b11 6
19
1>
1C
b11 G
#186960000000
0!
0*
09
0>
0C
#186970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#186980000000
0!
0*
09
0>
0C
#186990000000
1!
1*
b101 6
19
1>
1C
b101 G
#187000000000
0!
0*
09
0>
0C
#187010000000
1!
1*
b110 6
19
1>
1C
b110 G
#187020000000
0!
0*
09
0>
0C
#187030000000
1!
1*
b111 6
19
1>
1C
b111 G
#187040000000
0!
1"
0*
1+
09
1:
0>
0C
#187050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#187060000000
0!
0*
09
0>
0C
#187070000000
1!
1*
b1 6
19
1>
1C
b1 G
#187080000000
0!
0*
09
0>
0C
#187090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#187100000000
0!
0*
09
0>
0C
#187110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#187120000000
0!
0*
09
0>
0C
#187130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#187140000000
0!
0*
09
0>
0C
#187150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#187160000000
0!
0#
0*
0,
09
0>
0?
0C
#187170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#187180000000
0!
0*
09
0>
0C
#187190000000
1!
1*
19
1>
1C
#187200000000
0!
0*
09
0>
0C
#187210000000
1!
1*
19
1>
1C
#187220000000
0!
0*
09
0>
0C
#187230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#187240000000
0!
0*
09
0>
0C
#187250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#187260000000
0!
0*
09
0>
0C
#187270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#187280000000
0!
0*
09
0>
0C
#187290000000
1!
1*
b10 6
19
1>
1C
b10 G
#187300000000
0!
0*
09
0>
0C
#187310000000
1!
1*
b11 6
19
1>
1C
b11 G
#187320000000
0!
0*
09
0>
0C
#187330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#187340000000
0!
0*
09
0>
0C
#187350000000
1!
1*
b101 6
19
1>
1C
b101 G
#187360000000
0!
0*
09
0>
0C
#187370000000
1!
1*
b110 6
19
1>
1C
b110 G
#187380000000
0!
0*
09
0>
0C
#187390000000
1!
1*
b111 6
19
1>
1C
b111 G
#187400000000
0!
0*
09
0>
0C
#187410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#187420000000
0!
0*
09
0>
0C
#187430000000
1!
1*
b1 6
19
1>
1C
b1 G
#187440000000
0!
0*
09
0>
0C
#187450000000
1!
1*
b10 6
19
1>
1C
b10 G
#187460000000
0!
0*
09
0>
0C
#187470000000
1!
1*
b11 6
19
1>
1C
b11 G
#187480000000
0!
0*
09
0>
0C
#187490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#187500000000
0!
0*
09
0>
0C
#187510000000
1!
1*
b101 6
19
1>
1C
b101 G
#187520000000
0!
0*
09
0>
0C
#187530000000
1!
1*
b110 6
19
1>
1C
b110 G
#187540000000
0!
0*
09
0>
0C
#187550000000
1!
1*
b111 6
19
1>
1C
b111 G
#187560000000
0!
0*
09
0>
0C
#187570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#187580000000
0!
0*
09
0>
0C
#187590000000
1!
1*
b1 6
19
1>
1C
b1 G
#187600000000
0!
0*
09
0>
0C
#187610000000
1!
1*
b10 6
19
1>
1C
b10 G
#187620000000
0!
0*
09
0>
0C
#187630000000
1!
1*
b11 6
19
1>
1C
b11 G
#187640000000
0!
0*
09
0>
0C
#187650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#187660000000
0!
0*
09
0>
0C
#187670000000
1!
1*
b101 6
19
1>
1C
b101 G
#187680000000
0!
0*
09
0>
0C
#187690000000
1!
1*
b110 6
19
1>
1C
b110 G
#187700000000
0!
0*
09
0>
0C
#187710000000
1!
1*
b111 6
19
1>
1C
b111 G
#187720000000
0!
1"
0*
1+
09
1:
0>
0C
#187730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#187740000000
0!
0*
09
0>
0C
#187750000000
1!
1*
b1 6
19
1>
1C
b1 G
#187760000000
0!
0*
09
0>
0C
#187770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#187780000000
0!
0*
09
0>
0C
#187790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#187800000000
0!
0*
09
0>
0C
#187810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#187820000000
0!
0*
09
0>
0C
#187830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#187840000000
0!
0#
0*
0,
09
0>
0?
0C
#187850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#187860000000
0!
0*
09
0>
0C
#187870000000
1!
1*
19
1>
1C
#187880000000
0!
0*
09
0>
0C
#187890000000
1!
1*
19
1>
1C
#187900000000
0!
0*
09
0>
0C
#187910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#187920000000
0!
0*
09
0>
0C
#187930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#187940000000
0!
0*
09
0>
0C
#187950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#187960000000
0!
0*
09
0>
0C
#187970000000
1!
1*
b10 6
19
1>
1C
b10 G
#187980000000
0!
0*
09
0>
0C
#187990000000
1!
1*
b11 6
19
1>
1C
b11 G
#188000000000
0!
0*
09
0>
0C
#188010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#188020000000
0!
0*
09
0>
0C
#188030000000
1!
1*
b101 6
19
1>
1C
b101 G
#188040000000
0!
0*
09
0>
0C
#188050000000
1!
1*
b110 6
19
1>
1C
b110 G
#188060000000
0!
0*
09
0>
0C
#188070000000
1!
1*
b111 6
19
1>
1C
b111 G
#188080000000
0!
0*
09
0>
0C
#188090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#188100000000
0!
0*
09
0>
0C
#188110000000
1!
1*
b1 6
19
1>
1C
b1 G
#188120000000
0!
0*
09
0>
0C
#188130000000
1!
1*
b10 6
19
1>
1C
b10 G
#188140000000
0!
0*
09
0>
0C
#188150000000
1!
1*
b11 6
19
1>
1C
b11 G
#188160000000
0!
0*
09
0>
0C
#188170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#188180000000
0!
0*
09
0>
0C
#188190000000
1!
1*
b101 6
19
1>
1C
b101 G
#188200000000
0!
0*
09
0>
0C
#188210000000
1!
1*
b110 6
19
1>
1C
b110 G
#188220000000
0!
0*
09
0>
0C
#188230000000
1!
1*
b111 6
19
1>
1C
b111 G
#188240000000
0!
0*
09
0>
0C
#188250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#188260000000
0!
0*
09
0>
0C
#188270000000
1!
1*
b1 6
19
1>
1C
b1 G
#188280000000
0!
0*
09
0>
0C
#188290000000
1!
1*
b10 6
19
1>
1C
b10 G
#188300000000
0!
0*
09
0>
0C
#188310000000
1!
1*
b11 6
19
1>
1C
b11 G
#188320000000
0!
0*
09
0>
0C
#188330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#188340000000
0!
0*
09
0>
0C
#188350000000
1!
1*
b101 6
19
1>
1C
b101 G
#188360000000
0!
0*
09
0>
0C
#188370000000
1!
1*
b110 6
19
1>
1C
b110 G
#188380000000
0!
0*
09
0>
0C
#188390000000
1!
1*
b111 6
19
1>
1C
b111 G
#188400000000
0!
1"
0*
1+
09
1:
0>
0C
#188410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#188420000000
0!
0*
09
0>
0C
#188430000000
1!
1*
b1 6
19
1>
1C
b1 G
#188440000000
0!
0*
09
0>
0C
#188450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#188460000000
0!
0*
09
0>
0C
#188470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#188480000000
0!
0*
09
0>
0C
#188490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#188500000000
0!
0*
09
0>
0C
#188510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#188520000000
0!
0#
0*
0,
09
0>
0?
0C
#188530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#188540000000
0!
0*
09
0>
0C
#188550000000
1!
1*
19
1>
1C
#188560000000
0!
0*
09
0>
0C
#188570000000
1!
1*
19
1>
1C
#188580000000
0!
0*
09
0>
0C
#188590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#188600000000
0!
0*
09
0>
0C
#188610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#188620000000
0!
0*
09
0>
0C
#188630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#188640000000
0!
0*
09
0>
0C
#188650000000
1!
1*
b10 6
19
1>
1C
b10 G
#188660000000
0!
0*
09
0>
0C
#188670000000
1!
1*
b11 6
19
1>
1C
b11 G
#188680000000
0!
0*
09
0>
0C
#188690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#188700000000
0!
0*
09
0>
0C
#188710000000
1!
1*
b101 6
19
1>
1C
b101 G
#188720000000
0!
0*
09
0>
0C
#188730000000
1!
1*
b110 6
19
1>
1C
b110 G
#188740000000
0!
0*
09
0>
0C
#188750000000
1!
1*
b111 6
19
1>
1C
b111 G
#188760000000
0!
0*
09
0>
0C
#188770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#188780000000
0!
0*
09
0>
0C
#188790000000
1!
1*
b1 6
19
1>
1C
b1 G
#188800000000
0!
0*
09
0>
0C
#188810000000
1!
1*
b10 6
19
1>
1C
b10 G
#188820000000
0!
0*
09
0>
0C
#188830000000
1!
1*
b11 6
19
1>
1C
b11 G
#188840000000
0!
0*
09
0>
0C
#188850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#188860000000
0!
0*
09
0>
0C
#188870000000
1!
1*
b101 6
19
1>
1C
b101 G
#188880000000
0!
0*
09
0>
0C
#188890000000
1!
1*
b110 6
19
1>
1C
b110 G
#188900000000
0!
0*
09
0>
0C
#188910000000
1!
1*
b111 6
19
1>
1C
b111 G
#188920000000
0!
0*
09
0>
0C
#188930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#188940000000
0!
0*
09
0>
0C
#188950000000
1!
1*
b1 6
19
1>
1C
b1 G
#188960000000
0!
0*
09
0>
0C
#188970000000
1!
1*
b10 6
19
1>
1C
b10 G
#188980000000
0!
0*
09
0>
0C
#188990000000
1!
1*
b11 6
19
1>
1C
b11 G
#189000000000
0!
0*
09
0>
0C
#189010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#189020000000
0!
0*
09
0>
0C
#189030000000
1!
1*
b101 6
19
1>
1C
b101 G
#189040000000
0!
0*
09
0>
0C
#189050000000
1!
1*
b110 6
19
1>
1C
b110 G
#189060000000
0!
0*
09
0>
0C
#189070000000
1!
1*
b111 6
19
1>
1C
b111 G
#189080000000
0!
1"
0*
1+
09
1:
0>
0C
#189090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#189100000000
0!
0*
09
0>
0C
#189110000000
1!
1*
b1 6
19
1>
1C
b1 G
#189120000000
0!
0*
09
0>
0C
#189130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#189140000000
0!
0*
09
0>
0C
#189150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#189160000000
0!
0*
09
0>
0C
#189170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#189180000000
0!
0*
09
0>
0C
#189190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#189200000000
0!
0#
0*
0,
09
0>
0?
0C
#189210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#189220000000
0!
0*
09
0>
0C
#189230000000
1!
1*
19
1>
1C
#189240000000
0!
0*
09
0>
0C
#189250000000
1!
1*
19
1>
1C
#189260000000
0!
0*
09
0>
0C
#189270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#189280000000
0!
0*
09
0>
0C
#189290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#189300000000
0!
0*
09
0>
0C
#189310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#189320000000
0!
0*
09
0>
0C
#189330000000
1!
1*
b10 6
19
1>
1C
b10 G
#189340000000
0!
0*
09
0>
0C
#189350000000
1!
1*
b11 6
19
1>
1C
b11 G
#189360000000
0!
0*
09
0>
0C
#189370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#189380000000
0!
0*
09
0>
0C
#189390000000
1!
1*
b101 6
19
1>
1C
b101 G
#189400000000
0!
0*
09
0>
0C
#189410000000
1!
1*
b110 6
19
1>
1C
b110 G
#189420000000
0!
0*
09
0>
0C
#189430000000
1!
1*
b111 6
19
1>
1C
b111 G
#189440000000
0!
0*
09
0>
0C
#189450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#189460000000
0!
0*
09
0>
0C
#189470000000
1!
1*
b1 6
19
1>
1C
b1 G
#189480000000
0!
0*
09
0>
0C
#189490000000
1!
1*
b10 6
19
1>
1C
b10 G
#189500000000
0!
0*
09
0>
0C
#189510000000
1!
1*
b11 6
19
1>
1C
b11 G
#189520000000
0!
0*
09
0>
0C
#189530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#189540000000
0!
0*
09
0>
0C
#189550000000
1!
1*
b101 6
19
1>
1C
b101 G
#189560000000
0!
0*
09
0>
0C
#189570000000
1!
1*
b110 6
19
1>
1C
b110 G
#189580000000
0!
0*
09
0>
0C
#189590000000
1!
1*
b111 6
19
1>
1C
b111 G
#189600000000
0!
0*
09
0>
0C
#189610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#189620000000
0!
0*
09
0>
0C
#189630000000
1!
1*
b1 6
19
1>
1C
b1 G
#189640000000
0!
0*
09
0>
0C
#189650000000
1!
1*
b10 6
19
1>
1C
b10 G
#189660000000
0!
0*
09
0>
0C
#189670000000
1!
1*
b11 6
19
1>
1C
b11 G
#189680000000
0!
0*
09
0>
0C
#189690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#189700000000
0!
0*
09
0>
0C
#189710000000
1!
1*
b101 6
19
1>
1C
b101 G
#189720000000
0!
0*
09
0>
0C
#189730000000
1!
1*
b110 6
19
1>
1C
b110 G
#189740000000
0!
0*
09
0>
0C
#189750000000
1!
1*
b111 6
19
1>
1C
b111 G
#189760000000
0!
1"
0*
1+
09
1:
0>
0C
#189770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#189780000000
0!
0*
09
0>
0C
#189790000000
1!
1*
b1 6
19
1>
1C
b1 G
#189800000000
0!
0*
09
0>
0C
#189810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#189820000000
0!
0*
09
0>
0C
#189830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#189840000000
0!
0*
09
0>
0C
#189850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#189860000000
0!
0*
09
0>
0C
#189870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#189880000000
0!
0#
0*
0,
09
0>
0?
0C
#189890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#189900000000
0!
0*
09
0>
0C
#189910000000
1!
1*
19
1>
1C
#189920000000
0!
0*
09
0>
0C
#189930000000
1!
1*
19
1>
1C
#189940000000
0!
0*
09
0>
0C
#189950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#189960000000
0!
0*
09
0>
0C
#189970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#189980000000
0!
0*
09
0>
0C
#189990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#190000000000
0!
0*
09
0>
0C
#190010000000
1!
1*
b10 6
19
1>
1C
b10 G
#190020000000
0!
0*
09
0>
0C
#190030000000
1!
1*
b11 6
19
1>
1C
b11 G
#190040000000
0!
0*
09
0>
0C
#190050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#190060000000
0!
0*
09
0>
0C
#190070000000
1!
1*
b101 6
19
1>
1C
b101 G
#190080000000
0!
0*
09
0>
0C
#190090000000
1!
1*
b110 6
19
1>
1C
b110 G
#190100000000
0!
0*
09
0>
0C
#190110000000
1!
1*
b111 6
19
1>
1C
b111 G
#190120000000
0!
0*
09
0>
0C
#190130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#190140000000
0!
0*
09
0>
0C
#190150000000
1!
1*
b1 6
19
1>
1C
b1 G
#190160000000
0!
0*
09
0>
0C
#190170000000
1!
1*
b10 6
19
1>
1C
b10 G
#190180000000
0!
0*
09
0>
0C
#190190000000
1!
1*
b11 6
19
1>
1C
b11 G
#190200000000
0!
0*
09
0>
0C
#190210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#190220000000
0!
0*
09
0>
0C
#190230000000
1!
1*
b101 6
19
1>
1C
b101 G
#190240000000
0!
0*
09
0>
0C
#190250000000
1!
1*
b110 6
19
1>
1C
b110 G
#190260000000
0!
0*
09
0>
0C
#190270000000
1!
1*
b111 6
19
1>
1C
b111 G
#190280000000
0!
0*
09
0>
0C
#190290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#190300000000
0!
0*
09
0>
0C
#190310000000
1!
1*
b1 6
19
1>
1C
b1 G
#190320000000
0!
0*
09
0>
0C
#190330000000
1!
1*
b10 6
19
1>
1C
b10 G
#190340000000
0!
0*
09
0>
0C
#190350000000
1!
1*
b11 6
19
1>
1C
b11 G
#190360000000
0!
0*
09
0>
0C
#190370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#190380000000
0!
0*
09
0>
0C
#190390000000
1!
1*
b101 6
19
1>
1C
b101 G
#190400000000
0!
0*
09
0>
0C
#190410000000
1!
1*
b110 6
19
1>
1C
b110 G
#190420000000
0!
0*
09
0>
0C
#190430000000
1!
1*
b111 6
19
1>
1C
b111 G
#190440000000
0!
1"
0*
1+
09
1:
0>
0C
#190450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#190460000000
0!
0*
09
0>
0C
#190470000000
1!
1*
b1 6
19
1>
1C
b1 G
#190480000000
0!
0*
09
0>
0C
#190490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#190500000000
0!
0*
09
0>
0C
#190510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#190520000000
0!
0*
09
0>
0C
#190530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#190540000000
0!
0*
09
0>
0C
#190550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#190560000000
0!
0#
0*
0,
09
0>
0?
0C
#190570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#190580000000
0!
0*
09
0>
0C
#190590000000
1!
1*
19
1>
1C
#190600000000
0!
0*
09
0>
0C
#190610000000
1!
1*
19
1>
1C
#190620000000
0!
0*
09
0>
0C
#190630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#190640000000
0!
0*
09
0>
0C
#190650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#190660000000
0!
0*
09
0>
0C
#190670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#190680000000
0!
0*
09
0>
0C
#190690000000
1!
1*
b10 6
19
1>
1C
b10 G
#190700000000
0!
0*
09
0>
0C
#190710000000
1!
1*
b11 6
19
1>
1C
b11 G
#190720000000
0!
0*
09
0>
0C
#190730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#190740000000
0!
0*
09
0>
0C
#190750000000
1!
1*
b101 6
19
1>
1C
b101 G
#190760000000
0!
0*
09
0>
0C
#190770000000
1!
1*
b110 6
19
1>
1C
b110 G
#190780000000
0!
0*
09
0>
0C
#190790000000
1!
1*
b111 6
19
1>
1C
b111 G
#190800000000
0!
0*
09
0>
0C
#190810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#190820000000
0!
0*
09
0>
0C
#190830000000
1!
1*
b1 6
19
1>
1C
b1 G
#190840000000
0!
0*
09
0>
0C
#190850000000
1!
1*
b10 6
19
1>
1C
b10 G
#190860000000
0!
0*
09
0>
0C
#190870000000
1!
1*
b11 6
19
1>
1C
b11 G
#190880000000
0!
0*
09
0>
0C
#190890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#190900000000
0!
0*
09
0>
0C
#190910000000
1!
1*
b101 6
19
1>
1C
b101 G
#190920000000
0!
0*
09
0>
0C
#190930000000
1!
1*
b110 6
19
1>
1C
b110 G
#190940000000
0!
0*
09
0>
0C
#190950000000
1!
1*
b111 6
19
1>
1C
b111 G
#190960000000
0!
0*
09
0>
0C
#190970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#190980000000
0!
0*
09
0>
0C
#190990000000
1!
1*
b1 6
19
1>
1C
b1 G
#191000000000
0!
0*
09
0>
0C
#191010000000
1!
1*
b10 6
19
1>
1C
b10 G
#191020000000
0!
0*
09
0>
0C
#191030000000
1!
1*
b11 6
19
1>
1C
b11 G
#191040000000
0!
0*
09
0>
0C
#191050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#191060000000
0!
0*
09
0>
0C
#191070000000
1!
1*
b101 6
19
1>
1C
b101 G
#191080000000
0!
0*
09
0>
0C
#191090000000
1!
1*
b110 6
19
1>
1C
b110 G
#191100000000
0!
0*
09
0>
0C
#191110000000
1!
1*
b111 6
19
1>
1C
b111 G
#191120000000
0!
1"
0*
1+
09
1:
0>
0C
#191130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#191140000000
0!
0*
09
0>
0C
#191150000000
1!
1*
b1 6
19
1>
1C
b1 G
#191160000000
0!
0*
09
0>
0C
#191170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#191180000000
0!
0*
09
0>
0C
#191190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#191200000000
0!
0*
09
0>
0C
#191210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#191220000000
0!
0*
09
0>
0C
#191230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#191240000000
0!
0#
0*
0,
09
0>
0?
0C
#191250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#191260000000
0!
0*
09
0>
0C
#191270000000
1!
1*
19
1>
1C
#191280000000
0!
0*
09
0>
0C
#191290000000
1!
1*
19
1>
1C
#191300000000
0!
0*
09
0>
0C
#191310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#191320000000
0!
0*
09
0>
0C
#191330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#191340000000
0!
0*
09
0>
0C
#191350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#191360000000
0!
0*
09
0>
0C
#191370000000
1!
1*
b10 6
19
1>
1C
b10 G
#191380000000
0!
0*
09
0>
0C
#191390000000
1!
1*
b11 6
19
1>
1C
b11 G
#191400000000
0!
0*
09
0>
0C
#191410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#191420000000
0!
0*
09
0>
0C
#191430000000
1!
1*
b101 6
19
1>
1C
b101 G
#191440000000
0!
0*
09
0>
0C
#191450000000
1!
1*
b110 6
19
1>
1C
b110 G
#191460000000
0!
0*
09
0>
0C
#191470000000
1!
1*
b111 6
19
1>
1C
b111 G
#191480000000
0!
0*
09
0>
0C
#191490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#191500000000
0!
0*
09
0>
0C
#191510000000
1!
1*
b1 6
19
1>
1C
b1 G
#191520000000
0!
0*
09
0>
0C
#191530000000
1!
1*
b10 6
19
1>
1C
b10 G
#191540000000
0!
0*
09
0>
0C
#191550000000
1!
1*
b11 6
19
1>
1C
b11 G
#191560000000
0!
0*
09
0>
0C
#191570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#191580000000
0!
0*
09
0>
0C
#191590000000
1!
1*
b101 6
19
1>
1C
b101 G
#191600000000
0!
0*
09
0>
0C
#191610000000
1!
1*
b110 6
19
1>
1C
b110 G
#191620000000
0!
0*
09
0>
0C
#191630000000
1!
1*
b111 6
19
1>
1C
b111 G
#191640000000
0!
0*
09
0>
0C
#191650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#191660000000
0!
0*
09
0>
0C
#191670000000
1!
1*
b1 6
19
1>
1C
b1 G
#191680000000
0!
0*
09
0>
0C
#191690000000
1!
1*
b10 6
19
1>
1C
b10 G
#191700000000
0!
0*
09
0>
0C
#191710000000
1!
1*
b11 6
19
1>
1C
b11 G
#191720000000
0!
0*
09
0>
0C
#191730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#191740000000
0!
0*
09
0>
0C
#191750000000
1!
1*
b101 6
19
1>
1C
b101 G
#191760000000
0!
0*
09
0>
0C
#191770000000
1!
1*
b110 6
19
1>
1C
b110 G
#191780000000
0!
0*
09
0>
0C
#191790000000
1!
1*
b111 6
19
1>
1C
b111 G
#191800000000
0!
1"
0*
1+
09
1:
0>
0C
#191810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#191820000000
0!
0*
09
0>
0C
#191830000000
1!
1*
b1 6
19
1>
1C
b1 G
#191840000000
0!
0*
09
0>
0C
#191850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#191860000000
0!
0*
09
0>
0C
#191870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#191880000000
0!
0*
09
0>
0C
#191890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#191900000000
0!
0*
09
0>
0C
#191910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#191920000000
0!
0#
0*
0,
09
0>
0?
0C
#191930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#191940000000
0!
0*
09
0>
0C
#191950000000
1!
1*
19
1>
1C
#191960000000
0!
0*
09
0>
0C
#191970000000
1!
1*
19
1>
1C
#191980000000
0!
0*
09
0>
0C
#191990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#192000000000
0!
0*
09
0>
0C
#192010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#192020000000
0!
0*
09
0>
0C
#192030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#192040000000
0!
0*
09
0>
0C
#192050000000
1!
1*
b10 6
19
1>
1C
b10 G
#192060000000
0!
0*
09
0>
0C
#192070000000
1!
1*
b11 6
19
1>
1C
b11 G
#192080000000
0!
0*
09
0>
0C
#192090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#192100000000
0!
0*
09
0>
0C
#192110000000
1!
1*
b101 6
19
1>
1C
b101 G
#192120000000
0!
0*
09
0>
0C
#192130000000
1!
1*
b110 6
19
1>
1C
b110 G
#192140000000
0!
0*
09
0>
0C
#192150000000
1!
1*
b111 6
19
1>
1C
b111 G
#192160000000
0!
0*
09
0>
0C
#192170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#192180000000
0!
0*
09
0>
0C
#192190000000
1!
1*
b1 6
19
1>
1C
b1 G
#192200000000
0!
0*
09
0>
0C
#192210000000
1!
1*
b10 6
19
1>
1C
b10 G
#192220000000
0!
0*
09
0>
0C
#192230000000
1!
1*
b11 6
19
1>
1C
b11 G
#192240000000
0!
0*
09
0>
0C
#192250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#192260000000
0!
0*
09
0>
0C
#192270000000
1!
1*
b101 6
19
1>
1C
b101 G
#192280000000
0!
0*
09
0>
0C
#192290000000
1!
1*
b110 6
19
1>
1C
b110 G
#192300000000
0!
0*
09
0>
0C
#192310000000
1!
1*
b111 6
19
1>
1C
b111 G
#192320000000
0!
0*
09
0>
0C
#192330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#192340000000
0!
0*
09
0>
0C
#192350000000
1!
1*
b1 6
19
1>
1C
b1 G
#192360000000
0!
0*
09
0>
0C
#192370000000
1!
1*
b10 6
19
1>
1C
b10 G
#192380000000
0!
0*
09
0>
0C
#192390000000
1!
1*
b11 6
19
1>
1C
b11 G
#192400000000
0!
0*
09
0>
0C
#192410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#192420000000
0!
0*
09
0>
0C
#192430000000
1!
1*
b101 6
19
1>
1C
b101 G
#192440000000
0!
0*
09
0>
0C
#192450000000
1!
1*
b110 6
19
1>
1C
b110 G
#192460000000
0!
0*
09
0>
0C
#192470000000
1!
1*
b111 6
19
1>
1C
b111 G
#192480000000
0!
1"
0*
1+
09
1:
0>
0C
#192490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#192500000000
0!
0*
09
0>
0C
#192510000000
1!
1*
b1 6
19
1>
1C
b1 G
#192520000000
0!
0*
09
0>
0C
#192530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#192540000000
0!
0*
09
0>
0C
#192550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#192560000000
0!
0*
09
0>
0C
#192570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#192580000000
0!
0*
09
0>
0C
#192590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#192600000000
0!
0#
0*
0,
09
0>
0?
0C
#192610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#192620000000
0!
0*
09
0>
0C
#192630000000
1!
1*
19
1>
1C
#192640000000
0!
0*
09
0>
0C
#192650000000
1!
1*
19
1>
1C
#192660000000
0!
0*
09
0>
0C
#192670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#192680000000
0!
0*
09
0>
0C
#192690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#192700000000
0!
0*
09
0>
0C
#192710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#192720000000
0!
0*
09
0>
0C
#192730000000
1!
1*
b10 6
19
1>
1C
b10 G
#192740000000
0!
0*
09
0>
0C
#192750000000
1!
1*
b11 6
19
1>
1C
b11 G
#192760000000
0!
0*
09
0>
0C
#192770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#192780000000
0!
0*
09
0>
0C
#192790000000
1!
1*
b101 6
19
1>
1C
b101 G
#192800000000
0!
0*
09
0>
0C
#192810000000
1!
1*
b110 6
19
1>
1C
b110 G
#192820000000
0!
0*
09
0>
0C
#192830000000
1!
1*
b111 6
19
1>
1C
b111 G
#192840000000
0!
0*
09
0>
0C
#192850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#192860000000
0!
0*
09
0>
0C
#192870000000
1!
1*
b1 6
19
1>
1C
b1 G
#192880000000
0!
0*
09
0>
0C
#192890000000
1!
1*
b10 6
19
1>
1C
b10 G
#192900000000
0!
0*
09
0>
0C
#192910000000
1!
1*
b11 6
19
1>
1C
b11 G
#192920000000
0!
0*
09
0>
0C
#192930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#192940000000
0!
0*
09
0>
0C
#192950000000
1!
1*
b101 6
19
1>
1C
b101 G
#192960000000
0!
0*
09
0>
0C
#192970000000
1!
1*
b110 6
19
1>
1C
b110 G
#192980000000
0!
0*
09
0>
0C
#192990000000
1!
1*
b111 6
19
1>
1C
b111 G
#193000000000
0!
0*
09
0>
0C
#193010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#193020000000
0!
0*
09
0>
0C
#193030000000
1!
1*
b1 6
19
1>
1C
b1 G
#193040000000
0!
0*
09
0>
0C
#193050000000
1!
1*
b10 6
19
1>
1C
b10 G
#193060000000
0!
0*
09
0>
0C
#193070000000
1!
1*
b11 6
19
1>
1C
b11 G
#193080000000
0!
0*
09
0>
0C
#193090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#193100000000
0!
0*
09
0>
0C
#193110000000
1!
1*
b101 6
19
1>
1C
b101 G
#193120000000
0!
0*
09
0>
0C
#193130000000
1!
1*
b110 6
19
1>
1C
b110 G
#193140000000
0!
0*
09
0>
0C
#193150000000
1!
1*
b111 6
19
1>
1C
b111 G
#193160000000
0!
1"
0*
1+
09
1:
0>
0C
#193170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#193180000000
0!
0*
09
0>
0C
#193190000000
1!
1*
b1 6
19
1>
1C
b1 G
#193200000000
0!
0*
09
0>
0C
#193210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#193220000000
0!
0*
09
0>
0C
#193230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#193240000000
0!
0*
09
0>
0C
#193250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#193260000000
0!
0*
09
0>
0C
#193270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#193280000000
0!
0#
0*
0,
09
0>
0?
0C
#193290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#193300000000
0!
0*
09
0>
0C
#193310000000
1!
1*
19
1>
1C
#193320000000
0!
0*
09
0>
0C
#193330000000
1!
1*
19
1>
1C
#193340000000
0!
0*
09
0>
0C
#193350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#193360000000
0!
0*
09
0>
0C
#193370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#193380000000
0!
0*
09
0>
0C
#193390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#193400000000
0!
0*
09
0>
0C
#193410000000
1!
1*
b10 6
19
1>
1C
b10 G
#193420000000
0!
0*
09
0>
0C
#193430000000
1!
1*
b11 6
19
1>
1C
b11 G
#193440000000
0!
0*
09
0>
0C
#193450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#193460000000
0!
0*
09
0>
0C
#193470000000
1!
1*
b101 6
19
1>
1C
b101 G
#193480000000
0!
0*
09
0>
0C
#193490000000
1!
1*
b110 6
19
1>
1C
b110 G
#193500000000
0!
0*
09
0>
0C
#193510000000
1!
1*
b111 6
19
1>
1C
b111 G
#193520000000
0!
0*
09
0>
0C
#193530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#193540000000
0!
0*
09
0>
0C
#193550000000
1!
1*
b1 6
19
1>
1C
b1 G
#193560000000
0!
0*
09
0>
0C
#193570000000
1!
1*
b10 6
19
1>
1C
b10 G
#193580000000
0!
0*
09
0>
0C
#193590000000
1!
1*
b11 6
19
1>
1C
b11 G
#193600000000
0!
0*
09
0>
0C
#193610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#193620000000
0!
0*
09
0>
0C
#193630000000
1!
1*
b101 6
19
1>
1C
b101 G
#193640000000
0!
0*
09
0>
0C
#193650000000
1!
1*
b110 6
19
1>
1C
b110 G
#193660000000
0!
0*
09
0>
0C
#193670000000
1!
1*
b111 6
19
1>
1C
b111 G
#193680000000
0!
0*
09
0>
0C
#193690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#193700000000
0!
0*
09
0>
0C
#193710000000
1!
1*
b1 6
19
1>
1C
b1 G
#193720000000
0!
0*
09
0>
0C
#193730000000
1!
1*
b10 6
19
1>
1C
b10 G
#193740000000
0!
0*
09
0>
0C
#193750000000
1!
1*
b11 6
19
1>
1C
b11 G
#193760000000
0!
0*
09
0>
0C
#193770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#193780000000
0!
0*
09
0>
0C
#193790000000
1!
1*
b101 6
19
1>
1C
b101 G
#193800000000
0!
0*
09
0>
0C
#193810000000
1!
1*
b110 6
19
1>
1C
b110 G
#193820000000
0!
0*
09
0>
0C
#193830000000
1!
1*
b111 6
19
1>
1C
b111 G
#193840000000
0!
1"
0*
1+
09
1:
0>
0C
#193850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#193860000000
0!
0*
09
0>
0C
#193870000000
1!
1*
b1 6
19
1>
1C
b1 G
#193880000000
0!
0*
09
0>
0C
#193890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#193900000000
0!
0*
09
0>
0C
#193910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#193920000000
0!
0*
09
0>
0C
#193930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#193940000000
0!
0*
09
0>
0C
#193950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#193960000000
0!
0#
0*
0,
09
0>
0?
0C
#193970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#193980000000
0!
0*
09
0>
0C
#193990000000
1!
1*
19
1>
1C
#194000000000
0!
0*
09
0>
0C
#194010000000
1!
1*
19
1>
1C
#194020000000
0!
0*
09
0>
0C
#194030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#194040000000
0!
0*
09
0>
0C
#194050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#194060000000
0!
0*
09
0>
0C
#194070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#194080000000
0!
0*
09
0>
0C
#194090000000
1!
1*
b10 6
19
1>
1C
b10 G
#194100000000
0!
0*
09
0>
0C
#194110000000
1!
1*
b11 6
19
1>
1C
b11 G
#194120000000
0!
0*
09
0>
0C
#194130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#194140000000
0!
0*
09
0>
0C
#194150000000
1!
1*
b101 6
19
1>
1C
b101 G
#194160000000
0!
0*
09
0>
0C
#194170000000
1!
1*
b110 6
19
1>
1C
b110 G
#194180000000
0!
0*
09
0>
0C
#194190000000
1!
1*
b111 6
19
1>
1C
b111 G
#194200000000
0!
0*
09
0>
0C
#194210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#194220000000
0!
0*
09
0>
0C
#194230000000
1!
1*
b1 6
19
1>
1C
b1 G
#194240000000
0!
0*
09
0>
0C
#194250000000
1!
1*
b10 6
19
1>
1C
b10 G
#194260000000
0!
0*
09
0>
0C
#194270000000
1!
1*
b11 6
19
1>
1C
b11 G
#194280000000
0!
0*
09
0>
0C
#194290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#194300000000
0!
0*
09
0>
0C
#194310000000
1!
1*
b101 6
19
1>
1C
b101 G
#194320000000
0!
0*
09
0>
0C
#194330000000
1!
1*
b110 6
19
1>
1C
b110 G
#194340000000
0!
0*
09
0>
0C
#194350000000
1!
1*
b111 6
19
1>
1C
b111 G
#194360000000
0!
0*
09
0>
0C
#194370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#194380000000
0!
0*
09
0>
0C
#194390000000
1!
1*
b1 6
19
1>
1C
b1 G
#194400000000
0!
0*
09
0>
0C
#194410000000
1!
1*
b10 6
19
1>
1C
b10 G
#194420000000
0!
0*
09
0>
0C
#194430000000
1!
1*
b11 6
19
1>
1C
b11 G
#194440000000
0!
0*
09
0>
0C
#194450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#194460000000
0!
0*
09
0>
0C
#194470000000
1!
1*
b101 6
19
1>
1C
b101 G
#194480000000
0!
0*
09
0>
0C
#194490000000
1!
1*
b110 6
19
1>
1C
b110 G
#194500000000
0!
0*
09
0>
0C
#194510000000
1!
1*
b111 6
19
1>
1C
b111 G
#194520000000
0!
1"
0*
1+
09
1:
0>
0C
#194530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#194540000000
0!
0*
09
0>
0C
#194550000000
1!
1*
b1 6
19
1>
1C
b1 G
#194560000000
0!
0*
09
0>
0C
#194570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#194580000000
0!
0*
09
0>
0C
#194590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#194600000000
0!
0*
09
0>
0C
#194610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#194620000000
0!
0*
09
0>
0C
#194630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#194640000000
0!
0#
0*
0,
09
0>
0?
0C
#194650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#194660000000
0!
0*
09
0>
0C
#194670000000
1!
1*
19
1>
1C
#194680000000
0!
0*
09
0>
0C
#194690000000
1!
1*
19
1>
1C
#194700000000
0!
0*
09
0>
0C
#194710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#194720000000
0!
0*
09
0>
0C
#194730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#194740000000
0!
0*
09
0>
0C
#194750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#194760000000
0!
0*
09
0>
0C
#194770000000
1!
1*
b10 6
19
1>
1C
b10 G
#194780000000
0!
0*
09
0>
0C
#194790000000
1!
1*
b11 6
19
1>
1C
b11 G
#194800000000
0!
0*
09
0>
0C
#194810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#194820000000
0!
0*
09
0>
0C
#194830000000
1!
1*
b101 6
19
1>
1C
b101 G
#194840000000
0!
0*
09
0>
0C
#194850000000
1!
1*
b110 6
19
1>
1C
b110 G
#194860000000
0!
0*
09
0>
0C
#194870000000
1!
1*
b111 6
19
1>
1C
b111 G
#194880000000
0!
0*
09
0>
0C
#194890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#194900000000
0!
0*
09
0>
0C
#194910000000
1!
1*
b1 6
19
1>
1C
b1 G
#194920000000
0!
0*
09
0>
0C
#194930000000
1!
1*
b10 6
19
1>
1C
b10 G
#194940000000
0!
0*
09
0>
0C
#194950000000
1!
1*
b11 6
19
1>
1C
b11 G
#194960000000
0!
0*
09
0>
0C
#194970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#194980000000
0!
0*
09
0>
0C
#194990000000
1!
1*
b101 6
19
1>
1C
b101 G
#195000000000
0!
0*
09
0>
0C
#195010000000
1!
1*
b110 6
19
1>
1C
b110 G
#195020000000
0!
0*
09
0>
0C
#195030000000
1!
1*
b111 6
19
1>
1C
b111 G
#195040000000
0!
0*
09
0>
0C
#195050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#195060000000
0!
0*
09
0>
0C
#195070000000
1!
1*
b1 6
19
1>
1C
b1 G
#195080000000
0!
0*
09
0>
0C
#195090000000
1!
1*
b10 6
19
1>
1C
b10 G
#195100000000
0!
0*
09
0>
0C
#195110000000
1!
1*
b11 6
19
1>
1C
b11 G
#195120000000
0!
0*
09
0>
0C
#195130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#195140000000
0!
0*
09
0>
0C
#195150000000
1!
1*
b101 6
19
1>
1C
b101 G
#195160000000
0!
0*
09
0>
0C
#195170000000
1!
1*
b110 6
19
1>
1C
b110 G
#195180000000
0!
0*
09
0>
0C
#195190000000
1!
1*
b111 6
19
1>
1C
b111 G
#195200000000
0!
1"
0*
1+
09
1:
0>
0C
#195210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#195220000000
0!
0*
09
0>
0C
#195230000000
1!
1*
b1 6
19
1>
1C
b1 G
#195240000000
0!
0*
09
0>
0C
#195250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#195260000000
0!
0*
09
0>
0C
#195270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#195280000000
0!
0*
09
0>
0C
#195290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#195300000000
0!
0*
09
0>
0C
#195310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#195320000000
0!
0#
0*
0,
09
0>
0?
0C
#195330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#195340000000
0!
0*
09
0>
0C
#195350000000
1!
1*
19
1>
1C
#195360000000
0!
0*
09
0>
0C
#195370000000
1!
1*
19
1>
1C
#195380000000
0!
0*
09
0>
0C
#195390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#195400000000
0!
0*
09
0>
0C
#195410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#195420000000
0!
0*
09
0>
0C
#195430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#195440000000
0!
0*
09
0>
0C
#195450000000
1!
1*
b10 6
19
1>
1C
b10 G
#195460000000
0!
0*
09
0>
0C
#195470000000
1!
1*
b11 6
19
1>
1C
b11 G
#195480000000
0!
0*
09
0>
0C
#195490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#195500000000
0!
0*
09
0>
0C
#195510000000
1!
1*
b101 6
19
1>
1C
b101 G
#195520000000
0!
0*
09
0>
0C
#195530000000
1!
1*
b110 6
19
1>
1C
b110 G
#195540000000
0!
0*
09
0>
0C
#195550000000
1!
1*
b111 6
19
1>
1C
b111 G
#195560000000
0!
0*
09
0>
0C
#195570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#195580000000
0!
0*
09
0>
0C
#195590000000
1!
1*
b1 6
19
1>
1C
b1 G
#195600000000
0!
0*
09
0>
0C
#195610000000
1!
1*
b10 6
19
1>
1C
b10 G
#195620000000
0!
0*
09
0>
0C
#195630000000
1!
1*
b11 6
19
1>
1C
b11 G
#195640000000
0!
0*
09
0>
0C
#195650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#195660000000
0!
0*
09
0>
0C
#195670000000
1!
1*
b101 6
19
1>
1C
b101 G
#195680000000
0!
0*
09
0>
0C
#195690000000
1!
1*
b110 6
19
1>
1C
b110 G
#195700000000
0!
0*
09
0>
0C
#195710000000
1!
1*
b111 6
19
1>
1C
b111 G
#195720000000
0!
0*
09
0>
0C
#195730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#195740000000
0!
0*
09
0>
0C
#195750000000
1!
1*
b1 6
19
1>
1C
b1 G
#195760000000
0!
0*
09
0>
0C
#195770000000
1!
1*
b10 6
19
1>
1C
b10 G
#195780000000
0!
0*
09
0>
0C
#195790000000
1!
1*
b11 6
19
1>
1C
b11 G
#195800000000
0!
0*
09
0>
0C
#195810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#195820000000
0!
0*
09
0>
0C
#195830000000
1!
1*
b101 6
19
1>
1C
b101 G
#195840000000
0!
0*
09
0>
0C
#195850000000
1!
1*
b110 6
19
1>
1C
b110 G
#195860000000
0!
0*
09
0>
0C
#195870000000
1!
1*
b111 6
19
1>
1C
b111 G
#195880000000
0!
1"
0*
1+
09
1:
0>
0C
#195890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#195900000000
0!
0*
09
0>
0C
#195910000000
1!
1*
b1 6
19
1>
1C
b1 G
#195920000000
0!
0*
09
0>
0C
#195930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#195940000000
0!
0*
09
0>
0C
#195950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#195960000000
0!
0*
09
0>
0C
#195970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#195980000000
0!
0*
09
0>
0C
#195990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#196000000000
0!
0#
0*
0,
09
0>
0?
0C
#196010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#196020000000
0!
0*
09
0>
0C
#196030000000
1!
1*
19
1>
1C
#196040000000
0!
0*
09
0>
0C
#196050000000
1!
1*
19
1>
1C
#196060000000
0!
0*
09
0>
0C
#196070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#196080000000
0!
0*
09
0>
0C
#196090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#196100000000
0!
0*
09
0>
0C
#196110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#196120000000
0!
0*
09
0>
0C
#196130000000
1!
1*
b10 6
19
1>
1C
b10 G
#196140000000
0!
0*
09
0>
0C
#196150000000
1!
1*
b11 6
19
1>
1C
b11 G
#196160000000
0!
0*
09
0>
0C
#196170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#196180000000
0!
0*
09
0>
0C
#196190000000
1!
1*
b101 6
19
1>
1C
b101 G
#196200000000
0!
0*
09
0>
0C
#196210000000
1!
1*
b110 6
19
1>
1C
b110 G
#196220000000
0!
0*
09
0>
0C
#196230000000
1!
1*
b111 6
19
1>
1C
b111 G
#196240000000
0!
0*
09
0>
0C
#196250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#196260000000
0!
0*
09
0>
0C
#196270000000
1!
1*
b1 6
19
1>
1C
b1 G
#196280000000
0!
0*
09
0>
0C
#196290000000
1!
1*
b10 6
19
1>
1C
b10 G
#196300000000
0!
0*
09
0>
0C
#196310000000
1!
1*
b11 6
19
1>
1C
b11 G
#196320000000
0!
0*
09
0>
0C
#196330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#196340000000
0!
0*
09
0>
0C
#196350000000
1!
1*
b101 6
19
1>
1C
b101 G
#196360000000
0!
0*
09
0>
0C
#196370000000
1!
1*
b110 6
19
1>
1C
b110 G
#196380000000
0!
0*
09
0>
0C
#196390000000
1!
1*
b111 6
19
1>
1C
b111 G
#196400000000
0!
0*
09
0>
0C
#196410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#196420000000
0!
0*
09
0>
0C
#196430000000
1!
1*
b1 6
19
1>
1C
b1 G
#196440000000
0!
0*
09
0>
0C
#196450000000
1!
1*
b10 6
19
1>
1C
b10 G
#196460000000
0!
0*
09
0>
0C
#196470000000
1!
1*
b11 6
19
1>
1C
b11 G
#196480000000
0!
0*
09
0>
0C
#196490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#196500000000
0!
0*
09
0>
0C
#196510000000
1!
1*
b101 6
19
1>
1C
b101 G
#196520000000
0!
0*
09
0>
0C
#196530000000
1!
1*
b110 6
19
1>
1C
b110 G
#196540000000
0!
0*
09
0>
0C
#196550000000
1!
1*
b111 6
19
1>
1C
b111 G
#196560000000
0!
1"
0*
1+
09
1:
0>
0C
#196570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#196580000000
0!
0*
09
0>
0C
#196590000000
1!
1*
b1 6
19
1>
1C
b1 G
#196600000000
0!
0*
09
0>
0C
#196610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#196620000000
0!
0*
09
0>
0C
#196630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#196640000000
0!
0*
09
0>
0C
#196650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#196660000000
0!
0*
09
0>
0C
#196670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#196680000000
0!
0#
0*
0,
09
0>
0?
0C
#196690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#196700000000
0!
0*
09
0>
0C
#196710000000
1!
1*
19
1>
1C
#196720000000
0!
0*
09
0>
0C
#196730000000
1!
1*
19
1>
1C
#196740000000
0!
0*
09
0>
0C
#196750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#196760000000
0!
0*
09
0>
0C
#196770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#196780000000
0!
0*
09
0>
0C
#196790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#196800000000
0!
0*
09
0>
0C
#196810000000
1!
1*
b10 6
19
1>
1C
b10 G
#196820000000
0!
0*
09
0>
0C
#196830000000
1!
1*
b11 6
19
1>
1C
b11 G
#196840000000
0!
0*
09
0>
0C
#196850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#196860000000
0!
0*
09
0>
0C
#196870000000
1!
1*
b101 6
19
1>
1C
b101 G
#196880000000
0!
0*
09
0>
0C
#196890000000
1!
1*
b110 6
19
1>
1C
b110 G
#196900000000
0!
0*
09
0>
0C
#196910000000
1!
1*
b111 6
19
1>
1C
b111 G
#196920000000
0!
0*
09
0>
0C
#196930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#196940000000
0!
0*
09
0>
0C
#196950000000
1!
1*
b1 6
19
1>
1C
b1 G
#196960000000
0!
0*
09
0>
0C
#196970000000
1!
1*
b10 6
19
1>
1C
b10 G
#196980000000
0!
0*
09
0>
0C
#196990000000
1!
1*
b11 6
19
1>
1C
b11 G
#197000000000
0!
0*
09
0>
0C
#197010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#197020000000
0!
0*
09
0>
0C
#197030000000
1!
1*
b101 6
19
1>
1C
b101 G
#197040000000
0!
0*
09
0>
0C
#197050000000
1!
1*
b110 6
19
1>
1C
b110 G
#197060000000
0!
0*
09
0>
0C
#197070000000
1!
1*
b111 6
19
1>
1C
b111 G
#197080000000
0!
0*
09
0>
0C
#197090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#197100000000
0!
0*
09
0>
0C
#197110000000
1!
1*
b1 6
19
1>
1C
b1 G
#197120000000
0!
0*
09
0>
0C
#197130000000
1!
1*
b10 6
19
1>
1C
b10 G
#197140000000
0!
0*
09
0>
0C
#197150000000
1!
1*
b11 6
19
1>
1C
b11 G
#197160000000
0!
0*
09
0>
0C
#197170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#197180000000
0!
0*
09
0>
0C
#197190000000
1!
1*
b101 6
19
1>
1C
b101 G
#197200000000
0!
0*
09
0>
0C
#197210000000
1!
1*
b110 6
19
1>
1C
b110 G
#197220000000
0!
0*
09
0>
0C
#197230000000
1!
1*
b111 6
19
1>
1C
b111 G
#197240000000
0!
1"
0*
1+
09
1:
0>
0C
#197250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#197260000000
0!
0*
09
0>
0C
#197270000000
1!
1*
b1 6
19
1>
1C
b1 G
#197280000000
0!
0*
09
0>
0C
#197290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#197300000000
0!
0*
09
0>
0C
#197310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#197320000000
0!
0*
09
0>
0C
#197330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#197340000000
0!
0*
09
0>
0C
#197350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#197360000000
0!
0#
0*
0,
09
0>
0?
0C
#197370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#197380000000
0!
0*
09
0>
0C
#197390000000
1!
1*
19
1>
1C
#197400000000
0!
0*
09
0>
0C
#197410000000
1!
1*
19
1>
1C
#197420000000
0!
0*
09
0>
0C
#197430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#197440000000
0!
0*
09
0>
0C
#197450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#197460000000
0!
0*
09
0>
0C
#197470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#197480000000
0!
0*
09
0>
0C
#197490000000
1!
1*
b10 6
19
1>
1C
b10 G
#197500000000
0!
0*
09
0>
0C
#197510000000
1!
1*
b11 6
19
1>
1C
b11 G
#197520000000
0!
0*
09
0>
0C
#197530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#197540000000
0!
0*
09
0>
0C
#197550000000
1!
1*
b101 6
19
1>
1C
b101 G
#197560000000
0!
0*
09
0>
0C
#197570000000
1!
1*
b110 6
19
1>
1C
b110 G
#197580000000
0!
0*
09
0>
0C
#197590000000
1!
1*
b111 6
19
1>
1C
b111 G
#197600000000
0!
0*
09
0>
0C
#197610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#197620000000
0!
0*
09
0>
0C
#197630000000
1!
1*
b1 6
19
1>
1C
b1 G
#197640000000
0!
0*
09
0>
0C
#197650000000
1!
1*
b10 6
19
1>
1C
b10 G
#197660000000
0!
0*
09
0>
0C
#197670000000
1!
1*
b11 6
19
1>
1C
b11 G
#197680000000
0!
0*
09
0>
0C
#197690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#197700000000
0!
0*
09
0>
0C
#197710000000
1!
1*
b101 6
19
1>
1C
b101 G
#197720000000
0!
0*
09
0>
0C
#197730000000
1!
1*
b110 6
19
1>
1C
b110 G
#197740000000
0!
0*
09
0>
0C
#197750000000
1!
1*
b111 6
19
1>
1C
b111 G
#197760000000
0!
0*
09
0>
0C
#197770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#197780000000
0!
0*
09
0>
0C
#197790000000
1!
1*
b1 6
19
1>
1C
b1 G
#197800000000
0!
0*
09
0>
0C
#197810000000
1!
1*
b10 6
19
1>
1C
b10 G
#197820000000
0!
0*
09
0>
0C
#197830000000
1!
1*
b11 6
19
1>
1C
b11 G
#197840000000
0!
0*
09
0>
0C
#197850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#197860000000
0!
0*
09
0>
0C
#197870000000
1!
1*
b101 6
19
1>
1C
b101 G
#197880000000
0!
0*
09
0>
0C
#197890000000
1!
1*
b110 6
19
1>
1C
b110 G
#197900000000
0!
0*
09
0>
0C
#197910000000
1!
1*
b111 6
19
1>
1C
b111 G
#197920000000
0!
1"
0*
1+
09
1:
0>
0C
#197930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#197940000000
0!
0*
09
0>
0C
#197950000000
1!
1*
b1 6
19
1>
1C
b1 G
#197960000000
0!
0*
09
0>
0C
#197970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#197980000000
0!
0*
09
0>
0C
#197990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#198000000000
0!
0*
09
0>
0C
#198010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#198020000000
0!
0*
09
0>
0C
#198030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#198040000000
0!
0#
0*
0,
09
0>
0?
0C
#198050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#198060000000
0!
0*
09
0>
0C
#198070000000
1!
1*
19
1>
1C
#198080000000
0!
0*
09
0>
0C
#198090000000
1!
1*
19
1>
1C
#198100000000
0!
0*
09
0>
0C
#198110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#198120000000
0!
0*
09
0>
0C
#198130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#198140000000
0!
0*
09
0>
0C
#198150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#198160000000
0!
0*
09
0>
0C
#198170000000
1!
1*
b10 6
19
1>
1C
b10 G
#198180000000
0!
0*
09
0>
0C
#198190000000
1!
1*
b11 6
19
1>
1C
b11 G
#198200000000
0!
0*
09
0>
0C
#198210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#198220000000
0!
0*
09
0>
0C
#198230000000
1!
1*
b101 6
19
1>
1C
b101 G
#198240000000
0!
0*
09
0>
0C
#198250000000
1!
1*
b110 6
19
1>
1C
b110 G
#198260000000
0!
0*
09
0>
0C
#198270000000
1!
1*
b111 6
19
1>
1C
b111 G
#198280000000
0!
0*
09
0>
0C
#198290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#198300000000
0!
0*
09
0>
0C
#198310000000
1!
1*
b1 6
19
1>
1C
b1 G
#198320000000
0!
0*
09
0>
0C
#198330000000
1!
1*
b10 6
19
1>
1C
b10 G
#198340000000
0!
0*
09
0>
0C
#198350000000
1!
1*
b11 6
19
1>
1C
b11 G
#198360000000
0!
0*
09
0>
0C
#198370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#198380000000
0!
0*
09
0>
0C
#198390000000
1!
1*
b101 6
19
1>
1C
b101 G
#198400000000
0!
0*
09
0>
0C
#198410000000
1!
1*
b110 6
19
1>
1C
b110 G
#198420000000
0!
0*
09
0>
0C
#198430000000
1!
1*
b111 6
19
1>
1C
b111 G
#198440000000
0!
0*
09
0>
0C
#198450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#198460000000
0!
0*
09
0>
0C
#198470000000
1!
1*
b1 6
19
1>
1C
b1 G
#198480000000
0!
0*
09
0>
0C
#198490000000
1!
1*
b10 6
19
1>
1C
b10 G
#198500000000
0!
0*
09
0>
0C
#198510000000
1!
1*
b11 6
19
1>
1C
b11 G
#198520000000
0!
0*
09
0>
0C
#198530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#198540000000
0!
0*
09
0>
0C
#198550000000
1!
1*
b101 6
19
1>
1C
b101 G
#198560000000
0!
0*
09
0>
0C
#198570000000
1!
1*
b110 6
19
1>
1C
b110 G
#198580000000
0!
0*
09
0>
0C
#198590000000
1!
1*
b111 6
19
1>
1C
b111 G
#198600000000
0!
1"
0*
1+
09
1:
0>
0C
#198610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#198620000000
0!
0*
09
0>
0C
#198630000000
1!
1*
b1 6
19
1>
1C
b1 G
#198640000000
0!
0*
09
0>
0C
#198650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#198660000000
0!
0*
09
0>
0C
#198670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#198680000000
0!
0*
09
0>
0C
#198690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#198700000000
0!
0*
09
0>
0C
#198710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#198720000000
0!
0#
0*
0,
09
0>
0?
0C
#198730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#198740000000
0!
0*
09
0>
0C
#198750000000
1!
1*
19
1>
1C
#198760000000
0!
0*
09
0>
0C
#198770000000
1!
1*
19
1>
1C
#198780000000
0!
0*
09
0>
0C
#198790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#198800000000
0!
0*
09
0>
0C
#198810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#198820000000
0!
0*
09
0>
0C
#198830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#198840000000
0!
0*
09
0>
0C
#198850000000
1!
1*
b10 6
19
1>
1C
b10 G
#198860000000
0!
0*
09
0>
0C
#198870000000
1!
1*
b11 6
19
1>
1C
b11 G
#198880000000
0!
0*
09
0>
0C
#198890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#198900000000
0!
0*
09
0>
0C
#198910000000
1!
1*
b101 6
19
1>
1C
b101 G
#198920000000
0!
0*
09
0>
0C
#198930000000
1!
1*
b110 6
19
1>
1C
b110 G
#198940000000
0!
0*
09
0>
0C
#198950000000
1!
1*
b111 6
19
1>
1C
b111 G
#198960000000
0!
0*
09
0>
0C
#198970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#198980000000
0!
0*
09
0>
0C
#198990000000
1!
1*
b1 6
19
1>
1C
b1 G
#199000000000
0!
0*
09
0>
0C
#199010000000
1!
1*
b10 6
19
1>
1C
b10 G
#199020000000
0!
0*
09
0>
0C
#199030000000
1!
1*
b11 6
19
1>
1C
b11 G
#199040000000
0!
0*
09
0>
0C
#199050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#199060000000
0!
0*
09
0>
0C
#199070000000
1!
1*
b101 6
19
1>
1C
b101 G
#199080000000
0!
0*
09
0>
0C
#199090000000
1!
1*
b110 6
19
1>
1C
b110 G
#199100000000
0!
0*
09
0>
0C
#199110000000
1!
1*
b111 6
19
1>
1C
b111 G
#199120000000
0!
0*
09
0>
0C
#199130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#199140000000
0!
0*
09
0>
0C
#199150000000
1!
1*
b1 6
19
1>
1C
b1 G
#199160000000
0!
0*
09
0>
0C
#199170000000
1!
1*
b10 6
19
1>
1C
b10 G
#199180000000
0!
0*
09
0>
0C
#199190000000
1!
1*
b11 6
19
1>
1C
b11 G
#199200000000
0!
0*
09
0>
0C
#199210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#199220000000
0!
0*
09
0>
0C
#199230000000
1!
1*
b101 6
19
1>
1C
b101 G
#199240000000
0!
0*
09
0>
0C
#199250000000
1!
1*
b110 6
19
1>
1C
b110 G
#199260000000
0!
0*
09
0>
0C
#199270000000
1!
1*
b111 6
19
1>
1C
b111 G
#199280000000
0!
1"
0*
1+
09
1:
0>
0C
#199290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#199300000000
0!
0*
09
0>
0C
#199310000000
1!
1*
b1 6
19
1>
1C
b1 G
#199320000000
0!
0*
09
0>
0C
#199330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#199340000000
0!
0*
09
0>
0C
#199350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#199360000000
0!
0*
09
0>
0C
#199370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#199380000000
0!
0*
09
0>
0C
#199390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#199400000000
0!
0#
0*
0,
09
0>
0?
0C
#199410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#199420000000
0!
0*
09
0>
0C
#199430000000
1!
1*
19
1>
1C
#199440000000
0!
0*
09
0>
0C
#199450000000
1!
1*
19
1>
1C
#199460000000
0!
0*
09
0>
0C
#199470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#199480000000
0!
0*
09
0>
0C
#199490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#199500000000
0!
0*
09
0>
0C
#199510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#199520000000
0!
0*
09
0>
0C
#199530000000
1!
1*
b10 6
19
1>
1C
b10 G
#199540000000
0!
0*
09
0>
0C
#199550000000
1!
1*
b11 6
19
1>
1C
b11 G
#199560000000
0!
0*
09
0>
0C
#199570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#199580000000
0!
0*
09
0>
0C
#199590000000
1!
1*
b101 6
19
1>
1C
b101 G
#199600000000
0!
0*
09
0>
0C
#199610000000
1!
1*
b110 6
19
1>
1C
b110 G
#199620000000
0!
0*
09
0>
0C
#199630000000
1!
1*
b111 6
19
1>
1C
b111 G
#199640000000
0!
0*
09
0>
0C
#199650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#199660000000
0!
0*
09
0>
0C
#199670000000
1!
1*
b1 6
19
1>
1C
b1 G
#199680000000
0!
0*
09
0>
0C
#199690000000
1!
1*
b10 6
19
1>
1C
b10 G
#199700000000
0!
0*
09
0>
0C
#199710000000
1!
1*
b11 6
19
1>
1C
b11 G
#199720000000
0!
0*
09
0>
0C
#199730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#199740000000
0!
0*
09
0>
0C
#199750000000
1!
1*
b101 6
19
1>
1C
b101 G
#199760000000
0!
0*
09
0>
0C
#199770000000
1!
1*
b110 6
19
1>
1C
b110 G
#199780000000
0!
0*
09
0>
0C
#199790000000
1!
1*
b111 6
19
1>
1C
b111 G
#199800000000
0!
0*
09
0>
0C
#199810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#199820000000
0!
0*
09
0>
0C
#199830000000
1!
1*
b1 6
19
1>
1C
b1 G
#199840000000
0!
0*
09
0>
0C
#199850000000
1!
1*
b10 6
19
1>
1C
b10 G
#199860000000
0!
0*
09
0>
0C
#199870000000
1!
1*
b11 6
19
1>
1C
b11 G
#199880000000
0!
0*
09
0>
0C
#199890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#199900000000
0!
0*
09
0>
0C
#199910000000
1!
1*
b101 6
19
1>
1C
b101 G
#199920000000
0!
0*
09
0>
0C
#199930000000
1!
1*
b110 6
19
1>
1C
b110 G
#199940000000
0!
0*
09
0>
0C
#199950000000
1!
1*
b111 6
19
1>
1C
b111 G
#199960000000
0!
1"
0*
1+
09
1:
0>
0C
#199970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#199980000000
0!
0*
09
0>
0C
#199990000000
1!
1*
b1 6
19
1>
1C
b1 G
#200000000000
0!
0*
09
0>
0C
#200010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#200020000000
0!
0*
09
0>
0C
#200030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#200040000000
0!
0*
09
0>
0C
#200050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#200060000000
0!
0*
09
0>
0C
#200070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#200080000000
0!
0#
0*
0,
09
0>
0?
0C
#200090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#200100000000
0!
0*
09
0>
0C
#200110000000
1!
1*
19
1>
1C
#200120000000
0!
0*
09
0>
0C
#200130000000
1!
1*
19
1>
1C
#200140000000
0!
0*
09
0>
0C
#200150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#200160000000
0!
0*
09
0>
0C
#200170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#200180000000
0!
0*
09
0>
0C
#200190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#200200000000
0!
0*
09
0>
0C
#200210000000
1!
1*
b10 6
19
1>
1C
b10 G
#200220000000
0!
0*
09
0>
0C
#200230000000
1!
1*
b11 6
19
1>
1C
b11 G
#200240000000
0!
0*
09
0>
0C
#200250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#200260000000
0!
0*
09
0>
0C
#200270000000
1!
1*
b101 6
19
1>
1C
b101 G
#200280000000
0!
0*
09
0>
0C
#200290000000
1!
1*
b110 6
19
1>
1C
b110 G
#200300000000
0!
0*
09
0>
0C
#200310000000
1!
1*
b111 6
19
1>
1C
b111 G
#200320000000
0!
0*
09
0>
0C
#200330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#200340000000
0!
0*
09
0>
0C
#200350000000
1!
1*
b1 6
19
1>
1C
b1 G
#200360000000
0!
0*
09
0>
0C
#200370000000
1!
1*
b10 6
19
1>
1C
b10 G
#200380000000
0!
0*
09
0>
0C
#200390000000
1!
1*
b11 6
19
1>
1C
b11 G
#200400000000
0!
0*
09
0>
0C
#200410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#200420000000
0!
0*
09
0>
0C
#200430000000
1!
1*
b101 6
19
1>
1C
b101 G
#200440000000
0!
0*
09
0>
0C
#200450000000
1!
1*
b110 6
19
1>
1C
b110 G
#200460000000
0!
0*
09
0>
0C
#200470000000
1!
1*
b111 6
19
1>
1C
b111 G
#200480000000
0!
0*
09
0>
0C
#200490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#200500000000
0!
0*
09
0>
0C
#200510000000
1!
1*
b1 6
19
1>
1C
b1 G
#200520000000
0!
0*
09
0>
0C
#200530000000
1!
1*
b10 6
19
1>
1C
b10 G
#200540000000
0!
0*
09
0>
0C
#200550000000
1!
1*
b11 6
19
1>
1C
b11 G
#200560000000
0!
0*
09
0>
0C
#200570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#200580000000
0!
0*
09
0>
0C
#200590000000
1!
1*
b101 6
19
1>
1C
b101 G
#200600000000
0!
0*
09
0>
0C
#200610000000
1!
1*
b110 6
19
1>
1C
b110 G
#200620000000
0!
0*
09
0>
0C
#200630000000
1!
1*
b111 6
19
1>
1C
b111 G
#200640000000
0!
1"
0*
1+
09
1:
0>
0C
#200650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#200660000000
0!
0*
09
0>
0C
#200670000000
1!
1*
b1 6
19
1>
1C
b1 G
#200680000000
0!
0*
09
0>
0C
#200690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#200700000000
0!
0*
09
0>
0C
#200710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#200720000000
0!
0*
09
0>
0C
#200730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#200740000000
0!
0*
09
0>
0C
#200750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#200760000000
0!
0#
0*
0,
09
0>
0?
0C
#200770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#200780000000
0!
0*
09
0>
0C
#200790000000
1!
1*
19
1>
1C
#200800000000
0!
0*
09
0>
0C
#200810000000
1!
1*
19
1>
1C
#200820000000
0!
0*
09
0>
0C
#200830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#200840000000
0!
0*
09
0>
0C
#200850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#200860000000
0!
0*
09
0>
0C
#200870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#200880000000
0!
0*
09
0>
0C
#200890000000
1!
1*
b10 6
19
1>
1C
b10 G
#200900000000
0!
0*
09
0>
0C
#200910000000
1!
1*
b11 6
19
1>
1C
b11 G
#200920000000
0!
0*
09
0>
0C
#200930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#200940000000
0!
0*
09
0>
0C
#200950000000
1!
1*
b101 6
19
1>
1C
b101 G
#200960000000
0!
0*
09
0>
0C
#200970000000
1!
1*
b110 6
19
1>
1C
b110 G
#200980000000
0!
0*
09
0>
0C
#200990000000
1!
1*
b111 6
19
1>
1C
b111 G
#201000000000
0!
0*
09
0>
0C
#201010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#201020000000
0!
0*
09
0>
0C
#201030000000
1!
1*
b1 6
19
1>
1C
b1 G
#201040000000
0!
0*
09
0>
0C
#201050000000
1!
1*
b10 6
19
1>
1C
b10 G
#201060000000
0!
0*
09
0>
0C
#201070000000
1!
1*
b11 6
19
1>
1C
b11 G
#201080000000
0!
0*
09
0>
0C
#201090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#201100000000
0!
0*
09
0>
0C
#201110000000
1!
1*
b101 6
19
1>
1C
b101 G
#201120000000
0!
0*
09
0>
0C
#201130000000
1!
1*
b110 6
19
1>
1C
b110 G
#201140000000
0!
0*
09
0>
0C
#201150000000
1!
1*
b111 6
19
1>
1C
b111 G
#201160000000
0!
0*
09
0>
0C
#201170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#201180000000
0!
0*
09
0>
0C
#201190000000
1!
1*
b1 6
19
1>
1C
b1 G
#201200000000
0!
0*
09
0>
0C
#201210000000
1!
1*
b10 6
19
1>
1C
b10 G
#201220000000
0!
0*
09
0>
0C
#201230000000
1!
1*
b11 6
19
1>
1C
b11 G
#201240000000
0!
0*
09
0>
0C
#201250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#201260000000
0!
0*
09
0>
0C
#201270000000
1!
1*
b101 6
19
1>
1C
b101 G
#201280000000
0!
0*
09
0>
0C
#201290000000
1!
1*
b110 6
19
1>
1C
b110 G
#201300000000
0!
0*
09
0>
0C
#201310000000
1!
1*
b111 6
19
1>
1C
b111 G
#201320000000
0!
1"
0*
1+
09
1:
0>
0C
#201330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#201340000000
0!
0*
09
0>
0C
#201350000000
1!
1*
b1 6
19
1>
1C
b1 G
#201360000000
0!
0*
09
0>
0C
#201370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#201380000000
0!
0*
09
0>
0C
#201390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#201400000000
0!
0*
09
0>
0C
#201410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#201420000000
0!
0*
09
0>
0C
#201430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#201440000000
0!
0#
0*
0,
09
0>
0?
0C
#201450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#201460000000
0!
0*
09
0>
0C
#201470000000
1!
1*
19
1>
1C
#201480000000
0!
0*
09
0>
0C
#201490000000
1!
1*
19
1>
1C
#201500000000
0!
0*
09
0>
0C
#201510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#201520000000
0!
0*
09
0>
0C
#201530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#201540000000
0!
0*
09
0>
0C
#201550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#201560000000
0!
0*
09
0>
0C
#201570000000
1!
1*
b10 6
19
1>
1C
b10 G
#201580000000
0!
0*
09
0>
0C
#201590000000
1!
1*
b11 6
19
1>
1C
b11 G
#201600000000
0!
0*
09
0>
0C
#201610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#201620000000
0!
0*
09
0>
0C
#201630000000
1!
1*
b101 6
19
1>
1C
b101 G
#201640000000
0!
0*
09
0>
0C
#201650000000
1!
1*
b110 6
19
1>
1C
b110 G
#201660000000
0!
0*
09
0>
0C
#201670000000
1!
1*
b111 6
19
1>
1C
b111 G
#201680000000
0!
0*
09
0>
0C
#201690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#201700000000
0!
0*
09
0>
0C
#201710000000
1!
1*
b1 6
19
1>
1C
b1 G
#201720000000
0!
0*
09
0>
0C
#201730000000
1!
1*
b10 6
19
1>
1C
b10 G
#201740000000
0!
0*
09
0>
0C
#201750000000
1!
1*
b11 6
19
1>
1C
b11 G
#201760000000
0!
0*
09
0>
0C
#201770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#201780000000
0!
0*
09
0>
0C
#201790000000
1!
1*
b101 6
19
1>
1C
b101 G
#201800000000
0!
0*
09
0>
0C
#201810000000
1!
1*
b110 6
19
1>
1C
b110 G
#201820000000
0!
0*
09
0>
0C
#201830000000
1!
1*
b111 6
19
1>
1C
b111 G
#201840000000
0!
0*
09
0>
0C
#201850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#201860000000
0!
0*
09
0>
0C
#201870000000
1!
1*
b1 6
19
1>
1C
b1 G
#201880000000
0!
0*
09
0>
0C
#201890000000
1!
1*
b10 6
19
1>
1C
b10 G
#201900000000
0!
0*
09
0>
0C
#201910000000
1!
1*
b11 6
19
1>
1C
b11 G
#201920000000
0!
0*
09
0>
0C
#201930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#201940000000
0!
0*
09
0>
0C
#201950000000
1!
1*
b101 6
19
1>
1C
b101 G
#201960000000
0!
0*
09
0>
0C
#201970000000
1!
1*
b110 6
19
1>
1C
b110 G
#201980000000
0!
0*
09
0>
0C
#201990000000
1!
1*
b111 6
19
1>
1C
b111 G
#202000000000
0!
1"
0*
1+
09
1:
0>
0C
#202010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#202020000000
0!
0*
09
0>
0C
#202030000000
1!
1*
b1 6
19
1>
1C
b1 G
#202040000000
0!
0*
09
0>
0C
#202050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#202060000000
0!
0*
09
0>
0C
#202070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#202080000000
0!
0*
09
0>
0C
#202090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#202100000000
0!
0*
09
0>
0C
#202110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#202120000000
0!
0#
0*
0,
09
0>
0?
0C
#202130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#202140000000
0!
0*
09
0>
0C
#202150000000
1!
1*
19
1>
1C
#202160000000
0!
0*
09
0>
0C
#202170000000
1!
1*
19
1>
1C
#202180000000
0!
0*
09
0>
0C
#202190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#202200000000
0!
0*
09
0>
0C
#202210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#202220000000
0!
0*
09
0>
0C
#202230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#202240000000
0!
0*
09
0>
0C
#202250000000
1!
1*
b10 6
19
1>
1C
b10 G
#202260000000
0!
0*
09
0>
0C
#202270000000
1!
1*
b11 6
19
1>
1C
b11 G
#202280000000
0!
0*
09
0>
0C
#202290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#202300000000
0!
0*
09
0>
0C
#202310000000
1!
1*
b101 6
19
1>
1C
b101 G
#202320000000
0!
0*
09
0>
0C
#202330000000
1!
1*
b110 6
19
1>
1C
b110 G
#202340000000
0!
0*
09
0>
0C
#202350000000
1!
1*
b111 6
19
1>
1C
b111 G
#202360000000
0!
0*
09
0>
0C
#202370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#202380000000
0!
0*
09
0>
0C
#202390000000
1!
1*
b1 6
19
1>
1C
b1 G
#202400000000
0!
0*
09
0>
0C
#202410000000
1!
1*
b10 6
19
1>
1C
b10 G
#202420000000
0!
0*
09
0>
0C
#202430000000
1!
1*
b11 6
19
1>
1C
b11 G
#202440000000
0!
0*
09
0>
0C
#202450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#202460000000
0!
0*
09
0>
0C
#202470000000
1!
1*
b101 6
19
1>
1C
b101 G
#202480000000
0!
0*
09
0>
0C
#202490000000
1!
1*
b110 6
19
1>
1C
b110 G
#202500000000
0!
0*
09
0>
0C
#202510000000
1!
1*
b111 6
19
1>
1C
b111 G
#202520000000
0!
0*
09
0>
0C
#202530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#202540000000
0!
0*
09
0>
0C
#202550000000
1!
1*
b1 6
19
1>
1C
b1 G
#202560000000
0!
0*
09
0>
0C
#202570000000
1!
1*
b10 6
19
1>
1C
b10 G
#202580000000
0!
0*
09
0>
0C
#202590000000
1!
1*
b11 6
19
1>
1C
b11 G
#202600000000
0!
0*
09
0>
0C
#202610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#202620000000
0!
0*
09
0>
0C
#202630000000
1!
1*
b101 6
19
1>
1C
b101 G
#202640000000
0!
0*
09
0>
0C
#202650000000
1!
1*
b110 6
19
1>
1C
b110 G
#202660000000
0!
0*
09
0>
0C
#202670000000
1!
1*
b111 6
19
1>
1C
b111 G
#202680000000
0!
1"
0*
1+
09
1:
0>
0C
#202690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#202700000000
0!
0*
09
0>
0C
#202710000000
1!
1*
b1 6
19
1>
1C
b1 G
#202720000000
0!
0*
09
0>
0C
#202730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#202740000000
0!
0*
09
0>
0C
#202750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#202760000000
0!
0*
09
0>
0C
#202770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#202780000000
0!
0*
09
0>
0C
#202790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#202800000000
0!
0#
0*
0,
09
0>
0?
0C
#202810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#202820000000
0!
0*
09
0>
0C
#202830000000
1!
1*
19
1>
1C
#202840000000
0!
0*
09
0>
0C
#202850000000
1!
1*
19
1>
1C
#202860000000
0!
0*
09
0>
0C
#202870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#202880000000
0!
0*
09
0>
0C
#202890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#202900000000
0!
0*
09
0>
0C
#202910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#202920000000
0!
0*
09
0>
0C
#202930000000
1!
1*
b10 6
19
1>
1C
b10 G
#202940000000
0!
0*
09
0>
0C
#202950000000
1!
1*
b11 6
19
1>
1C
b11 G
#202960000000
0!
0*
09
0>
0C
#202970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#202980000000
0!
0*
09
0>
0C
#202990000000
1!
1*
b101 6
19
1>
1C
b101 G
#203000000000
0!
0*
09
0>
0C
#203010000000
1!
1*
b110 6
19
1>
1C
b110 G
#203020000000
0!
0*
09
0>
0C
#203030000000
1!
1*
b111 6
19
1>
1C
b111 G
#203040000000
0!
0*
09
0>
0C
#203050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#203060000000
0!
0*
09
0>
0C
#203070000000
1!
1*
b1 6
19
1>
1C
b1 G
#203080000000
0!
0*
09
0>
0C
#203090000000
1!
1*
b10 6
19
1>
1C
b10 G
#203100000000
0!
0*
09
0>
0C
#203110000000
1!
1*
b11 6
19
1>
1C
b11 G
#203120000000
0!
0*
09
0>
0C
#203130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#203140000000
0!
0*
09
0>
0C
#203150000000
1!
1*
b101 6
19
1>
1C
b101 G
#203160000000
0!
0*
09
0>
0C
#203170000000
1!
1*
b110 6
19
1>
1C
b110 G
#203180000000
0!
0*
09
0>
0C
#203190000000
1!
1*
b111 6
19
1>
1C
b111 G
#203200000000
0!
0*
09
0>
0C
#203210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#203220000000
0!
0*
09
0>
0C
#203230000000
1!
1*
b1 6
19
1>
1C
b1 G
#203240000000
0!
0*
09
0>
0C
#203250000000
1!
1*
b10 6
19
1>
1C
b10 G
#203260000000
0!
0*
09
0>
0C
#203270000000
1!
1*
b11 6
19
1>
1C
b11 G
#203280000000
0!
0*
09
0>
0C
#203290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#203300000000
0!
0*
09
0>
0C
#203310000000
1!
1*
b101 6
19
1>
1C
b101 G
#203320000000
0!
0*
09
0>
0C
#203330000000
1!
1*
b110 6
19
1>
1C
b110 G
#203340000000
0!
0*
09
0>
0C
#203350000000
1!
1*
b111 6
19
1>
1C
b111 G
#203360000000
0!
1"
0*
1+
09
1:
0>
0C
#203370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#203380000000
0!
0*
09
0>
0C
#203390000000
1!
1*
b1 6
19
1>
1C
b1 G
#203400000000
0!
0*
09
0>
0C
#203410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#203420000000
0!
0*
09
0>
0C
#203430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#203440000000
0!
0*
09
0>
0C
#203450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#203460000000
0!
0*
09
0>
0C
#203470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#203480000000
0!
0#
0*
0,
09
0>
0?
0C
#203490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#203500000000
0!
0*
09
0>
0C
#203510000000
1!
1*
19
1>
1C
#203520000000
0!
0*
09
0>
0C
#203530000000
1!
1*
19
1>
1C
#203540000000
0!
0*
09
0>
0C
#203550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#203560000000
0!
0*
09
0>
0C
#203570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#203580000000
0!
0*
09
0>
0C
#203590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#203600000000
0!
0*
09
0>
0C
#203610000000
1!
1*
b10 6
19
1>
1C
b10 G
#203620000000
0!
0*
09
0>
0C
#203630000000
1!
1*
b11 6
19
1>
1C
b11 G
#203640000000
0!
0*
09
0>
0C
#203650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#203660000000
0!
0*
09
0>
0C
#203670000000
1!
1*
b101 6
19
1>
1C
b101 G
#203680000000
0!
0*
09
0>
0C
#203690000000
1!
1*
b110 6
19
1>
1C
b110 G
#203700000000
0!
0*
09
0>
0C
#203710000000
1!
1*
b111 6
19
1>
1C
b111 G
#203720000000
0!
0*
09
0>
0C
#203730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#203740000000
0!
0*
09
0>
0C
#203750000000
1!
1*
b1 6
19
1>
1C
b1 G
#203760000000
0!
0*
09
0>
0C
#203770000000
1!
1*
b10 6
19
1>
1C
b10 G
#203780000000
0!
0*
09
0>
0C
#203790000000
1!
1*
b11 6
19
1>
1C
b11 G
#203800000000
0!
0*
09
0>
0C
#203810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#203820000000
0!
0*
09
0>
0C
#203830000000
1!
1*
b101 6
19
1>
1C
b101 G
#203840000000
0!
0*
09
0>
0C
#203850000000
1!
1*
b110 6
19
1>
1C
b110 G
#203860000000
0!
0*
09
0>
0C
#203870000000
1!
1*
b111 6
19
1>
1C
b111 G
#203880000000
0!
0*
09
0>
0C
#203890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#203900000000
0!
0*
09
0>
0C
#203910000000
1!
1*
b1 6
19
1>
1C
b1 G
#203920000000
0!
0*
09
0>
0C
#203930000000
1!
1*
b10 6
19
1>
1C
b10 G
#203940000000
0!
0*
09
0>
0C
#203950000000
1!
1*
b11 6
19
1>
1C
b11 G
#203960000000
0!
0*
09
0>
0C
#203970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#203980000000
0!
0*
09
0>
0C
#203990000000
1!
1*
b101 6
19
1>
1C
b101 G
#204000000000
0!
0*
09
0>
0C
#204010000000
1!
1*
b110 6
19
1>
1C
b110 G
#204020000000
0!
0*
09
0>
0C
#204030000000
1!
1*
b111 6
19
1>
1C
b111 G
#204040000000
0!
1"
0*
1+
09
1:
0>
0C
#204050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#204060000000
0!
0*
09
0>
0C
#204070000000
1!
1*
b1 6
19
1>
1C
b1 G
#204080000000
0!
0*
09
0>
0C
#204090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#204100000000
0!
0*
09
0>
0C
#204110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#204120000000
0!
0*
09
0>
0C
#204130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#204140000000
0!
0*
09
0>
0C
#204150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#204160000000
0!
0#
0*
0,
09
0>
0?
0C
#204170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#204180000000
0!
0*
09
0>
0C
#204190000000
1!
1*
19
1>
1C
#204200000000
0!
0*
09
0>
0C
#204210000000
1!
1*
19
1>
1C
#204220000000
0!
0*
09
0>
0C
#204230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#204240000000
0!
0*
09
0>
0C
#204250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#204260000000
0!
0*
09
0>
0C
#204270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#204280000000
0!
0*
09
0>
0C
#204290000000
1!
1*
b10 6
19
1>
1C
b10 G
#204300000000
0!
0*
09
0>
0C
#204310000000
1!
1*
b11 6
19
1>
1C
b11 G
#204320000000
0!
0*
09
0>
0C
#204330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#204340000000
0!
0*
09
0>
0C
#204350000000
1!
1*
b101 6
19
1>
1C
b101 G
#204360000000
0!
0*
09
0>
0C
#204370000000
1!
1*
b110 6
19
1>
1C
b110 G
#204380000000
0!
0*
09
0>
0C
#204390000000
1!
1*
b111 6
19
1>
1C
b111 G
#204400000000
0!
0*
09
0>
0C
#204410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#204420000000
0!
0*
09
0>
0C
#204430000000
1!
1*
b1 6
19
1>
1C
b1 G
#204440000000
0!
0*
09
0>
0C
#204450000000
1!
1*
b10 6
19
1>
1C
b10 G
#204460000000
0!
0*
09
0>
0C
#204470000000
1!
1*
b11 6
19
1>
1C
b11 G
#204480000000
0!
0*
09
0>
0C
#204490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#204500000000
0!
0*
09
0>
0C
#204510000000
1!
1*
b101 6
19
1>
1C
b101 G
#204520000000
0!
0*
09
0>
0C
#204530000000
1!
1*
b110 6
19
1>
1C
b110 G
#204540000000
0!
0*
09
0>
0C
#204550000000
1!
1*
b111 6
19
1>
1C
b111 G
#204560000000
0!
0*
09
0>
0C
#204570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#204580000000
0!
0*
09
0>
0C
#204590000000
1!
1*
b1 6
19
1>
1C
b1 G
#204600000000
0!
0*
09
0>
0C
#204610000000
1!
1*
b10 6
19
1>
1C
b10 G
#204620000000
0!
0*
09
0>
0C
#204630000000
1!
1*
b11 6
19
1>
1C
b11 G
#204640000000
0!
0*
09
0>
0C
#204650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#204660000000
0!
0*
09
0>
0C
#204670000000
1!
1*
b101 6
19
1>
1C
b101 G
#204680000000
0!
0*
09
0>
0C
#204690000000
1!
1*
b110 6
19
1>
1C
b110 G
#204700000000
0!
0*
09
0>
0C
#204710000000
1!
1*
b111 6
19
1>
1C
b111 G
#204720000000
0!
1"
0*
1+
09
1:
0>
0C
#204730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#204740000000
0!
0*
09
0>
0C
#204750000000
1!
1*
b1 6
19
1>
1C
b1 G
#204760000000
0!
0*
09
0>
0C
#204770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#204780000000
0!
0*
09
0>
0C
#204790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#204800000000
0!
0*
09
0>
0C
#204810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#204820000000
0!
0*
09
0>
0C
#204830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#204840000000
0!
0#
0*
0,
09
0>
0?
0C
#204850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#204860000000
0!
0*
09
0>
0C
#204870000000
1!
1*
19
1>
1C
#204880000000
0!
0*
09
0>
0C
#204890000000
1!
1*
19
1>
1C
#204900000000
0!
0*
09
0>
0C
#204910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#204920000000
0!
0*
09
0>
0C
#204930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#204940000000
0!
0*
09
0>
0C
#204950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#204960000000
0!
0*
09
0>
0C
#204970000000
1!
1*
b10 6
19
1>
1C
b10 G
#204980000000
0!
0*
09
0>
0C
#204990000000
1!
1*
b11 6
19
1>
1C
b11 G
#205000000000
0!
0*
09
0>
0C
#205010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#205020000000
0!
0*
09
0>
0C
#205030000000
1!
1*
b101 6
19
1>
1C
b101 G
#205040000000
0!
0*
09
0>
0C
#205050000000
1!
1*
b110 6
19
1>
1C
b110 G
#205060000000
0!
0*
09
0>
0C
#205070000000
1!
1*
b111 6
19
1>
1C
b111 G
#205080000000
0!
0*
09
0>
0C
#205090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#205100000000
0!
0*
09
0>
0C
#205110000000
1!
1*
b1 6
19
1>
1C
b1 G
#205120000000
0!
0*
09
0>
0C
#205130000000
1!
1*
b10 6
19
1>
1C
b10 G
#205140000000
0!
0*
09
0>
0C
#205150000000
1!
1*
b11 6
19
1>
1C
b11 G
#205160000000
0!
0*
09
0>
0C
#205170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#205180000000
0!
0*
09
0>
0C
#205190000000
1!
1*
b101 6
19
1>
1C
b101 G
#205200000000
0!
0*
09
0>
0C
#205210000000
1!
1*
b110 6
19
1>
1C
b110 G
#205220000000
0!
0*
09
0>
0C
#205230000000
1!
1*
b111 6
19
1>
1C
b111 G
#205240000000
0!
0*
09
0>
0C
#205250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#205260000000
0!
0*
09
0>
0C
#205270000000
1!
1*
b1 6
19
1>
1C
b1 G
#205280000000
0!
0*
09
0>
0C
#205290000000
1!
1*
b10 6
19
1>
1C
b10 G
#205300000000
0!
0*
09
0>
0C
#205310000000
1!
1*
b11 6
19
1>
1C
b11 G
#205320000000
0!
0*
09
0>
0C
#205330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#205340000000
0!
0*
09
0>
0C
#205350000000
1!
1*
b101 6
19
1>
1C
b101 G
#205360000000
0!
0*
09
0>
0C
#205370000000
1!
1*
b110 6
19
1>
1C
b110 G
#205380000000
0!
0*
09
0>
0C
#205390000000
1!
1*
b111 6
19
1>
1C
b111 G
#205400000000
0!
1"
0*
1+
09
1:
0>
0C
#205410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#205420000000
0!
0*
09
0>
0C
#205430000000
1!
1*
b1 6
19
1>
1C
b1 G
#205440000000
0!
0*
09
0>
0C
#205450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#205460000000
0!
0*
09
0>
0C
#205470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#205480000000
0!
0*
09
0>
0C
#205490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#205500000000
0!
0*
09
0>
0C
#205510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#205520000000
0!
0#
0*
0,
09
0>
0?
0C
#205530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#205540000000
0!
0*
09
0>
0C
#205550000000
1!
1*
19
1>
1C
#205560000000
0!
0*
09
0>
0C
#205570000000
1!
1*
19
1>
1C
#205580000000
0!
0*
09
0>
0C
#205590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#205600000000
0!
0*
09
0>
0C
#205610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#205620000000
0!
0*
09
0>
0C
#205630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#205640000000
0!
0*
09
0>
0C
#205650000000
1!
1*
b10 6
19
1>
1C
b10 G
#205660000000
0!
0*
09
0>
0C
#205670000000
1!
1*
b11 6
19
1>
1C
b11 G
#205680000000
0!
0*
09
0>
0C
#205690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#205700000000
0!
0*
09
0>
0C
#205710000000
1!
1*
b101 6
19
1>
1C
b101 G
#205720000000
0!
0*
09
0>
0C
#205730000000
1!
1*
b110 6
19
1>
1C
b110 G
#205740000000
0!
0*
09
0>
0C
#205750000000
1!
1*
b111 6
19
1>
1C
b111 G
#205760000000
0!
0*
09
0>
0C
#205770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#205780000000
0!
0*
09
0>
0C
#205790000000
1!
1*
b1 6
19
1>
1C
b1 G
#205800000000
0!
0*
09
0>
0C
#205810000000
1!
1*
b10 6
19
1>
1C
b10 G
#205820000000
0!
0*
09
0>
0C
#205830000000
1!
1*
b11 6
19
1>
1C
b11 G
#205840000000
0!
0*
09
0>
0C
#205850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#205860000000
0!
0*
09
0>
0C
#205870000000
1!
1*
b101 6
19
1>
1C
b101 G
#205880000000
0!
0*
09
0>
0C
#205890000000
1!
1*
b110 6
19
1>
1C
b110 G
#205900000000
0!
0*
09
0>
0C
#205910000000
1!
1*
b111 6
19
1>
1C
b111 G
#205920000000
0!
0*
09
0>
0C
#205930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#205940000000
0!
0*
09
0>
0C
#205950000000
1!
1*
b1 6
19
1>
1C
b1 G
#205960000000
0!
0*
09
0>
0C
#205970000000
1!
1*
b10 6
19
1>
1C
b10 G
#205980000000
0!
0*
09
0>
0C
#205990000000
1!
1*
b11 6
19
1>
1C
b11 G
#206000000000
0!
0*
09
0>
0C
#206010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#206020000000
0!
0*
09
0>
0C
#206030000000
1!
1*
b101 6
19
1>
1C
b101 G
#206040000000
0!
0*
09
0>
0C
#206050000000
1!
1*
b110 6
19
1>
1C
b110 G
#206060000000
0!
0*
09
0>
0C
#206070000000
1!
1*
b111 6
19
1>
1C
b111 G
#206080000000
0!
1"
0*
1+
09
1:
0>
0C
#206090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#206100000000
0!
0*
09
0>
0C
#206110000000
1!
1*
b1 6
19
1>
1C
b1 G
#206120000000
0!
0*
09
0>
0C
#206130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#206140000000
0!
0*
09
0>
0C
#206150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#206160000000
0!
0*
09
0>
0C
#206170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#206180000000
0!
0*
09
0>
0C
#206190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#206200000000
0!
0#
0*
0,
09
0>
0?
0C
#206210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#206220000000
0!
0*
09
0>
0C
#206230000000
1!
1*
19
1>
1C
#206240000000
0!
0*
09
0>
0C
#206250000000
1!
1*
19
1>
1C
#206260000000
0!
0*
09
0>
0C
#206270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#206280000000
0!
0*
09
0>
0C
#206290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#206300000000
0!
0*
09
0>
0C
#206310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#206320000000
0!
0*
09
0>
0C
#206330000000
1!
1*
b10 6
19
1>
1C
b10 G
#206340000000
0!
0*
09
0>
0C
#206350000000
1!
1*
b11 6
19
1>
1C
b11 G
#206360000000
0!
0*
09
0>
0C
#206370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#206380000000
0!
0*
09
0>
0C
#206390000000
1!
1*
b101 6
19
1>
1C
b101 G
#206400000000
0!
0*
09
0>
0C
#206410000000
1!
1*
b110 6
19
1>
1C
b110 G
#206420000000
0!
0*
09
0>
0C
#206430000000
1!
1*
b111 6
19
1>
1C
b111 G
#206440000000
0!
0*
09
0>
0C
#206450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#206460000000
0!
0*
09
0>
0C
#206470000000
1!
1*
b1 6
19
1>
1C
b1 G
#206480000000
0!
0*
09
0>
0C
#206490000000
1!
1*
b10 6
19
1>
1C
b10 G
#206500000000
0!
0*
09
0>
0C
#206510000000
1!
1*
b11 6
19
1>
1C
b11 G
#206520000000
0!
0*
09
0>
0C
#206530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#206540000000
0!
0*
09
0>
0C
#206550000000
1!
1*
b101 6
19
1>
1C
b101 G
#206560000000
0!
0*
09
0>
0C
#206570000000
1!
1*
b110 6
19
1>
1C
b110 G
#206580000000
0!
0*
09
0>
0C
#206590000000
1!
1*
b111 6
19
1>
1C
b111 G
#206600000000
0!
0*
09
0>
0C
#206610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#206620000000
0!
0*
09
0>
0C
#206630000000
1!
1*
b1 6
19
1>
1C
b1 G
#206640000000
0!
0*
09
0>
0C
#206650000000
1!
1*
b10 6
19
1>
1C
b10 G
#206660000000
0!
0*
09
0>
0C
#206670000000
1!
1*
b11 6
19
1>
1C
b11 G
#206680000000
0!
0*
09
0>
0C
#206690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#206700000000
0!
0*
09
0>
0C
#206710000000
1!
1*
b101 6
19
1>
1C
b101 G
#206720000000
0!
0*
09
0>
0C
#206730000000
1!
1*
b110 6
19
1>
1C
b110 G
#206740000000
0!
0*
09
0>
0C
#206750000000
1!
1*
b111 6
19
1>
1C
b111 G
#206760000000
0!
1"
0*
1+
09
1:
0>
0C
#206770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#206780000000
0!
0*
09
0>
0C
#206790000000
1!
1*
b1 6
19
1>
1C
b1 G
#206800000000
0!
0*
09
0>
0C
#206810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#206820000000
0!
0*
09
0>
0C
#206830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#206840000000
0!
0*
09
0>
0C
#206850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#206860000000
0!
0*
09
0>
0C
#206870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#206880000000
0!
0#
0*
0,
09
0>
0?
0C
#206890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#206900000000
0!
0*
09
0>
0C
#206910000000
1!
1*
19
1>
1C
#206920000000
0!
0*
09
0>
0C
#206930000000
1!
1*
19
1>
1C
#206940000000
0!
0*
09
0>
0C
#206950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#206960000000
0!
0*
09
0>
0C
#206970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#206980000000
0!
0*
09
0>
0C
#206990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#207000000000
0!
0*
09
0>
0C
#207010000000
1!
1*
b10 6
19
1>
1C
b10 G
#207020000000
0!
0*
09
0>
0C
#207030000000
1!
1*
b11 6
19
1>
1C
b11 G
#207040000000
0!
0*
09
0>
0C
#207050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#207060000000
0!
0*
09
0>
0C
#207070000000
1!
1*
b101 6
19
1>
1C
b101 G
#207080000000
0!
0*
09
0>
0C
#207090000000
1!
1*
b110 6
19
1>
1C
b110 G
#207100000000
0!
0*
09
0>
0C
#207110000000
1!
1*
b111 6
19
1>
1C
b111 G
#207120000000
0!
0*
09
0>
0C
#207130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#207140000000
0!
0*
09
0>
0C
#207150000000
1!
1*
b1 6
19
1>
1C
b1 G
#207160000000
0!
0*
09
0>
0C
#207170000000
1!
1*
b10 6
19
1>
1C
b10 G
#207180000000
0!
0*
09
0>
0C
#207190000000
1!
1*
b11 6
19
1>
1C
b11 G
#207200000000
0!
0*
09
0>
0C
#207210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#207220000000
0!
0*
09
0>
0C
#207230000000
1!
1*
b101 6
19
1>
1C
b101 G
#207240000000
0!
0*
09
0>
0C
#207250000000
1!
1*
b110 6
19
1>
1C
b110 G
#207260000000
0!
0*
09
0>
0C
#207270000000
1!
1*
b111 6
19
1>
1C
b111 G
#207280000000
0!
0*
09
0>
0C
#207290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#207300000000
0!
0*
09
0>
0C
#207310000000
1!
1*
b1 6
19
1>
1C
b1 G
#207320000000
0!
0*
09
0>
0C
#207330000000
1!
1*
b10 6
19
1>
1C
b10 G
#207340000000
0!
0*
09
0>
0C
#207350000000
1!
1*
b11 6
19
1>
1C
b11 G
#207360000000
0!
0*
09
0>
0C
#207370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#207380000000
0!
0*
09
0>
0C
#207390000000
1!
1*
b101 6
19
1>
1C
b101 G
#207400000000
0!
0*
09
0>
0C
#207410000000
1!
1*
b110 6
19
1>
1C
b110 G
#207420000000
0!
0*
09
0>
0C
#207430000000
1!
1*
b111 6
19
1>
1C
b111 G
#207440000000
0!
1"
0*
1+
09
1:
0>
0C
#207450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#207460000000
0!
0*
09
0>
0C
#207470000000
1!
1*
b1 6
19
1>
1C
b1 G
#207480000000
0!
0*
09
0>
0C
#207490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#207500000000
0!
0*
09
0>
0C
#207510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#207520000000
0!
0*
09
0>
0C
#207530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#207540000000
0!
0*
09
0>
0C
#207550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#207560000000
0!
0#
0*
0,
09
0>
0?
0C
#207570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#207580000000
0!
0*
09
0>
0C
#207590000000
1!
1*
19
1>
1C
#207600000000
0!
0*
09
0>
0C
#207610000000
1!
1*
19
1>
1C
#207620000000
0!
0*
09
0>
0C
#207630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#207640000000
0!
0*
09
0>
0C
#207650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#207660000000
0!
0*
09
0>
0C
#207670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#207680000000
0!
0*
09
0>
0C
#207690000000
1!
1*
b10 6
19
1>
1C
b10 G
#207700000000
0!
0*
09
0>
0C
#207710000000
1!
1*
b11 6
19
1>
1C
b11 G
#207720000000
0!
0*
09
0>
0C
#207730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#207740000000
0!
0*
09
0>
0C
#207750000000
1!
1*
b101 6
19
1>
1C
b101 G
#207760000000
0!
0*
09
0>
0C
#207770000000
1!
1*
b110 6
19
1>
1C
b110 G
#207780000000
0!
0*
09
0>
0C
#207790000000
1!
1*
b111 6
19
1>
1C
b111 G
#207800000000
0!
0*
09
0>
0C
#207810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#207820000000
0!
0*
09
0>
0C
#207830000000
1!
1*
b1 6
19
1>
1C
b1 G
#207840000000
0!
0*
09
0>
0C
#207850000000
1!
1*
b10 6
19
1>
1C
b10 G
#207860000000
0!
0*
09
0>
0C
#207870000000
1!
1*
b11 6
19
1>
1C
b11 G
#207880000000
0!
0*
09
0>
0C
#207890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#207900000000
0!
0*
09
0>
0C
#207910000000
1!
1*
b101 6
19
1>
1C
b101 G
#207920000000
0!
0*
09
0>
0C
#207930000000
1!
1*
b110 6
19
1>
1C
b110 G
#207940000000
0!
0*
09
0>
0C
#207950000000
1!
1*
b111 6
19
1>
1C
b111 G
#207960000000
0!
0*
09
0>
0C
#207970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#207980000000
0!
0*
09
0>
0C
#207990000000
1!
1*
b1 6
19
1>
1C
b1 G
#208000000000
0!
0*
09
0>
0C
#208010000000
1!
1*
b10 6
19
1>
1C
b10 G
#208020000000
0!
0*
09
0>
0C
#208030000000
1!
1*
b11 6
19
1>
1C
b11 G
#208040000000
0!
0*
09
0>
0C
#208050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#208060000000
0!
0*
09
0>
0C
#208070000000
1!
1*
b101 6
19
1>
1C
b101 G
#208080000000
0!
0*
09
0>
0C
#208090000000
1!
1*
b110 6
19
1>
1C
b110 G
#208100000000
0!
0*
09
0>
0C
#208110000000
1!
1*
b111 6
19
1>
1C
b111 G
#208120000000
0!
1"
0*
1+
09
1:
0>
0C
#208130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#208140000000
0!
0*
09
0>
0C
#208150000000
1!
1*
b1 6
19
1>
1C
b1 G
#208160000000
0!
0*
09
0>
0C
#208170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#208180000000
0!
0*
09
0>
0C
#208190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#208200000000
0!
0*
09
0>
0C
#208210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#208220000000
0!
0*
09
0>
0C
#208230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#208240000000
0!
0#
0*
0,
09
0>
0?
0C
#208250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#208260000000
0!
0*
09
0>
0C
#208270000000
1!
1*
19
1>
1C
#208280000000
0!
0*
09
0>
0C
#208290000000
1!
1*
19
1>
1C
#208300000000
0!
0*
09
0>
0C
#208310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#208320000000
0!
0*
09
0>
0C
#208330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#208340000000
0!
0*
09
0>
0C
#208350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#208360000000
0!
0*
09
0>
0C
#208370000000
1!
1*
b10 6
19
1>
1C
b10 G
#208380000000
0!
0*
09
0>
0C
#208390000000
1!
1*
b11 6
19
1>
1C
b11 G
#208400000000
0!
0*
09
0>
0C
#208410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#208420000000
0!
0*
09
0>
0C
#208430000000
1!
1*
b101 6
19
1>
1C
b101 G
#208440000000
0!
0*
09
0>
0C
#208450000000
1!
1*
b110 6
19
1>
1C
b110 G
#208460000000
0!
0*
09
0>
0C
#208470000000
1!
1*
b111 6
19
1>
1C
b111 G
#208480000000
0!
0*
09
0>
0C
#208490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#208500000000
0!
0*
09
0>
0C
#208510000000
1!
1*
b1 6
19
1>
1C
b1 G
#208520000000
0!
0*
09
0>
0C
#208530000000
1!
1*
b10 6
19
1>
1C
b10 G
#208540000000
0!
0*
09
0>
0C
#208550000000
1!
1*
b11 6
19
1>
1C
b11 G
#208560000000
0!
0*
09
0>
0C
#208570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#208580000000
0!
0*
09
0>
0C
#208590000000
1!
1*
b101 6
19
1>
1C
b101 G
#208600000000
0!
0*
09
0>
0C
#208610000000
1!
1*
b110 6
19
1>
1C
b110 G
#208620000000
0!
0*
09
0>
0C
#208630000000
1!
1*
b111 6
19
1>
1C
b111 G
#208640000000
0!
0*
09
0>
0C
#208650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#208660000000
0!
0*
09
0>
0C
#208670000000
1!
1*
b1 6
19
1>
1C
b1 G
#208680000000
0!
0*
09
0>
0C
#208690000000
1!
1*
b10 6
19
1>
1C
b10 G
#208700000000
0!
0*
09
0>
0C
#208710000000
1!
1*
b11 6
19
1>
1C
b11 G
#208720000000
0!
0*
09
0>
0C
#208730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#208740000000
0!
0*
09
0>
0C
#208750000000
1!
1*
b101 6
19
1>
1C
b101 G
#208760000000
0!
0*
09
0>
0C
#208770000000
1!
1*
b110 6
19
1>
1C
b110 G
#208780000000
0!
0*
09
0>
0C
#208790000000
1!
1*
b111 6
19
1>
1C
b111 G
#208800000000
0!
1"
0*
1+
09
1:
0>
0C
#208810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#208820000000
0!
0*
09
0>
0C
#208830000000
1!
1*
b1 6
19
1>
1C
b1 G
#208840000000
0!
0*
09
0>
0C
#208850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#208860000000
0!
0*
09
0>
0C
#208870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#208880000000
0!
0*
09
0>
0C
#208890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#208900000000
0!
0*
09
0>
0C
#208910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#208920000000
0!
0#
0*
0,
09
0>
0?
0C
#208930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#208940000000
0!
0*
09
0>
0C
#208950000000
1!
1*
19
1>
1C
#208960000000
0!
0*
09
0>
0C
#208970000000
1!
1*
19
1>
1C
#208980000000
0!
0*
09
0>
0C
#208990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#209000000000
0!
0*
09
0>
0C
#209010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#209020000000
0!
0*
09
0>
0C
#209030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#209040000000
0!
0*
09
0>
0C
#209050000000
1!
1*
b10 6
19
1>
1C
b10 G
#209060000000
0!
0*
09
0>
0C
#209070000000
1!
1*
b11 6
19
1>
1C
b11 G
#209080000000
0!
0*
09
0>
0C
#209090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#209100000000
0!
0*
09
0>
0C
#209110000000
1!
1*
b101 6
19
1>
1C
b101 G
#209120000000
0!
0*
09
0>
0C
#209130000000
1!
1*
b110 6
19
1>
1C
b110 G
#209140000000
0!
0*
09
0>
0C
#209150000000
1!
1*
b111 6
19
1>
1C
b111 G
#209160000000
0!
0*
09
0>
0C
#209170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#209180000000
0!
0*
09
0>
0C
#209190000000
1!
1*
b1 6
19
1>
1C
b1 G
#209200000000
0!
0*
09
0>
0C
#209210000000
1!
1*
b10 6
19
1>
1C
b10 G
#209220000000
0!
0*
09
0>
0C
#209230000000
1!
1*
b11 6
19
1>
1C
b11 G
#209240000000
0!
0*
09
0>
0C
#209250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#209260000000
0!
0*
09
0>
0C
#209270000000
1!
1*
b101 6
19
1>
1C
b101 G
#209280000000
0!
0*
09
0>
0C
#209290000000
1!
1*
b110 6
19
1>
1C
b110 G
#209300000000
0!
0*
09
0>
0C
#209310000000
1!
1*
b111 6
19
1>
1C
b111 G
#209320000000
0!
0*
09
0>
0C
#209330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#209340000000
0!
0*
09
0>
0C
#209350000000
1!
1*
b1 6
19
1>
1C
b1 G
#209360000000
0!
0*
09
0>
0C
#209370000000
1!
1*
b10 6
19
1>
1C
b10 G
#209380000000
0!
0*
09
0>
0C
#209390000000
1!
1*
b11 6
19
1>
1C
b11 G
#209400000000
0!
0*
09
0>
0C
#209410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#209420000000
0!
0*
09
0>
0C
#209430000000
1!
1*
b101 6
19
1>
1C
b101 G
#209440000000
0!
0*
09
0>
0C
#209450000000
1!
1*
b110 6
19
1>
1C
b110 G
#209460000000
0!
0*
09
0>
0C
#209470000000
1!
1*
b111 6
19
1>
1C
b111 G
#209480000000
0!
1"
0*
1+
09
1:
0>
0C
#209490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#209500000000
0!
0*
09
0>
0C
#209510000000
1!
1*
b1 6
19
1>
1C
b1 G
#209520000000
0!
0*
09
0>
0C
#209530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#209540000000
0!
0*
09
0>
0C
#209550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#209560000000
0!
0*
09
0>
0C
#209570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#209580000000
0!
0*
09
0>
0C
#209590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#209600000000
0!
0#
0*
0,
09
0>
0?
0C
#209610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#209620000000
0!
0*
09
0>
0C
#209630000000
1!
1*
19
1>
1C
#209640000000
0!
0*
09
0>
0C
#209650000000
1!
1*
19
1>
1C
#209660000000
0!
0*
09
0>
0C
#209670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#209680000000
0!
0*
09
0>
0C
#209690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#209700000000
0!
0*
09
0>
0C
#209710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#209720000000
0!
0*
09
0>
0C
#209730000000
1!
1*
b10 6
19
1>
1C
b10 G
#209740000000
0!
0*
09
0>
0C
#209750000000
1!
1*
b11 6
19
1>
1C
b11 G
#209760000000
0!
0*
09
0>
0C
#209770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#209780000000
0!
0*
09
0>
0C
#209790000000
1!
1*
b101 6
19
1>
1C
b101 G
#209800000000
0!
0*
09
0>
0C
#209810000000
1!
1*
b110 6
19
1>
1C
b110 G
#209820000000
0!
0*
09
0>
0C
#209830000000
1!
1*
b111 6
19
1>
1C
b111 G
#209840000000
0!
0*
09
0>
0C
#209850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#209860000000
0!
0*
09
0>
0C
#209870000000
1!
1*
b1 6
19
1>
1C
b1 G
#209880000000
0!
0*
09
0>
0C
#209890000000
1!
1*
b10 6
19
1>
1C
b10 G
#209900000000
0!
0*
09
0>
0C
#209910000000
1!
1*
b11 6
19
1>
1C
b11 G
#209920000000
0!
0*
09
0>
0C
#209930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#209940000000
0!
0*
09
0>
0C
#209950000000
1!
1*
b101 6
19
1>
1C
b101 G
#209960000000
0!
0*
09
0>
0C
#209970000000
1!
1*
b110 6
19
1>
1C
b110 G
#209980000000
0!
0*
09
0>
0C
#209990000000
1!
1*
b111 6
19
1>
1C
b111 G
#210000000000
0!
0*
09
0>
0C
#210010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#210020000000
0!
0*
09
0>
0C
#210030000000
1!
1*
b1 6
19
1>
1C
b1 G
#210040000000
0!
0*
09
0>
0C
#210050000000
1!
1*
b10 6
19
1>
1C
b10 G
#210060000000
0!
0*
09
0>
0C
#210070000000
1!
1*
b11 6
19
1>
1C
b11 G
#210080000000
0!
0*
09
0>
0C
#210090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#210100000000
0!
0*
09
0>
0C
#210110000000
1!
1*
b101 6
19
1>
1C
b101 G
#210120000000
0!
0*
09
0>
0C
#210130000000
1!
1*
b110 6
19
1>
1C
b110 G
#210140000000
0!
0*
09
0>
0C
#210150000000
1!
1*
b111 6
19
1>
1C
b111 G
#210160000000
0!
1"
0*
1+
09
1:
0>
0C
#210170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#210180000000
0!
0*
09
0>
0C
#210190000000
1!
1*
b1 6
19
1>
1C
b1 G
#210200000000
0!
0*
09
0>
0C
#210210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#210220000000
0!
0*
09
0>
0C
#210230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#210240000000
0!
0*
09
0>
0C
#210250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#210260000000
0!
0*
09
0>
0C
#210270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#210280000000
0!
0#
0*
0,
09
0>
0?
0C
#210290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#210300000000
0!
0*
09
0>
0C
#210310000000
1!
1*
19
1>
1C
#210320000000
0!
0*
09
0>
0C
#210330000000
1!
1*
19
1>
1C
#210340000000
0!
0*
09
0>
0C
#210350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#210360000000
0!
0*
09
0>
0C
#210370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#210380000000
0!
0*
09
0>
0C
#210390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#210400000000
0!
0*
09
0>
0C
#210410000000
1!
1*
b10 6
19
1>
1C
b10 G
#210420000000
0!
0*
09
0>
0C
#210430000000
1!
1*
b11 6
19
1>
1C
b11 G
#210440000000
0!
0*
09
0>
0C
#210450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#210460000000
0!
0*
09
0>
0C
#210470000000
1!
1*
b101 6
19
1>
1C
b101 G
#210480000000
0!
0*
09
0>
0C
#210490000000
1!
1*
b110 6
19
1>
1C
b110 G
#210500000000
0!
0*
09
0>
0C
#210510000000
1!
1*
b111 6
19
1>
1C
b111 G
#210520000000
0!
0*
09
0>
0C
#210530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#210540000000
0!
0*
09
0>
0C
#210550000000
1!
1*
b1 6
19
1>
1C
b1 G
#210560000000
0!
0*
09
0>
0C
#210570000000
1!
1*
b10 6
19
1>
1C
b10 G
#210580000000
0!
0*
09
0>
0C
#210590000000
1!
1*
b11 6
19
1>
1C
b11 G
#210600000000
0!
0*
09
0>
0C
#210610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#210620000000
0!
0*
09
0>
0C
#210630000000
1!
1*
b101 6
19
1>
1C
b101 G
#210640000000
0!
0*
09
0>
0C
#210650000000
1!
1*
b110 6
19
1>
1C
b110 G
#210660000000
0!
0*
09
0>
0C
#210670000000
1!
1*
b111 6
19
1>
1C
b111 G
#210680000000
0!
0*
09
0>
0C
#210690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#210700000000
0!
0*
09
0>
0C
#210710000000
1!
1*
b1 6
19
1>
1C
b1 G
#210720000000
0!
0*
09
0>
0C
#210730000000
1!
1*
b10 6
19
1>
1C
b10 G
#210740000000
0!
0*
09
0>
0C
#210750000000
1!
1*
b11 6
19
1>
1C
b11 G
#210760000000
0!
0*
09
0>
0C
#210770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#210780000000
0!
0*
09
0>
0C
#210790000000
1!
1*
b101 6
19
1>
1C
b101 G
#210800000000
0!
0*
09
0>
0C
#210810000000
1!
1*
b110 6
19
1>
1C
b110 G
#210820000000
0!
0*
09
0>
0C
#210830000000
1!
1*
b111 6
19
1>
1C
b111 G
#210840000000
0!
1"
0*
1+
09
1:
0>
0C
#210850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#210860000000
0!
0*
09
0>
0C
#210870000000
1!
1*
b1 6
19
1>
1C
b1 G
#210880000000
0!
0*
09
0>
0C
#210890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#210900000000
0!
0*
09
0>
0C
#210910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#210920000000
0!
0*
09
0>
0C
#210930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#210940000000
0!
0*
09
0>
0C
#210950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#210960000000
0!
0#
0*
0,
09
0>
0?
0C
#210970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#210980000000
0!
0*
09
0>
0C
#210990000000
1!
1*
19
1>
1C
#211000000000
0!
0*
09
0>
0C
#211010000000
1!
1*
19
1>
1C
#211020000000
0!
0*
09
0>
0C
#211030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#211040000000
0!
0*
09
0>
0C
#211050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#211060000000
0!
0*
09
0>
0C
#211070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#211080000000
0!
0*
09
0>
0C
#211090000000
1!
1*
b10 6
19
1>
1C
b10 G
#211100000000
0!
0*
09
0>
0C
#211110000000
1!
1*
b11 6
19
1>
1C
b11 G
#211120000000
0!
0*
09
0>
0C
#211130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#211140000000
0!
0*
09
0>
0C
#211150000000
1!
1*
b101 6
19
1>
1C
b101 G
#211160000000
0!
0*
09
0>
0C
#211170000000
1!
1*
b110 6
19
1>
1C
b110 G
#211180000000
0!
0*
09
0>
0C
#211190000000
1!
1*
b111 6
19
1>
1C
b111 G
#211200000000
0!
0*
09
0>
0C
#211210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#211220000000
0!
0*
09
0>
0C
#211230000000
1!
1*
b1 6
19
1>
1C
b1 G
#211240000000
0!
0*
09
0>
0C
#211250000000
1!
1*
b10 6
19
1>
1C
b10 G
#211260000000
0!
0*
09
0>
0C
#211270000000
1!
1*
b11 6
19
1>
1C
b11 G
#211280000000
0!
0*
09
0>
0C
#211290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#211300000000
0!
0*
09
0>
0C
#211310000000
1!
1*
b101 6
19
1>
1C
b101 G
#211320000000
0!
0*
09
0>
0C
#211330000000
1!
1*
b110 6
19
1>
1C
b110 G
#211340000000
0!
0*
09
0>
0C
#211350000000
1!
1*
b111 6
19
1>
1C
b111 G
#211360000000
0!
0*
09
0>
0C
#211370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#211380000000
0!
0*
09
0>
0C
#211390000000
1!
1*
b1 6
19
1>
1C
b1 G
#211400000000
0!
0*
09
0>
0C
#211410000000
1!
1*
b10 6
19
1>
1C
b10 G
#211420000000
0!
0*
09
0>
0C
#211430000000
1!
1*
b11 6
19
1>
1C
b11 G
#211440000000
0!
0*
09
0>
0C
#211450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#211460000000
0!
0*
09
0>
0C
#211470000000
1!
1*
b101 6
19
1>
1C
b101 G
#211480000000
0!
0*
09
0>
0C
#211490000000
1!
1*
b110 6
19
1>
1C
b110 G
#211500000000
0!
0*
09
0>
0C
#211510000000
1!
1*
b111 6
19
1>
1C
b111 G
#211520000000
0!
1"
0*
1+
09
1:
0>
0C
#211530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#211540000000
0!
0*
09
0>
0C
#211550000000
1!
1*
b1 6
19
1>
1C
b1 G
#211560000000
0!
0*
09
0>
0C
#211570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#211580000000
0!
0*
09
0>
0C
#211590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#211600000000
0!
0*
09
0>
0C
#211610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#211620000000
0!
0*
09
0>
0C
#211630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#211640000000
0!
0#
0*
0,
09
0>
0?
0C
#211650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#211660000000
0!
0*
09
0>
0C
#211670000000
1!
1*
19
1>
1C
#211680000000
0!
0*
09
0>
0C
#211690000000
1!
1*
19
1>
1C
#211700000000
0!
0*
09
0>
0C
#211710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#211720000000
0!
0*
09
0>
0C
#211730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#211740000000
0!
0*
09
0>
0C
#211750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#211760000000
0!
0*
09
0>
0C
#211770000000
1!
1*
b10 6
19
1>
1C
b10 G
#211780000000
0!
0*
09
0>
0C
#211790000000
1!
1*
b11 6
19
1>
1C
b11 G
#211800000000
0!
0*
09
0>
0C
#211810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#211820000000
0!
0*
09
0>
0C
#211830000000
1!
1*
b101 6
19
1>
1C
b101 G
#211840000000
0!
0*
09
0>
0C
#211850000000
1!
1*
b110 6
19
1>
1C
b110 G
#211860000000
0!
0*
09
0>
0C
#211870000000
1!
1*
b111 6
19
1>
1C
b111 G
#211880000000
0!
0*
09
0>
0C
#211890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#211900000000
0!
0*
09
0>
0C
#211910000000
1!
1*
b1 6
19
1>
1C
b1 G
#211920000000
0!
0*
09
0>
0C
#211930000000
1!
1*
b10 6
19
1>
1C
b10 G
#211940000000
0!
0*
09
0>
0C
#211950000000
1!
1*
b11 6
19
1>
1C
b11 G
#211960000000
0!
0*
09
0>
0C
#211970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#211980000000
0!
0*
09
0>
0C
#211990000000
1!
1*
b101 6
19
1>
1C
b101 G
#212000000000
0!
0*
09
0>
0C
#212010000000
1!
1*
b110 6
19
1>
1C
b110 G
#212020000000
0!
0*
09
0>
0C
#212030000000
1!
1*
b111 6
19
1>
1C
b111 G
#212040000000
0!
0*
09
0>
0C
#212050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#212060000000
0!
0*
09
0>
0C
#212070000000
1!
1*
b1 6
19
1>
1C
b1 G
#212080000000
0!
0*
09
0>
0C
#212090000000
1!
1*
b10 6
19
1>
1C
b10 G
#212100000000
0!
0*
09
0>
0C
#212110000000
1!
1*
b11 6
19
1>
1C
b11 G
#212120000000
0!
0*
09
0>
0C
#212130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#212140000000
0!
0*
09
0>
0C
#212150000000
1!
1*
b101 6
19
1>
1C
b101 G
#212160000000
0!
0*
09
0>
0C
#212170000000
1!
1*
b110 6
19
1>
1C
b110 G
#212180000000
0!
0*
09
0>
0C
#212190000000
1!
1*
b111 6
19
1>
1C
b111 G
#212200000000
0!
1"
0*
1+
09
1:
0>
0C
#212210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#212220000000
0!
0*
09
0>
0C
#212230000000
1!
1*
b1 6
19
1>
1C
b1 G
#212240000000
0!
0*
09
0>
0C
#212250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#212260000000
0!
0*
09
0>
0C
#212270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#212280000000
0!
0*
09
0>
0C
#212290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#212300000000
0!
0*
09
0>
0C
#212310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#212320000000
0!
0#
0*
0,
09
0>
0?
0C
#212330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#212340000000
0!
0*
09
0>
0C
#212350000000
1!
1*
19
1>
1C
#212360000000
0!
0*
09
0>
0C
#212370000000
1!
1*
19
1>
1C
#212380000000
0!
0*
09
0>
0C
#212390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#212400000000
0!
0*
09
0>
0C
#212410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#212420000000
0!
0*
09
0>
0C
#212430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#212440000000
0!
0*
09
0>
0C
#212450000000
1!
1*
b10 6
19
1>
1C
b10 G
#212460000000
0!
0*
09
0>
0C
#212470000000
1!
1*
b11 6
19
1>
1C
b11 G
#212480000000
0!
0*
09
0>
0C
#212490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#212500000000
0!
0*
09
0>
0C
#212510000000
1!
1*
b101 6
19
1>
1C
b101 G
#212520000000
0!
0*
09
0>
0C
#212530000000
1!
1*
b110 6
19
1>
1C
b110 G
#212540000000
0!
0*
09
0>
0C
#212550000000
1!
1*
b111 6
19
1>
1C
b111 G
#212560000000
0!
0*
09
0>
0C
#212570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#212580000000
0!
0*
09
0>
0C
#212590000000
1!
1*
b1 6
19
1>
1C
b1 G
#212600000000
0!
0*
09
0>
0C
#212610000000
1!
1*
b10 6
19
1>
1C
b10 G
#212620000000
0!
0*
09
0>
0C
#212630000000
1!
1*
b11 6
19
1>
1C
b11 G
#212640000000
0!
0*
09
0>
0C
#212650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#212660000000
0!
0*
09
0>
0C
#212670000000
1!
1*
b101 6
19
1>
1C
b101 G
#212680000000
0!
0*
09
0>
0C
#212690000000
1!
1*
b110 6
19
1>
1C
b110 G
#212700000000
0!
0*
09
0>
0C
#212710000000
1!
1*
b111 6
19
1>
1C
b111 G
#212720000000
0!
0*
09
0>
0C
#212730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#212740000000
0!
0*
09
0>
0C
#212750000000
1!
1*
b1 6
19
1>
1C
b1 G
#212760000000
0!
0*
09
0>
0C
#212770000000
1!
1*
b10 6
19
1>
1C
b10 G
#212780000000
0!
0*
09
0>
0C
#212790000000
1!
1*
b11 6
19
1>
1C
b11 G
#212800000000
0!
0*
09
0>
0C
#212810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#212820000000
0!
0*
09
0>
0C
#212830000000
1!
1*
b101 6
19
1>
1C
b101 G
#212840000000
0!
0*
09
0>
0C
#212850000000
1!
1*
b110 6
19
1>
1C
b110 G
#212860000000
0!
0*
09
0>
0C
#212870000000
1!
1*
b111 6
19
1>
1C
b111 G
#212880000000
0!
1"
0*
1+
09
1:
0>
0C
#212890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#212900000000
0!
0*
09
0>
0C
#212910000000
1!
1*
b1 6
19
1>
1C
b1 G
#212920000000
0!
0*
09
0>
0C
#212930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#212940000000
0!
0*
09
0>
0C
#212950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#212960000000
0!
0*
09
0>
0C
#212970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#212980000000
0!
0*
09
0>
0C
#212990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#213000000000
0!
0#
0*
0,
09
0>
0?
0C
#213010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#213020000000
0!
0*
09
0>
0C
#213030000000
1!
1*
19
1>
1C
#213040000000
0!
0*
09
0>
0C
#213050000000
1!
1*
19
1>
1C
#213060000000
0!
0*
09
0>
0C
#213070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#213080000000
0!
0*
09
0>
0C
#213090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#213100000000
0!
0*
09
0>
0C
#213110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#213120000000
0!
0*
09
0>
0C
#213130000000
1!
1*
b10 6
19
1>
1C
b10 G
#213140000000
0!
0*
09
0>
0C
#213150000000
1!
1*
b11 6
19
1>
1C
b11 G
#213160000000
0!
0*
09
0>
0C
#213170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#213180000000
0!
0*
09
0>
0C
#213190000000
1!
1*
b101 6
19
1>
1C
b101 G
#213200000000
0!
0*
09
0>
0C
#213210000000
1!
1*
b110 6
19
1>
1C
b110 G
#213220000000
0!
0*
09
0>
0C
#213230000000
1!
1*
b111 6
19
1>
1C
b111 G
#213240000000
0!
0*
09
0>
0C
#213250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#213260000000
0!
0*
09
0>
0C
#213270000000
1!
1*
b1 6
19
1>
1C
b1 G
#213280000000
0!
0*
09
0>
0C
#213290000000
1!
1*
b10 6
19
1>
1C
b10 G
#213300000000
0!
0*
09
0>
0C
#213310000000
1!
1*
b11 6
19
1>
1C
b11 G
#213320000000
0!
0*
09
0>
0C
#213330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#213340000000
0!
0*
09
0>
0C
#213350000000
1!
1*
b101 6
19
1>
1C
b101 G
#213360000000
0!
0*
09
0>
0C
#213370000000
1!
1*
b110 6
19
1>
1C
b110 G
#213380000000
0!
0*
09
0>
0C
#213390000000
1!
1*
b111 6
19
1>
1C
b111 G
#213400000000
0!
0*
09
0>
0C
#213410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#213420000000
0!
0*
09
0>
0C
#213430000000
1!
1*
b1 6
19
1>
1C
b1 G
#213440000000
0!
0*
09
0>
0C
#213450000000
1!
1*
b10 6
19
1>
1C
b10 G
#213460000000
0!
0*
09
0>
0C
#213470000000
1!
1*
b11 6
19
1>
1C
b11 G
#213480000000
0!
0*
09
0>
0C
#213490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#213500000000
0!
0*
09
0>
0C
#213510000000
1!
1*
b101 6
19
1>
1C
b101 G
#213520000000
0!
0*
09
0>
0C
#213530000000
1!
1*
b110 6
19
1>
1C
b110 G
#213540000000
0!
0*
09
0>
0C
#213550000000
1!
1*
b111 6
19
1>
1C
b111 G
#213560000000
0!
1"
0*
1+
09
1:
0>
0C
#213570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#213580000000
0!
0*
09
0>
0C
#213590000000
1!
1*
b1 6
19
1>
1C
b1 G
#213600000000
0!
0*
09
0>
0C
#213610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#213620000000
0!
0*
09
0>
0C
#213630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#213640000000
0!
0*
09
0>
0C
#213650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#213660000000
0!
0*
09
0>
0C
#213670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#213680000000
0!
0#
0*
0,
09
0>
0?
0C
#213690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#213700000000
0!
0*
09
0>
0C
#213710000000
1!
1*
19
1>
1C
#213720000000
0!
0*
09
0>
0C
#213730000000
1!
1*
19
1>
1C
#213740000000
0!
0*
09
0>
0C
#213750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#213760000000
0!
0*
09
0>
0C
#213770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#213780000000
0!
0*
09
0>
0C
#213790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#213800000000
0!
0*
09
0>
0C
#213810000000
1!
1*
b10 6
19
1>
1C
b10 G
#213820000000
0!
0*
09
0>
0C
#213830000000
1!
1*
b11 6
19
1>
1C
b11 G
#213840000000
0!
0*
09
0>
0C
#213850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#213860000000
0!
0*
09
0>
0C
#213870000000
1!
1*
b101 6
19
1>
1C
b101 G
#213880000000
0!
0*
09
0>
0C
#213890000000
1!
1*
b110 6
19
1>
1C
b110 G
#213900000000
0!
0*
09
0>
0C
#213910000000
1!
1*
b111 6
19
1>
1C
b111 G
#213920000000
0!
0*
09
0>
0C
#213930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#213940000000
0!
0*
09
0>
0C
#213950000000
1!
1*
b1 6
19
1>
1C
b1 G
#213960000000
0!
0*
09
0>
0C
#213970000000
1!
1*
b10 6
19
1>
1C
b10 G
#213980000000
0!
0*
09
0>
0C
#213990000000
1!
1*
b11 6
19
1>
1C
b11 G
#214000000000
0!
0*
09
0>
0C
#214010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#214020000000
0!
0*
09
0>
0C
#214030000000
1!
1*
b101 6
19
1>
1C
b101 G
#214040000000
0!
0*
09
0>
0C
#214050000000
1!
1*
b110 6
19
1>
1C
b110 G
#214060000000
0!
0*
09
0>
0C
#214070000000
1!
1*
b111 6
19
1>
1C
b111 G
#214080000000
0!
0*
09
0>
0C
#214090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#214100000000
0!
0*
09
0>
0C
#214110000000
1!
1*
b1 6
19
1>
1C
b1 G
#214120000000
0!
0*
09
0>
0C
#214130000000
1!
1*
b10 6
19
1>
1C
b10 G
#214140000000
0!
0*
09
0>
0C
#214150000000
1!
1*
b11 6
19
1>
1C
b11 G
#214160000000
0!
0*
09
0>
0C
#214170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#214180000000
0!
0*
09
0>
0C
#214190000000
1!
1*
b101 6
19
1>
1C
b101 G
#214200000000
0!
0*
09
0>
0C
#214210000000
1!
1*
b110 6
19
1>
1C
b110 G
#214220000000
0!
0*
09
0>
0C
#214230000000
1!
1*
b111 6
19
1>
1C
b111 G
#214240000000
0!
1"
0*
1+
09
1:
0>
0C
#214250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#214260000000
0!
0*
09
0>
0C
#214270000000
1!
1*
b1 6
19
1>
1C
b1 G
#214280000000
0!
0*
09
0>
0C
#214290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#214300000000
0!
0*
09
0>
0C
#214310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#214320000000
0!
0*
09
0>
0C
#214330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#214340000000
0!
0*
09
0>
0C
#214350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#214360000000
0!
0#
0*
0,
09
0>
0?
0C
#214370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#214380000000
0!
0*
09
0>
0C
#214390000000
1!
1*
19
1>
1C
#214400000000
0!
0*
09
0>
0C
#214410000000
1!
1*
19
1>
1C
#214420000000
0!
0*
09
0>
0C
#214430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#214440000000
0!
0*
09
0>
0C
#214450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#214460000000
0!
0*
09
0>
0C
#214470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#214480000000
0!
0*
09
0>
0C
#214490000000
1!
1*
b10 6
19
1>
1C
b10 G
#214500000000
0!
0*
09
0>
0C
#214510000000
1!
1*
b11 6
19
1>
1C
b11 G
#214520000000
0!
0*
09
0>
0C
#214530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#214540000000
0!
0*
09
0>
0C
#214550000000
1!
1*
b101 6
19
1>
1C
b101 G
#214560000000
0!
0*
09
0>
0C
#214570000000
1!
1*
b110 6
19
1>
1C
b110 G
#214580000000
0!
0*
09
0>
0C
#214590000000
1!
1*
b111 6
19
1>
1C
b111 G
#214600000000
0!
0*
09
0>
0C
#214610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#214620000000
0!
0*
09
0>
0C
#214630000000
1!
1*
b1 6
19
1>
1C
b1 G
#214640000000
0!
0*
09
0>
0C
#214650000000
1!
1*
b10 6
19
1>
1C
b10 G
#214660000000
0!
0*
09
0>
0C
#214670000000
1!
1*
b11 6
19
1>
1C
b11 G
#214680000000
0!
0*
09
0>
0C
#214690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#214700000000
0!
0*
09
0>
0C
#214710000000
1!
1*
b101 6
19
1>
1C
b101 G
#214720000000
0!
0*
09
0>
0C
#214730000000
1!
1*
b110 6
19
1>
1C
b110 G
#214740000000
0!
0*
09
0>
0C
#214750000000
1!
1*
b111 6
19
1>
1C
b111 G
#214760000000
0!
0*
09
0>
0C
#214770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#214780000000
0!
0*
09
0>
0C
#214790000000
1!
1*
b1 6
19
1>
1C
b1 G
#214800000000
0!
0*
09
0>
0C
#214810000000
1!
1*
b10 6
19
1>
1C
b10 G
#214820000000
0!
0*
09
0>
0C
#214830000000
1!
1*
b11 6
19
1>
1C
b11 G
#214840000000
0!
0*
09
0>
0C
#214850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#214860000000
0!
0*
09
0>
0C
#214870000000
1!
1*
b101 6
19
1>
1C
b101 G
#214880000000
0!
0*
09
0>
0C
#214890000000
1!
1*
b110 6
19
1>
1C
b110 G
#214900000000
0!
0*
09
0>
0C
#214910000000
1!
1*
b111 6
19
1>
1C
b111 G
#214920000000
0!
1"
0*
1+
09
1:
0>
0C
#214930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#214940000000
0!
0*
09
0>
0C
#214950000000
1!
1*
b1 6
19
1>
1C
b1 G
#214960000000
0!
0*
09
0>
0C
#214970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#214980000000
0!
0*
09
0>
0C
#214990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#215000000000
0!
0*
09
0>
0C
#215010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#215020000000
0!
0*
09
0>
0C
#215030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#215040000000
0!
0#
0*
0,
09
0>
0?
0C
#215050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#215060000000
0!
0*
09
0>
0C
#215070000000
1!
1*
19
1>
1C
#215080000000
0!
0*
09
0>
0C
#215090000000
1!
1*
19
1>
1C
#215100000000
0!
0*
09
0>
0C
#215110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#215120000000
0!
0*
09
0>
0C
#215130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#215140000000
0!
0*
09
0>
0C
#215150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#215160000000
0!
0*
09
0>
0C
#215170000000
1!
1*
b10 6
19
1>
1C
b10 G
#215180000000
0!
0*
09
0>
0C
#215190000000
1!
1*
b11 6
19
1>
1C
b11 G
#215200000000
0!
0*
09
0>
0C
#215210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#215220000000
0!
0*
09
0>
0C
#215230000000
1!
1*
b101 6
19
1>
1C
b101 G
#215240000000
0!
0*
09
0>
0C
#215250000000
1!
1*
b110 6
19
1>
1C
b110 G
#215260000000
0!
0*
09
0>
0C
#215270000000
1!
1*
b111 6
19
1>
1C
b111 G
#215280000000
0!
0*
09
0>
0C
#215290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#215300000000
0!
0*
09
0>
0C
#215310000000
1!
1*
b1 6
19
1>
1C
b1 G
#215320000000
0!
0*
09
0>
0C
#215330000000
1!
1*
b10 6
19
1>
1C
b10 G
#215340000000
0!
0*
09
0>
0C
#215350000000
1!
1*
b11 6
19
1>
1C
b11 G
#215360000000
0!
0*
09
0>
0C
#215370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#215380000000
0!
0*
09
0>
0C
#215390000000
1!
1*
b101 6
19
1>
1C
b101 G
#215400000000
0!
0*
09
0>
0C
#215410000000
1!
1*
b110 6
19
1>
1C
b110 G
#215420000000
0!
0*
09
0>
0C
#215430000000
1!
1*
b111 6
19
1>
1C
b111 G
#215440000000
0!
0*
09
0>
0C
#215450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#215460000000
0!
0*
09
0>
0C
#215470000000
1!
1*
b1 6
19
1>
1C
b1 G
#215480000000
0!
0*
09
0>
0C
#215490000000
1!
1*
b10 6
19
1>
1C
b10 G
#215500000000
0!
0*
09
0>
0C
#215510000000
1!
1*
b11 6
19
1>
1C
b11 G
#215520000000
0!
0*
09
0>
0C
#215530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#215540000000
0!
0*
09
0>
0C
#215550000000
1!
1*
b101 6
19
1>
1C
b101 G
#215560000000
0!
0*
09
0>
0C
#215570000000
1!
1*
b110 6
19
1>
1C
b110 G
#215580000000
0!
0*
09
0>
0C
#215590000000
1!
1*
b111 6
19
1>
1C
b111 G
#215600000000
0!
1"
0*
1+
09
1:
0>
0C
#215610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#215620000000
0!
0*
09
0>
0C
#215630000000
1!
1*
b1 6
19
1>
1C
b1 G
#215640000000
0!
0*
09
0>
0C
#215650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#215660000000
0!
0*
09
0>
0C
#215670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#215680000000
0!
0*
09
0>
0C
#215690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#215700000000
0!
0*
09
0>
0C
#215710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#215720000000
0!
0#
0*
0,
09
0>
0?
0C
#215730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#215740000000
0!
0*
09
0>
0C
#215750000000
1!
1*
19
1>
1C
#215760000000
0!
0*
09
0>
0C
#215770000000
1!
1*
19
1>
1C
#215780000000
0!
0*
09
0>
0C
#215790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#215800000000
0!
0*
09
0>
0C
#215810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#215820000000
0!
0*
09
0>
0C
#215830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#215840000000
0!
0*
09
0>
0C
#215850000000
1!
1*
b10 6
19
1>
1C
b10 G
#215860000000
0!
0*
09
0>
0C
#215870000000
1!
1*
b11 6
19
1>
1C
b11 G
#215880000000
0!
0*
09
0>
0C
#215890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#215900000000
0!
0*
09
0>
0C
#215910000000
1!
1*
b101 6
19
1>
1C
b101 G
#215920000000
0!
0*
09
0>
0C
#215930000000
1!
1*
b110 6
19
1>
1C
b110 G
#215940000000
0!
0*
09
0>
0C
#215950000000
1!
1*
b111 6
19
1>
1C
b111 G
#215960000000
0!
0*
09
0>
0C
#215970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#215980000000
0!
0*
09
0>
0C
#215990000000
1!
1*
b1 6
19
1>
1C
b1 G
#216000000000
0!
0*
09
0>
0C
#216010000000
1!
1*
b10 6
19
1>
1C
b10 G
#216020000000
0!
0*
09
0>
0C
#216030000000
1!
1*
b11 6
19
1>
1C
b11 G
#216040000000
0!
0*
09
0>
0C
#216050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#216060000000
0!
0*
09
0>
0C
#216070000000
1!
1*
b101 6
19
1>
1C
b101 G
#216080000000
0!
0*
09
0>
0C
#216090000000
1!
1*
b110 6
19
1>
1C
b110 G
#216100000000
0!
0*
09
0>
0C
#216110000000
1!
1*
b111 6
19
1>
1C
b111 G
#216120000000
0!
0*
09
0>
0C
#216130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#216140000000
0!
0*
09
0>
0C
#216150000000
1!
1*
b1 6
19
1>
1C
b1 G
#216160000000
0!
0*
09
0>
0C
#216170000000
1!
1*
b10 6
19
1>
1C
b10 G
#216180000000
0!
0*
09
0>
0C
#216190000000
1!
1*
b11 6
19
1>
1C
b11 G
#216200000000
0!
0*
09
0>
0C
#216210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#216220000000
0!
0*
09
0>
0C
#216230000000
1!
1*
b101 6
19
1>
1C
b101 G
#216240000000
0!
0*
09
0>
0C
#216250000000
1!
1*
b110 6
19
1>
1C
b110 G
#216260000000
0!
0*
09
0>
0C
#216270000000
1!
1*
b111 6
19
1>
1C
b111 G
#216280000000
0!
1"
0*
1+
09
1:
0>
0C
#216290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#216300000000
0!
0*
09
0>
0C
#216310000000
1!
1*
b1 6
19
1>
1C
b1 G
#216320000000
0!
0*
09
0>
0C
#216330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#216340000000
0!
0*
09
0>
0C
#216350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#216360000000
0!
0*
09
0>
0C
#216370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#216380000000
0!
0*
09
0>
0C
#216390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#216400000000
0!
0#
0*
0,
09
0>
0?
0C
#216410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#216420000000
0!
0*
09
0>
0C
#216430000000
1!
1*
19
1>
1C
#216440000000
0!
0*
09
0>
0C
#216450000000
1!
1*
19
1>
1C
#216460000000
0!
0*
09
0>
0C
#216470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#216480000000
0!
0*
09
0>
0C
#216490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#216500000000
0!
0*
09
0>
0C
#216510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#216520000000
0!
0*
09
0>
0C
#216530000000
1!
1*
b10 6
19
1>
1C
b10 G
#216540000000
0!
0*
09
0>
0C
#216550000000
1!
1*
b11 6
19
1>
1C
b11 G
#216560000000
0!
0*
09
0>
0C
#216570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#216580000000
0!
0*
09
0>
0C
#216590000000
1!
1*
b101 6
19
1>
1C
b101 G
#216600000000
0!
0*
09
0>
0C
#216610000000
1!
1*
b110 6
19
1>
1C
b110 G
#216620000000
0!
0*
09
0>
0C
#216630000000
1!
1*
b111 6
19
1>
1C
b111 G
#216640000000
0!
0*
09
0>
0C
#216650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#216660000000
0!
0*
09
0>
0C
#216670000000
1!
1*
b1 6
19
1>
1C
b1 G
#216680000000
0!
0*
09
0>
0C
#216690000000
1!
1*
b10 6
19
1>
1C
b10 G
#216700000000
0!
0*
09
0>
0C
#216710000000
1!
1*
b11 6
19
1>
1C
b11 G
#216720000000
0!
0*
09
0>
0C
#216730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#216740000000
0!
0*
09
0>
0C
#216750000000
1!
1*
b101 6
19
1>
1C
b101 G
#216760000000
0!
0*
09
0>
0C
#216770000000
1!
1*
b110 6
19
1>
1C
b110 G
#216780000000
0!
0*
09
0>
0C
#216790000000
1!
1*
b111 6
19
1>
1C
b111 G
#216800000000
0!
0*
09
0>
0C
#216810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#216820000000
0!
0*
09
0>
0C
#216830000000
1!
1*
b1 6
19
1>
1C
b1 G
#216840000000
0!
0*
09
0>
0C
#216850000000
1!
1*
b10 6
19
1>
1C
b10 G
#216860000000
0!
0*
09
0>
0C
#216870000000
1!
1*
b11 6
19
1>
1C
b11 G
#216880000000
0!
0*
09
0>
0C
#216890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#216900000000
0!
0*
09
0>
0C
#216910000000
1!
1*
b101 6
19
1>
1C
b101 G
#216920000000
0!
0*
09
0>
0C
#216930000000
1!
1*
b110 6
19
1>
1C
b110 G
#216940000000
0!
0*
09
0>
0C
#216950000000
1!
1*
b111 6
19
1>
1C
b111 G
#216960000000
0!
1"
0*
1+
09
1:
0>
0C
#216970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#216980000000
0!
0*
09
0>
0C
#216990000000
1!
1*
b1 6
19
1>
1C
b1 G
#217000000000
0!
0*
09
0>
0C
#217010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#217020000000
0!
0*
09
0>
0C
#217030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#217040000000
0!
0*
09
0>
0C
#217050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#217060000000
0!
0*
09
0>
0C
#217070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#217080000000
0!
0#
0*
0,
09
0>
0?
0C
#217090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#217100000000
0!
0*
09
0>
0C
#217110000000
1!
1*
19
1>
1C
#217120000000
0!
0*
09
0>
0C
#217130000000
1!
1*
19
1>
1C
#217140000000
0!
0*
09
0>
0C
#217150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#217160000000
0!
0*
09
0>
0C
#217170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#217180000000
0!
0*
09
0>
0C
#217190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#217200000000
0!
0*
09
0>
0C
#217210000000
1!
1*
b10 6
19
1>
1C
b10 G
#217220000000
0!
0*
09
0>
0C
#217230000000
1!
1*
b11 6
19
1>
1C
b11 G
#217240000000
0!
0*
09
0>
0C
#217250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#217260000000
0!
0*
09
0>
0C
#217270000000
1!
1*
b101 6
19
1>
1C
b101 G
#217280000000
0!
0*
09
0>
0C
#217290000000
1!
1*
b110 6
19
1>
1C
b110 G
#217300000000
0!
0*
09
0>
0C
#217310000000
1!
1*
b111 6
19
1>
1C
b111 G
#217320000000
0!
0*
09
0>
0C
#217330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#217340000000
0!
0*
09
0>
0C
#217350000000
1!
1*
b1 6
19
1>
1C
b1 G
#217360000000
0!
0*
09
0>
0C
#217370000000
1!
1*
b10 6
19
1>
1C
b10 G
#217380000000
0!
0*
09
0>
0C
#217390000000
1!
1*
b11 6
19
1>
1C
b11 G
#217400000000
0!
0*
09
0>
0C
#217410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#217420000000
0!
0*
09
0>
0C
#217430000000
1!
1*
b101 6
19
1>
1C
b101 G
#217440000000
0!
0*
09
0>
0C
#217450000000
1!
1*
b110 6
19
1>
1C
b110 G
#217460000000
0!
0*
09
0>
0C
#217470000000
1!
1*
b111 6
19
1>
1C
b111 G
#217480000000
0!
0*
09
0>
0C
#217490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#217500000000
0!
0*
09
0>
0C
#217510000000
1!
1*
b1 6
19
1>
1C
b1 G
#217520000000
0!
0*
09
0>
0C
#217530000000
1!
1*
b10 6
19
1>
1C
b10 G
#217540000000
0!
0*
09
0>
0C
#217550000000
1!
1*
b11 6
19
1>
1C
b11 G
#217560000000
0!
0*
09
0>
0C
#217570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#217580000000
0!
0*
09
0>
0C
#217590000000
1!
1*
b101 6
19
1>
1C
b101 G
#217600000000
0!
0*
09
0>
0C
#217610000000
1!
1*
b110 6
19
1>
1C
b110 G
#217620000000
0!
0*
09
0>
0C
#217630000000
1!
1*
b111 6
19
1>
1C
b111 G
#217640000000
0!
1"
0*
1+
09
1:
0>
0C
#217650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#217660000000
0!
0*
09
0>
0C
#217670000000
1!
1*
b1 6
19
1>
1C
b1 G
#217680000000
0!
0*
09
0>
0C
#217690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#217700000000
0!
0*
09
0>
0C
#217710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#217720000000
0!
0*
09
0>
0C
#217730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#217740000000
0!
0*
09
0>
0C
#217750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#217760000000
0!
0#
0*
0,
09
0>
0?
0C
#217770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#217780000000
0!
0*
09
0>
0C
#217790000000
1!
1*
19
1>
1C
#217800000000
0!
0*
09
0>
0C
#217810000000
1!
1*
19
1>
1C
#217820000000
0!
0*
09
0>
0C
#217830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#217840000000
0!
0*
09
0>
0C
#217850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#217860000000
0!
0*
09
0>
0C
#217870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#217880000000
0!
0*
09
0>
0C
#217890000000
1!
1*
b10 6
19
1>
1C
b10 G
#217900000000
0!
0*
09
0>
0C
#217910000000
1!
1*
b11 6
19
1>
1C
b11 G
#217920000000
0!
0*
09
0>
0C
#217930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#217940000000
0!
0*
09
0>
0C
#217950000000
1!
1*
b101 6
19
1>
1C
b101 G
#217960000000
0!
0*
09
0>
0C
#217970000000
1!
1*
b110 6
19
1>
1C
b110 G
#217980000000
0!
0*
09
0>
0C
#217990000000
1!
1*
b111 6
19
1>
1C
b111 G
#218000000000
0!
0*
09
0>
0C
#218010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#218020000000
0!
0*
09
0>
0C
#218030000000
1!
1*
b1 6
19
1>
1C
b1 G
#218040000000
0!
0*
09
0>
0C
#218050000000
1!
1*
b10 6
19
1>
1C
b10 G
#218060000000
0!
0*
09
0>
0C
#218070000000
1!
1*
b11 6
19
1>
1C
b11 G
#218080000000
0!
0*
09
0>
0C
#218090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#218100000000
0!
0*
09
0>
0C
#218110000000
1!
1*
b101 6
19
1>
1C
b101 G
#218120000000
0!
0*
09
0>
0C
#218130000000
1!
1*
b110 6
19
1>
1C
b110 G
#218140000000
0!
0*
09
0>
0C
#218150000000
1!
1*
b111 6
19
1>
1C
b111 G
#218160000000
0!
0*
09
0>
0C
#218170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#218180000000
0!
0*
09
0>
0C
#218190000000
1!
1*
b1 6
19
1>
1C
b1 G
#218200000000
0!
0*
09
0>
0C
#218210000000
1!
1*
b10 6
19
1>
1C
b10 G
#218220000000
0!
0*
09
0>
0C
#218230000000
1!
1*
b11 6
19
1>
1C
b11 G
#218240000000
0!
0*
09
0>
0C
#218250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#218260000000
0!
0*
09
0>
0C
#218270000000
1!
1*
b101 6
19
1>
1C
b101 G
#218280000000
0!
0*
09
0>
0C
#218290000000
1!
1*
b110 6
19
1>
1C
b110 G
#218300000000
0!
0*
09
0>
0C
#218310000000
1!
1*
b111 6
19
1>
1C
b111 G
#218320000000
0!
1"
0*
1+
09
1:
0>
0C
#218330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#218340000000
0!
0*
09
0>
0C
#218350000000
1!
1*
b1 6
19
1>
1C
b1 G
#218360000000
0!
0*
09
0>
0C
#218370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#218380000000
0!
0*
09
0>
0C
#218390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#218400000000
0!
0*
09
0>
0C
#218410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#218420000000
0!
0*
09
0>
0C
#218430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#218440000000
0!
0#
0*
0,
09
0>
0?
0C
#218450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#218460000000
0!
0*
09
0>
0C
#218470000000
1!
1*
19
1>
1C
#218480000000
0!
0*
09
0>
0C
#218490000000
1!
1*
19
1>
1C
#218500000000
0!
0*
09
0>
0C
#218510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#218520000000
0!
0*
09
0>
0C
#218530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#218540000000
0!
0*
09
0>
0C
#218550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#218560000000
0!
0*
09
0>
0C
#218570000000
1!
1*
b10 6
19
1>
1C
b10 G
#218580000000
0!
0*
09
0>
0C
#218590000000
1!
1*
b11 6
19
1>
1C
b11 G
#218600000000
0!
0*
09
0>
0C
#218610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#218620000000
0!
0*
09
0>
0C
#218630000000
1!
1*
b101 6
19
1>
1C
b101 G
#218640000000
0!
0*
09
0>
0C
#218650000000
1!
1*
b110 6
19
1>
1C
b110 G
#218660000000
0!
0*
09
0>
0C
#218670000000
1!
1*
b111 6
19
1>
1C
b111 G
#218680000000
0!
0*
09
0>
0C
#218690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#218700000000
0!
0*
09
0>
0C
#218710000000
1!
1*
b1 6
19
1>
1C
b1 G
#218720000000
0!
0*
09
0>
0C
#218730000000
1!
1*
b10 6
19
1>
1C
b10 G
#218740000000
0!
0*
09
0>
0C
#218750000000
1!
1*
b11 6
19
1>
1C
b11 G
#218760000000
0!
0*
09
0>
0C
#218770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#218780000000
0!
0*
09
0>
0C
#218790000000
1!
1*
b101 6
19
1>
1C
b101 G
#218800000000
0!
0*
09
0>
0C
#218810000000
1!
1*
b110 6
19
1>
1C
b110 G
#218820000000
0!
0*
09
0>
0C
#218830000000
1!
1*
b111 6
19
1>
1C
b111 G
#218840000000
0!
0*
09
0>
0C
#218850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#218860000000
0!
0*
09
0>
0C
#218870000000
1!
1*
b1 6
19
1>
1C
b1 G
#218880000000
0!
0*
09
0>
0C
#218890000000
1!
1*
b10 6
19
1>
1C
b10 G
#218900000000
0!
0*
09
0>
0C
#218910000000
1!
1*
b11 6
19
1>
1C
b11 G
#218920000000
0!
0*
09
0>
0C
#218930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#218940000000
0!
0*
09
0>
0C
#218950000000
1!
1*
b101 6
19
1>
1C
b101 G
#218960000000
0!
0*
09
0>
0C
#218970000000
1!
1*
b110 6
19
1>
1C
b110 G
#218980000000
0!
0*
09
0>
0C
#218990000000
1!
1*
b111 6
19
1>
1C
b111 G
#219000000000
0!
1"
0*
1+
09
1:
0>
0C
#219010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#219020000000
0!
0*
09
0>
0C
#219030000000
1!
1*
b1 6
19
1>
1C
b1 G
#219040000000
0!
0*
09
0>
0C
#219050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#219060000000
0!
0*
09
0>
0C
#219070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#219080000000
0!
0*
09
0>
0C
#219090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#219100000000
0!
0*
09
0>
0C
#219110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#219120000000
0!
0#
0*
0,
09
0>
0?
0C
#219130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#219140000000
0!
0*
09
0>
0C
#219150000000
1!
1*
19
1>
1C
#219160000000
0!
0*
09
0>
0C
#219170000000
1!
1*
19
1>
1C
#219180000000
0!
0*
09
0>
0C
#219190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#219200000000
0!
0*
09
0>
0C
#219210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#219220000000
0!
0*
09
0>
0C
#219230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#219240000000
0!
0*
09
0>
0C
#219250000000
1!
1*
b10 6
19
1>
1C
b10 G
#219260000000
0!
0*
09
0>
0C
#219270000000
1!
1*
b11 6
19
1>
1C
b11 G
#219280000000
0!
0*
09
0>
0C
#219290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#219300000000
0!
0*
09
0>
0C
#219310000000
1!
1*
b101 6
19
1>
1C
b101 G
#219320000000
0!
0*
09
0>
0C
#219330000000
1!
1*
b110 6
19
1>
1C
b110 G
#219340000000
0!
0*
09
0>
0C
#219350000000
1!
1*
b111 6
19
1>
1C
b111 G
#219360000000
0!
0*
09
0>
0C
#219370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#219380000000
0!
0*
09
0>
0C
#219390000000
1!
1*
b1 6
19
1>
1C
b1 G
#219400000000
0!
0*
09
0>
0C
#219410000000
1!
1*
b10 6
19
1>
1C
b10 G
#219420000000
0!
0*
09
0>
0C
#219430000000
1!
1*
b11 6
19
1>
1C
b11 G
#219440000000
0!
0*
09
0>
0C
#219450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#219460000000
0!
0*
09
0>
0C
#219470000000
1!
1*
b101 6
19
1>
1C
b101 G
#219480000000
0!
0*
09
0>
0C
#219490000000
1!
1*
b110 6
19
1>
1C
b110 G
#219500000000
0!
0*
09
0>
0C
#219510000000
1!
1*
b111 6
19
1>
1C
b111 G
#219520000000
0!
0*
09
0>
0C
#219530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#219540000000
0!
0*
09
0>
0C
#219550000000
1!
1*
b1 6
19
1>
1C
b1 G
#219560000000
0!
0*
09
0>
0C
#219570000000
1!
1*
b10 6
19
1>
1C
b10 G
#219580000000
0!
0*
09
0>
0C
#219590000000
1!
1*
b11 6
19
1>
1C
b11 G
#219600000000
0!
0*
09
0>
0C
#219610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#219620000000
0!
0*
09
0>
0C
#219630000000
1!
1*
b101 6
19
1>
1C
b101 G
#219640000000
0!
0*
09
0>
0C
#219650000000
1!
1*
b110 6
19
1>
1C
b110 G
#219660000000
0!
0*
09
0>
0C
#219670000000
1!
1*
b111 6
19
1>
1C
b111 G
#219680000000
0!
1"
0*
1+
09
1:
0>
0C
#219690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#219700000000
0!
0*
09
0>
0C
#219710000000
1!
1*
b1 6
19
1>
1C
b1 G
#219720000000
0!
0*
09
0>
0C
#219730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#219740000000
0!
0*
09
0>
0C
#219750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#219760000000
0!
0*
09
0>
0C
#219770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#219780000000
0!
0*
09
0>
0C
#219790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#219800000000
0!
0#
0*
0,
09
0>
0?
0C
#219810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#219820000000
0!
0*
09
0>
0C
#219830000000
1!
1*
19
1>
1C
#219840000000
0!
0*
09
0>
0C
#219850000000
1!
1*
19
1>
1C
#219860000000
0!
0*
09
0>
0C
#219870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#219880000000
0!
0*
09
0>
0C
#219890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#219900000000
0!
0*
09
0>
0C
#219910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#219920000000
0!
0*
09
0>
0C
#219930000000
1!
1*
b10 6
19
1>
1C
b10 G
#219940000000
0!
0*
09
0>
0C
#219950000000
1!
1*
b11 6
19
1>
1C
b11 G
#219960000000
0!
0*
09
0>
0C
#219970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#219980000000
0!
0*
09
0>
0C
#219990000000
1!
1*
b101 6
19
1>
1C
b101 G
#220000000000
0!
0*
09
0>
0C
#220010000000
1!
1*
b110 6
19
1>
1C
b110 G
#220020000000
0!
0*
09
0>
0C
#220030000000
1!
1*
b111 6
19
1>
1C
b111 G
#220040000000
0!
0*
09
0>
0C
#220050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#220060000000
0!
0*
09
0>
0C
#220070000000
1!
1*
b1 6
19
1>
1C
b1 G
#220080000000
0!
0*
09
0>
0C
#220090000000
1!
1*
b10 6
19
1>
1C
b10 G
#220100000000
0!
0*
09
0>
0C
#220110000000
1!
1*
b11 6
19
1>
1C
b11 G
#220120000000
0!
0*
09
0>
0C
#220130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#220140000000
0!
0*
09
0>
0C
#220150000000
1!
1*
b101 6
19
1>
1C
b101 G
#220160000000
0!
0*
09
0>
0C
#220170000000
1!
1*
b110 6
19
1>
1C
b110 G
#220180000000
0!
0*
09
0>
0C
#220190000000
1!
1*
b111 6
19
1>
1C
b111 G
#220200000000
0!
0*
09
0>
0C
#220210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#220220000000
0!
0*
09
0>
0C
#220230000000
1!
1*
b1 6
19
1>
1C
b1 G
#220240000000
0!
0*
09
0>
0C
#220250000000
1!
1*
b10 6
19
1>
1C
b10 G
#220260000000
0!
0*
09
0>
0C
#220270000000
1!
1*
b11 6
19
1>
1C
b11 G
#220280000000
0!
0*
09
0>
0C
#220290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#220300000000
0!
0*
09
0>
0C
#220310000000
1!
1*
b101 6
19
1>
1C
b101 G
#220320000000
0!
0*
09
0>
0C
#220330000000
1!
1*
b110 6
19
1>
1C
b110 G
#220340000000
0!
0*
09
0>
0C
#220350000000
1!
1*
b111 6
19
1>
1C
b111 G
#220360000000
0!
1"
0*
1+
09
1:
0>
0C
#220370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#220380000000
0!
0*
09
0>
0C
#220390000000
1!
1*
b1 6
19
1>
1C
b1 G
#220400000000
0!
0*
09
0>
0C
#220410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#220420000000
0!
0*
09
0>
0C
#220430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#220440000000
0!
0*
09
0>
0C
#220450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#220460000000
0!
0*
09
0>
0C
#220470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#220480000000
0!
0#
0*
0,
09
0>
0?
0C
#220490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#220500000000
0!
0*
09
0>
0C
#220510000000
1!
1*
19
1>
1C
#220520000000
0!
0*
09
0>
0C
#220530000000
1!
1*
19
1>
1C
#220540000000
0!
0*
09
0>
0C
#220550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#220560000000
0!
0*
09
0>
0C
#220570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#220580000000
0!
0*
09
0>
0C
#220590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#220600000000
0!
0*
09
0>
0C
#220610000000
1!
1*
b10 6
19
1>
1C
b10 G
#220620000000
0!
0*
09
0>
0C
#220630000000
1!
1*
b11 6
19
1>
1C
b11 G
#220640000000
0!
0*
09
0>
0C
#220650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#220660000000
0!
0*
09
0>
0C
#220670000000
1!
1*
b101 6
19
1>
1C
b101 G
#220680000000
0!
0*
09
0>
0C
#220690000000
1!
1*
b110 6
19
1>
1C
b110 G
#220700000000
0!
0*
09
0>
0C
#220710000000
1!
1*
b111 6
19
1>
1C
b111 G
#220720000000
0!
0*
09
0>
0C
#220730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#220740000000
0!
0*
09
0>
0C
#220750000000
1!
1*
b1 6
19
1>
1C
b1 G
#220760000000
0!
0*
09
0>
0C
#220770000000
1!
1*
b10 6
19
1>
1C
b10 G
#220780000000
0!
0*
09
0>
0C
#220790000000
1!
1*
b11 6
19
1>
1C
b11 G
#220800000000
0!
0*
09
0>
0C
#220810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#220820000000
0!
0*
09
0>
0C
#220830000000
1!
1*
b101 6
19
1>
1C
b101 G
#220840000000
0!
0*
09
0>
0C
#220850000000
1!
1*
b110 6
19
1>
1C
b110 G
#220860000000
0!
0*
09
0>
0C
#220870000000
1!
1*
b111 6
19
1>
1C
b111 G
#220880000000
0!
0*
09
0>
0C
#220890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#220900000000
0!
0*
09
0>
0C
#220910000000
1!
1*
b1 6
19
1>
1C
b1 G
#220920000000
0!
0*
09
0>
0C
#220930000000
1!
1*
b10 6
19
1>
1C
b10 G
#220940000000
0!
0*
09
0>
0C
#220950000000
1!
1*
b11 6
19
1>
1C
b11 G
#220960000000
0!
0*
09
0>
0C
#220970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#220980000000
0!
0*
09
0>
0C
#220990000000
1!
1*
b101 6
19
1>
1C
b101 G
#221000000000
0!
0*
09
0>
0C
#221010000000
1!
1*
b110 6
19
1>
1C
b110 G
#221020000000
0!
0*
09
0>
0C
#221030000000
1!
1*
b111 6
19
1>
1C
b111 G
#221040000000
0!
1"
0*
1+
09
1:
0>
0C
#221050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#221060000000
0!
0*
09
0>
0C
#221070000000
1!
1*
b1 6
19
1>
1C
b1 G
#221080000000
0!
0*
09
0>
0C
#221090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#221100000000
0!
0*
09
0>
0C
#221110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#221120000000
0!
0*
09
0>
0C
#221130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#221140000000
0!
0*
09
0>
0C
#221150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#221160000000
0!
0#
0*
0,
09
0>
0?
0C
#221170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#221180000000
0!
0*
09
0>
0C
#221190000000
1!
1*
19
1>
1C
#221200000000
0!
0*
09
0>
0C
#221210000000
1!
1*
19
1>
1C
#221220000000
0!
0*
09
0>
0C
#221230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#221240000000
0!
0*
09
0>
0C
#221250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#221260000000
0!
0*
09
0>
0C
#221270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#221280000000
0!
0*
09
0>
0C
#221290000000
1!
1*
b10 6
19
1>
1C
b10 G
#221300000000
0!
0*
09
0>
0C
#221310000000
1!
1*
b11 6
19
1>
1C
b11 G
#221320000000
0!
0*
09
0>
0C
#221330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#221340000000
0!
0*
09
0>
0C
#221350000000
1!
1*
b101 6
19
1>
1C
b101 G
#221360000000
0!
0*
09
0>
0C
#221370000000
1!
1*
b110 6
19
1>
1C
b110 G
#221380000000
0!
0*
09
0>
0C
#221390000000
1!
1*
b111 6
19
1>
1C
b111 G
#221400000000
0!
0*
09
0>
0C
#221410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#221420000000
0!
0*
09
0>
0C
#221430000000
1!
1*
b1 6
19
1>
1C
b1 G
#221440000000
0!
0*
09
0>
0C
#221450000000
1!
1*
b10 6
19
1>
1C
b10 G
#221460000000
0!
0*
09
0>
0C
#221470000000
1!
1*
b11 6
19
1>
1C
b11 G
#221480000000
0!
0*
09
0>
0C
#221490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#221500000000
0!
0*
09
0>
0C
#221510000000
1!
1*
b101 6
19
1>
1C
b101 G
#221520000000
0!
0*
09
0>
0C
#221530000000
1!
1*
b110 6
19
1>
1C
b110 G
#221540000000
0!
0*
09
0>
0C
#221550000000
1!
1*
b111 6
19
1>
1C
b111 G
#221560000000
0!
0*
09
0>
0C
#221570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#221580000000
0!
0*
09
0>
0C
#221590000000
1!
1*
b1 6
19
1>
1C
b1 G
#221600000000
0!
0*
09
0>
0C
#221610000000
1!
1*
b10 6
19
1>
1C
b10 G
#221620000000
0!
0*
09
0>
0C
#221630000000
1!
1*
b11 6
19
1>
1C
b11 G
#221640000000
0!
0*
09
0>
0C
#221650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#221660000000
0!
0*
09
0>
0C
#221670000000
1!
1*
b101 6
19
1>
1C
b101 G
#221680000000
0!
0*
09
0>
0C
#221690000000
1!
1*
b110 6
19
1>
1C
b110 G
#221700000000
0!
0*
09
0>
0C
#221710000000
1!
1*
b111 6
19
1>
1C
b111 G
#221720000000
0!
1"
0*
1+
09
1:
0>
0C
#221730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#221740000000
0!
0*
09
0>
0C
#221750000000
1!
1*
b1 6
19
1>
1C
b1 G
#221760000000
0!
0*
09
0>
0C
#221770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#221780000000
0!
0*
09
0>
0C
#221790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#221800000000
0!
0*
09
0>
0C
#221810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#221820000000
0!
0*
09
0>
0C
#221830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#221840000000
0!
0#
0*
0,
09
0>
0?
0C
#221850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#221860000000
0!
0*
09
0>
0C
#221870000000
1!
1*
19
1>
1C
#221880000000
0!
0*
09
0>
0C
#221890000000
1!
1*
19
1>
1C
#221900000000
0!
0*
09
0>
0C
#221910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#221920000000
0!
0*
09
0>
0C
#221930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#221940000000
0!
0*
09
0>
0C
#221950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#221960000000
0!
0*
09
0>
0C
#221970000000
1!
1*
b10 6
19
1>
1C
b10 G
#221980000000
0!
0*
09
0>
0C
#221990000000
1!
1*
b11 6
19
1>
1C
b11 G
#222000000000
0!
0*
09
0>
0C
#222010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#222020000000
0!
0*
09
0>
0C
#222030000000
1!
1*
b101 6
19
1>
1C
b101 G
#222040000000
0!
0*
09
0>
0C
#222050000000
1!
1*
b110 6
19
1>
1C
b110 G
#222060000000
0!
0*
09
0>
0C
#222070000000
1!
1*
b111 6
19
1>
1C
b111 G
#222080000000
0!
0*
09
0>
0C
#222090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#222100000000
0!
0*
09
0>
0C
#222110000000
1!
1*
b1 6
19
1>
1C
b1 G
#222120000000
0!
0*
09
0>
0C
#222130000000
1!
1*
b10 6
19
1>
1C
b10 G
#222140000000
0!
0*
09
0>
0C
#222150000000
1!
1*
b11 6
19
1>
1C
b11 G
#222160000000
0!
0*
09
0>
0C
#222170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#222180000000
0!
0*
09
0>
0C
#222190000000
1!
1*
b101 6
19
1>
1C
b101 G
#222200000000
0!
0*
09
0>
0C
#222210000000
1!
1*
b110 6
19
1>
1C
b110 G
#222220000000
0!
0*
09
0>
0C
#222230000000
1!
1*
b111 6
19
1>
1C
b111 G
#222240000000
0!
0*
09
0>
0C
#222250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#222260000000
0!
0*
09
0>
0C
#222270000000
1!
1*
b1 6
19
1>
1C
b1 G
#222280000000
0!
0*
09
0>
0C
#222290000000
1!
1*
b10 6
19
1>
1C
b10 G
#222300000000
0!
0*
09
0>
0C
#222310000000
1!
1*
b11 6
19
1>
1C
b11 G
#222320000000
0!
0*
09
0>
0C
#222330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#222340000000
0!
0*
09
0>
0C
#222350000000
1!
1*
b101 6
19
1>
1C
b101 G
#222360000000
0!
0*
09
0>
0C
#222370000000
1!
1*
b110 6
19
1>
1C
b110 G
#222380000000
0!
0*
09
0>
0C
#222390000000
1!
1*
b111 6
19
1>
1C
b111 G
#222400000000
0!
1"
0*
1+
09
1:
0>
0C
#222410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#222420000000
0!
0*
09
0>
0C
#222430000000
1!
1*
b1 6
19
1>
1C
b1 G
#222440000000
0!
0*
09
0>
0C
#222450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#222460000000
0!
0*
09
0>
0C
#222470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#222480000000
0!
0*
09
0>
0C
#222490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#222500000000
0!
0*
09
0>
0C
#222510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#222520000000
0!
0#
0*
0,
09
0>
0?
0C
#222530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#222540000000
0!
0*
09
0>
0C
#222550000000
1!
1*
19
1>
1C
#222560000000
0!
0*
09
0>
0C
#222570000000
1!
1*
19
1>
1C
#222580000000
0!
0*
09
0>
0C
#222590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#222600000000
0!
0*
09
0>
0C
#222610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#222620000000
0!
0*
09
0>
0C
#222630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#222640000000
0!
0*
09
0>
0C
#222650000000
1!
1*
b10 6
19
1>
1C
b10 G
#222660000000
0!
0*
09
0>
0C
#222670000000
1!
1*
b11 6
19
1>
1C
b11 G
#222680000000
0!
0*
09
0>
0C
#222690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#222700000000
0!
0*
09
0>
0C
#222710000000
1!
1*
b101 6
19
1>
1C
b101 G
#222720000000
0!
0*
09
0>
0C
#222730000000
1!
1*
b110 6
19
1>
1C
b110 G
#222740000000
0!
0*
09
0>
0C
#222750000000
1!
1*
b111 6
19
1>
1C
b111 G
#222760000000
0!
0*
09
0>
0C
#222770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#222780000000
0!
0*
09
0>
0C
#222790000000
1!
1*
b1 6
19
1>
1C
b1 G
#222800000000
0!
0*
09
0>
0C
#222810000000
1!
1*
b10 6
19
1>
1C
b10 G
#222820000000
0!
0*
09
0>
0C
#222830000000
1!
1*
b11 6
19
1>
1C
b11 G
#222840000000
0!
0*
09
0>
0C
#222850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#222860000000
0!
0*
09
0>
0C
#222870000000
1!
1*
b101 6
19
1>
1C
b101 G
#222880000000
0!
0*
09
0>
0C
#222890000000
1!
1*
b110 6
19
1>
1C
b110 G
#222900000000
0!
0*
09
0>
0C
#222910000000
1!
1*
b111 6
19
1>
1C
b111 G
#222920000000
0!
0*
09
0>
0C
#222930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#222940000000
0!
0*
09
0>
0C
#222950000000
1!
1*
b1 6
19
1>
1C
b1 G
#222960000000
0!
0*
09
0>
0C
#222970000000
1!
1*
b10 6
19
1>
1C
b10 G
#222980000000
0!
0*
09
0>
0C
#222990000000
1!
1*
b11 6
19
1>
1C
b11 G
#223000000000
0!
0*
09
0>
0C
#223010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#223020000000
0!
0*
09
0>
0C
#223030000000
1!
1*
b101 6
19
1>
1C
b101 G
#223040000000
0!
0*
09
0>
0C
#223050000000
1!
1*
b110 6
19
1>
1C
b110 G
#223060000000
0!
0*
09
0>
0C
#223070000000
1!
1*
b111 6
19
1>
1C
b111 G
#223080000000
0!
1"
0*
1+
09
1:
0>
0C
#223090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#223100000000
0!
0*
09
0>
0C
#223110000000
1!
1*
b1 6
19
1>
1C
b1 G
#223120000000
0!
0*
09
0>
0C
#223130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#223140000000
0!
0*
09
0>
0C
#223150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#223160000000
0!
0*
09
0>
0C
#223170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#223180000000
0!
0*
09
0>
0C
#223190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#223200000000
0!
0#
0*
0,
09
0>
0?
0C
#223210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#223220000000
0!
0*
09
0>
0C
#223230000000
1!
1*
19
1>
1C
#223240000000
0!
0*
09
0>
0C
#223250000000
1!
1*
19
1>
1C
#223260000000
0!
0*
09
0>
0C
#223270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#223280000000
0!
0*
09
0>
0C
#223290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#223300000000
0!
0*
09
0>
0C
#223310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#223320000000
0!
0*
09
0>
0C
#223330000000
1!
1*
b10 6
19
1>
1C
b10 G
#223340000000
0!
0*
09
0>
0C
#223350000000
1!
1*
b11 6
19
1>
1C
b11 G
#223360000000
0!
0*
09
0>
0C
#223370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#223380000000
0!
0*
09
0>
0C
#223390000000
1!
1*
b101 6
19
1>
1C
b101 G
#223400000000
0!
0*
09
0>
0C
#223410000000
1!
1*
b110 6
19
1>
1C
b110 G
#223420000000
0!
0*
09
0>
0C
#223430000000
1!
1*
b111 6
19
1>
1C
b111 G
#223440000000
0!
0*
09
0>
0C
#223450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#223460000000
0!
0*
09
0>
0C
#223470000000
1!
1*
b1 6
19
1>
1C
b1 G
#223480000000
0!
0*
09
0>
0C
#223490000000
1!
1*
b10 6
19
1>
1C
b10 G
#223500000000
0!
0*
09
0>
0C
#223510000000
1!
1*
b11 6
19
1>
1C
b11 G
#223520000000
0!
0*
09
0>
0C
#223530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#223540000000
0!
0*
09
0>
0C
#223550000000
1!
1*
b101 6
19
1>
1C
b101 G
#223560000000
0!
0*
09
0>
0C
#223570000000
1!
1*
b110 6
19
1>
1C
b110 G
#223580000000
0!
0*
09
0>
0C
#223590000000
1!
1*
b111 6
19
1>
1C
b111 G
#223600000000
0!
0*
09
0>
0C
#223610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#223620000000
0!
0*
09
0>
0C
#223630000000
1!
1*
b1 6
19
1>
1C
b1 G
#223640000000
0!
0*
09
0>
0C
#223650000000
1!
1*
b10 6
19
1>
1C
b10 G
#223660000000
0!
0*
09
0>
0C
#223670000000
1!
1*
b11 6
19
1>
1C
b11 G
#223680000000
0!
0*
09
0>
0C
#223690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#223700000000
0!
0*
09
0>
0C
#223710000000
1!
1*
b101 6
19
1>
1C
b101 G
#223720000000
0!
0*
09
0>
0C
#223730000000
1!
1*
b110 6
19
1>
1C
b110 G
#223740000000
0!
0*
09
0>
0C
#223750000000
1!
1*
b111 6
19
1>
1C
b111 G
#223760000000
0!
1"
0*
1+
09
1:
0>
0C
#223770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#223780000000
0!
0*
09
0>
0C
#223790000000
1!
1*
b1 6
19
1>
1C
b1 G
#223800000000
0!
0*
09
0>
0C
#223810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#223820000000
0!
0*
09
0>
0C
#223830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#223840000000
0!
0*
09
0>
0C
#223850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#223860000000
0!
0*
09
0>
0C
#223870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#223880000000
0!
0#
0*
0,
09
0>
0?
0C
#223890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#223900000000
0!
0*
09
0>
0C
#223910000000
1!
1*
19
1>
1C
#223920000000
0!
0*
09
0>
0C
#223930000000
1!
1*
19
1>
1C
#223940000000
0!
0*
09
0>
0C
#223950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#223960000000
0!
0*
09
0>
0C
#223970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#223980000000
0!
0*
09
0>
0C
#223990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#224000000000
0!
0*
09
0>
0C
#224010000000
1!
1*
b10 6
19
1>
1C
b10 G
#224020000000
0!
0*
09
0>
0C
#224030000000
1!
1*
b11 6
19
1>
1C
b11 G
#224040000000
0!
0*
09
0>
0C
#224050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#224060000000
0!
0*
09
0>
0C
#224070000000
1!
1*
b101 6
19
1>
1C
b101 G
#224080000000
0!
0*
09
0>
0C
#224090000000
1!
1*
b110 6
19
1>
1C
b110 G
#224100000000
0!
0*
09
0>
0C
#224110000000
1!
1*
b111 6
19
1>
1C
b111 G
#224120000000
0!
0*
09
0>
0C
#224130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#224140000000
0!
0*
09
0>
0C
#224150000000
1!
1*
b1 6
19
1>
1C
b1 G
#224160000000
0!
0*
09
0>
0C
#224170000000
1!
1*
b10 6
19
1>
1C
b10 G
#224180000000
0!
0*
09
0>
0C
#224190000000
1!
1*
b11 6
19
1>
1C
b11 G
#224200000000
0!
0*
09
0>
0C
#224210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#224220000000
0!
0*
09
0>
0C
#224230000000
1!
1*
b101 6
19
1>
1C
b101 G
#224240000000
0!
0*
09
0>
0C
#224250000000
1!
1*
b110 6
19
1>
1C
b110 G
#224260000000
0!
0*
09
0>
0C
#224270000000
1!
1*
b111 6
19
1>
1C
b111 G
#224280000000
0!
0*
09
0>
0C
#224290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#224300000000
0!
0*
09
0>
0C
#224310000000
1!
1*
b1 6
19
1>
1C
b1 G
#224320000000
0!
0*
09
0>
0C
#224330000000
1!
1*
b10 6
19
1>
1C
b10 G
#224340000000
0!
0*
09
0>
0C
#224350000000
1!
1*
b11 6
19
1>
1C
b11 G
#224360000000
0!
0*
09
0>
0C
#224370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#224380000000
0!
0*
09
0>
0C
#224390000000
1!
1*
b101 6
19
1>
1C
b101 G
#224400000000
0!
0*
09
0>
0C
#224410000000
1!
1*
b110 6
19
1>
1C
b110 G
#224420000000
0!
0*
09
0>
0C
#224430000000
1!
1*
b111 6
19
1>
1C
b111 G
#224440000000
0!
1"
0*
1+
09
1:
0>
0C
#224450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#224460000000
0!
0*
09
0>
0C
#224470000000
1!
1*
b1 6
19
1>
1C
b1 G
#224480000000
0!
0*
09
0>
0C
#224490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#224500000000
0!
0*
09
0>
0C
#224510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#224520000000
0!
0*
09
0>
0C
#224530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#224540000000
0!
0*
09
0>
0C
#224550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#224560000000
0!
0#
0*
0,
09
0>
0?
0C
#224570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#224580000000
0!
0*
09
0>
0C
#224590000000
1!
1*
19
1>
1C
#224600000000
0!
0*
09
0>
0C
#224610000000
1!
1*
19
1>
1C
#224620000000
0!
0*
09
0>
0C
#224630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#224640000000
0!
0*
09
0>
0C
#224650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#224660000000
0!
0*
09
0>
0C
#224670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#224680000000
0!
0*
09
0>
0C
#224690000000
1!
1*
b10 6
19
1>
1C
b10 G
#224700000000
0!
0*
09
0>
0C
#224710000000
1!
1*
b11 6
19
1>
1C
b11 G
#224720000000
0!
0*
09
0>
0C
#224730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#224740000000
0!
0*
09
0>
0C
#224750000000
1!
1*
b101 6
19
1>
1C
b101 G
#224760000000
0!
0*
09
0>
0C
#224770000000
1!
1*
b110 6
19
1>
1C
b110 G
#224780000000
0!
0*
09
0>
0C
#224790000000
1!
1*
b111 6
19
1>
1C
b111 G
#224800000000
0!
0*
09
0>
0C
#224810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#224820000000
0!
0*
09
0>
0C
#224830000000
1!
1*
b1 6
19
1>
1C
b1 G
#224840000000
0!
0*
09
0>
0C
#224850000000
1!
1*
b10 6
19
1>
1C
b10 G
#224860000000
0!
0*
09
0>
0C
#224870000000
1!
1*
b11 6
19
1>
1C
b11 G
#224880000000
0!
0*
09
0>
0C
#224890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#224900000000
0!
0*
09
0>
0C
#224910000000
1!
1*
b101 6
19
1>
1C
b101 G
#224920000000
0!
0*
09
0>
0C
#224930000000
1!
1*
b110 6
19
1>
1C
b110 G
#224940000000
0!
0*
09
0>
0C
#224950000000
1!
1*
b111 6
19
1>
1C
b111 G
#224960000000
0!
0*
09
0>
0C
#224970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#224980000000
0!
0*
09
0>
0C
#224990000000
1!
1*
b1 6
19
1>
1C
b1 G
#225000000000
0!
0*
09
0>
0C
#225010000000
1!
1*
b10 6
19
1>
1C
b10 G
#225020000000
0!
0*
09
0>
0C
#225030000000
1!
1*
b11 6
19
1>
1C
b11 G
#225040000000
0!
0*
09
0>
0C
#225050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#225060000000
0!
0*
09
0>
0C
#225070000000
1!
1*
b101 6
19
1>
1C
b101 G
#225080000000
0!
0*
09
0>
0C
#225090000000
1!
1*
b110 6
19
1>
1C
b110 G
#225100000000
0!
0*
09
0>
0C
#225110000000
1!
1*
b111 6
19
1>
1C
b111 G
#225120000000
0!
1"
0*
1+
09
1:
0>
0C
#225130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#225140000000
0!
0*
09
0>
0C
#225150000000
1!
1*
b1 6
19
1>
1C
b1 G
#225160000000
0!
0*
09
0>
0C
#225170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#225180000000
0!
0*
09
0>
0C
#225190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#225200000000
0!
0*
09
0>
0C
#225210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#225220000000
0!
0*
09
0>
0C
#225230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#225240000000
0!
0#
0*
0,
09
0>
0?
0C
#225250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#225260000000
0!
0*
09
0>
0C
#225270000000
1!
1*
19
1>
1C
#225280000000
0!
0*
09
0>
0C
#225290000000
1!
1*
19
1>
1C
#225300000000
0!
0*
09
0>
0C
#225310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#225320000000
0!
0*
09
0>
0C
#225330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#225340000000
0!
0*
09
0>
0C
#225350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#225360000000
0!
0*
09
0>
0C
#225370000000
1!
1*
b10 6
19
1>
1C
b10 G
#225380000000
0!
0*
09
0>
0C
#225390000000
1!
1*
b11 6
19
1>
1C
b11 G
#225400000000
0!
0*
09
0>
0C
#225410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#225420000000
0!
0*
09
0>
0C
#225430000000
1!
1*
b101 6
19
1>
1C
b101 G
#225440000000
0!
0*
09
0>
0C
#225450000000
1!
1*
b110 6
19
1>
1C
b110 G
#225460000000
0!
0*
09
0>
0C
#225470000000
1!
1*
b111 6
19
1>
1C
b111 G
#225480000000
0!
0*
09
0>
0C
#225490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#225500000000
0!
0*
09
0>
0C
#225510000000
1!
1*
b1 6
19
1>
1C
b1 G
#225520000000
0!
0*
09
0>
0C
#225530000000
1!
1*
b10 6
19
1>
1C
b10 G
#225540000000
0!
0*
09
0>
0C
#225550000000
1!
1*
b11 6
19
1>
1C
b11 G
#225560000000
0!
0*
09
0>
0C
#225570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#225580000000
0!
0*
09
0>
0C
#225590000000
1!
1*
b101 6
19
1>
1C
b101 G
#225600000000
0!
0*
09
0>
0C
#225610000000
1!
1*
b110 6
19
1>
1C
b110 G
#225620000000
0!
0*
09
0>
0C
#225630000000
1!
1*
b111 6
19
1>
1C
b111 G
#225640000000
0!
0*
09
0>
0C
#225650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#225660000000
0!
0*
09
0>
0C
#225670000000
1!
1*
b1 6
19
1>
1C
b1 G
#225680000000
0!
0*
09
0>
0C
#225690000000
1!
1*
b10 6
19
1>
1C
b10 G
#225700000000
0!
0*
09
0>
0C
#225710000000
1!
1*
b11 6
19
1>
1C
b11 G
#225720000000
0!
0*
09
0>
0C
#225730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#225740000000
0!
0*
09
0>
0C
#225750000000
1!
1*
b101 6
19
1>
1C
b101 G
#225760000000
0!
0*
09
0>
0C
#225770000000
1!
1*
b110 6
19
1>
1C
b110 G
#225780000000
0!
0*
09
0>
0C
#225790000000
1!
1*
b111 6
19
1>
1C
b111 G
#225800000000
0!
1"
0*
1+
09
1:
0>
0C
#225810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#225820000000
0!
0*
09
0>
0C
#225830000000
1!
1*
b1 6
19
1>
1C
b1 G
#225840000000
0!
0*
09
0>
0C
#225850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#225860000000
0!
0*
09
0>
0C
#225870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#225880000000
0!
0*
09
0>
0C
#225890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#225900000000
0!
0*
09
0>
0C
#225910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#225920000000
0!
0#
0*
0,
09
0>
0?
0C
#225930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#225940000000
0!
0*
09
0>
0C
#225950000000
1!
1*
19
1>
1C
#225960000000
0!
0*
09
0>
0C
#225970000000
1!
1*
19
1>
1C
#225980000000
0!
0*
09
0>
0C
#225990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#226000000000
0!
0*
09
0>
0C
#226010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#226020000000
0!
0*
09
0>
0C
#226030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#226040000000
0!
0*
09
0>
0C
#226050000000
1!
1*
b10 6
19
1>
1C
b10 G
#226060000000
0!
0*
09
0>
0C
#226070000000
1!
1*
b11 6
19
1>
1C
b11 G
#226080000000
0!
0*
09
0>
0C
#226090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#226100000000
0!
0*
09
0>
0C
#226110000000
1!
1*
b101 6
19
1>
1C
b101 G
#226120000000
0!
0*
09
0>
0C
#226130000000
1!
1*
b110 6
19
1>
1C
b110 G
#226140000000
0!
0*
09
0>
0C
#226150000000
1!
1*
b111 6
19
1>
1C
b111 G
#226160000000
0!
0*
09
0>
0C
#226170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#226180000000
0!
0*
09
0>
0C
#226190000000
1!
1*
b1 6
19
1>
1C
b1 G
#226200000000
0!
0*
09
0>
0C
#226210000000
1!
1*
b10 6
19
1>
1C
b10 G
#226220000000
0!
0*
09
0>
0C
#226230000000
1!
1*
b11 6
19
1>
1C
b11 G
#226240000000
0!
0*
09
0>
0C
#226250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#226260000000
0!
0*
09
0>
0C
#226270000000
1!
1*
b101 6
19
1>
1C
b101 G
#226280000000
0!
0*
09
0>
0C
#226290000000
1!
1*
b110 6
19
1>
1C
b110 G
#226300000000
0!
0*
09
0>
0C
#226310000000
1!
1*
b111 6
19
1>
1C
b111 G
#226320000000
0!
0*
09
0>
0C
#226330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#226340000000
0!
0*
09
0>
0C
#226350000000
1!
1*
b1 6
19
1>
1C
b1 G
#226360000000
0!
0*
09
0>
0C
#226370000000
1!
1*
b10 6
19
1>
1C
b10 G
#226380000000
0!
0*
09
0>
0C
#226390000000
1!
1*
b11 6
19
1>
1C
b11 G
#226400000000
0!
0*
09
0>
0C
#226410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#226420000000
0!
0*
09
0>
0C
#226430000000
1!
1*
b101 6
19
1>
1C
b101 G
#226440000000
0!
0*
09
0>
0C
#226450000000
1!
1*
b110 6
19
1>
1C
b110 G
#226460000000
0!
0*
09
0>
0C
#226470000000
1!
1*
b111 6
19
1>
1C
b111 G
#226480000000
0!
1"
0*
1+
09
1:
0>
0C
#226490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#226500000000
0!
0*
09
0>
0C
#226510000000
1!
1*
b1 6
19
1>
1C
b1 G
#226520000000
0!
0*
09
0>
0C
#226530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#226540000000
0!
0*
09
0>
0C
#226550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#226560000000
0!
0*
09
0>
0C
#226570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#226580000000
0!
0*
09
0>
0C
#226590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#226600000000
0!
0#
0*
0,
09
0>
0?
0C
#226610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#226620000000
0!
0*
09
0>
0C
#226630000000
1!
1*
19
1>
1C
#226640000000
0!
0*
09
0>
0C
#226650000000
1!
1*
19
1>
1C
#226660000000
0!
0*
09
0>
0C
#226670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#226680000000
0!
0*
09
0>
0C
#226690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#226700000000
0!
0*
09
0>
0C
#226710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#226720000000
0!
0*
09
0>
0C
#226730000000
1!
1*
b10 6
19
1>
1C
b10 G
#226740000000
0!
0*
09
0>
0C
#226750000000
1!
1*
b11 6
19
1>
1C
b11 G
#226760000000
0!
0*
09
0>
0C
#226770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#226780000000
0!
0*
09
0>
0C
#226790000000
1!
1*
b101 6
19
1>
1C
b101 G
#226800000000
0!
0*
09
0>
0C
#226810000000
1!
1*
b110 6
19
1>
1C
b110 G
#226820000000
0!
0*
09
0>
0C
#226830000000
1!
1*
b111 6
19
1>
1C
b111 G
#226840000000
0!
0*
09
0>
0C
#226850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#226860000000
0!
0*
09
0>
0C
#226870000000
1!
1*
b1 6
19
1>
1C
b1 G
#226880000000
0!
0*
09
0>
0C
#226890000000
1!
1*
b10 6
19
1>
1C
b10 G
#226900000000
0!
0*
09
0>
0C
#226910000000
1!
1*
b11 6
19
1>
1C
b11 G
#226920000000
0!
0*
09
0>
0C
#226930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#226940000000
0!
0*
09
0>
0C
#226950000000
1!
1*
b101 6
19
1>
1C
b101 G
#226960000000
0!
0*
09
0>
0C
#226970000000
1!
1*
b110 6
19
1>
1C
b110 G
#226980000000
0!
0*
09
0>
0C
#226990000000
1!
1*
b111 6
19
1>
1C
b111 G
#227000000000
0!
0*
09
0>
0C
#227010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#227020000000
0!
0*
09
0>
0C
#227030000000
1!
1*
b1 6
19
1>
1C
b1 G
#227040000000
0!
0*
09
0>
0C
#227050000000
1!
1*
b10 6
19
1>
1C
b10 G
#227060000000
0!
0*
09
0>
0C
#227070000000
1!
1*
b11 6
19
1>
1C
b11 G
#227080000000
0!
0*
09
0>
0C
#227090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#227100000000
0!
0*
09
0>
0C
#227110000000
1!
1*
b101 6
19
1>
1C
b101 G
#227120000000
0!
0*
09
0>
0C
#227130000000
1!
1*
b110 6
19
1>
1C
b110 G
#227140000000
0!
0*
09
0>
0C
#227150000000
1!
1*
b111 6
19
1>
1C
b111 G
#227160000000
0!
1"
0*
1+
09
1:
0>
0C
#227170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#227180000000
0!
0*
09
0>
0C
#227190000000
1!
1*
b1 6
19
1>
1C
b1 G
#227200000000
0!
0*
09
0>
0C
#227210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#227220000000
0!
0*
09
0>
0C
#227230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#227240000000
0!
0*
09
0>
0C
#227250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#227260000000
0!
0*
09
0>
0C
#227270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#227280000000
0!
0#
0*
0,
09
0>
0?
0C
#227290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#227300000000
0!
0*
09
0>
0C
#227310000000
1!
1*
19
1>
1C
#227320000000
0!
0*
09
0>
0C
#227330000000
1!
1*
19
1>
1C
#227340000000
0!
0*
09
0>
0C
#227350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#227360000000
0!
0*
09
0>
0C
#227370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#227380000000
0!
0*
09
0>
0C
#227390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#227400000000
0!
0*
09
0>
0C
#227410000000
1!
1*
b10 6
19
1>
1C
b10 G
#227420000000
0!
0*
09
0>
0C
#227430000000
1!
1*
b11 6
19
1>
1C
b11 G
#227440000000
0!
0*
09
0>
0C
#227450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#227460000000
0!
0*
09
0>
0C
#227470000000
1!
1*
b101 6
19
1>
1C
b101 G
#227480000000
0!
0*
09
0>
0C
#227490000000
1!
1*
b110 6
19
1>
1C
b110 G
#227500000000
0!
0*
09
0>
0C
#227510000000
1!
1*
b111 6
19
1>
1C
b111 G
#227520000000
0!
0*
09
0>
0C
#227530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#227540000000
0!
0*
09
0>
0C
#227550000000
1!
1*
b1 6
19
1>
1C
b1 G
#227560000000
0!
0*
09
0>
0C
#227570000000
1!
1*
b10 6
19
1>
1C
b10 G
#227580000000
0!
0*
09
0>
0C
#227590000000
1!
1*
b11 6
19
1>
1C
b11 G
#227600000000
0!
0*
09
0>
0C
#227610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#227620000000
0!
0*
09
0>
0C
#227630000000
1!
1*
b101 6
19
1>
1C
b101 G
#227640000000
0!
0*
09
0>
0C
#227650000000
1!
1*
b110 6
19
1>
1C
b110 G
#227660000000
0!
0*
09
0>
0C
#227670000000
1!
1*
b111 6
19
1>
1C
b111 G
#227680000000
0!
0*
09
0>
0C
#227690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#227700000000
0!
0*
09
0>
0C
#227710000000
1!
1*
b1 6
19
1>
1C
b1 G
#227720000000
0!
0*
09
0>
0C
#227730000000
1!
1*
b10 6
19
1>
1C
b10 G
#227740000000
0!
0*
09
0>
0C
#227750000000
1!
1*
b11 6
19
1>
1C
b11 G
#227760000000
0!
0*
09
0>
0C
#227770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#227780000000
0!
0*
09
0>
0C
#227790000000
1!
1*
b101 6
19
1>
1C
b101 G
#227800000000
0!
0*
09
0>
0C
#227810000000
1!
1*
b110 6
19
1>
1C
b110 G
#227820000000
0!
0*
09
0>
0C
#227830000000
1!
1*
b111 6
19
1>
1C
b111 G
#227840000000
0!
1"
0*
1+
09
1:
0>
0C
#227850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#227860000000
0!
0*
09
0>
0C
#227870000000
1!
1*
b1 6
19
1>
1C
b1 G
#227880000000
0!
0*
09
0>
0C
#227890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#227900000000
0!
0*
09
0>
0C
#227910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#227920000000
0!
0*
09
0>
0C
#227930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#227940000000
0!
0*
09
0>
0C
#227950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#227960000000
0!
0#
0*
0,
09
0>
0?
0C
#227970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#227980000000
0!
0*
09
0>
0C
#227990000000
1!
1*
19
1>
1C
#228000000000
0!
0*
09
0>
0C
#228010000000
1!
1*
19
1>
1C
#228020000000
0!
0*
09
0>
0C
#228030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#228040000000
0!
0*
09
0>
0C
#228050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#228060000000
0!
0*
09
0>
0C
#228070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#228080000000
0!
0*
09
0>
0C
#228090000000
1!
1*
b10 6
19
1>
1C
b10 G
#228100000000
0!
0*
09
0>
0C
#228110000000
1!
1*
b11 6
19
1>
1C
b11 G
#228120000000
0!
0*
09
0>
0C
#228130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#228140000000
0!
0*
09
0>
0C
#228150000000
1!
1*
b101 6
19
1>
1C
b101 G
#228160000000
0!
0*
09
0>
0C
#228170000000
1!
1*
b110 6
19
1>
1C
b110 G
#228180000000
0!
0*
09
0>
0C
#228190000000
1!
1*
b111 6
19
1>
1C
b111 G
#228200000000
0!
0*
09
0>
0C
#228210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#228220000000
0!
0*
09
0>
0C
#228230000000
1!
1*
b1 6
19
1>
1C
b1 G
#228240000000
0!
0*
09
0>
0C
#228250000000
1!
1*
b10 6
19
1>
1C
b10 G
#228260000000
0!
0*
09
0>
0C
#228270000000
1!
1*
b11 6
19
1>
1C
b11 G
#228280000000
0!
0*
09
0>
0C
#228290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#228300000000
0!
0*
09
0>
0C
#228310000000
1!
1*
b101 6
19
1>
1C
b101 G
#228320000000
0!
0*
09
0>
0C
#228330000000
1!
1*
b110 6
19
1>
1C
b110 G
#228340000000
0!
0*
09
0>
0C
#228350000000
1!
1*
b111 6
19
1>
1C
b111 G
#228360000000
0!
0*
09
0>
0C
#228370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#228380000000
0!
0*
09
0>
0C
#228390000000
1!
1*
b1 6
19
1>
1C
b1 G
#228400000000
0!
0*
09
0>
0C
#228410000000
1!
1*
b10 6
19
1>
1C
b10 G
#228420000000
0!
0*
09
0>
0C
#228430000000
1!
1*
b11 6
19
1>
1C
b11 G
#228440000000
0!
0*
09
0>
0C
#228450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#228460000000
0!
0*
09
0>
0C
#228470000000
1!
1*
b101 6
19
1>
1C
b101 G
#228480000000
0!
0*
09
0>
0C
#228490000000
1!
1*
b110 6
19
1>
1C
b110 G
#228500000000
0!
0*
09
0>
0C
#228510000000
1!
1*
b111 6
19
1>
1C
b111 G
#228520000000
0!
1"
0*
1+
09
1:
0>
0C
#228530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#228540000000
0!
0*
09
0>
0C
#228550000000
1!
1*
b1 6
19
1>
1C
b1 G
#228560000000
0!
0*
09
0>
0C
#228570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#228580000000
0!
0*
09
0>
0C
#228590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#228600000000
0!
0*
09
0>
0C
#228610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#228620000000
0!
0*
09
0>
0C
#228630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#228640000000
0!
0#
0*
0,
09
0>
0?
0C
#228650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#228660000000
0!
0*
09
0>
0C
#228670000000
1!
1*
19
1>
1C
#228680000000
0!
0*
09
0>
0C
#228690000000
1!
1*
19
1>
1C
#228700000000
0!
0*
09
0>
0C
#228710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#228720000000
0!
0*
09
0>
0C
#228730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#228740000000
0!
0*
09
0>
0C
#228750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#228760000000
0!
0*
09
0>
0C
#228770000000
1!
1*
b10 6
19
1>
1C
b10 G
#228780000000
0!
0*
09
0>
0C
#228790000000
1!
1*
b11 6
19
1>
1C
b11 G
#228800000000
0!
0*
09
0>
0C
#228810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#228820000000
0!
0*
09
0>
0C
#228830000000
1!
1*
b101 6
19
1>
1C
b101 G
#228840000000
0!
0*
09
0>
0C
#228850000000
1!
1*
b110 6
19
1>
1C
b110 G
#228860000000
0!
0*
09
0>
0C
#228870000000
1!
1*
b111 6
19
1>
1C
b111 G
#228880000000
0!
0*
09
0>
0C
#228890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#228900000000
0!
0*
09
0>
0C
#228910000000
1!
1*
b1 6
19
1>
1C
b1 G
#228920000000
0!
0*
09
0>
0C
#228930000000
1!
1*
b10 6
19
1>
1C
b10 G
#228940000000
0!
0*
09
0>
0C
#228950000000
1!
1*
b11 6
19
1>
1C
b11 G
#228960000000
0!
0*
09
0>
0C
#228970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#228980000000
0!
0*
09
0>
0C
#228990000000
1!
1*
b101 6
19
1>
1C
b101 G
#229000000000
0!
0*
09
0>
0C
#229010000000
1!
1*
b110 6
19
1>
1C
b110 G
#229020000000
0!
0*
09
0>
0C
#229030000000
1!
1*
b111 6
19
1>
1C
b111 G
#229040000000
0!
0*
09
0>
0C
#229050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#229060000000
0!
0*
09
0>
0C
#229070000000
1!
1*
b1 6
19
1>
1C
b1 G
#229080000000
0!
0*
09
0>
0C
#229090000000
1!
1*
b10 6
19
1>
1C
b10 G
#229100000000
0!
0*
09
0>
0C
#229110000000
1!
1*
b11 6
19
1>
1C
b11 G
#229120000000
0!
0*
09
0>
0C
#229130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#229140000000
0!
0*
09
0>
0C
#229150000000
1!
1*
b101 6
19
1>
1C
b101 G
#229160000000
0!
0*
09
0>
0C
#229170000000
1!
1*
b110 6
19
1>
1C
b110 G
#229180000000
0!
0*
09
0>
0C
#229190000000
1!
1*
b111 6
19
1>
1C
b111 G
#229200000000
0!
1"
0*
1+
09
1:
0>
0C
#229210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#229220000000
0!
0*
09
0>
0C
#229230000000
1!
1*
b1 6
19
1>
1C
b1 G
#229240000000
0!
0*
09
0>
0C
#229250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#229260000000
0!
0*
09
0>
0C
#229270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#229280000000
0!
0*
09
0>
0C
#229290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#229300000000
0!
0*
09
0>
0C
#229310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#229320000000
0!
0#
0*
0,
09
0>
0?
0C
#229330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#229340000000
0!
0*
09
0>
0C
#229350000000
1!
1*
19
1>
1C
#229360000000
0!
0*
09
0>
0C
#229370000000
1!
1*
19
1>
1C
#229380000000
0!
0*
09
0>
0C
#229390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#229400000000
0!
0*
09
0>
0C
#229410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#229420000000
0!
0*
09
0>
0C
#229430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#229440000000
0!
0*
09
0>
0C
#229450000000
1!
1*
b10 6
19
1>
1C
b10 G
#229460000000
0!
0*
09
0>
0C
#229470000000
1!
1*
b11 6
19
1>
1C
b11 G
#229480000000
0!
0*
09
0>
0C
#229490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#229500000000
0!
0*
09
0>
0C
#229510000000
1!
1*
b101 6
19
1>
1C
b101 G
#229520000000
0!
0*
09
0>
0C
#229530000000
1!
1*
b110 6
19
1>
1C
b110 G
#229540000000
0!
0*
09
0>
0C
#229550000000
1!
1*
b111 6
19
1>
1C
b111 G
#229560000000
0!
0*
09
0>
0C
#229570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#229580000000
0!
0*
09
0>
0C
#229590000000
1!
1*
b1 6
19
1>
1C
b1 G
#229600000000
0!
0*
09
0>
0C
#229610000000
1!
1*
b10 6
19
1>
1C
b10 G
#229620000000
0!
0*
09
0>
0C
#229630000000
1!
1*
b11 6
19
1>
1C
b11 G
#229640000000
0!
0*
09
0>
0C
#229650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#229660000000
0!
0*
09
0>
0C
#229670000000
1!
1*
b101 6
19
1>
1C
b101 G
#229680000000
0!
0*
09
0>
0C
#229690000000
1!
1*
b110 6
19
1>
1C
b110 G
#229700000000
0!
0*
09
0>
0C
#229710000000
1!
1*
b111 6
19
1>
1C
b111 G
#229720000000
0!
0*
09
0>
0C
#229730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#229740000000
0!
0*
09
0>
0C
#229750000000
1!
1*
b1 6
19
1>
1C
b1 G
#229760000000
0!
0*
09
0>
0C
#229770000000
1!
1*
b10 6
19
1>
1C
b10 G
#229780000000
0!
0*
09
0>
0C
#229790000000
1!
1*
b11 6
19
1>
1C
b11 G
#229800000000
0!
0*
09
0>
0C
#229810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#229820000000
0!
0*
09
0>
0C
#229830000000
1!
1*
b101 6
19
1>
1C
b101 G
#229840000000
0!
0*
09
0>
0C
#229850000000
1!
1*
b110 6
19
1>
1C
b110 G
#229860000000
0!
0*
09
0>
0C
#229870000000
1!
1*
b111 6
19
1>
1C
b111 G
#229880000000
0!
1"
0*
1+
09
1:
0>
0C
#229890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#229900000000
0!
0*
09
0>
0C
#229910000000
1!
1*
b1 6
19
1>
1C
b1 G
#229920000000
0!
0*
09
0>
0C
#229930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#229940000000
0!
0*
09
0>
0C
#229950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#229960000000
0!
0*
09
0>
0C
#229970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#229980000000
0!
0*
09
0>
0C
#229990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#230000000000
0!
0#
0*
0,
09
0>
0?
0C
#230010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#230020000000
0!
0*
09
0>
0C
#230030000000
1!
1*
19
1>
1C
#230040000000
0!
0*
09
0>
0C
#230050000000
1!
1*
19
1>
1C
#230060000000
0!
0*
09
0>
0C
#230070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#230080000000
0!
0*
09
0>
0C
#230090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#230100000000
0!
0*
09
0>
0C
#230110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#230120000000
0!
0*
09
0>
0C
#230130000000
1!
1*
b10 6
19
1>
1C
b10 G
#230140000000
0!
0*
09
0>
0C
#230150000000
1!
1*
b11 6
19
1>
1C
b11 G
#230160000000
0!
0*
09
0>
0C
#230170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#230180000000
0!
0*
09
0>
0C
#230190000000
1!
1*
b101 6
19
1>
1C
b101 G
#230200000000
0!
0*
09
0>
0C
#230210000000
1!
1*
b110 6
19
1>
1C
b110 G
#230220000000
0!
0*
09
0>
0C
#230230000000
1!
1*
b111 6
19
1>
1C
b111 G
#230240000000
0!
0*
09
0>
0C
#230250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#230260000000
0!
0*
09
0>
0C
#230270000000
1!
1*
b1 6
19
1>
1C
b1 G
#230280000000
0!
0*
09
0>
0C
#230290000000
1!
1*
b10 6
19
1>
1C
b10 G
#230300000000
0!
0*
09
0>
0C
#230310000000
1!
1*
b11 6
19
1>
1C
b11 G
#230320000000
0!
0*
09
0>
0C
#230330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#230340000000
0!
0*
09
0>
0C
#230350000000
1!
1*
b101 6
19
1>
1C
b101 G
#230360000000
0!
0*
09
0>
0C
#230370000000
1!
1*
b110 6
19
1>
1C
b110 G
#230380000000
0!
0*
09
0>
0C
#230390000000
1!
1*
b111 6
19
1>
1C
b111 G
#230400000000
0!
0*
09
0>
0C
#230410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#230420000000
0!
0*
09
0>
0C
#230430000000
1!
1*
b1 6
19
1>
1C
b1 G
#230440000000
0!
0*
09
0>
0C
#230450000000
1!
1*
b10 6
19
1>
1C
b10 G
#230460000000
0!
0*
09
0>
0C
#230470000000
1!
1*
b11 6
19
1>
1C
b11 G
#230480000000
0!
0*
09
0>
0C
#230490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#230500000000
0!
0*
09
0>
0C
#230510000000
1!
1*
b101 6
19
1>
1C
b101 G
#230520000000
0!
0*
09
0>
0C
#230530000000
1!
1*
b110 6
19
1>
1C
b110 G
#230540000000
0!
0*
09
0>
0C
#230550000000
1!
1*
b111 6
19
1>
1C
b111 G
#230560000000
0!
1"
0*
1+
09
1:
0>
0C
#230570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#230580000000
0!
0*
09
0>
0C
#230590000000
1!
1*
b1 6
19
1>
1C
b1 G
#230600000000
0!
0*
09
0>
0C
#230610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#230620000000
0!
0*
09
0>
0C
#230630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#230640000000
0!
0*
09
0>
0C
#230650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#230660000000
0!
0*
09
0>
0C
#230670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#230680000000
0!
0#
0*
0,
09
0>
0?
0C
#230690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#230700000000
0!
0*
09
0>
0C
#230710000000
1!
1*
19
1>
1C
#230720000000
0!
0*
09
0>
0C
#230730000000
1!
1*
19
1>
1C
#230740000000
0!
0*
09
0>
0C
#230750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#230760000000
0!
0*
09
0>
0C
#230770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#230780000000
0!
0*
09
0>
0C
#230790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#230800000000
0!
0*
09
0>
0C
#230810000000
1!
1*
b10 6
19
1>
1C
b10 G
#230820000000
0!
0*
09
0>
0C
#230830000000
1!
1*
b11 6
19
1>
1C
b11 G
#230840000000
0!
0*
09
0>
0C
#230850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#230860000000
0!
0*
09
0>
0C
#230870000000
1!
1*
b101 6
19
1>
1C
b101 G
#230880000000
0!
0*
09
0>
0C
#230890000000
1!
1*
b110 6
19
1>
1C
b110 G
#230900000000
0!
0*
09
0>
0C
#230910000000
1!
1*
b111 6
19
1>
1C
b111 G
#230920000000
0!
0*
09
0>
0C
#230930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#230940000000
0!
0*
09
0>
0C
#230950000000
1!
1*
b1 6
19
1>
1C
b1 G
#230960000000
0!
0*
09
0>
0C
#230970000000
1!
1*
b10 6
19
1>
1C
b10 G
#230980000000
0!
0*
09
0>
0C
#230990000000
1!
1*
b11 6
19
1>
1C
b11 G
#231000000000
0!
0*
09
0>
0C
#231010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#231020000000
0!
0*
09
0>
0C
#231030000000
1!
1*
b101 6
19
1>
1C
b101 G
#231040000000
0!
0*
09
0>
0C
#231050000000
1!
1*
b110 6
19
1>
1C
b110 G
#231060000000
0!
0*
09
0>
0C
#231070000000
1!
1*
b111 6
19
1>
1C
b111 G
#231080000000
0!
0*
09
0>
0C
#231090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#231100000000
0!
0*
09
0>
0C
#231110000000
1!
1*
b1 6
19
1>
1C
b1 G
#231120000000
0!
0*
09
0>
0C
#231130000000
1!
1*
b10 6
19
1>
1C
b10 G
#231140000000
0!
0*
09
0>
0C
#231150000000
1!
1*
b11 6
19
1>
1C
b11 G
#231160000000
0!
0*
09
0>
0C
#231170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#231180000000
0!
0*
09
0>
0C
#231190000000
1!
1*
b101 6
19
1>
1C
b101 G
#231200000000
0!
0*
09
0>
0C
#231210000000
1!
1*
b110 6
19
1>
1C
b110 G
#231220000000
0!
0*
09
0>
0C
#231230000000
1!
1*
b111 6
19
1>
1C
b111 G
#231240000000
0!
1"
0*
1+
09
1:
0>
0C
#231250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#231260000000
0!
0*
09
0>
0C
#231270000000
1!
1*
b1 6
19
1>
1C
b1 G
#231280000000
0!
0*
09
0>
0C
#231290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#231300000000
0!
0*
09
0>
0C
#231310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#231320000000
0!
0*
09
0>
0C
#231330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#231340000000
0!
0*
09
0>
0C
#231350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#231360000000
0!
0#
0*
0,
09
0>
0?
0C
#231370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#231380000000
0!
0*
09
0>
0C
#231390000000
1!
1*
19
1>
1C
#231400000000
0!
0*
09
0>
0C
#231410000000
1!
1*
19
1>
1C
#231420000000
0!
0*
09
0>
0C
#231430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#231440000000
0!
0*
09
0>
0C
#231450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#231460000000
0!
0*
09
0>
0C
#231470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#231480000000
0!
0*
09
0>
0C
#231490000000
1!
1*
b10 6
19
1>
1C
b10 G
#231500000000
0!
0*
09
0>
0C
#231510000000
1!
1*
b11 6
19
1>
1C
b11 G
#231520000000
0!
0*
09
0>
0C
#231530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#231540000000
0!
0*
09
0>
0C
#231550000000
1!
1*
b101 6
19
1>
1C
b101 G
#231560000000
0!
0*
09
0>
0C
#231570000000
1!
1*
b110 6
19
1>
1C
b110 G
#231580000000
0!
0*
09
0>
0C
#231590000000
1!
1*
b111 6
19
1>
1C
b111 G
#231600000000
0!
0*
09
0>
0C
#231610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#231620000000
0!
0*
09
0>
0C
#231630000000
1!
1*
b1 6
19
1>
1C
b1 G
#231640000000
0!
0*
09
0>
0C
#231650000000
1!
1*
b10 6
19
1>
1C
b10 G
#231660000000
0!
0*
09
0>
0C
#231670000000
1!
1*
b11 6
19
1>
1C
b11 G
#231680000000
0!
0*
09
0>
0C
#231690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#231700000000
0!
0*
09
0>
0C
#231710000000
1!
1*
b101 6
19
1>
1C
b101 G
#231720000000
0!
0*
09
0>
0C
#231730000000
1!
1*
b110 6
19
1>
1C
b110 G
#231740000000
0!
0*
09
0>
0C
#231750000000
1!
1*
b111 6
19
1>
1C
b111 G
#231760000000
0!
0*
09
0>
0C
#231770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#231780000000
0!
0*
09
0>
0C
#231790000000
1!
1*
b1 6
19
1>
1C
b1 G
#231800000000
0!
0*
09
0>
0C
#231810000000
1!
1*
b10 6
19
1>
1C
b10 G
#231820000000
0!
0*
09
0>
0C
#231830000000
1!
1*
b11 6
19
1>
1C
b11 G
#231840000000
0!
0*
09
0>
0C
#231850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#231860000000
0!
0*
09
0>
0C
#231870000000
1!
1*
b101 6
19
1>
1C
b101 G
#231880000000
0!
0*
09
0>
0C
#231890000000
1!
1*
b110 6
19
1>
1C
b110 G
#231900000000
0!
0*
09
0>
0C
#231910000000
1!
1*
b111 6
19
1>
1C
b111 G
#231920000000
0!
1"
0*
1+
09
1:
0>
0C
#231930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#231940000000
0!
0*
09
0>
0C
#231950000000
1!
1*
b1 6
19
1>
1C
b1 G
#231960000000
0!
0*
09
0>
0C
#231970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#231980000000
0!
0*
09
0>
0C
#231990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#232000000000
0!
0*
09
0>
0C
#232010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#232020000000
0!
0*
09
0>
0C
#232030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#232040000000
0!
0#
0*
0,
09
0>
0?
0C
#232050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#232060000000
0!
0*
09
0>
0C
#232070000000
1!
1*
19
1>
1C
#232080000000
0!
0*
09
0>
0C
#232090000000
1!
1*
19
1>
1C
#232100000000
0!
0*
09
0>
0C
#232110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#232120000000
0!
0*
09
0>
0C
#232130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#232140000000
0!
0*
09
0>
0C
#232150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#232160000000
0!
0*
09
0>
0C
#232170000000
1!
1*
b10 6
19
1>
1C
b10 G
#232180000000
0!
0*
09
0>
0C
#232190000000
1!
1*
b11 6
19
1>
1C
b11 G
#232200000000
0!
0*
09
0>
0C
#232210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#232220000000
0!
0*
09
0>
0C
#232230000000
1!
1*
b101 6
19
1>
1C
b101 G
#232240000000
0!
0*
09
0>
0C
#232250000000
1!
1*
b110 6
19
1>
1C
b110 G
#232260000000
0!
0*
09
0>
0C
#232270000000
1!
1*
b111 6
19
1>
1C
b111 G
#232280000000
0!
0*
09
0>
0C
#232290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#232300000000
0!
0*
09
0>
0C
#232310000000
1!
1*
b1 6
19
1>
1C
b1 G
#232320000000
0!
0*
09
0>
0C
#232330000000
1!
1*
b10 6
19
1>
1C
b10 G
#232340000000
0!
0*
09
0>
0C
#232350000000
1!
1*
b11 6
19
1>
1C
b11 G
#232360000000
0!
0*
09
0>
0C
#232370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#232380000000
0!
0*
09
0>
0C
#232390000000
1!
1*
b101 6
19
1>
1C
b101 G
#232400000000
0!
0*
09
0>
0C
#232410000000
1!
1*
b110 6
19
1>
1C
b110 G
#232420000000
0!
0*
09
0>
0C
#232430000000
1!
1*
b111 6
19
1>
1C
b111 G
#232440000000
0!
0*
09
0>
0C
#232450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#232460000000
0!
0*
09
0>
0C
#232470000000
1!
1*
b1 6
19
1>
1C
b1 G
#232480000000
0!
0*
09
0>
0C
#232490000000
1!
1*
b10 6
19
1>
1C
b10 G
#232500000000
0!
0*
09
0>
0C
#232510000000
1!
1*
b11 6
19
1>
1C
b11 G
#232520000000
0!
0*
09
0>
0C
#232530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#232540000000
0!
0*
09
0>
0C
#232550000000
1!
1*
b101 6
19
1>
1C
b101 G
#232560000000
0!
0*
09
0>
0C
#232570000000
1!
1*
b110 6
19
1>
1C
b110 G
#232580000000
0!
0*
09
0>
0C
#232590000000
1!
1*
b111 6
19
1>
1C
b111 G
#232600000000
0!
1"
0*
1+
09
1:
0>
0C
#232610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#232620000000
0!
0*
09
0>
0C
#232630000000
1!
1*
b1 6
19
1>
1C
b1 G
#232640000000
0!
0*
09
0>
0C
#232650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#232660000000
0!
0*
09
0>
0C
#232670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#232680000000
0!
0*
09
0>
0C
#232690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#232700000000
0!
0*
09
0>
0C
#232710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#232720000000
0!
0#
0*
0,
09
0>
0?
0C
#232730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#232740000000
0!
0*
09
0>
0C
#232750000000
1!
1*
19
1>
1C
#232760000000
0!
0*
09
0>
0C
#232770000000
1!
1*
19
1>
1C
#232780000000
0!
0*
09
0>
0C
#232790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#232800000000
0!
0*
09
0>
0C
#232810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#232820000000
0!
0*
09
0>
0C
#232830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#232840000000
0!
0*
09
0>
0C
#232850000000
1!
1*
b10 6
19
1>
1C
b10 G
#232860000000
0!
0*
09
0>
0C
#232870000000
1!
1*
b11 6
19
1>
1C
b11 G
#232880000000
0!
0*
09
0>
0C
#232890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#232900000000
0!
0*
09
0>
0C
#232910000000
1!
1*
b101 6
19
1>
1C
b101 G
#232920000000
0!
0*
09
0>
0C
#232930000000
1!
1*
b110 6
19
1>
1C
b110 G
#232940000000
0!
0*
09
0>
0C
#232950000000
1!
1*
b111 6
19
1>
1C
b111 G
#232960000000
0!
0*
09
0>
0C
#232970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#232980000000
0!
0*
09
0>
0C
#232990000000
1!
1*
b1 6
19
1>
1C
b1 G
#233000000000
0!
0*
09
0>
0C
#233010000000
1!
1*
b10 6
19
1>
1C
b10 G
#233020000000
0!
0*
09
0>
0C
#233030000000
1!
1*
b11 6
19
1>
1C
b11 G
#233040000000
0!
0*
09
0>
0C
#233050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#233060000000
0!
0*
09
0>
0C
#233070000000
1!
1*
b101 6
19
1>
1C
b101 G
#233080000000
0!
0*
09
0>
0C
#233090000000
1!
1*
b110 6
19
1>
1C
b110 G
#233100000000
0!
0*
09
0>
0C
#233110000000
1!
1*
b111 6
19
1>
1C
b111 G
#233120000000
0!
0*
09
0>
0C
#233130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#233140000000
0!
0*
09
0>
0C
#233150000000
1!
1*
b1 6
19
1>
1C
b1 G
#233160000000
0!
0*
09
0>
0C
#233170000000
1!
1*
b10 6
19
1>
1C
b10 G
#233180000000
0!
0*
09
0>
0C
#233190000000
1!
1*
b11 6
19
1>
1C
b11 G
#233200000000
0!
0*
09
0>
0C
#233210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#233220000000
0!
0*
09
0>
0C
#233230000000
1!
1*
b101 6
19
1>
1C
b101 G
#233240000000
0!
0*
09
0>
0C
#233250000000
1!
1*
b110 6
19
1>
1C
b110 G
#233260000000
0!
0*
09
0>
0C
#233270000000
1!
1*
b111 6
19
1>
1C
b111 G
#233280000000
0!
1"
0*
1+
09
1:
0>
0C
#233290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#233300000000
0!
0*
09
0>
0C
#233310000000
1!
1*
b1 6
19
1>
1C
b1 G
#233320000000
0!
0*
09
0>
0C
#233330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#233340000000
0!
0*
09
0>
0C
#233350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#233360000000
0!
0*
09
0>
0C
#233370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#233380000000
0!
0*
09
0>
0C
#233390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#233400000000
0!
0#
0*
0,
09
0>
0?
0C
#233410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#233420000000
0!
0*
09
0>
0C
#233430000000
1!
1*
19
1>
1C
#233440000000
0!
0*
09
0>
0C
#233450000000
1!
1*
19
1>
1C
#233460000000
0!
0*
09
0>
0C
#233470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#233480000000
0!
0*
09
0>
0C
#233490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#233500000000
0!
0*
09
0>
0C
#233510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#233520000000
0!
0*
09
0>
0C
#233530000000
1!
1*
b10 6
19
1>
1C
b10 G
#233540000000
0!
0*
09
0>
0C
#233550000000
1!
1*
b11 6
19
1>
1C
b11 G
#233560000000
0!
0*
09
0>
0C
#233570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#233580000000
0!
0*
09
0>
0C
#233590000000
1!
1*
b101 6
19
1>
1C
b101 G
#233600000000
0!
0*
09
0>
0C
#233610000000
1!
1*
b110 6
19
1>
1C
b110 G
#233620000000
0!
0*
09
0>
0C
#233630000000
1!
1*
b111 6
19
1>
1C
b111 G
#233640000000
0!
0*
09
0>
0C
#233650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#233660000000
0!
0*
09
0>
0C
#233670000000
1!
1*
b1 6
19
1>
1C
b1 G
#233680000000
0!
0*
09
0>
0C
#233690000000
1!
1*
b10 6
19
1>
1C
b10 G
#233700000000
0!
0*
09
0>
0C
#233710000000
1!
1*
b11 6
19
1>
1C
b11 G
#233720000000
0!
0*
09
0>
0C
#233730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#233740000000
0!
0*
09
0>
0C
#233750000000
1!
1*
b101 6
19
1>
1C
b101 G
#233760000000
0!
0*
09
0>
0C
#233770000000
1!
1*
b110 6
19
1>
1C
b110 G
#233780000000
0!
0*
09
0>
0C
#233790000000
1!
1*
b111 6
19
1>
1C
b111 G
#233800000000
0!
0*
09
0>
0C
#233810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#233820000000
0!
0*
09
0>
0C
#233830000000
1!
1*
b1 6
19
1>
1C
b1 G
#233840000000
0!
0*
09
0>
0C
#233850000000
1!
1*
b10 6
19
1>
1C
b10 G
#233860000000
0!
0*
09
0>
0C
#233870000000
1!
1*
b11 6
19
1>
1C
b11 G
#233880000000
0!
0*
09
0>
0C
#233890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#233900000000
0!
0*
09
0>
0C
#233910000000
1!
1*
b101 6
19
1>
1C
b101 G
#233920000000
0!
0*
09
0>
0C
#233930000000
1!
1*
b110 6
19
1>
1C
b110 G
#233940000000
0!
0*
09
0>
0C
#233950000000
1!
1*
b111 6
19
1>
1C
b111 G
#233960000000
0!
1"
0*
1+
09
1:
0>
0C
#233970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#233980000000
0!
0*
09
0>
0C
#233990000000
1!
1*
b1 6
19
1>
1C
b1 G
#234000000000
0!
0*
09
0>
0C
#234010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#234020000000
0!
0*
09
0>
0C
#234030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#234040000000
0!
0*
09
0>
0C
#234050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#234060000000
0!
0*
09
0>
0C
#234070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#234080000000
0!
0#
0*
0,
09
0>
0?
0C
#234090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#234100000000
0!
0*
09
0>
0C
#234110000000
1!
1*
19
1>
1C
#234120000000
0!
0*
09
0>
0C
#234130000000
1!
1*
19
1>
1C
#234140000000
0!
0*
09
0>
0C
#234150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#234160000000
0!
0*
09
0>
0C
#234170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#234180000000
0!
0*
09
0>
0C
#234190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#234200000000
0!
0*
09
0>
0C
#234210000000
1!
1*
b10 6
19
1>
1C
b10 G
#234220000000
0!
0*
09
0>
0C
#234230000000
1!
1*
b11 6
19
1>
1C
b11 G
#234240000000
0!
0*
09
0>
0C
#234250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#234260000000
0!
0*
09
0>
0C
#234270000000
1!
1*
b101 6
19
1>
1C
b101 G
#234280000000
0!
0*
09
0>
0C
#234290000000
1!
1*
b110 6
19
1>
1C
b110 G
#234300000000
0!
0*
09
0>
0C
#234310000000
1!
1*
b111 6
19
1>
1C
b111 G
#234320000000
0!
0*
09
0>
0C
#234330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#234340000000
0!
0*
09
0>
0C
#234350000000
1!
1*
b1 6
19
1>
1C
b1 G
#234360000000
0!
0*
09
0>
0C
#234370000000
1!
1*
b10 6
19
1>
1C
b10 G
#234380000000
0!
0*
09
0>
0C
#234390000000
1!
1*
b11 6
19
1>
1C
b11 G
#234400000000
0!
0*
09
0>
0C
#234410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#234420000000
0!
0*
09
0>
0C
#234430000000
1!
1*
b101 6
19
1>
1C
b101 G
#234440000000
0!
0*
09
0>
0C
#234450000000
1!
1*
b110 6
19
1>
1C
b110 G
#234460000000
0!
0*
09
0>
0C
#234470000000
1!
1*
b111 6
19
1>
1C
b111 G
#234480000000
0!
0*
09
0>
0C
#234490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#234500000000
0!
0*
09
0>
0C
#234510000000
1!
1*
b1 6
19
1>
1C
b1 G
#234520000000
0!
0*
09
0>
0C
#234530000000
1!
1*
b10 6
19
1>
1C
b10 G
#234540000000
0!
0*
09
0>
0C
#234550000000
1!
1*
b11 6
19
1>
1C
b11 G
#234560000000
0!
0*
09
0>
0C
#234570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#234580000000
0!
0*
09
0>
0C
#234590000000
1!
1*
b101 6
19
1>
1C
b101 G
#234600000000
0!
0*
09
0>
0C
#234610000000
1!
1*
b110 6
19
1>
1C
b110 G
#234620000000
0!
0*
09
0>
0C
#234630000000
1!
1*
b111 6
19
1>
1C
b111 G
#234640000000
0!
1"
0*
1+
09
1:
0>
0C
#234650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#234660000000
0!
0*
09
0>
0C
#234670000000
1!
1*
b1 6
19
1>
1C
b1 G
#234680000000
0!
0*
09
0>
0C
#234690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#234700000000
0!
0*
09
0>
0C
#234710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#234720000000
0!
0*
09
0>
0C
#234730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#234740000000
0!
0*
09
0>
0C
#234750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#234760000000
0!
0#
0*
0,
09
0>
0?
0C
#234770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#234780000000
0!
0*
09
0>
0C
#234790000000
1!
1*
19
1>
1C
#234800000000
0!
0*
09
0>
0C
#234810000000
1!
1*
19
1>
1C
#234820000000
0!
0*
09
0>
0C
#234830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#234840000000
0!
0*
09
0>
0C
#234850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#234860000000
0!
0*
09
0>
0C
#234870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#234880000000
0!
0*
09
0>
0C
#234890000000
1!
1*
b10 6
19
1>
1C
b10 G
#234900000000
0!
0*
09
0>
0C
#234910000000
1!
1*
b11 6
19
1>
1C
b11 G
#234920000000
0!
0*
09
0>
0C
#234930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#234940000000
0!
0*
09
0>
0C
#234950000000
1!
1*
b101 6
19
1>
1C
b101 G
#234960000000
0!
0*
09
0>
0C
#234970000000
1!
1*
b110 6
19
1>
1C
b110 G
#234980000000
0!
0*
09
0>
0C
#234990000000
1!
1*
b111 6
19
1>
1C
b111 G
#235000000000
0!
0*
09
0>
0C
#235010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#235020000000
0!
0*
09
0>
0C
#235030000000
1!
1*
b1 6
19
1>
1C
b1 G
#235040000000
0!
0*
09
0>
0C
#235050000000
1!
1*
b10 6
19
1>
1C
b10 G
#235060000000
0!
0*
09
0>
0C
#235070000000
1!
1*
b11 6
19
1>
1C
b11 G
#235080000000
0!
0*
09
0>
0C
#235090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#235100000000
0!
0*
09
0>
0C
#235110000000
1!
1*
b101 6
19
1>
1C
b101 G
#235120000000
0!
0*
09
0>
0C
#235130000000
1!
1*
b110 6
19
1>
1C
b110 G
#235140000000
0!
0*
09
0>
0C
#235150000000
1!
1*
b111 6
19
1>
1C
b111 G
#235160000000
0!
0*
09
0>
0C
#235170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#235180000000
0!
0*
09
0>
0C
#235190000000
1!
1*
b1 6
19
1>
1C
b1 G
#235200000000
0!
0*
09
0>
0C
#235210000000
1!
1*
b10 6
19
1>
1C
b10 G
#235220000000
0!
0*
09
0>
0C
#235230000000
1!
1*
b11 6
19
1>
1C
b11 G
#235240000000
0!
0*
09
0>
0C
#235250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#235260000000
0!
0*
09
0>
0C
#235270000000
1!
1*
b101 6
19
1>
1C
b101 G
#235280000000
0!
0*
09
0>
0C
#235290000000
1!
1*
b110 6
19
1>
1C
b110 G
#235300000000
0!
0*
09
0>
0C
#235310000000
1!
1*
b111 6
19
1>
1C
b111 G
#235320000000
0!
1"
0*
1+
09
1:
0>
0C
#235330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#235340000000
0!
0*
09
0>
0C
#235350000000
1!
1*
b1 6
19
1>
1C
b1 G
#235360000000
0!
0*
09
0>
0C
#235370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#235380000000
0!
0*
09
0>
0C
#235390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#235400000000
0!
0*
09
0>
0C
#235410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#235420000000
0!
0*
09
0>
0C
#235430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#235440000000
0!
0#
0*
0,
09
0>
0?
0C
#235450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#235460000000
0!
0*
09
0>
0C
#235470000000
1!
1*
19
1>
1C
#235480000000
0!
0*
09
0>
0C
#235490000000
1!
1*
19
1>
1C
#235500000000
0!
0*
09
0>
0C
#235510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#235520000000
0!
0*
09
0>
0C
#235530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#235540000000
0!
0*
09
0>
0C
#235550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#235560000000
0!
0*
09
0>
0C
#235570000000
1!
1*
b10 6
19
1>
1C
b10 G
#235580000000
0!
0*
09
0>
0C
#235590000000
1!
1*
b11 6
19
1>
1C
b11 G
#235600000000
0!
0*
09
0>
0C
#235610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#235620000000
0!
0*
09
0>
0C
#235630000000
1!
1*
b101 6
19
1>
1C
b101 G
#235640000000
0!
0*
09
0>
0C
#235650000000
1!
1*
b110 6
19
1>
1C
b110 G
#235660000000
0!
0*
09
0>
0C
#235670000000
1!
1*
b111 6
19
1>
1C
b111 G
#235680000000
0!
0*
09
0>
0C
#235690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#235700000000
0!
0*
09
0>
0C
#235710000000
1!
1*
b1 6
19
1>
1C
b1 G
#235720000000
0!
0*
09
0>
0C
#235730000000
1!
1*
b10 6
19
1>
1C
b10 G
#235740000000
0!
0*
09
0>
0C
#235750000000
1!
1*
b11 6
19
1>
1C
b11 G
#235760000000
0!
0*
09
0>
0C
#235770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#235780000000
0!
0*
09
0>
0C
#235790000000
1!
1*
b101 6
19
1>
1C
b101 G
#235800000000
0!
0*
09
0>
0C
#235810000000
1!
1*
b110 6
19
1>
1C
b110 G
#235820000000
0!
0*
09
0>
0C
#235830000000
1!
1*
b111 6
19
1>
1C
b111 G
#235840000000
0!
0*
09
0>
0C
#235850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#235860000000
0!
0*
09
0>
0C
#235870000000
1!
1*
b1 6
19
1>
1C
b1 G
#235880000000
0!
0*
09
0>
0C
#235890000000
1!
1*
b10 6
19
1>
1C
b10 G
#235900000000
0!
0*
09
0>
0C
#235910000000
1!
1*
b11 6
19
1>
1C
b11 G
#235920000000
0!
0*
09
0>
0C
#235930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#235940000000
0!
0*
09
0>
0C
#235950000000
1!
1*
b101 6
19
1>
1C
b101 G
#235960000000
0!
0*
09
0>
0C
#235970000000
1!
1*
b110 6
19
1>
1C
b110 G
#235980000000
0!
0*
09
0>
0C
#235990000000
1!
1*
b111 6
19
1>
1C
b111 G
#236000000000
0!
1"
0*
1+
09
1:
0>
0C
#236010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#236020000000
0!
0*
09
0>
0C
#236030000000
1!
1*
b1 6
19
1>
1C
b1 G
#236040000000
0!
0*
09
0>
0C
#236050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#236060000000
0!
0*
09
0>
0C
#236070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#236080000000
0!
0*
09
0>
0C
#236090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#236100000000
0!
0*
09
0>
0C
#236110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#236120000000
0!
0#
0*
0,
09
0>
0?
0C
#236130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#236140000000
0!
0*
09
0>
0C
#236150000000
1!
1*
19
1>
1C
#236160000000
0!
0*
09
0>
0C
#236170000000
1!
1*
19
1>
1C
#236180000000
0!
0*
09
0>
0C
#236190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#236200000000
0!
0*
09
0>
0C
#236210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#236220000000
0!
0*
09
0>
0C
#236230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#236240000000
0!
0*
09
0>
0C
#236250000000
1!
1*
b10 6
19
1>
1C
b10 G
#236260000000
0!
0*
09
0>
0C
#236270000000
1!
1*
b11 6
19
1>
1C
b11 G
#236280000000
0!
0*
09
0>
0C
#236290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#236300000000
0!
0*
09
0>
0C
#236310000000
1!
1*
b101 6
19
1>
1C
b101 G
#236320000000
0!
0*
09
0>
0C
#236330000000
1!
1*
b110 6
19
1>
1C
b110 G
#236340000000
0!
0*
09
0>
0C
#236350000000
1!
1*
b111 6
19
1>
1C
b111 G
#236360000000
0!
0*
09
0>
0C
#236370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#236380000000
0!
0*
09
0>
0C
#236390000000
1!
1*
b1 6
19
1>
1C
b1 G
#236400000000
0!
0*
09
0>
0C
#236410000000
1!
1*
b10 6
19
1>
1C
b10 G
#236420000000
0!
0*
09
0>
0C
#236430000000
1!
1*
b11 6
19
1>
1C
b11 G
#236440000000
0!
0*
09
0>
0C
#236450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#236460000000
0!
0*
09
0>
0C
#236470000000
1!
1*
b101 6
19
1>
1C
b101 G
#236480000000
0!
0*
09
0>
0C
#236490000000
1!
1*
b110 6
19
1>
1C
b110 G
#236500000000
0!
0*
09
0>
0C
#236510000000
1!
1*
b111 6
19
1>
1C
b111 G
#236520000000
0!
0*
09
0>
0C
#236530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#236540000000
0!
0*
09
0>
0C
#236550000000
1!
1*
b1 6
19
1>
1C
b1 G
#236560000000
0!
0*
09
0>
0C
#236570000000
1!
1*
b10 6
19
1>
1C
b10 G
#236580000000
0!
0*
09
0>
0C
#236590000000
1!
1*
b11 6
19
1>
1C
b11 G
#236600000000
0!
0*
09
0>
0C
#236610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#236620000000
0!
0*
09
0>
0C
#236630000000
1!
1*
b101 6
19
1>
1C
b101 G
#236640000000
0!
0*
09
0>
0C
#236650000000
1!
1*
b110 6
19
1>
1C
b110 G
#236660000000
0!
0*
09
0>
0C
#236670000000
1!
1*
b111 6
19
1>
1C
b111 G
#236680000000
0!
1"
0*
1+
09
1:
0>
0C
#236690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#236700000000
0!
0*
09
0>
0C
#236710000000
1!
1*
b1 6
19
1>
1C
b1 G
#236720000000
0!
0*
09
0>
0C
#236730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#236740000000
0!
0*
09
0>
0C
#236750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#236760000000
0!
0*
09
0>
0C
#236770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#236780000000
0!
0*
09
0>
0C
#236790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#236800000000
0!
0#
0*
0,
09
0>
0?
0C
#236810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#236820000000
0!
0*
09
0>
0C
#236830000000
1!
1*
19
1>
1C
#236840000000
0!
0*
09
0>
0C
#236850000000
1!
1*
19
1>
1C
#236860000000
0!
0*
09
0>
0C
#236870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#236880000000
0!
0*
09
0>
0C
#236890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#236900000000
0!
0*
09
0>
0C
#236910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#236920000000
0!
0*
09
0>
0C
#236930000000
1!
1*
b10 6
19
1>
1C
b10 G
#236940000000
0!
0*
09
0>
0C
#236950000000
1!
1*
b11 6
19
1>
1C
b11 G
#236960000000
0!
0*
09
0>
0C
#236970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#236980000000
0!
0*
09
0>
0C
#236990000000
1!
1*
b101 6
19
1>
1C
b101 G
#237000000000
0!
0*
09
0>
0C
#237010000000
1!
1*
b110 6
19
1>
1C
b110 G
#237020000000
0!
0*
09
0>
0C
#237030000000
1!
1*
b111 6
19
1>
1C
b111 G
#237040000000
0!
0*
09
0>
0C
#237050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#237060000000
0!
0*
09
0>
0C
#237070000000
1!
1*
b1 6
19
1>
1C
b1 G
#237080000000
0!
0*
09
0>
0C
#237090000000
1!
1*
b10 6
19
1>
1C
b10 G
#237100000000
0!
0*
09
0>
0C
#237110000000
1!
1*
b11 6
19
1>
1C
b11 G
#237120000000
0!
0*
09
0>
0C
#237130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#237140000000
0!
0*
09
0>
0C
#237150000000
1!
1*
b101 6
19
1>
1C
b101 G
#237160000000
0!
0*
09
0>
0C
#237170000000
1!
1*
b110 6
19
1>
1C
b110 G
#237180000000
0!
0*
09
0>
0C
#237190000000
1!
1*
b111 6
19
1>
1C
b111 G
#237200000000
0!
0*
09
0>
0C
#237210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#237220000000
0!
0*
09
0>
0C
#237230000000
1!
1*
b1 6
19
1>
1C
b1 G
#237240000000
0!
0*
09
0>
0C
#237250000000
1!
1*
b10 6
19
1>
1C
b10 G
#237260000000
0!
0*
09
0>
0C
#237270000000
1!
1*
b11 6
19
1>
1C
b11 G
#237280000000
0!
0*
09
0>
0C
#237290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#237300000000
0!
0*
09
0>
0C
#237310000000
1!
1*
b101 6
19
1>
1C
b101 G
#237320000000
0!
0*
09
0>
0C
#237330000000
1!
1*
b110 6
19
1>
1C
b110 G
#237340000000
0!
0*
09
0>
0C
#237350000000
1!
1*
b111 6
19
1>
1C
b111 G
#237360000000
0!
1"
0*
1+
09
1:
0>
0C
#237370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#237380000000
0!
0*
09
0>
0C
#237390000000
1!
1*
b1 6
19
1>
1C
b1 G
#237400000000
0!
0*
09
0>
0C
#237410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#237420000000
0!
0*
09
0>
0C
#237430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#237440000000
0!
0*
09
0>
0C
#237450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#237460000000
0!
0*
09
0>
0C
#237470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#237480000000
0!
0#
0*
0,
09
0>
0?
0C
#237490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#237500000000
0!
0*
09
0>
0C
#237510000000
1!
1*
19
1>
1C
#237520000000
0!
0*
09
0>
0C
#237530000000
1!
1*
19
1>
1C
#237540000000
0!
0*
09
0>
0C
#237550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#237560000000
0!
0*
09
0>
0C
#237570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#237580000000
0!
0*
09
0>
0C
#237590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#237600000000
0!
0*
09
0>
0C
#237610000000
1!
1*
b10 6
19
1>
1C
b10 G
#237620000000
0!
0*
09
0>
0C
#237630000000
1!
1*
b11 6
19
1>
1C
b11 G
#237640000000
0!
0*
09
0>
0C
#237650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#237660000000
0!
0*
09
0>
0C
#237670000000
1!
1*
b101 6
19
1>
1C
b101 G
#237680000000
0!
0*
09
0>
0C
#237690000000
1!
1*
b110 6
19
1>
1C
b110 G
#237700000000
0!
0*
09
0>
0C
#237710000000
1!
1*
b111 6
19
1>
1C
b111 G
#237720000000
0!
0*
09
0>
0C
#237730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#237740000000
0!
0*
09
0>
0C
#237750000000
1!
1*
b1 6
19
1>
1C
b1 G
#237760000000
0!
0*
09
0>
0C
#237770000000
1!
1*
b10 6
19
1>
1C
b10 G
#237780000000
0!
0*
09
0>
0C
#237790000000
1!
1*
b11 6
19
1>
1C
b11 G
#237800000000
0!
0*
09
0>
0C
#237810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#237820000000
0!
0*
09
0>
0C
#237830000000
1!
1*
b101 6
19
1>
1C
b101 G
#237840000000
0!
0*
09
0>
0C
#237850000000
1!
1*
b110 6
19
1>
1C
b110 G
#237860000000
0!
0*
09
0>
0C
#237870000000
1!
1*
b111 6
19
1>
1C
b111 G
#237880000000
0!
0*
09
0>
0C
#237890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#237900000000
0!
0*
09
0>
0C
#237910000000
1!
1*
b1 6
19
1>
1C
b1 G
#237920000000
0!
0*
09
0>
0C
#237930000000
1!
1*
b10 6
19
1>
1C
b10 G
#237940000000
0!
0*
09
0>
0C
#237950000000
1!
1*
b11 6
19
1>
1C
b11 G
#237960000000
0!
0*
09
0>
0C
#237970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#237980000000
0!
0*
09
0>
0C
#237990000000
1!
1*
b101 6
19
1>
1C
b101 G
#238000000000
0!
0*
09
0>
0C
#238010000000
1!
1*
b110 6
19
1>
1C
b110 G
#238020000000
0!
0*
09
0>
0C
#238030000000
1!
1*
b111 6
19
1>
1C
b111 G
#238040000000
0!
1"
0*
1+
09
1:
0>
0C
#238050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#238060000000
0!
0*
09
0>
0C
#238070000000
1!
1*
b1 6
19
1>
1C
b1 G
#238080000000
0!
0*
09
0>
0C
#238090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#238100000000
0!
0*
09
0>
0C
#238110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#238120000000
0!
0*
09
0>
0C
#238130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#238140000000
0!
0*
09
0>
0C
#238150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#238160000000
0!
0#
0*
0,
09
0>
0?
0C
#238170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#238180000000
0!
0*
09
0>
0C
#238190000000
1!
1*
19
1>
1C
#238200000000
0!
0*
09
0>
0C
#238210000000
1!
1*
19
1>
1C
#238220000000
0!
0*
09
0>
0C
#238230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#238240000000
0!
0*
09
0>
0C
#238250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#238260000000
0!
0*
09
0>
0C
#238270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#238280000000
0!
0*
09
0>
0C
#238290000000
1!
1*
b10 6
19
1>
1C
b10 G
#238300000000
0!
0*
09
0>
0C
#238310000000
1!
1*
b11 6
19
1>
1C
b11 G
#238320000000
0!
0*
09
0>
0C
#238330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#238340000000
0!
0*
09
0>
0C
#238350000000
1!
1*
b101 6
19
1>
1C
b101 G
#238360000000
0!
0*
09
0>
0C
#238370000000
1!
1*
b110 6
19
1>
1C
b110 G
#238380000000
0!
0*
09
0>
0C
#238390000000
1!
1*
b111 6
19
1>
1C
b111 G
#238400000000
0!
0*
09
0>
0C
#238410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#238420000000
0!
0*
09
0>
0C
#238430000000
1!
1*
b1 6
19
1>
1C
b1 G
#238440000000
0!
0*
09
0>
0C
#238450000000
1!
1*
b10 6
19
1>
1C
b10 G
#238460000000
0!
0*
09
0>
0C
#238470000000
1!
1*
b11 6
19
1>
1C
b11 G
#238480000000
0!
0*
09
0>
0C
#238490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#238500000000
0!
0*
09
0>
0C
#238510000000
1!
1*
b101 6
19
1>
1C
b101 G
#238520000000
0!
0*
09
0>
0C
#238530000000
1!
1*
b110 6
19
1>
1C
b110 G
#238540000000
0!
0*
09
0>
0C
#238550000000
1!
1*
b111 6
19
1>
1C
b111 G
#238560000000
0!
0*
09
0>
0C
#238570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#238580000000
0!
0*
09
0>
0C
#238590000000
1!
1*
b1 6
19
1>
1C
b1 G
#238600000000
0!
0*
09
0>
0C
#238610000000
1!
1*
b10 6
19
1>
1C
b10 G
#238620000000
0!
0*
09
0>
0C
#238630000000
1!
1*
b11 6
19
1>
1C
b11 G
#238640000000
0!
0*
09
0>
0C
#238650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#238660000000
0!
0*
09
0>
0C
#238670000000
1!
1*
b101 6
19
1>
1C
b101 G
#238680000000
0!
0*
09
0>
0C
#238690000000
1!
1*
b110 6
19
1>
1C
b110 G
#238700000000
0!
0*
09
0>
0C
#238710000000
1!
1*
b111 6
19
1>
1C
b111 G
#238720000000
0!
1"
0*
1+
09
1:
0>
0C
#238730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#238740000000
0!
0*
09
0>
0C
#238750000000
1!
1*
b1 6
19
1>
1C
b1 G
#238760000000
0!
0*
09
0>
0C
#238770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#238780000000
0!
0*
09
0>
0C
#238790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#238800000000
0!
0*
09
0>
0C
#238810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#238820000000
0!
0*
09
0>
0C
#238830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#238840000000
0!
0#
0*
0,
09
0>
0?
0C
#238850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#238860000000
0!
0*
09
0>
0C
#238870000000
1!
1*
19
1>
1C
#238880000000
0!
0*
09
0>
0C
#238890000000
1!
1*
19
1>
1C
#238900000000
0!
0*
09
0>
0C
#238910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#238920000000
0!
0*
09
0>
0C
#238930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#238940000000
0!
0*
09
0>
0C
#238950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#238960000000
0!
0*
09
0>
0C
#238970000000
1!
1*
b10 6
19
1>
1C
b10 G
#238980000000
0!
0*
09
0>
0C
#238990000000
1!
1*
b11 6
19
1>
1C
b11 G
#239000000000
0!
0*
09
0>
0C
#239010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#239020000000
0!
0*
09
0>
0C
#239030000000
1!
1*
b101 6
19
1>
1C
b101 G
#239040000000
0!
0*
09
0>
0C
#239050000000
1!
1*
b110 6
19
1>
1C
b110 G
#239060000000
0!
0*
09
0>
0C
#239070000000
1!
1*
b111 6
19
1>
1C
b111 G
#239080000000
0!
0*
09
0>
0C
#239090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#239100000000
0!
0*
09
0>
0C
#239110000000
1!
1*
b1 6
19
1>
1C
b1 G
#239120000000
0!
0*
09
0>
0C
#239130000000
1!
1*
b10 6
19
1>
1C
b10 G
#239140000000
0!
0*
09
0>
0C
#239150000000
1!
1*
b11 6
19
1>
1C
b11 G
#239160000000
0!
0*
09
0>
0C
#239170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#239180000000
0!
0*
09
0>
0C
#239190000000
1!
1*
b101 6
19
1>
1C
b101 G
#239200000000
0!
0*
09
0>
0C
#239210000000
1!
1*
b110 6
19
1>
1C
b110 G
#239220000000
0!
0*
09
0>
0C
#239230000000
1!
1*
b111 6
19
1>
1C
b111 G
#239240000000
0!
0*
09
0>
0C
#239250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#239260000000
0!
0*
09
0>
0C
#239270000000
1!
1*
b1 6
19
1>
1C
b1 G
#239280000000
0!
0*
09
0>
0C
#239290000000
1!
1*
b10 6
19
1>
1C
b10 G
#239300000000
0!
0*
09
0>
0C
#239310000000
1!
1*
b11 6
19
1>
1C
b11 G
#239320000000
0!
0*
09
0>
0C
#239330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#239340000000
0!
0*
09
0>
0C
#239350000000
1!
1*
b101 6
19
1>
1C
b101 G
#239360000000
0!
0*
09
0>
0C
#239370000000
1!
1*
b110 6
19
1>
1C
b110 G
#239380000000
0!
0*
09
0>
0C
#239390000000
1!
1*
b111 6
19
1>
1C
b111 G
#239400000000
0!
1"
0*
1+
09
1:
0>
0C
#239410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#239420000000
0!
0*
09
0>
0C
#239430000000
1!
1*
b1 6
19
1>
1C
b1 G
#239440000000
0!
0*
09
0>
0C
#239450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#239460000000
0!
0*
09
0>
0C
#239470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#239480000000
0!
0*
09
0>
0C
#239490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#239500000000
0!
0*
09
0>
0C
#239510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#239520000000
0!
0#
0*
0,
09
0>
0?
0C
#239530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#239540000000
0!
0*
09
0>
0C
#239550000000
1!
1*
19
1>
1C
#239560000000
0!
0*
09
0>
0C
#239570000000
1!
1*
19
1>
1C
#239580000000
0!
0*
09
0>
0C
#239590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#239600000000
0!
0*
09
0>
0C
#239610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#239620000000
0!
0*
09
0>
0C
#239630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#239640000000
0!
0*
09
0>
0C
#239650000000
1!
1*
b10 6
19
1>
1C
b10 G
#239660000000
0!
0*
09
0>
0C
#239670000000
1!
1*
b11 6
19
1>
1C
b11 G
#239680000000
0!
0*
09
0>
0C
#239690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#239700000000
0!
0*
09
0>
0C
#239710000000
1!
1*
b101 6
19
1>
1C
b101 G
#239720000000
0!
0*
09
0>
0C
#239730000000
1!
1*
b110 6
19
1>
1C
b110 G
#239740000000
0!
0*
09
0>
0C
#239750000000
1!
1*
b111 6
19
1>
1C
b111 G
#239760000000
0!
0*
09
0>
0C
#239770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#239780000000
0!
0*
09
0>
0C
#239790000000
1!
1*
b1 6
19
1>
1C
b1 G
#239800000000
0!
0*
09
0>
0C
#239810000000
1!
1*
b10 6
19
1>
1C
b10 G
#239820000000
0!
0*
09
0>
0C
#239830000000
1!
1*
b11 6
19
1>
1C
b11 G
#239840000000
0!
0*
09
0>
0C
#239850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#239860000000
0!
0*
09
0>
0C
#239870000000
1!
1*
b101 6
19
1>
1C
b101 G
#239880000000
0!
0*
09
0>
0C
#239890000000
1!
1*
b110 6
19
1>
1C
b110 G
#239900000000
0!
0*
09
0>
0C
#239910000000
1!
1*
b111 6
19
1>
1C
b111 G
#239920000000
0!
0*
09
0>
0C
#239930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#239940000000
0!
0*
09
0>
0C
#239950000000
1!
1*
b1 6
19
1>
1C
b1 G
#239960000000
0!
0*
09
0>
0C
#239970000000
1!
1*
b10 6
19
1>
1C
b10 G
#239980000000
0!
0*
09
0>
0C
#239990000000
1!
1*
b11 6
19
1>
1C
b11 G
#240000000000
0!
0*
09
0>
0C
#240010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#240020000000
0!
0*
09
0>
0C
#240030000000
1!
1*
b101 6
19
1>
1C
b101 G
#240040000000
0!
0*
09
0>
0C
#240050000000
1!
1*
b110 6
19
1>
1C
b110 G
#240060000000
0!
0*
09
0>
0C
#240070000000
1!
1*
b111 6
19
1>
1C
b111 G
#240080000000
0!
1"
0*
1+
09
1:
0>
0C
#240090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#240100000000
0!
0*
09
0>
0C
#240110000000
1!
1*
b1 6
19
1>
1C
b1 G
#240120000000
0!
0*
09
0>
0C
#240130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#240140000000
0!
0*
09
0>
0C
#240150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#240160000000
0!
0*
09
0>
0C
#240170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#240180000000
0!
0*
09
0>
0C
#240190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#240200000000
0!
0#
0*
0,
09
0>
0?
0C
#240210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#240220000000
0!
0*
09
0>
0C
#240230000000
1!
1*
19
1>
1C
#240240000000
0!
0*
09
0>
0C
#240250000000
1!
1*
19
1>
1C
#240260000000
0!
0*
09
0>
0C
#240270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#240280000000
0!
0*
09
0>
0C
#240290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#240300000000
0!
0*
09
0>
0C
#240310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#240320000000
0!
0*
09
0>
0C
#240330000000
1!
1*
b10 6
19
1>
1C
b10 G
#240340000000
0!
0*
09
0>
0C
#240350000000
1!
1*
b11 6
19
1>
1C
b11 G
#240360000000
0!
0*
09
0>
0C
#240370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#240380000000
0!
0*
09
0>
0C
#240390000000
1!
1*
b101 6
19
1>
1C
b101 G
#240400000000
0!
0*
09
0>
0C
#240410000000
1!
1*
b110 6
19
1>
1C
b110 G
#240420000000
0!
0*
09
0>
0C
#240430000000
1!
1*
b111 6
19
1>
1C
b111 G
#240440000000
0!
0*
09
0>
0C
#240450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#240460000000
0!
0*
09
0>
0C
#240470000000
1!
1*
b1 6
19
1>
1C
b1 G
#240480000000
0!
0*
09
0>
0C
#240490000000
1!
1*
b10 6
19
1>
1C
b10 G
#240500000000
0!
0*
09
0>
0C
#240510000000
1!
1*
b11 6
19
1>
1C
b11 G
#240520000000
0!
0*
09
0>
0C
#240530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#240540000000
0!
0*
09
0>
0C
#240550000000
1!
1*
b101 6
19
1>
1C
b101 G
#240560000000
0!
0*
09
0>
0C
#240570000000
1!
1*
b110 6
19
1>
1C
b110 G
#240580000000
0!
0*
09
0>
0C
#240590000000
1!
1*
b111 6
19
1>
1C
b111 G
#240600000000
0!
0*
09
0>
0C
#240610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#240620000000
0!
0*
09
0>
0C
#240630000000
1!
1*
b1 6
19
1>
1C
b1 G
#240640000000
0!
0*
09
0>
0C
#240650000000
1!
1*
b10 6
19
1>
1C
b10 G
#240660000000
0!
0*
09
0>
0C
#240670000000
1!
1*
b11 6
19
1>
1C
b11 G
#240680000000
0!
0*
09
0>
0C
#240690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#240700000000
0!
0*
09
0>
0C
#240710000000
1!
1*
b101 6
19
1>
1C
b101 G
#240720000000
0!
0*
09
0>
0C
#240730000000
1!
1*
b110 6
19
1>
1C
b110 G
#240740000000
0!
0*
09
0>
0C
#240750000000
1!
1*
b111 6
19
1>
1C
b111 G
#240760000000
0!
1"
0*
1+
09
1:
0>
0C
#240770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#240780000000
0!
0*
09
0>
0C
#240790000000
1!
1*
b1 6
19
1>
1C
b1 G
#240800000000
0!
0*
09
0>
0C
#240810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#240820000000
0!
0*
09
0>
0C
#240830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#240840000000
0!
0*
09
0>
0C
#240850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#240860000000
0!
0*
09
0>
0C
#240870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#240880000000
0!
0#
0*
0,
09
0>
0?
0C
#240890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#240900000000
0!
0*
09
0>
0C
#240910000000
1!
1*
19
1>
1C
#240920000000
0!
0*
09
0>
0C
#240930000000
1!
1*
19
1>
1C
#240940000000
0!
0*
09
0>
0C
#240950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#240960000000
0!
0*
09
0>
0C
#240970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#240980000000
0!
0*
09
0>
0C
#240990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#241000000000
0!
0*
09
0>
0C
#241010000000
1!
1*
b10 6
19
1>
1C
b10 G
#241020000000
0!
0*
09
0>
0C
#241030000000
1!
1*
b11 6
19
1>
1C
b11 G
#241040000000
0!
0*
09
0>
0C
#241050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#241060000000
0!
0*
09
0>
0C
#241070000000
1!
1*
b101 6
19
1>
1C
b101 G
#241080000000
0!
0*
09
0>
0C
#241090000000
1!
1*
b110 6
19
1>
1C
b110 G
#241100000000
0!
0*
09
0>
0C
#241110000000
1!
1*
b111 6
19
1>
1C
b111 G
#241120000000
0!
0*
09
0>
0C
#241130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#241140000000
0!
0*
09
0>
0C
#241150000000
1!
1*
b1 6
19
1>
1C
b1 G
#241160000000
0!
0*
09
0>
0C
#241170000000
1!
1*
b10 6
19
1>
1C
b10 G
#241180000000
0!
0*
09
0>
0C
#241190000000
1!
1*
b11 6
19
1>
1C
b11 G
#241200000000
0!
0*
09
0>
0C
#241210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#241220000000
0!
0*
09
0>
0C
#241230000000
1!
1*
b101 6
19
1>
1C
b101 G
#241240000000
0!
0*
09
0>
0C
#241250000000
1!
1*
b110 6
19
1>
1C
b110 G
#241260000000
0!
0*
09
0>
0C
#241270000000
1!
1*
b111 6
19
1>
1C
b111 G
#241280000000
0!
0*
09
0>
0C
#241290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#241300000000
0!
0*
09
0>
0C
#241310000000
1!
1*
b1 6
19
1>
1C
b1 G
#241320000000
0!
0*
09
0>
0C
#241330000000
1!
1*
b10 6
19
1>
1C
b10 G
#241340000000
0!
0*
09
0>
0C
#241350000000
1!
1*
b11 6
19
1>
1C
b11 G
#241360000000
0!
0*
09
0>
0C
#241370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#241380000000
0!
0*
09
0>
0C
#241390000000
1!
1*
b101 6
19
1>
1C
b101 G
#241400000000
0!
0*
09
0>
0C
#241410000000
1!
1*
b110 6
19
1>
1C
b110 G
#241420000000
0!
0*
09
0>
0C
#241430000000
1!
1*
b111 6
19
1>
1C
b111 G
#241440000000
0!
1"
0*
1+
09
1:
0>
0C
#241450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#241460000000
0!
0*
09
0>
0C
#241470000000
1!
1*
b1 6
19
1>
1C
b1 G
#241480000000
0!
0*
09
0>
0C
#241490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#241500000000
0!
0*
09
0>
0C
#241510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#241520000000
0!
0*
09
0>
0C
#241530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#241540000000
0!
0*
09
0>
0C
#241550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#241560000000
0!
0#
0*
0,
09
0>
0?
0C
#241570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#241580000000
0!
0*
09
0>
0C
#241590000000
1!
1*
19
1>
1C
#241600000000
0!
0*
09
0>
0C
#241610000000
1!
1*
19
1>
1C
#241620000000
0!
0*
09
0>
0C
#241630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#241640000000
0!
0*
09
0>
0C
#241650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#241660000000
0!
0*
09
0>
0C
#241670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#241680000000
0!
0*
09
0>
0C
#241690000000
1!
1*
b10 6
19
1>
1C
b10 G
#241700000000
0!
0*
09
0>
0C
#241710000000
1!
1*
b11 6
19
1>
1C
b11 G
#241720000000
0!
0*
09
0>
0C
#241730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#241740000000
0!
0*
09
0>
0C
#241750000000
1!
1*
b101 6
19
1>
1C
b101 G
#241760000000
0!
0*
09
0>
0C
#241770000000
1!
1*
b110 6
19
1>
1C
b110 G
#241780000000
0!
0*
09
0>
0C
#241790000000
1!
1*
b111 6
19
1>
1C
b111 G
#241800000000
0!
0*
09
0>
0C
#241810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#241820000000
0!
0*
09
0>
0C
#241830000000
1!
1*
b1 6
19
1>
1C
b1 G
#241840000000
0!
0*
09
0>
0C
#241850000000
1!
1*
b10 6
19
1>
1C
b10 G
#241860000000
0!
0*
09
0>
0C
#241870000000
1!
1*
b11 6
19
1>
1C
b11 G
#241880000000
0!
0*
09
0>
0C
#241890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#241900000000
0!
0*
09
0>
0C
#241910000000
1!
1*
b101 6
19
1>
1C
b101 G
#241920000000
0!
0*
09
0>
0C
#241930000000
1!
1*
b110 6
19
1>
1C
b110 G
#241940000000
0!
0*
09
0>
0C
#241950000000
1!
1*
b111 6
19
1>
1C
b111 G
#241960000000
0!
0*
09
0>
0C
#241970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#241980000000
0!
0*
09
0>
0C
#241990000000
1!
1*
b1 6
19
1>
1C
b1 G
#242000000000
0!
0*
09
0>
0C
#242010000000
1!
1*
b10 6
19
1>
1C
b10 G
#242020000000
0!
0*
09
0>
0C
#242030000000
1!
1*
b11 6
19
1>
1C
b11 G
#242040000000
0!
0*
09
0>
0C
#242050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#242060000000
0!
0*
09
0>
0C
#242070000000
1!
1*
b101 6
19
1>
1C
b101 G
#242080000000
0!
0*
09
0>
0C
#242090000000
1!
1*
b110 6
19
1>
1C
b110 G
#242100000000
0!
0*
09
0>
0C
#242110000000
1!
1*
b111 6
19
1>
1C
b111 G
#242120000000
0!
1"
0*
1+
09
1:
0>
0C
#242130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#242140000000
0!
0*
09
0>
0C
#242150000000
1!
1*
b1 6
19
1>
1C
b1 G
#242160000000
0!
0*
09
0>
0C
#242170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#242180000000
0!
0*
09
0>
0C
#242190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#242200000000
0!
0*
09
0>
0C
#242210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#242220000000
0!
0*
09
0>
0C
#242230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#242240000000
0!
0#
0*
0,
09
0>
0?
0C
#242250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#242260000000
0!
0*
09
0>
0C
#242270000000
1!
1*
19
1>
1C
#242280000000
0!
0*
09
0>
0C
#242290000000
1!
1*
19
1>
1C
#242300000000
0!
0*
09
0>
0C
#242310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#242320000000
0!
0*
09
0>
0C
#242330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#242340000000
0!
0*
09
0>
0C
#242350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#242360000000
0!
0*
09
0>
0C
#242370000000
1!
1*
b10 6
19
1>
1C
b10 G
#242380000000
0!
0*
09
0>
0C
#242390000000
1!
1*
b11 6
19
1>
1C
b11 G
#242400000000
0!
0*
09
0>
0C
#242410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#242420000000
0!
0*
09
0>
0C
#242430000000
1!
1*
b101 6
19
1>
1C
b101 G
#242440000000
0!
0*
09
0>
0C
#242450000000
1!
1*
b110 6
19
1>
1C
b110 G
#242460000000
0!
0*
09
0>
0C
#242470000000
1!
1*
b111 6
19
1>
1C
b111 G
#242480000000
0!
0*
09
0>
0C
#242490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#242500000000
0!
0*
09
0>
0C
#242510000000
1!
1*
b1 6
19
1>
1C
b1 G
#242520000000
0!
0*
09
0>
0C
#242530000000
1!
1*
b10 6
19
1>
1C
b10 G
#242540000000
0!
0*
09
0>
0C
#242550000000
1!
1*
b11 6
19
1>
1C
b11 G
#242560000000
0!
0*
09
0>
0C
#242570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#242580000000
0!
0*
09
0>
0C
#242590000000
1!
1*
b101 6
19
1>
1C
b101 G
#242600000000
0!
0*
09
0>
0C
#242610000000
1!
1*
b110 6
19
1>
1C
b110 G
#242620000000
0!
0*
09
0>
0C
#242630000000
1!
1*
b111 6
19
1>
1C
b111 G
#242640000000
0!
0*
09
0>
0C
#242650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#242660000000
0!
0*
09
0>
0C
#242670000000
1!
1*
b1 6
19
1>
1C
b1 G
#242680000000
0!
0*
09
0>
0C
#242690000000
1!
1*
b10 6
19
1>
1C
b10 G
#242700000000
0!
0*
09
0>
0C
#242710000000
1!
1*
b11 6
19
1>
1C
b11 G
#242720000000
0!
0*
09
0>
0C
#242730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#242740000000
0!
0*
09
0>
0C
#242750000000
1!
1*
b101 6
19
1>
1C
b101 G
#242760000000
0!
0*
09
0>
0C
#242770000000
1!
1*
b110 6
19
1>
1C
b110 G
#242780000000
0!
0*
09
0>
0C
#242790000000
1!
1*
b111 6
19
1>
1C
b111 G
#242800000000
0!
1"
0*
1+
09
1:
0>
0C
#242810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#242820000000
0!
0*
09
0>
0C
#242830000000
1!
1*
b1 6
19
1>
1C
b1 G
#242840000000
0!
0*
09
0>
0C
#242850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#242860000000
0!
0*
09
0>
0C
#242870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#242880000000
0!
0*
09
0>
0C
#242890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#242900000000
0!
0*
09
0>
0C
#242910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#242920000000
0!
0#
0*
0,
09
0>
0?
0C
#242930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#242940000000
0!
0*
09
0>
0C
#242950000000
1!
1*
19
1>
1C
#242960000000
0!
0*
09
0>
0C
#242970000000
1!
1*
19
1>
1C
#242980000000
0!
0*
09
0>
0C
#242990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#243000000000
0!
0*
09
0>
0C
#243010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#243020000000
0!
0*
09
0>
0C
#243030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#243040000000
0!
0*
09
0>
0C
#243050000000
1!
1*
b10 6
19
1>
1C
b10 G
#243060000000
0!
0*
09
0>
0C
#243070000000
1!
1*
b11 6
19
1>
1C
b11 G
#243080000000
0!
0*
09
0>
0C
#243090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#243100000000
0!
0*
09
0>
0C
#243110000000
1!
1*
b101 6
19
1>
1C
b101 G
#243120000000
0!
0*
09
0>
0C
#243130000000
1!
1*
b110 6
19
1>
1C
b110 G
#243140000000
0!
0*
09
0>
0C
#243150000000
1!
1*
b111 6
19
1>
1C
b111 G
#243160000000
0!
0*
09
0>
0C
#243170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#243180000000
0!
0*
09
0>
0C
#243190000000
1!
1*
b1 6
19
1>
1C
b1 G
#243200000000
0!
0*
09
0>
0C
#243210000000
1!
1*
b10 6
19
1>
1C
b10 G
#243220000000
0!
0*
09
0>
0C
#243230000000
1!
1*
b11 6
19
1>
1C
b11 G
#243240000000
0!
0*
09
0>
0C
#243250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#243260000000
0!
0*
09
0>
0C
#243270000000
1!
1*
b101 6
19
1>
1C
b101 G
#243280000000
0!
0*
09
0>
0C
#243290000000
1!
1*
b110 6
19
1>
1C
b110 G
#243300000000
0!
0*
09
0>
0C
#243310000000
1!
1*
b111 6
19
1>
1C
b111 G
#243320000000
0!
0*
09
0>
0C
#243330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#243340000000
0!
0*
09
0>
0C
#243350000000
1!
1*
b1 6
19
1>
1C
b1 G
#243360000000
0!
0*
09
0>
0C
#243370000000
1!
1*
b10 6
19
1>
1C
b10 G
#243380000000
0!
0*
09
0>
0C
#243390000000
1!
1*
b11 6
19
1>
1C
b11 G
#243400000000
0!
0*
09
0>
0C
#243410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#243420000000
0!
0*
09
0>
0C
#243430000000
1!
1*
b101 6
19
1>
1C
b101 G
#243440000000
0!
0*
09
0>
0C
#243450000000
1!
1*
b110 6
19
1>
1C
b110 G
#243460000000
0!
0*
09
0>
0C
#243470000000
1!
1*
b111 6
19
1>
1C
b111 G
#243480000000
0!
1"
0*
1+
09
1:
0>
0C
#243490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#243500000000
0!
0*
09
0>
0C
#243510000000
1!
1*
b1 6
19
1>
1C
b1 G
#243520000000
0!
0*
09
0>
0C
#243530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#243540000000
0!
0*
09
0>
0C
#243550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#243560000000
0!
0*
09
0>
0C
#243570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#243580000000
0!
0*
09
0>
0C
#243590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#243600000000
0!
0#
0*
0,
09
0>
0?
0C
#243610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#243620000000
0!
0*
09
0>
0C
#243630000000
1!
1*
19
1>
1C
#243640000000
0!
0*
09
0>
0C
#243650000000
1!
1*
19
1>
1C
#243660000000
0!
0*
09
0>
0C
#243670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#243680000000
0!
0*
09
0>
0C
#243690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#243700000000
0!
0*
09
0>
0C
#243710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#243720000000
0!
0*
09
0>
0C
#243730000000
1!
1*
b10 6
19
1>
1C
b10 G
#243740000000
0!
0*
09
0>
0C
#243750000000
1!
1*
b11 6
19
1>
1C
b11 G
#243760000000
0!
0*
09
0>
0C
#243770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#243780000000
0!
0*
09
0>
0C
#243790000000
1!
1*
b101 6
19
1>
1C
b101 G
#243800000000
0!
0*
09
0>
0C
#243810000000
1!
1*
b110 6
19
1>
1C
b110 G
#243820000000
0!
0*
09
0>
0C
#243830000000
1!
1*
b111 6
19
1>
1C
b111 G
#243840000000
0!
0*
09
0>
0C
#243850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#243860000000
0!
0*
09
0>
0C
#243870000000
1!
1*
b1 6
19
1>
1C
b1 G
#243880000000
0!
0*
09
0>
0C
#243890000000
1!
1*
b10 6
19
1>
1C
b10 G
#243900000000
0!
0*
09
0>
0C
#243910000000
1!
1*
b11 6
19
1>
1C
b11 G
#243920000000
0!
0*
09
0>
0C
#243930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#243940000000
0!
0*
09
0>
0C
#243950000000
1!
1*
b101 6
19
1>
1C
b101 G
#243960000000
0!
0*
09
0>
0C
#243970000000
1!
1*
b110 6
19
1>
1C
b110 G
#243980000000
0!
0*
09
0>
0C
#243990000000
1!
1*
b111 6
19
1>
1C
b111 G
#244000000000
0!
0*
09
0>
0C
#244010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#244020000000
0!
0*
09
0>
0C
#244030000000
1!
1*
b1 6
19
1>
1C
b1 G
#244040000000
0!
0*
09
0>
0C
#244050000000
1!
1*
b10 6
19
1>
1C
b10 G
#244060000000
0!
0*
09
0>
0C
#244070000000
1!
1*
b11 6
19
1>
1C
b11 G
#244080000000
0!
0*
09
0>
0C
#244090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#244100000000
0!
0*
09
0>
0C
#244110000000
1!
1*
b101 6
19
1>
1C
b101 G
#244120000000
0!
0*
09
0>
0C
#244130000000
1!
1*
b110 6
19
1>
1C
b110 G
#244140000000
0!
0*
09
0>
0C
#244150000000
1!
1*
b111 6
19
1>
1C
b111 G
#244160000000
0!
1"
0*
1+
09
1:
0>
0C
#244170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#244180000000
0!
0*
09
0>
0C
#244190000000
1!
1*
b1 6
19
1>
1C
b1 G
#244200000000
0!
0*
09
0>
0C
#244210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#244220000000
0!
0*
09
0>
0C
#244230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#244240000000
0!
0*
09
0>
0C
#244250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#244260000000
0!
0*
09
0>
0C
#244270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#244280000000
0!
0#
0*
0,
09
0>
0?
0C
#244290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#244300000000
0!
0*
09
0>
0C
#244310000000
1!
1*
19
1>
1C
#244320000000
0!
0*
09
0>
0C
#244330000000
1!
1*
19
1>
1C
#244340000000
0!
0*
09
0>
0C
#244350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#244360000000
0!
0*
09
0>
0C
#244370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#244380000000
0!
0*
09
0>
0C
#244390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#244400000000
0!
0*
09
0>
0C
#244410000000
1!
1*
b10 6
19
1>
1C
b10 G
#244420000000
0!
0*
09
0>
0C
#244430000000
1!
1*
b11 6
19
1>
1C
b11 G
#244440000000
0!
0*
09
0>
0C
#244450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#244460000000
0!
0*
09
0>
0C
#244470000000
1!
1*
b101 6
19
1>
1C
b101 G
#244480000000
0!
0*
09
0>
0C
#244490000000
1!
1*
b110 6
19
1>
1C
b110 G
#244500000000
0!
0*
09
0>
0C
#244510000000
1!
1*
b111 6
19
1>
1C
b111 G
#244520000000
0!
0*
09
0>
0C
#244530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#244540000000
0!
0*
09
0>
0C
#244550000000
1!
1*
b1 6
19
1>
1C
b1 G
#244560000000
0!
0*
09
0>
0C
#244570000000
1!
1*
b10 6
19
1>
1C
b10 G
#244580000000
0!
0*
09
0>
0C
#244590000000
1!
1*
b11 6
19
1>
1C
b11 G
#244600000000
0!
0*
09
0>
0C
#244610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#244620000000
0!
0*
09
0>
0C
#244630000000
1!
1*
b101 6
19
1>
1C
b101 G
#244640000000
0!
0*
09
0>
0C
#244650000000
1!
1*
b110 6
19
1>
1C
b110 G
#244660000000
0!
0*
09
0>
0C
#244670000000
1!
1*
b111 6
19
1>
1C
b111 G
#244680000000
0!
0*
09
0>
0C
#244690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#244700000000
0!
0*
09
0>
0C
#244710000000
1!
1*
b1 6
19
1>
1C
b1 G
#244720000000
0!
0*
09
0>
0C
#244730000000
1!
1*
b10 6
19
1>
1C
b10 G
#244740000000
0!
0*
09
0>
0C
#244750000000
1!
1*
b11 6
19
1>
1C
b11 G
#244760000000
0!
0*
09
0>
0C
#244770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#244780000000
0!
0*
09
0>
0C
#244790000000
1!
1*
b101 6
19
1>
1C
b101 G
#244800000000
0!
0*
09
0>
0C
#244810000000
1!
1*
b110 6
19
1>
1C
b110 G
#244820000000
0!
0*
09
0>
0C
#244830000000
1!
1*
b111 6
19
1>
1C
b111 G
#244840000000
0!
1"
0*
1+
09
1:
0>
0C
#244850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#244860000000
0!
0*
09
0>
0C
#244870000000
1!
1*
b1 6
19
1>
1C
b1 G
#244880000000
0!
0*
09
0>
0C
#244890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#244900000000
0!
0*
09
0>
0C
#244910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#244920000000
0!
0*
09
0>
0C
#244930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#244940000000
0!
0*
09
0>
0C
#244950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#244960000000
0!
0#
0*
0,
09
0>
0?
0C
#244970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#244980000000
0!
0*
09
0>
0C
#244990000000
1!
1*
19
1>
1C
#245000000000
0!
0*
09
0>
0C
#245010000000
1!
1*
19
1>
1C
#245020000000
0!
0*
09
0>
0C
#245030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#245040000000
0!
0*
09
0>
0C
#245050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#245060000000
0!
0*
09
0>
0C
#245070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#245080000000
0!
0*
09
0>
0C
#245090000000
1!
1*
b10 6
19
1>
1C
b10 G
#245100000000
0!
0*
09
0>
0C
#245110000000
1!
1*
b11 6
19
1>
1C
b11 G
#245120000000
0!
0*
09
0>
0C
#245130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#245140000000
0!
0*
09
0>
0C
#245150000000
1!
1*
b101 6
19
1>
1C
b101 G
#245160000000
0!
0*
09
0>
0C
#245170000000
1!
1*
b110 6
19
1>
1C
b110 G
#245180000000
0!
0*
09
0>
0C
#245190000000
1!
1*
b111 6
19
1>
1C
b111 G
#245200000000
0!
0*
09
0>
0C
#245210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#245220000000
0!
0*
09
0>
0C
#245230000000
1!
1*
b1 6
19
1>
1C
b1 G
#245240000000
0!
0*
09
0>
0C
#245250000000
1!
1*
b10 6
19
1>
1C
b10 G
#245260000000
0!
0*
09
0>
0C
#245270000000
1!
1*
b11 6
19
1>
1C
b11 G
#245280000000
0!
0*
09
0>
0C
#245290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#245300000000
0!
0*
09
0>
0C
#245310000000
1!
1*
b101 6
19
1>
1C
b101 G
#245320000000
0!
0*
09
0>
0C
#245330000000
1!
1*
b110 6
19
1>
1C
b110 G
#245340000000
0!
0*
09
0>
0C
#245350000000
1!
1*
b111 6
19
1>
1C
b111 G
#245360000000
0!
0*
09
0>
0C
#245370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#245380000000
0!
0*
09
0>
0C
#245390000000
1!
1*
b1 6
19
1>
1C
b1 G
#245400000000
0!
0*
09
0>
0C
#245410000000
1!
1*
b10 6
19
1>
1C
b10 G
#245420000000
0!
0*
09
0>
0C
#245430000000
1!
1*
b11 6
19
1>
1C
b11 G
#245440000000
0!
0*
09
0>
0C
#245450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#245460000000
0!
0*
09
0>
0C
#245470000000
1!
1*
b101 6
19
1>
1C
b101 G
#245480000000
0!
0*
09
0>
0C
#245490000000
1!
1*
b110 6
19
1>
1C
b110 G
#245500000000
0!
0*
09
0>
0C
#245510000000
1!
1*
b111 6
19
1>
1C
b111 G
#245520000000
0!
1"
0*
1+
09
1:
0>
0C
#245530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#245540000000
0!
0*
09
0>
0C
#245550000000
1!
1*
b1 6
19
1>
1C
b1 G
#245560000000
0!
0*
09
0>
0C
#245570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#245580000000
0!
0*
09
0>
0C
#245590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#245600000000
0!
0*
09
0>
0C
#245610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#245620000000
0!
0*
09
0>
0C
#245630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#245640000000
0!
0#
0*
0,
09
0>
0?
0C
#245650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#245660000000
0!
0*
09
0>
0C
#245670000000
1!
1*
19
1>
1C
#245680000000
0!
0*
09
0>
0C
#245690000000
1!
1*
19
1>
1C
#245700000000
0!
0*
09
0>
0C
#245710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#245720000000
0!
0*
09
0>
0C
#245730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#245740000000
0!
0*
09
0>
0C
#245750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#245760000000
0!
0*
09
0>
0C
#245770000000
1!
1*
b10 6
19
1>
1C
b10 G
#245780000000
0!
0*
09
0>
0C
#245790000000
1!
1*
b11 6
19
1>
1C
b11 G
#245800000000
0!
0*
09
0>
0C
#245810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#245820000000
0!
0*
09
0>
0C
#245830000000
1!
1*
b101 6
19
1>
1C
b101 G
#245840000000
0!
0*
09
0>
0C
#245850000000
1!
1*
b110 6
19
1>
1C
b110 G
#245860000000
0!
0*
09
0>
0C
#245870000000
1!
1*
b111 6
19
1>
1C
b111 G
#245880000000
0!
0*
09
0>
0C
#245890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#245900000000
0!
0*
09
0>
0C
#245910000000
1!
1*
b1 6
19
1>
1C
b1 G
#245920000000
0!
0*
09
0>
0C
#245930000000
1!
1*
b10 6
19
1>
1C
b10 G
#245940000000
0!
0*
09
0>
0C
#245950000000
1!
1*
b11 6
19
1>
1C
b11 G
#245960000000
0!
0*
09
0>
0C
#245970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#245980000000
0!
0*
09
0>
0C
#245990000000
1!
1*
b101 6
19
1>
1C
b101 G
#246000000000
0!
0*
09
0>
0C
#246010000000
1!
1*
b110 6
19
1>
1C
b110 G
#246020000000
0!
0*
09
0>
0C
#246030000000
1!
1*
b111 6
19
1>
1C
b111 G
#246040000000
0!
0*
09
0>
0C
#246050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#246060000000
0!
0*
09
0>
0C
#246070000000
1!
1*
b1 6
19
1>
1C
b1 G
#246080000000
0!
0*
09
0>
0C
#246090000000
1!
1*
b10 6
19
1>
1C
b10 G
#246100000000
0!
0*
09
0>
0C
#246110000000
1!
1*
b11 6
19
1>
1C
b11 G
#246120000000
0!
0*
09
0>
0C
#246130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#246140000000
0!
0*
09
0>
0C
#246150000000
1!
1*
b101 6
19
1>
1C
b101 G
#246160000000
0!
0*
09
0>
0C
#246170000000
1!
1*
b110 6
19
1>
1C
b110 G
#246180000000
0!
0*
09
0>
0C
#246190000000
1!
1*
b111 6
19
1>
1C
b111 G
#246200000000
0!
1"
0*
1+
09
1:
0>
0C
#246210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#246220000000
0!
0*
09
0>
0C
#246230000000
1!
1*
b1 6
19
1>
1C
b1 G
#246240000000
0!
0*
09
0>
0C
#246250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#246260000000
0!
0*
09
0>
0C
#246270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#246280000000
0!
0*
09
0>
0C
#246290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#246300000000
0!
0*
09
0>
0C
#246310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#246320000000
0!
0#
0*
0,
09
0>
0?
0C
#246330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#246340000000
0!
0*
09
0>
0C
#246350000000
1!
1*
19
1>
1C
#246360000000
0!
0*
09
0>
0C
#246370000000
1!
1*
19
1>
1C
#246380000000
0!
0*
09
0>
0C
#246390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#246400000000
0!
0*
09
0>
0C
#246410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#246420000000
0!
0*
09
0>
0C
#246430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#246440000000
0!
0*
09
0>
0C
#246450000000
1!
1*
b10 6
19
1>
1C
b10 G
#246460000000
0!
0*
09
0>
0C
#246470000000
1!
1*
b11 6
19
1>
1C
b11 G
#246480000000
0!
0*
09
0>
0C
#246490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#246500000000
0!
0*
09
0>
0C
#246510000000
1!
1*
b101 6
19
1>
1C
b101 G
#246520000000
0!
0*
09
0>
0C
#246530000000
1!
1*
b110 6
19
1>
1C
b110 G
#246540000000
0!
0*
09
0>
0C
#246550000000
1!
1*
b111 6
19
1>
1C
b111 G
#246560000000
0!
0*
09
0>
0C
#246570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#246580000000
0!
0*
09
0>
0C
#246590000000
1!
1*
b1 6
19
1>
1C
b1 G
#246600000000
0!
0*
09
0>
0C
#246610000000
1!
1*
b10 6
19
1>
1C
b10 G
#246620000000
0!
0*
09
0>
0C
#246630000000
1!
1*
b11 6
19
1>
1C
b11 G
#246640000000
0!
0*
09
0>
0C
#246650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#246660000000
0!
0*
09
0>
0C
#246670000000
1!
1*
b101 6
19
1>
1C
b101 G
#246680000000
0!
0*
09
0>
0C
#246690000000
1!
1*
b110 6
19
1>
1C
b110 G
#246700000000
0!
0*
09
0>
0C
#246710000000
1!
1*
b111 6
19
1>
1C
b111 G
#246720000000
0!
0*
09
0>
0C
#246730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#246740000000
0!
0*
09
0>
0C
#246750000000
1!
1*
b1 6
19
1>
1C
b1 G
#246760000000
0!
0*
09
0>
0C
#246770000000
1!
1*
b10 6
19
1>
1C
b10 G
#246780000000
0!
0*
09
0>
0C
#246790000000
1!
1*
b11 6
19
1>
1C
b11 G
#246800000000
0!
0*
09
0>
0C
#246810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#246820000000
0!
0*
09
0>
0C
#246830000000
1!
1*
b101 6
19
1>
1C
b101 G
#246840000000
0!
0*
09
0>
0C
#246850000000
1!
1*
b110 6
19
1>
1C
b110 G
#246860000000
0!
0*
09
0>
0C
#246870000000
1!
1*
b111 6
19
1>
1C
b111 G
#246880000000
0!
1"
0*
1+
09
1:
0>
0C
#246890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#246900000000
0!
0*
09
0>
0C
#246910000000
1!
1*
b1 6
19
1>
1C
b1 G
#246920000000
0!
0*
09
0>
0C
#246930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#246940000000
0!
0*
09
0>
0C
#246950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#246960000000
0!
0*
09
0>
0C
#246970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#246980000000
0!
0*
09
0>
0C
#246990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#247000000000
0!
0#
0*
0,
09
0>
0?
0C
#247010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#247020000000
0!
0*
09
0>
0C
#247030000000
1!
1*
19
1>
1C
#247040000000
0!
0*
09
0>
0C
#247050000000
1!
1*
19
1>
1C
#247060000000
0!
0*
09
0>
0C
#247070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#247080000000
0!
0*
09
0>
0C
#247090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#247100000000
0!
0*
09
0>
0C
#247110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#247120000000
0!
0*
09
0>
0C
#247130000000
1!
1*
b10 6
19
1>
1C
b10 G
#247140000000
0!
0*
09
0>
0C
#247150000000
1!
1*
b11 6
19
1>
1C
b11 G
#247160000000
0!
0*
09
0>
0C
#247170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#247180000000
0!
0*
09
0>
0C
#247190000000
1!
1*
b101 6
19
1>
1C
b101 G
#247200000000
0!
0*
09
0>
0C
#247210000000
1!
1*
b110 6
19
1>
1C
b110 G
#247220000000
0!
0*
09
0>
0C
#247230000000
1!
1*
b111 6
19
1>
1C
b111 G
#247240000000
0!
0*
09
0>
0C
#247250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#247260000000
0!
0*
09
0>
0C
#247270000000
1!
1*
b1 6
19
1>
1C
b1 G
#247280000000
0!
0*
09
0>
0C
#247290000000
1!
1*
b10 6
19
1>
1C
b10 G
#247300000000
0!
0*
09
0>
0C
#247310000000
1!
1*
b11 6
19
1>
1C
b11 G
#247320000000
0!
0*
09
0>
0C
#247330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#247340000000
0!
0*
09
0>
0C
#247350000000
1!
1*
b101 6
19
1>
1C
b101 G
#247360000000
0!
0*
09
0>
0C
#247370000000
1!
1*
b110 6
19
1>
1C
b110 G
#247380000000
0!
0*
09
0>
0C
#247390000000
1!
1*
b111 6
19
1>
1C
b111 G
#247400000000
0!
0*
09
0>
0C
#247410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#247420000000
0!
0*
09
0>
0C
#247430000000
1!
1*
b1 6
19
1>
1C
b1 G
#247440000000
0!
0*
09
0>
0C
#247450000000
1!
1*
b10 6
19
1>
1C
b10 G
#247460000000
0!
0*
09
0>
0C
#247470000000
1!
1*
b11 6
19
1>
1C
b11 G
#247480000000
0!
0*
09
0>
0C
#247490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#247500000000
0!
0*
09
0>
0C
#247510000000
1!
1*
b101 6
19
1>
1C
b101 G
#247520000000
0!
0*
09
0>
0C
#247530000000
1!
1*
b110 6
19
1>
1C
b110 G
#247540000000
0!
0*
09
0>
0C
#247550000000
1!
1*
b111 6
19
1>
1C
b111 G
#247560000000
0!
1"
0*
1+
09
1:
0>
0C
#247570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#247580000000
0!
0*
09
0>
0C
#247590000000
1!
1*
b1 6
19
1>
1C
b1 G
#247600000000
0!
0*
09
0>
0C
#247610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#247620000000
0!
0*
09
0>
0C
#247630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#247640000000
0!
0*
09
0>
0C
#247650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#247660000000
0!
0*
09
0>
0C
#247670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#247680000000
0!
0#
0*
0,
09
0>
0?
0C
#247690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#247700000000
0!
0*
09
0>
0C
#247710000000
1!
1*
19
1>
1C
#247720000000
0!
0*
09
0>
0C
#247730000000
1!
1*
19
1>
1C
#247740000000
0!
0*
09
0>
0C
#247750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#247760000000
0!
0*
09
0>
0C
#247770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#247780000000
0!
0*
09
0>
0C
#247790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#247800000000
0!
0*
09
0>
0C
#247810000000
1!
1*
b10 6
19
1>
1C
b10 G
#247820000000
0!
0*
09
0>
0C
#247830000000
1!
1*
b11 6
19
1>
1C
b11 G
#247840000000
0!
0*
09
0>
0C
#247850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#247860000000
0!
0*
09
0>
0C
#247870000000
1!
1*
b101 6
19
1>
1C
b101 G
#247880000000
0!
0*
09
0>
0C
#247890000000
1!
1*
b110 6
19
1>
1C
b110 G
#247900000000
0!
0*
09
0>
0C
#247910000000
1!
1*
b111 6
19
1>
1C
b111 G
#247920000000
0!
0*
09
0>
0C
#247930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#247940000000
0!
0*
09
0>
0C
#247950000000
1!
1*
b1 6
19
1>
1C
b1 G
#247960000000
0!
0*
09
0>
0C
#247970000000
1!
1*
b10 6
19
1>
1C
b10 G
#247980000000
0!
0*
09
0>
0C
#247990000000
1!
1*
b11 6
19
1>
1C
b11 G
#248000000000
0!
0*
09
0>
0C
#248010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#248020000000
0!
0*
09
0>
0C
#248030000000
1!
1*
b101 6
19
1>
1C
b101 G
#248040000000
0!
0*
09
0>
0C
#248050000000
1!
1*
b110 6
19
1>
1C
b110 G
#248060000000
0!
0*
09
0>
0C
#248070000000
1!
1*
b111 6
19
1>
1C
b111 G
#248080000000
0!
0*
09
0>
0C
#248090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#248100000000
0!
0*
09
0>
0C
#248110000000
1!
1*
b1 6
19
1>
1C
b1 G
#248120000000
0!
0*
09
0>
0C
#248130000000
1!
1*
b10 6
19
1>
1C
b10 G
#248140000000
0!
0*
09
0>
0C
#248150000000
1!
1*
b11 6
19
1>
1C
b11 G
#248160000000
0!
0*
09
0>
0C
#248170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#248180000000
0!
0*
09
0>
0C
#248190000000
1!
1*
b101 6
19
1>
1C
b101 G
#248200000000
0!
0*
09
0>
0C
#248210000000
1!
1*
b110 6
19
1>
1C
b110 G
#248220000000
0!
0*
09
0>
0C
#248230000000
1!
1*
b111 6
19
1>
1C
b111 G
#248240000000
0!
1"
0*
1+
09
1:
0>
0C
#248250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#248260000000
0!
0*
09
0>
0C
#248270000000
1!
1*
b1 6
19
1>
1C
b1 G
#248280000000
0!
0*
09
0>
0C
#248290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#248300000000
0!
0*
09
0>
0C
#248310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#248320000000
0!
0*
09
0>
0C
#248330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#248340000000
0!
0*
09
0>
0C
#248350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#248360000000
0!
0#
0*
0,
09
0>
0?
0C
#248370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#248380000000
0!
0*
09
0>
0C
#248390000000
1!
1*
19
1>
1C
#248400000000
0!
0*
09
0>
0C
#248410000000
1!
1*
19
1>
1C
#248420000000
0!
0*
09
0>
0C
#248430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#248440000000
0!
0*
09
0>
0C
#248450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#248460000000
0!
0*
09
0>
0C
#248470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#248480000000
0!
0*
09
0>
0C
#248490000000
1!
1*
b10 6
19
1>
1C
b10 G
#248500000000
0!
0*
09
0>
0C
#248510000000
1!
1*
b11 6
19
1>
1C
b11 G
#248520000000
0!
0*
09
0>
0C
#248530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#248540000000
0!
0*
09
0>
0C
#248550000000
1!
1*
b101 6
19
1>
1C
b101 G
#248560000000
0!
0*
09
0>
0C
#248570000000
1!
1*
b110 6
19
1>
1C
b110 G
#248580000000
0!
0*
09
0>
0C
#248590000000
1!
1*
b111 6
19
1>
1C
b111 G
#248600000000
0!
0*
09
0>
0C
#248610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#248620000000
0!
0*
09
0>
0C
#248630000000
1!
1*
b1 6
19
1>
1C
b1 G
#248640000000
0!
0*
09
0>
0C
#248650000000
1!
1*
b10 6
19
1>
1C
b10 G
#248660000000
0!
0*
09
0>
0C
#248670000000
1!
1*
b11 6
19
1>
1C
b11 G
#248680000000
0!
0*
09
0>
0C
#248690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#248700000000
0!
0*
09
0>
0C
#248710000000
1!
1*
b101 6
19
1>
1C
b101 G
#248720000000
0!
0*
09
0>
0C
#248730000000
1!
1*
b110 6
19
1>
1C
b110 G
#248740000000
0!
0*
09
0>
0C
#248750000000
1!
1*
b111 6
19
1>
1C
b111 G
#248760000000
0!
0*
09
0>
0C
#248770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#248780000000
0!
0*
09
0>
0C
#248790000000
1!
1*
b1 6
19
1>
1C
b1 G
#248800000000
0!
0*
09
0>
0C
#248810000000
1!
1*
b10 6
19
1>
1C
b10 G
#248820000000
0!
0*
09
0>
0C
#248830000000
1!
1*
b11 6
19
1>
1C
b11 G
#248840000000
0!
0*
09
0>
0C
#248850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#248860000000
0!
0*
09
0>
0C
#248870000000
1!
1*
b101 6
19
1>
1C
b101 G
#248880000000
0!
0*
09
0>
0C
#248890000000
1!
1*
b110 6
19
1>
1C
b110 G
#248900000000
0!
0*
09
0>
0C
#248910000000
1!
1*
b111 6
19
1>
1C
b111 G
#248920000000
0!
1"
0*
1+
09
1:
0>
0C
#248930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#248940000000
0!
0*
09
0>
0C
#248950000000
1!
1*
b1 6
19
1>
1C
b1 G
#248960000000
0!
0*
09
0>
0C
#248970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#248980000000
0!
0*
09
0>
0C
#248990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#249000000000
0!
0*
09
0>
0C
#249010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#249020000000
0!
0*
09
0>
0C
#249030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#249040000000
0!
0#
0*
0,
09
0>
0?
0C
#249050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#249060000000
0!
0*
09
0>
0C
#249070000000
1!
1*
19
1>
1C
#249080000000
0!
0*
09
0>
0C
#249090000000
1!
1*
19
1>
1C
#249100000000
0!
0*
09
0>
0C
#249110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#249120000000
0!
0*
09
0>
0C
#249130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#249140000000
0!
0*
09
0>
0C
#249150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#249160000000
0!
0*
09
0>
0C
#249170000000
1!
1*
b10 6
19
1>
1C
b10 G
#249180000000
0!
0*
09
0>
0C
#249190000000
1!
1*
b11 6
19
1>
1C
b11 G
#249200000000
0!
0*
09
0>
0C
#249210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#249220000000
0!
0*
09
0>
0C
#249230000000
1!
1*
b101 6
19
1>
1C
b101 G
#249240000000
0!
0*
09
0>
0C
#249250000000
1!
1*
b110 6
19
1>
1C
b110 G
#249260000000
0!
0*
09
0>
0C
#249270000000
1!
1*
b111 6
19
1>
1C
b111 G
#249280000000
0!
0*
09
0>
0C
#249290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#249300000000
0!
0*
09
0>
0C
#249310000000
1!
1*
b1 6
19
1>
1C
b1 G
#249320000000
0!
0*
09
0>
0C
#249330000000
1!
1*
b10 6
19
1>
1C
b10 G
#249340000000
0!
0*
09
0>
0C
#249350000000
1!
1*
b11 6
19
1>
1C
b11 G
#249360000000
0!
0*
09
0>
0C
#249370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#249380000000
0!
0*
09
0>
0C
#249390000000
1!
1*
b101 6
19
1>
1C
b101 G
#249400000000
0!
0*
09
0>
0C
#249410000000
1!
1*
b110 6
19
1>
1C
b110 G
#249420000000
0!
0*
09
0>
0C
#249430000000
1!
1*
b111 6
19
1>
1C
b111 G
#249440000000
0!
0*
09
0>
0C
#249450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#249460000000
0!
0*
09
0>
0C
#249470000000
1!
1*
b1 6
19
1>
1C
b1 G
#249480000000
0!
0*
09
0>
0C
#249490000000
1!
1*
b10 6
19
1>
1C
b10 G
#249500000000
0!
0*
09
0>
0C
#249510000000
1!
1*
b11 6
19
1>
1C
b11 G
#249520000000
0!
0*
09
0>
0C
#249530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#249540000000
0!
0*
09
0>
0C
#249550000000
1!
1*
b101 6
19
1>
1C
b101 G
#249560000000
0!
0*
09
0>
0C
#249570000000
1!
1*
b110 6
19
1>
1C
b110 G
#249580000000
0!
0*
09
0>
0C
#249590000000
1!
1*
b111 6
19
1>
1C
b111 G
#249600000000
0!
1"
0*
1+
09
1:
0>
0C
#249610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#249620000000
0!
0*
09
0>
0C
#249630000000
1!
1*
b1 6
19
1>
1C
b1 G
#249640000000
0!
0*
09
0>
0C
#249650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#249660000000
0!
0*
09
0>
0C
#249670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#249680000000
0!
0*
09
0>
0C
#249690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#249700000000
0!
0*
09
0>
0C
#249710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#249720000000
0!
0#
0*
0,
09
0>
0?
0C
#249730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#249740000000
0!
0*
09
0>
0C
#249750000000
1!
1*
19
1>
1C
#249760000000
0!
0*
09
0>
0C
#249770000000
1!
1*
19
1>
1C
#249780000000
0!
0*
09
0>
0C
#249790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#249800000000
0!
0*
09
0>
0C
#249810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#249820000000
0!
0*
09
0>
0C
#249830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#249840000000
0!
0*
09
0>
0C
#249850000000
1!
1*
b10 6
19
1>
1C
b10 G
#249860000000
0!
0*
09
0>
0C
#249870000000
1!
1*
b11 6
19
1>
1C
b11 G
#249880000000
0!
0*
09
0>
0C
#249890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#249900000000
0!
0*
09
0>
0C
#249910000000
1!
1*
b101 6
19
1>
1C
b101 G
#249920000000
0!
0*
09
0>
0C
#249930000000
1!
1*
b110 6
19
1>
1C
b110 G
#249940000000
0!
0*
09
0>
0C
#249950000000
1!
1*
b111 6
19
1>
1C
b111 G
#249960000000
0!
0*
09
0>
0C
#249970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#249980000000
0!
0*
09
0>
0C
#249990000000
1!
1*
b1 6
19
1>
1C
b1 G
#250000000000
0!
0*
09
0>
0C
#250010000000
1!
1*
b10 6
19
1>
1C
b10 G
#250020000000
0!
0*
09
0>
0C
#250030000000
1!
1*
b11 6
19
1>
1C
b11 G
#250040000000
0!
0*
09
0>
0C
#250050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#250060000000
0!
0*
09
0>
0C
#250070000000
1!
1*
b101 6
19
1>
1C
b101 G
#250080000000
0!
0*
09
0>
0C
#250090000000
1!
1*
b110 6
19
1>
1C
b110 G
#250100000000
0!
0*
09
0>
0C
#250110000000
1!
1*
b111 6
19
1>
1C
b111 G
#250120000000
0!
0*
09
0>
0C
#250130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#250140000000
0!
0*
09
0>
0C
#250150000000
1!
1*
b1 6
19
1>
1C
b1 G
#250160000000
0!
0*
09
0>
0C
#250170000000
1!
1*
b10 6
19
1>
1C
b10 G
#250180000000
0!
0*
09
0>
0C
#250190000000
1!
1*
b11 6
19
1>
1C
b11 G
#250200000000
0!
0*
09
0>
0C
#250210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#250220000000
0!
0*
09
0>
0C
#250230000000
1!
1*
b101 6
19
1>
1C
b101 G
#250240000000
0!
0*
09
0>
0C
#250250000000
1!
1*
b110 6
19
1>
1C
b110 G
#250260000000
0!
0*
09
0>
0C
#250270000000
1!
1*
b111 6
19
1>
1C
b111 G
#250280000000
0!
1"
0*
1+
09
1:
0>
0C
#250290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#250300000000
0!
0*
09
0>
0C
#250310000000
1!
1*
b1 6
19
1>
1C
b1 G
#250320000000
0!
0*
09
0>
0C
#250330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#250340000000
0!
0*
09
0>
0C
#250350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#250360000000
0!
0*
09
0>
0C
#250370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#250380000000
0!
0*
09
0>
0C
#250390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#250400000000
0!
0#
0*
0,
09
0>
0?
0C
#250410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#250420000000
0!
0*
09
0>
0C
#250430000000
1!
1*
19
1>
1C
#250440000000
0!
0*
09
0>
0C
#250450000000
1!
1*
19
1>
1C
#250460000000
0!
0*
09
0>
0C
#250470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#250480000000
0!
0*
09
0>
0C
#250490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#250500000000
0!
0*
09
0>
0C
#250510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#250520000000
0!
0*
09
0>
0C
#250530000000
1!
1*
b10 6
19
1>
1C
b10 G
#250540000000
0!
0*
09
0>
0C
#250550000000
1!
1*
b11 6
19
1>
1C
b11 G
#250560000000
0!
0*
09
0>
0C
#250570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#250580000000
0!
0*
09
0>
0C
#250590000000
1!
1*
b101 6
19
1>
1C
b101 G
#250600000000
0!
0*
09
0>
0C
#250610000000
1!
1*
b110 6
19
1>
1C
b110 G
#250620000000
0!
0*
09
0>
0C
#250630000000
1!
1*
b111 6
19
1>
1C
b111 G
#250640000000
0!
0*
09
0>
0C
#250650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#250660000000
0!
0*
09
0>
0C
#250670000000
1!
1*
b1 6
19
1>
1C
b1 G
#250680000000
0!
0*
09
0>
0C
#250690000000
1!
1*
b10 6
19
1>
1C
b10 G
#250700000000
0!
0*
09
0>
0C
#250710000000
1!
1*
b11 6
19
1>
1C
b11 G
#250720000000
0!
0*
09
0>
0C
#250730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#250740000000
0!
0*
09
0>
0C
#250750000000
1!
1*
b101 6
19
1>
1C
b101 G
#250760000000
0!
0*
09
0>
0C
#250770000000
1!
1*
b110 6
19
1>
1C
b110 G
#250780000000
0!
0*
09
0>
0C
#250790000000
1!
1*
b111 6
19
1>
1C
b111 G
#250800000000
0!
0*
09
0>
0C
#250810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#250820000000
0!
0*
09
0>
0C
#250830000000
1!
1*
b1 6
19
1>
1C
b1 G
#250840000000
0!
0*
09
0>
0C
#250850000000
1!
1*
b10 6
19
1>
1C
b10 G
#250860000000
0!
0*
09
0>
0C
#250870000000
1!
1*
b11 6
19
1>
1C
b11 G
#250880000000
0!
0*
09
0>
0C
#250890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#250900000000
0!
0*
09
0>
0C
#250910000000
1!
1*
b101 6
19
1>
1C
b101 G
#250920000000
0!
0*
09
0>
0C
#250930000000
1!
1*
b110 6
19
1>
1C
b110 G
#250940000000
0!
0*
09
0>
0C
#250950000000
1!
1*
b111 6
19
1>
1C
b111 G
#250960000000
0!
1"
0*
1+
09
1:
0>
0C
#250970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#250980000000
0!
0*
09
0>
0C
#250990000000
1!
1*
b1 6
19
1>
1C
b1 G
#251000000000
0!
0*
09
0>
0C
#251010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#251020000000
0!
0*
09
0>
0C
#251030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#251040000000
0!
0*
09
0>
0C
#251050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#251060000000
0!
0*
09
0>
0C
#251070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#251080000000
0!
0#
0*
0,
09
0>
0?
0C
#251090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#251100000000
0!
0*
09
0>
0C
#251110000000
1!
1*
19
1>
1C
#251120000000
0!
0*
09
0>
0C
#251130000000
1!
1*
19
1>
1C
#251140000000
0!
0*
09
0>
0C
#251150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#251160000000
0!
0*
09
0>
0C
#251170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#251180000000
0!
0*
09
0>
0C
#251190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#251200000000
0!
0*
09
0>
0C
#251210000000
1!
1*
b10 6
19
1>
1C
b10 G
#251220000000
0!
0*
09
0>
0C
#251230000000
1!
1*
b11 6
19
1>
1C
b11 G
#251240000000
0!
0*
09
0>
0C
#251250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#251260000000
0!
0*
09
0>
0C
#251270000000
1!
1*
b101 6
19
1>
1C
b101 G
#251280000000
0!
0*
09
0>
0C
#251290000000
1!
1*
b110 6
19
1>
1C
b110 G
#251300000000
0!
0*
09
0>
0C
#251310000000
1!
1*
b111 6
19
1>
1C
b111 G
#251320000000
0!
0*
09
0>
0C
#251330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#251340000000
0!
0*
09
0>
0C
#251350000000
1!
1*
b1 6
19
1>
1C
b1 G
#251360000000
0!
0*
09
0>
0C
#251370000000
1!
1*
b10 6
19
1>
1C
b10 G
#251380000000
0!
0*
09
0>
0C
#251390000000
1!
1*
b11 6
19
1>
1C
b11 G
#251400000000
0!
0*
09
0>
0C
#251410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#251420000000
0!
0*
09
0>
0C
#251430000000
1!
1*
b101 6
19
1>
1C
b101 G
#251440000000
0!
0*
09
0>
0C
#251450000000
1!
1*
b110 6
19
1>
1C
b110 G
#251460000000
0!
0*
09
0>
0C
#251470000000
1!
1*
b111 6
19
1>
1C
b111 G
#251480000000
0!
0*
09
0>
0C
#251490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#251500000000
0!
0*
09
0>
0C
#251510000000
1!
1*
b1 6
19
1>
1C
b1 G
#251520000000
0!
0*
09
0>
0C
#251530000000
1!
1*
b10 6
19
1>
1C
b10 G
#251540000000
0!
0*
09
0>
0C
#251550000000
1!
1*
b11 6
19
1>
1C
b11 G
#251560000000
0!
0*
09
0>
0C
#251570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#251580000000
0!
0*
09
0>
0C
#251590000000
1!
1*
b101 6
19
1>
1C
b101 G
#251600000000
0!
0*
09
0>
0C
#251610000000
1!
1*
b110 6
19
1>
1C
b110 G
#251620000000
0!
0*
09
0>
0C
#251630000000
1!
1*
b111 6
19
1>
1C
b111 G
#251640000000
0!
1"
0*
1+
09
1:
0>
0C
#251650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#251660000000
0!
0*
09
0>
0C
#251670000000
1!
1*
b1 6
19
1>
1C
b1 G
#251680000000
0!
0*
09
0>
0C
#251690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#251700000000
0!
0*
09
0>
0C
#251710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#251720000000
0!
0*
09
0>
0C
#251730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#251740000000
0!
0*
09
0>
0C
#251750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#251760000000
0!
0#
0*
0,
09
0>
0?
0C
#251770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#251780000000
0!
0*
09
0>
0C
#251790000000
1!
1*
19
1>
1C
#251800000000
0!
0*
09
0>
0C
#251810000000
1!
1*
19
1>
1C
#251820000000
0!
0*
09
0>
0C
#251830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#251840000000
0!
0*
09
0>
0C
#251850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#251860000000
0!
0*
09
0>
0C
#251870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#251880000000
0!
0*
09
0>
0C
#251890000000
1!
1*
b10 6
19
1>
1C
b10 G
#251900000000
0!
0*
09
0>
0C
#251910000000
1!
1*
b11 6
19
1>
1C
b11 G
#251920000000
0!
0*
09
0>
0C
#251930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#251940000000
0!
0*
09
0>
0C
#251950000000
1!
1*
b101 6
19
1>
1C
b101 G
#251960000000
0!
0*
09
0>
0C
#251970000000
1!
1*
b110 6
19
1>
1C
b110 G
#251980000000
0!
0*
09
0>
0C
#251990000000
1!
1*
b111 6
19
1>
1C
b111 G
#252000000000
0!
0*
09
0>
0C
#252010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#252020000000
0!
0*
09
0>
0C
#252030000000
1!
1*
b1 6
19
1>
1C
b1 G
#252040000000
0!
0*
09
0>
0C
#252050000000
1!
1*
b10 6
19
1>
1C
b10 G
#252060000000
0!
0*
09
0>
0C
#252070000000
1!
1*
b11 6
19
1>
1C
b11 G
#252080000000
0!
0*
09
0>
0C
#252090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#252100000000
0!
0*
09
0>
0C
#252110000000
1!
1*
b101 6
19
1>
1C
b101 G
#252120000000
0!
0*
09
0>
0C
#252130000000
1!
1*
b110 6
19
1>
1C
b110 G
#252140000000
0!
0*
09
0>
0C
#252150000000
1!
1*
b111 6
19
1>
1C
b111 G
#252160000000
0!
0*
09
0>
0C
#252170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#252180000000
0!
0*
09
0>
0C
#252190000000
1!
1*
b1 6
19
1>
1C
b1 G
#252200000000
0!
0*
09
0>
0C
#252210000000
1!
1*
b10 6
19
1>
1C
b10 G
#252220000000
0!
0*
09
0>
0C
#252230000000
1!
1*
b11 6
19
1>
1C
b11 G
#252240000000
0!
0*
09
0>
0C
#252250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#252260000000
0!
0*
09
0>
0C
#252270000000
1!
1*
b101 6
19
1>
1C
b101 G
#252280000000
0!
0*
09
0>
0C
#252290000000
1!
1*
b110 6
19
1>
1C
b110 G
#252300000000
0!
0*
09
0>
0C
#252310000000
1!
1*
b111 6
19
1>
1C
b111 G
#252320000000
0!
1"
0*
1+
09
1:
0>
0C
#252330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#252340000000
0!
0*
09
0>
0C
#252350000000
1!
1*
b1 6
19
1>
1C
b1 G
#252360000000
0!
0*
09
0>
0C
#252370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#252380000000
0!
0*
09
0>
0C
#252390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#252400000000
0!
0*
09
0>
0C
#252410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#252420000000
0!
0*
09
0>
0C
#252430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#252440000000
0!
0#
0*
0,
09
0>
0?
0C
#252450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#252460000000
0!
0*
09
0>
0C
#252470000000
1!
1*
19
1>
1C
#252480000000
0!
0*
09
0>
0C
#252490000000
1!
1*
19
1>
1C
#252500000000
0!
0*
09
0>
0C
#252510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#252520000000
0!
0*
09
0>
0C
#252530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#252540000000
0!
0*
09
0>
0C
#252550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#252560000000
0!
0*
09
0>
0C
#252570000000
1!
1*
b10 6
19
1>
1C
b10 G
#252580000000
0!
0*
09
0>
0C
#252590000000
1!
1*
b11 6
19
1>
1C
b11 G
#252600000000
0!
0*
09
0>
0C
#252610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#252620000000
0!
0*
09
0>
0C
#252630000000
1!
1*
b101 6
19
1>
1C
b101 G
#252640000000
0!
0*
09
0>
0C
#252650000000
1!
1*
b110 6
19
1>
1C
b110 G
#252660000000
0!
0*
09
0>
0C
#252670000000
1!
1*
b111 6
19
1>
1C
b111 G
#252680000000
0!
0*
09
0>
0C
#252690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#252700000000
0!
0*
09
0>
0C
#252710000000
1!
1*
b1 6
19
1>
1C
b1 G
#252720000000
0!
0*
09
0>
0C
#252730000000
1!
1*
b10 6
19
1>
1C
b10 G
#252740000000
0!
0*
09
0>
0C
#252750000000
1!
1*
b11 6
19
1>
1C
b11 G
#252760000000
0!
0*
09
0>
0C
#252770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#252780000000
0!
0*
09
0>
0C
#252790000000
1!
1*
b101 6
19
1>
1C
b101 G
#252800000000
0!
0*
09
0>
0C
#252810000000
1!
1*
b110 6
19
1>
1C
b110 G
#252820000000
0!
0*
09
0>
0C
#252830000000
1!
1*
b111 6
19
1>
1C
b111 G
#252840000000
0!
0*
09
0>
0C
#252850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#252860000000
0!
0*
09
0>
0C
#252870000000
1!
1*
b1 6
19
1>
1C
b1 G
#252880000000
0!
0*
09
0>
0C
#252890000000
1!
1*
b10 6
19
1>
1C
b10 G
#252900000000
0!
0*
09
0>
0C
#252910000000
1!
1*
b11 6
19
1>
1C
b11 G
#252920000000
0!
0*
09
0>
0C
#252930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#252940000000
0!
0*
09
0>
0C
#252950000000
1!
1*
b101 6
19
1>
1C
b101 G
#252960000000
0!
0*
09
0>
0C
#252970000000
1!
1*
b110 6
19
1>
1C
b110 G
#252980000000
0!
0*
09
0>
0C
#252990000000
1!
1*
b111 6
19
1>
1C
b111 G
#253000000000
0!
1"
0*
1+
09
1:
0>
0C
#253010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#253020000000
0!
0*
09
0>
0C
#253030000000
1!
1*
b1 6
19
1>
1C
b1 G
#253040000000
0!
0*
09
0>
0C
#253050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#253060000000
0!
0*
09
0>
0C
#253070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#253080000000
0!
0*
09
0>
0C
#253090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#253100000000
0!
0*
09
0>
0C
#253110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#253120000000
0!
0#
0*
0,
09
0>
0?
0C
#253130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#253140000000
0!
0*
09
0>
0C
#253150000000
1!
1*
19
1>
1C
#253160000000
0!
0*
09
0>
0C
#253170000000
1!
1*
19
1>
1C
#253180000000
0!
0*
09
0>
0C
#253190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#253200000000
0!
0*
09
0>
0C
#253210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#253220000000
0!
0*
09
0>
0C
#253230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#253240000000
0!
0*
09
0>
0C
#253250000000
1!
1*
b10 6
19
1>
1C
b10 G
#253260000000
0!
0*
09
0>
0C
#253270000000
1!
1*
b11 6
19
1>
1C
b11 G
#253280000000
0!
0*
09
0>
0C
#253290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#253300000000
0!
0*
09
0>
0C
#253310000000
1!
1*
b101 6
19
1>
1C
b101 G
#253320000000
0!
0*
09
0>
0C
#253330000000
1!
1*
b110 6
19
1>
1C
b110 G
#253340000000
0!
0*
09
0>
0C
#253350000000
1!
1*
b111 6
19
1>
1C
b111 G
#253360000000
0!
0*
09
0>
0C
#253370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#253380000000
0!
0*
09
0>
0C
#253390000000
1!
1*
b1 6
19
1>
1C
b1 G
#253400000000
0!
0*
09
0>
0C
#253410000000
1!
1*
b10 6
19
1>
1C
b10 G
#253420000000
0!
0*
09
0>
0C
#253430000000
1!
1*
b11 6
19
1>
1C
b11 G
#253440000000
0!
0*
09
0>
0C
#253450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#253460000000
0!
0*
09
0>
0C
#253470000000
1!
1*
b101 6
19
1>
1C
b101 G
#253480000000
0!
0*
09
0>
0C
#253490000000
1!
1*
b110 6
19
1>
1C
b110 G
#253500000000
0!
0*
09
0>
0C
#253510000000
1!
1*
b111 6
19
1>
1C
b111 G
#253520000000
0!
0*
09
0>
0C
#253530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#253540000000
0!
0*
09
0>
0C
#253550000000
1!
1*
b1 6
19
1>
1C
b1 G
#253560000000
0!
0*
09
0>
0C
#253570000000
1!
1*
b10 6
19
1>
1C
b10 G
#253580000000
0!
0*
09
0>
0C
#253590000000
1!
1*
b11 6
19
1>
1C
b11 G
#253600000000
0!
0*
09
0>
0C
#253610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#253620000000
0!
0*
09
0>
0C
#253630000000
1!
1*
b101 6
19
1>
1C
b101 G
#253640000000
0!
0*
09
0>
0C
#253650000000
1!
1*
b110 6
19
1>
1C
b110 G
#253660000000
0!
0*
09
0>
0C
#253670000000
1!
1*
b111 6
19
1>
1C
b111 G
#253680000000
0!
1"
0*
1+
09
1:
0>
0C
#253690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#253700000000
0!
0*
09
0>
0C
#253710000000
1!
1*
b1 6
19
1>
1C
b1 G
#253720000000
0!
0*
09
0>
0C
#253730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#253740000000
0!
0*
09
0>
0C
#253750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#253760000000
0!
0*
09
0>
0C
#253770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#253780000000
0!
0*
09
0>
0C
#253790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#253800000000
0!
0#
0*
0,
09
0>
0?
0C
#253810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#253820000000
0!
0*
09
0>
0C
#253830000000
1!
1*
19
1>
1C
#253840000000
0!
0*
09
0>
0C
#253850000000
1!
1*
19
1>
1C
#253860000000
0!
0*
09
0>
0C
#253870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#253880000000
0!
0*
09
0>
0C
#253890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#253900000000
0!
0*
09
0>
0C
#253910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#253920000000
0!
0*
09
0>
0C
#253930000000
1!
1*
b10 6
19
1>
1C
b10 G
#253940000000
0!
0*
09
0>
0C
#253950000000
1!
1*
b11 6
19
1>
1C
b11 G
#253960000000
0!
0*
09
0>
0C
#253970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#253980000000
0!
0*
09
0>
0C
#253990000000
1!
1*
b101 6
19
1>
1C
b101 G
#254000000000
0!
0*
09
0>
0C
#254010000000
1!
1*
b110 6
19
1>
1C
b110 G
#254020000000
0!
0*
09
0>
0C
#254030000000
1!
1*
b111 6
19
1>
1C
b111 G
#254040000000
0!
0*
09
0>
0C
#254050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#254060000000
0!
0*
09
0>
0C
#254070000000
1!
1*
b1 6
19
1>
1C
b1 G
#254080000000
0!
0*
09
0>
0C
#254090000000
1!
1*
b10 6
19
1>
1C
b10 G
#254100000000
0!
0*
09
0>
0C
#254110000000
1!
1*
b11 6
19
1>
1C
b11 G
#254120000000
0!
0*
09
0>
0C
#254130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#254140000000
0!
0*
09
0>
0C
#254150000000
1!
1*
b101 6
19
1>
1C
b101 G
#254160000000
0!
0*
09
0>
0C
#254170000000
1!
1*
b110 6
19
1>
1C
b110 G
#254180000000
0!
0*
09
0>
0C
#254190000000
1!
1*
b111 6
19
1>
1C
b111 G
#254200000000
0!
0*
09
0>
0C
#254210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#254220000000
0!
0*
09
0>
0C
#254230000000
1!
1*
b1 6
19
1>
1C
b1 G
#254240000000
0!
0*
09
0>
0C
#254250000000
1!
1*
b10 6
19
1>
1C
b10 G
#254260000000
0!
0*
09
0>
0C
#254270000000
1!
1*
b11 6
19
1>
1C
b11 G
#254280000000
0!
0*
09
0>
0C
#254290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#254300000000
0!
0*
09
0>
0C
#254310000000
1!
1*
b101 6
19
1>
1C
b101 G
#254320000000
0!
0*
09
0>
0C
#254330000000
1!
1*
b110 6
19
1>
1C
b110 G
#254340000000
0!
0*
09
0>
0C
#254350000000
1!
1*
b111 6
19
1>
1C
b111 G
#254360000000
0!
1"
0*
1+
09
1:
0>
0C
#254370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#254380000000
0!
0*
09
0>
0C
#254390000000
1!
1*
b1 6
19
1>
1C
b1 G
#254400000000
0!
0*
09
0>
0C
#254410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#254420000000
0!
0*
09
0>
0C
#254430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#254440000000
0!
0*
09
0>
0C
#254450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#254460000000
0!
0*
09
0>
0C
#254470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#254480000000
0!
0#
0*
0,
09
0>
0?
0C
#254490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#254500000000
0!
0*
09
0>
0C
#254510000000
1!
1*
19
1>
1C
#254520000000
0!
0*
09
0>
0C
#254530000000
1!
1*
19
1>
1C
#254540000000
0!
0*
09
0>
0C
#254550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#254560000000
0!
0*
09
0>
0C
#254570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#254580000000
0!
0*
09
0>
0C
#254590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#254600000000
0!
0*
09
0>
0C
#254610000000
1!
1*
b10 6
19
1>
1C
b10 G
#254620000000
0!
0*
09
0>
0C
#254630000000
1!
1*
b11 6
19
1>
1C
b11 G
#254640000000
0!
0*
09
0>
0C
#254650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#254660000000
0!
0*
09
0>
0C
#254670000000
1!
1*
b101 6
19
1>
1C
b101 G
#254680000000
0!
0*
09
0>
0C
#254690000000
1!
1*
b110 6
19
1>
1C
b110 G
#254700000000
0!
0*
09
0>
0C
#254710000000
1!
1*
b111 6
19
1>
1C
b111 G
#254720000000
0!
0*
09
0>
0C
#254730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#254740000000
0!
0*
09
0>
0C
#254750000000
1!
1*
b1 6
19
1>
1C
b1 G
#254760000000
0!
0*
09
0>
0C
#254770000000
1!
1*
b10 6
19
1>
1C
b10 G
#254780000000
0!
0*
09
0>
0C
#254790000000
1!
1*
b11 6
19
1>
1C
b11 G
#254800000000
0!
0*
09
0>
0C
#254810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#254820000000
0!
0*
09
0>
0C
#254830000000
1!
1*
b101 6
19
1>
1C
b101 G
#254840000000
0!
0*
09
0>
0C
#254850000000
1!
1*
b110 6
19
1>
1C
b110 G
#254860000000
0!
0*
09
0>
0C
#254870000000
1!
1*
b111 6
19
1>
1C
b111 G
#254880000000
0!
0*
09
0>
0C
#254890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#254900000000
0!
0*
09
0>
0C
#254910000000
1!
1*
b1 6
19
1>
1C
b1 G
#254920000000
0!
0*
09
0>
0C
#254930000000
1!
1*
b10 6
19
1>
1C
b10 G
#254940000000
0!
0*
09
0>
0C
#254950000000
1!
1*
b11 6
19
1>
1C
b11 G
#254960000000
0!
0*
09
0>
0C
#254970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#254980000000
0!
0*
09
0>
0C
#254990000000
1!
1*
b101 6
19
1>
1C
b101 G
#255000000000
0!
0*
09
0>
0C
#255010000000
1!
1*
b110 6
19
1>
1C
b110 G
#255020000000
0!
0*
09
0>
0C
#255030000000
1!
1*
b111 6
19
1>
1C
b111 G
#255040000000
0!
1"
0*
1+
09
1:
0>
0C
#255050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#255060000000
0!
0*
09
0>
0C
#255070000000
1!
1*
b1 6
19
1>
1C
b1 G
#255080000000
0!
0*
09
0>
0C
#255090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#255100000000
0!
0*
09
0>
0C
#255110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#255120000000
0!
0*
09
0>
0C
#255130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#255140000000
0!
0*
09
0>
0C
#255150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#255160000000
0!
0#
0*
0,
09
0>
0?
0C
#255170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#255180000000
0!
0*
09
0>
0C
#255190000000
1!
1*
19
1>
1C
#255200000000
0!
0*
09
0>
0C
#255210000000
1!
1*
19
1>
1C
#255220000000
0!
0*
09
0>
0C
#255230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#255240000000
0!
0*
09
0>
0C
#255250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#255260000000
0!
0*
09
0>
0C
#255270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#255280000000
0!
0*
09
0>
0C
#255290000000
1!
1*
b10 6
19
1>
1C
b10 G
#255300000000
0!
0*
09
0>
0C
#255310000000
1!
1*
b11 6
19
1>
1C
b11 G
#255320000000
0!
0*
09
0>
0C
#255330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#255340000000
0!
0*
09
0>
0C
#255350000000
1!
1*
b101 6
19
1>
1C
b101 G
#255360000000
0!
0*
09
0>
0C
#255370000000
1!
1*
b110 6
19
1>
1C
b110 G
#255380000000
0!
0*
09
0>
0C
#255390000000
1!
1*
b111 6
19
1>
1C
b111 G
#255400000000
0!
0*
09
0>
0C
#255410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#255420000000
0!
0*
09
0>
0C
#255430000000
1!
1*
b1 6
19
1>
1C
b1 G
#255440000000
0!
0*
09
0>
0C
#255450000000
1!
1*
b10 6
19
1>
1C
b10 G
#255460000000
0!
0*
09
0>
0C
#255470000000
1!
1*
b11 6
19
1>
1C
b11 G
#255480000000
0!
0*
09
0>
0C
#255490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#255500000000
0!
0*
09
0>
0C
#255510000000
1!
1*
b101 6
19
1>
1C
b101 G
#255520000000
0!
0*
09
0>
0C
#255530000000
1!
1*
b110 6
19
1>
1C
b110 G
#255540000000
0!
0*
09
0>
0C
#255550000000
1!
1*
b111 6
19
1>
1C
b111 G
#255560000000
0!
0*
09
0>
0C
#255570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#255580000000
0!
0*
09
0>
0C
#255590000000
1!
1*
b1 6
19
1>
1C
b1 G
#255600000000
0!
0*
09
0>
0C
#255610000000
1!
1*
b10 6
19
1>
1C
b10 G
#255620000000
0!
0*
09
0>
0C
#255630000000
1!
1*
b11 6
19
1>
1C
b11 G
#255640000000
0!
0*
09
0>
0C
#255650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#255660000000
0!
0*
09
0>
0C
#255670000000
1!
1*
b101 6
19
1>
1C
b101 G
#255680000000
0!
0*
09
0>
0C
#255690000000
1!
1*
b110 6
19
1>
1C
b110 G
#255700000000
0!
0*
09
0>
0C
#255710000000
1!
1*
b111 6
19
1>
1C
b111 G
#255720000000
0!
1"
0*
1+
09
1:
0>
0C
#255730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#255740000000
0!
0*
09
0>
0C
#255750000000
1!
1*
b1 6
19
1>
1C
b1 G
#255760000000
0!
0*
09
0>
0C
#255770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#255780000000
0!
0*
09
0>
0C
#255790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#255800000000
0!
0*
09
0>
0C
#255810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#255820000000
0!
0*
09
0>
0C
#255830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#255840000000
0!
0#
0*
0,
09
0>
0?
0C
#255850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#255860000000
0!
0*
09
0>
0C
#255870000000
1!
1*
19
1>
1C
#255880000000
0!
0*
09
0>
0C
#255890000000
1!
1*
19
1>
1C
#255900000000
0!
0*
09
0>
0C
#255910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#255920000000
0!
0*
09
0>
0C
#255930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#255940000000
0!
0*
09
0>
0C
#255950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#255960000000
0!
0*
09
0>
0C
#255970000000
1!
1*
b10 6
19
1>
1C
b10 G
#255980000000
0!
0*
09
0>
0C
#255990000000
1!
1*
b11 6
19
1>
1C
b11 G
#256000000000
0!
0*
09
0>
0C
#256010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#256020000000
0!
0*
09
0>
0C
#256030000000
1!
1*
b101 6
19
1>
1C
b101 G
#256040000000
0!
0*
09
0>
0C
#256050000000
1!
1*
b110 6
19
1>
1C
b110 G
#256060000000
0!
0*
09
0>
0C
#256070000000
1!
1*
b111 6
19
1>
1C
b111 G
#256080000000
0!
0*
09
0>
0C
#256090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#256100000000
0!
0*
09
0>
0C
#256110000000
1!
1*
b1 6
19
1>
1C
b1 G
#256120000000
0!
0*
09
0>
0C
#256130000000
1!
1*
b10 6
19
1>
1C
b10 G
#256140000000
0!
0*
09
0>
0C
#256150000000
1!
1*
b11 6
19
1>
1C
b11 G
#256160000000
0!
0*
09
0>
0C
#256170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#256180000000
0!
0*
09
0>
0C
#256190000000
1!
1*
b101 6
19
1>
1C
b101 G
#256200000000
0!
0*
09
0>
0C
#256210000000
1!
1*
b110 6
19
1>
1C
b110 G
#256220000000
0!
0*
09
0>
0C
#256230000000
1!
1*
b111 6
19
1>
1C
b111 G
#256240000000
0!
0*
09
0>
0C
#256250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#256260000000
0!
0*
09
0>
0C
#256270000000
1!
1*
b1 6
19
1>
1C
b1 G
#256280000000
0!
0*
09
0>
0C
#256290000000
1!
1*
b10 6
19
1>
1C
b10 G
#256300000000
0!
0*
09
0>
0C
#256310000000
1!
1*
b11 6
19
1>
1C
b11 G
#256320000000
0!
0*
09
0>
0C
#256330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#256340000000
0!
0*
09
0>
0C
#256350000000
1!
1*
b101 6
19
1>
1C
b101 G
#256360000000
0!
0*
09
0>
0C
#256370000000
1!
1*
b110 6
19
1>
1C
b110 G
#256380000000
0!
0*
09
0>
0C
#256390000000
1!
1*
b111 6
19
1>
1C
b111 G
#256400000000
0!
1"
0*
1+
09
1:
0>
0C
#256410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#256420000000
0!
0*
09
0>
0C
#256430000000
1!
1*
b1 6
19
1>
1C
b1 G
#256440000000
0!
0*
09
0>
0C
#256450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#256460000000
0!
0*
09
0>
0C
#256470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#256480000000
0!
0*
09
0>
0C
#256490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#256500000000
0!
0*
09
0>
0C
#256510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#256520000000
0!
0#
0*
0,
09
0>
0?
0C
#256530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#256540000000
0!
0*
09
0>
0C
#256550000000
1!
1*
19
1>
1C
#256560000000
0!
0*
09
0>
0C
#256570000000
1!
1*
19
1>
1C
#256580000000
0!
0*
09
0>
0C
#256590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#256600000000
0!
0*
09
0>
0C
#256610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#256620000000
0!
0*
09
0>
0C
#256630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#256640000000
0!
0*
09
0>
0C
#256650000000
1!
1*
b10 6
19
1>
1C
b10 G
#256660000000
0!
0*
09
0>
0C
#256670000000
1!
1*
b11 6
19
1>
1C
b11 G
#256680000000
0!
0*
09
0>
0C
#256690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#256700000000
0!
0*
09
0>
0C
#256710000000
1!
1*
b101 6
19
1>
1C
b101 G
#256720000000
0!
0*
09
0>
0C
#256730000000
1!
1*
b110 6
19
1>
1C
b110 G
#256740000000
0!
0*
09
0>
0C
#256750000000
1!
1*
b111 6
19
1>
1C
b111 G
#256760000000
0!
0*
09
0>
0C
#256770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#256780000000
0!
0*
09
0>
0C
#256790000000
1!
1*
b1 6
19
1>
1C
b1 G
#256800000000
0!
0*
09
0>
0C
#256810000000
1!
1*
b10 6
19
1>
1C
b10 G
#256820000000
0!
0*
09
0>
0C
#256830000000
1!
1*
b11 6
19
1>
1C
b11 G
#256840000000
0!
0*
09
0>
0C
#256850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#256860000000
0!
0*
09
0>
0C
#256870000000
1!
1*
b101 6
19
1>
1C
b101 G
#256880000000
0!
0*
09
0>
0C
#256890000000
1!
1*
b110 6
19
1>
1C
b110 G
#256900000000
0!
0*
09
0>
0C
#256910000000
1!
1*
b111 6
19
1>
1C
b111 G
#256920000000
0!
0*
09
0>
0C
#256930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#256940000000
0!
0*
09
0>
0C
#256950000000
1!
1*
b1 6
19
1>
1C
b1 G
#256960000000
0!
0*
09
0>
0C
#256970000000
1!
1*
b10 6
19
1>
1C
b10 G
#256980000000
0!
0*
09
0>
0C
#256990000000
1!
1*
b11 6
19
1>
1C
b11 G
#257000000000
0!
0*
09
0>
0C
#257010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#257020000000
0!
0*
09
0>
0C
#257030000000
1!
1*
b101 6
19
1>
1C
b101 G
#257040000000
0!
0*
09
0>
0C
#257050000000
1!
1*
b110 6
19
1>
1C
b110 G
#257060000000
0!
0*
09
0>
0C
#257070000000
1!
1*
b111 6
19
1>
1C
b111 G
#257080000000
0!
1"
0*
1+
09
1:
0>
0C
#257090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#257100000000
0!
0*
09
0>
0C
#257110000000
1!
1*
b1 6
19
1>
1C
b1 G
#257120000000
0!
0*
09
0>
0C
#257130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#257140000000
0!
0*
09
0>
0C
#257150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#257160000000
0!
0*
09
0>
0C
#257170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#257180000000
0!
0*
09
0>
0C
#257190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#257200000000
0!
0#
0*
0,
09
0>
0?
0C
#257210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#257220000000
0!
0*
09
0>
0C
#257230000000
1!
1*
19
1>
1C
#257240000000
0!
0*
09
0>
0C
#257250000000
1!
1*
19
1>
1C
#257260000000
0!
0*
09
0>
0C
#257270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#257280000000
0!
0*
09
0>
0C
#257290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#257300000000
0!
0*
09
0>
0C
#257310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#257320000000
0!
0*
09
0>
0C
#257330000000
1!
1*
b10 6
19
1>
1C
b10 G
#257340000000
0!
0*
09
0>
0C
#257350000000
1!
1*
b11 6
19
1>
1C
b11 G
#257360000000
0!
0*
09
0>
0C
#257370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#257380000000
0!
0*
09
0>
0C
#257390000000
1!
1*
b101 6
19
1>
1C
b101 G
#257400000000
0!
0*
09
0>
0C
#257410000000
1!
1*
b110 6
19
1>
1C
b110 G
#257420000000
0!
0*
09
0>
0C
#257430000000
1!
1*
b111 6
19
1>
1C
b111 G
#257440000000
0!
0*
09
0>
0C
#257450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#257460000000
0!
0*
09
0>
0C
#257470000000
1!
1*
b1 6
19
1>
1C
b1 G
#257480000000
0!
0*
09
0>
0C
#257490000000
1!
1*
b10 6
19
1>
1C
b10 G
#257500000000
0!
0*
09
0>
0C
#257510000000
1!
1*
b11 6
19
1>
1C
b11 G
#257520000000
0!
0*
09
0>
0C
#257530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#257540000000
0!
0*
09
0>
0C
#257550000000
1!
1*
b101 6
19
1>
1C
b101 G
#257560000000
0!
0*
09
0>
0C
#257570000000
1!
1*
b110 6
19
1>
1C
b110 G
#257580000000
0!
0*
09
0>
0C
#257590000000
1!
1*
b111 6
19
1>
1C
b111 G
#257600000000
0!
0*
09
0>
0C
#257610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#257620000000
0!
0*
09
0>
0C
#257630000000
1!
1*
b1 6
19
1>
1C
b1 G
#257640000000
0!
0*
09
0>
0C
#257650000000
1!
1*
b10 6
19
1>
1C
b10 G
#257660000000
0!
0*
09
0>
0C
#257670000000
1!
1*
b11 6
19
1>
1C
b11 G
#257680000000
0!
0*
09
0>
0C
#257690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#257700000000
0!
0*
09
0>
0C
#257710000000
1!
1*
b101 6
19
1>
1C
b101 G
#257720000000
0!
0*
09
0>
0C
#257730000000
1!
1*
b110 6
19
1>
1C
b110 G
#257740000000
0!
0*
09
0>
0C
#257750000000
1!
1*
b111 6
19
1>
1C
b111 G
#257760000000
0!
1"
0*
1+
09
1:
0>
0C
#257770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#257780000000
0!
0*
09
0>
0C
#257790000000
1!
1*
b1 6
19
1>
1C
b1 G
#257800000000
0!
0*
09
0>
0C
#257810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#257820000000
0!
0*
09
0>
0C
#257830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#257840000000
0!
0*
09
0>
0C
#257850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#257860000000
0!
0*
09
0>
0C
#257870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#257880000000
0!
0#
0*
0,
09
0>
0?
0C
#257890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#257900000000
0!
0*
09
0>
0C
#257910000000
1!
1*
19
1>
1C
#257920000000
0!
0*
09
0>
0C
#257930000000
1!
1*
19
1>
1C
#257940000000
0!
0*
09
0>
0C
#257950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#257960000000
0!
0*
09
0>
0C
#257970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#257980000000
0!
0*
09
0>
0C
#257990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#258000000000
0!
0*
09
0>
0C
#258010000000
1!
1*
b10 6
19
1>
1C
b10 G
#258020000000
0!
0*
09
0>
0C
#258030000000
1!
1*
b11 6
19
1>
1C
b11 G
#258040000000
0!
0*
09
0>
0C
#258050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#258060000000
0!
0*
09
0>
0C
#258070000000
1!
1*
b101 6
19
1>
1C
b101 G
#258080000000
0!
0*
09
0>
0C
#258090000000
1!
1*
b110 6
19
1>
1C
b110 G
#258100000000
0!
0*
09
0>
0C
#258110000000
1!
1*
b111 6
19
1>
1C
b111 G
#258120000000
0!
0*
09
0>
0C
#258130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#258140000000
0!
0*
09
0>
0C
#258150000000
1!
1*
b1 6
19
1>
1C
b1 G
#258160000000
0!
0*
09
0>
0C
#258170000000
1!
1*
b10 6
19
1>
1C
b10 G
#258180000000
0!
0*
09
0>
0C
#258190000000
1!
1*
b11 6
19
1>
1C
b11 G
#258200000000
0!
0*
09
0>
0C
#258210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#258220000000
0!
0*
09
0>
0C
#258230000000
1!
1*
b101 6
19
1>
1C
b101 G
#258240000000
0!
0*
09
0>
0C
#258250000000
1!
1*
b110 6
19
1>
1C
b110 G
#258260000000
0!
0*
09
0>
0C
#258270000000
1!
1*
b111 6
19
1>
1C
b111 G
#258280000000
0!
0*
09
0>
0C
#258290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#258300000000
0!
0*
09
0>
0C
#258310000000
1!
1*
b1 6
19
1>
1C
b1 G
#258320000000
0!
0*
09
0>
0C
#258330000000
1!
1*
b10 6
19
1>
1C
b10 G
#258340000000
0!
0*
09
0>
0C
#258350000000
1!
1*
b11 6
19
1>
1C
b11 G
#258360000000
0!
0*
09
0>
0C
#258370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#258380000000
0!
0*
09
0>
0C
#258390000000
1!
1*
b101 6
19
1>
1C
b101 G
#258400000000
0!
0*
09
0>
0C
#258410000000
1!
1*
b110 6
19
1>
1C
b110 G
#258420000000
0!
0*
09
0>
0C
#258430000000
1!
1*
b111 6
19
1>
1C
b111 G
#258440000000
0!
1"
0*
1+
09
1:
0>
0C
#258450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#258460000000
0!
0*
09
0>
0C
#258470000000
1!
1*
b1 6
19
1>
1C
b1 G
#258480000000
0!
0*
09
0>
0C
#258490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#258500000000
0!
0*
09
0>
0C
#258510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#258520000000
0!
0*
09
0>
0C
#258530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#258540000000
0!
0*
09
0>
0C
#258550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#258560000000
0!
0#
0*
0,
09
0>
0?
0C
#258570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#258580000000
0!
0*
09
0>
0C
#258590000000
1!
1*
19
1>
1C
#258600000000
0!
0*
09
0>
0C
#258610000000
1!
1*
19
1>
1C
#258620000000
0!
0*
09
0>
0C
#258630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#258640000000
0!
0*
09
0>
0C
#258650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#258660000000
0!
0*
09
0>
0C
#258670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#258680000000
0!
0*
09
0>
0C
#258690000000
1!
1*
b10 6
19
1>
1C
b10 G
#258700000000
0!
0*
09
0>
0C
#258710000000
1!
1*
b11 6
19
1>
1C
b11 G
#258720000000
0!
0*
09
0>
0C
#258730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#258740000000
0!
0*
09
0>
0C
#258750000000
1!
1*
b101 6
19
1>
1C
b101 G
#258760000000
0!
0*
09
0>
0C
#258770000000
1!
1*
b110 6
19
1>
1C
b110 G
#258780000000
0!
0*
09
0>
0C
#258790000000
1!
1*
b111 6
19
1>
1C
b111 G
#258800000000
0!
0*
09
0>
0C
#258810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#258820000000
0!
0*
09
0>
0C
#258830000000
1!
1*
b1 6
19
1>
1C
b1 G
#258840000000
0!
0*
09
0>
0C
#258850000000
1!
1*
b10 6
19
1>
1C
b10 G
#258860000000
0!
0*
09
0>
0C
#258870000000
1!
1*
b11 6
19
1>
1C
b11 G
#258880000000
0!
0*
09
0>
0C
#258890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#258900000000
0!
0*
09
0>
0C
#258910000000
1!
1*
b101 6
19
1>
1C
b101 G
#258920000000
0!
0*
09
0>
0C
#258930000000
1!
1*
b110 6
19
1>
1C
b110 G
#258940000000
0!
0*
09
0>
0C
#258950000000
1!
1*
b111 6
19
1>
1C
b111 G
#258960000000
0!
0*
09
0>
0C
#258970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#258980000000
0!
0*
09
0>
0C
#258990000000
1!
1*
b1 6
19
1>
1C
b1 G
#259000000000
0!
0*
09
0>
0C
#259010000000
1!
1*
b10 6
19
1>
1C
b10 G
#259020000000
0!
0*
09
0>
0C
#259030000000
1!
1*
b11 6
19
1>
1C
b11 G
#259040000000
0!
0*
09
0>
0C
#259050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#259060000000
0!
0*
09
0>
0C
#259070000000
1!
1*
b101 6
19
1>
1C
b101 G
#259080000000
0!
0*
09
0>
0C
#259090000000
1!
1*
b110 6
19
1>
1C
b110 G
#259100000000
0!
0*
09
0>
0C
#259110000000
1!
1*
b111 6
19
1>
1C
b111 G
#259120000000
0!
1"
0*
1+
09
1:
0>
0C
#259130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#259140000000
0!
0*
09
0>
0C
#259150000000
1!
1*
b1 6
19
1>
1C
b1 G
#259160000000
0!
0*
09
0>
0C
#259170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#259180000000
0!
0*
09
0>
0C
#259190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#259200000000
0!
0*
09
0>
0C
#259210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#259220000000
0!
0*
09
0>
0C
#259230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#259240000000
0!
0#
0*
0,
09
0>
0?
0C
#259250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#259260000000
0!
0*
09
0>
0C
#259270000000
1!
1*
19
1>
1C
#259280000000
0!
0*
09
0>
0C
#259290000000
1!
1*
19
1>
1C
#259300000000
0!
0*
09
0>
0C
#259310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#259320000000
0!
0*
09
0>
0C
#259330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#259340000000
0!
0*
09
0>
0C
#259350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#259360000000
0!
0*
09
0>
0C
#259370000000
1!
1*
b10 6
19
1>
1C
b10 G
#259380000000
0!
0*
09
0>
0C
#259390000000
1!
1*
b11 6
19
1>
1C
b11 G
#259400000000
0!
0*
09
0>
0C
#259410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#259420000000
0!
0*
09
0>
0C
#259430000000
1!
1*
b101 6
19
1>
1C
b101 G
#259440000000
0!
0*
09
0>
0C
#259450000000
1!
1*
b110 6
19
1>
1C
b110 G
#259460000000
0!
0*
09
0>
0C
#259470000000
1!
1*
b111 6
19
1>
1C
b111 G
#259480000000
0!
0*
09
0>
0C
#259490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#259500000000
0!
0*
09
0>
0C
#259510000000
1!
1*
b1 6
19
1>
1C
b1 G
#259520000000
0!
0*
09
0>
0C
#259530000000
1!
1*
b10 6
19
1>
1C
b10 G
#259540000000
0!
0*
09
0>
0C
#259550000000
1!
1*
b11 6
19
1>
1C
b11 G
#259560000000
0!
0*
09
0>
0C
#259570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#259580000000
0!
0*
09
0>
0C
#259590000000
1!
1*
b101 6
19
1>
1C
b101 G
#259600000000
0!
0*
09
0>
0C
#259610000000
1!
1*
b110 6
19
1>
1C
b110 G
#259620000000
0!
0*
09
0>
0C
#259630000000
1!
1*
b111 6
19
1>
1C
b111 G
#259640000000
0!
0*
09
0>
0C
#259650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#259660000000
0!
0*
09
0>
0C
#259670000000
1!
1*
b1 6
19
1>
1C
b1 G
#259680000000
0!
0*
09
0>
0C
#259690000000
1!
1*
b10 6
19
1>
1C
b10 G
#259700000000
0!
0*
09
0>
0C
#259710000000
1!
1*
b11 6
19
1>
1C
b11 G
#259720000000
0!
0*
09
0>
0C
#259730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#259740000000
0!
0*
09
0>
0C
#259750000000
1!
1*
b101 6
19
1>
1C
b101 G
#259760000000
0!
0*
09
0>
0C
#259770000000
1!
1*
b110 6
19
1>
1C
b110 G
#259780000000
0!
0*
09
0>
0C
#259790000000
1!
1*
b111 6
19
1>
1C
b111 G
#259800000000
0!
1"
0*
1+
09
1:
0>
0C
#259810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#259820000000
0!
0*
09
0>
0C
#259830000000
1!
1*
b1 6
19
1>
1C
b1 G
#259840000000
0!
0*
09
0>
0C
#259850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#259860000000
0!
0*
09
0>
0C
#259870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#259880000000
0!
0*
09
0>
0C
#259890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#259900000000
0!
0*
09
0>
0C
#259910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#259920000000
0!
0#
0*
0,
09
0>
0?
0C
#259930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#259940000000
0!
0*
09
0>
0C
#259950000000
1!
1*
19
1>
1C
#259960000000
0!
0*
09
0>
0C
#259970000000
1!
1*
19
1>
1C
#259980000000
0!
0*
09
0>
0C
#259990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#260000000000
0!
0*
09
0>
0C
#260010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#260020000000
0!
0*
09
0>
0C
#260030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#260040000000
0!
0*
09
0>
0C
#260050000000
1!
1*
b10 6
19
1>
1C
b10 G
#260060000000
0!
0*
09
0>
0C
#260070000000
1!
1*
b11 6
19
1>
1C
b11 G
#260080000000
0!
0*
09
0>
0C
#260090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#260100000000
0!
0*
09
0>
0C
#260110000000
1!
1*
b101 6
19
1>
1C
b101 G
#260120000000
0!
0*
09
0>
0C
#260130000000
1!
1*
b110 6
19
1>
1C
b110 G
#260140000000
0!
0*
09
0>
0C
#260150000000
1!
1*
b111 6
19
1>
1C
b111 G
#260160000000
0!
0*
09
0>
0C
#260170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#260180000000
0!
0*
09
0>
0C
#260190000000
1!
1*
b1 6
19
1>
1C
b1 G
#260200000000
0!
0*
09
0>
0C
#260210000000
1!
1*
b10 6
19
1>
1C
b10 G
#260220000000
0!
0*
09
0>
0C
#260230000000
1!
1*
b11 6
19
1>
1C
b11 G
#260240000000
0!
0*
09
0>
0C
#260250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#260260000000
0!
0*
09
0>
0C
#260270000000
1!
1*
b101 6
19
1>
1C
b101 G
#260280000000
0!
0*
09
0>
0C
#260290000000
1!
1*
b110 6
19
1>
1C
b110 G
#260300000000
0!
0*
09
0>
0C
#260310000000
1!
1*
b111 6
19
1>
1C
b111 G
#260320000000
0!
0*
09
0>
0C
#260330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#260340000000
0!
0*
09
0>
0C
#260350000000
1!
1*
b1 6
19
1>
1C
b1 G
#260360000000
0!
0*
09
0>
0C
#260370000000
1!
1*
b10 6
19
1>
1C
b10 G
#260380000000
0!
0*
09
0>
0C
#260390000000
1!
1*
b11 6
19
1>
1C
b11 G
#260400000000
0!
0*
09
0>
0C
#260410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#260420000000
0!
0*
09
0>
0C
#260430000000
1!
1*
b101 6
19
1>
1C
b101 G
#260440000000
0!
0*
09
0>
0C
#260450000000
1!
1*
b110 6
19
1>
1C
b110 G
#260460000000
0!
0*
09
0>
0C
#260470000000
1!
1*
b111 6
19
1>
1C
b111 G
#260480000000
0!
1"
0*
1+
09
1:
0>
0C
#260490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#260500000000
0!
0*
09
0>
0C
#260510000000
1!
1*
b1 6
19
1>
1C
b1 G
#260520000000
0!
0*
09
0>
0C
#260530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#260540000000
0!
0*
09
0>
0C
#260550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#260560000000
0!
0*
09
0>
0C
#260570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#260580000000
0!
0*
09
0>
0C
#260590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#260600000000
0!
0#
0*
0,
09
0>
0?
0C
#260610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#260620000000
0!
0*
09
0>
0C
#260630000000
1!
1*
19
1>
1C
#260640000000
0!
0*
09
0>
0C
#260650000000
1!
1*
19
1>
1C
#260660000000
0!
0*
09
0>
0C
#260670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#260680000000
0!
0*
09
0>
0C
#260690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#260700000000
0!
0*
09
0>
0C
#260710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#260720000000
0!
0*
09
0>
0C
#260730000000
1!
1*
b10 6
19
1>
1C
b10 G
#260740000000
0!
0*
09
0>
0C
#260750000000
1!
1*
b11 6
19
1>
1C
b11 G
#260760000000
0!
0*
09
0>
0C
#260770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#260780000000
0!
0*
09
0>
0C
#260790000000
1!
1*
b101 6
19
1>
1C
b101 G
#260800000000
0!
0*
09
0>
0C
#260810000000
1!
1*
b110 6
19
1>
1C
b110 G
#260820000000
0!
0*
09
0>
0C
#260830000000
1!
1*
b111 6
19
1>
1C
b111 G
#260840000000
0!
0*
09
0>
0C
#260850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#260860000000
0!
0*
09
0>
0C
#260870000000
1!
1*
b1 6
19
1>
1C
b1 G
#260880000000
0!
0*
09
0>
0C
#260890000000
1!
1*
b10 6
19
1>
1C
b10 G
#260900000000
0!
0*
09
0>
0C
#260910000000
1!
1*
b11 6
19
1>
1C
b11 G
#260920000000
0!
0*
09
0>
0C
#260930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#260940000000
0!
0*
09
0>
0C
#260950000000
1!
1*
b101 6
19
1>
1C
b101 G
#260960000000
0!
0*
09
0>
0C
#260970000000
1!
1*
b110 6
19
1>
1C
b110 G
#260980000000
0!
0*
09
0>
0C
#260990000000
1!
1*
b111 6
19
1>
1C
b111 G
#261000000000
0!
0*
09
0>
0C
#261010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#261020000000
0!
0*
09
0>
0C
#261030000000
1!
1*
b1 6
19
1>
1C
b1 G
#261040000000
0!
0*
09
0>
0C
#261050000000
1!
1*
b10 6
19
1>
1C
b10 G
#261060000000
0!
0*
09
0>
0C
#261070000000
1!
1*
b11 6
19
1>
1C
b11 G
#261080000000
0!
0*
09
0>
0C
#261090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#261100000000
0!
0*
09
0>
0C
#261110000000
1!
1*
b101 6
19
1>
1C
b101 G
#261120000000
0!
0*
09
0>
0C
#261130000000
1!
1*
b110 6
19
1>
1C
b110 G
#261140000000
0!
0*
09
0>
0C
#261150000000
1!
1*
b111 6
19
1>
1C
b111 G
#261160000000
0!
1"
0*
1+
09
1:
0>
0C
#261170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#261180000000
0!
0*
09
0>
0C
#261190000000
1!
1*
b1 6
19
1>
1C
b1 G
#261200000000
0!
0*
09
0>
0C
#261210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#261220000000
0!
0*
09
0>
0C
#261230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#261240000000
0!
0*
09
0>
0C
#261250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#261260000000
0!
0*
09
0>
0C
#261270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#261280000000
0!
0#
0*
0,
09
0>
0?
0C
#261290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#261300000000
0!
0*
09
0>
0C
#261310000000
1!
1*
19
1>
1C
#261320000000
0!
0*
09
0>
0C
#261330000000
1!
1*
19
1>
1C
#261340000000
0!
0*
09
0>
0C
#261350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#261360000000
0!
0*
09
0>
0C
#261370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#261380000000
0!
0*
09
0>
0C
#261390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#261400000000
0!
0*
09
0>
0C
#261410000000
1!
1*
b10 6
19
1>
1C
b10 G
#261420000000
0!
0*
09
0>
0C
#261430000000
1!
1*
b11 6
19
1>
1C
b11 G
#261440000000
0!
0*
09
0>
0C
#261450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#261460000000
0!
0*
09
0>
0C
#261470000000
1!
1*
b101 6
19
1>
1C
b101 G
#261480000000
0!
0*
09
0>
0C
#261490000000
1!
1*
b110 6
19
1>
1C
b110 G
#261500000000
0!
0*
09
0>
0C
#261510000000
1!
1*
b111 6
19
1>
1C
b111 G
#261520000000
0!
0*
09
0>
0C
#261530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#261540000000
0!
0*
09
0>
0C
#261550000000
1!
1*
b1 6
19
1>
1C
b1 G
#261560000000
0!
0*
09
0>
0C
#261570000000
1!
1*
b10 6
19
1>
1C
b10 G
#261580000000
0!
0*
09
0>
0C
#261590000000
1!
1*
b11 6
19
1>
1C
b11 G
#261600000000
0!
0*
09
0>
0C
#261610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#261620000000
0!
0*
09
0>
0C
#261630000000
1!
1*
b101 6
19
1>
1C
b101 G
#261640000000
0!
0*
09
0>
0C
#261650000000
1!
1*
b110 6
19
1>
1C
b110 G
#261660000000
0!
0*
09
0>
0C
#261670000000
1!
1*
b111 6
19
1>
1C
b111 G
#261680000000
0!
0*
09
0>
0C
#261690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#261700000000
0!
0*
09
0>
0C
#261710000000
1!
1*
b1 6
19
1>
1C
b1 G
#261720000000
0!
0*
09
0>
0C
#261730000000
1!
1*
b10 6
19
1>
1C
b10 G
#261740000000
0!
0*
09
0>
0C
#261750000000
1!
1*
b11 6
19
1>
1C
b11 G
#261760000000
0!
0*
09
0>
0C
#261770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#261780000000
0!
0*
09
0>
0C
#261790000000
1!
1*
b101 6
19
1>
1C
b101 G
#261800000000
0!
0*
09
0>
0C
#261810000000
1!
1*
b110 6
19
1>
1C
b110 G
#261820000000
0!
0*
09
0>
0C
#261830000000
1!
1*
b111 6
19
1>
1C
b111 G
#261840000000
0!
1"
0*
1+
09
1:
0>
0C
#261850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#261860000000
0!
0*
09
0>
0C
#261870000000
1!
1*
b1 6
19
1>
1C
b1 G
#261880000000
0!
0*
09
0>
0C
#261890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#261900000000
0!
0*
09
0>
0C
#261910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#261920000000
0!
0*
09
0>
0C
#261930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#261940000000
0!
0*
09
0>
0C
#261950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#261960000000
0!
0#
0*
0,
09
0>
0?
0C
#261970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#261980000000
0!
0*
09
0>
0C
#261990000000
1!
1*
19
1>
1C
#262000000000
0!
0*
09
0>
0C
#262010000000
1!
1*
19
1>
1C
#262020000000
0!
0*
09
0>
0C
#262030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#262040000000
0!
0*
09
0>
0C
#262050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#262060000000
0!
0*
09
0>
0C
#262070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#262080000000
0!
0*
09
0>
0C
#262090000000
1!
1*
b10 6
19
1>
1C
b10 G
#262100000000
0!
0*
09
0>
0C
#262110000000
1!
1*
b11 6
19
1>
1C
b11 G
#262120000000
0!
0*
09
0>
0C
#262130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#262140000000
0!
0*
09
0>
0C
#262150000000
1!
1*
b101 6
19
1>
1C
b101 G
#262160000000
0!
0*
09
0>
0C
#262170000000
1!
1*
b110 6
19
1>
1C
b110 G
#262180000000
0!
0*
09
0>
0C
#262190000000
1!
1*
b111 6
19
1>
1C
b111 G
#262200000000
0!
0*
09
0>
0C
#262210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#262220000000
0!
0*
09
0>
0C
#262230000000
1!
1*
b1 6
19
1>
1C
b1 G
#262240000000
0!
0*
09
0>
0C
#262250000000
1!
1*
b10 6
19
1>
1C
b10 G
#262260000000
0!
0*
09
0>
0C
#262270000000
1!
1*
b11 6
19
1>
1C
b11 G
#262280000000
0!
0*
09
0>
0C
#262290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#262300000000
0!
0*
09
0>
0C
#262310000000
1!
1*
b101 6
19
1>
1C
b101 G
#262320000000
0!
0*
09
0>
0C
#262330000000
1!
1*
b110 6
19
1>
1C
b110 G
#262340000000
0!
0*
09
0>
0C
#262350000000
1!
1*
b111 6
19
1>
1C
b111 G
#262360000000
0!
0*
09
0>
0C
#262370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#262380000000
0!
0*
09
0>
0C
#262390000000
1!
1*
b1 6
19
1>
1C
b1 G
#262400000000
0!
0*
09
0>
0C
#262410000000
1!
1*
b10 6
19
1>
1C
b10 G
#262420000000
0!
0*
09
0>
0C
#262430000000
1!
1*
b11 6
19
1>
1C
b11 G
#262440000000
0!
0*
09
0>
0C
#262450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#262460000000
0!
0*
09
0>
0C
#262470000000
1!
1*
b101 6
19
1>
1C
b101 G
#262480000000
0!
0*
09
0>
0C
#262490000000
1!
1*
b110 6
19
1>
1C
b110 G
#262500000000
0!
0*
09
0>
0C
#262510000000
1!
1*
b111 6
19
1>
1C
b111 G
#262520000000
0!
1"
0*
1+
09
1:
0>
0C
#262530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#262540000000
0!
0*
09
0>
0C
#262550000000
1!
1*
b1 6
19
1>
1C
b1 G
#262560000000
0!
0*
09
0>
0C
#262570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#262580000000
0!
0*
09
0>
0C
#262590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#262600000000
0!
0*
09
0>
0C
#262610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#262620000000
0!
0*
09
0>
0C
#262630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#262640000000
0!
0#
0*
0,
09
0>
0?
0C
#262650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#262660000000
0!
0*
09
0>
0C
#262670000000
1!
1*
19
1>
1C
#262680000000
0!
0*
09
0>
0C
#262690000000
1!
1*
19
1>
1C
#262700000000
0!
0*
09
0>
0C
#262710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#262720000000
0!
0*
09
0>
0C
#262730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#262740000000
0!
0*
09
0>
0C
#262750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#262760000000
0!
0*
09
0>
0C
#262770000000
1!
1*
b10 6
19
1>
1C
b10 G
#262780000000
0!
0*
09
0>
0C
#262790000000
1!
1*
b11 6
19
1>
1C
b11 G
#262800000000
0!
0*
09
0>
0C
#262810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#262820000000
0!
0*
09
0>
0C
#262830000000
1!
1*
b101 6
19
1>
1C
b101 G
#262840000000
0!
0*
09
0>
0C
#262850000000
1!
1*
b110 6
19
1>
1C
b110 G
#262860000000
0!
0*
09
0>
0C
#262870000000
1!
1*
b111 6
19
1>
1C
b111 G
#262880000000
0!
0*
09
0>
0C
#262890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#262900000000
0!
0*
09
0>
0C
#262910000000
1!
1*
b1 6
19
1>
1C
b1 G
#262920000000
0!
0*
09
0>
0C
#262930000000
1!
1*
b10 6
19
1>
1C
b10 G
#262940000000
0!
0*
09
0>
0C
#262950000000
1!
1*
b11 6
19
1>
1C
b11 G
#262960000000
0!
0*
09
0>
0C
#262970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#262980000000
0!
0*
09
0>
0C
#262990000000
1!
1*
b101 6
19
1>
1C
b101 G
#263000000000
0!
0*
09
0>
0C
#263010000000
1!
1*
b110 6
19
1>
1C
b110 G
#263020000000
0!
0*
09
0>
0C
#263030000000
1!
1*
b111 6
19
1>
1C
b111 G
#263040000000
0!
0*
09
0>
0C
#263050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#263060000000
0!
0*
09
0>
0C
#263070000000
1!
1*
b1 6
19
1>
1C
b1 G
#263080000000
0!
0*
09
0>
0C
#263090000000
1!
1*
b10 6
19
1>
1C
b10 G
#263100000000
0!
0*
09
0>
0C
#263110000000
1!
1*
b11 6
19
1>
1C
b11 G
#263120000000
0!
0*
09
0>
0C
#263130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#263140000000
0!
0*
09
0>
0C
#263150000000
1!
1*
b101 6
19
1>
1C
b101 G
#263160000000
0!
0*
09
0>
0C
#263170000000
1!
1*
b110 6
19
1>
1C
b110 G
#263180000000
0!
0*
09
0>
0C
#263190000000
1!
1*
b111 6
19
1>
1C
b111 G
#263200000000
0!
1"
0*
1+
09
1:
0>
0C
#263210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#263220000000
0!
0*
09
0>
0C
#263230000000
1!
1*
b1 6
19
1>
1C
b1 G
#263240000000
0!
0*
09
0>
0C
#263250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#263260000000
0!
0*
09
0>
0C
#263270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#263280000000
0!
0*
09
0>
0C
#263290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#263300000000
0!
0*
09
0>
0C
#263310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#263320000000
0!
0#
0*
0,
09
0>
0?
0C
#263330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#263340000000
0!
0*
09
0>
0C
#263350000000
1!
1*
19
1>
1C
#263360000000
0!
0*
09
0>
0C
#263370000000
1!
1*
19
1>
1C
#263380000000
0!
0*
09
0>
0C
#263390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#263400000000
0!
0*
09
0>
0C
#263410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#263420000000
0!
0*
09
0>
0C
#263430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#263440000000
0!
0*
09
0>
0C
#263450000000
1!
1*
b10 6
19
1>
1C
b10 G
#263460000000
0!
0*
09
0>
0C
#263470000000
1!
1*
b11 6
19
1>
1C
b11 G
#263480000000
0!
0*
09
0>
0C
#263490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#263500000000
0!
0*
09
0>
0C
#263510000000
1!
1*
b101 6
19
1>
1C
b101 G
#263520000000
0!
0*
09
0>
0C
#263530000000
1!
1*
b110 6
19
1>
1C
b110 G
#263540000000
0!
0*
09
0>
0C
#263550000000
1!
1*
b111 6
19
1>
1C
b111 G
#263560000000
0!
0*
09
0>
0C
#263570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#263580000000
0!
0*
09
0>
0C
#263590000000
1!
1*
b1 6
19
1>
1C
b1 G
#263600000000
0!
0*
09
0>
0C
#263610000000
1!
1*
b10 6
19
1>
1C
b10 G
#263620000000
0!
0*
09
0>
0C
#263630000000
1!
1*
b11 6
19
1>
1C
b11 G
#263640000000
0!
0*
09
0>
0C
#263650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#263660000000
0!
0*
09
0>
0C
#263670000000
1!
1*
b101 6
19
1>
1C
b101 G
#263680000000
0!
0*
09
0>
0C
#263690000000
1!
1*
b110 6
19
1>
1C
b110 G
#263700000000
0!
0*
09
0>
0C
#263710000000
1!
1*
b111 6
19
1>
1C
b111 G
#263720000000
0!
0*
09
0>
0C
#263730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#263740000000
0!
0*
09
0>
0C
#263750000000
1!
1*
b1 6
19
1>
1C
b1 G
#263760000000
0!
0*
09
0>
0C
#263770000000
1!
1*
b10 6
19
1>
1C
b10 G
#263780000000
0!
0*
09
0>
0C
#263790000000
1!
1*
b11 6
19
1>
1C
b11 G
#263800000000
0!
0*
09
0>
0C
#263810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#263820000000
0!
0*
09
0>
0C
#263830000000
1!
1*
b101 6
19
1>
1C
b101 G
#263840000000
0!
0*
09
0>
0C
#263850000000
1!
1*
b110 6
19
1>
1C
b110 G
#263860000000
0!
0*
09
0>
0C
#263870000000
1!
1*
b111 6
19
1>
1C
b111 G
#263880000000
0!
1"
0*
1+
09
1:
0>
0C
#263890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#263900000000
0!
0*
09
0>
0C
#263910000000
1!
1*
b1 6
19
1>
1C
b1 G
#263920000000
0!
0*
09
0>
0C
#263930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#263940000000
0!
0*
09
0>
0C
#263950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#263960000000
0!
0*
09
0>
0C
#263970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#263980000000
0!
0*
09
0>
0C
#263990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#264000000000
0!
0#
0*
0,
09
0>
0?
0C
#264010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#264020000000
0!
0*
09
0>
0C
#264030000000
1!
1*
19
1>
1C
#264040000000
0!
0*
09
0>
0C
#264050000000
1!
1*
19
1>
1C
#264060000000
0!
0*
09
0>
0C
#264070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#264080000000
0!
0*
09
0>
0C
#264090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#264100000000
0!
0*
09
0>
0C
#264110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#264120000000
0!
0*
09
0>
0C
#264130000000
1!
1*
b10 6
19
1>
1C
b10 G
#264140000000
0!
0*
09
0>
0C
#264150000000
1!
1*
b11 6
19
1>
1C
b11 G
#264160000000
0!
0*
09
0>
0C
#264170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#264180000000
0!
0*
09
0>
0C
#264190000000
1!
1*
b101 6
19
1>
1C
b101 G
#264200000000
0!
0*
09
0>
0C
#264210000000
1!
1*
b110 6
19
1>
1C
b110 G
#264220000000
0!
0*
09
0>
0C
#264230000000
1!
1*
b111 6
19
1>
1C
b111 G
#264240000000
0!
0*
09
0>
0C
#264250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#264260000000
0!
0*
09
0>
0C
#264270000000
1!
1*
b1 6
19
1>
1C
b1 G
#264280000000
0!
0*
09
0>
0C
#264290000000
1!
1*
b10 6
19
1>
1C
b10 G
#264300000000
0!
0*
09
0>
0C
#264310000000
1!
1*
b11 6
19
1>
1C
b11 G
#264320000000
0!
0*
09
0>
0C
#264330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#264340000000
0!
0*
09
0>
0C
#264350000000
1!
1*
b101 6
19
1>
1C
b101 G
#264360000000
0!
0*
09
0>
0C
#264370000000
1!
1*
b110 6
19
1>
1C
b110 G
#264380000000
0!
0*
09
0>
0C
#264390000000
1!
1*
b111 6
19
1>
1C
b111 G
#264400000000
0!
0*
09
0>
0C
#264410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#264420000000
0!
0*
09
0>
0C
#264430000000
1!
1*
b1 6
19
1>
1C
b1 G
#264440000000
0!
0*
09
0>
0C
#264450000000
1!
1*
b10 6
19
1>
1C
b10 G
#264460000000
0!
0*
09
0>
0C
#264470000000
1!
1*
b11 6
19
1>
1C
b11 G
#264480000000
0!
0*
09
0>
0C
#264490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#264500000000
0!
0*
09
0>
0C
#264510000000
1!
1*
b101 6
19
1>
1C
b101 G
#264520000000
0!
0*
09
0>
0C
#264530000000
1!
1*
b110 6
19
1>
1C
b110 G
#264540000000
0!
0*
09
0>
0C
#264550000000
1!
1*
b111 6
19
1>
1C
b111 G
#264560000000
0!
1"
0*
1+
09
1:
0>
0C
#264570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#264580000000
0!
0*
09
0>
0C
#264590000000
1!
1*
b1 6
19
1>
1C
b1 G
#264600000000
0!
0*
09
0>
0C
#264610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#264620000000
0!
0*
09
0>
0C
#264630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#264640000000
0!
0*
09
0>
0C
#264650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#264660000000
0!
0*
09
0>
0C
#264670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#264680000000
0!
0#
0*
0,
09
0>
0?
0C
#264690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#264700000000
0!
0*
09
0>
0C
#264710000000
1!
1*
19
1>
1C
#264720000000
0!
0*
09
0>
0C
#264730000000
1!
1*
19
1>
1C
#264740000000
0!
0*
09
0>
0C
#264750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#264760000000
0!
0*
09
0>
0C
#264770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#264780000000
0!
0*
09
0>
0C
#264790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#264800000000
0!
0*
09
0>
0C
#264810000000
1!
1*
b10 6
19
1>
1C
b10 G
#264820000000
0!
0*
09
0>
0C
#264830000000
1!
1*
b11 6
19
1>
1C
b11 G
#264840000000
0!
0*
09
0>
0C
#264850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#264860000000
0!
0*
09
0>
0C
#264870000000
1!
1*
b101 6
19
1>
1C
b101 G
#264880000000
0!
0*
09
0>
0C
#264890000000
1!
1*
b110 6
19
1>
1C
b110 G
#264900000000
0!
0*
09
0>
0C
#264910000000
1!
1*
b111 6
19
1>
1C
b111 G
#264920000000
0!
0*
09
0>
0C
#264930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#264940000000
0!
0*
09
0>
0C
#264950000000
1!
1*
b1 6
19
1>
1C
b1 G
#264960000000
0!
0*
09
0>
0C
#264970000000
1!
1*
b10 6
19
1>
1C
b10 G
#264980000000
0!
0*
09
0>
0C
#264990000000
1!
1*
b11 6
19
1>
1C
b11 G
#265000000000
0!
0*
09
0>
0C
#265010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#265020000000
0!
0*
09
0>
0C
#265030000000
1!
1*
b101 6
19
1>
1C
b101 G
#265040000000
0!
0*
09
0>
0C
#265050000000
1!
1*
b110 6
19
1>
1C
b110 G
#265060000000
0!
0*
09
0>
0C
#265070000000
1!
1*
b111 6
19
1>
1C
b111 G
#265080000000
0!
0*
09
0>
0C
#265090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#265100000000
0!
0*
09
0>
0C
#265110000000
1!
1*
b1 6
19
1>
1C
b1 G
#265120000000
0!
0*
09
0>
0C
#265130000000
1!
1*
b10 6
19
1>
1C
b10 G
#265140000000
0!
0*
09
0>
0C
#265150000000
1!
1*
b11 6
19
1>
1C
b11 G
#265160000000
0!
0*
09
0>
0C
#265170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#265180000000
0!
0*
09
0>
0C
#265190000000
1!
1*
b101 6
19
1>
1C
b101 G
#265200000000
0!
0*
09
0>
0C
#265210000000
1!
1*
b110 6
19
1>
1C
b110 G
#265220000000
0!
0*
09
0>
0C
#265230000000
1!
1*
b111 6
19
1>
1C
b111 G
#265240000000
0!
1"
0*
1+
09
1:
0>
0C
#265250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#265260000000
0!
0*
09
0>
0C
#265270000000
1!
1*
b1 6
19
1>
1C
b1 G
#265280000000
0!
0*
09
0>
0C
#265290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#265300000000
0!
0*
09
0>
0C
#265310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#265320000000
0!
0*
09
0>
0C
#265330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#265340000000
0!
0*
09
0>
0C
#265350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#265360000000
0!
0#
0*
0,
09
0>
0?
0C
#265370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#265380000000
0!
0*
09
0>
0C
#265390000000
1!
1*
19
1>
1C
#265400000000
0!
0*
09
0>
0C
#265410000000
1!
1*
19
1>
1C
#265420000000
0!
0*
09
0>
0C
#265430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#265440000000
0!
0*
09
0>
0C
#265450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#265460000000
0!
0*
09
0>
0C
#265470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#265480000000
0!
0*
09
0>
0C
#265490000000
1!
1*
b10 6
19
1>
1C
b10 G
#265500000000
0!
0*
09
0>
0C
#265510000000
1!
1*
b11 6
19
1>
1C
b11 G
#265520000000
0!
0*
09
0>
0C
#265530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#265540000000
0!
0*
09
0>
0C
#265550000000
1!
1*
b101 6
19
1>
1C
b101 G
#265560000000
0!
0*
09
0>
0C
#265570000000
1!
1*
b110 6
19
1>
1C
b110 G
#265580000000
0!
0*
09
0>
0C
#265590000000
1!
1*
b111 6
19
1>
1C
b111 G
#265600000000
0!
0*
09
0>
0C
#265610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#265620000000
0!
0*
09
0>
0C
#265630000000
1!
1*
b1 6
19
1>
1C
b1 G
#265640000000
0!
0*
09
0>
0C
#265650000000
1!
1*
b10 6
19
1>
1C
b10 G
#265660000000
0!
0*
09
0>
0C
#265670000000
1!
1*
b11 6
19
1>
1C
b11 G
#265680000000
0!
0*
09
0>
0C
#265690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#265700000000
0!
0*
09
0>
0C
#265710000000
1!
1*
b101 6
19
1>
1C
b101 G
#265720000000
0!
0*
09
0>
0C
#265730000000
1!
1*
b110 6
19
1>
1C
b110 G
#265740000000
0!
0*
09
0>
0C
#265750000000
1!
1*
b111 6
19
1>
1C
b111 G
#265760000000
0!
0*
09
0>
0C
#265770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#265780000000
0!
0*
09
0>
0C
#265790000000
1!
1*
b1 6
19
1>
1C
b1 G
#265800000000
0!
0*
09
0>
0C
#265810000000
1!
1*
b10 6
19
1>
1C
b10 G
#265820000000
0!
0*
09
0>
0C
#265830000000
1!
1*
b11 6
19
1>
1C
b11 G
#265840000000
0!
0*
09
0>
0C
#265850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#265860000000
0!
0*
09
0>
0C
#265870000000
1!
1*
b101 6
19
1>
1C
b101 G
#265880000000
0!
0*
09
0>
0C
#265890000000
1!
1*
b110 6
19
1>
1C
b110 G
#265900000000
0!
0*
09
0>
0C
#265910000000
1!
1*
b111 6
19
1>
1C
b111 G
#265920000000
0!
1"
0*
1+
09
1:
0>
0C
#265930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#265940000000
0!
0*
09
0>
0C
#265950000000
1!
1*
b1 6
19
1>
1C
b1 G
#265960000000
0!
0*
09
0>
0C
#265970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#265980000000
0!
0*
09
0>
0C
#265990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#266000000000
0!
0*
09
0>
0C
#266010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#266020000000
0!
0*
09
0>
0C
#266030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#266040000000
0!
0#
0*
0,
09
0>
0?
0C
#266050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#266060000000
0!
0*
09
0>
0C
#266070000000
1!
1*
19
1>
1C
#266080000000
0!
0*
09
0>
0C
#266090000000
1!
1*
19
1>
1C
#266100000000
0!
0*
09
0>
0C
#266110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#266120000000
0!
0*
09
0>
0C
#266130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#266140000000
0!
0*
09
0>
0C
#266150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#266160000000
0!
0*
09
0>
0C
#266170000000
1!
1*
b10 6
19
1>
1C
b10 G
#266180000000
0!
0*
09
0>
0C
#266190000000
1!
1*
b11 6
19
1>
1C
b11 G
#266200000000
0!
0*
09
0>
0C
#266210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#266220000000
0!
0*
09
0>
0C
#266230000000
1!
1*
b101 6
19
1>
1C
b101 G
#266240000000
0!
0*
09
0>
0C
#266250000000
1!
1*
b110 6
19
1>
1C
b110 G
#266260000000
0!
0*
09
0>
0C
#266270000000
1!
1*
b111 6
19
1>
1C
b111 G
#266280000000
0!
0*
09
0>
0C
#266290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#266300000000
0!
0*
09
0>
0C
#266310000000
1!
1*
b1 6
19
1>
1C
b1 G
#266320000000
0!
0*
09
0>
0C
#266330000000
1!
1*
b10 6
19
1>
1C
b10 G
#266340000000
0!
0*
09
0>
0C
#266350000000
1!
1*
b11 6
19
1>
1C
b11 G
#266360000000
0!
0*
09
0>
0C
#266370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#266380000000
0!
0*
09
0>
0C
#266390000000
1!
1*
b101 6
19
1>
1C
b101 G
#266400000000
0!
0*
09
0>
0C
#266410000000
1!
1*
b110 6
19
1>
1C
b110 G
#266420000000
0!
0*
09
0>
0C
#266430000000
1!
1*
b111 6
19
1>
1C
b111 G
#266440000000
0!
0*
09
0>
0C
#266450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#266460000000
0!
0*
09
0>
0C
#266470000000
1!
1*
b1 6
19
1>
1C
b1 G
#266480000000
0!
0*
09
0>
0C
#266490000000
1!
1*
b10 6
19
1>
1C
b10 G
#266500000000
0!
0*
09
0>
0C
#266510000000
1!
1*
b11 6
19
1>
1C
b11 G
#266520000000
0!
0*
09
0>
0C
#266530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#266540000000
0!
0*
09
0>
0C
#266550000000
1!
1*
b101 6
19
1>
1C
b101 G
#266560000000
0!
0*
09
0>
0C
#266570000000
1!
1*
b110 6
19
1>
1C
b110 G
#266580000000
0!
0*
09
0>
0C
#266590000000
1!
1*
b111 6
19
1>
1C
b111 G
#266600000000
0!
1"
0*
1+
09
1:
0>
0C
#266610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#266620000000
0!
0*
09
0>
0C
#266630000000
1!
1*
b1 6
19
1>
1C
b1 G
#266640000000
0!
0*
09
0>
0C
#266650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#266660000000
0!
0*
09
0>
0C
#266670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#266680000000
0!
0*
09
0>
0C
#266690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#266700000000
0!
0*
09
0>
0C
#266710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#266720000000
0!
0#
0*
0,
09
0>
0?
0C
#266730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#266740000000
0!
0*
09
0>
0C
#266750000000
1!
1*
19
1>
1C
#266760000000
0!
0*
09
0>
0C
#266770000000
1!
1*
19
1>
1C
#266780000000
0!
0*
09
0>
0C
#266790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#266800000000
0!
0*
09
0>
0C
#266810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#266820000000
0!
0*
09
0>
0C
#266830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#266840000000
0!
0*
09
0>
0C
#266850000000
1!
1*
b10 6
19
1>
1C
b10 G
#266860000000
0!
0*
09
0>
0C
#266870000000
1!
1*
b11 6
19
1>
1C
b11 G
#266880000000
0!
0*
09
0>
0C
#266890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#266900000000
0!
0*
09
0>
0C
#266910000000
1!
1*
b101 6
19
1>
1C
b101 G
#266920000000
0!
0*
09
0>
0C
#266930000000
1!
1*
b110 6
19
1>
1C
b110 G
#266940000000
0!
0*
09
0>
0C
#266950000000
1!
1*
b111 6
19
1>
1C
b111 G
#266960000000
0!
0*
09
0>
0C
#266970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#266980000000
0!
0*
09
0>
0C
#266990000000
1!
1*
b1 6
19
1>
1C
b1 G
#267000000000
0!
0*
09
0>
0C
#267010000000
1!
1*
b10 6
19
1>
1C
b10 G
#267020000000
0!
0*
09
0>
0C
#267030000000
1!
1*
b11 6
19
1>
1C
b11 G
#267040000000
0!
0*
09
0>
0C
#267050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#267060000000
0!
0*
09
0>
0C
#267070000000
1!
1*
b101 6
19
1>
1C
b101 G
#267080000000
0!
0*
09
0>
0C
#267090000000
1!
1*
b110 6
19
1>
1C
b110 G
#267100000000
0!
0*
09
0>
0C
#267110000000
1!
1*
b111 6
19
1>
1C
b111 G
#267120000000
0!
0*
09
0>
0C
#267130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#267140000000
0!
0*
09
0>
0C
#267150000000
1!
1*
b1 6
19
1>
1C
b1 G
#267160000000
0!
0*
09
0>
0C
#267170000000
1!
1*
b10 6
19
1>
1C
b10 G
#267180000000
0!
0*
09
0>
0C
#267190000000
1!
1*
b11 6
19
1>
1C
b11 G
#267200000000
0!
0*
09
0>
0C
#267210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#267220000000
0!
0*
09
0>
0C
#267230000000
1!
1*
b101 6
19
1>
1C
b101 G
#267240000000
0!
0*
09
0>
0C
#267250000000
1!
1*
b110 6
19
1>
1C
b110 G
#267260000000
0!
0*
09
0>
0C
#267270000000
1!
1*
b111 6
19
1>
1C
b111 G
#267280000000
0!
1"
0*
1+
09
1:
0>
0C
#267290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#267300000000
0!
0*
09
0>
0C
#267310000000
1!
1*
b1 6
19
1>
1C
b1 G
#267320000000
0!
0*
09
0>
0C
#267330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#267340000000
0!
0*
09
0>
0C
#267350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#267360000000
0!
0*
09
0>
0C
#267370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#267380000000
0!
0*
09
0>
0C
#267390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#267400000000
0!
0#
0*
0,
09
0>
0?
0C
#267410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#267420000000
0!
0*
09
0>
0C
#267430000000
1!
1*
19
1>
1C
#267440000000
0!
0*
09
0>
0C
#267450000000
1!
1*
19
1>
1C
#267460000000
0!
0*
09
0>
0C
#267470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#267480000000
0!
0*
09
0>
0C
#267490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#267500000000
0!
0*
09
0>
0C
#267510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#267520000000
0!
0*
09
0>
0C
#267530000000
1!
1*
b10 6
19
1>
1C
b10 G
#267540000000
0!
0*
09
0>
0C
#267550000000
1!
1*
b11 6
19
1>
1C
b11 G
#267560000000
0!
0*
09
0>
0C
#267570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#267580000000
0!
0*
09
0>
0C
#267590000000
1!
1*
b101 6
19
1>
1C
b101 G
#267600000000
0!
0*
09
0>
0C
#267610000000
1!
1*
b110 6
19
1>
1C
b110 G
#267620000000
0!
0*
09
0>
0C
#267630000000
1!
1*
b111 6
19
1>
1C
b111 G
#267640000000
0!
0*
09
0>
0C
#267650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#267660000000
0!
0*
09
0>
0C
#267670000000
1!
1*
b1 6
19
1>
1C
b1 G
#267680000000
0!
0*
09
0>
0C
#267690000000
1!
1*
b10 6
19
1>
1C
b10 G
#267700000000
0!
0*
09
0>
0C
#267710000000
1!
1*
b11 6
19
1>
1C
b11 G
#267720000000
0!
0*
09
0>
0C
#267730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#267740000000
0!
0*
09
0>
0C
#267750000000
1!
1*
b101 6
19
1>
1C
b101 G
#267760000000
0!
0*
09
0>
0C
#267770000000
1!
1*
b110 6
19
1>
1C
b110 G
#267780000000
0!
0*
09
0>
0C
#267790000000
1!
1*
b111 6
19
1>
1C
b111 G
#267800000000
0!
0*
09
0>
0C
#267810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#267820000000
0!
0*
09
0>
0C
#267830000000
1!
1*
b1 6
19
1>
1C
b1 G
#267840000000
0!
0*
09
0>
0C
#267850000000
1!
1*
b10 6
19
1>
1C
b10 G
#267860000000
0!
0*
09
0>
0C
#267870000000
1!
1*
b11 6
19
1>
1C
b11 G
#267880000000
0!
0*
09
0>
0C
#267890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#267900000000
0!
0*
09
0>
0C
#267910000000
1!
1*
b101 6
19
1>
1C
b101 G
#267920000000
0!
0*
09
0>
0C
#267930000000
1!
1*
b110 6
19
1>
1C
b110 G
#267940000000
0!
0*
09
0>
0C
#267950000000
1!
1*
b111 6
19
1>
1C
b111 G
#267960000000
0!
1"
0*
1+
09
1:
0>
0C
#267970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#267980000000
0!
0*
09
0>
0C
#267990000000
1!
1*
b1 6
19
1>
1C
b1 G
#268000000000
0!
0*
09
0>
0C
#268010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#268020000000
0!
0*
09
0>
0C
#268030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#268040000000
0!
0*
09
0>
0C
#268050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#268060000000
0!
0*
09
0>
0C
#268070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#268080000000
0!
0#
0*
0,
09
0>
0?
0C
#268090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#268100000000
0!
0*
09
0>
0C
#268110000000
1!
1*
19
1>
1C
#268120000000
0!
0*
09
0>
0C
#268130000000
1!
1*
19
1>
1C
#268140000000
0!
0*
09
0>
0C
#268150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#268160000000
0!
0*
09
0>
0C
#268170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#268180000000
0!
0*
09
0>
0C
#268190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#268200000000
0!
0*
09
0>
0C
#268210000000
1!
1*
b10 6
19
1>
1C
b10 G
#268220000000
0!
0*
09
0>
0C
#268230000000
1!
1*
b11 6
19
1>
1C
b11 G
#268240000000
0!
0*
09
0>
0C
#268250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#268260000000
0!
0*
09
0>
0C
#268270000000
1!
1*
b101 6
19
1>
1C
b101 G
#268280000000
0!
0*
09
0>
0C
#268290000000
1!
1*
b110 6
19
1>
1C
b110 G
#268300000000
0!
0*
09
0>
0C
#268310000000
1!
1*
b111 6
19
1>
1C
b111 G
#268320000000
0!
0*
09
0>
0C
#268330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#268340000000
0!
0*
09
0>
0C
#268350000000
1!
1*
b1 6
19
1>
1C
b1 G
#268360000000
0!
0*
09
0>
0C
#268370000000
1!
1*
b10 6
19
1>
1C
b10 G
#268380000000
0!
0*
09
0>
0C
#268390000000
1!
1*
b11 6
19
1>
1C
b11 G
#268400000000
0!
0*
09
0>
0C
#268410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#268420000000
0!
0*
09
0>
0C
#268430000000
1!
1*
b101 6
19
1>
1C
b101 G
#268440000000
0!
0*
09
0>
0C
#268450000000
1!
1*
b110 6
19
1>
1C
b110 G
#268460000000
0!
0*
09
0>
0C
#268470000000
1!
1*
b111 6
19
1>
1C
b111 G
#268480000000
0!
0*
09
0>
0C
#268490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#268500000000
0!
0*
09
0>
0C
#268510000000
1!
1*
b1 6
19
1>
1C
b1 G
#268520000000
0!
0*
09
0>
0C
#268530000000
1!
1*
b10 6
19
1>
1C
b10 G
#268540000000
0!
0*
09
0>
0C
#268550000000
1!
1*
b11 6
19
1>
1C
b11 G
#268560000000
0!
0*
09
0>
0C
#268570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#268580000000
0!
0*
09
0>
0C
#268590000000
1!
1*
b101 6
19
1>
1C
b101 G
#268600000000
0!
0*
09
0>
0C
#268610000000
1!
1*
b110 6
19
1>
1C
b110 G
#268620000000
0!
0*
09
0>
0C
#268630000000
1!
1*
b111 6
19
1>
1C
b111 G
#268640000000
0!
1"
0*
1+
09
1:
0>
0C
#268650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#268660000000
0!
0*
09
0>
0C
#268670000000
1!
1*
b1 6
19
1>
1C
b1 G
#268680000000
0!
0*
09
0>
0C
#268690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#268700000000
0!
0*
09
0>
0C
#268710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#268720000000
0!
0*
09
0>
0C
#268730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#268740000000
0!
0*
09
0>
0C
#268750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#268760000000
0!
0#
0*
0,
09
0>
0?
0C
#268770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#268780000000
0!
0*
09
0>
0C
#268790000000
1!
1*
19
1>
1C
#268800000000
0!
0*
09
0>
0C
#268810000000
1!
1*
19
1>
1C
#268820000000
0!
0*
09
0>
0C
#268830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#268840000000
0!
0*
09
0>
0C
#268850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#268860000000
0!
0*
09
0>
0C
#268870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#268880000000
0!
0*
09
0>
0C
#268890000000
1!
1*
b10 6
19
1>
1C
b10 G
#268900000000
0!
0*
09
0>
0C
#268910000000
1!
1*
b11 6
19
1>
1C
b11 G
#268920000000
0!
0*
09
0>
0C
#268930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#268940000000
0!
0*
09
0>
0C
#268950000000
1!
1*
b101 6
19
1>
1C
b101 G
#268960000000
0!
0*
09
0>
0C
#268970000000
1!
1*
b110 6
19
1>
1C
b110 G
#268980000000
0!
0*
09
0>
0C
#268990000000
1!
1*
b111 6
19
1>
1C
b111 G
#269000000000
0!
0*
09
0>
0C
#269010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#269020000000
0!
0*
09
0>
0C
#269030000000
1!
1*
b1 6
19
1>
1C
b1 G
#269040000000
0!
0*
09
0>
0C
#269050000000
1!
1*
b10 6
19
1>
1C
b10 G
#269060000000
0!
0*
09
0>
0C
#269070000000
1!
1*
b11 6
19
1>
1C
b11 G
#269080000000
0!
0*
09
0>
0C
#269090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#269100000000
0!
0*
09
0>
0C
#269110000000
1!
1*
b101 6
19
1>
1C
b101 G
#269120000000
0!
0*
09
0>
0C
#269130000000
1!
1*
b110 6
19
1>
1C
b110 G
#269140000000
0!
0*
09
0>
0C
#269150000000
1!
1*
b111 6
19
1>
1C
b111 G
#269160000000
0!
0*
09
0>
0C
#269170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#269180000000
0!
0*
09
0>
0C
#269190000000
1!
1*
b1 6
19
1>
1C
b1 G
#269200000000
0!
0*
09
0>
0C
#269210000000
1!
1*
b10 6
19
1>
1C
b10 G
#269220000000
0!
0*
09
0>
0C
#269230000000
1!
1*
b11 6
19
1>
1C
b11 G
#269240000000
0!
0*
09
0>
0C
#269250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#269260000000
0!
0*
09
0>
0C
#269270000000
1!
1*
b101 6
19
1>
1C
b101 G
#269280000000
0!
0*
09
0>
0C
#269290000000
1!
1*
b110 6
19
1>
1C
b110 G
#269300000000
0!
0*
09
0>
0C
#269310000000
1!
1*
b111 6
19
1>
1C
b111 G
#269320000000
0!
1"
0*
1+
09
1:
0>
0C
#269330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#269340000000
0!
0*
09
0>
0C
#269350000000
1!
1*
b1 6
19
1>
1C
b1 G
#269360000000
0!
0*
09
0>
0C
#269370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#269380000000
0!
0*
09
0>
0C
#269390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#269400000000
0!
0*
09
0>
0C
#269410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#269420000000
0!
0*
09
0>
0C
#269430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#269440000000
0!
0#
0*
0,
09
0>
0?
0C
#269450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#269460000000
0!
0*
09
0>
0C
#269470000000
1!
1*
19
1>
1C
#269480000000
0!
0*
09
0>
0C
#269490000000
1!
1*
19
1>
1C
#269500000000
0!
0*
09
0>
0C
#269510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#269520000000
0!
0*
09
0>
0C
#269530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#269540000000
0!
0*
09
0>
0C
#269550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#269560000000
0!
0*
09
0>
0C
#269570000000
1!
1*
b10 6
19
1>
1C
b10 G
#269580000000
0!
0*
09
0>
0C
#269590000000
1!
1*
b11 6
19
1>
1C
b11 G
#269600000000
0!
0*
09
0>
0C
#269610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#269620000000
0!
0*
09
0>
0C
#269630000000
1!
1*
b101 6
19
1>
1C
b101 G
#269640000000
0!
0*
09
0>
0C
#269650000000
1!
1*
b110 6
19
1>
1C
b110 G
#269660000000
0!
0*
09
0>
0C
#269670000000
1!
1*
b111 6
19
1>
1C
b111 G
#269680000000
0!
0*
09
0>
0C
#269690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#269700000000
0!
0*
09
0>
0C
#269710000000
1!
1*
b1 6
19
1>
1C
b1 G
#269720000000
0!
0*
09
0>
0C
#269730000000
1!
1*
b10 6
19
1>
1C
b10 G
#269740000000
0!
0*
09
0>
0C
#269750000000
1!
1*
b11 6
19
1>
1C
b11 G
#269760000000
0!
0*
09
0>
0C
#269770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#269780000000
0!
0*
09
0>
0C
#269790000000
1!
1*
b101 6
19
1>
1C
b101 G
#269800000000
0!
0*
09
0>
0C
#269810000000
1!
1*
b110 6
19
1>
1C
b110 G
#269820000000
0!
0*
09
0>
0C
#269830000000
1!
1*
b111 6
19
1>
1C
b111 G
#269840000000
0!
0*
09
0>
0C
#269850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#269860000000
0!
0*
09
0>
0C
#269870000000
1!
1*
b1 6
19
1>
1C
b1 G
#269880000000
0!
0*
09
0>
0C
#269890000000
1!
1*
b10 6
19
1>
1C
b10 G
#269900000000
0!
0*
09
0>
0C
#269910000000
1!
1*
b11 6
19
1>
1C
b11 G
#269920000000
0!
0*
09
0>
0C
#269930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#269940000000
0!
0*
09
0>
0C
#269950000000
1!
1*
b101 6
19
1>
1C
b101 G
#269960000000
0!
0*
09
0>
0C
#269970000000
1!
1*
b110 6
19
1>
1C
b110 G
#269980000000
0!
0*
09
0>
0C
#269990000000
1!
1*
b111 6
19
1>
1C
b111 G
#270000000000
0!
1"
0*
1+
09
1:
0>
0C
#270010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#270020000000
0!
0*
09
0>
0C
#270030000000
1!
1*
b1 6
19
1>
1C
b1 G
#270040000000
0!
0*
09
0>
0C
#270050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#270060000000
0!
0*
09
0>
0C
#270070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#270080000000
0!
0*
09
0>
0C
#270090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#270100000000
0!
0*
09
0>
0C
#270110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#270120000000
0!
0#
0*
0,
09
0>
0?
0C
#270130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#270140000000
0!
0*
09
0>
0C
#270150000000
1!
1*
19
1>
1C
#270160000000
0!
0*
09
0>
0C
#270170000000
1!
1*
19
1>
1C
#270180000000
0!
0*
09
0>
0C
#270190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#270200000000
0!
0*
09
0>
0C
#270210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#270220000000
0!
0*
09
0>
0C
#270230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#270240000000
0!
0*
09
0>
0C
#270250000000
1!
1*
b10 6
19
1>
1C
b10 G
#270260000000
0!
0*
09
0>
0C
#270270000000
1!
1*
b11 6
19
1>
1C
b11 G
#270280000000
0!
0*
09
0>
0C
#270290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#270300000000
0!
0*
09
0>
0C
#270310000000
1!
1*
b101 6
19
1>
1C
b101 G
#270320000000
0!
0*
09
0>
0C
#270330000000
1!
1*
b110 6
19
1>
1C
b110 G
#270340000000
0!
0*
09
0>
0C
#270350000000
1!
1*
b111 6
19
1>
1C
b111 G
#270360000000
0!
0*
09
0>
0C
#270370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#270380000000
0!
0*
09
0>
0C
#270390000000
1!
1*
b1 6
19
1>
1C
b1 G
#270400000000
0!
0*
09
0>
0C
#270410000000
1!
1*
b10 6
19
1>
1C
b10 G
#270420000000
0!
0*
09
0>
0C
#270430000000
1!
1*
b11 6
19
1>
1C
b11 G
#270440000000
0!
0*
09
0>
0C
#270450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#270460000000
0!
0*
09
0>
0C
#270470000000
1!
1*
b101 6
19
1>
1C
b101 G
#270480000000
0!
0*
09
0>
0C
#270490000000
1!
1*
b110 6
19
1>
1C
b110 G
#270500000000
0!
0*
09
0>
0C
#270510000000
1!
1*
b111 6
19
1>
1C
b111 G
#270520000000
0!
0*
09
0>
0C
#270530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#270540000000
0!
0*
09
0>
0C
#270550000000
1!
1*
b1 6
19
1>
1C
b1 G
#270560000000
0!
0*
09
0>
0C
#270570000000
1!
1*
b10 6
19
1>
1C
b10 G
#270580000000
0!
0*
09
0>
0C
#270590000000
1!
1*
b11 6
19
1>
1C
b11 G
#270600000000
0!
0*
09
0>
0C
#270610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#270620000000
0!
0*
09
0>
0C
#270630000000
1!
1*
b101 6
19
1>
1C
b101 G
#270640000000
0!
0*
09
0>
0C
#270650000000
1!
1*
b110 6
19
1>
1C
b110 G
#270660000000
0!
0*
09
0>
0C
#270670000000
1!
1*
b111 6
19
1>
1C
b111 G
#270680000000
0!
1"
0*
1+
09
1:
0>
0C
#270690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#270700000000
0!
0*
09
0>
0C
#270710000000
1!
1*
b1 6
19
1>
1C
b1 G
#270720000000
0!
0*
09
0>
0C
#270730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#270740000000
0!
0*
09
0>
0C
#270750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#270760000000
0!
0*
09
0>
0C
#270770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#270780000000
0!
0*
09
0>
0C
#270790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#270800000000
0!
0#
0*
0,
09
0>
0?
0C
#270810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#270820000000
0!
0*
09
0>
0C
#270830000000
1!
1*
19
1>
1C
#270840000000
0!
0*
09
0>
0C
#270850000000
1!
1*
19
1>
1C
#270860000000
0!
0*
09
0>
0C
#270870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#270880000000
0!
0*
09
0>
0C
#270890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#270900000000
0!
0*
09
0>
0C
#270910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#270920000000
0!
0*
09
0>
0C
#270930000000
1!
1*
b10 6
19
1>
1C
b10 G
#270940000000
0!
0*
09
0>
0C
#270950000000
1!
1*
b11 6
19
1>
1C
b11 G
#270960000000
0!
0*
09
0>
0C
#270970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#270980000000
0!
0*
09
0>
0C
#270990000000
1!
1*
b101 6
19
1>
1C
b101 G
#271000000000
0!
0*
09
0>
0C
#271010000000
1!
1*
b110 6
19
1>
1C
b110 G
#271020000000
0!
0*
09
0>
0C
#271030000000
1!
1*
b111 6
19
1>
1C
b111 G
#271040000000
0!
0*
09
0>
0C
#271050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#271060000000
0!
0*
09
0>
0C
#271070000000
1!
1*
b1 6
19
1>
1C
b1 G
#271080000000
0!
0*
09
0>
0C
#271090000000
1!
1*
b10 6
19
1>
1C
b10 G
#271100000000
0!
0*
09
0>
0C
#271110000000
1!
1*
b11 6
19
1>
1C
b11 G
#271120000000
0!
0*
09
0>
0C
#271130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#271140000000
0!
0*
09
0>
0C
#271150000000
1!
1*
b101 6
19
1>
1C
b101 G
#271160000000
0!
0*
09
0>
0C
#271170000000
1!
1*
b110 6
19
1>
1C
b110 G
#271180000000
0!
0*
09
0>
0C
#271190000000
1!
1*
b111 6
19
1>
1C
b111 G
#271200000000
0!
0*
09
0>
0C
#271210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#271220000000
0!
0*
09
0>
0C
#271230000000
1!
1*
b1 6
19
1>
1C
b1 G
#271240000000
0!
0*
09
0>
0C
#271250000000
1!
1*
b10 6
19
1>
1C
b10 G
#271260000000
0!
0*
09
0>
0C
#271270000000
1!
1*
b11 6
19
1>
1C
b11 G
#271280000000
0!
0*
09
0>
0C
#271290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#271300000000
0!
0*
09
0>
0C
#271310000000
1!
1*
b101 6
19
1>
1C
b101 G
#271320000000
0!
0*
09
0>
0C
#271330000000
1!
1*
b110 6
19
1>
1C
b110 G
#271340000000
0!
0*
09
0>
0C
#271350000000
1!
1*
b111 6
19
1>
1C
b111 G
#271360000000
0!
1"
0*
1+
09
1:
0>
0C
#271370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#271380000000
0!
0*
09
0>
0C
#271390000000
1!
1*
b1 6
19
1>
1C
b1 G
#271400000000
0!
0*
09
0>
0C
#271410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#271420000000
0!
0*
09
0>
0C
#271430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#271440000000
0!
0*
09
0>
0C
#271450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#271460000000
0!
0*
09
0>
0C
#271470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#271480000000
0!
0#
0*
0,
09
0>
0?
0C
#271490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#271500000000
0!
0*
09
0>
0C
#271510000000
1!
1*
19
1>
1C
#271520000000
0!
0*
09
0>
0C
#271530000000
1!
1*
19
1>
1C
#271540000000
0!
0*
09
0>
0C
#271550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#271560000000
0!
0*
09
0>
0C
#271570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#271580000000
0!
0*
09
0>
0C
#271590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#271600000000
0!
0*
09
0>
0C
#271610000000
1!
1*
b10 6
19
1>
1C
b10 G
#271620000000
0!
0*
09
0>
0C
#271630000000
1!
1*
b11 6
19
1>
1C
b11 G
#271640000000
0!
0*
09
0>
0C
#271650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#271660000000
0!
0*
09
0>
0C
#271670000000
1!
1*
b101 6
19
1>
1C
b101 G
#271680000000
0!
0*
09
0>
0C
#271690000000
1!
1*
b110 6
19
1>
1C
b110 G
#271700000000
0!
0*
09
0>
0C
#271710000000
1!
1*
b111 6
19
1>
1C
b111 G
#271720000000
0!
0*
09
0>
0C
#271730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#271740000000
0!
0*
09
0>
0C
#271750000000
1!
1*
b1 6
19
1>
1C
b1 G
#271760000000
0!
0*
09
0>
0C
#271770000000
1!
1*
b10 6
19
1>
1C
b10 G
#271780000000
0!
0*
09
0>
0C
#271790000000
1!
1*
b11 6
19
1>
1C
b11 G
#271800000000
0!
0*
09
0>
0C
#271810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#271820000000
0!
0*
09
0>
0C
#271830000000
1!
1*
b101 6
19
1>
1C
b101 G
#271840000000
0!
0*
09
0>
0C
#271850000000
1!
1*
b110 6
19
1>
1C
b110 G
#271860000000
0!
0*
09
0>
0C
#271870000000
1!
1*
b111 6
19
1>
1C
b111 G
#271880000000
0!
0*
09
0>
0C
#271890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#271900000000
0!
0*
09
0>
0C
#271910000000
1!
1*
b1 6
19
1>
1C
b1 G
#271920000000
0!
0*
09
0>
0C
#271930000000
1!
1*
b10 6
19
1>
1C
b10 G
#271940000000
0!
0*
09
0>
0C
#271950000000
1!
1*
b11 6
19
1>
1C
b11 G
#271960000000
0!
0*
09
0>
0C
#271970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#271980000000
0!
0*
09
0>
0C
#271990000000
1!
1*
b101 6
19
1>
1C
b101 G
#272000000000
0!
0*
09
0>
0C
#272010000000
1!
1*
b110 6
19
1>
1C
b110 G
#272020000000
0!
0*
09
0>
0C
#272030000000
1!
1*
b111 6
19
1>
1C
b111 G
#272040000000
0!
1"
0*
1+
09
1:
0>
0C
#272050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#272060000000
0!
0*
09
0>
0C
#272070000000
1!
1*
b1 6
19
1>
1C
b1 G
#272080000000
0!
0*
09
0>
0C
#272090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#272100000000
0!
0*
09
0>
0C
#272110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#272120000000
0!
0*
09
0>
0C
#272130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#272140000000
0!
0*
09
0>
0C
#272150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#272160000000
0!
0#
0*
0,
09
0>
0?
0C
#272170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#272180000000
0!
0*
09
0>
0C
#272190000000
1!
1*
19
1>
1C
#272200000000
0!
0*
09
0>
0C
#272210000000
1!
1*
19
1>
1C
#272220000000
0!
0*
09
0>
0C
#272230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#272240000000
0!
0*
09
0>
0C
#272250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#272260000000
0!
0*
09
0>
0C
#272270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#272280000000
0!
0*
09
0>
0C
#272290000000
1!
1*
b10 6
19
1>
1C
b10 G
#272300000000
0!
0*
09
0>
0C
#272310000000
1!
1*
b11 6
19
1>
1C
b11 G
#272320000000
0!
0*
09
0>
0C
#272330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#272340000000
0!
0*
09
0>
0C
#272350000000
1!
1*
b101 6
19
1>
1C
b101 G
#272360000000
0!
0*
09
0>
0C
#272370000000
1!
1*
b110 6
19
1>
1C
b110 G
#272380000000
0!
0*
09
0>
0C
#272390000000
1!
1*
b111 6
19
1>
1C
b111 G
#272400000000
0!
0*
09
0>
0C
#272410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#272420000000
0!
0*
09
0>
0C
#272430000000
1!
1*
b1 6
19
1>
1C
b1 G
#272440000000
0!
0*
09
0>
0C
#272450000000
1!
1*
b10 6
19
1>
1C
b10 G
#272460000000
0!
0*
09
0>
0C
#272470000000
1!
1*
b11 6
19
1>
1C
b11 G
#272480000000
0!
0*
09
0>
0C
#272490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#272500000000
0!
0*
09
0>
0C
#272510000000
1!
1*
b101 6
19
1>
1C
b101 G
#272520000000
0!
0*
09
0>
0C
#272530000000
1!
1*
b110 6
19
1>
1C
b110 G
#272540000000
0!
0*
09
0>
0C
#272550000000
1!
1*
b111 6
19
1>
1C
b111 G
#272560000000
0!
0*
09
0>
0C
#272570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#272580000000
0!
0*
09
0>
0C
#272590000000
1!
1*
b1 6
19
1>
1C
b1 G
#272600000000
0!
0*
09
0>
0C
#272610000000
1!
1*
b10 6
19
1>
1C
b10 G
#272620000000
0!
0*
09
0>
0C
#272630000000
1!
1*
b11 6
19
1>
1C
b11 G
#272640000000
0!
0*
09
0>
0C
#272650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#272660000000
0!
0*
09
0>
0C
#272670000000
1!
1*
b101 6
19
1>
1C
b101 G
#272680000000
0!
0*
09
0>
0C
#272690000000
1!
1*
b110 6
19
1>
1C
b110 G
#272700000000
0!
0*
09
0>
0C
#272710000000
1!
1*
b111 6
19
1>
1C
b111 G
#272720000000
0!
1"
0*
1+
09
1:
0>
0C
#272730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#272740000000
0!
0*
09
0>
0C
#272750000000
1!
1*
b1 6
19
1>
1C
b1 G
#272760000000
0!
0*
09
0>
0C
#272770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#272780000000
0!
0*
09
0>
0C
#272790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#272800000000
0!
0*
09
0>
0C
#272810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#272820000000
0!
0*
09
0>
0C
#272830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#272840000000
0!
0#
0*
0,
09
0>
0?
0C
#272850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#272860000000
0!
0*
09
0>
0C
#272870000000
1!
1*
19
1>
1C
#272880000000
0!
0*
09
0>
0C
#272890000000
1!
1*
19
1>
1C
#272900000000
0!
0*
09
0>
0C
#272910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#272920000000
0!
0*
09
0>
0C
#272930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#272940000000
0!
0*
09
0>
0C
#272950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#272960000000
0!
0*
09
0>
0C
#272970000000
1!
1*
b10 6
19
1>
1C
b10 G
#272980000000
0!
0*
09
0>
0C
#272990000000
1!
1*
b11 6
19
1>
1C
b11 G
#273000000000
0!
0*
09
0>
0C
#273010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#273020000000
0!
0*
09
0>
0C
#273030000000
1!
1*
b101 6
19
1>
1C
b101 G
#273040000000
0!
0*
09
0>
0C
#273050000000
1!
1*
b110 6
19
1>
1C
b110 G
#273060000000
0!
0*
09
0>
0C
#273070000000
1!
1*
b111 6
19
1>
1C
b111 G
#273080000000
0!
0*
09
0>
0C
#273090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#273100000000
0!
0*
09
0>
0C
#273110000000
1!
1*
b1 6
19
1>
1C
b1 G
#273120000000
0!
0*
09
0>
0C
#273130000000
1!
1*
b10 6
19
1>
1C
b10 G
#273140000000
0!
0*
09
0>
0C
#273150000000
1!
1*
b11 6
19
1>
1C
b11 G
#273160000000
0!
0*
09
0>
0C
#273170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#273180000000
0!
0*
09
0>
0C
#273190000000
1!
1*
b101 6
19
1>
1C
b101 G
#273200000000
0!
0*
09
0>
0C
#273210000000
1!
1*
b110 6
19
1>
1C
b110 G
#273220000000
0!
0*
09
0>
0C
#273230000000
1!
1*
b111 6
19
1>
1C
b111 G
#273240000000
0!
0*
09
0>
0C
#273250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#273260000000
0!
0*
09
0>
0C
#273270000000
1!
1*
b1 6
19
1>
1C
b1 G
#273280000000
0!
0*
09
0>
0C
#273290000000
1!
1*
b10 6
19
1>
1C
b10 G
#273300000000
0!
0*
09
0>
0C
#273310000000
1!
1*
b11 6
19
1>
1C
b11 G
#273320000000
0!
0*
09
0>
0C
#273330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#273340000000
0!
0*
09
0>
0C
#273350000000
1!
1*
b101 6
19
1>
1C
b101 G
#273360000000
0!
0*
09
0>
0C
#273370000000
1!
1*
b110 6
19
1>
1C
b110 G
#273380000000
0!
0*
09
0>
0C
#273390000000
1!
1*
b111 6
19
1>
1C
b111 G
#273400000000
0!
1"
0*
1+
09
1:
0>
0C
#273410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#273420000000
0!
0*
09
0>
0C
#273430000000
1!
1*
b1 6
19
1>
1C
b1 G
#273440000000
0!
0*
09
0>
0C
#273450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#273460000000
0!
0*
09
0>
0C
#273470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#273480000000
0!
0*
09
0>
0C
#273490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#273500000000
0!
0*
09
0>
0C
#273510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#273520000000
0!
0#
0*
0,
09
0>
0?
0C
#273530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#273540000000
0!
0*
09
0>
0C
#273550000000
1!
1*
19
1>
1C
#273560000000
0!
0*
09
0>
0C
#273570000000
1!
1*
19
1>
1C
#273580000000
0!
0*
09
0>
0C
#273590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#273600000000
0!
0*
09
0>
0C
#273610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#273620000000
0!
0*
09
0>
0C
#273630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#273640000000
0!
0*
09
0>
0C
#273650000000
1!
1*
b10 6
19
1>
1C
b10 G
#273660000000
0!
0*
09
0>
0C
#273670000000
1!
1*
b11 6
19
1>
1C
b11 G
#273680000000
0!
0*
09
0>
0C
#273690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#273700000000
0!
0*
09
0>
0C
#273710000000
1!
1*
b101 6
19
1>
1C
b101 G
#273720000000
0!
0*
09
0>
0C
#273730000000
1!
1*
b110 6
19
1>
1C
b110 G
#273740000000
0!
0*
09
0>
0C
#273750000000
1!
1*
b111 6
19
1>
1C
b111 G
#273760000000
0!
0*
09
0>
0C
#273770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#273780000000
0!
0*
09
0>
0C
#273790000000
1!
1*
b1 6
19
1>
1C
b1 G
#273800000000
0!
0*
09
0>
0C
#273810000000
1!
1*
b10 6
19
1>
1C
b10 G
#273820000000
0!
0*
09
0>
0C
#273830000000
1!
1*
b11 6
19
1>
1C
b11 G
#273840000000
0!
0*
09
0>
0C
#273850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#273860000000
0!
0*
09
0>
0C
#273870000000
1!
1*
b101 6
19
1>
1C
b101 G
#273880000000
0!
0*
09
0>
0C
#273890000000
1!
1*
b110 6
19
1>
1C
b110 G
#273900000000
0!
0*
09
0>
0C
#273910000000
1!
1*
b111 6
19
1>
1C
b111 G
#273920000000
0!
0*
09
0>
0C
#273930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#273940000000
0!
0*
09
0>
0C
#273950000000
1!
1*
b1 6
19
1>
1C
b1 G
#273960000000
0!
0*
09
0>
0C
#273970000000
1!
1*
b10 6
19
1>
1C
b10 G
#273980000000
0!
0*
09
0>
0C
#273990000000
1!
1*
b11 6
19
1>
1C
b11 G
#274000000000
0!
0*
09
0>
0C
#274010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#274020000000
0!
0*
09
0>
0C
#274030000000
1!
1*
b101 6
19
1>
1C
b101 G
#274040000000
0!
0*
09
0>
0C
#274050000000
1!
1*
b110 6
19
1>
1C
b110 G
#274060000000
0!
0*
09
0>
0C
#274070000000
1!
1*
b111 6
19
1>
1C
b111 G
#274080000000
0!
1"
0*
1+
09
1:
0>
0C
#274090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#274100000000
0!
0*
09
0>
0C
#274110000000
1!
1*
b1 6
19
1>
1C
b1 G
#274120000000
0!
0*
09
0>
0C
#274130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#274140000000
0!
0*
09
0>
0C
#274150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#274160000000
0!
0*
09
0>
0C
#274170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#274180000000
0!
0*
09
0>
0C
#274190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#274200000000
0!
0#
0*
0,
09
0>
0?
0C
#274210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#274220000000
0!
0*
09
0>
0C
#274230000000
1!
1*
19
1>
1C
#274240000000
0!
0*
09
0>
0C
#274250000000
1!
1*
19
1>
1C
#274260000000
0!
0*
09
0>
0C
#274270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#274280000000
0!
0*
09
0>
0C
#274290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#274300000000
0!
0*
09
0>
0C
#274310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#274320000000
0!
0*
09
0>
0C
#274330000000
1!
1*
b10 6
19
1>
1C
b10 G
#274340000000
0!
0*
09
0>
0C
#274350000000
1!
1*
b11 6
19
1>
1C
b11 G
#274360000000
0!
0*
09
0>
0C
#274370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#274380000000
0!
0*
09
0>
0C
#274390000000
1!
1*
b101 6
19
1>
1C
b101 G
#274400000000
0!
0*
09
0>
0C
#274410000000
1!
1*
b110 6
19
1>
1C
b110 G
#274420000000
0!
0*
09
0>
0C
#274430000000
1!
1*
b111 6
19
1>
1C
b111 G
#274440000000
0!
0*
09
0>
0C
#274450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#274460000000
0!
0*
09
0>
0C
#274470000000
1!
1*
b1 6
19
1>
1C
b1 G
#274480000000
0!
0*
09
0>
0C
#274490000000
1!
1*
b10 6
19
1>
1C
b10 G
#274500000000
0!
0*
09
0>
0C
#274510000000
1!
1*
b11 6
19
1>
1C
b11 G
#274520000000
0!
0*
09
0>
0C
#274530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#274540000000
0!
0*
09
0>
0C
#274550000000
1!
1*
b101 6
19
1>
1C
b101 G
#274560000000
0!
0*
09
0>
0C
#274570000000
1!
1*
b110 6
19
1>
1C
b110 G
#274580000000
0!
0*
09
0>
0C
#274590000000
1!
1*
b111 6
19
1>
1C
b111 G
#274600000000
0!
0*
09
0>
0C
#274610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#274620000000
0!
0*
09
0>
0C
#274630000000
1!
1*
b1 6
19
1>
1C
b1 G
#274640000000
0!
0*
09
0>
0C
#274650000000
1!
1*
b10 6
19
1>
1C
b10 G
#274660000000
0!
0*
09
0>
0C
#274670000000
1!
1*
b11 6
19
1>
1C
b11 G
#274680000000
0!
0*
09
0>
0C
#274690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#274700000000
0!
0*
09
0>
0C
#274710000000
1!
1*
b101 6
19
1>
1C
b101 G
#274720000000
0!
0*
09
0>
0C
#274730000000
1!
1*
b110 6
19
1>
1C
b110 G
#274740000000
0!
0*
09
0>
0C
#274750000000
1!
1*
b111 6
19
1>
1C
b111 G
#274760000000
0!
1"
0*
1+
09
1:
0>
0C
#274770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#274780000000
0!
0*
09
0>
0C
#274790000000
1!
1*
b1 6
19
1>
1C
b1 G
#274800000000
0!
0*
09
0>
0C
#274810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#274820000000
0!
0*
09
0>
0C
#274830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#274840000000
0!
0*
09
0>
0C
#274850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#274860000000
0!
0*
09
0>
0C
#274870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#274880000000
0!
0#
0*
0,
09
0>
0?
0C
#274890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#274900000000
0!
0*
09
0>
0C
#274910000000
1!
1*
19
1>
1C
#274920000000
0!
0*
09
0>
0C
#274930000000
1!
1*
19
1>
1C
#274940000000
0!
0*
09
0>
0C
#274950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#274960000000
0!
0*
09
0>
0C
#274970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#274980000000
0!
0*
09
0>
0C
#274990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#275000000000
0!
0*
09
0>
0C
#275010000000
1!
1*
b10 6
19
1>
1C
b10 G
#275020000000
0!
0*
09
0>
0C
#275030000000
1!
1*
b11 6
19
1>
1C
b11 G
#275040000000
0!
0*
09
0>
0C
#275050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#275060000000
0!
0*
09
0>
0C
#275070000000
1!
1*
b101 6
19
1>
1C
b101 G
#275080000000
0!
0*
09
0>
0C
#275090000000
1!
1*
b110 6
19
1>
1C
b110 G
#275100000000
0!
0*
09
0>
0C
#275110000000
1!
1*
b111 6
19
1>
1C
b111 G
#275120000000
0!
0*
09
0>
0C
#275130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#275140000000
0!
0*
09
0>
0C
#275150000000
1!
1*
b1 6
19
1>
1C
b1 G
#275160000000
0!
0*
09
0>
0C
#275170000000
1!
1*
b10 6
19
1>
1C
b10 G
#275180000000
0!
0*
09
0>
0C
#275190000000
1!
1*
b11 6
19
1>
1C
b11 G
#275200000000
0!
0*
09
0>
0C
#275210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#275220000000
0!
0*
09
0>
0C
#275230000000
1!
1*
b101 6
19
1>
1C
b101 G
#275240000000
0!
0*
09
0>
0C
#275250000000
1!
1*
b110 6
19
1>
1C
b110 G
#275260000000
0!
0*
09
0>
0C
#275270000000
1!
1*
b111 6
19
1>
1C
b111 G
#275280000000
0!
0*
09
0>
0C
#275290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#275300000000
0!
0*
09
0>
0C
#275310000000
1!
1*
b1 6
19
1>
1C
b1 G
#275320000000
0!
0*
09
0>
0C
#275330000000
1!
1*
b10 6
19
1>
1C
b10 G
#275340000000
0!
0*
09
0>
0C
#275350000000
1!
1*
b11 6
19
1>
1C
b11 G
#275360000000
0!
0*
09
0>
0C
#275370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#275380000000
0!
0*
09
0>
0C
#275390000000
1!
1*
b101 6
19
1>
1C
b101 G
#275400000000
0!
0*
09
0>
0C
#275410000000
1!
1*
b110 6
19
1>
1C
b110 G
#275420000000
0!
0*
09
0>
0C
#275430000000
1!
1*
b111 6
19
1>
1C
b111 G
#275440000000
0!
1"
0*
1+
09
1:
0>
0C
#275450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#275460000000
0!
0*
09
0>
0C
#275470000000
1!
1*
b1 6
19
1>
1C
b1 G
#275480000000
0!
0*
09
0>
0C
#275490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#275500000000
0!
0*
09
0>
0C
#275510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#275520000000
0!
0*
09
0>
0C
#275530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#275540000000
0!
0*
09
0>
0C
#275550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#275560000000
0!
0#
0*
0,
09
0>
0?
0C
#275570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#275580000000
0!
0*
09
0>
0C
#275590000000
1!
1*
19
1>
1C
#275600000000
0!
0*
09
0>
0C
#275610000000
1!
1*
19
1>
1C
#275620000000
0!
0*
09
0>
0C
#275630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#275640000000
0!
0*
09
0>
0C
#275650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#275660000000
0!
0*
09
0>
0C
#275670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#275680000000
0!
0*
09
0>
0C
#275690000000
1!
1*
b10 6
19
1>
1C
b10 G
#275700000000
0!
0*
09
0>
0C
#275710000000
1!
1*
b11 6
19
1>
1C
b11 G
#275720000000
0!
0*
09
0>
0C
#275730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#275740000000
0!
0*
09
0>
0C
#275750000000
1!
1*
b101 6
19
1>
1C
b101 G
#275760000000
0!
0*
09
0>
0C
#275770000000
1!
1*
b110 6
19
1>
1C
b110 G
#275780000000
0!
0*
09
0>
0C
#275790000000
1!
1*
b111 6
19
1>
1C
b111 G
#275800000000
0!
0*
09
0>
0C
#275810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#275820000000
0!
0*
09
0>
0C
#275830000000
1!
1*
b1 6
19
1>
1C
b1 G
#275840000000
0!
0*
09
0>
0C
#275850000000
1!
1*
b10 6
19
1>
1C
b10 G
#275860000000
0!
0*
09
0>
0C
#275870000000
1!
1*
b11 6
19
1>
1C
b11 G
#275880000000
0!
0*
09
0>
0C
#275890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#275900000000
0!
0*
09
0>
0C
#275910000000
1!
1*
b101 6
19
1>
1C
b101 G
#275920000000
0!
0*
09
0>
0C
#275930000000
1!
1*
b110 6
19
1>
1C
b110 G
#275940000000
0!
0*
09
0>
0C
#275950000000
1!
1*
b111 6
19
1>
1C
b111 G
#275960000000
0!
0*
09
0>
0C
#275970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#275980000000
0!
0*
09
0>
0C
#275990000000
1!
1*
b1 6
19
1>
1C
b1 G
#276000000000
0!
0*
09
0>
0C
#276010000000
1!
1*
b10 6
19
1>
1C
b10 G
#276020000000
0!
0*
09
0>
0C
#276030000000
1!
1*
b11 6
19
1>
1C
b11 G
#276040000000
0!
0*
09
0>
0C
#276050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#276060000000
0!
0*
09
0>
0C
#276070000000
1!
1*
b101 6
19
1>
1C
b101 G
#276080000000
0!
0*
09
0>
0C
#276090000000
1!
1*
b110 6
19
1>
1C
b110 G
#276100000000
0!
0*
09
0>
0C
#276110000000
1!
1*
b111 6
19
1>
1C
b111 G
#276120000000
0!
1"
0*
1+
09
1:
0>
0C
#276130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#276140000000
0!
0*
09
0>
0C
#276150000000
1!
1*
b1 6
19
1>
1C
b1 G
#276160000000
0!
0*
09
0>
0C
#276170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#276180000000
0!
0*
09
0>
0C
#276190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#276200000000
0!
0*
09
0>
0C
#276210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#276220000000
0!
0*
09
0>
0C
#276230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#276240000000
0!
0#
0*
0,
09
0>
0?
0C
#276250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#276260000000
0!
0*
09
0>
0C
#276270000000
1!
1*
19
1>
1C
#276280000000
0!
0*
09
0>
0C
#276290000000
1!
1*
19
1>
1C
#276300000000
0!
0*
09
0>
0C
#276310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#276320000000
0!
0*
09
0>
0C
#276330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#276340000000
0!
0*
09
0>
0C
#276350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#276360000000
0!
0*
09
0>
0C
#276370000000
1!
1*
b10 6
19
1>
1C
b10 G
#276380000000
0!
0*
09
0>
0C
#276390000000
1!
1*
b11 6
19
1>
1C
b11 G
#276400000000
0!
0*
09
0>
0C
#276410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#276420000000
0!
0*
09
0>
0C
#276430000000
1!
1*
b101 6
19
1>
1C
b101 G
#276440000000
0!
0*
09
0>
0C
#276450000000
1!
1*
b110 6
19
1>
1C
b110 G
#276460000000
0!
0*
09
0>
0C
#276470000000
1!
1*
b111 6
19
1>
1C
b111 G
#276480000000
0!
0*
09
0>
0C
#276490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#276500000000
0!
0*
09
0>
0C
#276510000000
1!
1*
b1 6
19
1>
1C
b1 G
#276520000000
0!
0*
09
0>
0C
#276530000000
1!
1*
b10 6
19
1>
1C
b10 G
#276540000000
0!
0*
09
0>
0C
#276550000000
1!
1*
b11 6
19
1>
1C
b11 G
#276560000000
0!
0*
09
0>
0C
#276570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#276580000000
0!
0*
09
0>
0C
#276590000000
1!
1*
b101 6
19
1>
1C
b101 G
#276600000000
0!
0*
09
0>
0C
#276610000000
1!
1*
b110 6
19
1>
1C
b110 G
#276620000000
0!
0*
09
0>
0C
#276630000000
1!
1*
b111 6
19
1>
1C
b111 G
#276640000000
0!
0*
09
0>
0C
#276650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#276660000000
0!
0*
09
0>
0C
#276670000000
1!
1*
b1 6
19
1>
1C
b1 G
#276680000000
0!
0*
09
0>
0C
#276690000000
1!
1*
b10 6
19
1>
1C
b10 G
#276700000000
0!
0*
09
0>
0C
#276710000000
1!
1*
b11 6
19
1>
1C
b11 G
#276720000000
0!
0*
09
0>
0C
#276730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#276740000000
0!
0*
09
0>
0C
#276750000000
1!
1*
b101 6
19
1>
1C
b101 G
#276760000000
0!
0*
09
0>
0C
#276770000000
1!
1*
b110 6
19
1>
1C
b110 G
#276780000000
0!
0*
09
0>
0C
#276790000000
1!
1*
b111 6
19
1>
1C
b111 G
#276800000000
0!
1"
0*
1+
09
1:
0>
0C
#276810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#276820000000
0!
0*
09
0>
0C
#276830000000
1!
1*
b1 6
19
1>
1C
b1 G
#276840000000
0!
0*
09
0>
0C
#276850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#276860000000
0!
0*
09
0>
0C
#276870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#276880000000
0!
0*
09
0>
0C
#276890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#276900000000
0!
0*
09
0>
0C
#276910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#276920000000
0!
0#
0*
0,
09
0>
0?
0C
#276930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#276940000000
0!
0*
09
0>
0C
#276950000000
1!
1*
19
1>
1C
#276960000000
0!
0*
09
0>
0C
#276970000000
1!
1*
19
1>
1C
#276980000000
0!
0*
09
0>
0C
#276990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#277000000000
0!
0*
09
0>
0C
#277010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#277020000000
0!
0*
09
0>
0C
#277030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#277040000000
0!
0*
09
0>
0C
#277050000000
1!
1*
b10 6
19
1>
1C
b10 G
#277060000000
0!
0*
09
0>
0C
#277070000000
1!
1*
b11 6
19
1>
1C
b11 G
#277080000000
0!
0*
09
0>
0C
#277090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#277100000000
0!
0*
09
0>
0C
#277110000000
1!
1*
b101 6
19
1>
1C
b101 G
#277120000000
0!
0*
09
0>
0C
#277130000000
1!
1*
b110 6
19
1>
1C
b110 G
#277140000000
0!
0*
09
0>
0C
#277150000000
1!
1*
b111 6
19
1>
1C
b111 G
#277160000000
0!
0*
09
0>
0C
#277170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#277180000000
0!
0*
09
0>
0C
#277190000000
1!
1*
b1 6
19
1>
1C
b1 G
#277200000000
0!
0*
09
0>
0C
#277210000000
1!
1*
b10 6
19
1>
1C
b10 G
#277220000000
0!
0*
09
0>
0C
#277230000000
1!
1*
b11 6
19
1>
1C
b11 G
#277240000000
0!
0*
09
0>
0C
#277250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#277260000000
0!
0*
09
0>
0C
#277270000000
1!
1*
b101 6
19
1>
1C
b101 G
#277280000000
0!
0*
09
0>
0C
#277290000000
1!
1*
b110 6
19
1>
1C
b110 G
#277300000000
0!
0*
09
0>
0C
#277310000000
1!
1*
b111 6
19
1>
1C
b111 G
#277320000000
0!
0*
09
0>
0C
#277330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#277340000000
0!
0*
09
0>
0C
#277350000000
1!
1*
b1 6
19
1>
1C
b1 G
#277360000000
0!
0*
09
0>
0C
#277370000000
1!
1*
b10 6
19
1>
1C
b10 G
#277380000000
0!
0*
09
0>
0C
#277390000000
1!
1*
b11 6
19
1>
1C
b11 G
#277400000000
0!
0*
09
0>
0C
#277410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#277420000000
0!
0*
09
0>
0C
#277430000000
1!
1*
b101 6
19
1>
1C
b101 G
#277440000000
0!
0*
09
0>
0C
#277450000000
1!
1*
b110 6
19
1>
1C
b110 G
#277460000000
0!
0*
09
0>
0C
#277470000000
1!
1*
b111 6
19
1>
1C
b111 G
#277480000000
0!
1"
0*
1+
09
1:
0>
0C
#277490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#277500000000
0!
0*
09
0>
0C
#277510000000
1!
1*
b1 6
19
1>
1C
b1 G
#277520000000
0!
0*
09
0>
0C
#277530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#277540000000
0!
0*
09
0>
0C
#277550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#277560000000
0!
0*
09
0>
0C
#277570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#277580000000
0!
0*
09
0>
0C
#277590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#277600000000
0!
0#
0*
0,
09
0>
0?
0C
#277610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#277620000000
0!
0*
09
0>
0C
#277630000000
1!
1*
19
1>
1C
#277640000000
0!
0*
09
0>
0C
#277650000000
1!
1*
19
1>
1C
#277660000000
0!
0*
09
0>
0C
#277670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#277680000000
0!
0*
09
0>
0C
#277690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#277700000000
0!
0*
09
0>
0C
#277710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#277720000000
0!
0*
09
0>
0C
#277730000000
1!
1*
b10 6
19
1>
1C
b10 G
#277740000000
0!
0*
09
0>
0C
#277750000000
1!
1*
b11 6
19
1>
1C
b11 G
#277760000000
0!
0*
09
0>
0C
#277770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#277780000000
0!
0*
09
0>
0C
#277790000000
1!
1*
b101 6
19
1>
1C
b101 G
#277800000000
0!
0*
09
0>
0C
#277810000000
1!
1*
b110 6
19
1>
1C
b110 G
#277820000000
0!
0*
09
0>
0C
#277830000000
1!
1*
b111 6
19
1>
1C
b111 G
#277840000000
0!
0*
09
0>
0C
#277850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#277860000000
0!
0*
09
0>
0C
#277870000000
1!
1*
b1 6
19
1>
1C
b1 G
#277880000000
0!
0*
09
0>
0C
#277890000000
1!
1*
b10 6
19
1>
1C
b10 G
#277900000000
0!
0*
09
0>
0C
#277910000000
1!
1*
b11 6
19
1>
1C
b11 G
#277920000000
0!
0*
09
0>
0C
#277930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#277940000000
0!
0*
09
0>
0C
#277950000000
1!
1*
b101 6
19
1>
1C
b101 G
#277960000000
0!
0*
09
0>
0C
#277970000000
1!
1*
b110 6
19
1>
1C
b110 G
#277980000000
0!
0*
09
0>
0C
#277990000000
1!
1*
b111 6
19
1>
1C
b111 G
#278000000000
0!
0*
09
0>
0C
#278010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#278020000000
0!
0*
09
0>
0C
#278030000000
1!
1*
b1 6
19
1>
1C
b1 G
#278040000000
0!
0*
09
0>
0C
#278050000000
1!
1*
b10 6
19
1>
1C
b10 G
#278060000000
0!
0*
09
0>
0C
#278070000000
1!
1*
b11 6
19
1>
1C
b11 G
#278080000000
0!
0*
09
0>
0C
#278090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#278100000000
0!
0*
09
0>
0C
#278110000000
1!
1*
b101 6
19
1>
1C
b101 G
#278120000000
0!
0*
09
0>
0C
#278130000000
1!
1*
b110 6
19
1>
1C
b110 G
#278140000000
0!
0*
09
0>
0C
#278150000000
1!
1*
b111 6
19
1>
1C
b111 G
#278160000000
0!
1"
0*
1+
09
1:
0>
0C
#278170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#278180000000
0!
0*
09
0>
0C
#278190000000
1!
1*
b1 6
19
1>
1C
b1 G
#278200000000
0!
0*
09
0>
0C
#278210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#278220000000
0!
0*
09
0>
0C
#278230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#278240000000
0!
0*
09
0>
0C
#278250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#278260000000
0!
0*
09
0>
0C
#278270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#278280000000
0!
0#
0*
0,
09
0>
0?
0C
#278290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#278300000000
0!
0*
09
0>
0C
#278310000000
1!
1*
19
1>
1C
#278320000000
0!
0*
09
0>
0C
#278330000000
1!
1*
19
1>
1C
#278340000000
0!
0*
09
0>
0C
#278350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#278360000000
0!
0*
09
0>
0C
#278370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#278380000000
0!
0*
09
0>
0C
#278390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#278400000000
0!
0*
09
0>
0C
#278410000000
1!
1*
b10 6
19
1>
1C
b10 G
#278420000000
0!
0*
09
0>
0C
#278430000000
1!
1*
b11 6
19
1>
1C
b11 G
#278440000000
0!
0*
09
0>
0C
#278450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#278460000000
0!
0*
09
0>
0C
#278470000000
1!
1*
b101 6
19
1>
1C
b101 G
#278480000000
0!
0*
09
0>
0C
#278490000000
1!
1*
b110 6
19
1>
1C
b110 G
#278500000000
0!
0*
09
0>
0C
#278510000000
1!
1*
b111 6
19
1>
1C
b111 G
#278520000000
0!
0*
09
0>
0C
#278530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#278540000000
0!
0*
09
0>
0C
#278550000000
1!
1*
b1 6
19
1>
1C
b1 G
#278560000000
0!
0*
09
0>
0C
#278570000000
1!
1*
b10 6
19
1>
1C
b10 G
#278580000000
0!
0*
09
0>
0C
#278590000000
1!
1*
b11 6
19
1>
1C
b11 G
#278600000000
0!
0*
09
0>
0C
#278610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#278620000000
0!
0*
09
0>
0C
#278630000000
1!
1*
b101 6
19
1>
1C
b101 G
#278640000000
0!
0*
09
0>
0C
#278650000000
1!
1*
b110 6
19
1>
1C
b110 G
#278660000000
0!
0*
09
0>
0C
#278670000000
1!
1*
b111 6
19
1>
1C
b111 G
#278680000000
0!
0*
09
0>
0C
#278690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#278700000000
0!
0*
09
0>
0C
#278710000000
1!
1*
b1 6
19
1>
1C
b1 G
#278720000000
0!
0*
09
0>
0C
#278730000000
1!
1*
b10 6
19
1>
1C
b10 G
#278740000000
0!
0*
09
0>
0C
#278750000000
1!
1*
b11 6
19
1>
1C
b11 G
#278760000000
0!
0*
09
0>
0C
#278770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#278780000000
0!
0*
09
0>
0C
#278790000000
1!
1*
b101 6
19
1>
1C
b101 G
#278800000000
0!
0*
09
0>
0C
#278810000000
1!
1*
b110 6
19
1>
1C
b110 G
#278820000000
0!
0*
09
0>
0C
#278830000000
1!
1*
b111 6
19
1>
1C
b111 G
#278840000000
0!
1"
0*
1+
09
1:
0>
0C
#278850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#278860000000
0!
0*
09
0>
0C
#278870000000
1!
1*
b1 6
19
1>
1C
b1 G
#278880000000
0!
0*
09
0>
0C
#278890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#278900000000
0!
0*
09
0>
0C
#278910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#278920000000
0!
0*
09
0>
0C
#278930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#278940000000
0!
0*
09
0>
0C
#278950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#278960000000
0!
0#
0*
0,
09
0>
0?
0C
#278970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#278980000000
0!
0*
09
0>
0C
#278990000000
1!
1*
19
1>
1C
#279000000000
0!
0*
09
0>
0C
#279010000000
1!
1*
19
1>
1C
#279020000000
0!
0*
09
0>
0C
#279030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#279040000000
0!
0*
09
0>
0C
#279050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#279060000000
0!
0*
09
0>
0C
#279070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#279080000000
0!
0*
09
0>
0C
#279090000000
1!
1*
b10 6
19
1>
1C
b10 G
#279100000000
0!
0*
09
0>
0C
#279110000000
1!
1*
b11 6
19
1>
1C
b11 G
#279120000000
0!
0*
09
0>
0C
#279130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#279140000000
0!
0*
09
0>
0C
#279150000000
1!
1*
b101 6
19
1>
1C
b101 G
#279160000000
0!
0*
09
0>
0C
#279170000000
1!
1*
b110 6
19
1>
1C
b110 G
#279180000000
0!
0*
09
0>
0C
#279190000000
1!
1*
b111 6
19
1>
1C
b111 G
#279200000000
0!
0*
09
0>
0C
#279210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#279220000000
0!
0*
09
0>
0C
#279230000000
1!
1*
b1 6
19
1>
1C
b1 G
#279240000000
0!
0*
09
0>
0C
#279250000000
1!
1*
b10 6
19
1>
1C
b10 G
#279260000000
0!
0*
09
0>
0C
#279270000000
1!
1*
b11 6
19
1>
1C
b11 G
#279280000000
0!
0*
09
0>
0C
#279290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#279300000000
0!
0*
09
0>
0C
#279310000000
1!
1*
b101 6
19
1>
1C
b101 G
#279320000000
0!
0*
09
0>
0C
#279330000000
1!
1*
b110 6
19
1>
1C
b110 G
#279340000000
0!
0*
09
0>
0C
#279350000000
1!
1*
b111 6
19
1>
1C
b111 G
#279360000000
0!
0*
09
0>
0C
#279370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#279380000000
0!
0*
09
0>
0C
#279390000000
1!
1*
b1 6
19
1>
1C
b1 G
#279400000000
0!
0*
09
0>
0C
#279410000000
1!
1*
b10 6
19
1>
1C
b10 G
#279420000000
0!
0*
09
0>
0C
#279430000000
1!
1*
b11 6
19
1>
1C
b11 G
#279440000000
0!
0*
09
0>
0C
#279450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#279460000000
0!
0*
09
0>
0C
#279470000000
1!
1*
b101 6
19
1>
1C
b101 G
#279480000000
0!
0*
09
0>
0C
#279490000000
1!
1*
b110 6
19
1>
1C
b110 G
#279500000000
0!
0*
09
0>
0C
#279510000000
1!
1*
b111 6
19
1>
1C
b111 G
#279520000000
0!
1"
0*
1+
09
1:
0>
0C
#279530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#279540000000
0!
0*
09
0>
0C
#279550000000
1!
1*
b1 6
19
1>
1C
b1 G
#279560000000
0!
0*
09
0>
0C
#279570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#279580000000
0!
0*
09
0>
0C
#279590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#279600000000
0!
0*
09
0>
0C
#279610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#279620000000
0!
0*
09
0>
0C
#279630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#279640000000
0!
0#
0*
0,
09
0>
0?
0C
#279650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#279660000000
0!
0*
09
0>
0C
#279670000000
1!
1*
19
1>
1C
#279680000000
0!
0*
09
0>
0C
#279690000000
1!
1*
19
1>
1C
#279700000000
0!
0*
09
0>
0C
#279710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#279720000000
0!
0*
09
0>
0C
#279730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#279740000000
0!
0*
09
0>
0C
#279750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#279760000000
0!
0*
09
0>
0C
#279770000000
1!
1*
b10 6
19
1>
1C
b10 G
#279780000000
0!
0*
09
0>
0C
#279790000000
1!
1*
b11 6
19
1>
1C
b11 G
#279800000000
0!
0*
09
0>
0C
#279810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#279820000000
0!
0*
09
0>
0C
#279830000000
1!
1*
b101 6
19
1>
1C
b101 G
#279840000000
0!
0*
09
0>
0C
#279850000000
1!
1*
b110 6
19
1>
1C
b110 G
#279860000000
0!
0*
09
0>
0C
#279870000000
1!
1*
b111 6
19
1>
1C
b111 G
#279880000000
0!
0*
09
0>
0C
#279890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#279900000000
0!
0*
09
0>
0C
#279910000000
1!
1*
b1 6
19
1>
1C
b1 G
#279920000000
0!
0*
09
0>
0C
#279930000000
1!
1*
b10 6
19
1>
1C
b10 G
#279940000000
0!
0*
09
0>
0C
#279950000000
1!
1*
b11 6
19
1>
1C
b11 G
#279960000000
0!
0*
09
0>
0C
#279970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#279980000000
0!
0*
09
0>
0C
#279990000000
1!
1*
b101 6
19
1>
1C
b101 G
#280000000000
0!
0*
09
0>
0C
#280010000000
1!
1*
b110 6
19
1>
1C
b110 G
#280020000000
0!
0*
09
0>
0C
#280030000000
1!
1*
b111 6
19
1>
1C
b111 G
#280040000000
0!
0*
09
0>
0C
#280050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#280060000000
0!
0*
09
0>
0C
#280070000000
1!
1*
b1 6
19
1>
1C
b1 G
#280080000000
0!
0*
09
0>
0C
#280090000000
1!
1*
b10 6
19
1>
1C
b10 G
#280100000000
0!
0*
09
0>
0C
#280110000000
1!
1*
b11 6
19
1>
1C
b11 G
#280120000000
0!
0*
09
0>
0C
#280130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#280140000000
0!
0*
09
0>
0C
#280150000000
1!
1*
b101 6
19
1>
1C
b101 G
#280160000000
0!
0*
09
0>
0C
#280170000000
1!
1*
b110 6
19
1>
1C
b110 G
#280180000000
0!
0*
09
0>
0C
#280190000000
1!
1*
b111 6
19
1>
1C
b111 G
#280200000000
0!
1"
0*
1+
09
1:
0>
0C
#280210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#280220000000
0!
0*
09
0>
0C
#280230000000
1!
1*
b1 6
19
1>
1C
b1 G
#280240000000
0!
0*
09
0>
0C
#280250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#280260000000
0!
0*
09
0>
0C
#280270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#280280000000
0!
0*
09
0>
0C
#280290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#280300000000
0!
0*
09
0>
0C
#280310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#280320000000
0!
0#
0*
0,
09
0>
0?
0C
#280330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#280340000000
0!
0*
09
0>
0C
#280350000000
1!
1*
19
1>
1C
#280360000000
0!
0*
09
0>
0C
#280370000000
1!
1*
19
1>
1C
#280380000000
0!
0*
09
0>
0C
#280390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#280400000000
0!
0*
09
0>
0C
#280410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#280420000000
0!
0*
09
0>
0C
#280430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#280440000000
0!
0*
09
0>
0C
#280450000000
1!
1*
b10 6
19
1>
1C
b10 G
#280460000000
0!
0*
09
0>
0C
#280470000000
1!
1*
b11 6
19
1>
1C
b11 G
#280480000000
0!
0*
09
0>
0C
#280490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#280500000000
0!
0*
09
0>
0C
#280510000000
1!
1*
b101 6
19
1>
1C
b101 G
#280520000000
0!
0*
09
0>
0C
#280530000000
1!
1*
b110 6
19
1>
1C
b110 G
#280540000000
0!
0*
09
0>
0C
#280550000000
1!
1*
b111 6
19
1>
1C
b111 G
#280560000000
0!
0*
09
0>
0C
#280570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#280580000000
0!
0*
09
0>
0C
#280590000000
1!
1*
b1 6
19
1>
1C
b1 G
#280600000000
0!
0*
09
0>
0C
#280610000000
1!
1*
b10 6
19
1>
1C
b10 G
#280620000000
0!
0*
09
0>
0C
#280630000000
1!
1*
b11 6
19
1>
1C
b11 G
#280640000000
0!
0*
09
0>
0C
#280650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#280660000000
0!
0*
09
0>
0C
#280670000000
1!
1*
b101 6
19
1>
1C
b101 G
#280680000000
0!
0*
09
0>
0C
#280690000000
1!
1*
b110 6
19
1>
1C
b110 G
#280700000000
0!
0*
09
0>
0C
#280710000000
1!
1*
b111 6
19
1>
1C
b111 G
#280720000000
0!
0*
09
0>
0C
#280730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#280740000000
0!
0*
09
0>
0C
#280750000000
1!
1*
b1 6
19
1>
1C
b1 G
#280760000000
0!
0*
09
0>
0C
#280770000000
1!
1*
b10 6
19
1>
1C
b10 G
#280780000000
0!
0*
09
0>
0C
#280790000000
1!
1*
b11 6
19
1>
1C
b11 G
#280800000000
0!
0*
09
0>
0C
#280810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#280820000000
0!
0*
09
0>
0C
#280830000000
1!
1*
b101 6
19
1>
1C
b101 G
#280840000000
0!
0*
09
0>
0C
#280850000000
1!
1*
b110 6
19
1>
1C
b110 G
#280860000000
0!
0*
09
0>
0C
#280870000000
1!
1*
b111 6
19
1>
1C
b111 G
#280880000000
0!
1"
0*
1+
09
1:
0>
0C
#280890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#280900000000
0!
0*
09
0>
0C
#280910000000
1!
1*
b1 6
19
1>
1C
b1 G
#280920000000
0!
0*
09
0>
0C
#280930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#280940000000
0!
0*
09
0>
0C
#280950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#280960000000
0!
0*
09
0>
0C
#280970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#280980000000
0!
0*
09
0>
0C
#280990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#281000000000
0!
0#
0*
0,
09
0>
0?
0C
#281010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#281020000000
0!
0*
09
0>
0C
#281030000000
1!
1*
19
1>
1C
#281040000000
0!
0*
09
0>
0C
#281050000000
1!
1*
19
1>
1C
#281060000000
0!
0*
09
0>
0C
#281070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#281080000000
0!
0*
09
0>
0C
#281090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#281100000000
0!
0*
09
0>
0C
#281110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#281120000000
0!
0*
09
0>
0C
#281130000000
1!
1*
b10 6
19
1>
1C
b10 G
#281140000000
0!
0*
09
0>
0C
#281150000000
1!
1*
b11 6
19
1>
1C
b11 G
#281160000000
0!
0*
09
0>
0C
#281170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#281180000000
0!
0*
09
0>
0C
#281190000000
1!
1*
b101 6
19
1>
1C
b101 G
#281200000000
0!
0*
09
0>
0C
#281210000000
1!
1*
b110 6
19
1>
1C
b110 G
#281220000000
0!
0*
09
0>
0C
#281230000000
1!
1*
b111 6
19
1>
1C
b111 G
#281240000000
0!
0*
09
0>
0C
#281250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#281260000000
0!
0*
09
0>
0C
#281270000000
1!
1*
b1 6
19
1>
1C
b1 G
#281280000000
0!
0*
09
0>
0C
#281290000000
1!
1*
b10 6
19
1>
1C
b10 G
#281300000000
0!
0*
09
0>
0C
#281310000000
1!
1*
b11 6
19
1>
1C
b11 G
#281320000000
0!
0*
09
0>
0C
#281330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#281340000000
0!
0*
09
0>
0C
#281350000000
1!
1*
b101 6
19
1>
1C
b101 G
#281360000000
0!
0*
09
0>
0C
#281370000000
1!
1*
b110 6
19
1>
1C
b110 G
#281380000000
0!
0*
09
0>
0C
#281390000000
1!
1*
b111 6
19
1>
1C
b111 G
#281400000000
0!
0*
09
0>
0C
#281410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#281420000000
0!
0*
09
0>
0C
#281430000000
1!
1*
b1 6
19
1>
1C
b1 G
#281440000000
0!
0*
09
0>
0C
#281450000000
1!
1*
b10 6
19
1>
1C
b10 G
#281460000000
0!
0*
09
0>
0C
#281470000000
1!
1*
b11 6
19
1>
1C
b11 G
#281480000000
0!
0*
09
0>
0C
#281490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#281500000000
0!
0*
09
0>
0C
#281510000000
1!
1*
b101 6
19
1>
1C
b101 G
#281520000000
0!
0*
09
0>
0C
#281530000000
1!
1*
b110 6
19
1>
1C
b110 G
#281540000000
0!
0*
09
0>
0C
#281550000000
1!
1*
b111 6
19
1>
1C
b111 G
#281560000000
0!
1"
0*
1+
09
1:
0>
0C
#281570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#281580000000
0!
0*
09
0>
0C
#281590000000
1!
1*
b1 6
19
1>
1C
b1 G
#281600000000
0!
0*
09
0>
0C
#281610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#281620000000
0!
0*
09
0>
0C
#281630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#281640000000
0!
0*
09
0>
0C
#281650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#281660000000
0!
0*
09
0>
0C
#281670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#281680000000
0!
0#
0*
0,
09
0>
0?
0C
#281690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#281700000000
0!
0*
09
0>
0C
#281710000000
1!
1*
19
1>
1C
#281720000000
0!
0*
09
0>
0C
#281730000000
1!
1*
19
1>
1C
#281740000000
0!
0*
09
0>
0C
#281750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#281760000000
0!
0*
09
0>
0C
#281770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#281780000000
0!
0*
09
0>
0C
#281790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#281800000000
0!
0*
09
0>
0C
#281810000000
1!
1*
b10 6
19
1>
1C
b10 G
#281820000000
0!
0*
09
0>
0C
#281830000000
1!
1*
b11 6
19
1>
1C
b11 G
#281840000000
0!
0*
09
0>
0C
#281850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#281860000000
0!
0*
09
0>
0C
#281870000000
1!
1*
b101 6
19
1>
1C
b101 G
#281880000000
0!
0*
09
0>
0C
#281890000000
1!
1*
b110 6
19
1>
1C
b110 G
#281900000000
0!
0*
09
0>
0C
#281910000000
1!
1*
b111 6
19
1>
1C
b111 G
#281920000000
0!
0*
09
0>
0C
#281930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#281940000000
0!
0*
09
0>
0C
#281950000000
1!
1*
b1 6
19
1>
1C
b1 G
#281960000000
0!
0*
09
0>
0C
#281970000000
1!
1*
b10 6
19
1>
1C
b10 G
#281980000000
0!
0*
09
0>
0C
#281990000000
1!
1*
b11 6
19
1>
1C
b11 G
#282000000000
0!
0*
09
0>
0C
#282010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#282020000000
0!
0*
09
0>
0C
#282030000000
1!
1*
b101 6
19
1>
1C
b101 G
#282040000000
0!
0*
09
0>
0C
#282050000000
1!
1*
b110 6
19
1>
1C
b110 G
#282060000000
0!
0*
09
0>
0C
#282070000000
1!
1*
b111 6
19
1>
1C
b111 G
#282080000000
0!
0*
09
0>
0C
#282090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#282100000000
0!
0*
09
0>
0C
#282110000000
1!
1*
b1 6
19
1>
1C
b1 G
#282120000000
0!
0*
09
0>
0C
#282130000000
1!
1*
b10 6
19
1>
1C
b10 G
#282140000000
0!
0*
09
0>
0C
#282150000000
1!
1*
b11 6
19
1>
1C
b11 G
#282160000000
0!
0*
09
0>
0C
#282170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#282180000000
0!
0*
09
0>
0C
#282190000000
1!
1*
b101 6
19
1>
1C
b101 G
#282200000000
0!
0*
09
0>
0C
#282210000000
1!
1*
b110 6
19
1>
1C
b110 G
#282220000000
0!
0*
09
0>
0C
#282230000000
1!
1*
b111 6
19
1>
1C
b111 G
#282240000000
0!
1"
0*
1+
09
1:
0>
0C
#282250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#282260000000
0!
0*
09
0>
0C
#282270000000
1!
1*
b1 6
19
1>
1C
b1 G
#282280000000
0!
0*
09
0>
0C
#282290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#282300000000
0!
0*
09
0>
0C
#282310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#282320000000
0!
0*
09
0>
0C
#282330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#282340000000
0!
0*
09
0>
0C
#282350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#282360000000
0!
0#
0*
0,
09
0>
0?
0C
#282370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#282380000000
0!
0*
09
0>
0C
#282390000000
1!
1*
19
1>
1C
#282400000000
0!
0*
09
0>
0C
#282410000000
1!
1*
19
1>
1C
#282420000000
0!
0*
09
0>
0C
#282430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#282440000000
0!
0*
09
0>
0C
#282450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#282460000000
0!
0*
09
0>
0C
#282470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#282480000000
0!
0*
09
0>
0C
#282490000000
1!
1*
b10 6
19
1>
1C
b10 G
#282500000000
0!
0*
09
0>
0C
#282510000000
1!
1*
b11 6
19
1>
1C
b11 G
#282520000000
0!
0*
09
0>
0C
#282530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#282540000000
0!
0*
09
0>
0C
#282550000000
1!
1*
b101 6
19
1>
1C
b101 G
#282560000000
0!
0*
09
0>
0C
#282570000000
1!
1*
b110 6
19
1>
1C
b110 G
#282580000000
0!
0*
09
0>
0C
#282590000000
1!
1*
b111 6
19
1>
1C
b111 G
#282600000000
0!
0*
09
0>
0C
#282610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#282620000000
0!
0*
09
0>
0C
#282630000000
1!
1*
b1 6
19
1>
1C
b1 G
#282640000000
0!
0*
09
0>
0C
#282650000000
1!
1*
b10 6
19
1>
1C
b10 G
#282660000000
0!
0*
09
0>
0C
#282670000000
1!
1*
b11 6
19
1>
1C
b11 G
#282680000000
0!
0*
09
0>
0C
#282690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#282700000000
0!
0*
09
0>
0C
#282710000000
1!
1*
b101 6
19
1>
1C
b101 G
#282720000000
0!
0*
09
0>
0C
#282730000000
1!
1*
b110 6
19
1>
1C
b110 G
#282740000000
0!
0*
09
0>
0C
#282750000000
1!
1*
b111 6
19
1>
1C
b111 G
#282760000000
0!
0*
09
0>
0C
#282770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#282780000000
0!
0*
09
0>
0C
#282790000000
1!
1*
b1 6
19
1>
1C
b1 G
#282800000000
0!
0*
09
0>
0C
#282810000000
1!
1*
b10 6
19
1>
1C
b10 G
#282820000000
0!
0*
09
0>
0C
#282830000000
1!
1*
b11 6
19
1>
1C
b11 G
#282840000000
0!
0*
09
0>
0C
#282850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#282860000000
0!
0*
09
0>
0C
#282870000000
1!
1*
b101 6
19
1>
1C
b101 G
#282880000000
0!
0*
09
0>
0C
#282890000000
1!
1*
b110 6
19
1>
1C
b110 G
#282900000000
0!
0*
09
0>
0C
#282910000000
1!
1*
b111 6
19
1>
1C
b111 G
#282920000000
0!
1"
0*
1+
09
1:
0>
0C
#282930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#282940000000
0!
0*
09
0>
0C
#282950000000
1!
1*
b1 6
19
1>
1C
b1 G
#282960000000
0!
0*
09
0>
0C
#282970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#282980000000
0!
0*
09
0>
0C
#282990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#283000000000
0!
0*
09
0>
0C
#283010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#283020000000
0!
0*
09
0>
0C
#283030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#283040000000
0!
0#
0*
0,
09
0>
0?
0C
#283050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#283060000000
0!
0*
09
0>
0C
#283070000000
1!
1*
19
1>
1C
#283080000000
0!
0*
09
0>
0C
#283090000000
1!
1*
19
1>
1C
#283100000000
0!
0*
09
0>
0C
#283110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#283120000000
0!
0*
09
0>
0C
#283130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#283140000000
0!
0*
09
0>
0C
#283150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#283160000000
0!
0*
09
0>
0C
#283170000000
1!
1*
b10 6
19
1>
1C
b10 G
#283180000000
0!
0*
09
0>
0C
#283190000000
1!
1*
b11 6
19
1>
1C
b11 G
#283200000000
0!
0*
09
0>
0C
#283210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#283220000000
0!
0*
09
0>
0C
#283230000000
1!
1*
b101 6
19
1>
1C
b101 G
#283240000000
0!
0*
09
0>
0C
#283250000000
1!
1*
b110 6
19
1>
1C
b110 G
#283260000000
0!
0*
09
0>
0C
#283270000000
1!
1*
b111 6
19
1>
1C
b111 G
#283280000000
0!
0*
09
0>
0C
#283290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#283300000000
0!
0*
09
0>
0C
#283310000000
1!
1*
b1 6
19
1>
1C
b1 G
#283320000000
0!
0*
09
0>
0C
#283330000000
1!
1*
b10 6
19
1>
1C
b10 G
#283340000000
0!
0*
09
0>
0C
#283350000000
1!
1*
b11 6
19
1>
1C
b11 G
#283360000000
0!
0*
09
0>
0C
#283370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#283380000000
0!
0*
09
0>
0C
#283390000000
1!
1*
b101 6
19
1>
1C
b101 G
#283400000000
0!
0*
09
0>
0C
#283410000000
1!
1*
b110 6
19
1>
1C
b110 G
#283420000000
0!
0*
09
0>
0C
#283430000000
1!
1*
b111 6
19
1>
1C
b111 G
#283440000000
0!
0*
09
0>
0C
#283450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#283460000000
0!
0*
09
0>
0C
#283470000000
1!
1*
b1 6
19
1>
1C
b1 G
#283480000000
0!
0*
09
0>
0C
#283490000000
1!
1*
b10 6
19
1>
1C
b10 G
#283500000000
0!
0*
09
0>
0C
#283510000000
1!
1*
b11 6
19
1>
1C
b11 G
#283520000000
0!
0*
09
0>
0C
#283530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#283540000000
0!
0*
09
0>
0C
#283550000000
1!
1*
b101 6
19
1>
1C
b101 G
#283560000000
0!
0*
09
0>
0C
#283570000000
1!
1*
b110 6
19
1>
1C
b110 G
#283580000000
0!
0*
09
0>
0C
#283590000000
1!
1*
b111 6
19
1>
1C
b111 G
#283600000000
0!
1"
0*
1+
09
1:
0>
0C
#283610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#283620000000
0!
0*
09
0>
0C
#283630000000
1!
1*
b1 6
19
1>
1C
b1 G
#283640000000
0!
0*
09
0>
0C
#283650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#283660000000
0!
0*
09
0>
0C
#283670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#283680000000
0!
0*
09
0>
0C
#283690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#283700000000
0!
0*
09
0>
0C
#283710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#283720000000
0!
0#
0*
0,
09
0>
0?
0C
#283730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#283740000000
0!
0*
09
0>
0C
#283750000000
1!
1*
19
1>
1C
#283760000000
0!
0*
09
0>
0C
#283770000000
1!
1*
19
1>
1C
#283780000000
0!
0*
09
0>
0C
#283790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#283800000000
0!
0*
09
0>
0C
#283810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#283820000000
0!
0*
09
0>
0C
#283830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#283840000000
0!
0*
09
0>
0C
#283850000000
1!
1*
b10 6
19
1>
1C
b10 G
#283860000000
0!
0*
09
0>
0C
#283870000000
1!
1*
b11 6
19
1>
1C
b11 G
#283880000000
0!
0*
09
0>
0C
#283890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#283900000000
0!
0*
09
0>
0C
#283910000000
1!
1*
b101 6
19
1>
1C
b101 G
#283920000000
0!
0*
09
0>
0C
#283930000000
1!
1*
b110 6
19
1>
1C
b110 G
#283940000000
0!
0*
09
0>
0C
#283950000000
1!
1*
b111 6
19
1>
1C
b111 G
#283960000000
0!
0*
09
0>
0C
#283970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#283980000000
0!
0*
09
0>
0C
#283990000000
1!
1*
b1 6
19
1>
1C
b1 G
#284000000000
0!
0*
09
0>
0C
#284010000000
1!
1*
b10 6
19
1>
1C
b10 G
#284020000000
0!
0*
09
0>
0C
#284030000000
1!
1*
b11 6
19
1>
1C
b11 G
#284040000000
0!
0*
09
0>
0C
#284050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#284060000000
0!
0*
09
0>
0C
#284070000000
1!
1*
b101 6
19
1>
1C
b101 G
#284080000000
0!
0*
09
0>
0C
#284090000000
1!
1*
b110 6
19
1>
1C
b110 G
#284100000000
0!
0*
09
0>
0C
#284110000000
1!
1*
b111 6
19
1>
1C
b111 G
#284120000000
0!
0*
09
0>
0C
#284130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#284140000000
0!
0*
09
0>
0C
#284150000000
1!
1*
b1 6
19
1>
1C
b1 G
#284160000000
0!
0*
09
0>
0C
#284170000000
1!
1*
b10 6
19
1>
1C
b10 G
#284180000000
0!
0*
09
0>
0C
#284190000000
1!
1*
b11 6
19
1>
1C
b11 G
#284200000000
0!
0*
09
0>
0C
#284210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#284220000000
0!
0*
09
0>
0C
#284230000000
1!
1*
b101 6
19
1>
1C
b101 G
#284240000000
0!
0*
09
0>
0C
#284250000000
1!
1*
b110 6
19
1>
1C
b110 G
#284260000000
0!
0*
09
0>
0C
#284270000000
1!
1*
b111 6
19
1>
1C
b111 G
#284280000000
0!
1"
0*
1+
09
1:
0>
0C
#284290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#284300000000
0!
0*
09
0>
0C
#284310000000
1!
1*
b1 6
19
1>
1C
b1 G
#284320000000
0!
0*
09
0>
0C
#284330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#284340000000
0!
0*
09
0>
0C
#284350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#284360000000
0!
0*
09
0>
0C
#284370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#284380000000
0!
0*
09
0>
0C
#284390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#284400000000
0!
0#
0*
0,
09
0>
0?
0C
#284410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#284420000000
0!
0*
09
0>
0C
#284430000000
1!
1*
19
1>
1C
#284440000000
0!
0*
09
0>
0C
#284450000000
1!
1*
19
1>
1C
#284460000000
0!
0*
09
0>
0C
#284470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#284480000000
0!
0*
09
0>
0C
#284490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#284500000000
0!
0*
09
0>
0C
#284510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#284520000000
0!
0*
09
0>
0C
#284530000000
1!
1*
b10 6
19
1>
1C
b10 G
#284540000000
0!
0*
09
0>
0C
#284550000000
1!
1*
b11 6
19
1>
1C
b11 G
#284560000000
0!
0*
09
0>
0C
#284570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#284580000000
0!
0*
09
0>
0C
#284590000000
1!
1*
b101 6
19
1>
1C
b101 G
#284600000000
0!
0*
09
0>
0C
#284610000000
1!
1*
b110 6
19
1>
1C
b110 G
#284620000000
0!
0*
09
0>
0C
#284630000000
1!
1*
b111 6
19
1>
1C
b111 G
#284640000000
0!
0*
09
0>
0C
#284650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#284660000000
0!
0*
09
0>
0C
#284670000000
1!
1*
b1 6
19
1>
1C
b1 G
#284680000000
0!
0*
09
0>
0C
#284690000000
1!
1*
b10 6
19
1>
1C
b10 G
#284700000000
0!
0*
09
0>
0C
#284710000000
1!
1*
b11 6
19
1>
1C
b11 G
#284720000000
0!
0*
09
0>
0C
#284730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#284740000000
0!
0*
09
0>
0C
#284750000000
1!
1*
b101 6
19
1>
1C
b101 G
#284760000000
0!
0*
09
0>
0C
#284770000000
1!
1*
b110 6
19
1>
1C
b110 G
#284780000000
0!
0*
09
0>
0C
#284790000000
1!
1*
b111 6
19
1>
1C
b111 G
#284800000000
0!
0*
09
0>
0C
#284810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#284820000000
0!
0*
09
0>
0C
#284830000000
1!
1*
b1 6
19
1>
1C
b1 G
#284840000000
0!
0*
09
0>
0C
#284850000000
1!
1*
b10 6
19
1>
1C
b10 G
#284860000000
0!
0*
09
0>
0C
#284870000000
1!
1*
b11 6
19
1>
1C
b11 G
#284880000000
0!
0*
09
0>
0C
#284890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#284900000000
0!
0*
09
0>
0C
#284910000000
1!
1*
b101 6
19
1>
1C
b101 G
#284920000000
0!
0*
09
0>
0C
#284930000000
1!
1*
b110 6
19
1>
1C
b110 G
#284940000000
0!
0*
09
0>
0C
#284950000000
1!
1*
b111 6
19
1>
1C
b111 G
#284960000000
0!
1"
0*
1+
09
1:
0>
0C
#284970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#284980000000
0!
0*
09
0>
0C
#284990000000
1!
1*
b1 6
19
1>
1C
b1 G
#285000000000
0!
0*
09
0>
0C
#285010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#285020000000
0!
0*
09
0>
0C
#285030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#285040000000
0!
0*
09
0>
0C
#285050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#285060000000
0!
0*
09
0>
0C
#285070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#285080000000
0!
0#
0*
0,
09
0>
0?
0C
#285090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#285100000000
0!
0*
09
0>
0C
#285110000000
1!
1*
19
1>
1C
#285120000000
0!
0*
09
0>
0C
#285130000000
1!
1*
19
1>
1C
#285140000000
0!
0*
09
0>
0C
#285150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#285160000000
0!
0*
09
0>
0C
#285170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#285180000000
0!
0*
09
0>
0C
#285190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#285200000000
0!
0*
09
0>
0C
#285210000000
1!
1*
b10 6
19
1>
1C
b10 G
#285220000000
0!
0*
09
0>
0C
#285230000000
1!
1*
b11 6
19
1>
1C
b11 G
#285240000000
0!
0*
09
0>
0C
#285250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#285260000000
0!
0*
09
0>
0C
#285270000000
1!
1*
b101 6
19
1>
1C
b101 G
#285280000000
0!
0*
09
0>
0C
#285290000000
1!
1*
b110 6
19
1>
1C
b110 G
#285300000000
0!
0*
09
0>
0C
#285310000000
1!
1*
b111 6
19
1>
1C
b111 G
#285320000000
0!
0*
09
0>
0C
#285330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#285340000000
0!
0*
09
0>
0C
#285350000000
1!
1*
b1 6
19
1>
1C
b1 G
#285360000000
0!
0*
09
0>
0C
#285370000000
1!
1*
b10 6
19
1>
1C
b10 G
#285380000000
0!
0*
09
0>
0C
#285390000000
1!
1*
b11 6
19
1>
1C
b11 G
#285400000000
0!
0*
09
0>
0C
#285410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#285420000000
0!
0*
09
0>
0C
#285430000000
1!
1*
b101 6
19
1>
1C
b101 G
#285440000000
0!
0*
09
0>
0C
#285450000000
1!
1*
b110 6
19
1>
1C
b110 G
#285460000000
0!
0*
09
0>
0C
#285470000000
1!
1*
b111 6
19
1>
1C
b111 G
#285480000000
0!
0*
09
0>
0C
#285490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#285500000000
0!
0*
09
0>
0C
#285510000000
1!
1*
b1 6
19
1>
1C
b1 G
#285520000000
0!
0*
09
0>
0C
#285530000000
1!
1*
b10 6
19
1>
1C
b10 G
#285540000000
0!
0*
09
0>
0C
#285550000000
1!
1*
b11 6
19
1>
1C
b11 G
#285560000000
0!
0*
09
0>
0C
#285570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#285580000000
0!
0*
09
0>
0C
#285590000000
1!
1*
b101 6
19
1>
1C
b101 G
#285600000000
0!
0*
09
0>
0C
#285610000000
1!
1*
b110 6
19
1>
1C
b110 G
#285620000000
0!
0*
09
0>
0C
#285630000000
1!
1*
b111 6
19
1>
1C
b111 G
#285640000000
0!
1"
0*
1+
09
1:
0>
0C
#285650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#285660000000
0!
0*
09
0>
0C
#285670000000
1!
1*
b1 6
19
1>
1C
b1 G
#285680000000
0!
0*
09
0>
0C
#285690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#285700000000
0!
0*
09
0>
0C
#285710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#285720000000
0!
0*
09
0>
0C
#285730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#285740000000
0!
0*
09
0>
0C
#285750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#285760000000
0!
0#
0*
0,
09
0>
0?
0C
#285770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#285780000000
0!
0*
09
0>
0C
#285790000000
1!
1*
19
1>
1C
#285800000000
0!
0*
09
0>
0C
#285810000000
1!
1*
19
1>
1C
#285820000000
0!
0*
09
0>
0C
#285830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#285840000000
0!
0*
09
0>
0C
#285850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#285860000000
0!
0*
09
0>
0C
#285870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#285880000000
0!
0*
09
0>
0C
#285890000000
1!
1*
b10 6
19
1>
1C
b10 G
#285900000000
0!
0*
09
0>
0C
#285910000000
1!
1*
b11 6
19
1>
1C
b11 G
#285920000000
0!
0*
09
0>
0C
#285930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#285940000000
0!
0*
09
0>
0C
#285950000000
1!
1*
b101 6
19
1>
1C
b101 G
#285960000000
0!
0*
09
0>
0C
#285970000000
1!
1*
b110 6
19
1>
1C
b110 G
#285980000000
0!
0*
09
0>
0C
#285990000000
1!
1*
b111 6
19
1>
1C
b111 G
#286000000000
0!
0*
09
0>
0C
#286010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#286020000000
0!
0*
09
0>
0C
#286030000000
1!
1*
b1 6
19
1>
1C
b1 G
#286040000000
0!
0*
09
0>
0C
#286050000000
1!
1*
b10 6
19
1>
1C
b10 G
#286060000000
0!
0*
09
0>
0C
#286070000000
1!
1*
b11 6
19
1>
1C
b11 G
#286080000000
0!
0*
09
0>
0C
#286090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#286100000000
0!
0*
09
0>
0C
#286110000000
1!
1*
b101 6
19
1>
1C
b101 G
#286120000000
0!
0*
09
0>
0C
#286130000000
1!
1*
b110 6
19
1>
1C
b110 G
#286140000000
0!
0*
09
0>
0C
#286150000000
1!
1*
b111 6
19
1>
1C
b111 G
#286160000000
0!
0*
09
0>
0C
#286170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#286180000000
0!
0*
09
0>
0C
#286190000000
1!
1*
b1 6
19
1>
1C
b1 G
#286200000000
0!
0*
09
0>
0C
#286210000000
1!
1*
b10 6
19
1>
1C
b10 G
#286220000000
0!
0*
09
0>
0C
#286230000000
1!
1*
b11 6
19
1>
1C
b11 G
#286240000000
0!
0*
09
0>
0C
#286250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#286260000000
0!
0*
09
0>
0C
#286270000000
1!
1*
b101 6
19
1>
1C
b101 G
#286280000000
0!
0*
09
0>
0C
#286290000000
1!
1*
b110 6
19
1>
1C
b110 G
#286300000000
0!
0*
09
0>
0C
#286310000000
1!
1*
b111 6
19
1>
1C
b111 G
#286320000000
0!
1"
0*
1+
09
1:
0>
0C
#286330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#286340000000
0!
0*
09
0>
0C
#286350000000
1!
1*
b1 6
19
1>
1C
b1 G
#286360000000
0!
0*
09
0>
0C
#286370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#286380000000
0!
0*
09
0>
0C
#286390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#286400000000
0!
0*
09
0>
0C
#286410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#286420000000
0!
0*
09
0>
0C
#286430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#286440000000
0!
0#
0*
0,
09
0>
0?
0C
#286450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#286460000000
0!
0*
09
0>
0C
#286470000000
1!
1*
19
1>
1C
#286480000000
0!
0*
09
0>
0C
#286490000000
1!
1*
19
1>
1C
#286500000000
0!
0*
09
0>
0C
#286510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#286520000000
0!
0*
09
0>
0C
#286530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#286540000000
0!
0*
09
0>
0C
#286550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#286560000000
0!
0*
09
0>
0C
#286570000000
1!
1*
b10 6
19
1>
1C
b10 G
#286580000000
0!
0*
09
0>
0C
#286590000000
1!
1*
b11 6
19
1>
1C
b11 G
#286600000000
0!
0*
09
0>
0C
#286610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#286620000000
0!
0*
09
0>
0C
#286630000000
1!
1*
b101 6
19
1>
1C
b101 G
#286640000000
0!
0*
09
0>
0C
#286650000000
1!
1*
b110 6
19
1>
1C
b110 G
#286660000000
0!
0*
09
0>
0C
#286670000000
1!
1*
b111 6
19
1>
1C
b111 G
#286680000000
0!
0*
09
0>
0C
#286690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#286700000000
0!
0*
09
0>
0C
#286710000000
1!
1*
b1 6
19
1>
1C
b1 G
#286720000000
0!
0*
09
0>
0C
#286730000000
1!
1*
b10 6
19
1>
1C
b10 G
#286740000000
0!
0*
09
0>
0C
#286750000000
1!
1*
b11 6
19
1>
1C
b11 G
#286760000000
0!
0*
09
0>
0C
#286770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#286780000000
0!
0*
09
0>
0C
#286790000000
1!
1*
b101 6
19
1>
1C
b101 G
#286800000000
0!
0*
09
0>
0C
#286810000000
1!
1*
b110 6
19
1>
1C
b110 G
#286820000000
0!
0*
09
0>
0C
#286830000000
1!
1*
b111 6
19
1>
1C
b111 G
#286840000000
0!
0*
09
0>
0C
#286850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#286860000000
0!
0*
09
0>
0C
#286870000000
1!
1*
b1 6
19
1>
1C
b1 G
#286880000000
0!
0*
09
0>
0C
#286890000000
1!
1*
b10 6
19
1>
1C
b10 G
#286900000000
0!
0*
09
0>
0C
#286910000000
1!
1*
b11 6
19
1>
1C
b11 G
#286920000000
0!
0*
09
0>
0C
#286930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#286940000000
0!
0*
09
0>
0C
#286950000000
1!
1*
b101 6
19
1>
1C
b101 G
#286960000000
0!
0*
09
0>
0C
#286970000000
1!
1*
b110 6
19
1>
1C
b110 G
#286980000000
0!
0*
09
0>
0C
#286990000000
1!
1*
b111 6
19
1>
1C
b111 G
#287000000000
0!
1"
0*
1+
09
1:
0>
0C
#287010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#287020000000
0!
0*
09
0>
0C
#287030000000
1!
1*
b1 6
19
1>
1C
b1 G
#287040000000
0!
0*
09
0>
0C
#287050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#287060000000
0!
0*
09
0>
0C
#287070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#287080000000
0!
0*
09
0>
0C
#287090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#287100000000
0!
0*
09
0>
0C
#287110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#287120000000
0!
0#
0*
0,
09
0>
0?
0C
#287130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#287140000000
0!
0*
09
0>
0C
#287150000000
1!
1*
19
1>
1C
#287160000000
0!
0*
09
0>
0C
#287170000000
1!
1*
19
1>
1C
#287180000000
0!
0*
09
0>
0C
#287190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#287200000000
0!
0*
09
0>
0C
#287210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#287220000000
0!
0*
09
0>
0C
#287230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#287240000000
0!
0*
09
0>
0C
#287250000000
1!
1*
b10 6
19
1>
1C
b10 G
#287260000000
0!
0*
09
0>
0C
#287270000000
1!
1*
b11 6
19
1>
1C
b11 G
#287280000000
0!
0*
09
0>
0C
#287290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#287300000000
0!
0*
09
0>
0C
#287310000000
1!
1*
b101 6
19
1>
1C
b101 G
#287320000000
0!
0*
09
0>
0C
#287330000000
1!
1*
b110 6
19
1>
1C
b110 G
#287340000000
0!
0*
09
0>
0C
#287350000000
1!
1*
b111 6
19
1>
1C
b111 G
#287360000000
0!
0*
09
0>
0C
#287370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#287380000000
0!
0*
09
0>
0C
#287390000000
1!
1*
b1 6
19
1>
1C
b1 G
#287400000000
0!
0*
09
0>
0C
#287410000000
1!
1*
b10 6
19
1>
1C
b10 G
#287420000000
0!
0*
09
0>
0C
#287430000000
1!
1*
b11 6
19
1>
1C
b11 G
#287440000000
0!
0*
09
0>
0C
#287450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#287460000000
0!
0*
09
0>
0C
#287470000000
1!
1*
b101 6
19
1>
1C
b101 G
#287480000000
0!
0*
09
0>
0C
#287490000000
1!
1*
b110 6
19
1>
1C
b110 G
#287500000000
0!
0*
09
0>
0C
#287510000000
1!
1*
b111 6
19
1>
1C
b111 G
#287520000000
0!
0*
09
0>
0C
#287530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#287540000000
0!
0*
09
0>
0C
#287550000000
1!
1*
b1 6
19
1>
1C
b1 G
#287560000000
0!
0*
09
0>
0C
#287570000000
1!
1*
b10 6
19
1>
1C
b10 G
#287580000000
0!
0*
09
0>
0C
#287590000000
1!
1*
b11 6
19
1>
1C
b11 G
#287600000000
0!
0*
09
0>
0C
#287610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#287620000000
0!
0*
09
0>
0C
#287630000000
1!
1*
b101 6
19
1>
1C
b101 G
#287640000000
0!
0*
09
0>
0C
#287650000000
1!
1*
b110 6
19
1>
1C
b110 G
#287660000000
0!
0*
09
0>
0C
#287670000000
1!
1*
b111 6
19
1>
1C
b111 G
#287680000000
0!
1"
0*
1+
09
1:
0>
0C
#287690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#287700000000
0!
0*
09
0>
0C
#287710000000
1!
1*
b1 6
19
1>
1C
b1 G
#287720000000
0!
0*
09
0>
0C
#287730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#287740000000
0!
0*
09
0>
0C
#287750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#287760000000
0!
0*
09
0>
0C
#287770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#287780000000
0!
0*
09
0>
0C
#287790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#287800000000
0!
0#
0*
0,
09
0>
0?
0C
#287810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#287820000000
0!
0*
09
0>
0C
#287830000000
1!
1*
19
1>
1C
#287840000000
0!
0*
09
0>
0C
#287850000000
1!
1*
19
1>
1C
#287860000000
0!
0*
09
0>
0C
#287870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#287880000000
0!
0*
09
0>
0C
#287890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#287900000000
0!
0*
09
0>
0C
#287910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#287920000000
0!
0*
09
0>
0C
#287930000000
1!
1*
b10 6
19
1>
1C
b10 G
#287940000000
0!
0*
09
0>
0C
#287950000000
1!
1*
b11 6
19
1>
1C
b11 G
#287960000000
0!
0*
09
0>
0C
#287970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#287980000000
0!
0*
09
0>
0C
#287990000000
1!
1*
b101 6
19
1>
1C
b101 G
#288000000000
0!
0*
09
0>
0C
#288010000000
1!
1*
b110 6
19
1>
1C
b110 G
#288020000000
0!
0*
09
0>
0C
#288030000000
1!
1*
b111 6
19
1>
1C
b111 G
#288040000000
0!
0*
09
0>
0C
#288050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#288060000000
0!
0*
09
0>
0C
#288070000000
1!
1*
b1 6
19
1>
1C
b1 G
#288080000000
0!
0*
09
0>
0C
#288090000000
1!
1*
b10 6
19
1>
1C
b10 G
#288100000000
0!
0*
09
0>
0C
#288110000000
1!
1*
b11 6
19
1>
1C
b11 G
#288120000000
0!
0*
09
0>
0C
#288130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#288140000000
0!
0*
09
0>
0C
#288150000000
1!
1*
b101 6
19
1>
1C
b101 G
#288160000000
0!
0*
09
0>
0C
#288170000000
1!
1*
b110 6
19
1>
1C
b110 G
#288180000000
0!
0*
09
0>
0C
#288190000000
1!
1*
b111 6
19
1>
1C
b111 G
#288200000000
0!
0*
09
0>
0C
#288210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#288220000000
0!
0*
09
0>
0C
#288230000000
1!
1*
b1 6
19
1>
1C
b1 G
#288240000000
0!
0*
09
0>
0C
#288250000000
1!
1*
b10 6
19
1>
1C
b10 G
#288260000000
0!
0*
09
0>
0C
#288270000000
1!
1*
b11 6
19
1>
1C
b11 G
#288280000000
0!
0*
09
0>
0C
#288290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#288300000000
0!
0*
09
0>
0C
#288310000000
1!
1*
b101 6
19
1>
1C
b101 G
#288320000000
0!
0*
09
0>
0C
#288330000000
1!
1*
b110 6
19
1>
1C
b110 G
#288340000000
0!
0*
09
0>
0C
#288350000000
1!
1*
b111 6
19
1>
1C
b111 G
#288360000000
0!
1"
0*
1+
09
1:
0>
0C
#288370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#288380000000
0!
0*
09
0>
0C
#288390000000
1!
1*
b1 6
19
1>
1C
b1 G
#288400000000
0!
0*
09
0>
0C
#288410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#288420000000
0!
0*
09
0>
0C
#288430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#288440000000
0!
0*
09
0>
0C
#288450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#288460000000
0!
0*
09
0>
0C
#288470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#288480000000
0!
0#
0*
0,
09
0>
0?
0C
#288490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#288500000000
0!
0*
09
0>
0C
#288510000000
1!
1*
19
1>
1C
#288520000000
0!
0*
09
0>
0C
#288530000000
1!
1*
19
1>
1C
#288540000000
0!
0*
09
0>
0C
#288550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#288560000000
0!
0*
09
0>
0C
#288570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#288580000000
0!
0*
09
0>
0C
#288590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#288600000000
0!
0*
09
0>
0C
#288610000000
1!
1*
b10 6
19
1>
1C
b10 G
#288620000000
0!
0*
09
0>
0C
#288630000000
1!
1*
b11 6
19
1>
1C
b11 G
#288640000000
0!
0*
09
0>
0C
#288650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#288660000000
0!
0*
09
0>
0C
#288670000000
1!
1*
b101 6
19
1>
1C
b101 G
#288680000000
0!
0*
09
0>
0C
#288690000000
1!
1*
b110 6
19
1>
1C
b110 G
#288700000000
0!
0*
09
0>
0C
#288710000000
1!
1*
b111 6
19
1>
1C
b111 G
#288720000000
0!
0*
09
0>
0C
#288730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#288740000000
0!
0*
09
0>
0C
#288750000000
1!
1*
b1 6
19
1>
1C
b1 G
#288760000000
0!
0*
09
0>
0C
#288770000000
1!
1*
b10 6
19
1>
1C
b10 G
#288780000000
0!
0*
09
0>
0C
#288790000000
1!
1*
b11 6
19
1>
1C
b11 G
#288800000000
0!
0*
09
0>
0C
#288810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#288820000000
0!
0*
09
0>
0C
#288830000000
1!
1*
b101 6
19
1>
1C
b101 G
#288840000000
0!
0*
09
0>
0C
#288850000000
1!
1*
b110 6
19
1>
1C
b110 G
#288860000000
0!
0*
09
0>
0C
#288870000000
1!
1*
b111 6
19
1>
1C
b111 G
#288880000000
0!
0*
09
0>
0C
#288890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#288900000000
0!
0*
09
0>
0C
#288910000000
1!
1*
b1 6
19
1>
1C
b1 G
#288920000000
0!
0*
09
0>
0C
#288930000000
1!
1*
b10 6
19
1>
1C
b10 G
#288940000000
0!
0*
09
0>
0C
#288950000000
1!
1*
b11 6
19
1>
1C
b11 G
#288960000000
0!
0*
09
0>
0C
#288970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#288980000000
0!
0*
09
0>
0C
#288990000000
1!
1*
b101 6
19
1>
1C
b101 G
#289000000000
0!
0*
09
0>
0C
#289010000000
1!
1*
b110 6
19
1>
1C
b110 G
#289020000000
0!
0*
09
0>
0C
#289030000000
1!
1*
b111 6
19
1>
1C
b111 G
#289040000000
0!
1"
0*
1+
09
1:
0>
0C
#289050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#289060000000
0!
0*
09
0>
0C
#289070000000
1!
1*
b1 6
19
1>
1C
b1 G
#289080000000
0!
0*
09
0>
0C
#289090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#289100000000
0!
0*
09
0>
0C
#289110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#289120000000
0!
0*
09
0>
0C
#289130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#289140000000
0!
0*
09
0>
0C
#289150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#289160000000
0!
0#
0*
0,
09
0>
0?
0C
#289170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#289180000000
0!
0*
09
0>
0C
#289190000000
1!
1*
19
1>
1C
#289200000000
0!
0*
09
0>
0C
#289210000000
1!
1*
19
1>
1C
#289220000000
0!
0*
09
0>
0C
#289230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#289240000000
0!
0*
09
0>
0C
#289250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#289260000000
0!
0*
09
0>
0C
#289270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#289280000000
0!
0*
09
0>
0C
#289290000000
1!
1*
b10 6
19
1>
1C
b10 G
#289300000000
0!
0*
09
0>
0C
#289310000000
1!
1*
b11 6
19
1>
1C
b11 G
#289320000000
0!
0*
09
0>
0C
#289330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#289340000000
0!
0*
09
0>
0C
#289350000000
1!
1*
b101 6
19
1>
1C
b101 G
#289360000000
0!
0*
09
0>
0C
#289370000000
1!
1*
b110 6
19
1>
1C
b110 G
#289380000000
0!
0*
09
0>
0C
#289390000000
1!
1*
b111 6
19
1>
1C
b111 G
#289400000000
0!
0*
09
0>
0C
#289410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#289420000000
0!
0*
09
0>
0C
#289430000000
1!
1*
b1 6
19
1>
1C
b1 G
#289440000000
0!
0*
09
0>
0C
#289450000000
1!
1*
b10 6
19
1>
1C
b10 G
#289460000000
0!
0*
09
0>
0C
#289470000000
1!
1*
b11 6
19
1>
1C
b11 G
#289480000000
0!
0*
09
0>
0C
#289490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#289500000000
0!
0*
09
0>
0C
#289510000000
1!
1*
b101 6
19
1>
1C
b101 G
#289520000000
0!
0*
09
0>
0C
#289530000000
1!
1*
b110 6
19
1>
1C
b110 G
#289540000000
0!
0*
09
0>
0C
#289550000000
1!
1*
b111 6
19
1>
1C
b111 G
#289560000000
0!
0*
09
0>
0C
#289570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#289580000000
0!
0*
09
0>
0C
#289590000000
1!
1*
b1 6
19
1>
1C
b1 G
#289600000000
0!
0*
09
0>
0C
#289610000000
1!
1*
b10 6
19
1>
1C
b10 G
#289620000000
0!
0*
09
0>
0C
#289630000000
1!
1*
b11 6
19
1>
1C
b11 G
#289640000000
0!
0*
09
0>
0C
#289650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#289660000000
0!
0*
09
0>
0C
#289670000000
1!
1*
b101 6
19
1>
1C
b101 G
#289680000000
0!
0*
09
0>
0C
#289690000000
1!
1*
b110 6
19
1>
1C
b110 G
#289700000000
0!
0*
09
0>
0C
#289710000000
1!
1*
b111 6
19
1>
1C
b111 G
#289720000000
0!
1"
0*
1+
09
1:
0>
0C
#289730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#289740000000
0!
0*
09
0>
0C
#289750000000
1!
1*
b1 6
19
1>
1C
b1 G
#289760000000
0!
0*
09
0>
0C
#289770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#289780000000
0!
0*
09
0>
0C
#289790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#289800000000
0!
0*
09
0>
0C
#289810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#289820000000
0!
0*
09
0>
0C
#289830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#289840000000
0!
0#
0*
0,
09
0>
0?
0C
#289850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#289860000000
0!
0*
09
0>
0C
#289870000000
1!
1*
19
1>
1C
#289880000000
0!
0*
09
0>
0C
#289890000000
1!
1*
19
1>
1C
#289900000000
0!
0*
09
0>
0C
#289910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#289920000000
0!
0*
09
0>
0C
#289930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#289940000000
0!
0*
09
0>
0C
#289950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#289960000000
0!
0*
09
0>
0C
#289970000000
1!
1*
b10 6
19
1>
1C
b10 G
#289980000000
0!
0*
09
0>
0C
#289990000000
1!
1*
b11 6
19
1>
1C
b11 G
#290000000000
0!
0*
09
0>
0C
#290010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#290020000000
0!
0*
09
0>
0C
#290030000000
1!
1*
b101 6
19
1>
1C
b101 G
#290040000000
0!
0*
09
0>
0C
#290050000000
1!
1*
b110 6
19
1>
1C
b110 G
#290060000000
0!
0*
09
0>
0C
#290070000000
1!
1*
b111 6
19
1>
1C
b111 G
#290080000000
0!
0*
09
0>
0C
#290090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#290100000000
0!
0*
09
0>
0C
#290110000000
1!
1*
b1 6
19
1>
1C
b1 G
#290120000000
0!
0*
09
0>
0C
#290130000000
1!
1*
b10 6
19
1>
1C
b10 G
#290140000000
0!
0*
09
0>
0C
#290150000000
1!
1*
b11 6
19
1>
1C
b11 G
#290160000000
0!
0*
09
0>
0C
#290170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#290180000000
0!
0*
09
0>
0C
#290190000000
1!
1*
b101 6
19
1>
1C
b101 G
#290200000000
0!
0*
09
0>
0C
#290210000000
1!
1*
b110 6
19
1>
1C
b110 G
#290220000000
0!
0*
09
0>
0C
#290230000000
1!
1*
b111 6
19
1>
1C
b111 G
#290240000000
0!
0*
09
0>
0C
#290250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#290260000000
0!
0*
09
0>
0C
#290270000000
1!
1*
b1 6
19
1>
1C
b1 G
#290280000000
0!
0*
09
0>
0C
#290290000000
1!
1*
b10 6
19
1>
1C
b10 G
#290300000000
0!
0*
09
0>
0C
#290310000000
1!
1*
b11 6
19
1>
1C
b11 G
#290320000000
0!
0*
09
0>
0C
#290330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#290340000000
0!
0*
09
0>
0C
#290350000000
1!
1*
b101 6
19
1>
1C
b101 G
#290360000000
0!
0*
09
0>
0C
#290370000000
1!
1*
b110 6
19
1>
1C
b110 G
#290380000000
0!
0*
09
0>
0C
#290390000000
1!
1*
b111 6
19
1>
1C
b111 G
#290400000000
0!
1"
0*
1+
09
1:
0>
0C
#290410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#290420000000
0!
0*
09
0>
0C
#290430000000
1!
1*
b1 6
19
1>
1C
b1 G
#290440000000
0!
0*
09
0>
0C
#290450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#290460000000
0!
0*
09
0>
0C
#290470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#290480000000
0!
0*
09
0>
0C
#290490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#290500000000
0!
0*
09
0>
0C
#290510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#290520000000
0!
0#
0*
0,
09
0>
0?
0C
#290530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#290540000000
0!
0*
09
0>
0C
#290550000000
1!
1*
19
1>
1C
#290560000000
0!
0*
09
0>
0C
#290570000000
1!
1*
19
1>
1C
#290580000000
0!
0*
09
0>
0C
#290590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#290600000000
0!
0*
09
0>
0C
#290610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#290620000000
0!
0*
09
0>
0C
#290630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#290640000000
0!
0*
09
0>
0C
#290650000000
1!
1*
b10 6
19
1>
1C
b10 G
#290660000000
0!
0*
09
0>
0C
#290670000000
1!
1*
b11 6
19
1>
1C
b11 G
#290680000000
0!
0*
09
0>
0C
#290690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#290700000000
0!
0*
09
0>
0C
#290710000000
1!
1*
b101 6
19
1>
1C
b101 G
#290720000000
0!
0*
09
0>
0C
#290730000000
1!
1*
b110 6
19
1>
1C
b110 G
#290740000000
0!
0*
09
0>
0C
#290750000000
1!
1*
b111 6
19
1>
1C
b111 G
#290760000000
0!
0*
09
0>
0C
#290770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#290780000000
0!
0*
09
0>
0C
#290790000000
1!
1*
b1 6
19
1>
1C
b1 G
#290800000000
0!
0*
09
0>
0C
#290810000000
1!
1*
b10 6
19
1>
1C
b10 G
#290820000000
0!
0*
09
0>
0C
#290830000000
1!
1*
b11 6
19
1>
1C
b11 G
#290840000000
0!
0*
09
0>
0C
#290850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#290860000000
0!
0*
09
0>
0C
#290870000000
1!
1*
b101 6
19
1>
1C
b101 G
#290880000000
0!
0*
09
0>
0C
#290890000000
1!
1*
b110 6
19
1>
1C
b110 G
#290900000000
0!
0*
09
0>
0C
#290910000000
1!
1*
b111 6
19
1>
1C
b111 G
#290920000000
0!
0*
09
0>
0C
#290930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#290940000000
0!
0*
09
0>
0C
#290950000000
1!
1*
b1 6
19
1>
1C
b1 G
#290960000000
0!
0*
09
0>
0C
#290970000000
1!
1*
b10 6
19
1>
1C
b10 G
#290980000000
0!
0*
09
0>
0C
#290990000000
1!
1*
b11 6
19
1>
1C
b11 G
#291000000000
0!
0*
09
0>
0C
#291010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#291020000000
0!
0*
09
0>
0C
#291030000000
1!
1*
b101 6
19
1>
1C
b101 G
#291040000000
0!
0*
09
0>
0C
#291050000000
1!
1*
b110 6
19
1>
1C
b110 G
#291060000000
0!
0*
09
0>
0C
#291070000000
1!
1*
b111 6
19
1>
1C
b111 G
#291080000000
0!
1"
0*
1+
09
1:
0>
0C
#291090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#291100000000
0!
0*
09
0>
0C
#291110000000
1!
1*
b1 6
19
1>
1C
b1 G
#291120000000
0!
0*
09
0>
0C
#291130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#291140000000
0!
0*
09
0>
0C
#291150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#291160000000
0!
0*
09
0>
0C
#291170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#291180000000
0!
0*
09
0>
0C
#291190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#291200000000
0!
0#
0*
0,
09
0>
0?
0C
#291210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#291220000000
0!
0*
09
0>
0C
#291230000000
1!
1*
19
1>
1C
#291240000000
0!
0*
09
0>
0C
#291250000000
1!
1*
19
1>
1C
#291260000000
0!
0*
09
0>
0C
#291270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#291280000000
0!
0*
09
0>
0C
#291290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#291300000000
0!
0*
09
0>
0C
#291310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#291320000000
0!
0*
09
0>
0C
#291330000000
1!
1*
b10 6
19
1>
1C
b10 G
#291340000000
0!
0*
09
0>
0C
#291350000000
1!
1*
b11 6
19
1>
1C
b11 G
#291360000000
0!
0*
09
0>
0C
#291370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#291380000000
0!
0*
09
0>
0C
#291390000000
1!
1*
b101 6
19
1>
1C
b101 G
#291400000000
0!
0*
09
0>
0C
#291410000000
1!
1*
b110 6
19
1>
1C
b110 G
#291420000000
0!
0*
09
0>
0C
#291430000000
1!
1*
b111 6
19
1>
1C
b111 G
#291440000000
0!
0*
09
0>
0C
#291450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#291460000000
0!
0*
09
0>
0C
#291470000000
1!
1*
b1 6
19
1>
1C
b1 G
#291480000000
0!
0*
09
0>
0C
#291490000000
1!
1*
b10 6
19
1>
1C
b10 G
#291500000000
0!
0*
09
0>
0C
#291510000000
1!
1*
b11 6
19
1>
1C
b11 G
#291520000000
0!
0*
09
0>
0C
#291530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#291540000000
0!
0*
09
0>
0C
#291550000000
1!
1*
b101 6
19
1>
1C
b101 G
#291560000000
0!
0*
09
0>
0C
#291570000000
1!
1*
b110 6
19
1>
1C
b110 G
#291580000000
0!
0*
09
0>
0C
#291590000000
1!
1*
b111 6
19
1>
1C
b111 G
#291600000000
0!
0*
09
0>
0C
#291610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#291620000000
0!
0*
09
0>
0C
#291630000000
1!
1*
b1 6
19
1>
1C
b1 G
#291640000000
0!
0*
09
0>
0C
#291650000000
1!
1*
b10 6
19
1>
1C
b10 G
#291660000000
0!
0*
09
0>
0C
#291670000000
1!
1*
b11 6
19
1>
1C
b11 G
#291680000000
0!
0*
09
0>
0C
#291690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#291700000000
0!
0*
09
0>
0C
#291710000000
1!
1*
b101 6
19
1>
1C
b101 G
#291720000000
0!
0*
09
0>
0C
#291730000000
1!
1*
b110 6
19
1>
1C
b110 G
#291740000000
0!
0*
09
0>
0C
#291750000000
1!
1*
b111 6
19
1>
1C
b111 G
#291760000000
0!
1"
0*
1+
09
1:
0>
0C
#291770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#291780000000
0!
0*
09
0>
0C
#291790000000
1!
1*
b1 6
19
1>
1C
b1 G
#291800000000
0!
0*
09
0>
0C
#291810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#291820000000
0!
0*
09
0>
0C
#291830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#291840000000
0!
0*
09
0>
0C
#291850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#291860000000
0!
0*
09
0>
0C
#291870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#291880000000
0!
0#
0*
0,
09
0>
0?
0C
#291890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#291900000000
0!
0*
09
0>
0C
#291910000000
1!
1*
19
1>
1C
#291920000000
0!
0*
09
0>
0C
#291930000000
1!
1*
19
1>
1C
#291940000000
0!
0*
09
0>
0C
#291950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#291960000000
0!
0*
09
0>
0C
#291970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#291980000000
0!
0*
09
0>
0C
#291990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#292000000000
0!
0*
09
0>
0C
#292010000000
1!
1*
b10 6
19
1>
1C
b10 G
#292020000000
0!
0*
09
0>
0C
#292030000000
1!
1*
b11 6
19
1>
1C
b11 G
#292040000000
0!
0*
09
0>
0C
#292050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#292060000000
0!
0*
09
0>
0C
#292070000000
1!
1*
b101 6
19
1>
1C
b101 G
#292080000000
0!
0*
09
0>
0C
#292090000000
1!
1*
b110 6
19
1>
1C
b110 G
#292100000000
0!
0*
09
0>
0C
#292110000000
1!
1*
b111 6
19
1>
1C
b111 G
#292120000000
0!
0*
09
0>
0C
#292130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#292140000000
0!
0*
09
0>
0C
#292150000000
1!
1*
b1 6
19
1>
1C
b1 G
#292160000000
0!
0*
09
0>
0C
#292170000000
1!
1*
b10 6
19
1>
1C
b10 G
#292180000000
0!
0*
09
0>
0C
#292190000000
1!
1*
b11 6
19
1>
1C
b11 G
#292200000000
0!
0*
09
0>
0C
#292210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#292220000000
0!
0*
09
0>
0C
#292230000000
1!
1*
b101 6
19
1>
1C
b101 G
#292240000000
0!
0*
09
0>
0C
#292250000000
1!
1*
b110 6
19
1>
1C
b110 G
#292260000000
0!
0*
09
0>
0C
#292270000000
1!
1*
b111 6
19
1>
1C
b111 G
#292280000000
0!
0*
09
0>
0C
#292290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#292300000000
0!
0*
09
0>
0C
#292310000000
1!
1*
b1 6
19
1>
1C
b1 G
#292320000000
0!
0*
09
0>
0C
#292330000000
1!
1*
b10 6
19
1>
1C
b10 G
#292340000000
0!
0*
09
0>
0C
#292350000000
1!
1*
b11 6
19
1>
1C
b11 G
#292360000000
0!
0*
09
0>
0C
#292370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#292380000000
0!
0*
09
0>
0C
#292390000000
1!
1*
b101 6
19
1>
1C
b101 G
#292400000000
0!
0*
09
0>
0C
#292410000000
1!
1*
b110 6
19
1>
1C
b110 G
#292420000000
0!
0*
09
0>
0C
#292430000000
1!
1*
b111 6
19
1>
1C
b111 G
#292440000000
0!
1"
0*
1+
09
1:
0>
0C
#292450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#292460000000
0!
0*
09
0>
0C
#292470000000
1!
1*
b1 6
19
1>
1C
b1 G
#292480000000
0!
0*
09
0>
0C
#292490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#292500000000
0!
0*
09
0>
0C
#292510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#292520000000
0!
0*
09
0>
0C
#292530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#292540000000
0!
0*
09
0>
0C
#292550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#292560000000
0!
0#
0*
0,
09
0>
0?
0C
#292570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#292580000000
0!
0*
09
0>
0C
#292590000000
1!
1*
19
1>
1C
#292600000000
0!
0*
09
0>
0C
#292610000000
1!
1*
19
1>
1C
#292620000000
0!
0*
09
0>
0C
#292630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#292640000000
0!
0*
09
0>
0C
#292650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#292660000000
0!
0*
09
0>
0C
#292670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#292680000000
0!
0*
09
0>
0C
#292690000000
1!
1*
b10 6
19
1>
1C
b10 G
#292700000000
0!
0*
09
0>
0C
#292710000000
1!
1*
b11 6
19
1>
1C
b11 G
#292720000000
0!
0*
09
0>
0C
#292730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#292740000000
0!
0*
09
0>
0C
#292750000000
1!
1*
b101 6
19
1>
1C
b101 G
#292760000000
0!
0*
09
0>
0C
#292770000000
1!
1*
b110 6
19
1>
1C
b110 G
#292780000000
0!
0*
09
0>
0C
#292790000000
1!
1*
b111 6
19
1>
1C
b111 G
#292800000000
0!
0*
09
0>
0C
#292810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#292820000000
0!
0*
09
0>
0C
#292830000000
1!
1*
b1 6
19
1>
1C
b1 G
#292840000000
0!
0*
09
0>
0C
#292850000000
1!
1*
b10 6
19
1>
1C
b10 G
#292860000000
0!
0*
09
0>
0C
#292870000000
1!
1*
b11 6
19
1>
1C
b11 G
#292880000000
0!
0*
09
0>
0C
#292890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#292900000000
0!
0*
09
0>
0C
#292910000000
1!
1*
b101 6
19
1>
1C
b101 G
#292920000000
0!
0*
09
0>
0C
#292930000000
1!
1*
b110 6
19
1>
1C
b110 G
#292940000000
0!
0*
09
0>
0C
#292950000000
1!
1*
b111 6
19
1>
1C
b111 G
#292960000000
0!
0*
09
0>
0C
#292970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#292980000000
0!
0*
09
0>
0C
#292990000000
1!
1*
b1 6
19
1>
1C
b1 G
#293000000000
0!
0*
09
0>
0C
#293010000000
1!
1*
b10 6
19
1>
1C
b10 G
#293020000000
0!
0*
09
0>
0C
#293030000000
1!
1*
b11 6
19
1>
1C
b11 G
#293040000000
0!
0*
09
0>
0C
#293050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#293060000000
0!
0*
09
0>
0C
#293070000000
1!
1*
b101 6
19
1>
1C
b101 G
#293080000000
0!
0*
09
0>
0C
#293090000000
1!
1*
b110 6
19
1>
1C
b110 G
#293100000000
0!
0*
09
0>
0C
#293110000000
1!
1*
b111 6
19
1>
1C
b111 G
#293120000000
0!
1"
0*
1+
09
1:
0>
0C
#293130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#293140000000
0!
0*
09
0>
0C
#293150000000
1!
1*
b1 6
19
1>
1C
b1 G
#293160000000
0!
0*
09
0>
0C
#293170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#293180000000
0!
0*
09
0>
0C
#293190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#293200000000
0!
0*
09
0>
0C
#293210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#293220000000
0!
0*
09
0>
0C
#293230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#293240000000
0!
0#
0*
0,
09
0>
0?
0C
#293250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#293260000000
0!
0*
09
0>
0C
#293270000000
1!
1*
19
1>
1C
#293280000000
0!
0*
09
0>
0C
#293290000000
1!
1*
19
1>
1C
#293300000000
0!
0*
09
0>
0C
#293310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#293320000000
0!
0*
09
0>
0C
#293330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#293340000000
0!
0*
09
0>
0C
#293350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#293360000000
0!
0*
09
0>
0C
#293370000000
1!
1*
b10 6
19
1>
1C
b10 G
#293380000000
0!
0*
09
0>
0C
#293390000000
1!
1*
b11 6
19
1>
1C
b11 G
#293400000000
0!
0*
09
0>
0C
#293410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#293420000000
0!
0*
09
0>
0C
#293430000000
1!
1*
b101 6
19
1>
1C
b101 G
#293440000000
0!
0*
09
0>
0C
#293450000000
1!
1*
b110 6
19
1>
1C
b110 G
#293460000000
0!
0*
09
0>
0C
#293470000000
1!
1*
b111 6
19
1>
1C
b111 G
#293480000000
0!
0*
09
0>
0C
#293490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#293500000000
0!
0*
09
0>
0C
#293510000000
1!
1*
b1 6
19
1>
1C
b1 G
#293520000000
0!
0*
09
0>
0C
#293530000000
1!
1*
b10 6
19
1>
1C
b10 G
#293540000000
0!
0*
09
0>
0C
#293550000000
1!
1*
b11 6
19
1>
1C
b11 G
#293560000000
0!
0*
09
0>
0C
#293570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#293580000000
0!
0*
09
0>
0C
#293590000000
1!
1*
b101 6
19
1>
1C
b101 G
#293600000000
0!
0*
09
0>
0C
#293610000000
1!
1*
b110 6
19
1>
1C
b110 G
#293620000000
0!
0*
09
0>
0C
#293630000000
1!
1*
b111 6
19
1>
1C
b111 G
#293640000000
0!
0*
09
0>
0C
#293650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#293660000000
0!
0*
09
0>
0C
#293670000000
1!
1*
b1 6
19
1>
1C
b1 G
#293680000000
0!
0*
09
0>
0C
#293690000000
1!
1*
b10 6
19
1>
1C
b10 G
#293700000000
0!
0*
09
0>
0C
#293710000000
1!
1*
b11 6
19
1>
1C
b11 G
#293720000000
0!
0*
09
0>
0C
#293730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#293740000000
0!
0*
09
0>
0C
#293750000000
1!
1*
b101 6
19
1>
1C
b101 G
#293760000000
0!
0*
09
0>
0C
#293770000000
1!
1*
b110 6
19
1>
1C
b110 G
#293780000000
0!
0*
09
0>
0C
#293790000000
1!
1*
b111 6
19
1>
1C
b111 G
#293800000000
0!
1"
0*
1+
09
1:
0>
0C
#293810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#293820000000
0!
0*
09
0>
0C
#293830000000
1!
1*
b1 6
19
1>
1C
b1 G
#293840000000
0!
0*
09
0>
0C
#293850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#293860000000
0!
0*
09
0>
0C
#293870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#293880000000
0!
0*
09
0>
0C
#293890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#293900000000
0!
0*
09
0>
0C
#293910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#293920000000
0!
0#
0*
0,
09
0>
0?
0C
#293930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#293940000000
0!
0*
09
0>
0C
#293950000000
1!
1*
19
1>
1C
#293960000000
0!
0*
09
0>
0C
#293970000000
1!
1*
19
1>
1C
#293980000000
0!
0*
09
0>
0C
#293990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#294000000000
0!
0*
09
0>
0C
#294010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#294020000000
0!
0*
09
0>
0C
#294030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#294040000000
0!
0*
09
0>
0C
#294050000000
1!
1*
b10 6
19
1>
1C
b10 G
#294060000000
0!
0*
09
0>
0C
#294070000000
1!
1*
b11 6
19
1>
1C
b11 G
#294080000000
0!
0*
09
0>
0C
#294090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#294100000000
0!
0*
09
0>
0C
#294110000000
1!
1*
b101 6
19
1>
1C
b101 G
#294120000000
0!
0*
09
0>
0C
#294130000000
1!
1*
b110 6
19
1>
1C
b110 G
#294140000000
0!
0*
09
0>
0C
#294150000000
1!
1*
b111 6
19
1>
1C
b111 G
#294160000000
0!
0*
09
0>
0C
#294170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#294180000000
0!
0*
09
0>
0C
#294190000000
1!
1*
b1 6
19
1>
1C
b1 G
#294200000000
0!
0*
09
0>
0C
#294210000000
1!
1*
b10 6
19
1>
1C
b10 G
#294220000000
0!
0*
09
0>
0C
#294230000000
1!
1*
b11 6
19
1>
1C
b11 G
#294240000000
0!
0*
09
0>
0C
#294250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#294260000000
0!
0*
09
0>
0C
#294270000000
1!
1*
b101 6
19
1>
1C
b101 G
#294280000000
0!
0*
09
0>
0C
#294290000000
1!
1*
b110 6
19
1>
1C
b110 G
#294300000000
0!
0*
09
0>
0C
#294310000000
1!
1*
b111 6
19
1>
1C
b111 G
#294320000000
0!
0*
09
0>
0C
#294330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#294340000000
0!
0*
09
0>
0C
#294350000000
1!
1*
b1 6
19
1>
1C
b1 G
#294360000000
0!
0*
09
0>
0C
#294370000000
1!
1*
b10 6
19
1>
1C
b10 G
#294380000000
0!
0*
09
0>
0C
#294390000000
1!
1*
b11 6
19
1>
1C
b11 G
#294400000000
0!
0*
09
0>
0C
#294410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#294420000000
0!
0*
09
0>
0C
#294430000000
1!
1*
b101 6
19
1>
1C
b101 G
#294440000000
0!
0*
09
0>
0C
#294450000000
1!
1*
b110 6
19
1>
1C
b110 G
#294460000000
0!
0*
09
0>
0C
#294470000000
1!
1*
b111 6
19
1>
1C
b111 G
#294480000000
0!
1"
0*
1+
09
1:
0>
0C
#294490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#294500000000
0!
0*
09
0>
0C
#294510000000
1!
1*
b1 6
19
1>
1C
b1 G
#294520000000
0!
0*
09
0>
0C
#294530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#294540000000
0!
0*
09
0>
0C
#294550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#294560000000
0!
0*
09
0>
0C
#294570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#294580000000
0!
0*
09
0>
0C
#294590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#294600000000
0!
0#
0*
0,
09
0>
0?
0C
#294610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#294620000000
0!
0*
09
0>
0C
#294630000000
1!
1*
19
1>
1C
#294640000000
0!
0*
09
0>
0C
#294650000000
1!
1*
19
1>
1C
#294660000000
0!
0*
09
0>
0C
#294670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#294680000000
0!
0*
09
0>
0C
#294690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#294700000000
0!
0*
09
0>
0C
#294710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#294720000000
0!
0*
09
0>
0C
#294730000000
1!
1*
b10 6
19
1>
1C
b10 G
#294740000000
0!
0*
09
0>
0C
#294750000000
1!
1*
b11 6
19
1>
1C
b11 G
#294760000000
0!
0*
09
0>
0C
#294770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#294780000000
0!
0*
09
0>
0C
#294790000000
1!
1*
b101 6
19
1>
1C
b101 G
#294800000000
0!
0*
09
0>
0C
#294810000000
1!
1*
b110 6
19
1>
1C
b110 G
#294820000000
0!
0*
09
0>
0C
#294830000000
1!
1*
b111 6
19
1>
1C
b111 G
#294840000000
0!
0*
09
0>
0C
#294850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#294860000000
0!
0*
09
0>
0C
#294870000000
1!
1*
b1 6
19
1>
1C
b1 G
#294880000000
0!
0*
09
0>
0C
#294890000000
1!
1*
b10 6
19
1>
1C
b10 G
#294900000000
0!
0*
09
0>
0C
#294910000000
1!
1*
b11 6
19
1>
1C
b11 G
#294920000000
0!
0*
09
0>
0C
#294930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#294940000000
0!
0*
09
0>
0C
#294950000000
1!
1*
b101 6
19
1>
1C
b101 G
#294960000000
0!
0*
09
0>
0C
#294970000000
1!
1*
b110 6
19
1>
1C
b110 G
#294980000000
0!
0*
09
0>
0C
#294990000000
1!
1*
b111 6
19
1>
1C
b111 G
#295000000000
0!
0*
09
0>
0C
#295010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#295020000000
0!
0*
09
0>
0C
#295030000000
1!
1*
b1 6
19
1>
1C
b1 G
#295040000000
0!
0*
09
0>
0C
#295050000000
1!
1*
b10 6
19
1>
1C
b10 G
#295060000000
0!
0*
09
0>
0C
#295070000000
1!
1*
b11 6
19
1>
1C
b11 G
#295080000000
0!
0*
09
0>
0C
#295090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#295100000000
0!
0*
09
0>
0C
#295110000000
1!
1*
b101 6
19
1>
1C
b101 G
#295120000000
0!
0*
09
0>
0C
#295130000000
1!
1*
b110 6
19
1>
1C
b110 G
#295140000000
0!
0*
09
0>
0C
#295150000000
1!
1*
b111 6
19
1>
1C
b111 G
#295160000000
0!
1"
0*
1+
09
1:
0>
0C
#295170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#295180000000
0!
0*
09
0>
0C
#295190000000
1!
1*
b1 6
19
1>
1C
b1 G
#295200000000
0!
0*
09
0>
0C
#295210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#295220000000
0!
0*
09
0>
0C
#295230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#295240000000
0!
0*
09
0>
0C
#295250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#295260000000
0!
0*
09
0>
0C
#295270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#295280000000
0!
0#
0*
0,
09
0>
0?
0C
#295290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#295300000000
0!
0*
09
0>
0C
#295310000000
1!
1*
19
1>
1C
#295320000000
0!
0*
09
0>
0C
#295330000000
1!
1*
19
1>
1C
#295340000000
0!
0*
09
0>
0C
#295350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#295360000000
0!
0*
09
0>
0C
#295370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#295380000000
0!
0*
09
0>
0C
#295390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#295400000000
0!
0*
09
0>
0C
#295410000000
1!
1*
b10 6
19
1>
1C
b10 G
#295420000000
0!
0*
09
0>
0C
#295430000000
1!
1*
b11 6
19
1>
1C
b11 G
#295440000000
0!
0*
09
0>
0C
#295450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#295460000000
0!
0*
09
0>
0C
#295470000000
1!
1*
b101 6
19
1>
1C
b101 G
#295480000000
0!
0*
09
0>
0C
#295490000000
1!
1*
b110 6
19
1>
1C
b110 G
#295500000000
0!
0*
09
0>
0C
#295510000000
1!
1*
b111 6
19
1>
1C
b111 G
#295520000000
0!
0*
09
0>
0C
#295530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#295540000000
0!
0*
09
0>
0C
#295550000000
1!
1*
b1 6
19
1>
1C
b1 G
#295560000000
0!
0*
09
0>
0C
#295570000000
1!
1*
b10 6
19
1>
1C
b10 G
#295580000000
0!
0*
09
0>
0C
#295590000000
1!
1*
b11 6
19
1>
1C
b11 G
#295600000000
0!
0*
09
0>
0C
#295610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#295620000000
0!
0*
09
0>
0C
#295630000000
1!
1*
b101 6
19
1>
1C
b101 G
#295640000000
0!
0*
09
0>
0C
#295650000000
1!
1*
b110 6
19
1>
1C
b110 G
#295660000000
0!
0*
09
0>
0C
#295670000000
1!
1*
b111 6
19
1>
1C
b111 G
#295680000000
0!
0*
09
0>
0C
#295690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#295700000000
0!
0*
09
0>
0C
#295710000000
1!
1*
b1 6
19
1>
1C
b1 G
#295720000000
0!
0*
09
0>
0C
#295730000000
1!
1*
b10 6
19
1>
1C
b10 G
#295740000000
0!
0*
09
0>
0C
#295750000000
1!
1*
b11 6
19
1>
1C
b11 G
#295760000000
0!
0*
09
0>
0C
#295770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#295780000000
0!
0*
09
0>
0C
#295790000000
1!
1*
b101 6
19
1>
1C
b101 G
#295800000000
0!
0*
09
0>
0C
#295810000000
1!
1*
b110 6
19
1>
1C
b110 G
#295820000000
0!
0*
09
0>
0C
#295830000000
1!
1*
b111 6
19
1>
1C
b111 G
#295840000000
0!
1"
0*
1+
09
1:
0>
0C
#295850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#295860000000
0!
0*
09
0>
0C
#295870000000
1!
1*
b1 6
19
1>
1C
b1 G
#295880000000
0!
0*
09
0>
0C
#295890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#295900000000
0!
0*
09
0>
0C
#295910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#295920000000
0!
0*
09
0>
0C
#295930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#295940000000
0!
0*
09
0>
0C
#295950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#295960000000
0!
0#
0*
0,
09
0>
0?
0C
#295970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#295980000000
0!
0*
09
0>
0C
#295990000000
1!
1*
19
1>
1C
#296000000000
0!
0*
09
0>
0C
#296010000000
1!
1*
19
1>
1C
#296020000000
0!
0*
09
0>
0C
#296030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#296040000000
0!
0*
09
0>
0C
#296050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#296060000000
0!
0*
09
0>
0C
#296070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#296080000000
0!
0*
09
0>
0C
#296090000000
1!
1*
b10 6
19
1>
1C
b10 G
#296100000000
0!
0*
09
0>
0C
#296110000000
1!
1*
b11 6
19
1>
1C
b11 G
#296120000000
0!
0*
09
0>
0C
#296130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#296140000000
0!
0*
09
0>
0C
#296150000000
1!
1*
b101 6
19
1>
1C
b101 G
#296160000000
0!
0*
09
0>
0C
#296170000000
1!
1*
b110 6
19
1>
1C
b110 G
#296180000000
0!
0*
09
0>
0C
#296190000000
1!
1*
b111 6
19
1>
1C
b111 G
#296200000000
0!
0*
09
0>
0C
#296210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#296220000000
0!
0*
09
0>
0C
#296230000000
1!
1*
b1 6
19
1>
1C
b1 G
#296240000000
0!
0*
09
0>
0C
#296250000000
1!
1*
b10 6
19
1>
1C
b10 G
#296260000000
0!
0*
09
0>
0C
#296270000000
1!
1*
b11 6
19
1>
1C
b11 G
#296280000000
0!
0*
09
0>
0C
#296290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#296300000000
0!
0*
09
0>
0C
#296310000000
1!
1*
b101 6
19
1>
1C
b101 G
#296320000000
0!
0*
09
0>
0C
#296330000000
1!
1*
b110 6
19
1>
1C
b110 G
#296340000000
0!
0*
09
0>
0C
#296350000000
1!
1*
b111 6
19
1>
1C
b111 G
#296360000000
0!
0*
09
0>
0C
#296370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#296380000000
0!
0*
09
0>
0C
#296390000000
1!
1*
b1 6
19
1>
1C
b1 G
#296400000000
0!
0*
09
0>
0C
#296410000000
1!
1*
b10 6
19
1>
1C
b10 G
#296420000000
0!
0*
09
0>
0C
#296430000000
1!
1*
b11 6
19
1>
1C
b11 G
#296440000000
0!
0*
09
0>
0C
#296450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#296460000000
0!
0*
09
0>
0C
#296470000000
1!
1*
b101 6
19
1>
1C
b101 G
#296480000000
0!
0*
09
0>
0C
#296490000000
1!
1*
b110 6
19
1>
1C
b110 G
#296500000000
0!
0*
09
0>
0C
#296510000000
1!
1*
b111 6
19
1>
1C
b111 G
#296520000000
0!
1"
0*
1+
09
1:
0>
0C
#296530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#296540000000
0!
0*
09
0>
0C
#296550000000
1!
1*
b1 6
19
1>
1C
b1 G
#296560000000
0!
0*
09
0>
0C
#296570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#296580000000
0!
0*
09
0>
0C
#296590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#296600000000
0!
0*
09
0>
0C
#296610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#296620000000
0!
0*
09
0>
0C
#296630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#296640000000
0!
0#
0*
0,
09
0>
0?
0C
#296650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#296660000000
0!
0*
09
0>
0C
#296670000000
1!
1*
19
1>
1C
#296680000000
0!
0*
09
0>
0C
#296690000000
1!
1*
19
1>
1C
#296700000000
0!
0*
09
0>
0C
#296710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#296720000000
0!
0*
09
0>
0C
#296730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#296740000000
0!
0*
09
0>
0C
#296750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#296760000000
0!
0*
09
0>
0C
#296770000000
1!
1*
b10 6
19
1>
1C
b10 G
#296780000000
0!
0*
09
0>
0C
#296790000000
1!
1*
b11 6
19
1>
1C
b11 G
#296800000000
0!
0*
09
0>
0C
#296810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#296820000000
0!
0*
09
0>
0C
#296830000000
1!
1*
b101 6
19
1>
1C
b101 G
#296840000000
0!
0*
09
0>
0C
#296850000000
1!
1*
b110 6
19
1>
1C
b110 G
#296860000000
0!
0*
09
0>
0C
#296870000000
1!
1*
b111 6
19
1>
1C
b111 G
#296880000000
0!
0*
09
0>
0C
#296890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#296900000000
0!
0*
09
0>
0C
#296910000000
1!
1*
b1 6
19
1>
1C
b1 G
#296920000000
0!
0*
09
0>
0C
#296930000000
1!
1*
b10 6
19
1>
1C
b10 G
#296940000000
0!
0*
09
0>
0C
#296950000000
1!
1*
b11 6
19
1>
1C
b11 G
#296960000000
0!
0*
09
0>
0C
#296970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#296980000000
0!
0*
09
0>
0C
#296990000000
1!
1*
b101 6
19
1>
1C
b101 G
#297000000000
0!
0*
09
0>
0C
#297010000000
1!
1*
b110 6
19
1>
1C
b110 G
#297020000000
0!
0*
09
0>
0C
#297030000000
1!
1*
b111 6
19
1>
1C
b111 G
#297040000000
0!
0*
09
0>
0C
#297050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#297060000000
0!
0*
09
0>
0C
#297070000000
1!
1*
b1 6
19
1>
1C
b1 G
#297080000000
0!
0*
09
0>
0C
#297090000000
1!
1*
b10 6
19
1>
1C
b10 G
#297100000000
0!
0*
09
0>
0C
#297110000000
1!
1*
b11 6
19
1>
1C
b11 G
#297120000000
0!
0*
09
0>
0C
#297130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#297140000000
0!
0*
09
0>
0C
#297150000000
1!
1*
b101 6
19
1>
1C
b101 G
#297160000000
0!
0*
09
0>
0C
#297170000000
1!
1*
b110 6
19
1>
1C
b110 G
#297180000000
0!
0*
09
0>
0C
#297190000000
1!
1*
b111 6
19
1>
1C
b111 G
#297200000000
0!
1"
0*
1+
09
1:
0>
0C
#297210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#297220000000
0!
0*
09
0>
0C
#297230000000
1!
1*
b1 6
19
1>
1C
b1 G
#297240000000
0!
0*
09
0>
0C
#297250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#297260000000
0!
0*
09
0>
0C
#297270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#297280000000
0!
0*
09
0>
0C
#297290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#297300000000
0!
0*
09
0>
0C
#297310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#297320000000
0!
0#
0*
0,
09
0>
0?
0C
#297330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#297340000000
0!
0*
09
0>
0C
#297350000000
1!
1*
19
1>
1C
#297360000000
0!
0*
09
0>
0C
#297370000000
1!
1*
19
1>
1C
#297380000000
0!
0*
09
0>
0C
#297390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#297400000000
0!
0*
09
0>
0C
#297410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#297420000000
0!
0*
09
0>
0C
#297430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#297440000000
0!
0*
09
0>
0C
#297450000000
1!
1*
b10 6
19
1>
1C
b10 G
#297460000000
0!
0*
09
0>
0C
#297470000000
1!
1*
b11 6
19
1>
1C
b11 G
#297480000000
0!
0*
09
0>
0C
#297490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#297500000000
0!
0*
09
0>
0C
#297510000000
1!
1*
b101 6
19
1>
1C
b101 G
#297520000000
0!
0*
09
0>
0C
#297530000000
1!
1*
b110 6
19
1>
1C
b110 G
#297540000000
0!
0*
09
0>
0C
#297550000000
1!
1*
b111 6
19
1>
1C
b111 G
#297560000000
0!
0*
09
0>
0C
#297570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#297580000000
0!
0*
09
0>
0C
#297590000000
1!
1*
b1 6
19
1>
1C
b1 G
#297600000000
0!
0*
09
0>
0C
#297610000000
1!
1*
b10 6
19
1>
1C
b10 G
#297620000000
0!
0*
09
0>
0C
#297630000000
1!
1*
b11 6
19
1>
1C
b11 G
#297640000000
0!
0*
09
0>
0C
#297650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#297660000000
0!
0*
09
0>
0C
#297670000000
1!
1*
b101 6
19
1>
1C
b101 G
#297680000000
0!
0*
09
0>
0C
#297690000000
1!
1*
b110 6
19
1>
1C
b110 G
#297700000000
0!
0*
09
0>
0C
#297710000000
1!
1*
b111 6
19
1>
1C
b111 G
#297720000000
0!
0*
09
0>
0C
#297730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#297740000000
0!
0*
09
0>
0C
#297750000000
1!
1*
b1 6
19
1>
1C
b1 G
#297760000000
0!
0*
09
0>
0C
#297770000000
1!
1*
b10 6
19
1>
1C
b10 G
#297780000000
0!
0*
09
0>
0C
#297790000000
1!
1*
b11 6
19
1>
1C
b11 G
#297800000000
0!
0*
09
0>
0C
#297810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#297820000000
0!
0*
09
0>
0C
#297830000000
1!
1*
b101 6
19
1>
1C
b101 G
#297840000000
0!
0*
09
0>
0C
#297850000000
1!
1*
b110 6
19
1>
1C
b110 G
#297860000000
0!
0*
09
0>
0C
#297870000000
1!
1*
b111 6
19
1>
1C
b111 G
#297880000000
0!
1"
0*
1+
09
1:
0>
0C
#297890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#297900000000
0!
0*
09
0>
0C
#297910000000
1!
1*
b1 6
19
1>
1C
b1 G
#297920000000
0!
0*
09
0>
0C
#297930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#297940000000
0!
0*
09
0>
0C
#297950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#297960000000
0!
0*
09
0>
0C
#297970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#297980000000
0!
0*
09
0>
0C
#297990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#298000000000
0!
0#
0*
0,
09
0>
0?
0C
#298010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#298020000000
0!
0*
09
0>
0C
#298030000000
1!
1*
19
1>
1C
#298040000000
0!
0*
09
0>
0C
#298050000000
1!
1*
19
1>
1C
#298060000000
0!
0*
09
0>
0C
#298070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#298080000000
0!
0*
09
0>
0C
#298090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#298100000000
0!
0*
09
0>
0C
#298110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#298120000000
0!
0*
09
0>
0C
#298130000000
1!
1*
b10 6
19
1>
1C
b10 G
#298140000000
0!
0*
09
0>
0C
#298150000000
1!
1*
b11 6
19
1>
1C
b11 G
#298160000000
0!
0*
09
0>
0C
#298170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#298180000000
0!
0*
09
0>
0C
#298190000000
1!
1*
b101 6
19
1>
1C
b101 G
#298200000000
0!
0*
09
0>
0C
#298210000000
1!
1*
b110 6
19
1>
1C
b110 G
#298220000000
0!
0*
09
0>
0C
#298230000000
1!
1*
b111 6
19
1>
1C
b111 G
#298240000000
0!
0*
09
0>
0C
#298250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#298260000000
0!
0*
09
0>
0C
#298270000000
1!
1*
b1 6
19
1>
1C
b1 G
#298280000000
0!
0*
09
0>
0C
#298290000000
1!
1*
b10 6
19
1>
1C
b10 G
#298300000000
0!
0*
09
0>
0C
#298310000000
1!
1*
b11 6
19
1>
1C
b11 G
#298320000000
0!
0*
09
0>
0C
#298330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#298340000000
0!
0*
09
0>
0C
#298350000000
1!
1*
b101 6
19
1>
1C
b101 G
#298360000000
0!
0*
09
0>
0C
#298370000000
1!
1*
b110 6
19
1>
1C
b110 G
#298380000000
0!
0*
09
0>
0C
#298390000000
1!
1*
b111 6
19
1>
1C
b111 G
#298400000000
0!
0*
09
0>
0C
#298410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#298420000000
0!
0*
09
0>
0C
#298430000000
1!
1*
b1 6
19
1>
1C
b1 G
#298440000000
0!
0*
09
0>
0C
#298450000000
1!
1*
b10 6
19
1>
1C
b10 G
#298460000000
0!
0*
09
0>
0C
#298470000000
1!
1*
b11 6
19
1>
1C
b11 G
#298480000000
0!
0*
09
0>
0C
#298490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#298500000000
0!
0*
09
0>
0C
#298510000000
1!
1*
b101 6
19
1>
1C
b101 G
#298520000000
0!
0*
09
0>
0C
#298530000000
1!
1*
b110 6
19
1>
1C
b110 G
#298540000000
0!
0*
09
0>
0C
#298550000000
1!
1*
b111 6
19
1>
1C
b111 G
#298560000000
0!
1"
0*
1+
09
1:
0>
0C
#298570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#298580000000
0!
0*
09
0>
0C
#298590000000
1!
1*
b1 6
19
1>
1C
b1 G
#298600000000
0!
0*
09
0>
0C
#298610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#298620000000
0!
0*
09
0>
0C
#298630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#298640000000
0!
0*
09
0>
0C
#298650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#298660000000
0!
0*
09
0>
0C
#298670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#298680000000
0!
0#
0*
0,
09
0>
0?
0C
#298690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#298700000000
0!
0*
09
0>
0C
#298710000000
1!
1*
19
1>
1C
#298720000000
0!
0*
09
0>
0C
#298730000000
1!
1*
19
1>
1C
#298740000000
0!
0*
09
0>
0C
#298750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#298760000000
0!
0*
09
0>
0C
#298770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#298780000000
0!
0*
09
0>
0C
#298790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#298800000000
0!
0*
09
0>
0C
#298810000000
1!
1*
b10 6
19
1>
1C
b10 G
#298820000000
0!
0*
09
0>
0C
#298830000000
1!
1*
b11 6
19
1>
1C
b11 G
#298840000000
0!
0*
09
0>
0C
#298850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#298860000000
0!
0*
09
0>
0C
#298870000000
1!
1*
b101 6
19
1>
1C
b101 G
#298880000000
0!
0*
09
0>
0C
#298890000000
1!
1*
b110 6
19
1>
1C
b110 G
#298900000000
0!
0*
09
0>
0C
#298910000000
1!
1*
b111 6
19
1>
1C
b111 G
#298920000000
0!
0*
09
0>
0C
#298930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#298940000000
0!
0*
09
0>
0C
#298950000000
1!
1*
b1 6
19
1>
1C
b1 G
#298960000000
0!
0*
09
0>
0C
#298970000000
1!
1*
b10 6
19
1>
1C
b10 G
#298980000000
0!
0*
09
0>
0C
#298990000000
1!
1*
b11 6
19
1>
1C
b11 G
#299000000000
0!
0*
09
0>
0C
#299010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#299020000000
0!
0*
09
0>
0C
#299030000000
1!
1*
b101 6
19
1>
1C
b101 G
#299040000000
0!
0*
09
0>
0C
#299050000000
1!
1*
b110 6
19
1>
1C
b110 G
#299060000000
0!
0*
09
0>
0C
#299070000000
1!
1*
b111 6
19
1>
1C
b111 G
#299080000000
0!
0*
09
0>
0C
#299090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#299100000000
0!
0*
09
0>
0C
#299110000000
1!
1*
b1 6
19
1>
1C
b1 G
#299120000000
0!
0*
09
0>
0C
#299130000000
1!
1*
b10 6
19
1>
1C
b10 G
#299140000000
0!
0*
09
0>
0C
#299150000000
1!
1*
b11 6
19
1>
1C
b11 G
#299160000000
0!
0*
09
0>
0C
#299170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#299180000000
0!
0*
09
0>
0C
#299190000000
1!
1*
b101 6
19
1>
1C
b101 G
#299200000000
0!
0*
09
0>
0C
#299210000000
1!
1*
b110 6
19
1>
1C
b110 G
#299220000000
0!
0*
09
0>
0C
#299230000000
1!
1*
b111 6
19
1>
1C
b111 G
#299240000000
0!
1"
0*
1+
09
1:
0>
0C
#299250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#299260000000
0!
0*
09
0>
0C
#299270000000
1!
1*
b1 6
19
1>
1C
b1 G
#299280000000
0!
0*
09
0>
0C
#299290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#299300000000
0!
0*
09
0>
0C
#299310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#299320000000
0!
0*
09
0>
0C
#299330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#299340000000
0!
0*
09
0>
0C
#299350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#299360000000
0!
0#
0*
0,
09
0>
0?
0C
#299370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#299380000000
0!
0*
09
0>
0C
#299390000000
1!
1*
19
1>
1C
#299400000000
0!
0*
09
0>
0C
#299410000000
1!
1*
19
1>
1C
#299420000000
0!
0*
09
0>
0C
#299430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#299440000000
0!
0*
09
0>
0C
#299450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#299460000000
0!
0*
09
0>
0C
#299470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#299480000000
0!
0*
09
0>
0C
#299490000000
1!
1*
b10 6
19
1>
1C
b10 G
#299500000000
0!
0*
09
0>
0C
#299510000000
1!
1*
b11 6
19
1>
1C
b11 G
#299520000000
0!
0*
09
0>
0C
#299530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#299540000000
0!
0*
09
0>
0C
#299550000000
1!
1*
b101 6
19
1>
1C
b101 G
#299560000000
0!
0*
09
0>
0C
#299570000000
1!
1*
b110 6
19
1>
1C
b110 G
#299580000000
0!
0*
09
0>
0C
#299590000000
1!
1*
b111 6
19
1>
1C
b111 G
#299600000000
0!
0*
09
0>
0C
#299610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#299620000000
0!
0*
09
0>
0C
#299630000000
1!
1*
b1 6
19
1>
1C
b1 G
#299640000000
0!
0*
09
0>
0C
#299650000000
1!
1*
b10 6
19
1>
1C
b10 G
#299660000000
0!
0*
09
0>
0C
#299670000000
1!
1*
b11 6
19
1>
1C
b11 G
#299680000000
0!
0*
09
0>
0C
#299690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#299700000000
0!
0*
09
0>
0C
#299710000000
1!
1*
b101 6
19
1>
1C
b101 G
#299720000000
0!
0*
09
0>
0C
#299730000000
1!
1*
b110 6
19
1>
1C
b110 G
#299740000000
0!
0*
09
0>
0C
#299750000000
1!
1*
b111 6
19
1>
1C
b111 G
#299760000000
0!
0*
09
0>
0C
#299770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#299780000000
0!
0*
09
0>
0C
#299790000000
1!
1*
b1 6
19
1>
1C
b1 G
#299800000000
0!
0*
09
0>
0C
#299810000000
1!
1*
b10 6
19
1>
1C
b10 G
#299820000000
0!
0*
09
0>
0C
#299830000000
1!
1*
b11 6
19
1>
1C
b11 G
#299840000000
0!
0*
09
0>
0C
#299850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#299860000000
0!
0*
09
0>
0C
#299870000000
1!
1*
b101 6
19
1>
1C
b101 G
#299880000000
0!
0*
09
0>
0C
#299890000000
1!
1*
b110 6
19
1>
1C
b110 G
#299900000000
0!
0*
09
0>
0C
#299910000000
1!
1*
b111 6
19
1>
1C
b111 G
#299920000000
0!
1"
0*
1+
09
1:
0>
0C
#299930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#299940000000
0!
0*
09
0>
0C
#299950000000
1!
1*
b1 6
19
1>
1C
b1 G
#299960000000
0!
0*
09
0>
0C
#299970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#299980000000
0!
0*
09
0>
0C
#299990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#300000000000
0!
0*
09
0>
0C
#300010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#300020000000
0!
0*
09
0>
0C
#300030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#300040000000
0!
0#
0*
0,
09
0>
0?
0C
#300050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#300060000000
0!
0*
09
0>
0C
#300070000000
1!
1*
19
1>
1C
#300080000000
0!
0*
09
0>
0C
#300090000000
1!
1*
19
1>
1C
#300100000000
0!
0*
09
0>
0C
#300110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#300120000000
0!
0*
09
0>
0C
#300130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#300140000000
0!
0*
09
0>
0C
#300150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#300160000000
0!
0*
09
0>
0C
#300170000000
1!
1*
b10 6
19
1>
1C
b10 G
#300180000000
0!
0*
09
0>
0C
#300190000000
1!
1*
b11 6
19
1>
1C
b11 G
#300200000000
0!
0*
09
0>
0C
#300210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#300220000000
0!
0*
09
0>
0C
#300230000000
1!
1*
b101 6
19
1>
1C
b101 G
#300240000000
0!
0*
09
0>
0C
#300250000000
1!
1*
b110 6
19
1>
1C
b110 G
#300260000000
0!
0*
09
0>
0C
#300270000000
1!
1*
b111 6
19
1>
1C
b111 G
#300280000000
0!
0*
09
0>
0C
#300290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#300300000000
0!
0*
09
0>
0C
#300310000000
1!
1*
b1 6
19
1>
1C
b1 G
#300320000000
0!
0*
09
0>
0C
#300330000000
1!
1*
b10 6
19
1>
1C
b10 G
#300340000000
0!
0*
09
0>
0C
#300350000000
1!
1*
b11 6
19
1>
1C
b11 G
#300360000000
0!
0*
09
0>
0C
#300370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#300380000000
0!
0*
09
0>
0C
#300390000000
1!
1*
b101 6
19
1>
1C
b101 G
#300400000000
0!
0*
09
0>
0C
#300410000000
1!
1*
b110 6
19
1>
1C
b110 G
#300420000000
0!
0*
09
0>
0C
#300430000000
1!
1*
b111 6
19
1>
1C
b111 G
#300440000000
0!
0*
09
0>
0C
#300450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#300460000000
0!
0*
09
0>
0C
#300470000000
1!
1*
b1 6
19
1>
1C
b1 G
#300480000000
0!
0*
09
0>
0C
#300490000000
1!
1*
b10 6
19
1>
1C
b10 G
#300500000000
0!
0*
09
0>
0C
#300510000000
1!
1*
b11 6
19
1>
1C
b11 G
#300520000000
0!
0*
09
0>
0C
#300530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#300540000000
0!
0*
09
0>
0C
#300550000000
1!
1*
b101 6
19
1>
1C
b101 G
#300560000000
0!
0*
09
0>
0C
#300570000000
1!
1*
b110 6
19
1>
1C
b110 G
#300580000000
0!
0*
09
0>
0C
#300590000000
1!
1*
b111 6
19
1>
1C
b111 G
#300600000000
0!
1"
0*
1+
09
1:
0>
0C
#300610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#300620000000
0!
0*
09
0>
0C
#300630000000
1!
1*
b1 6
19
1>
1C
b1 G
#300640000000
0!
0*
09
0>
0C
#300650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#300660000000
0!
0*
09
0>
0C
#300670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#300680000000
0!
0*
09
0>
0C
#300690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#300700000000
0!
0*
09
0>
0C
#300710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#300720000000
0!
0#
0*
0,
09
0>
0?
0C
#300730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#300740000000
0!
0*
09
0>
0C
#300750000000
1!
1*
19
1>
1C
#300760000000
0!
0*
09
0>
0C
#300770000000
1!
1*
19
1>
1C
#300780000000
0!
0*
09
0>
0C
#300790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#300800000000
0!
0*
09
0>
0C
#300810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#300820000000
0!
0*
09
0>
0C
#300830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#300840000000
0!
0*
09
0>
0C
#300850000000
1!
1*
b10 6
19
1>
1C
b10 G
#300860000000
0!
0*
09
0>
0C
#300870000000
1!
1*
b11 6
19
1>
1C
b11 G
#300880000000
0!
0*
09
0>
0C
#300890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#300900000000
0!
0*
09
0>
0C
#300910000000
1!
1*
b101 6
19
1>
1C
b101 G
#300920000000
0!
0*
09
0>
0C
#300930000000
1!
1*
b110 6
19
1>
1C
b110 G
#300940000000
0!
0*
09
0>
0C
#300950000000
1!
1*
b111 6
19
1>
1C
b111 G
#300960000000
0!
0*
09
0>
0C
#300970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#300980000000
0!
0*
09
0>
0C
#300990000000
1!
1*
b1 6
19
1>
1C
b1 G
#301000000000
0!
0*
09
0>
0C
#301010000000
1!
1*
b10 6
19
1>
1C
b10 G
#301020000000
0!
0*
09
0>
0C
#301030000000
1!
1*
b11 6
19
1>
1C
b11 G
#301040000000
0!
0*
09
0>
0C
#301050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#301060000000
0!
0*
09
0>
0C
#301070000000
1!
1*
b101 6
19
1>
1C
b101 G
#301080000000
0!
0*
09
0>
0C
#301090000000
1!
1*
b110 6
19
1>
1C
b110 G
#301100000000
0!
0*
09
0>
0C
#301110000000
1!
1*
b111 6
19
1>
1C
b111 G
#301120000000
0!
0*
09
0>
0C
#301130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#301140000000
0!
0*
09
0>
0C
#301150000000
1!
1*
b1 6
19
1>
1C
b1 G
#301160000000
0!
0*
09
0>
0C
#301170000000
1!
1*
b10 6
19
1>
1C
b10 G
#301180000000
0!
0*
09
0>
0C
#301190000000
1!
1*
b11 6
19
1>
1C
b11 G
#301200000000
0!
0*
09
0>
0C
#301210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#301220000000
0!
0*
09
0>
0C
#301230000000
1!
1*
b101 6
19
1>
1C
b101 G
#301240000000
0!
0*
09
0>
0C
#301250000000
1!
1*
b110 6
19
1>
1C
b110 G
#301260000000
0!
0*
09
0>
0C
#301270000000
1!
1*
b111 6
19
1>
1C
b111 G
#301280000000
0!
1"
0*
1+
09
1:
0>
0C
#301290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#301300000000
0!
0*
09
0>
0C
#301310000000
1!
1*
b1 6
19
1>
1C
b1 G
#301320000000
0!
0*
09
0>
0C
#301330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#301340000000
0!
0*
09
0>
0C
#301350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#301360000000
0!
0*
09
0>
0C
#301370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#301380000000
0!
0*
09
0>
0C
#301390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#301400000000
0!
0#
0*
0,
09
0>
0?
0C
#301410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#301420000000
0!
0*
09
0>
0C
#301430000000
1!
1*
19
1>
1C
#301440000000
0!
0*
09
0>
0C
#301450000000
1!
1*
19
1>
1C
#301460000000
0!
0*
09
0>
0C
#301470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#301480000000
0!
0*
09
0>
0C
#301490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#301500000000
0!
0*
09
0>
0C
#301510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#301520000000
0!
0*
09
0>
0C
#301530000000
1!
1*
b10 6
19
1>
1C
b10 G
#301540000000
0!
0*
09
0>
0C
#301550000000
1!
1*
b11 6
19
1>
1C
b11 G
#301560000000
0!
0*
09
0>
0C
#301570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#301580000000
0!
0*
09
0>
0C
#301590000000
1!
1*
b101 6
19
1>
1C
b101 G
#301600000000
0!
0*
09
0>
0C
#301610000000
1!
1*
b110 6
19
1>
1C
b110 G
#301620000000
0!
0*
09
0>
0C
#301630000000
1!
1*
b111 6
19
1>
1C
b111 G
#301640000000
0!
0*
09
0>
0C
#301650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#301660000000
0!
0*
09
0>
0C
#301670000000
1!
1*
b1 6
19
1>
1C
b1 G
#301680000000
0!
0*
09
0>
0C
#301690000000
1!
1*
b10 6
19
1>
1C
b10 G
#301700000000
0!
0*
09
0>
0C
#301710000000
1!
1*
b11 6
19
1>
1C
b11 G
#301720000000
0!
0*
09
0>
0C
#301730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#301740000000
0!
0*
09
0>
0C
#301750000000
1!
1*
b101 6
19
1>
1C
b101 G
#301760000000
0!
0*
09
0>
0C
#301770000000
1!
1*
b110 6
19
1>
1C
b110 G
#301780000000
0!
0*
09
0>
0C
#301790000000
1!
1*
b111 6
19
1>
1C
b111 G
#301800000000
0!
0*
09
0>
0C
#301810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#301820000000
0!
0*
09
0>
0C
#301830000000
1!
1*
b1 6
19
1>
1C
b1 G
#301840000000
0!
0*
09
0>
0C
#301850000000
1!
1*
b10 6
19
1>
1C
b10 G
#301860000000
0!
0*
09
0>
0C
#301870000000
1!
1*
b11 6
19
1>
1C
b11 G
#301880000000
0!
0*
09
0>
0C
#301890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#301900000000
0!
0*
09
0>
0C
#301910000000
1!
1*
b101 6
19
1>
1C
b101 G
#301920000000
0!
0*
09
0>
0C
#301930000000
1!
1*
b110 6
19
1>
1C
b110 G
#301940000000
0!
0*
09
0>
0C
#301950000000
1!
1*
b111 6
19
1>
1C
b111 G
#301960000000
0!
1"
0*
1+
09
1:
0>
0C
#301970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#301980000000
0!
0*
09
0>
0C
#301990000000
1!
1*
b1 6
19
1>
1C
b1 G
#302000000000
0!
0*
09
0>
0C
#302010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#302020000000
0!
0*
09
0>
0C
#302030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#302040000000
0!
0*
09
0>
0C
#302050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#302060000000
0!
0*
09
0>
0C
#302070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#302080000000
0!
0#
0*
0,
09
0>
0?
0C
#302090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#302100000000
0!
0*
09
0>
0C
#302110000000
1!
1*
19
1>
1C
#302120000000
0!
0*
09
0>
0C
#302130000000
1!
1*
19
1>
1C
#302140000000
0!
0*
09
0>
0C
#302150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#302160000000
0!
0*
09
0>
0C
#302170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#302180000000
0!
0*
09
0>
0C
#302190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#302200000000
0!
0*
09
0>
0C
#302210000000
1!
1*
b10 6
19
1>
1C
b10 G
#302220000000
0!
0*
09
0>
0C
#302230000000
1!
1*
b11 6
19
1>
1C
b11 G
#302240000000
0!
0*
09
0>
0C
#302250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#302260000000
0!
0*
09
0>
0C
#302270000000
1!
1*
b101 6
19
1>
1C
b101 G
#302280000000
0!
0*
09
0>
0C
#302290000000
1!
1*
b110 6
19
1>
1C
b110 G
#302300000000
0!
0*
09
0>
0C
#302310000000
1!
1*
b111 6
19
1>
1C
b111 G
#302320000000
0!
0*
09
0>
0C
#302330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#302340000000
0!
0*
09
0>
0C
#302350000000
1!
1*
b1 6
19
1>
1C
b1 G
#302360000000
0!
0*
09
0>
0C
#302370000000
1!
1*
b10 6
19
1>
1C
b10 G
#302380000000
0!
0*
09
0>
0C
#302390000000
1!
1*
b11 6
19
1>
1C
b11 G
#302400000000
0!
0*
09
0>
0C
#302410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#302420000000
0!
0*
09
0>
0C
#302430000000
1!
1*
b101 6
19
1>
1C
b101 G
#302440000000
0!
0*
09
0>
0C
#302450000000
1!
1*
b110 6
19
1>
1C
b110 G
#302460000000
0!
0*
09
0>
0C
#302470000000
1!
1*
b111 6
19
1>
1C
b111 G
#302480000000
0!
0*
09
0>
0C
#302490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#302500000000
0!
0*
09
0>
0C
#302510000000
1!
1*
b1 6
19
1>
1C
b1 G
#302520000000
0!
0*
09
0>
0C
#302530000000
1!
1*
b10 6
19
1>
1C
b10 G
#302540000000
0!
0*
09
0>
0C
#302550000000
1!
1*
b11 6
19
1>
1C
b11 G
#302560000000
0!
0*
09
0>
0C
#302570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#302580000000
0!
0*
09
0>
0C
#302590000000
1!
1*
b101 6
19
1>
1C
b101 G
#302600000000
0!
0*
09
0>
0C
#302610000000
1!
1*
b110 6
19
1>
1C
b110 G
#302620000000
0!
0*
09
0>
0C
#302630000000
1!
1*
b111 6
19
1>
1C
b111 G
#302640000000
0!
1"
0*
1+
09
1:
0>
0C
#302650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#302660000000
0!
0*
09
0>
0C
#302670000000
1!
1*
b1 6
19
1>
1C
b1 G
#302680000000
0!
0*
09
0>
0C
#302690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#302700000000
0!
0*
09
0>
0C
#302710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#302720000000
0!
0*
09
0>
0C
#302730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#302740000000
0!
0*
09
0>
0C
#302750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#302760000000
0!
0#
0*
0,
09
0>
0?
0C
#302770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#302780000000
0!
0*
09
0>
0C
#302790000000
1!
1*
19
1>
1C
#302800000000
0!
0*
09
0>
0C
#302810000000
1!
1*
19
1>
1C
#302820000000
0!
0*
09
0>
0C
#302830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#302840000000
0!
0*
09
0>
0C
#302850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#302860000000
0!
0*
09
0>
0C
#302870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#302880000000
0!
0*
09
0>
0C
#302890000000
1!
1*
b10 6
19
1>
1C
b10 G
#302900000000
0!
0*
09
0>
0C
#302910000000
1!
1*
b11 6
19
1>
1C
b11 G
#302920000000
0!
0*
09
0>
0C
#302930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#302940000000
0!
0*
09
0>
0C
#302950000000
1!
1*
b101 6
19
1>
1C
b101 G
#302960000000
0!
0*
09
0>
0C
#302970000000
1!
1*
b110 6
19
1>
1C
b110 G
#302980000000
0!
0*
09
0>
0C
#302990000000
1!
1*
b111 6
19
1>
1C
b111 G
#303000000000
0!
0*
09
0>
0C
#303010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#303020000000
0!
0*
09
0>
0C
#303030000000
1!
1*
b1 6
19
1>
1C
b1 G
#303040000000
0!
0*
09
0>
0C
#303050000000
1!
1*
b10 6
19
1>
1C
b10 G
#303060000000
0!
0*
09
0>
0C
#303070000000
1!
1*
b11 6
19
1>
1C
b11 G
#303080000000
0!
0*
09
0>
0C
#303090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#303100000000
0!
0*
09
0>
0C
#303110000000
1!
1*
b101 6
19
1>
1C
b101 G
#303120000000
0!
0*
09
0>
0C
#303130000000
1!
1*
b110 6
19
1>
1C
b110 G
#303140000000
0!
0*
09
0>
0C
#303150000000
1!
1*
b111 6
19
1>
1C
b111 G
#303160000000
0!
0*
09
0>
0C
#303170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#303180000000
0!
0*
09
0>
0C
#303190000000
1!
1*
b1 6
19
1>
1C
b1 G
#303200000000
0!
0*
09
0>
0C
#303210000000
1!
1*
b10 6
19
1>
1C
b10 G
#303220000000
0!
0*
09
0>
0C
#303230000000
1!
1*
b11 6
19
1>
1C
b11 G
#303240000000
0!
0*
09
0>
0C
#303250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#303260000000
0!
0*
09
0>
0C
#303270000000
1!
1*
b101 6
19
1>
1C
b101 G
#303280000000
0!
0*
09
0>
0C
#303290000000
1!
1*
b110 6
19
1>
1C
b110 G
#303300000000
0!
0*
09
0>
0C
#303310000000
1!
1*
b111 6
19
1>
1C
b111 G
#303320000000
0!
1"
0*
1+
09
1:
0>
0C
#303330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#303340000000
0!
0*
09
0>
0C
#303350000000
1!
1*
b1 6
19
1>
1C
b1 G
#303360000000
0!
0*
09
0>
0C
#303370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#303380000000
0!
0*
09
0>
0C
#303390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#303400000000
0!
0*
09
0>
0C
#303410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#303420000000
0!
0*
09
0>
0C
#303430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#303440000000
0!
0#
0*
0,
09
0>
0?
0C
#303450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#303460000000
0!
0*
09
0>
0C
#303470000000
1!
1*
19
1>
1C
#303480000000
0!
0*
09
0>
0C
#303490000000
1!
1*
19
1>
1C
#303500000000
0!
0*
09
0>
0C
#303510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#303520000000
0!
0*
09
0>
0C
#303530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#303540000000
0!
0*
09
0>
0C
#303550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#303560000000
0!
0*
09
0>
0C
#303570000000
1!
1*
b10 6
19
1>
1C
b10 G
#303580000000
0!
0*
09
0>
0C
#303590000000
1!
1*
b11 6
19
1>
1C
b11 G
#303600000000
0!
0*
09
0>
0C
#303610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#303620000000
0!
0*
09
0>
0C
#303630000000
1!
1*
b101 6
19
1>
1C
b101 G
#303640000000
0!
0*
09
0>
0C
#303650000000
1!
1*
b110 6
19
1>
1C
b110 G
#303660000000
0!
0*
09
0>
0C
#303670000000
1!
1*
b111 6
19
1>
1C
b111 G
#303680000000
0!
0*
09
0>
0C
#303690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#303700000000
0!
0*
09
0>
0C
#303710000000
1!
1*
b1 6
19
1>
1C
b1 G
#303720000000
0!
0*
09
0>
0C
#303730000000
1!
1*
b10 6
19
1>
1C
b10 G
#303740000000
0!
0*
09
0>
0C
#303750000000
1!
1*
b11 6
19
1>
1C
b11 G
#303760000000
0!
0*
09
0>
0C
#303770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#303780000000
0!
0*
09
0>
0C
#303790000000
1!
1*
b101 6
19
1>
1C
b101 G
#303800000000
0!
0*
09
0>
0C
#303810000000
1!
1*
b110 6
19
1>
1C
b110 G
#303820000000
0!
0*
09
0>
0C
#303830000000
1!
1*
b111 6
19
1>
1C
b111 G
#303840000000
0!
0*
09
0>
0C
#303850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#303860000000
0!
0*
09
0>
0C
#303870000000
1!
1*
b1 6
19
1>
1C
b1 G
#303880000000
0!
0*
09
0>
0C
#303890000000
1!
1*
b10 6
19
1>
1C
b10 G
#303900000000
0!
0*
09
0>
0C
#303910000000
1!
1*
b11 6
19
1>
1C
b11 G
#303920000000
0!
0*
09
0>
0C
#303930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#303940000000
0!
0*
09
0>
0C
#303950000000
1!
1*
b101 6
19
1>
1C
b101 G
#303960000000
0!
0*
09
0>
0C
#303970000000
1!
1*
b110 6
19
1>
1C
b110 G
#303980000000
0!
0*
09
0>
0C
#303990000000
1!
1*
b111 6
19
1>
1C
b111 G
#304000000000
0!
1"
0*
1+
09
1:
0>
0C
#304010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#304020000000
0!
0*
09
0>
0C
#304030000000
1!
1*
b1 6
19
1>
1C
b1 G
#304040000000
0!
0*
09
0>
0C
#304050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#304060000000
0!
0*
09
0>
0C
#304070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#304080000000
0!
0*
09
0>
0C
#304090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#304100000000
0!
0*
09
0>
0C
#304110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#304120000000
0!
0#
0*
0,
09
0>
0?
0C
#304130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#304140000000
0!
0*
09
0>
0C
#304150000000
1!
1*
19
1>
1C
#304160000000
0!
0*
09
0>
0C
#304170000000
1!
1*
19
1>
1C
#304180000000
0!
0*
09
0>
0C
#304190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#304200000000
0!
0*
09
0>
0C
#304210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#304220000000
0!
0*
09
0>
0C
#304230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#304240000000
0!
0*
09
0>
0C
#304250000000
1!
1*
b10 6
19
1>
1C
b10 G
#304260000000
0!
0*
09
0>
0C
#304270000000
1!
1*
b11 6
19
1>
1C
b11 G
#304280000000
0!
0*
09
0>
0C
#304290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#304300000000
0!
0*
09
0>
0C
#304310000000
1!
1*
b101 6
19
1>
1C
b101 G
#304320000000
0!
0*
09
0>
0C
#304330000000
1!
1*
b110 6
19
1>
1C
b110 G
#304340000000
0!
0*
09
0>
0C
#304350000000
1!
1*
b111 6
19
1>
1C
b111 G
#304360000000
0!
0*
09
0>
0C
#304370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#304380000000
0!
0*
09
0>
0C
#304390000000
1!
1*
b1 6
19
1>
1C
b1 G
#304400000000
0!
0*
09
0>
0C
#304410000000
1!
1*
b10 6
19
1>
1C
b10 G
#304420000000
0!
0*
09
0>
0C
#304430000000
1!
1*
b11 6
19
1>
1C
b11 G
#304440000000
0!
0*
09
0>
0C
#304450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#304460000000
0!
0*
09
0>
0C
#304470000000
1!
1*
b101 6
19
1>
1C
b101 G
#304480000000
0!
0*
09
0>
0C
#304490000000
1!
1*
b110 6
19
1>
1C
b110 G
#304500000000
0!
0*
09
0>
0C
#304510000000
1!
1*
b111 6
19
1>
1C
b111 G
#304520000000
0!
0*
09
0>
0C
#304530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#304540000000
0!
0*
09
0>
0C
#304550000000
1!
1*
b1 6
19
1>
1C
b1 G
#304560000000
0!
0*
09
0>
0C
#304570000000
1!
1*
b10 6
19
1>
1C
b10 G
#304580000000
0!
0*
09
0>
0C
#304590000000
1!
1*
b11 6
19
1>
1C
b11 G
#304600000000
0!
0*
09
0>
0C
#304610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#304620000000
0!
0*
09
0>
0C
#304630000000
1!
1*
b101 6
19
1>
1C
b101 G
#304640000000
0!
0*
09
0>
0C
#304650000000
1!
1*
b110 6
19
1>
1C
b110 G
#304660000000
0!
0*
09
0>
0C
#304670000000
1!
1*
b111 6
19
1>
1C
b111 G
#304680000000
0!
1"
0*
1+
09
1:
0>
0C
#304690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#304700000000
0!
0*
09
0>
0C
#304710000000
1!
1*
b1 6
19
1>
1C
b1 G
#304720000000
0!
0*
09
0>
0C
#304730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#304740000000
0!
0*
09
0>
0C
#304750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#304760000000
0!
0*
09
0>
0C
#304770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#304780000000
0!
0*
09
0>
0C
#304790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#304800000000
0!
0#
0*
0,
09
0>
0?
0C
#304810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#304820000000
0!
0*
09
0>
0C
#304830000000
1!
1*
19
1>
1C
#304840000000
0!
0*
09
0>
0C
#304850000000
1!
1*
19
1>
1C
#304860000000
0!
0*
09
0>
0C
#304870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#304880000000
0!
0*
09
0>
0C
#304890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#304900000000
0!
0*
09
0>
0C
#304910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#304920000000
0!
0*
09
0>
0C
#304930000000
1!
1*
b10 6
19
1>
1C
b10 G
#304940000000
0!
0*
09
0>
0C
#304950000000
1!
1*
b11 6
19
1>
1C
b11 G
#304960000000
0!
0*
09
0>
0C
#304970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#304980000000
0!
0*
09
0>
0C
#304990000000
1!
1*
b101 6
19
1>
1C
b101 G
#305000000000
0!
0*
09
0>
0C
#305010000000
1!
1*
b110 6
19
1>
1C
b110 G
#305020000000
0!
0*
09
0>
0C
#305030000000
1!
1*
b111 6
19
1>
1C
b111 G
#305040000000
0!
0*
09
0>
0C
#305050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#305060000000
0!
0*
09
0>
0C
#305070000000
1!
1*
b1 6
19
1>
1C
b1 G
#305080000000
0!
0*
09
0>
0C
#305090000000
1!
1*
b10 6
19
1>
1C
b10 G
#305100000000
0!
0*
09
0>
0C
#305110000000
1!
1*
b11 6
19
1>
1C
b11 G
#305120000000
0!
0*
09
0>
0C
#305130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#305140000000
0!
0*
09
0>
0C
#305150000000
1!
1*
b101 6
19
1>
1C
b101 G
#305160000000
0!
0*
09
0>
0C
#305170000000
1!
1*
b110 6
19
1>
1C
b110 G
#305180000000
0!
0*
09
0>
0C
#305190000000
1!
1*
b111 6
19
1>
1C
b111 G
#305200000000
0!
0*
09
0>
0C
#305210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#305220000000
0!
0*
09
0>
0C
#305230000000
1!
1*
b1 6
19
1>
1C
b1 G
#305240000000
0!
0*
09
0>
0C
#305250000000
1!
1*
b10 6
19
1>
1C
b10 G
#305260000000
0!
0*
09
0>
0C
#305270000000
1!
1*
b11 6
19
1>
1C
b11 G
#305280000000
0!
0*
09
0>
0C
#305290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#305300000000
0!
0*
09
0>
0C
#305310000000
1!
1*
b101 6
19
1>
1C
b101 G
#305320000000
0!
0*
09
0>
0C
#305330000000
1!
1*
b110 6
19
1>
1C
b110 G
#305340000000
0!
0*
09
0>
0C
#305350000000
1!
1*
b111 6
19
1>
1C
b111 G
#305360000000
0!
1"
0*
1+
09
1:
0>
0C
#305370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#305380000000
0!
0*
09
0>
0C
#305390000000
1!
1*
b1 6
19
1>
1C
b1 G
#305400000000
0!
0*
09
0>
0C
#305410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#305420000000
0!
0*
09
0>
0C
#305430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#305440000000
0!
0*
09
0>
0C
#305450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#305460000000
0!
0*
09
0>
0C
#305470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#305480000000
0!
0#
0*
0,
09
0>
0?
0C
#305490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#305500000000
0!
0*
09
0>
0C
#305510000000
1!
1*
19
1>
1C
#305520000000
0!
0*
09
0>
0C
#305530000000
1!
1*
19
1>
1C
#305540000000
0!
0*
09
0>
0C
#305550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#305560000000
0!
0*
09
0>
0C
#305570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#305580000000
0!
0*
09
0>
0C
#305590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#305600000000
0!
0*
09
0>
0C
#305610000000
1!
1*
b10 6
19
1>
1C
b10 G
#305620000000
0!
0*
09
0>
0C
#305630000000
1!
1*
b11 6
19
1>
1C
b11 G
#305640000000
0!
0*
09
0>
0C
#305650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#305660000000
0!
0*
09
0>
0C
#305670000000
1!
1*
b101 6
19
1>
1C
b101 G
#305680000000
0!
0*
09
0>
0C
#305690000000
1!
1*
b110 6
19
1>
1C
b110 G
#305700000000
0!
0*
09
0>
0C
#305710000000
1!
1*
b111 6
19
1>
1C
b111 G
#305720000000
0!
0*
09
0>
0C
#305730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#305740000000
0!
0*
09
0>
0C
#305750000000
1!
1*
b1 6
19
1>
1C
b1 G
#305760000000
0!
0*
09
0>
0C
#305770000000
1!
1*
b10 6
19
1>
1C
b10 G
#305780000000
0!
0*
09
0>
0C
#305790000000
1!
1*
b11 6
19
1>
1C
b11 G
#305800000000
0!
0*
09
0>
0C
#305810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#305820000000
0!
0*
09
0>
0C
#305830000000
1!
1*
b101 6
19
1>
1C
b101 G
#305840000000
0!
0*
09
0>
0C
#305850000000
1!
1*
b110 6
19
1>
1C
b110 G
#305860000000
0!
0*
09
0>
0C
#305870000000
1!
1*
b111 6
19
1>
1C
b111 G
#305880000000
0!
0*
09
0>
0C
#305890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#305900000000
0!
0*
09
0>
0C
#305910000000
1!
1*
b1 6
19
1>
1C
b1 G
#305920000000
0!
0*
09
0>
0C
#305930000000
1!
1*
b10 6
19
1>
1C
b10 G
#305940000000
0!
0*
09
0>
0C
#305950000000
1!
1*
b11 6
19
1>
1C
b11 G
#305960000000
0!
0*
09
0>
0C
#305970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#305980000000
0!
0*
09
0>
0C
#305990000000
1!
1*
b101 6
19
1>
1C
b101 G
#306000000000
0!
0*
09
0>
0C
#306010000000
1!
1*
b110 6
19
1>
1C
b110 G
#306020000000
0!
0*
09
0>
0C
#306030000000
1!
1*
b111 6
19
1>
1C
b111 G
#306040000000
0!
1"
0*
1+
09
1:
0>
0C
#306050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#306060000000
0!
0*
09
0>
0C
#306070000000
1!
1*
b1 6
19
1>
1C
b1 G
#306080000000
0!
0*
09
0>
0C
#306090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#306100000000
0!
0*
09
0>
0C
#306110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#306120000000
0!
0*
09
0>
0C
#306130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#306140000000
0!
0*
09
0>
0C
#306150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#306160000000
0!
0#
0*
0,
09
0>
0?
0C
#306170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#306180000000
0!
0*
09
0>
0C
#306190000000
1!
1*
19
1>
1C
#306200000000
0!
0*
09
0>
0C
#306210000000
1!
1*
19
1>
1C
#306220000000
0!
0*
09
0>
0C
#306230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#306240000000
0!
0*
09
0>
0C
#306250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#306260000000
0!
0*
09
0>
0C
#306270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#306280000000
0!
0*
09
0>
0C
#306290000000
1!
1*
b10 6
19
1>
1C
b10 G
#306300000000
0!
0*
09
0>
0C
#306310000000
1!
1*
b11 6
19
1>
1C
b11 G
#306320000000
0!
0*
09
0>
0C
#306330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#306340000000
0!
0*
09
0>
0C
#306350000000
1!
1*
b101 6
19
1>
1C
b101 G
#306360000000
0!
0*
09
0>
0C
#306370000000
1!
1*
b110 6
19
1>
1C
b110 G
#306380000000
0!
0*
09
0>
0C
#306390000000
1!
1*
b111 6
19
1>
1C
b111 G
#306400000000
0!
0*
09
0>
0C
#306410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#306420000000
0!
0*
09
0>
0C
#306430000000
1!
1*
b1 6
19
1>
1C
b1 G
#306440000000
0!
0*
09
0>
0C
#306450000000
1!
1*
b10 6
19
1>
1C
b10 G
#306460000000
0!
0*
09
0>
0C
#306470000000
1!
1*
b11 6
19
1>
1C
b11 G
#306480000000
0!
0*
09
0>
0C
#306490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#306500000000
0!
0*
09
0>
0C
#306510000000
1!
1*
b101 6
19
1>
1C
b101 G
#306520000000
0!
0*
09
0>
0C
#306530000000
1!
1*
b110 6
19
1>
1C
b110 G
#306540000000
0!
0*
09
0>
0C
#306550000000
1!
1*
b111 6
19
1>
1C
b111 G
#306560000000
0!
0*
09
0>
0C
#306570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#306580000000
0!
0*
09
0>
0C
#306590000000
1!
1*
b1 6
19
1>
1C
b1 G
#306600000000
0!
0*
09
0>
0C
#306610000000
1!
1*
b10 6
19
1>
1C
b10 G
#306620000000
0!
0*
09
0>
0C
#306630000000
1!
1*
b11 6
19
1>
1C
b11 G
#306640000000
0!
0*
09
0>
0C
#306650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#306660000000
0!
0*
09
0>
0C
#306670000000
1!
1*
b101 6
19
1>
1C
b101 G
#306680000000
0!
0*
09
0>
0C
#306690000000
1!
1*
b110 6
19
1>
1C
b110 G
#306700000000
0!
0*
09
0>
0C
#306710000000
1!
1*
b111 6
19
1>
1C
b111 G
#306720000000
0!
1"
0*
1+
09
1:
0>
0C
#306730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#306740000000
0!
0*
09
0>
0C
#306750000000
1!
1*
b1 6
19
1>
1C
b1 G
#306760000000
0!
0*
09
0>
0C
#306770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#306780000000
0!
0*
09
0>
0C
#306790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#306800000000
0!
0*
09
0>
0C
#306810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#306820000000
0!
0*
09
0>
0C
#306830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#306840000000
0!
0#
0*
0,
09
0>
0?
0C
#306850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#306860000000
0!
0*
09
0>
0C
#306870000000
1!
1*
19
1>
1C
#306880000000
0!
0*
09
0>
0C
#306890000000
1!
1*
19
1>
1C
#306900000000
0!
0*
09
0>
0C
#306910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#306920000000
0!
0*
09
0>
0C
#306930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#306940000000
0!
0*
09
0>
0C
#306950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#306960000000
0!
0*
09
0>
0C
#306970000000
1!
1*
b10 6
19
1>
1C
b10 G
#306980000000
0!
0*
09
0>
0C
#306990000000
1!
1*
b11 6
19
1>
1C
b11 G
#307000000000
0!
0*
09
0>
0C
#307010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#307020000000
0!
0*
09
0>
0C
#307030000000
1!
1*
b101 6
19
1>
1C
b101 G
#307040000000
0!
0*
09
0>
0C
#307050000000
1!
1*
b110 6
19
1>
1C
b110 G
#307060000000
0!
0*
09
0>
0C
#307070000000
1!
1*
b111 6
19
1>
1C
b111 G
#307080000000
0!
0*
09
0>
0C
#307090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#307100000000
0!
0*
09
0>
0C
#307110000000
1!
1*
b1 6
19
1>
1C
b1 G
#307120000000
0!
0*
09
0>
0C
#307130000000
1!
1*
b10 6
19
1>
1C
b10 G
#307140000000
0!
0*
09
0>
0C
#307150000000
1!
1*
b11 6
19
1>
1C
b11 G
#307160000000
0!
0*
09
0>
0C
#307170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#307180000000
0!
0*
09
0>
0C
#307190000000
1!
1*
b101 6
19
1>
1C
b101 G
#307200000000
0!
0*
09
0>
0C
#307210000000
1!
1*
b110 6
19
1>
1C
b110 G
#307220000000
0!
0*
09
0>
0C
#307230000000
1!
1*
b111 6
19
1>
1C
b111 G
#307240000000
0!
0*
09
0>
0C
#307250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#307260000000
0!
0*
09
0>
0C
#307270000000
1!
1*
b1 6
19
1>
1C
b1 G
#307280000000
0!
0*
09
0>
0C
#307290000000
1!
1*
b10 6
19
1>
1C
b10 G
#307300000000
0!
0*
09
0>
0C
#307310000000
1!
1*
b11 6
19
1>
1C
b11 G
#307320000000
0!
0*
09
0>
0C
#307330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#307340000000
0!
0*
09
0>
0C
#307350000000
1!
1*
b101 6
19
1>
1C
b101 G
#307360000000
0!
0*
09
0>
0C
#307370000000
1!
1*
b110 6
19
1>
1C
b110 G
#307380000000
0!
0*
09
0>
0C
#307390000000
1!
1*
b111 6
19
1>
1C
b111 G
#307400000000
0!
1"
0*
1+
09
1:
0>
0C
#307410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#307420000000
0!
0*
09
0>
0C
#307430000000
1!
1*
b1 6
19
1>
1C
b1 G
#307440000000
0!
0*
09
0>
0C
#307450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#307460000000
0!
0*
09
0>
0C
#307470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#307480000000
0!
0*
09
0>
0C
#307490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#307500000000
0!
0*
09
0>
0C
#307510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#307520000000
0!
0#
0*
0,
09
0>
0?
0C
#307530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#307540000000
0!
0*
09
0>
0C
#307550000000
1!
1*
19
1>
1C
#307560000000
0!
0*
09
0>
0C
#307570000000
1!
1*
19
1>
1C
#307580000000
0!
0*
09
0>
0C
#307590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#307600000000
0!
0*
09
0>
0C
#307610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#307620000000
0!
0*
09
0>
0C
#307630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#307640000000
0!
0*
09
0>
0C
#307650000000
1!
1*
b10 6
19
1>
1C
b10 G
#307660000000
0!
0*
09
0>
0C
#307670000000
1!
1*
b11 6
19
1>
1C
b11 G
#307680000000
0!
0*
09
0>
0C
#307690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#307700000000
0!
0*
09
0>
0C
#307710000000
1!
1*
b101 6
19
1>
1C
b101 G
#307720000000
0!
0*
09
0>
0C
#307730000000
1!
1*
b110 6
19
1>
1C
b110 G
#307740000000
0!
0*
09
0>
0C
#307750000000
1!
1*
b111 6
19
1>
1C
b111 G
#307760000000
0!
0*
09
0>
0C
#307770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#307780000000
0!
0*
09
0>
0C
#307790000000
1!
1*
b1 6
19
1>
1C
b1 G
#307800000000
0!
0*
09
0>
0C
#307810000000
1!
1*
b10 6
19
1>
1C
b10 G
#307820000000
0!
0*
09
0>
0C
#307830000000
1!
1*
b11 6
19
1>
1C
b11 G
#307840000000
0!
0*
09
0>
0C
#307850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#307860000000
0!
0*
09
0>
0C
#307870000000
1!
1*
b101 6
19
1>
1C
b101 G
#307880000000
0!
0*
09
0>
0C
#307890000000
1!
1*
b110 6
19
1>
1C
b110 G
#307900000000
0!
0*
09
0>
0C
#307910000000
1!
1*
b111 6
19
1>
1C
b111 G
#307920000000
0!
0*
09
0>
0C
#307930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#307940000000
0!
0*
09
0>
0C
#307950000000
1!
1*
b1 6
19
1>
1C
b1 G
#307960000000
0!
0*
09
0>
0C
#307970000000
1!
1*
b10 6
19
1>
1C
b10 G
#307980000000
0!
0*
09
0>
0C
#307990000000
1!
1*
b11 6
19
1>
1C
b11 G
#308000000000
0!
0*
09
0>
0C
#308010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#308020000000
0!
0*
09
0>
0C
#308030000000
1!
1*
b101 6
19
1>
1C
b101 G
#308040000000
0!
0*
09
0>
0C
#308050000000
1!
1*
b110 6
19
1>
1C
b110 G
#308060000000
0!
0*
09
0>
0C
#308070000000
1!
1*
b111 6
19
1>
1C
b111 G
#308080000000
0!
1"
0*
1+
09
1:
0>
0C
#308090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#308100000000
0!
0*
09
0>
0C
#308110000000
1!
1*
b1 6
19
1>
1C
b1 G
#308120000000
0!
0*
09
0>
0C
#308130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#308140000000
0!
0*
09
0>
0C
#308150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#308160000000
0!
0*
09
0>
0C
#308170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#308180000000
0!
0*
09
0>
0C
#308190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#308200000000
0!
0#
0*
0,
09
0>
0?
0C
#308210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#308220000000
0!
0*
09
0>
0C
#308230000000
1!
1*
19
1>
1C
#308240000000
0!
0*
09
0>
0C
#308250000000
1!
1*
19
1>
1C
#308260000000
0!
0*
09
0>
0C
#308270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#308280000000
0!
0*
09
0>
0C
#308290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#308300000000
0!
0*
09
0>
0C
#308310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#308320000000
0!
0*
09
0>
0C
#308330000000
1!
1*
b10 6
19
1>
1C
b10 G
#308340000000
0!
0*
09
0>
0C
#308350000000
1!
1*
b11 6
19
1>
1C
b11 G
#308360000000
0!
0*
09
0>
0C
#308370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#308380000000
0!
0*
09
0>
0C
#308390000000
1!
1*
b101 6
19
1>
1C
b101 G
#308400000000
0!
0*
09
0>
0C
#308410000000
1!
1*
b110 6
19
1>
1C
b110 G
#308420000000
0!
0*
09
0>
0C
#308430000000
1!
1*
b111 6
19
1>
1C
b111 G
#308440000000
0!
0*
09
0>
0C
#308450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#308460000000
0!
0*
09
0>
0C
#308470000000
1!
1*
b1 6
19
1>
1C
b1 G
#308480000000
0!
0*
09
0>
0C
#308490000000
1!
1*
b10 6
19
1>
1C
b10 G
#308500000000
0!
0*
09
0>
0C
#308510000000
1!
1*
b11 6
19
1>
1C
b11 G
#308520000000
0!
0*
09
0>
0C
#308530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#308540000000
0!
0*
09
0>
0C
#308550000000
1!
1*
b101 6
19
1>
1C
b101 G
#308560000000
0!
0*
09
0>
0C
#308570000000
1!
1*
b110 6
19
1>
1C
b110 G
#308580000000
0!
0*
09
0>
0C
#308590000000
1!
1*
b111 6
19
1>
1C
b111 G
#308600000000
0!
0*
09
0>
0C
#308610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#308620000000
0!
0*
09
0>
0C
#308630000000
1!
1*
b1 6
19
1>
1C
b1 G
#308640000000
0!
0*
09
0>
0C
#308650000000
1!
1*
b10 6
19
1>
1C
b10 G
#308660000000
0!
0*
09
0>
0C
#308670000000
1!
1*
b11 6
19
1>
1C
b11 G
#308680000000
0!
0*
09
0>
0C
#308690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#308700000000
0!
0*
09
0>
0C
#308710000000
1!
1*
b101 6
19
1>
1C
b101 G
#308720000000
0!
0*
09
0>
0C
#308730000000
1!
1*
b110 6
19
1>
1C
b110 G
#308740000000
0!
0*
09
0>
0C
#308750000000
1!
1*
b111 6
19
1>
1C
b111 G
#308760000000
0!
1"
0*
1+
09
1:
0>
0C
#308770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#308780000000
0!
0*
09
0>
0C
#308790000000
1!
1*
b1 6
19
1>
1C
b1 G
#308800000000
0!
0*
09
0>
0C
#308810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#308820000000
0!
0*
09
0>
0C
#308830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#308840000000
0!
0*
09
0>
0C
#308850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#308860000000
0!
0*
09
0>
0C
#308870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#308880000000
0!
0#
0*
0,
09
0>
0?
0C
#308890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#308900000000
0!
0*
09
0>
0C
#308910000000
1!
1*
19
1>
1C
#308920000000
0!
0*
09
0>
0C
#308930000000
1!
1*
19
1>
1C
#308940000000
0!
0*
09
0>
0C
#308950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#308960000000
0!
0*
09
0>
0C
#308970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#308980000000
0!
0*
09
0>
0C
#308990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#309000000000
0!
0*
09
0>
0C
#309010000000
1!
1*
b10 6
19
1>
1C
b10 G
#309020000000
0!
0*
09
0>
0C
#309030000000
1!
1*
b11 6
19
1>
1C
b11 G
#309040000000
0!
0*
09
0>
0C
#309050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#309060000000
0!
0*
09
0>
0C
#309070000000
1!
1*
b101 6
19
1>
1C
b101 G
#309080000000
0!
0*
09
0>
0C
#309090000000
1!
1*
b110 6
19
1>
1C
b110 G
#309100000000
0!
0*
09
0>
0C
#309110000000
1!
1*
b111 6
19
1>
1C
b111 G
#309120000000
0!
0*
09
0>
0C
#309130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#309140000000
0!
0*
09
0>
0C
#309150000000
1!
1*
b1 6
19
1>
1C
b1 G
#309160000000
0!
0*
09
0>
0C
#309170000000
1!
1*
b10 6
19
1>
1C
b10 G
#309180000000
0!
0*
09
0>
0C
#309190000000
1!
1*
b11 6
19
1>
1C
b11 G
#309200000000
0!
0*
09
0>
0C
#309210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#309220000000
0!
0*
09
0>
0C
#309230000000
1!
1*
b101 6
19
1>
1C
b101 G
#309240000000
0!
0*
09
0>
0C
#309250000000
1!
1*
b110 6
19
1>
1C
b110 G
#309260000000
0!
0*
09
0>
0C
#309270000000
1!
1*
b111 6
19
1>
1C
b111 G
#309280000000
0!
0*
09
0>
0C
#309290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#309300000000
0!
0*
09
0>
0C
#309310000000
1!
1*
b1 6
19
1>
1C
b1 G
#309320000000
0!
0*
09
0>
0C
#309330000000
1!
1*
b10 6
19
1>
1C
b10 G
#309340000000
0!
0*
09
0>
0C
#309350000000
1!
1*
b11 6
19
1>
1C
b11 G
#309360000000
0!
0*
09
0>
0C
#309370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#309380000000
0!
0*
09
0>
0C
#309390000000
1!
1*
b101 6
19
1>
1C
b101 G
#309400000000
0!
0*
09
0>
0C
#309410000000
1!
1*
b110 6
19
1>
1C
b110 G
#309420000000
0!
0*
09
0>
0C
#309430000000
1!
1*
b111 6
19
1>
1C
b111 G
#309440000000
0!
1"
0*
1+
09
1:
0>
0C
#309450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#309460000000
0!
0*
09
0>
0C
#309470000000
1!
1*
b1 6
19
1>
1C
b1 G
#309480000000
0!
0*
09
0>
0C
#309490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#309500000000
0!
0*
09
0>
0C
#309510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#309520000000
0!
0*
09
0>
0C
#309530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#309540000000
0!
0*
09
0>
0C
#309550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#309560000000
0!
0#
0*
0,
09
0>
0?
0C
#309570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#309580000000
0!
0*
09
0>
0C
#309590000000
1!
1*
19
1>
1C
#309600000000
0!
0*
09
0>
0C
#309610000000
1!
1*
19
1>
1C
#309620000000
0!
0*
09
0>
0C
#309630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#309640000000
0!
0*
09
0>
0C
#309650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#309660000000
0!
0*
09
0>
0C
#309670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#309680000000
0!
0*
09
0>
0C
#309690000000
1!
1*
b10 6
19
1>
1C
b10 G
#309700000000
0!
0*
09
0>
0C
#309710000000
1!
1*
b11 6
19
1>
1C
b11 G
#309720000000
0!
0*
09
0>
0C
#309730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#309740000000
0!
0*
09
0>
0C
#309750000000
1!
1*
b101 6
19
1>
1C
b101 G
#309760000000
0!
0*
09
0>
0C
#309770000000
1!
1*
b110 6
19
1>
1C
b110 G
#309780000000
0!
0*
09
0>
0C
#309790000000
1!
1*
b111 6
19
1>
1C
b111 G
#309800000000
0!
0*
09
0>
0C
#309810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#309820000000
0!
0*
09
0>
0C
#309830000000
1!
1*
b1 6
19
1>
1C
b1 G
#309840000000
0!
0*
09
0>
0C
#309850000000
1!
1*
b10 6
19
1>
1C
b10 G
#309860000000
0!
0*
09
0>
0C
#309870000000
1!
1*
b11 6
19
1>
1C
b11 G
#309880000000
0!
0*
09
0>
0C
#309890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#309900000000
0!
0*
09
0>
0C
#309910000000
1!
1*
b101 6
19
1>
1C
b101 G
#309920000000
0!
0*
09
0>
0C
#309930000000
1!
1*
b110 6
19
1>
1C
b110 G
#309940000000
0!
0*
09
0>
0C
#309950000000
1!
1*
b111 6
19
1>
1C
b111 G
#309960000000
0!
0*
09
0>
0C
#309970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#309980000000
0!
0*
09
0>
0C
#309990000000
1!
1*
b1 6
19
1>
1C
b1 G
#310000000000
0!
0*
09
0>
0C
#310010000000
1!
1*
b10 6
19
1>
1C
b10 G
#310020000000
0!
0*
09
0>
0C
#310030000000
1!
1*
b11 6
19
1>
1C
b11 G
#310040000000
0!
0*
09
0>
0C
#310050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#310060000000
0!
0*
09
0>
0C
#310070000000
1!
1*
b101 6
19
1>
1C
b101 G
#310080000000
0!
0*
09
0>
0C
#310090000000
1!
1*
b110 6
19
1>
1C
b110 G
#310100000000
0!
0*
09
0>
0C
#310110000000
1!
1*
b111 6
19
1>
1C
b111 G
#310120000000
0!
1"
0*
1+
09
1:
0>
0C
#310130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#310140000000
0!
0*
09
0>
0C
#310150000000
1!
1*
b1 6
19
1>
1C
b1 G
#310160000000
0!
0*
09
0>
0C
#310170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#310180000000
0!
0*
09
0>
0C
#310190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#310200000000
0!
0*
09
0>
0C
#310210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#310220000000
0!
0*
09
0>
0C
#310230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#310240000000
0!
0#
0*
0,
09
0>
0?
0C
#310250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#310260000000
0!
0*
09
0>
0C
#310270000000
1!
1*
19
1>
1C
#310280000000
0!
0*
09
0>
0C
#310290000000
1!
1*
19
1>
1C
#310300000000
0!
0*
09
0>
0C
#310310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#310320000000
0!
0*
09
0>
0C
#310330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#310340000000
0!
0*
09
0>
0C
#310350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#310360000000
0!
0*
09
0>
0C
#310370000000
1!
1*
b10 6
19
1>
1C
b10 G
#310380000000
0!
0*
09
0>
0C
#310390000000
1!
1*
b11 6
19
1>
1C
b11 G
#310400000000
0!
0*
09
0>
0C
#310410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#310420000000
0!
0*
09
0>
0C
#310430000000
1!
1*
b101 6
19
1>
1C
b101 G
#310440000000
0!
0*
09
0>
0C
#310450000000
1!
1*
b110 6
19
1>
1C
b110 G
#310460000000
0!
0*
09
0>
0C
#310470000000
1!
1*
b111 6
19
1>
1C
b111 G
#310480000000
0!
0*
09
0>
0C
#310490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#310500000000
0!
0*
09
0>
0C
#310510000000
1!
1*
b1 6
19
1>
1C
b1 G
#310520000000
0!
0*
09
0>
0C
#310530000000
1!
1*
b10 6
19
1>
1C
b10 G
#310540000000
0!
0*
09
0>
0C
#310550000000
1!
1*
b11 6
19
1>
1C
b11 G
#310560000000
0!
0*
09
0>
0C
#310570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#310580000000
0!
0*
09
0>
0C
#310590000000
1!
1*
b101 6
19
1>
1C
b101 G
#310600000000
0!
0*
09
0>
0C
#310610000000
1!
1*
b110 6
19
1>
1C
b110 G
#310620000000
0!
0*
09
0>
0C
#310630000000
1!
1*
b111 6
19
1>
1C
b111 G
#310640000000
0!
0*
09
0>
0C
#310650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#310660000000
0!
0*
09
0>
0C
#310670000000
1!
1*
b1 6
19
1>
1C
b1 G
#310680000000
0!
0*
09
0>
0C
#310690000000
1!
1*
b10 6
19
1>
1C
b10 G
#310700000000
0!
0*
09
0>
0C
#310710000000
1!
1*
b11 6
19
1>
1C
b11 G
#310720000000
0!
0*
09
0>
0C
#310730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#310740000000
0!
0*
09
0>
0C
#310750000000
1!
1*
b101 6
19
1>
1C
b101 G
#310760000000
0!
0*
09
0>
0C
#310770000000
1!
1*
b110 6
19
1>
1C
b110 G
#310780000000
0!
0*
09
0>
0C
#310790000000
1!
1*
b111 6
19
1>
1C
b111 G
#310800000000
0!
1"
0*
1+
09
1:
0>
0C
#310810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#310820000000
0!
0*
09
0>
0C
#310830000000
1!
1*
b1 6
19
1>
1C
b1 G
#310840000000
0!
0*
09
0>
0C
#310850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#310860000000
0!
0*
09
0>
0C
#310870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#310880000000
0!
0*
09
0>
0C
#310890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#310900000000
0!
0*
09
0>
0C
#310910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#310920000000
0!
0#
0*
0,
09
0>
0?
0C
#310930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#310940000000
0!
0*
09
0>
0C
#310950000000
1!
1*
19
1>
1C
#310960000000
0!
0*
09
0>
0C
#310970000000
1!
1*
19
1>
1C
#310980000000
0!
0*
09
0>
0C
#310990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#311000000000
0!
0*
09
0>
0C
#311010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#311020000000
0!
0*
09
0>
0C
#311030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#311040000000
0!
0*
09
0>
0C
#311050000000
1!
1*
b10 6
19
1>
1C
b10 G
#311060000000
0!
0*
09
0>
0C
#311070000000
1!
1*
b11 6
19
1>
1C
b11 G
#311080000000
0!
0*
09
0>
0C
#311090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#311100000000
0!
0*
09
0>
0C
#311110000000
1!
1*
b101 6
19
1>
1C
b101 G
#311120000000
0!
0*
09
0>
0C
#311130000000
1!
1*
b110 6
19
1>
1C
b110 G
#311140000000
0!
0*
09
0>
0C
#311150000000
1!
1*
b111 6
19
1>
1C
b111 G
#311160000000
0!
0*
09
0>
0C
#311170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#311180000000
0!
0*
09
0>
0C
#311190000000
1!
1*
b1 6
19
1>
1C
b1 G
#311200000000
0!
0*
09
0>
0C
#311210000000
1!
1*
b10 6
19
1>
1C
b10 G
#311220000000
0!
0*
09
0>
0C
#311230000000
1!
1*
b11 6
19
1>
1C
b11 G
#311240000000
0!
0*
09
0>
0C
#311250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#311260000000
0!
0*
09
0>
0C
#311270000000
1!
1*
b101 6
19
1>
1C
b101 G
#311280000000
0!
0*
09
0>
0C
#311290000000
1!
1*
b110 6
19
1>
1C
b110 G
#311300000000
0!
0*
09
0>
0C
#311310000000
1!
1*
b111 6
19
1>
1C
b111 G
#311320000000
0!
0*
09
0>
0C
#311330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#311340000000
0!
0*
09
0>
0C
#311350000000
1!
1*
b1 6
19
1>
1C
b1 G
#311360000000
0!
0*
09
0>
0C
#311370000000
1!
1*
b10 6
19
1>
1C
b10 G
#311380000000
0!
0*
09
0>
0C
#311390000000
1!
1*
b11 6
19
1>
1C
b11 G
#311400000000
0!
0*
09
0>
0C
#311410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#311420000000
0!
0*
09
0>
0C
#311430000000
1!
1*
b101 6
19
1>
1C
b101 G
#311440000000
0!
0*
09
0>
0C
#311450000000
1!
1*
b110 6
19
1>
1C
b110 G
#311460000000
0!
0*
09
0>
0C
#311470000000
1!
1*
b111 6
19
1>
1C
b111 G
#311480000000
0!
1"
0*
1+
09
1:
0>
0C
#311490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#311500000000
0!
0*
09
0>
0C
#311510000000
1!
1*
b1 6
19
1>
1C
b1 G
#311520000000
0!
0*
09
0>
0C
#311530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#311540000000
0!
0*
09
0>
0C
#311550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#311560000000
0!
0*
09
0>
0C
#311570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#311580000000
0!
0*
09
0>
0C
#311590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#311600000000
0!
0#
0*
0,
09
0>
0?
0C
#311610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#311620000000
0!
0*
09
0>
0C
#311630000000
1!
1*
19
1>
1C
#311640000000
0!
0*
09
0>
0C
#311650000000
1!
1*
19
1>
1C
#311660000000
0!
0*
09
0>
0C
#311670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#311680000000
0!
0*
09
0>
0C
#311690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#311700000000
0!
0*
09
0>
0C
#311710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#311720000000
0!
0*
09
0>
0C
#311730000000
1!
1*
b10 6
19
1>
1C
b10 G
#311740000000
0!
0*
09
0>
0C
#311750000000
1!
1*
b11 6
19
1>
1C
b11 G
#311760000000
0!
0*
09
0>
0C
#311770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#311780000000
0!
0*
09
0>
0C
#311790000000
1!
1*
b101 6
19
1>
1C
b101 G
#311800000000
0!
0*
09
0>
0C
#311810000000
1!
1*
b110 6
19
1>
1C
b110 G
#311820000000
0!
0*
09
0>
0C
#311830000000
1!
1*
b111 6
19
1>
1C
b111 G
#311840000000
0!
0*
09
0>
0C
#311850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#311860000000
0!
0*
09
0>
0C
#311870000000
1!
1*
b1 6
19
1>
1C
b1 G
#311880000000
0!
0*
09
0>
0C
#311890000000
1!
1*
b10 6
19
1>
1C
b10 G
#311900000000
0!
0*
09
0>
0C
#311910000000
1!
1*
b11 6
19
1>
1C
b11 G
#311920000000
0!
0*
09
0>
0C
#311930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#311940000000
0!
0*
09
0>
0C
#311950000000
1!
1*
b101 6
19
1>
1C
b101 G
#311960000000
0!
0*
09
0>
0C
#311970000000
1!
1*
b110 6
19
1>
1C
b110 G
#311980000000
0!
0*
09
0>
0C
#311990000000
1!
1*
b111 6
19
1>
1C
b111 G
#312000000000
0!
0*
09
0>
0C
#312010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#312020000000
0!
0*
09
0>
0C
#312030000000
1!
1*
b1 6
19
1>
1C
b1 G
#312040000000
0!
0*
09
0>
0C
#312050000000
1!
1*
b10 6
19
1>
1C
b10 G
#312060000000
0!
0*
09
0>
0C
#312070000000
1!
1*
b11 6
19
1>
1C
b11 G
#312080000000
0!
0*
09
0>
0C
#312090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#312100000000
0!
0*
09
0>
0C
#312110000000
1!
1*
b101 6
19
1>
1C
b101 G
#312120000000
0!
0*
09
0>
0C
#312130000000
1!
1*
b110 6
19
1>
1C
b110 G
#312140000000
0!
0*
09
0>
0C
#312150000000
1!
1*
b111 6
19
1>
1C
b111 G
#312160000000
0!
1"
0*
1+
09
1:
0>
0C
#312170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#312180000000
0!
0*
09
0>
0C
#312190000000
1!
1*
b1 6
19
1>
1C
b1 G
#312200000000
0!
0*
09
0>
0C
#312210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#312220000000
0!
0*
09
0>
0C
#312230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#312240000000
0!
0*
09
0>
0C
#312250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#312260000000
0!
0*
09
0>
0C
#312270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#312280000000
0!
0#
0*
0,
09
0>
0?
0C
#312290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#312300000000
0!
0*
09
0>
0C
#312310000000
1!
1*
19
1>
1C
#312320000000
0!
0*
09
0>
0C
#312330000000
1!
1*
19
1>
1C
#312340000000
0!
0*
09
0>
0C
#312350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#312360000000
0!
0*
09
0>
0C
#312370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#312380000000
0!
0*
09
0>
0C
#312390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#312400000000
0!
0*
09
0>
0C
#312410000000
1!
1*
b10 6
19
1>
1C
b10 G
#312420000000
0!
0*
09
0>
0C
#312430000000
1!
1*
b11 6
19
1>
1C
b11 G
#312440000000
0!
0*
09
0>
0C
#312450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#312460000000
0!
0*
09
0>
0C
#312470000000
1!
1*
b101 6
19
1>
1C
b101 G
#312480000000
0!
0*
09
0>
0C
#312490000000
1!
1*
b110 6
19
1>
1C
b110 G
#312500000000
0!
0*
09
0>
0C
#312510000000
1!
1*
b111 6
19
1>
1C
b111 G
#312520000000
0!
0*
09
0>
0C
#312530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#312540000000
0!
0*
09
0>
0C
#312550000000
1!
1*
b1 6
19
1>
1C
b1 G
#312560000000
0!
0*
09
0>
0C
#312570000000
1!
1*
b10 6
19
1>
1C
b10 G
#312580000000
0!
0*
09
0>
0C
#312590000000
1!
1*
b11 6
19
1>
1C
b11 G
#312600000000
0!
0*
09
0>
0C
#312610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#312620000000
0!
0*
09
0>
0C
#312630000000
1!
1*
b101 6
19
1>
1C
b101 G
#312640000000
0!
0*
09
0>
0C
#312650000000
1!
1*
b110 6
19
1>
1C
b110 G
#312660000000
0!
0*
09
0>
0C
#312670000000
1!
1*
b111 6
19
1>
1C
b111 G
#312680000000
0!
0*
09
0>
0C
#312690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#312700000000
0!
0*
09
0>
0C
#312710000000
1!
1*
b1 6
19
1>
1C
b1 G
#312720000000
0!
0*
09
0>
0C
#312730000000
1!
1*
b10 6
19
1>
1C
b10 G
#312740000000
0!
0*
09
0>
0C
#312750000000
1!
1*
b11 6
19
1>
1C
b11 G
#312760000000
0!
0*
09
0>
0C
#312770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#312780000000
0!
0*
09
0>
0C
#312790000000
1!
1*
b101 6
19
1>
1C
b101 G
#312800000000
0!
0*
09
0>
0C
#312810000000
1!
1*
b110 6
19
1>
1C
b110 G
#312820000000
0!
0*
09
0>
0C
#312830000000
1!
1*
b111 6
19
1>
1C
b111 G
#312840000000
0!
1"
0*
1+
09
1:
0>
0C
#312850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#312860000000
0!
0*
09
0>
0C
#312870000000
1!
1*
b1 6
19
1>
1C
b1 G
#312880000000
0!
0*
09
0>
0C
#312890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#312900000000
0!
0*
09
0>
0C
#312910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#312920000000
0!
0*
09
0>
0C
#312930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#312940000000
0!
0*
09
0>
0C
#312950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#312960000000
0!
0#
0*
0,
09
0>
0?
0C
#312970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#312980000000
0!
0*
09
0>
0C
#312990000000
1!
1*
19
1>
1C
#313000000000
0!
0*
09
0>
0C
#313010000000
1!
1*
19
1>
1C
#313020000000
0!
0*
09
0>
0C
#313030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#313040000000
0!
0*
09
0>
0C
#313050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#313060000000
0!
0*
09
0>
0C
#313070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#313080000000
0!
0*
09
0>
0C
#313090000000
1!
1*
b10 6
19
1>
1C
b10 G
#313100000000
0!
0*
09
0>
0C
#313110000000
1!
1*
b11 6
19
1>
1C
b11 G
#313120000000
0!
0*
09
0>
0C
#313130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#313140000000
0!
0*
09
0>
0C
#313150000000
1!
1*
b101 6
19
1>
1C
b101 G
#313160000000
0!
0*
09
0>
0C
#313170000000
1!
1*
b110 6
19
1>
1C
b110 G
#313180000000
0!
0*
09
0>
0C
#313190000000
1!
1*
b111 6
19
1>
1C
b111 G
#313200000000
0!
0*
09
0>
0C
#313210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#313220000000
0!
0*
09
0>
0C
#313230000000
1!
1*
b1 6
19
1>
1C
b1 G
#313240000000
0!
0*
09
0>
0C
#313250000000
1!
1*
b10 6
19
1>
1C
b10 G
#313260000000
0!
0*
09
0>
0C
#313270000000
1!
1*
b11 6
19
1>
1C
b11 G
#313280000000
0!
0*
09
0>
0C
#313290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#313300000000
0!
0*
09
0>
0C
#313310000000
1!
1*
b101 6
19
1>
1C
b101 G
#313320000000
0!
0*
09
0>
0C
#313330000000
1!
1*
b110 6
19
1>
1C
b110 G
#313340000000
0!
0*
09
0>
0C
#313350000000
1!
1*
b111 6
19
1>
1C
b111 G
#313360000000
0!
0*
09
0>
0C
#313370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#313380000000
0!
0*
09
0>
0C
#313390000000
1!
1*
b1 6
19
1>
1C
b1 G
#313400000000
0!
0*
09
0>
0C
#313410000000
1!
1*
b10 6
19
1>
1C
b10 G
#313420000000
0!
0*
09
0>
0C
#313430000000
1!
1*
b11 6
19
1>
1C
b11 G
#313440000000
0!
0*
09
0>
0C
#313450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#313460000000
0!
0*
09
0>
0C
#313470000000
1!
1*
b101 6
19
1>
1C
b101 G
#313480000000
0!
0*
09
0>
0C
#313490000000
1!
1*
b110 6
19
1>
1C
b110 G
#313500000000
0!
0*
09
0>
0C
#313510000000
1!
1*
b111 6
19
1>
1C
b111 G
#313520000000
0!
1"
0*
1+
09
1:
0>
0C
#313530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#313540000000
0!
0*
09
0>
0C
#313550000000
1!
1*
b1 6
19
1>
1C
b1 G
#313560000000
0!
0*
09
0>
0C
#313570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#313580000000
0!
0*
09
0>
0C
#313590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#313600000000
0!
0*
09
0>
0C
#313610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#313620000000
0!
0*
09
0>
0C
#313630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#313640000000
0!
0#
0*
0,
09
0>
0?
0C
#313650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#313660000000
0!
0*
09
0>
0C
#313670000000
1!
1*
19
1>
1C
#313680000000
0!
0*
09
0>
0C
#313690000000
1!
1*
19
1>
1C
#313700000000
0!
0*
09
0>
0C
#313710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#313720000000
0!
0*
09
0>
0C
#313730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#313740000000
0!
0*
09
0>
0C
#313750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#313760000000
0!
0*
09
0>
0C
#313770000000
1!
1*
b10 6
19
1>
1C
b10 G
#313780000000
0!
0*
09
0>
0C
#313790000000
1!
1*
b11 6
19
1>
1C
b11 G
#313800000000
0!
0*
09
0>
0C
#313810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#313820000000
0!
0*
09
0>
0C
#313830000000
1!
1*
b101 6
19
1>
1C
b101 G
#313840000000
0!
0*
09
0>
0C
#313850000000
1!
1*
b110 6
19
1>
1C
b110 G
#313860000000
0!
0*
09
0>
0C
#313870000000
1!
1*
b111 6
19
1>
1C
b111 G
#313880000000
0!
0*
09
0>
0C
#313890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#313900000000
0!
0*
09
0>
0C
#313910000000
1!
1*
b1 6
19
1>
1C
b1 G
#313920000000
0!
0*
09
0>
0C
#313930000000
1!
1*
b10 6
19
1>
1C
b10 G
#313940000000
0!
0*
09
0>
0C
#313950000000
1!
1*
b11 6
19
1>
1C
b11 G
#313960000000
0!
0*
09
0>
0C
#313970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#313980000000
0!
0*
09
0>
0C
#313990000000
1!
1*
b101 6
19
1>
1C
b101 G
#314000000000
0!
0*
09
0>
0C
#314010000000
1!
1*
b110 6
19
1>
1C
b110 G
#314020000000
0!
0*
09
0>
0C
#314030000000
1!
1*
b111 6
19
1>
1C
b111 G
#314040000000
0!
0*
09
0>
0C
#314050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#314060000000
0!
0*
09
0>
0C
#314070000000
1!
1*
b1 6
19
1>
1C
b1 G
#314080000000
0!
0*
09
0>
0C
#314090000000
1!
1*
b10 6
19
1>
1C
b10 G
#314100000000
0!
0*
09
0>
0C
#314110000000
1!
1*
b11 6
19
1>
1C
b11 G
#314120000000
0!
0*
09
0>
0C
#314130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#314140000000
0!
0*
09
0>
0C
#314150000000
1!
1*
b101 6
19
1>
1C
b101 G
#314160000000
0!
0*
09
0>
0C
#314170000000
1!
1*
b110 6
19
1>
1C
b110 G
#314180000000
0!
0*
09
0>
0C
#314190000000
1!
1*
b111 6
19
1>
1C
b111 G
#314200000000
0!
1"
0*
1+
09
1:
0>
0C
#314210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#314220000000
0!
0*
09
0>
0C
#314230000000
1!
1*
b1 6
19
1>
1C
b1 G
#314240000000
0!
0*
09
0>
0C
#314250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#314260000000
0!
0*
09
0>
0C
#314270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#314280000000
0!
0*
09
0>
0C
#314290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#314300000000
0!
0*
09
0>
0C
#314310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#314320000000
0!
0#
0*
0,
09
0>
0?
0C
#314330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#314340000000
0!
0*
09
0>
0C
#314350000000
1!
1*
19
1>
1C
#314360000000
0!
0*
09
0>
0C
#314370000000
1!
1*
19
1>
1C
#314380000000
0!
0*
09
0>
0C
#314390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#314400000000
0!
0*
09
0>
0C
#314410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#314420000000
0!
0*
09
0>
0C
#314430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#314440000000
0!
0*
09
0>
0C
#314450000000
1!
1*
b10 6
19
1>
1C
b10 G
#314460000000
0!
0*
09
0>
0C
#314470000000
1!
1*
b11 6
19
1>
1C
b11 G
#314480000000
0!
0*
09
0>
0C
#314490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#314500000000
0!
0*
09
0>
0C
#314510000000
1!
1*
b101 6
19
1>
1C
b101 G
#314520000000
0!
0*
09
0>
0C
#314530000000
1!
1*
b110 6
19
1>
1C
b110 G
#314540000000
0!
0*
09
0>
0C
#314550000000
1!
1*
b111 6
19
1>
1C
b111 G
#314560000000
0!
0*
09
0>
0C
#314570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#314580000000
0!
0*
09
0>
0C
#314590000000
1!
1*
b1 6
19
1>
1C
b1 G
#314600000000
0!
0*
09
0>
0C
#314610000000
1!
1*
b10 6
19
1>
1C
b10 G
#314620000000
0!
0*
09
0>
0C
#314630000000
1!
1*
b11 6
19
1>
1C
b11 G
#314640000000
0!
0*
09
0>
0C
#314650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#314660000000
0!
0*
09
0>
0C
#314670000000
1!
1*
b101 6
19
1>
1C
b101 G
#314680000000
0!
0*
09
0>
0C
#314690000000
1!
1*
b110 6
19
1>
1C
b110 G
#314700000000
0!
0*
09
0>
0C
#314710000000
1!
1*
b111 6
19
1>
1C
b111 G
#314720000000
0!
0*
09
0>
0C
#314730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#314740000000
0!
0*
09
0>
0C
#314750000000
1!
1*
b1 6
19
1>
1C
b1 G
#314760000000
0!
0*
09
0>
0C
#314770000000
1!
1*
b10 6
19
1>
1C
b10 G
#314780000000
0!
0*
09
0>
0C
#314790000000
1!
1*
b11 6
19
1>
1C
b11 G
#314800000000
0!
0*
09
0>
0C
#314810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#314820000000
0!
0*
09
0>
0C
#314830000000
1!
1*
b101 6
19
1>
1C
b101 G
#314840000000
0!
0*
09
0>
0C
#314850000000
1!
1*
b110 6
19
1>
1C
b110 G
#314860000000
0!
0*
09
0>
0C
#314870000000
1!
1*
b111 6
19
1>
1C
b111 G
#314880000000
0!
1"
0*
1+
09
1:
0>
0C
#314890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#314900000000
0!
0*
09
0>
0C
#314910000000
1!
1*
b1 6
19
1>
1C
b1 G
#314920000000
0!
0*
09
0>
0C
#314930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#314940000000
0!
0*
09
0>
0C
#314950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#314960000000
0!
0*
09
0>
0C
#314970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#314980000000
0!
0*
09
0>
0C
#314990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#315000000000
0!
0#
0*
0,
09
0>
0?
0C
#315010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#315020000000
0!
0*
09
0>
0C
#315030000000
1!
1*
19
1>
1C
#315040000000
0!
0*
09
0>
0C
#315050000000
1!
1*
19
1>
1C
#315060000000
0!
0*
09
0>
0C
#315070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#315080000000
0!
0*
09
0>
0C
#315090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#315100000000
0!
0*
09
0>
0C
#315110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#315120000000
0!
0*
09
0>
0C
#315130000000
1!
1*
b10 6
19
1>
1C
b10 G
#315140000000
0!
0*
09
0>
0C
#315150000000
1!
1*
b11 6
19
1>
1C
b11 G
#315160000000
0!
0*
09
0>
0C
#315170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#315180000000
0!
0*
09
0>
0C
#315190000000
1!
1*
b101 6
19
1>
1C
b101 G
#315200000000
0!
0*
09
0>
0C
#315210000000
1!
1*
b110 6
19
1>
1C
b110 G
#315220000000
0!
0*
09
0>
0C
#315230000000
1!
1*
b111 6
19
1>
1C
b111 G
#315240000000
0!
0*
09
0>
0C
#315250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#315260000000
0!
0*
09
0>
0C
#315270000000
1!
1*
b1 6
19
1>
1C
b1 G
#315280000000
0!
0*
09
0>
0C
#315290000000
1!
1*
b10 6
19
1>
1C
b10 G
#315300000000
0!
0*
09
0>
0C
#315310000000
1!
1*
b11 6
19
1>
1C
b11 G
#315320000000
0!
0*
09
0>
0C
#315330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#315340000000
0!
0*
09
0>
0C
#315350000000
1!
1*
b101 6
19
1>
1C
b101 G
#315360000000
0!
0*
09
0>
0C
#315370000000
1!
1*
b110 6
19
1>
1C
b110 G
#315380000000
0!
0*
09
0>
0C
#315390000000
1!
1*
b111 6
19
1>
1C
b111 G
#315400000000
0!
0*
09
0>
0C
#315410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#315420000000
0!
0*
09
0>
0C
#315430000000
1!
1*
b1 6
19
1>
1C
b1 G
#315440000000
0!
0*
09
0>
0C
#315450000000
1!
1*
b10 6
19
1>
1C
b10 G
#315460000000
0!
0*
09
0>
0C
#315470000000
1!
1*
b11 6
19
1>
1C
b11 G
#315480000000
0!
0*
09
0>
0C
#315490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#315500000000
0!
0*
09
0>
0C
#315510000000
1!
1*
b101 6
19
1>
1C
b101 G
#315520000000
0!
0*
09
0>
0C
#315530000000
1!
1*
b110 6
19
1>
1C
b110 G
#315540000000
0!
0*
09
0>
0C
#315550000000
1!
1*
b111 6
19
1>
1C
b111 G
#315560000000
0!
1"
0*
1+
09
1:
0>
0C
#315570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#315580000000
0!
0*
09
0>
0C
#315590000000
1!
1*
b1 6
19
1>
1C
b1 G
#315600000000
0!
0*
09
0>
0C
#315610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#315620000000
0!
0*
09
0>
0C
#315630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#315640000000
0!
0*
09
0>
0C
#315650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#315660000000
0!
0*
09
0>
0C
#315670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#315680000000
0!
0#
0*
0,
09
0>
0?
0C
#315690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#315700000000
0!
0*
09
0>
0C
#315710000000
1!
1*
19
1>
1C
#315720000000
0!
0*
09
0>
0C
#315730000000
1!
1*
19
1>
1C
#315740000000
0!
0*
09
0>
0C
#315750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#315760000000
0!
0*
09
0>
0C
#315770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#315780000000
0!
0*
09
0>
0C
#315790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#315800000000
0!
0*
09
0>
0C
#315810000000
1!
1*
b10 6
19
1>
1C
b10 G
#315820000000
0!
0*
09
0>
0C
#315830000000
1!
1*
b11 6
19
1>
1C
b11 G
#315840000000
0!
0*
09
0>
0C
#315850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#315860000000
0!
0*
09
0>
0C
#315870000000
1!
1*
b101 6
19
1>
1C
b101 G
#315880000000
0!
0*
09
0>
0C
#315890000000
1!
1*
b110 6
19
1>
1C
b110 G
#315900000000
0!
0*
09
0>
0C
#315910000000
1!
1*
b111 6
19
1>
1C
b111 G
#315920000000
0!
0*
09
0>
0C
#315930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#315940000000
0!
0*
09
0>
0C
#315950000000
1!
1*
b1 6
19
1>
1C
b1 G
#315960000000
0!
0*
09
0>
0C
#315970000000
1!
1*
b10 6
19
1>
1C
b10 G
#315980000000
0!
0*
09
0>
0C
#315990000000
1!
1*
b11 6
19
1>
1C
b11 G
#316000000000
0!
0*
09
0>
0C
#316010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#316020000000
0!
0*
09
0>
0C
#316030000000
1!
1*
b101 6
19
1>
1C
b101 G
#316040000000
0!
0*
09
0>
0C
#316050000000
1!
1*
b110 6
19
1>
1C
b110 G
#316060000000
0!
0*
09
0>
0C
#316070000000
1!
1*
b111 6
19
1>
1C
b111 G
#316080000000
0!
0*
09
0>
0C
#316090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#316100000000
0!
0*
09
0>
0C
#316110000000
1!
1*
b1 6
19
1>
1C
b1 G
#316120000000
0!
0*
09
0>
0C
#316130000000
1!
1*
b10 6
19
1>
1C
b10 G
#316140000000
0!
0*
09
0>
0C
#316150000000
1!
1*
b11 6
19
1>
1C
b11 G
#316160000000
0!
0*
09
0>
0C
#316170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#316180000000
0!
0*
09
0>
0C
#316190000000
1!
1*
b101 6
19
1>
1C
b101 G
#316200000000
0!
0*
09
0>
0C
#316210000000
1!
1*
b110 6
19
1>
1C
b110 G
#316220000000
0!
0*
09
0>
0C
#316230000000
1!
1*
b111 6
19
1>
1C
b111 G
#316240000000
0!
1"
0*
1+
09
1:
0>
0C
#316250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#316260000000
0!
0*
09
0>
0C
#316270000000
1!
1*
b1 6
19
1>
1C
b1 G
#316280000000
0!
0*
09
0>
0C
#316290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#316300000000
0!
0*
09
0>
0C
#316310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#316320000000
0!
0*
09
0>
0C
#316330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#316340000000
0!
0*
09
0>
0C
#316350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#316360000000
0!
0#
0*
0,
09
0>
0?
0C
#316370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#316380000000
0!
0*
09
0>
0C
#316390000000
1!
1*
19
1>
1C
#316400000000
0!
0*
09
0>
0C
#316410000000
1!
1*
19
1>
1C
#316420000000
0!
0*
09
0>
0C
#316430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#316440000000
0!
0*
09
0>
0C
#316450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#316460000000
0!
0*
09
0>
0C
#316470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#316480000000
0!
0*
09
0>
0C
#316490000000
1!
1*
b10 6
19
1>
1C
b10 G
#316500000000
0!
0*
09
0>
0C
#316510000000
1!
1*
b11 6
19
1>
1C
b11 G
#316520000000
0!
0*
09
0>
0C
#316530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#316540000000
0!
0*
09
0>
0C
#316550000000
1!
1*
b101 6
19
1>
1C
b101 G
#316560000000
0!
0*
09
0>
0C
#316570000000
1!
1*
b110 6
19
1>
1C
b110 G
#316580000000
0!
0*
09
0>
0C
#316590000000
1!
1*
b111 6
19
1>
1C
b111 G
#316600000000
0!
0*
09
0>
0C
#316610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#316620000000
0!
0*
09
0>
0C
#316630000000
1!
1*
b1 6
19
1>
1C
b1 G
#316640000000
0!
0*
09
0>
0C
#316650000000
1!
1*
b10 6
19
1>
1C
b10 G
#316660000000
0!
0*
09
0>
0C
#316670000000
1!
1*
b11 6
19
1>
1C
b11 G
#316680000000
0!
0*
09
0>
0C
#316690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#316700000000
0!
0*
09
0>
0C
#316710000000
1!
1*
b101 6
19
1>
1C
b101 G
#316720000000
0!
0*
09
0>
0C
#316730000000
1!
1*
b110 6
19
1>
1C
b110 G
#316740000000
0!
0*
09
0>
0C
#316750000000
1!
1*
b111 6
19
1>
1C
b111 G
#316760000000
0!
0*
09
0>
0C
#316770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#316780000000
0!
0*
09
0>
0C
#316790000000
1!
1*
b1 6
19
1>
1C
b1 G
#316800000000
0!
0*
09
0>
0C
#316810000000
1!
1*
b10 6
19
1>
1C
b10 G
#316820000000
0!
0*
09
0>
0C
#316830000000
1!
1*
b11 6
19
1>
1C
b11 G
#316840000000
0!
0*
09
0>
0C
#316850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#316860000000
0!
0*
09
0>
0C
#316870000000
1!
1*
b101 6
19
1>
1C
b101 G
#316880000000
0!
0*
09
0>
0C
#316890000000
1!
1*
b110 6
19
1>
1C
b110 G
#316900000000
0!
0*
09
0>
0C
#316910000000
1!
1*
b111 6
19
1>
1C
b111 G
#316920000000
0!
1"
0*
1+
09
1:
0>
0C
#316930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#316940000000
0!
0*
09
0>
0C
#316950000000
1!
1*
b1 6
19
1>
1C
b1 G
#316960000000
0!
0*
09
0>
0C
#316970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#316980000000
0!
0*
09
0>
0C
#316990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#317000000000
0!
0*
09
0>
0C
#317010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#317020000000
0!
0*
09
0>
0C
#317030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#317040000000
0!
0#
0*
0,
09
0>
0?
0C
#317050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#317060000000
0!
0*
09
0>
0C
#317070000000
1!
1*
19
1>
1C
#317080000000
0!
0*
09
0>
0C
#317090000000
1!
1*
19
1>
1C
#317100000000
0!
0*
09
0>
0C
#317110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#317120000000
0!
0*
09
0>
0C
#317130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#317140000000
0!
0*
09
0>
0C
#317150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#317160000000
0!
0*
09
0>
0C
#317170000000
1!
1*
b10 6
19
1>
1C
b10 G
#317180000000
0!
0*
09
0>
0C
#317190000000
1!
1*
b11 6
19
1>
1C
b11 G
#317200000000
0!
0*
09
0>
0C
#317210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#317220000000
0!
0*
09
0>
0C
#317230000000
1!
1*
b101 6
19
1>
1C
b101 G
#317240000000
0!
0*
09
0>
0C
#317250000000
1!
1*
b110 6
19
1>
1C
b110 G
#317260000000
0!
0*
09
0>
0C
#317270000000
1!
1*
b111 6
19
1>
1C
b111 G
#317280000000
0!
0*
09
0>
0C
#317290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#317300000000
0!
0*
09
0>
0C
#317310000000
1!
1*
b1 6
19
1>
1C
b1 G
#317320000000
0!
0*
09
0>
0C
#317330000000
1!
1*
b10 6
19
1>
1C
b10 G
#317340000000
0!
0*
09
0>
0C
#317350000000
1!
1*
b11 6
19
1>
1C
b11 G
#317360000000
0!
0*
09
0>
0C
#317370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#317380000000
0!
0*
09
0>
0C
#317390000000
1!
1*
b101 6
19
1>
1C
b101 G
#317400000000
0!
0*
09
0>
0C
#317410000000
1!
1*
b110 6
19
1>
1C
b110 G
#317420000000
0!
0*
09
0>
0C
#317430000000
1!
1*
b111 6
19
1>
1C
b111 G
#317440000000
0!
0*
09
0>
0C
#317450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#317460000000
0!
0*
09
0>
0C
#317470000000
1!
1*
b1 6
19
1>
1C
b1 G
#317480000000
0!
0*
09
0>
0C
#317490000000
1!
1*
b10 6
19
1>
1C
b10 G
#317500000000
0!
0*
09
0>
0C
#317510000000
1!
1*
b11 6
19
1>
1C
b11 G
#317520000000
0!
0*
09
0>
0C
#317530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#317540000000
0!
0*
09
0>
0C
#317550000000
1!
1*
b101 6
19
1>
1C
b101 G
#317560000000
0!
0*
09
0>
0C
#317570000000
1!
1*
b110 6
19
1>
1C
b110 G
#317580000000
0!
0*
09
0>
0C
#317590000000
1!
1*
b111 6
19
1>
1C
b111 G
#317600000000
0!
1"
0*
1+
09
1:
0>
0C
#317610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#317620000000
0!
0*
09
0>
0C
#317630000000
1!
1*
b1 6
19
1>
1C
b1 G
#317640000000
0!
0*
09
0>
0C
#317650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#317660000000
0!
0*
09
0>
0C
#317670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#317680000000
0!
0*
09
0>
0C
#317690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#317700000000
0!
0*
09
0>
0C
#317710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#317720000000
0!
0#
0*
0,
09
0>
0?
0C
#317730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#317740000000
0!
0*
09
0>
0C
#317750000000
1!
1*
19
1>
1C
#317760000000
0!
0*
09
0>
0C
#317770000000
1!
1*
19
1>
1C
#317780000000
0!
0*
09
0>
0C
#317790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#317800000000
0!
0*
09
0>
0C
#317810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#317820000000
0!
0*
09
0>
0C
#317830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#317840000000
0!
0*
09
0>
0C
#317850000000
1!
1*
b10 6
19
1>
1C
b10 G
#317860000000
0!
0*
09
0>
0C
#317870000000
1!
1*
b11 6
19
1>
1C
b11 G
#317880000000
0!
0*
09
0>
0C
#317890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#317900000000
0!
0*
09
0>
0C
#317910000000
1!
1*
b101 6
19
1>
1C
b101 G
#317920000000
0!
0*
09
0>
0C
#317930000000
1!
1*
b110 6
19
1>
1C
b110 G
#317940000000
0!
0*
09
0>
0C
#317950000000
1!
1*
b111 6
19
1>
1C
b111 G
#317960000000
0!
0*
09
0>
0C
#317970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#317980000000
0!
0*
09
0>
0C
#317990000000
1!
1*
b1 6
19
1>
1C
b1 G
#318000000000
0!
0*
09
0>
0C
#318010000000
1!
1*
b10 6
19
1>
1C
b10 G
#318020000000
0!
0*
09
0>
0C
#318030000000
1!
1*
b11 6
19
1>
1C
b11 G
#318040000000
0!
0*
09
0>
0C
#318050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#318060000000
0!
0*
09
0>
0C
#318070000000
1!
1*
b101 6
19
1>
1C
b101 G
#318080000000
0!
0*
09
0>
0C
#318090000000
1!
1*
b110 6
19
1>
1C
b110 G
#318100000000
0!
0*
09
0>
0C
#318110000000
1!
1*
b111 6
19
1>
1C
b111 G
#318120000000
0!
0*
09
0>
0C
#318130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#318140000000
0!
0*
09
0>
0C
#318150000000
1!
1*
b1 6
19
1>
1C
b1 G
#318160000000
0!
0*
09
0>
0C
#318170000000
1!
1*
b10 6
19
1>
1C
b10 G
#318180000000
0!
0*
09
0>
0C
#318190000000
1!
1*
b11 6
19
1>
1C
b11 G
#318200000000
0!
0*
09
0>
0C
#318210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#318220000000
0!
0*
09
0>
0C
#318230000000
1!
1*
b101 6
19
1>
1C
b101 G
#318240000000
0!
0*
09
0>
0C
#318250000000
1!
1*
b110 6
19
1>
1C
b110 G
#318260000000
0!
0*
09
0>
0C
#318270000000
1!
1*
b111 6
19
1>
1C
b111 G
#318280000000
0!
1"
0*
1+
09
1:
0>
0C
#318290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#318300000000
0!
0*
09
0>
0C
#318310000000
1!
1*
b1 6
19
1>
1C
b1 G
#318320000000
0!
0*
09
0>
0C
#318330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#318340000000
0!
0*
09
0>
0C
#318350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#318360000000
0!
0*
09
0>
0C
#318370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#318380000000
0!
0*
09
0>
0C
#318390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#318400000000
0!
0#
0*
0,
09
0>
0?
0C
#318410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#318420000000
0!
0*
09
0>
0C
#318430000000
1!
1*
19
1>
1C
#318440000000
0!
0*
09
0>
0C
#318450000000
1!
1*
19
1>
1C
#318460000000
0!
0*
09
0>
0C
#318470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#318480000000
0!
0*
09
0>
0C
#318490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#318500000000
0!
0*
09
0>
0C
#318510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#318520000000
0!
0*
09
0>
0C
#318530000000
1!
1*
b10 6
19
1>
1C
b10 G
#318540000000
0!
0*
09
0>
0C
#318550000000
1!
1*
b11 6
19
1>
1C
b11 G
#318560000000
0!
0*
09
0>
0C
#318570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#318580000000
0!
0*
09
0>
0C
#318590000000
1!
1*
b101 6
19
1>
1C
b101 G
#318600000000
0!
0*
09
0>
0C
#318610000000
1!
1*
b110 6
19
1>
1C
b110 G
#318620000000
0!
0*
09
0>
0C
#318630000000
1!
1*
b111 6
19
1>
1C
b111 G
#318640000000
0!
0*
09
0>
0C
#318650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#318660000000
0!
0*
09
0>
0C
#318670000000
1!
1*
b1 6
19
1>
1C
b1 G
#318680000000
0!
0*
09
0>
0C
#318690000000
1!
1*
b10 6
19
1>
1C
b10 G
#318700000000
0!
0*
09
0>
0C
#318710000000
1!
1*
b11 6
19
1>
1C
b11 G
#318720000000
0!
0*
09
0>
0C
#318730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#318740000000
0!
0*
09
0>
0C
#318750000000
1!
1*
b101 6
19
1>
1C
b101 G
#318760000000
0!
0*
09
0>
0C
#318770000000
1!
1*
b110 6
19
1>
1C
b110 G
#318780000000
0!
0*
09
0>
0C
#318790000000
1!
1*
b111 6
19
1>
1C
b111 G
#318800000000
0!
0*
09
0>
0C
#318810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#318820000000
0!
0*
09
0>
0C
#318830000000
1!
1*
b1 6
19
1>
1C
b1 G
#318840000000
0!
0*
09
0>
0C
#318850000000
1!
1*
b10 6
19
1>
1C
b10 G
#318860000000
0!
0*
09
0>
0C
#318870000000
1!
1*
b11 6
19
1>
1C
b11 G
#318880000000
0!
0*
09
0>
0C
#318890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#318900000000
0!
0*
09
0>
0C
#318910000000
1!
1*
b101 6
19
1>
1C
b101 G
#318920000000
0!
0*
09
0>
0C
#318930000000
1!
1*
b110 6
19
1>
1C
b110 G
#318940000000
0!
0*
09
0>
0C
#318950000000
1!
1*
b111 6
19
1>
1C
b111 G
#318960000000
0!
1"
0*
1+
09
1:
0>
0C
#318970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#318980000000
0!
0*
09
0>
0C
#318990000000
1!
1*
b1 6
19
1>
1C
b1 G
#319000000000
0!
0*
09
0>
0C
#319010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#319020000000
0!
0*
09
0>
0C
#319030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#319040000000
0!
0*
09
0>
0C
#319050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#319060000000
0!
0*
09
0>
0C
#319070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#319080000000
0!
0#
0*
0,
09
0>
0?
0C
#319090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#319100000000
0!
0*
09
0>
0C
#319110000000
1!
1*
19
1>
1C
#319120000000
0!
0*
09
0>
0C
#319130000000
1!
1*
19
1>
1C
#319140000000
0!
0*
09
0>
0C
#319150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#319160000000
0!
0*
09
0>
0C
#319170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#319180000000
0!
0*
09
0>
0C
#319190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#319200000000
0!
0*
09
0>
0C
#319210000000
1!
1*
b10 6
19
1>
1C
b10 G
#319220000000
0!
0*
09
0>
0C
#319230000000
1!
1*
b11 6
19
1>
1C
b11 G
#319240000000
0!
0*
09
0>
0C
#319250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#319260000000
0!
0*
09
0>
0C
#319270000000
1!
1*
b101 6
19
1>
1C
b101 G
#319280000000
0!
0*
09
0>
0C
#319290000000
1!
1*
b110 6
19
1>
1C
b110 G
#319300000000
0!
0*
09
0>
0C
#319310000000
1!
1*
b111 6
19
1>
1C
b111 G
#319320000000
0!
0*
09
0>
0C
#319330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#319340000000
0!
0*
09
0>
0C
#319350000000
1!
1*
b1 6
19
1>
1C
b1 G
#319360000000
0!
0*
09
0>
0C
#319370000000
1!
1*
b10 6
19
1>
1C
b10 G
#319380000000
0!
0*
09
0>
0C
#319390000000
1!
1*
b11 6
19
1>
1C
b11 G
#319400000000
0!
0*
09
0>
0C
#319410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#319420000000
0!
0*
09
0>
0C
#319430000000
1!
1*
b101 6
19
1>
1C
b101 G
#319440000000
0!
0*
09
0>
0C
#319450000000
1!
1*
b110 6
19
1>
1C
b110 G
#319460000000
0!
0*
09
0>
0C
#319470000000
1!
1*
b111 6
19
1>
1C
b111 G
#319480000000
0!
0*
09
0>
0C
#319490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#319500000000
0!
0*
09
0>
0C
#319510000000
1!
1*
b1 6
19
1>
1C
b1 G
#319520000000
0!
0*
09
0>
0C
#319530000000
1!
1*
b10 6
19
1>
1C
b10 G
#319540000000
0!
0*
09
0>
0C
#319550000000
1!
1*
b11 6
19
1>
1C
b11 G
#319560000000
0!
0*
09
0>
0C
#319570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#319580000000
0!
0*
09
0>
0C
#319590000000
1!
1*
b101 6
19
1>
1C
b101 G
#319600000000
0!
0*
09
0>
0C
#319610000000
1!
1*
b110 6
19
1>
1C
b110 G
#319620000000
0!
0*
09
0>
0C
#319630000000
1!
1*
b111 6
19
1>
1C
b111 G
#319640000000
0!
1"
0*
1+
09
1:
0>
0C
#319650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#319660000000
0!
0*
09
0>
0C
#319670000000
1!
1*
b1 6
19
1>
1C
b1 G
#319680000000
0!
0*
09
0>
0C
#319690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#319700000000
0!
0*
09
0>
0C
#319710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#319720000000
0!
0*
09
0>
0C
#319730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#319740000000
0!
0*
09
0>
0C
#319750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#319760000000
0!
0#
0*
0,
09
0>
0?
0C
#319770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#319780000000
0!
0*
09
0>
0C
#319790000000
1!
1*
19
1>
1C
#319800000000
0!
0*
09
0>
0C
#319810000000
1!
1*
19
1>
1C
#319820000000
0!
0*
09
0>
0C
#319830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#319840000000
0!
0*
09
0>
0C
#319850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#319860000000
0!
0*
09
0>
0C
#319870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#319880000000
0!
0*
09
0>
0C
#319890000000
1!
1*
b10 6
19
1>
1C
b10 G
#319900000000
0!
0*
09
0>
0C
#319910000000
1!
1*
b11 6
19
1>
1C
b11 G
#319920000000
0!
0*
09
0>
0C
#319930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#319940000000
0!
0*
09
0>
0C
#319950000000
1!
1*
b101 6
19
1>
1C
b101 G
#319960000000
0!
0*
09
0>
0C
#319970000000
1!
1*
b110 6
19
1>
1C
b110 G
#319980000000
0!
0*
09
0>
0C
#319990000000
1!
1*
b111 6
19
1>
1C
b111 G
#320000000000
0!
0*
09
0>
0C
#320010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#320020000000
0!
0*
09
0>
0C
#320030000000
1!
1*
b1 6
19
1>
1C
b1 G
#320040000000
0!
0*
09
0>
0C
#320050000000
1!
1*
b10 6
19
1>
1C
b10 G
#320060000000
0!
0*
09
0>
0C
#320070000000
1!
1*
b11 6
19
1>
1C
b11 G
#320080000000
0!
0*
09
0>
0C
#320090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#320100000000
0!
0*
09
0>
0C
#320110000000
1!
1*
b101 6
19
1>
1C
b101 G
#320120000000
0!
0*
09
0>
0C
#320130000000
1!
1*
b110 6
19
1>
1C
b110 G
#320140000000
0!
0*
09
0>
0C
#320150000000
1!
1*
b111 6
19
1>
1C
b111 G
#320160000000
0!
0*
09
0>
0C
#320170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#320180000000
0!
0*
09
0>
0C
#320190000000
1!
1*
b1 6
19
1>
1C
b1 G
#320200000000
0!
0*
09
0>
0C
#320210000000
1!
1*
b10 6
19
1>
1C
b10 G
#320220000000
0!
0*
09
0>
0C
#320230000000
1!
1*
b11 6
19
1>
1C
b11 G
#320240000000
0!
0*
09
0>
0C
#320250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#320260000000
0!
0*
09
0>
0C
#320270000000
1!
1*
b101 6
19
1>
1C
b101 G
#320280000000
0!
0*
09
0>
0C
#320290000000
1!
1*
b110 6
19
1>
1C
b110 G
#320300000000
0!
0*
09
0>
0C
#320310000000
1!
1*
b111 6
19
1>
1C
b111 G
#320320000000
0!
1"
0*
1+
09
1:
0>
0C
#320330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#320340000000
0!
0*
09
0>
0C
#320350000000
1!
1*
b1 6
19
1>
1C
b1 G
#320360000000
0!
0*
09
0>
0C
#320370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#320380000000
0!
0*
09
0>
0C
#320390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#320400000000
0!
0*
09
0>
0C
#320410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#320420000000
0!
0*
09
0>
0C
#320430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#320440000000
0!
0#
0*
0,
09
0>
0?
0C
#320450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#320460000000
0!
0*
09
0>
0C
#320470000000
1!
1*
19
1>
1C
#320480000000
0!
0*
09
0>
0C
#320490000000
1!
1*
19
1>
1C
#320500000000
0!
0*
09
0>
0C
#320510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#320520000000
0!
0*
09
0>
0C
#320530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#320540000000
0!
0*
09
0>
0C
#320550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#320560000000
0!
0*
09
0>
0C
#320570000000
1!
1*
b10 6
19
1>
1C
b10 G
#320580000000
0!
0*
09
0>
0C
#320590000000
1!
1*
b11 6
19
1>
1C
b11 G
#320600000000
0!
0*
09
0>
0C
#320610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#320620000000
0!
0*
09
0>
0C
#320630000000
1!
1*
b101 6
19
1>
1C
b101 G
#320640000000
0!
0*
09
0>
0C
#320650000000
1!
1*
b110 6
19
1>
1C
b110 G
#320660000000
0!
0*
09
0>
0C
#320670000000
1!
1*
b111 6
19
1>
1C
b111 G
#320680000000
0!
0*
09
0>
0C
#320690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#320700000000
0!
0*
09
0>
0C
#320710000000
1!
1*
b1 6
19
1>
1C
b1 G
#320720000000
0!
0*
09
0>
0C
#320730000000
1!
1*
b10 6
19
1>
1C
b10 G
#320740000000
0!
0*
09
0>
0C
#320750000000
1!
1*
b11 6
19
1>
1C
b11 G
#320760000000
0!
0*
09
0>
0C
#320770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#320780000000
0!
0*
09
0>
0C
#320790000000
1!
1*
b101 6
19
1>
1C
b101 G
#320800000000
0!
0*
09
0>
0C
#320810000000
1!
1*
b110 6
19
1>
1C
b110 G
#320820000000
0!
0*
09
0>
0C
#320830000000
1!
1*
b111 6
19
1>
1C
b111 G
#320840000000
0!
0*
09
0>
0C
#320850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#320860000000
0!
0*
09
0>
0C
#320870000000
1!
1*
b1 6
19
1>
1C
b1 G
#320880000000
0!
0*
09
0>
0C
#320890000000
1!
1*
b10 6
19
1>
1C
b10 G
#320900000000
0!
0*
09
0>
0C
#320910000000
1!
1*
b11 6
19
1>
1C
b11 G
#320920000000
0!
0*
09
0>
0C
#320930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#320940000000
0!
0*
09
0>
0C
#320950000000
1!
1*
b101 6
19
1>
1C
b101 G
#320960000000
0!
0*
09
0>
0C
#320970000000
1!
1*
b110 6
19
1>
1C
b110 G
#320980000000
0!
0*
09
0>
0C
#320990000000
1!
1*
b111 6
19
1>
1C
b111 G
#321000000000
0!
1"
0*
1+
09
1:
0>
0C
#321010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#321020000000
0!
0*
09
0>
0C
#321030000000
1!
1*
b1 6
19
1>
1C
b1 G
#321040000000
0!
0*
09
0>
0C
#321050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#321060000000
0!
0*
09
0>
0C
#321070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#321080000000
0!
0*
09
0>
0C
#321090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#321100000000
0!
0*
09
0>
0C
#321110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#321120000000
0!
0#
0*
0,
09
0>
0?
0C
#321130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#321140000000
0!
0*
09
0>
0C
#321150000000
1!
1*
19
1>
1C
#321160000000
0!
0*
09
0>
0C
#321170000000
1!
1*
19
1>
1C
#321180000000
0!
0*
09
0>
0C
#321190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#321200000000
0!
0*
09
0>
0C
#321210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#321220000000
0!
0*
09
0>
0C
#321230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#321240000000
0!
0*
09
0>
0C
#321250000000
1!
1*
b10 6
19
1>
1C
b10 G
#321260000000
0!
0*
09
0>
0C
#321270000000
1!
1*
b11 6
19
1>
1C
b11 G
#321280000000
0!
0*
09
0>
0C
#321290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#321300000000
0!
0*
09
0>
0C
#321310000000
1!
1*
b101 6
19
1>
1C
b101 G
#321320000000
0!
0*
09
0>
0C
#321330000000
1!
1*
b110 6
19
1>
1C
b110 G
#321340000000
0!
0*
09
0>
0C
#321350000000
1!
1*
b111 6
19
1>
1C
b111 G
#321360000000
0!
0*
09
0>
0C
#321370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#321380000000
0!
0*
09
0>
0C
#321390000000
1!
1*
b1 6
19
1>
1C
b1 G
#321400000000
0!
0*
09
0>
0C
#321410000000
1!
1*
b10 6
19
1>
1C
b10 G
#321420000000
0!
0*
09
0>
0C
#321430000000
1!
1*
b11 6
19
1>
1C
b11 G
#321440000000
0!
0*
09
0>
0C
#321450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#321460000000
0!
0*
09
0>
0C
#321470000000
1!
1*
b101 6
19
1>
1C
b101 G
#321480000000
0!
0*
09
0>
0C
#321490000000
1!
1*
b110 6
19
1>
1C
b110 G
#321500000000
0!
0*
09
0>
0C
#321510000000
1!
1*
b111 6
19
1>
1C
b111 G
#321520000000
0!
0*
09
0>
0C
#321530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#321540000000
0!
0*
09
0>
0C
#321550000000
1!
1*
b1 6
19
1>
1C
b1 G
#321560000000
0!
0*
09
0>
0C
#321570000000
1!
1*
b10 6
19
1>
1C
b10 G
#321580000000
0!
0*
09
0>
0C
#321590000000
1!
1*
b11 6
19
1>
1C
b11 G
#321600000000
0!
0*
09
0>
0C
#321610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#321620000000
0!
0*
09
0>
0C
#321630000000
1!
1*
b101 6
19
1>
1C
b101 G
#321640000000
0!
0*
09
0>
0C
#321650000000
1!
1*
b110 6
19
1>
1C
b110 G
#321660000000
0!
0*
09
0>
0C
#321670000000
1!
1*
b111 6
19
1>
1C
b111 G
#321680000000
0!
1"
0*
1+
09
1:
0>
0C
#321690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#321700000000
0!
0*
09
0>
0C
#321710000000
1!
1*
b1 6
19
1>
1C
b1 G
#321720000000
0!
0*
09
0>
0C
#321730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#321740000000
0!
0*
09
0>
0C
#321750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#321760000000
0!
0*
09
0>
0C
#321770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#321780000000
0!
0*
09
0>
0C
#321790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#321800000000
0!
0#
0*
0,
09
0>
0?
0C
#321810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#321820000000
0!
0*
09
0>
0C
#321830000000
1!
1*
19
1>
1C
#321840000000
0!
0*
09
0>
0C
#321850000000
1!
1*
19
1>
1C
#321860000000
0!
0*
09
0>
0C
#321870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#321880000000
0!
0*
09
0>
0C
#321890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#321900000000
0!
0*
09
0>
0C
#321910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#321920000000
0!
0*
09
0>
0C
#321930000000
1!
1*
b10 6
19
1>
1C
b10 G
#321940000000
0!
0*
09
0>
0C
#321950000000
1!
1*
b11 6
19
1>
1C
b11 G
#321960000000
0!
0*
09
0>
0C
#321970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#321980000000
0!
0*
09
0>
0C
#321990000000
1!
1*
b101 6
19
1>
1C
b101 G
#322000000000
0!
0*
09
0>
0C
#322010000000
1!
1*
b110 6
19
1>
1C
b110 G
#322020000000
0!
0*
09
0>
0C
#322030000000
1!
1*
b111 6
19
1>
1C
b111 G
#322040000000
0!
0*
09
0>
0C
#322050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#322060000000
0!
0*
09
0>
0C
#322070000000
1!
1*
b1 6
19
1>
1C
b1 G
#322080000000
0!
0*
09
0>
0C
#322090000000
1!
1*
b10 6
19
1>
1C
b10 G
#322100000000
0!
0*
09
0>
0C
#322110000000
1!
1*
b11 6
19
1>
1C
b11 G
#322120000000
0!
0*
09
0>
0C
#322130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#322140000000
0!
0*
09
0>
0C
#322150000000
1!
1*
b101 6
19
1>
1C
b101 G
#322160000000
0!
0*
09
0>
0C
#322170000000
1!
1*
b110 6
19
1>
1C
b110 G
#322180000000
0!
0*
09
0>
0C
#322190000000
1!
1*
b111 6
19
1>
1C
b111 G
#322200000000
0!
0*
09
0>
0C
#322210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#322220000000
0!
0*
09
0>
0C
#322230000000
1!
1*
b1 6
19
1>
1C
b1 G
#322240000000
0!
0*
09
0>
0C
#322250000000
1!
1*
b10 6
19
1>
1C
b10 G
#322260000000
0!
0*
09
0>
0C
#322270000000
1!
1*
b11 6
19
1>
1C
b11 G
#322280000000
0!
0*
09
0>
0C
#322290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#322300000000
0!
0*
09
0>
0C
#322310000000
1!
1*
b101 6
19
1>
1C
b101 G
#322320000000
0!
0*
09
0>
0C
#322330000000
1!
1*
b110 6
19
1>
1C
b110 G
#322340000000
0!
0*
09
0>
0C
#322350000000
1!
1*
b111 6
19
1>
1C
b111 G
#322360000000
0!
1"
0*
1+
09
1:
0>
0C
#322370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#322380000000
0!
0*
09
0>
0C
#322390000000
1!
1*
b1 6
19
1>
1C
b1 G
#322400000000
0!
0*
09
0>
0C
#322410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#322420000000
0!
0*
09
0>
0C
#322430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#322440000000
0!
0*
09
0>
0C
#322450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#322460000000
0!
0*
09
0>
0C
#322470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#322480000000
0!
0#
0*
0,
09
0>
0?
0C
#322490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#322500000000
0!
0*
09
0>
0C
#322510000000
1!
1*
19
1>
1C
#322520000000
0!
0*
09
0>
0C
#322530000000
1!
1*
19
1>
1C
#322540000000
0!
0*
09
0>
0C
#322550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#322560000000
0!
0*
09
0>
0C
#322570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#322580000000
0!
0*
09
0>
0C
#322590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#322600000000
0!
0*
09
0>
0C
#322610000000
1!
1*
b10 6
19
1>
1C
b10 G
#322620000000
0!
0*
09
0>
0C
#322630000000
1!
1*
b11 6
19
1>
1C
b11 G
#322640000000
0!
0*
09
0>
0C
#322650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#322660000000
0!
0*
09
0>
0C
#322670000000
1!
1*
b101 6
19
1>
1C
b101 G
#322680000000
0!
0*
09
0>
0C
#322690000000
1!
1*
b110 6
19
1>
1C
b110 G
#322700000000
0!
0*
09
0>
0C
#322710000000
1!
1*
b111 6
19
1>
1C
b111 G
#322720000000
0!
0*
09
0>
0C
#322730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#322740000000
0!
0*
09
0>
0C
#322750000000
1!
1*
b1 6
19
1>
1C
b1 G
#322760000000
0!
0*
09
0>
0C
#322770000000
1!
1*
b10 6
19
1>
1C
b10 G
#322780000000
0!
0*
09
0>
0C
#322790000000
1!
1*
b11 6
19
1>
1C
b11 G
#322800000000
0!
0*
09
0>
0C
#322810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#322820000000
0!
0*
09
0>
0C
#322830000000
1!
1*
b101 6
19
1>
1C
b101 G
#322840000000
0!
0*
09
0>
0C
#322850000000
1!
1*
b110 6
19
1>
1C
b110 G
#322860000000
0!
0*
09
0>
0C
#322870000000
1!
1*
b111 6
19
1>
1C
b111 G
#322880000000
0!
0*
09
0>
0C
#322890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#322900000000
0!
0*
09
0>
0C
#322910000000
1!
1*
b1 6
19
1>
1C
b1 G
#322920000000
0!
0*
09
0>
0C
#322930000000
1!
1*
b10 6
19
1>
1C
b10 G
#322940000000
0!
0*
09
0>
0C
#322950000000
1!
1*
b11 6
19
1>
1C
b11 G
#322960000000
0!
0*
09
0>
0C
#322970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#322980000000
0!
0*
09
0>
0C
#322990000000
1!
1*
b101 6
19
1>
1C
b101 G
#323000000000
0!
0*
09
0>
0C
#323010000000
1!
1*
b110 6
19
1>
1C
b110 G
#323020000000
0!
0*
09
0>
0C
#323030000000
1!
1*
b111 6
19
1>
1C
b111 G
#323040000000
0!
1"
0*
1+
09
1:
0>
0C
#323050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#323060000000
0!
0*
09
0>
0C
#323070000000
1!
1*
b1 6
19
1>
1C
b1 G
#323080000000
0!
0*
09
0>
0C
#323090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#323100000000
0!
0*
09
0>
0C
#323110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#323120000000
0!
0*
09
0>
0C
#323130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#323140000000
0!
0*
09
0>
0C
#323150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#323160000000
0!
0#
0*
0,
09
0>
0?
0C
#323170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#323180000000
0!
0*
09
0>
0C
#323190000000
1!
1*
19
1>
1C
#323200000000
0!
0*
09
0>
0C
#323210000000
1!
1*
19
1>
1C
#323220000000
0!
0*
09
0>
0C
#323230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#323240000000
0!
0*
09
0>
0C
#323250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#323260000000
0!
0*
09
0>
0C
#323270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#323280000000
0!
0*
09
0>
0C
#323290000000
1!
1*
b10 6
19
1>
1C
b10 G
#323300000000
0!
0*
09
0>
0C
#323310000000
1!
1*
b11 6
19
1>
1C
b11 G
#323320000000
0!
0*
09
0>
0C
#323330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#323340000000
0!
0*
09
0>
0C
#323350000000
1!
1*
b101 6
19
1>
1C
b101 G
#323360000000
0!
0*
09
0>
0C
#323370000000
1!
1*
b110 6
19
1>
1C
b110 G
#323380000000
0!
0*
09
0>
0C
#323390000000
1!
1*
b111 6
19
1>
1C
b111 G
#323400000000
0!
0*
09
0>
0C
#323410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#323420000000
0!
0*
09
0>
0C
#323430000000
1!
1*
b1 6
19
1>
1C
b1 G
#323440000000
0!
0*
09
0>
0C
#323450000000
1!
1*
b10 6
19
1>
1C
b10 G
#323460000000
0!
0*
09
0>
0C
#323470000000
1!
1*
b11 6
19
1>
1C
b11 G
#323480000000
0!
0*
09
0>
0C
#323490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#323500000000
0!
0*
09
0>
0C
#323510000000
1!
1*
b101 6
19
1>
1C
b101 G
#323520000000
0!
0*
09
0>
0C
#323530000000
1!
1*
b110 6
19
1>
1C
b110 G
#323540000000
0!
0*
09
0>
0C
#323550000000
1!
1*
b111 6
19
1>
1C
b111 G
#323560000000
0!
0*
09
0>
0C
#323570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#323580000000
0!
0*
09
0>
0C
#323590000000
1!
1*
b1 6
19
1>
1C
b1 G
#323600000000
0!
0*
09
0>
0C
#323610000000
1!
1*
b10 6
19
1>
1C
b10 G
#323620000000
0!
0*
09
0>
0C
#323630000000
1!
1*
b11 6
19
1>
1C
b11 G
#323640000000
0!
0*
09
0>
0C
#323650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#323660000000
0!
0*
09
0>
0C
#323670000000
1!
1*
b101 6
19
1>
1C
b101 G
#323680000000
0!
0*
09
0>
0C
#323690000000
1!
1*
b110 6
19
1>
1C
b110 G
#323700000000
0!
0*
09
0>
0C
#323710000000
1!
1*
b111 6
19
1>
1C
b111 G
#323720000000
0!
1"
0*
1+
09
1:
0>
0C
#323730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#323740000000
0!
0*
09
0>
0C
#323750000000
1!
1*
b1 6
19
1>
1C
b1 G
#323760000000
0!
0*
09
0>
0C
#323770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#323780000000
0!
0*
09
0>
0C
#323790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#323800000000
0!
0*
09
0>
0C
#323810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#323820000000
0!
0*
09
0>
0C
#323830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#323840000000
0!
0#
0*
0,
09
0>
0?
0C
#323850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#323860000000
0!
0*
09
0>
0C
#323870000000
1!
1*
19
1>
1C
#323880000000
0!
0*
09
0>
0C
#323890000000
1!
1*
19
1>
1C
#323900000000
0!
0*
09
0>
0C
#323910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#323920000000
0!
0*
09
0>
0C
#323930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#323940000000
0!
0*
09
0>
0C
#323950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#323960000000
0!
0*
09
0>
0C
#323970000000
1!
1*
b10 6
19
1>
1C
b10 G
#323980000000
0!
0*
09
0>
0C
#323990000000
1!
1*
b11 6
19
1>
1C
b11 G
#324000000000
0!
0*
09
0>
0C
#324010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#324020000000
0!
0*
09
0>
0C
#324030000000
1!
1*
b101 6
19
1>
1C
b101 G
#324040000000
0!
0*
09
0>
0C
#324050000000
1!
1*
b110 6
19
1>
1C
b110 G
#324060000000
0!
0*
09
0>
0C
#324070000000
1!
1*
b111 6
19
1>
1C
b111 G
#324080000000
0!
0*
09
0>
0C
#324090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#324100000000
0!
0*
09
0>
0C
#324110000000
1!
1*
b1 6
19
1>
1C
b1 G
#324120000000
0!
0*
09
0>
0C
#324130000000
1!
1*
b10 6
19
1>
1C
b10 G
#324140000000
0!
0*
09
0>
0C
#324150000000
1!
1*
b11 6
19
1>
1C
b11 G
#324160000000
0!
0*
09
0>
0C
#324170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#324180000000
0!
0*
09
0>
0C
#324190000000
1!
1*
b101 6
19
1>
1C
b101 G
#324200000000
0!
0*
09
0>
0C
#324210000000
1!
1*
b110 6
19
1>
1C
b110 G
#324220000000
0!
0*
09
0>
0C
#324230000000
1!
1*
b111 6
19
1>
1C
b111 G
#324240000000
0!
0*
09
0>
0C
#324250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#324260000000
0!
0*
09
0>
0C
#324270000000
1!
1*
b1 6
19
1>
1C
b1 G
#324280000000
0!
0*
09
0>
0C
#324290000000
1!
1*
b10 6
19
1>
1C
b10 G
#324300000000
0!
0*
09
0>
0C
#324310000000
1!
1*
b11 6
19
1>
1C
b11 G
#324320000000
0!
0*
09
0>
0C
#324330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#324340000000
0!
0*
09
0>
0C
#324350000000
1!
1*
b101 6
19
1>
1C
b101 G
#324360000000
0!
0*
09
0>
0C
#324370000000
1!
1*
b110 6
19
1>
1C
b110 G
#324380000000
0!
0*
09
0>
0C
#324390000000
1!
1*
b111 6
19
1>
1C
b111 G
#324400000000
0!
1"
0*
1+
09
1:
0>
0C
#324410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#324420000000
0!
0*
09
0>
0C
#324430000000
1!
1*
b1 6
19
1>
1C
b1 G
#324440000000
0!
0*
09
0>
0C
#324450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#324460000000
0!
0*
09
0>
0C
#324470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#324480000000
0!
0*
09
0>
0C
#324490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#324500000000
0!
0*
09
0>
0C
#324510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#324520000000
0!
0#
0*
0,
09
0>
0?
0C
#324530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#324540000000
0!
0*
09
0>
0C
#324550000000
1!
1*
19
1>
1C
#324560000000
0!
0*
09
0>
0C
#324570000000
1!
1*
19
1>
1C
#324580000000
0!
0*
09
0>
0C
#324590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#324600000000
0!
0*
09
0>
0C
#324610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#324620000000
0!
0*
09
0>
0C
#324630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#324640000000
0!
0*
09
0>
0C
#324650000000
1!
1*
b10 6
19
1>
1C
b10 G
#324660000000
0!
0*
09
0>
0C
#324670000000
1!
1*
b11 6
19
1>
1C
b11 G
#324680000000
0!
0*
09
0>
0C
#324690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#324700000000
0!
0*
09
0>
0C
#324710000000
1!
1*
b101 6
19
1>
1C
b101 G
#324720000000
0!
0*
09
0>
0C
#324730000000
1!
1*
b110 6
19
1>
1C
b110 G
#324740000000
0!
0*
09
0>
0C
#324750000000
1!
1*
b111 6
19
1>
1C
b111 G
#324760000000
0!
0*
09
0>
0C
#324770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#324780000000
0!
0*
09
0>
0C
#324790000000
1!
1*
b1 6
19
1>
1C
b1 G
#324800000000
0!
0*
09
0>
0C
#324810000000
1!
1*
b10 6
19
1>
1C
b10 G
#324820000000
0!
0*
09
0>
0C
#324830000000
1!
1*
b11 6
19
1>
1C
b11 G
#324840000000
0!
0*
09
0>
0C
#324850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#324860000000
0!
0*
09
0>
0C
#324870000000
1!
1*
b101 6
19
1>
1C
b101 G
#324880000000
0!
0*
09
0>
0C
#324890000000
1!
1*
b110 6
19
1>
1C
b110 G
#324900000000
0!
0*
09
0>
0C
#324910000000
1!
1*
b111 6
19
1>
1C
b111 G
#324920000000
0!
0*
09
0>
0C
#324930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#324940000000
0!
0*
09
0>
0C
#324950000000
1!
1*
b1 6
19
1>
1C
b1 G
#324960000000
0!
0*
09
0>
0C
#324970000000
1!
1*
b10 6
19
1>
1C
b10 G
#324980000000
0!
0*
09
0>
0C
#324990000000
1!
1*
b11 6
19
1>
1C
b11 G
#325000000000
0!
0*
09
0>
0C
#325010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#325020000000
0!
0*
09
0>
0C
#325030000000
1!
1*
b101 6
19
1>
1C
b101 G
#325040000000
0!
0*
09
0>
0C
#325050000000
1!
1*
b110 6
19
1>
1C
b110 G
#325060000000
0!
0*
09
0>
0C
#325070000000
1!
1*
b111 6
19
1>
1C
b111 G
#325080000000
0!
1"
0*
1+
09
1:
0>
0C
#325090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#325100000000
0!
0*
09
0>
0C
#325110000000
1!
1*
b1 6
19
1>
1C
b1 G
#325120000000
0!
0*
09
0>
0C
#325130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#325140000000
0!
0*
09
0>
0C
#325150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#325160000000
0!
0*
09
0>
0C
#325170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#325180000000
0!
0*
09
0>
0C
#325190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#325200000000
0!
0#
0*
0,
09
0>
0?
0C
#325210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#325220000000
0!
0*
09
0>
0C
#325230000000
1!
1*
19
1>
1C
#325240000000
0!
0*
09
0>
0C
#325250000000
1!
1*
19
1>
1C
#325260000000
0!
0*
09
0>
0C
#325270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#325280000000
0!
0*
09
0>
0C
#325290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#325300000000
0!
0*
09
0>
0C
#325310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#325320000000
0!
0*
09
0>
0C
#325330000000
1!
1*
b10 6
19
1>
1C
b10 G
#325340000000
0!
0*
09
0>
0C
#325350000000
1!
1*
b11 6
19
1>
1C
b11 G
#325360000000
0!
0*
09
0>
0C
#325370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#325380000000
0!
0*
09
0>
0C
#325390000000
1!
1*
b101 6
19
1>
1C
b101 G
#325400000000
0!
0*
09
0>
0C
#325410000000
1!
1*
b110 6
19
1>
1C
b110 G
#325420000000
0!
0*
09
0>
0C
#325430000000
1!
1*
b111 6
19
1>
1C
b111 G
#325440000000
0!
0*
09
0>
0C
#325450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#325460000000
0!
0*
09
0>
0C
#325470000000
1!
1*
b1 6
19
1>
1C
b1 G
#325480000000
0!
0*
09
0>
0C
#325490000000
1!
1*
b10 6
19
1>
1C
b10 G
#325500000000
0!
0*
09
0>
0C
#325510000000
1!
1*
b11 6
19
1>
1C
b11 G
#325520000000
0!
0*
09
0>
0C
#325530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#325540000000
0!
0*
09
0>
0C
#325550000000
1!
1*
b101 6
19
1>
1C
b101 G
#325560000000
0!
0*
09
0>
0C
#325570000000
1!
1*
b110 6
19
1>
1C
b110 G
#325580000000
0!
0*
09
0>
0C
#325590000000
1!
1*
b111 6
19
1>
1C
b111 G
#325600000000
0!
0*
09
0>
0C
#325610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#325620000000
0!
0*
09
0>
0C
#325630000000
1!
1*
b1 6
19
1>
1C
b1 G
#325640000000
0!
0*
09
0>
0C
#325650000000
1!
1*
b10 6
19
1>
1C
b10 G
#325660000000
0!
0*
09
0>
0C
#325670000000
1!
1*
b11 6
19
1>
1C
b11 G
#325680000000
0!
0*
09
0>
0C
#325690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#325700000000
0!
0*
09
0>
0C
#325710000000
1!
1*
b101 6
19
1>
1C
b101 G
#325720000000
0!
0*
09
0>
0C
#325730000000
1!
1*
b110 6
19
1>
1C
b110 G
#325740000000
0!
0*
09
0>
0C
#325750000000
1!
1*
b111 6
19
1>
1C
b111 G
#325760000000
0!
1"
0*
1+
09
1:
0>
0C
#325770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#325780000000
0!
0*
09
0>
0C
#325790000000
1!
1*
b1 6
19
1>
1C
b1 G
#325800000000
0!
0*
09
0>
0C
#325810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#325820000000
0!
0*
09
0>
0C
#325830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#325840000000
0!
0*
09
0>
0C
#325850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#325860000000
0!
0*
09
0>
0C
#325870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#325880000000
0!
0#
0*
0,
09
0>
0?
0C
#325890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#325900000000
0!
0*
09
0>
0C
#325910000000
1!
1*
19
1>
1C
#325920000000
0!
0*
09
0>
0C
#325930000000
1!
1*
19
1>
1C
#325940000000
0!
0*
09
0>
0C
#325950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#325960000000
0!
0*
09
0>
0C
#325970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#325980000000
0!
0*
09
0>
0C
#325990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#326000000000
0!
0*
09
0>
0C
#326010000000
1!
1*
b10 6
19
1>
1C
b10 G
#326020000000
0!
0*
09
0>
0C
#326030000000
1!
1*
b11 6
19
1>
1C
b11 G
#326040000000
0!
0*
09
0>
0C
#326050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#326060000000
0!
0*
09
0>
0C
#326070000000
1!
1*
b101 6
19
1>
1C
b101 G
#326080000000
0!
0*
09
0>
0C
#326090000000
1!
1*
b110 6
19
1>
1C
b110 G
#326100000000
0!
0*
09
0>
0C
#326110000000
1!
1*
b111 6
19
1>
1C
b111 G
#326120000000
0!
0*
09
0>
0C
#326130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#326140000000
0!
0*
09
0>
0C
#326150000000
1!
1*
b1 6
19
1>
1C
b1 G
#326160000000
0!
0*
09
0>
0C
#326170000000
1!
1*
b10 6
19
1>
1C
b10 G
#326180000000
0!
0*
09
0>
0C
#326190000000
1!
1*
b11 6
19
1>
1C
b11 G
#326200000000
0!
0*
09
0>
0C
#326210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#326220000000
0!
0*
09
0>
0C
#326230000000
1!
1*
b101 6
19
1>
1C
b101 G
#326240000000
0!
0*
09
0>
0C
#326250000000
1!
1*
b110 6
19
1>
1C
b110 G
#326260000000
0!
0*
09
0>
0C
#326270000000
1!
1*
b111 6
19
1>
1C
b111 G
#326280000000
0!
0*
09
0>
0C
#326290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#326300000000
0!
0*
09
0>
0C
#326310000000
1!
1*
b1 6
19
1>
1C
b1 G
#326320000000
0!
0*
09
0>
0C
#326330000000
1!
1*
b10 6
19
1>
1C
b10 G
#326340000000
0!
0*
09
0>
0C
#326350000000
1!
1*
b11 6
19
1>
1C
b11 G
#326360000000
0!
0*
09
0>
0C
#326370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#326380000000
0!
0*
09
0>
0C
#326390000000
1!
1*
b101 6
19
1>
1C
b101 G
#326400000000
0!
0*
09
0>
0C
#326410000000
1!
1*
b110 6
19
1>
1C
b110 G
#326420000000
0!
0*
09
0>
0C
#326430000000
1!
1*
b111 6
19
1>
1C
b111 G
#326440000000
0!
1"
0*
1+
09
1:
0>
0C
#326450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#326460000000
0!
0*
09
0>
0C
#326470000000
1!
1*
b1 6
19
1>
1C
b1 G
#326480000000
0!
0*
09
0>
0C
#326490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#326500000000
0!
0*
09
0>
0C
#326510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#326520000000
0!
0*
09
0>
0C
#326530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#326540000000
0!
0*
09
0>
0C
#326550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#326560000000
0!
0#
0*
0,
09
0>
0?
0C
#326570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#326580000000
0!
0*
09
0>
0C
#326590000000
1!
1*
19
1>
1C
#326600000000
0!
0*
09
0>
0C
#326610000000
1!
1*
19
1>
1C
#326620000000
0!
0*
09
0>
0C
#326630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#326640000000
0!
0*
09
0>
0C
#326650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#326660000000
0!
0*
09
0>
0C
#326670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#326680000000
0!
0*
09
0>
0C
#326690000000
1!
1*
b10 6
19
1>
1C
b10 G
#326700000000
0!
0*
09
0>
0C
#326710000000
1!
1*
b11 6
19
1>
1C
b11 G
#326720000000
0!
0*
09
0>
0C
#326730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#326740000000
0!
0*
09
0>
0C
#326750000000
1!
1*
b101 6
19
1>
1C
b101 G
#326760000000
0!
0*
09
0>
0C
#326770000000
1!
1*
b110 6
19
1>
1C
b110 G
#326780000000
0!
0*
09
0>
0C
#326790000000
1!
1*
b111 6
19
1>
1C
b111 G
#326800000000
0!
0*
09
0>
0C
#326810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#326820000000
0!
0*
09
0>
0C
#326830000000
1!
1*
b1 6
19
1>
1C
b1 G
#326840000000
0!
0*
09
0>
0C
#326850000000
1!
1*
b10 6
19
1>
1C
b10 G
#326860000000
0!
0*
09
0>
0C
#326870000000
1!
1*
b11 6
19
1>
1C
b11 G
#326880000000
0!
0*
09
0>
0C
#326890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#326900000000
0!
0*
09
0>
0C
#326910000000
1!
1*
b101 6
19
1>
1C
b101 G
#326920000000
0!
0*
09
0>
0C
#326930000000
1!
1*
b110 6
19
1>
1C
b110 G
#326940000000
0!
0*
09
0>
0C
#326950000000
1!
1*
b111 6
19
1>
1C
b111 G
#326960000000
0!
0*
09
0>
0C
#326970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#326980000000
0!
0*
09
0>
0C
#326990000000
1!
1*
b1 6
19
1>
1C
b1 G
#327000000000
0!
0*
09
0>
0C
#327010000000
1!
1*
b10 6
19
1>
1C
b10 G
#327020000000
0!
0*
09
0>
0C
#327030000000
1!
1*
b11 6
19
1>
1C
b11 G
#327040000000
0!
0*
09
0>
0C
#327050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#327060000000
0!
0*
09
0>
0C
#327070000000
1!
1*
b101 6
19
1>
1C
b101 G
#327080000000
0!
0*
09
0>
0C
#327090000000
1!
1*
b110 6
19
1>
1C
b110 G
#327100000000
0!
0*
09
0>
0C
#327110000000
1!
1*
b111 6
19
1>
1C
b111 G
#327120000000
0!
1"
0*
1+
09
1:
0>
0C
#327130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#327140000000
0!
0*
09
0>
0C
#327150000000
1!
1*
b1 6
19
1>
1C
b1 G
#327160000000
0!
0*
09
0>
0C
#327170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#327180000000
0!
0*
09
0>
0C
#327190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#327200000000
0!
0*
09
0>
0C
#327210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#327220000000
0!
0*
09
0>
0C
#327230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#327240000000
0!
0#
0*
0,
09
0>
0?
0C
#327250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#327260000000
0!
0*
09
0>
0C
#327270000000
1!
1*
19
1>
1C
#327280000000
0!
0*
09
0>
0C
#327290000000
1!
1*
19
1>
1C
#327300000000
0!
0*
09
0>
0C
#327310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#327320000000
0!
0*
09
0>
0C
#327330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#327340000000
0!
0*
09
0>
0C
#327350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#327360000000
0!
0*
09
0>
0C
#327370000000
1!
1*
b10 6
19
1>
1C
b10 G
#327380000000
0!
0*
09
0>
0C
#327390000000
1!
1*
b11 6
19
1>
1C
b11 G
#327400000000
0!
0*
09
0>
0C
#327410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#327420000000
0!
0*
09
0>
0C
#327430000000
1!
1*
b101 6
19
1>
1C
b101 G
#327440000000
0!
0*
09
0>
0C
#327450000000
1!
1*
b110 6
19
1>
1C
b110 G
#327460000000
0!
0*
09
0>
0C
#327470000000
1!
1*
b111 6
19
1>
1C
b111 G
#327480000000
0!
0*
09
0>
0C
#327490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#327500000000
0!
0*
09
0>
0C
#327510000000
1!
1*
b1 6
19
1>
1C
b1 G
#327520000000
0!
0*
09
0>
0C
#327530000000
1!
1*
b10 6
19
1>
1C
b10 G
#327540000000
0!
0*
09
0>
0C
#327550000000
1!
1*
b11 6
19
1>
1C
b11 G
#327560000000
0!
0*
09
0>
0C
#327570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#327580000000
0!
0*
09
0>
0C
#327590000000
1!
1*
b101 6
19
1>
1C
b101 G
#327600000000
0!
0*
09
0>
0C
#327610000000
1!
1*
b110 6
19
1>
1C
b110 G
#327620000000
0!
0*
09
0>
0C
#327630000000
1!
1*
b111 6
19
1>
1C
b111 G
#327640000000
0!
0*
09
0>
0C
#327650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#327660000000
0!
0*
09
0>
0C
#327670000000
1!
1*
b1 6
19
1>
1C
b1 G
#327680000000
0!
0*
09
0>
0C
#327690000000
1!
1*
b10 6
19
1>
1C
b10 G
#327700000000
0!
0*
09
0>
0C
#327710000000
1!
1*
b11 6
19
1>
1C
b11 G
#327720000000
0!
0*
09
0>
0C
#327730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#327740000000
0!
0*
09
0>
0C
#327750000000
1!
1*
b101 6
19
1>
1C
b101 G
#327760000000
0!
0*
09
0>
0C
#327770000000
1!
1*
b110 6
19
1>
1C
b110 G
#327780000000
0!
0*
09
0>
0C
#327790000000
1!
1*
b111 6
19
1>
1C
b111 G
#327800000000
0!
1"
0*
1+
09
1:
0>
0C
#327810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#327820000000
0!
0*
09
0>
0C
#327830000000
1!
1*
b1 6
19
1>
1C
b1 G
#327840000000
0!
0*
09
0>
0C
#327850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#327860000000
0!
0*
09
0>
0C
#327870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#327880000000
0!
0*
09
0>
0C
#327890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#327900000000
0!
0*
09
0>
0C
#327910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#327920000000
0!
0#
0*
0,
09
0>
0?
0C
#327930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#327940000000
0!
0*
09
0>
0C
#327950000000
1!
1*
19
1>
1C
#327960000000
0!
0*
09
0>
0C
#327970000000
1!
1*
19
1>
1C
#327980000000
0!
0*
09
0>
0C
#327990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#328000000000
0!
0*
09
0>
0C
#328010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#328020000000
0!
0*
09
0>
0C
#328030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#328040000000
0!
0*
09
0>
0C
#328050000000
1!
1*
b10 6
19
1>
1C
b10 G
#328060000000
0!
0*
09
0>
0C
#328070000000
1!
1*
b11 6
19
1>
1C
b11 G
#328080000000
0!
0*
09
0>
0C
#328090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#328100000000
0!
0*
09
0>
0C
#328110000000
1!
1*
b101 6
19
1>
1C
b101 G
#328120000000
0!
0*
09
0>
0C
#328130000000
1!
1*
b110 6
19
1>
1C
b110 G
#328140000000
0!
0*
09
0>
0C
#328150000000
1!
1*
b111 6
19
1>
1C
b111 G
#328160000000
0!
0*
09
0>
0C
#328170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#328180000000
0!
0*
09
0>
0C
#328190000000
1!
1*
b1 6
19
1>
1C
b1 G
#328200000000
0!
0*
09
0>
0C
#328210000000
1!
1*
b10 6
19
1>
1C
b10 G
#328220000000
0!
0*
09
0>
0C
#328230000000
1!
1*
b11 6
19
1>
1C
b11 G
#328240000000
0!
0*
09
0>
0C
#328250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#328260000000
0!
0*
09
0>
0C
#328270000000
1!
1*
b101 6
19
1>
1C
b101 G
#328280000000
0!
0*
09
0>
0C
#328290000000
1!
1*
b110 6
19
1>
1C
b110 G
#328300000000
0!
0*
09
0>
0C
#328310000000
1!
1*
b111 6
19
1>
1C
b111 G
#328320000000
0!
0*
09
0>
0C
#328330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#328340000000
0!
0*
09
0>
0C
#328350000000
1!
1*
b1 6
19
1>
1C
b1 G
#328360000000
0!
0*
09
0>
0C
#328370000000
1!
1*
b10 6
19
1>
1C
b10 G
#328380000000
0!
0*
09
0>
0C
#328390000000
1!
1*
b11 6
19
1>
1C
b11 G
#328400000000
0!
0*
09
0>
0C
#328410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#328420000000
0!
0*
09
0>
0C
#328430000000
1!
1*
b101 6
19
1>
1C
b101 G
#328440000000
0!
0*
09
0>
0C
#328450000000
1!
1*
b110 6
19
1>
1C
b110 G
#328460000000
0!
0*
09
0>
0C
#328470000000
1!
1*
b111 6
19
1>
1C
b111 G
#328480000000
0!
1"
0*
1+
09
1:
0>
0C
#328490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#328500000000
0!
0*
09
0>
0C
#328510000000
1!
1*
b1 6
19
1>
1C
b1 G
#328520000000
0!
0*
09
0>
0C
#328530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#328540000000
0!
0*
09
0>
0C
#328550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#328560000000
0!
0*
09
0>
0C
#328570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#328580000000
0!
0*
09
0>
0C
#328590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#328600000000
0!
0#
0*
0,
09
0>
0?
0C
#328610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#328620000000
0!
0*
09
0>
0C
#328630000000
1!
1*
19
1>
1C
#328640000000
0!
0*
09
0>
0C
#328650000000
1!
1*
19
1>
1C
#328660000000
0!
0*
09
0>
0C
#328670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#328680000000
0!
0*
09
0>
0C
#328690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#328700000000
0!
0*
09
0>
0C
#328710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#328720000000
0!
0*
09
0>
0C
#328730000000
1!
1*
b10 6
19
1>
1C
b10 G
#328740000000
0!
0*
09
0>
0C
#328750000000
1!
1*
b11 6
19
1>
1C
b11 G
#328760000000
0!
0*
09
0>
0C
#328770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#328780000000
0!
0*
09
0>
0C
#328790000000
1!
1*
b101 6
19
1>
1C
b101 G
#328800000000
0!
0*
09
0>
0C
#328810000000
1!
1*
b110 6
19
1>
1C
b110 G
#328820000000
0!
0*
09
0>
0C
#328830000000
1!
1*
b111 6
19
1>
1C
b111 G
#328840000000
0!
0*
09
0>
0C
#328850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#328860000000
0!
0*
09
0>
0C
#328870000000
1!
1*
b1 6
19
1>
1C
b1 G
#328880000000
0!
0*
09
0>
0C
#328890000000
1!
1*
b10 6
19
1>
1C
b10 G
#328900000000
0!
0*
09
0>
0C
#328910000000
1!
1*
b11 6
19
1>
1C
b11 G
#328920000000
0!
0*
09
0>
0C
#328930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#328940000000
0!
0*
09
0>
0C
#328950000000
1!
1*
b101 6
19
1>
1C
b101 G
#328960000000
0!
0*
09
0>
0C
#328970000000
1!
1*
b110 6
19
1>
1C
b110 G
#328980000000
0!
0*
09
0>
0C
#328990000000
1!
1*
b111 6
19
1>
1C
b111 G
#329000000000
0!
0*
09
0>
0C
#329010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#329020000000
0!
0*
09
0>
0C
#329030000000
1!
1*
b1 6
19
1>
1C
b1 G
#329040000000
0!
0*
09
0>
0C
#329050000000
1!
1*
b10 6
19
1>
1C
b10 G
#329060000000
0!
0*
09
0>
0C
#329070000000
1!
1*
b11 6
19
1>
1C
b11 G
#329080000000
0!
0*
09
0>
0C
#329090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#329100000000
0!
0*
09
0>
0C
#329110000000
1!
1*
b101 6
19
1>
1C
b101 G
#329120000000
0!
0*
09
0>
0C
#329130000000
1!
1*
b110 6
19
1>
1C
b110 G
#329140000000
0!
0*
09
0>
0C
#329150000000
1!
1*
b111 6
19
1>
1C
b111 G
#329160000000
0!
1"
0*
1+
09
1:
0>
0C
#329170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#329180000000
0!
0*
09
0>
0C
#329190000000
1!
1*
b1 6
19
1>
1C
b1 G
#329200000000
0!
0*
09
0>
0C
#329210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#329220000000
0!
0*
09
0>
0C
#329230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#329240000000
0!
0*
09
0>
0C
#329250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#329260000000
0!
0*
09
0>
0C
#329270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#329280000000
0!
0#
0*
0,
09
0>
0?
0C
#329290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#329300000000
0!
0*
09
0>
0C
#329310000000
1!
1*
19
1>
1C
#329320000000
0!
0*
09
0>
0C
#329330000000
1!
1*
19
1>
1C
#329340000000
0!
0*
09
0>
0C
#329350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#329360000000
0!
0*
09
0>
0C
#329370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#329380000000
0!
0*
09
0>
0C
#329390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#329400000000
0!
0*
09
0>
0C
#329410000000
1!
1*
b10 6
19
1>
1C
b10 G
#329420000000
0!
0*
09
0>
0C
#329430000000
1!
1*
b11 6
19
1>
1C
b11 G
#329440000000
0!
0*
09
0>
0C
#329450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#329460000000
0!
0*
09
0>
0C
#329470000000
1!
1*
b101 6
19
1>
1C
b101 G
#329480000000
0!
0*
09
0>
0C
#329490000000
1!
1*
b110 6
19
1>
1C
b110 G
#329500000000
0!
0*
09
0>
0C
#329510000000
1!
1*
b111 6
19
1>
1C
b111 G
#329520000000
0!
0*
09
0>
0C
#329530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#329540000000
0!
0*
09
0>
0C
#329550000000
1!
1*
b1 6
19
1>
1C
b1 G
#329560000000
0!
0*
09
0>
0C
#329570000000
1!
1*
b10 6
19
1>
1C
b10 G
#329580000000
0!
0*
09
0>
0C
#329590000000
1!
1*
b11 6
19
1>
1C
b11 G
#329600000000
0!
0*
09
0>
0C
#329610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#329620000000
0!
0*
09
0>
0C
#329630000000
1!
1*
b101 6
19
1>
1C
b101 G
#329640000000
0!
0*
09
0>
0C
#329650000000
1!
1*
b110 6
19
1>
1C
b110 G
#329660000000
0!
0*
09
0>
0C
#329670000000
1!
1*
b111 6
19
1>
1C
b111 G
#329680000000
0!
0*
09
0>
0C
#329690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#329700000000
0!
0*
09
0>
0C
#329710000000
1!
1*
b1 6
19
1>
1C
b1 G
#329720000000
0!
0*
09
0>
0C
#329730000000
1!
1*
b10 6
19
1>
1C
b10 G
#329740000000
0!
0*
09
0>
0C
#329750000000
1!
1*
b11 6
19
1>
1C
b11 G
#329760000000
0!
0*
09
0>
0C
#329770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#329780000000
0!
0*
09
0>
0C
#329790000000
1!
1*
b101 6
19
1>
1C
b101 G
#329800000000
0!
0*
09
0>
0C
#329810000000
1!
1*
b110 6
19
1>
1C
b110 G
#329820000000
0!
0*
09
0>
0C
#329830000000
1!
1*
b111 6
19
1>
1C
b111 G
#329840000000
0!
1"
0*
1+
09
1:
0>
0C
#329850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#329860000000
0!
0*
09
0>
0C
#329870000000
1!
1*
b1 6
19
1>
1C
b1 G
#329880000000
0!
0*
09
0>
0C
#329890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#329900000000
0!
0*
09
0>
0C
#329910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#329920000000
0!
0*
09
0>
0C
#329930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#329940000000
0!
0*
09
0>
0C
#329950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#329960000000
0!
0#
0*
0,
09
0>
0?
0C
#329970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#329980000000
0!
0*
09
0>
0C
#329990000000
1!
1*
19
1>
1C
#330000000000
0!
0*
09
0>
0C
#330010000000
1!
1*
19
1>
1C
#330020000000
0!
0*
09
0>
0C
#330030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#330040000000
0!
0*
09
0>
0C
#330050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#330060000000
0!
0*
09
0>
0C
#330070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#330080000000
0!
0*
09
0>
0C
#330090000000
1!
1*
b10 6
19
1>
1C
b10 G
#330100000000
0!
0*
09
0>
0C
#330110000000
1!
1*
b11 6
19
1>
1C
b11 G
#330120000000
0!
0*
09
0>
0C
#330130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#330140000000
0!
0*
09
0>
0C
#330150000000
1!
1*
b101 6
19
1>
1C
b101 G
#330160000000
0!
0*
09
0>
0C
#330170000000
1!
1*
b110 6
19
1>
1C
b110 G
#330180000000
0!
0*
09
0>
0C
#330190000000
1!
1*
b111 6
19
1>
1C
b111 G
#330200000000
0!
0*
09
0>
0C
#330210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#330220000000
0!
0*
09
0>
0C
#330230000000
1!
1*
b1 6
19
1>
1C
b1 G
#330240000000
0!
0*
09
0>
0C
#330250000000
1!
1*
b10 6
19
1>
1C
b10 G
#330260000000
0!
0*
09
0>
0C
#330270000000
1!
1*
b11 6
19
1>
1C
b11 G
#330280000000
0!
0*
09
0>
0C
#330290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#330300000000
0!
0*
09
0>
0C
#330310000000
1!
1*
b101 6
19
1>
1C
b101 G
#330320000000
0!
0*
09
0>
0C
#330330000000
1!
1*
b110 6
19
1>
1C
b110 G
#330340000000
0!
0*
09
0>
0C
#330350000000
1!
1*
b111 6
19
1>
1C
b111 G
#330360000000
0!
0*
09
0>
0C
#330370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#330380000000
0!
0*
09
0>
0C
#330390000000
1!
1*
b1 6
19
1>
1C
b1 G
#330400000000
0!
0*
09
0>
0C
#330410000000
1!
1*
b10 6
19
1>
1C
b10 G
#330420000000
0!
0*
09
0>
0C
#330430000000
1!
1*
b11 6
19
1>
1C
b11 G
#330440000000
0!
0*
09
0>
0C
#330450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#330460000000
0!
0*
09
0>
0C
#330470000000
1!
1*
b101 6
19
1>
1C
b101 G
#330480000000
0!
0*
09
0>
0C
#330490000000
1!
1*
b110 6
19
1>
1C
b110 G
#330500000000
0!
0*
09
0>
0C
#330510000000
1!
1*
b111 6
19
1>
1C
b111 G
#330520000000
0!
1"
0*
1+
09
1:
0>
0C
#330530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#330540000000
0!
0*
09
0>
0C
#330550000000
1!
1*
b1 6
19
1>
1C
b1 G
#330560000000
0!
0*
09
0>
0C
#330570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#330580000000
0!
0*
09
0>
0C
#330590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#330600000000
0!
0*
09
0>
0C
#330610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#330620000000
0!
0*
09
0>
0C
#330630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#330640000000
0!
0#
0*
0,
09
0>
0?
0C
#330650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#330660000000
0!
0*
09
0>
0C
#330670000000
1!
1*
19
1>
1C
#330680000000
0!
0*
09
0>
0C
#330690000000
1!
1*
19
1>
1C
#330700000000
0!
0*
09
0>
0C
#330710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#330720000000
0!
0*
09
0>
0C
#330730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#330740000000
0!
0*
09
0>
0C
#330750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#330760000000
0!
0*
09
0>
0C
#330770000000
1!
1*
b10 6
19
1>
1C
b10 G
#330780000000
0!
0*
09
0>
0C
#330790000000
1!
1*
b11 6
19
1>
1C
b11 G
#330800000000
0!
0*
09
0>
0C
#330810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#330820000000
0!
0*
09
0>
0C
#330830000000
1!
1*
b101 6
19
1>
1C
b101 G
#330840000000
0!
0*
09
0>
0C
#330850000000
1!
1*
b110 6
19
1>
1C
b110 G
#330860000000
0!
0*
09
0>
0C
#330870000000
1!
1*
b111 6
19
1>
1C
b111 G
#330880000000
0!
0*
09
0>
0C
#330890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#330900000000
0!
0*
09
0>
0C
#330910000000
1!
1*
b1 6
19
1>
1C
b1 G
#330920000000
0!
0*
09
0>
0C
#330930000000
1!
1*
b10 6
19
1>
1C
b10 G
#330940000000
0!
0*
09
0>
0C
#330950000000
1!
1*
b11 6
19
1>
1C
b11 G
#330960000000
0!
0*
09
0>
0C
#330970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#330980000000
0!
0*
09
0>
0C
#330990000000
1!
1*
b101 6
19
1>
1C
b101 G
#331000000000
0!
0*
09
0>
0C
#331010000000
1!
1*
b110 6
19
1>
1C
b110 G
#331020000000
0!
0*
09
0>
0C
#331030000000
1!
1*
b111 6
19
1>
1C
b111 G
#331040000000
0!
0*
09
0>
0C
#331050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#331060000000
0!
0*
09
0>
0C
#331070000000
1!
1*
b1 6
19
1>
1C
b1 G
#331080000000
0!
0*
09
0>
0C
#331090000000
1!
1*
b10 6
19
1>
1C
b10 G
#331100000000
0!
0*
09
0>
0C
#331110000000
1!
1*
b11 6
19
1>
1C
b11 G
#331120000000
0!
0*
09
0>
0C
#331130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#331140000000
0!
0*
09
0>
0C
#331150000000
1!
1*
b101 6
19
1>
1C
b101 G
#331160000000
0!
0*
09
0>
0C
#331170000000
1!
1*
b110 6
19
1>
1C
b110 G
#331180000000
0!
0*
09
0>
0C
#331190000000
1!
1*
b111 6
19
1>
1C
b111 G
#331200000000
0!
1"
0*
1+
09
1:
0>
0C
#331210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#331220000000
0!
0*
09
0>
0C
#331230000000
1!
1*
b1 6
19
1>
1C
b1 G
#331240000000
0!
0*
09
0>
0C
#331250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#331260000000
0!
0*
09
0>
0C
#331270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#331280000000
0!
0*
09
0>
0C
#331290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#331300000000
0!
0*
09
0>
0C
#331310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#331320000000
0!
0#
0*
0,
09
0>
0?
0C
#331330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#331340000000
0!
0*
09
0>
0C
#331350000000
1!
1*
19
1>
1C
#331360000000
0!
0*
09
0>
0C
#331370000000
1!
1*
19
1>
1C
#331380000000
0!
0*
09
0>
0C
#331390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#331400000000
0!
0*
09
0>
0C
#331410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#331420000000
0!
0*
09
0>
0C
#331430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#331440000000
0!
0*
09
0>
0C
#331450000000
1!
1*
b10 6
19
1>
1C
b10 G
#331460000000
0!
0*
09
0>
0C
#331470000000
1!
1*
b11 6
19
1>
1C
b11 G
#331480000000
0!
0*
09
0>
0C
#331490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#331500000000
0!
0*
09
0>
0C
#331510000000
1!
1*
b101 6
19
1>
1C
b101 G
#331520000000
0!
0*
09
0>
0C
#331530000000
1!
1*
b110 6
19
1>
1C
b110 G
#331540000000
0!
0*
09
0>
0C
#331550000000
1!
1*
b111 6
19
1>
1C
b111 G
#331560000000
0!
0*
09
0>
0C
#331570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#331580000000
0!
0*
09
0>
0C
#331590000000
1!
1*
b1 6
19
1>
1C
b1 G
#331600000000
0!
0*
09
0>
0C
#331610000000
1!
1*
b10 6
19
1>
1C
b10 G
#331620000000
0!
0*
09
0>
0C
#331630000000
1!
1*
b11 6
19
1>
1C
b11 G
#331640000000
0!
0*
09
0>
0C
#331650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#331660000000
0!
0*
09
0>
0C
#331670000000
1!
1*
b101 6
19
1>
1C
b101 G
#331680000000
0!
0*
09
0>
0C
#331690000000
1!
1*
b110 6
19
1>
1C
b110 G
#331700000000
0!
0*
09
0>
0C
#331710000000
1!
1*
b111 6
19
1>
1C
b111 G
#331720000000
0!
0*
09
0>
0C
#331730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#331740000000
0!
0*
09
0>
0C
#331750000000
1!
1*
b1 6
19
1>
1C
b1 G
#331760000000
0!
0*
09
0>
0C
#331770000000
1!
1*
b10 6
19
1>
1C
b10 G
#331780000000
0!
0*
09
0>
0C
#331790000000
1!
1*
b11 6
19
1>
1C
b11 G
#331800000000
0!
0*
09
0>
0C
#331810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#331820000000
0!
0*
09
0>
0C
#331830000000
1!
1*
b101 6
19
1>
1C
b101 G
#331840000000
0!
0*
09
0>
0C
#331850000000
1!
1*
b110 6
19
1>
1C
b110 G
#331860000000
0!
0*
09
0>
0C
#331870000000
1!
1*
b111 6
19
1>
1C
b111 G
#331880000000
0!
1"
0*
1+
09
1:
0>
0C
#331890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#331900000000
0!
0*
09
0>
0C
#331910000000
1!
1*
b1 6
19
1>
1C
b1 G
#331920000000
0!
0*
09
0>
0C
#331930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#331940000000
0!
0*
09
0>
0C
#331950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#331960000000
0!
0*
09
0>
0C
#331970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#331980000000
0!
0*
09
0>
0C
#331990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#332000000000
0!
0#
0*
0,
09
0>
0?
0C
#332010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#332020000000
0!
0*
09
0>
0C
#332030000000
1!
1*
19
1>
1C
#332040000000
0!
0*
09
0>
0C
#332050000000
1!
1*
19
1>
1C
#332060000000
0!
0*
09
0>
0C
#332070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#332080000000
0!
0*
09
0>
0C
#332090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#332100000000
0!
0*
09
0>
0C
#332110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#332120000000
0!
0*
09
0>
0C
#332130000000
1!
1*
b10 6
19
1>
1C
b10 G
#332140000000
0!
0*
09
0>
0C
#332150000000
1!
1*
b11 6
19
1>
1C
b11 G
#332160000000
0!
0*
09
0>
0C
#332170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#332180000000
0!
0*
09
0>
0C
#332190000000
1!
1*
b101 6
19
1>
1C
b101 G
#332200000000
0!
0*
09
0>
0C
#332210000000
1!
1*
b110 6
19
1>
1C
b110 G
#332220000000
0!
0*
09
0>
0C
#332230000000
1!
1*
b111 6
19
1>
1C
b111 G
#332240000000
0!
0*
09
0>
0C
#332250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#332260000000
0!
0*
09
0>
0C
#332270000000
1!
1*
b1 6
19
1>
1C
b1 G
#332280000000
0!
0*
09
0>
0C
#332290000000
1!
1*
b10 6
19
1>
1C
b10 G
#332300000000
0!
0*
09
0>
0C
#332310000000
1!
1*
b11 6
19
1>
1C
b11 G
#332320000000
0!
0*
09
0>
0C
#332330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#332340000000
0!
0*
09
0>
0C
#332350000000
1!
1*
b101 6
19
1>
1C
b101 G
#332360000000
0!
0*
09
0>
0C
#332370000000
1!
1*
b110 6
19
1>
1C
b110 G
#332380000000
0!
0*
09
0>
0C
#332390000000
1!
1*
b111 6
19
1>
1C
b111 G
#332400000000
0!
0*
09
0>
0C
#332410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#332420000000
0!
0*
09
0>
0C
#332430000000
1!
1*
b1 6
19
1>
1C
b1 G
#332440000000
0!
0*
09
0>
0C
#332450000000
1!
1*
b10 6
19
1>
1C
b10 G
#332460000000
0!
0*
09
0>
0C
#332470000000
1!
1*
b11 6
19
1>
1C
b11 G
#332480000000
0!
0*
09
0>
0C
#332490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#332500000000
0!
0*
09
0>
0C
#332510000000
1!
1*
b101 6
19
1>
1C
b101 G
#332520000000
0!
0*
09
0>
0C
#332530000000
1!
1*
b110 6
19
1>
1C
b110 G
#332540000000
0!
0*
09
0>
0C
#332550000000
1!
1*
b111 6
19
1>
1C
b111 G
#332560000000
0!
1"
0*
1+
09
1:
0>
0C
#332570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#332580000000
0!
0*
09
0>
0C
#332590000000
1!
1*
b1 6
19
1>
1C
b1 G
#332600000000
0!
0*
09
0>
0C
#332610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#332620000000
0!
0*
09
0>
0C
#332630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#332640000000
0!
0*
09
0>
0C
#332650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#332660000000
0!
0*
09
0>
0C
#332670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#332680000000
0!
0#
0*
0,
09
0>
0?
0C
#332690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#332700000000
0!
0*
09
0>
0C
#332710000000
1!
1*
19
1>
1C
#332720000000
0!
0*
09
0>
0C
#332730000000
1!
1*
19
1>
1C
#332740000000
0!
0*
09
0>
0C
#332750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#332760000000
0!
0*
09
0>
0C
#332770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#332780000000
0!
0*
09
0>
0C
#332790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#332800000000
0!
0*
09
0>
0C
#332810000000
1!
1*
b10 6
19
1>
1C
b10 G
#332820000000
0!
0*
09
0>
0C
#332830000000
1!
1*
b11 6
19
1>
1C
b11 G
#332840000000
0!
0*
09
0>
0C
#332850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#332860000000
0!
0*
09
0>
0C
#332870000000
1!
1*
b101 6
19
1>
1C
b101 G
#332880000000
0!
0*
09
0>
0C
#332890000000
1!
1*
b110 6
19
1>
1C
b110 G
#332900000000
0!
0*
09
0>
0C
#332910000000
1!
1*
b111 6
19
1>
1C
b111 G
#332920000000
0!
0*
09
0>
0C
#332930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#332940000000
0!
0*
09
0>
0C
#332950000000
1!
1*
b1 6
19
1>
1C
b1 G
#332960000000
0!
0*
09
0>
0C
#332970000000
1!
1*
b10 6
19
1>
1C
b10 G
#332980000000
0!
0*
09
0>
0C
#332990000000
1!
1*
b11 6
19
1>
1C
b11 G
#333000000000
0!
0*
09
0>
0C
#333010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#333020000000
0!
0*
09
0>
0C
#333030000000
1!
1*
b101 6
19
1>
1C
b101 G
#333040000000
0!
0*
09
0>
0C
#333050000000
1!
1*
b110 6
19
1>
1C
b110 G
#333060000000
0!
0*
09
0>
0C
#333070000000
1!
1*
b111 6
19
1>
1C
b111 G
#333080000000
0!
0*
09
0>
0C
#333090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#333100000000
0!
0*
09
0>
0C
#333110000000
1!
1*
b1 6
19
1>
1C
b1 G
#333120000000
0!
0*
09
0>
0C
#333130000000
1!
1*
b10 6
19
1>
1C
b10 G
#333140000000
0!
0*
09
0>
0C
#333150000000
1!
1*
b11 6
19
1>
1C
b11 G
#333160000000
0!
0*
09
0>
0C
#333170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#333180000000
0!
0*
09
0>
0C
#333190000000
1!
1*
b101 6
19
1>
1C
b101 G
#333200000000
0!
0*
09
0>
0C
#333210000000
1!
1*
b110 6
19
1>
1C
b110 G
#333220000000
0!
0*
09
0>
0C
#333230000000
1!
1*
b111 6
19
1>
1C
b111 G
#333240000000
0!
1"
0*
1+
09
1:
0>
0C
#333250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#333260000000
0!
0*
09
0>
0C
#333270000000
1!
1*
b1 6
19
1>
1C
b1 G
#333280000000
0!
0*
09
0>
0C
#333290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#333300000000
0!
0*
09
0>
0C
#333310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#333320000000
0!
0*
09
0>
0C
#333330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#333340000000
0!
0*
09
0>
0C
#333350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#333360000000
0!
0#
0*
0,
09
0>
0?
0C
#333370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#333380000000
0!
0*
09
0>
0C
#333390000000
1!
1*
19
1>
1C
#333400000000
0!
0*
09
0>
0C
#333410000000
1!
1*
19
1>
1C
#333420000000
0!
0*
09
0>
0C
#333430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#333440000000
0!
0*
09
0>
0C
#333450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#333460000000
0!
0*
09
0>
0C
#333470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#333480000000
0!
0*
09
0>
0C
#333490000000
1!
1*
b10 6
19
1>
1C
b10 G
#333500000000
0!
0*
09
0>
0C
#333510000000
1!
1*
b11 6
19
1>
1C
b11 G
#333520000000
0!
0*
09
0>
0C
#333530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#333540000000
0!
0*
09
0>
0C
#333550000000
1!
1*
b101 6
19
1>
1C
b101 G
#333560000000
0!
0*
09
0>
0C
#333570000000
1!
1*
b110 6
19
1>
1C
b110 G
#333580000000
0!
0*
09
0>
0C
#333590000000
1!
1*
b111 6
19
1>
1C
b111 G
#333600000000
0!
0*
09
0>
0C
#333610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#333620000000
0!
0*
09
0>
0C
#333630000000
1!
1*
b1 6
19
1>
1C
b1 G
#333640000000
0!
0*
09
0>
0C
#333650000000
1!
1*
b10 6
19
1>
1C
b10 G
#333660000000
0!
0*
09
0>
0C
#333670000000
1!
1*
b11 6
19
1>
1C
b11 G
#333680000000
0!
0*
09
0>
0C
#333690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#333700000000
0!
0*
09
0>
0C
#333710000000
1!
1*
b101 6
19
1>
1C
b101 G
#333720000000
0!
0*
09
0>
0C
#333730000000
1!
1*
b110 6
19
1>
1C
b110 G
#333740000000
0!
0*
09
0>
0C
#333750000000
1!
1*
b111 6
19
1>
1C
b111 G
#333760000000
0!
0*
09
0>
0C
#333770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#333780000000
0!
0*
09
0>
0C
#333790000000
1!
1*
b1 6
19
1>
1C
b1 G
#333800000000
0!
0*
09
0>
0C
#333810000000
1!
1*
b10 6
19
1>
1C
b10 G
#333820000000
0!
0*
09
0>
0C
#333830000000
1!
1*
b11 6
19
1>
1C
b11 G
#333840000000
0!
0*
09
0>
0C
#333850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#333860000000
0!
0*
09
0>
0C
#333870000000
1!
1*
b101 6
19
1>
1C
b101 G
#333880000000
0!
0*
09
0>
0C
#333890000000
1!
1*
b110 6
19
1>
1C
b110 G
#333900000000
0!
0*
09
0>
0C
#333910000000
1!
1*
b111 6
19
1>
1C
b111 G
#333920000000
0!
1"
0*
1+
09
1:
0>
0C
#333930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#333940000000
0!
0*
09
0>
0C
#333950000000
1!
1*
b1 6
19
1>
1C
b1 G
#333960000000
0!
0*
09
0>
0C
#333970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#333980000000
0!
0*
09
0>
0C
#333990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#334000000000
0!
0*
09
0>
0C
#334010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#334020000000
0!
0*
09
0>
0C
#334030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#334040000000
0!
0#
0*
0,
09
0>
0?
0C
#334050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#334060000000
0!
0*
09
0>
0C
#334070000000
1!
1*
19
1>
1C
#334080000000
0!
0*
09
0>
0C
#334090000000
1!
1*
19
1>
1C
#334100000000
0!
0*
09
0>
0C
#334110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#334120000000
0!
0*
09
0>
0C
#334130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#334140000000
0!
0*
09
0>
0C
#334150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#334160000000
0!
0*
09
0>
0C
#334170000000
1!
1*
b10 6
19
1>
1C
b10 G
#334180000000
0!
0*
09
0>
0C
#334190000000
1!
1*
b11 6
19
1>
1C
b11 G
#334200000000
0!
0*
09
0>
0C
#334210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#334220000000
0!
0*
09
0>
0C
#334230000000
1!
1*
b101 6
19
1>
1C
b101 G
#334240000000
0!
0*
09
0>
0C
#334250000000
1!
1*
b110 6
19
1>
1C
b110 G
#334260000000
0!
0*
09
0>
0C
#334270000000
1!
1*
b111 6
19
1>
1C
b111 G
#334280000000
0!
0*
09
0>
0C
#334290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#334300000000
0!
0*
09
0>
0C
#334310000000
1!
1*
b1 6
19
1>
1C
b1 G
#334320000000
0!
0*
09
0>
0C
#334330000000
1!
1*
b10 6
19
1>
1C
b10 G
#334340000000
0!
0*
09
0>
0C
#334350000000
1!
1*
b11 6
19
1>
1C
b11 G
#334360000000
0!
0*
09
0>
0C
#334370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#334380000000
0!
0*
09
0>
0C
#334390000000
1!
1*
b101 6
19
1>
1C
b101 G
#334400000000
0!
0*
09
0>
0C
#334410000000
1!
1*
b110 6
19
1>
1C
b110 G
#334420000000
0!
0*
09
0>
0C
#334430000000
1!
1*
b111 6
19
1>
1C
b111 G
#334440000000
0!
0*
09
0>
0C
#334450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#334460000000
0!
0*
09
0>
0C
#334470000000
1!
1*
b1 6
19
1>
1C
b1 G
#334480000000
0!
0*
09
0>
0C
#334490000000
1!
1*
b10 6
19
1>
1C
b10 G
#334500000000
0!
0*
09
0>
0C
#334510000000
1!
1*
b11 6
19
1>
1C
b11 G
#334520000000
0!
0*
09
0>
0C
#334530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#334540000000
0!
0*
09
0>
0C
#334550000000
1!
1*
b101 6
19
1>
1C
b101 G
#334560000000
0!
0*
09
0>
0C
#334570000000
1!
1*
b110 6
19
1>
1C
b110 G
#334580000000
0!
0*
09
0>
0C
#334590000000
1!
1*
b111 6
19
1>
1C
b111 G
#334600000000
0!
1"
0*
1+
09
1:
0>
0C
#334610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#334620000000
0!
0*
09
0>
0C
#334630000000
1!
1*
b1 6
19
1>
1C
b1 G
#334640000000
0!
0*
09
0>
0C
#334650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#334660000000
0!
0*
09
0>
0C
#334670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#334680000000
0!
0*
09
0>
0C
#334690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#334700000000
0!
0*
09
0>
0C
#334710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#334720000000
0!
0#
0*
0,
09
0>
0?
0C
#334730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#334740000000
0!
0*
09
0>
0C
#334750000000
1!
1*
19
1>
1C
#334760000000
0!
0*
09
0>
0C
#334770000000
1!
1*
19
1>
1C
#334780000000
0!
0*
09
0>
0C
#334790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#334800000000
0!
0*
09
0>
0C
#334810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#334820000000
0!
0*
09
0>
0C
#334830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#334840000000
0!
0*
09
0>
0C
#334850000000
1!
1*
b10 6
19
1>
1C
b10 G
#334860000000
0!
0*
09
0>
0C
#334870000000
1!
1*
b11 6
19
1>
1C
b11 G
#334880000000
0!
0*
09
0>
0C
#334890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#334900000000
0!
0*
09
0>
0C
#334910000000
1!
1*
b101 6
19
1>
1C
b101 G
#334920000000
0!
0*
09
0>
0C
#334930000000
1!
1*
b110 6
19
1>
1C
b110 G
#334940000000
0!
0*
09
0>
0C
#334950000000
1!
1*
b111 6
19
1>
1C
b111 G
#334960000000
0!
0*
09
0>
0C
#334970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#334980000000
0!
0*
09
0>
0C
#334990000000
1!
1*
b1 6
19
1>
1C
b1 G
#335000000000
0!
0*
09
0>
0C
#335010000000
1!
1*
b10 6
19
1>
1C
b10 G
#335020000000
0!
0*
09
0>
0C
#335030000000
1!
1*
b11 6
19
1>
1C
b11 G
#335040000000
0!
0*
09
0>
0C
#335050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#335060000000
0!
0*
09
0>
0C
#335070000000
1!
1*
b101 6
19
1>
1C
b101 G
#335080000000
0!
0*
09
0>
0C
#335090000000
1!
1*
b110 6
19
1>
1C
b110 G
#335100000000
0!
0*
09
0>
0C
#335110000000
1!
1*
b111 6
19
1>
1C
b111 G
#335120000000
0!
0*
09
0>
0C
#335130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#335140000000
0!
0*
09
0>
0C
#335150000000
1!
1*
b1 6
19
1>
1C
b1 G
#335160000000
0!
0*
09
0>
0C
#335170000000
1!
1*
b10 6
19
1>
1C
b10 G
#335180000000
0!
0*
09
0>
0C
#335190000000
1!
1*
b11 6
19
1>
1C
b11 G
#335200000000
0!
0*
09
0>
0C
#335210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#335220000000
0!
0*
09
0>
0C
#335230000000
1!
1*
b101 6
19
1>
1C
b101 G
#335240000000
0!
0*
09
0>
0C
#335250000000
1!
1*
b110 6
19
1>
1C
b110 G
#335260000000
0!
0*
09
0>
0C
#335270000000
1!
1*
b111 6
19
1>
1C
b111 G
#335280000000
0!
1"
0*
1+
09
1:
0>
0C
#335290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#335300000000
0!
0*
09
0>
0C
#335310000000
1!
1*
b1 6
19
1>
1C
b1 G
#335320000000
0!
0*
09
0>
0C
#335330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#335340000000
0!
0*
09
0>
0C
#335350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#335360000000
0!
0*
09
0>
0C
#335370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#335380000000
0!
0*
09
0>
0C
#335390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#335400000000
0!
0#
0*
0,
09
0>
0?
0C
#335410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#335420000000
0!
0*
09
0>
0C
#335430000000
1!
1*
19
1>
1C
#335440000000
0!
0*
09
0>
0C
#335450000000
1!
1*
19
1>
1C
#335460000000
0!
0*
09
0>
0C
#335470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#335480000000
0!
0*
09
0>
0C
#335490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#335500000000
0!
0*
09
0>
0C
#335510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#335520000000
0!
0*
09
0>
0C
#335530000000
1!
1*
b10 6
19
1>
1C
b10 G
#335540000000
0!
0*
09
0>
0C
#335550000000
1!
1*
b11 6
19
1>
1C
b11 G
#335560000000
0!
0*
09
0>
0C
#335570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#335580000000
0!
0*
09
0>
0C
#335590000000
1!
1*
b101 6
19
1>
1C
b101 G
#335600000000
0!
0*
09
0>
0C
#335610000000
1!
1*
b110 6
19
1>
1C
b110 G
#335620000000
0!
0*
09
0>
0C
#335630000000
1!
1*
b111 6
19
1>
1C
b111 G
#335640000000
0!
0*
09
0>
0C
#335650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#335660000000
0!
0*
09
0>
0C
#335670000000
1!
1*
b1 6
19
1>
1C
b1 G
#335680000000
0!
0*
09
0>
0C
#335690000000
1!
1*
b10 6
19
1>
1C
b10 G
#335700000000
0!
0*
09
0>
0C
#335710000000
1!
1*
b11 6
19
1>
1C
b11 G
#335720000000
0!
0*
09
0>
0C
#335730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#335740000000
0!
0*
09
0>
0C
#335750000000
1!
1*
b101 6
19
1>
1C
b101 G
#335760000000
0!
0*
09
0>
0C
#335770000000
1!
1*
b110 6
19
1>
1C
b110 G
#335780000000
0!
0*
09
0>
0C
#335790000000
1!
1*
b111 6
19
1>
1C
b111 G
#335800000000
0!
0*
09
0>
0C
#335810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#335820000000
0!
0*
09
0>
0C
#335830000000
1!
1*
b1 6
19
1>
1C
b1 G
#335840000000
0!
0*
09
0>
0C
#335850000000
1!
1*
b10 6
19
1>
1C
b10 G
#335860000000
0!
0*
09
0>
0C
#335870000000
1!
1*
b11 6
19
1>
1C
b11 G
#335880000000
0!
0*
09
0>
0C
#335890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#335900000000
0!
0*
09
0>
0C
#335910000000
1!
1*
b101 6
19
1>
1C
b101 G
#335920000000
0!
0*
09
0>
0C
#335930000000
1!
1*
b110 6
19
1>
1C
b110 G
#335940000000
0!
0*
09
0>
0C
#335950000000
1!
1*
b111 6
19
1>
1C
b111 G
#335960000000
0!
1"
0*
1+
09
1:
0>
0C
#335970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#335980000000
0!
0*
09
0>
0C
#335990000000
1!
1*
b1 6
19
1>
1C
b1 G
#336000000000
0!
0*
09
0>
0C
#336010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#336020000000
0!
0*
09
0>
0C
#336030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#336040000000
0!
0*
09
0>
0C
#336050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#336060000000
0!
0*
09
0>
0C
#336070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#336080000000
0!
0#
0*
0,
09
0>
0?
0C
#336090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#336100000000
0!
0*
09
0>
0C
#336110000000
1!
1*
19
1>
1C
#336120000000
0!
0*
09
0>
0C
#336130000000
1!
1*
19
1>
1C
#336140000000
0!
0*
09
0>
0C
#336150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#336160000000
0!
0*
09
0>
0C
#336170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#336180000000
0!
0*
09
0>
0C
#336190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#336200000000
0!
0*
09
0>
0C
#336210000000
1!
1*
b10 6
19
1>
1C
b10 G
#336220000000
0!
0*
09
0>
0C
#336230000000
1!
1*
b11 6
19
1>
1C
b11 G
#336240000000
0!
0*
09
0>
0C
#336250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#336260000000
0!
0*
09
0>
0C
#336270000000
1!
1*
b101 6
19
1>
1C
b101 G
#336280000000
0!
0*
09
0>
0C
#336290000000
1!
1*
b110 6
19
1>
1C
b110 G
#336300000000
0!
0*
09
0>
0C
#336310000000
1!
1*
b111 6
19
1>
1C
b111 G
#336320000000
0!
0*
09
0>
0C
#336330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#336340000000
0!
0*
09
0>
0C
#336350000000
1!
1*
b1 6
19
1>
1C
b1 G
#336360000000
0!
0*
09
0>
0C
#336370000000
1!
1*
b10 6
19
1>
1C
b10 G
#336380000000
0!
0*
09
0>
0C
#336390000000
1!
1*
b11 6
19
1>
1C
b11 G
#336400000000
0!
0*
09
0>
0C
#336410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#336420000000
0!
0*
09
0>
0C
#336430000000
1!
1*
b101 6
19
1>
1C
b101 G
#336440000000
0!
0*
09
0>
0C
#336450000000
1!
1*
b110 6
19
1>
1C
b110 G
#336460000000
0!
0*
09
0>
0C
#336470000000
1!
1*
b111 6
19
1>
1C
b111 G
#336480000000
0!
0*
09
0>
0C
#336490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#336500000000
0!
0*
09
0>
0C
#336510000000
1!
1*
b1 6
19
1>
1C
b1 G
#336520000000
0!
0*
09
0>
0C
#336530000000
1!
1*
b10 6
19
1>
1C
b10 G
#336540000000
0!
0*
09
0>
0C
#336550000000
1!
1*
b11 6
19
1>
1C
b11 G
#336560000000
0!
0*
09
0>
0C
#336570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#336580000000
0!
0*
09
0>
0C
#336590000000
1!
1*
b101 6
19
1>
1C
b101 G
#336600000000
0!
0*
09
0>
0C
#336610000000
1!
1*
b110 6
19
1>
1C
b110 G
#336620000000
0!
0*
09
0>
0C
#336630000000
1!
1*
b111 6
19
1>
1C
b111 G
#336640000000
0!
1"
0*
1+
09
1:
0>
0C
#336650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#336660000000
0!
0*
09
0>
0C
#336670000000
1!
1*
b1 6
19
1>
1C
b1 G
#336680000000
0!
0*
09
0>
0C
#336690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#336700000000
0!
0*
09
0>
0C
#336710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#336720000000
0!
0*
09
0>
0C
#336730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#336740000000
0!
0*
09
0>
0C
#336750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#336760000000
0!
0#
0*
0,
09
0>
0?
0C
#336770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#336780000000
0!
0*
09
0>
0C
#336790000000
1!
1*
19
1>
1C
#336800000000
0!
0*
09
0>
0C
#336810000000
1!
1*
19
1>
1C
#336820000000
0!
0*
09
0>
0C
#336830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#336840000000
0!
0*
09
0>
0C
#336850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#336860000000
0!
0*
09
0>
0C
#336870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#336880000000
0!
0*
09
0>
0C
#336890000000
1!
1*
b10 6
19
1>
1C
b10 G
#336900000000
0!
0*
09
0>
0C
#336910000000
1!
1*
b11 6
19
1>
1C
b11 G
#336920000000
0!
0*
09
0>
0C
#336930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#336940000000
0!
0*
09
0>
0C
#336950000000
1!
1*
b101 6
19
1>
1C
b101 G
#336960000000
0!
0*
09
0>
0C
#336970000000
1!
1*
b110 6
19
1>
1C
b110 G
#336980000000
0!
0*
09
0>
0C
#336990000000
1!
1*
b111 6
19
1>
1C
b111 G
#337000000000
0!
0*
09
0>
0C
#337010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#337020000000
0!
0*
09
0>
0C
#337030000000
1!
1*
b1 6
19
1>
1C
b1 G
#337040000000
0!
0*
09
0>
0C
#337050000000
1!
1*
b10 6
19
1>
1C
b10 G
#337060000000
0!
0*
09
0>
0C
#337070000000
1!
1*
b11 6
19
1>
1C
b11 G
#337080000000
0!
0*
09
0>
0C
#337090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#337100000000
0!
0*
09
0>
0C
#337110000000
1!
1*
b101 6
19
1>
1C
b101 G
#337120000000
0!
0*
09
0>
0C
#337130000000
1!
1*
b110 6
19
1>
1C
b110 G
#337140000000
0!
0*
09
0>
0C
#337150000000
1!
1*
b111 6
19
1>
1C
b111 G
#337160000000
0!
0*
09
0>
0C
#337170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#337180000000
0!
0*
09
0>
0C
#337190000000
1!
1*
b1 6
19
1>
1C
b1 G
#337200000000
0!
0*
09
0>
0C
#337210000000
1!
1*
b10 6
19
1>
1C
b10 G
#337220000000
0!
0*
09
0>
0C
#337230000000
1!
1*
b11 6
19
1>
1C
b11 G
#337240000000
0!
0*
09
0>
0C
#337250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#337260000000
0!
0*
09
0>
0C
#337270000000
1!
1*
b101 6
19
1>
1C
b101 G
#337280000000
0!
0*
09
0>
0C
#337290000000
1!
1*
b110 6
19
1>
1C
b110 G
#337300000000
0!
0*
09
0>
0C
#337310000000
1!
1*
b111 6
19
1>
1C
b111 G
#337320000000
0!
1"
0*
1+
09
1:
0>
0C
#337330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#337340000000
0!
0*
09
0>
0C
#337350000000
1!
1*
b1 6
19
1>
1C
b1 G
#337360000000
0!
0*
09
0>
0C
#337370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#337380000000
0!
0*
09
0>
0C
#337390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#337400000000
0!
0*
09
0>
0C
#337410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#337420000000
0!
0*
09
0>
0C
#337430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#337440000000
0!
0#
0*
0,
09
0>
0?
0C
#337450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#337460000000
0!
0*
09
0>
0C
#337470000000
1!
1*
19
1>
1C
#337480000000
0!
0*
09
0>
0C
#337490000000
1!
1*
19
1>
1C
#337500000000
0!
0*
09
0>
0C
#337510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#337520000000
0!
0*
09
0>
0C
#337530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#337540000000
0!
0*
09
0>
0C
#337550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#337560000000
0!
0*
09
0>
0C
#337570000000
1!
1*
b10 6
19
1>
1C
b10 G
#337580000000
0!
0*
09
0>
0C
#337590000000
1!
1*
b11 6
19
1>
1C
b11 G
#337600000000
0!
0*
09
0>
0C
#337610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#337620000000
0!
0*
09
0>
0C
#337630000000
1!
1*
b101 6
19
1>
1C
b101 G
#337640000000
0!
0*
09
0>
0C
#337650000000
1!
1*
b110 6
19
1>
1C
b110 G
#337660000000
0!
0*
09
0>
0C
#337670000000
1!
1*
b111 6
19
1>
1C
b111 G
#337680000000
0!
0*
09
0>
0C
#337690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#337700000000
0!
0*
09
0>
0C
#337710000000
1!
1*
b1 6
19
1>
1C
b1 G
#337720000000
0!
0*
09
0>
0C
#337730000000
1!
1*
b10 6
19
1>
1C
b10 G
#337740000000
0!
0*
09
0>
0C
#337750000000
1!
1*
b11 6
19
1>
1C
b11 G
#337760000000
0!
0*
09
0>
0C
#337770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#337780000000
0!
0*
09
0>
0C
#337790000000
1!
1*
b101 6
19
1>
1C
b101 G
#337800000000
0!
0*
09
0>
0C
#337810000000
1!
1*
b110 6
19
1>
1C
b110 G
#337820000000
0!
0*
09
0>
0C
#337830000000
1!
1*
b111 6
19
1>
1C
b111 G
#337840000000
0!
0*
09
0>
0C
#337850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#337860000000
0!
0*
09
0>
0C
#337870000000
1!
1*
b1 6
19
1>
1C
b1 G
#337880000000
0!
0*
09
0>
0C
#337890000000
1!
1*
b10 6
19
1>
1C
b10 G
#337900000000
0!
0*
09
0>
0C
#337910000000
1!
1*
b11 6
19
1>
1C
b11 G
#337920000000
0!
0*
09
0>
0C
#337930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#337940000000
0!
0*
09
0>
0C
#337950000000
1!
1*
b101 6
19
1>
1C
b101 G
#337960000000
0!
0*
09
0>
0C
#337970000000
1!
1*
b110 6
19
1>
1C
b110 G
#337980000000
0!
0*
09
0>
0C
#337990000000
1!
1*
b111 6
19
1>
1C
b111 G
#338000000000
0!
1"
0*
1+
09
1:
0>
0C
#338010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#338020000000
0!
0*
09
0>
0C
#338030000000
1!
1*
b1 6
19
1>
1C
b1 G
#338040000000
0!
0*
09
0>
0C
#338050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#338060000000
0!
0*
09
0>
0C
#338070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#338080000000
0!
0*
09
0>
0C
#338090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#338100000000
0!
0*
09
0>
0C
#338110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#338120000000
0!
0#
0*
0,
09
0>
0?
0C
#338130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#338140000000
0!
0*
09
0>
0C
#338150000000
1!
1*
19
1>
1C
#338160000000
0!
0*
09
0>
0C
#338170000000
1!
1*
19
1>
1C
#338180000000
0!
0*
09
0>
0C
#338190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#338200000000
0!
0*
09
0>
0C
#338210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#338220000000
0!
0*
09
0>
0C
#338230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#338240000000
0!
0*
09
0>
0C
#338250000000
1!
1*
b10 6
19
1>
1C
b10 G
#338260000000
0!
0*
09
0>
0C
#338270000000
1!
1*
b11 6
19
1>
1C
b11 G
#338280000000
0!
0*
09
0>
0C
#338290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#338300000000
0!
0*
09
0>
0C
#338310000000
1!
1*
b101 6
19
1>
1C
b101 G
#338320000000
0!
0*
09
0>
0C
#338330000000
1!
1*
b110 6
19
1>
1C
b110 G
#338340000000
0!
0*
09
0>
0C
#338350000000
1!
1*
b111 6
19
1>
1C
b111 G
#338360000000
0!
0*
09
0>
0C
#338370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#338380000000
0!
0*
09
0>
0C
#338390000000
1!
1*
b1 6
19
1>
1C
b1 G
#338400000000
0!
0*
09
0>
0C
#338410000000
1!
1*
b10 6
19
1>
1C
b10 G
#338420000000
0!
0*
09
0>
0C
#338430000000
1!
1*
b11 6
19
1>
1C
b11 G
#338440000000
0!
0*
09
0>
0C
#338450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#338460000000
0!
0*
09
0>
0C
#338470000000
1!
1*
b101 6
19
1>
1C
b101 G
#338480000000
0!
0*
09
0>
0C
#338490000000
1!
1*
b110 6
19
1>
1C
b110 G
#338500000000
0!
0*
09
0>
0C
#338510000000
1!
1*
b111 6
19
1>
1C
b111 G
#338520000000
0!
0*
09
0>
0C
#338530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#338540000000
0!
0*
09
0>
0C
#338550000000
1!
1*
b1 6
19
1>
1C
b1 G
#338560000000
0!
0*
09
0>
0C
#338570000000
1!
1*
b10 6
19
1>
1C
b10 G
#338580000000
0!
0*
09
0>
0C
#338590000000
1!
1*
b11 6
19
1>
1C
b11 G
#338600000000
0!
0*
09
0>
0C
#338610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#338620000000
0!
0*
09
0>
0C
#338630000000
1!
1*
b101 6
19
1>
1C
b101 G
#338640000000
0!
0*
09
0>
0C
#338650000000
1!
1*
b110 6
19
1>
1C
b110 G
#338660000000
0!
0*
09
0>
0C
#338670000000
1!
1*
b111 6
19
1>
1C
b111 G
#338680000000
0!
1"
0*
1+
09
1:
0>
0C
#338690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#338700000000
0!
0*
09
0>
0C
#338710000000
1!
1*
b1 6
19
1>
1C
b1 G
#338720000000
0!
0*
09
0>
0C
#338730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#338740000000
0!
0*
09
0>
0C
#338750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#338760000000
0!
0*
09
0>
0C
#338770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#338780000000
0!
0*
09
0>
0C
#338790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#338800000000
0!
0#
0*
0,
09
0>
0?
0C
#338810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#338820000000
0!
0*
09
0>
0C
#338830000000
1!
1*
19
1>
1C
#338840000000
0!
0*
09
0>
0C
#338850000000
1!
1*
19
1>
1C
#338860000000
0!
0*
09
0>
0C
#338870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#338880000000
0!
0*
09
0>
0C
#338890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#338900000000
0!
0*
09
0>
0C
#338910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#338920000000
0!
0*
09
0>
0C
#338930000000
1!
1*
b10 6
19
1>
1C
b10 G
#338940000000
0!
0*
09
0>
0C
#338950000000
1!
1*
b11 6
19
1>
1C
b11 G
#338960000000
0!
0*
09
0>
0C
#338970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#338980000000
0!
0*
09
0>
0C
#338990000000
1!
1*
b101 6
19
1>
1C
b101 G
#339000000000
0!
0*
09
0>
0C
#339010000000
1!
1*
b110 6
19
1>
1C
b110 G
#339020000000
0!
0*
09
0>
0C
#339030000000
1!
1*
b111 6
19
1>
1C
b111 G
#339040000000
0!
0*
09
0>
0C
#339050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#339060000000
0!
0*
09
0>
0C
#339070000000
1!
1*
b1 6
19
1>
1C
b1 G
#339080000000
0!
0*
09
0>
0C
#339090000000
1!
1*
b10 6
19
1>
1C
b10 G
#339100000000
0!
0*
09
0>
0C
#339110000000
1!
1*
b11 6
19
1>
1C
b11 G
#339120000000
0!
0*
09
0>
0C
#339130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#339140000000
0!
0*
09
0>
0C
#339150000000
1!
1*
b101 6
19
1>
1C
b101 G
#339160000000
0!
0*
09
0>
0C
#339170000000
1!
1*
b110 6
19
1>
1C
b110 G
#339180000000
0!
0*
09
0>
0C
#339190000000
1!
1*
b111 6
19
1>
1C
b111 G
#339200000000
0!
0*
09
0>
0C
#339210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#339220000000
0!
0*
09
0>
0C
#339230000000
1!
1*
b1 6
19
1>
1C
b1 G
#339240000000
0!
0*
09
0>
0C
#339250000000
1!
1*
b10 6
19
1>
1C
b10 G
#339260000000
0!
0*
09
0>
0C
#339270000000
1!
1*
b11 6
19
1>
1C
b11 G
#339280000000
0!
0*
09
0>
0C
#339290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#339300000000
0!
0*
09
0>
0C
#339310000000
1!
1*
b101 6
19
1>
1C
b101 G
#339320000000
0!
0*
09
0>
0C
#339330000000
1!
1*
b110 6
19
1>
1C
b110 G
#339340000000
0!
0*
09
0>
0C
#339350000000
1!
1*
b111 6
19
1>
1C
b111 G
#339360000000
0!
1"
0*
1+
09
1:
0>
0C
#339370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#339380000000
0!
0*
09
0>
0C
#339390000000
1!
1*
b1 6
19
1>
1C
b1 G
#339400000000
0!
0*
09
0>
0C
#339410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#339420000000
0!
0*
09
0>
0C
#339430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#339440000000
0!
0*
09
0>
0C
#339450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#339460000000
0!
0*
09
0>
0C
#339470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#339480000000
0!
0#
0*
0,
09
0>
0?
0C
#339490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#339500000000
0!
0*
09
0>
0C
#339510000000
1!
1*
19
1>
1C
#339520000000
0!
0*
09
0>
0C
#339530000000
1!
1*
19
1>
1C
#339540000000
0!
0*
09
0>
0C
#339550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#339560000000
0!
0*
09
0>
0C
#339570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#339580000000
0!
0*
09
0>
0C
#339590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#339600000000
0!
0*
09
0>
0C
#339610000000
1!
1*
b10 6
19
1>
1C
b10 G
#339620000000
0!
0*
09
0>
0C
#339630000000
1!
1*
b11 6
19
1>
1C
b11 G
#339640000000
0!
0*
09
0>
0C
#339650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#339660000000
0!
0*
09
0>
0C
#339670000000
1!
1*
b101 6
19
1>
1C
b101 G
#339680000000
0!
0*
09
0>
0C
#339690000000
1!
1*
b110 6
19
1>
1C
b110 G
#339700000000
0!
0*
09
0>
0C
#339710000000
1!
1*
b111 6
19
1>
1C
b111 G
#339720000000
0!
0*
09
0>
0C
#339730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#339740000000
0!
0*
09
0>
0C
#339750000000
1!
1*
b1 6
19
1>
1C
b1 G
#339760000000
0!
0*
09
0>
0C
#339770000000
1!
1*
b10 6
19
1>
1C
b10 G
#339780000000
0!
0*
09
0>
0C
#339790000000
1!
1*
b11 6
19
1>
1C
b11 G
#339800000000
0!
0*
09
0>
0C
#339810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#339820000000
0!
0*
09
0>
0C
#339830000000
1!
1*
b101 6
19
1>
1C
b101 G
#339840000000
0!
0*
09
0>
0C
#339850000000
1!
1*
b110 6
19
1>
1C
b110 G
#339860000000
0!
0*
09
0>
0C
#339870000000
1!
1*
b111 6
19
1>
1C
b111 G
#339880000000
0!
0*
09
0>
0C
#339890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#339900000000
0!
0*
09
0>
0C
#339910000000
1!
1*
b1 6
19
1>
1C
b1 G
#339920000000
0!
0*
09
0>
0C
#339930000000
1!
1*
b10 6
19
1>
1C
b10 G
#339940000000
0!
0*
09
0>
0C
#339950000000
1!
1*
b11 6
19
1>
1C
b11 G
#339960000000
0!
0*
09
0>
0C
#339970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#339980000000
0!
0*
09
0>
0C
#339990000000
1!
1*
b101 6
19
1>
1C
b101 G
#340000000000
0!
0*
09
0>
0C
#340010000000
1!
1*
b110 6
19
1>
1C
b110 G
#340020000000
0!
0*
09
0>
0C
#340030000000
1!
1*
b111 6
19
1>
1C
b111 G
#340040000000
0!
1"
0*
1+
09
1:
0>
0C
#340050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#340060000000
0!
0*
09
0>
0C
#340070000000
1!
1*
b1 6
19
1>
1C
b1 G
#340080000000
0!
0*
09
0>
0C
#340090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#340100000000
0!
0*
09
0>
0C
#340110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#340120000000
0!
0*
09
0>
0C
#340130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#340140000000
0!
0*
09
0>
0C
#340150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#340160000000
0!
0#
0*
0,
09
0>
0?
0C
#340170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#340180000000
0!
0*
09
0>
0C
#340190000000
1!
1*
19
1>
1C
#340200000000
0!
0*
09
0>
0C
#340210000000
1!
1*
19
1>
1C
#340220000000
0!
0*
09
0>
0C
#340230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#340240000000
0!
0*
09
0>
0C
#340250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#340260000000
0!
0*
09
0>
0C
#340270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#340280000000
0!
0*
09
0>
0C
#340290000000
1!
1*
b10 6
19
1>
1C
b10 G
#340300000000
0!
0*
09
0>
0C
#340310000000
1!
1*
b11 6
19
1>
1C
b11 G
#340320000000
0!
0*
09
0>
0C
#340330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#340340000000
0!
0*
09
0>
0C
#340350000000
1!
1*
b101 6
19
1>
1C
b101 G
#340360000000
0!
0*
09
0>
0C
#340370000000
1!
1*
b110 6
19
1>
1C
b110 G
#340380000000
0!
0*
09
0>
0C
#340390000000
1!
1*
b111 6
19
1>
1C
b111 G
#340400000000
0!
0*
09
0>
0C
#340410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#340420000000
0!
0*
09
0>
0C
#340430000000
1!
1*
b1 6
19
1>
1C
b1 G
#340440000000
0!
0*
09
0>
0C
#340450000000
1!
1*
b10 6
19
1>
1C
b10 G
#340460000000
0!
0*
09
0>
0C
#340470000000
1!
1*
b11 6
19
1>
1C
b11 G
#340480000000
0!
0*
09
0>
0C
#340490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#340500000000
0!
0*
09
0>
0C
#340510000000
1!
1*
b101 6
19
1>
1C
b101 G
#340520000000
0!
0*
09
0>
0C
#340530000000
1!
1*
b110 6
19
1>
1C
b110 G
#340540000000
0!
0*
09
0>
0C
#340550000000
1!
1*
b111 6
19
1>
1C
b111 G
#340560000000
0!
0*
09
0>
0C
#340570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#340580000000
0!
0*
09
0>
0C
#340590000000
1!
1*
b1 6
19
1>
1C
b1 G
#340600000000
0!
0*
09
0>
0C
#340610000000
1!
1*
b10 6
19
1>
1C
b10 G
#340620000000
0!
0*
09
0>
0C
#340630000000
1!
1*
b11 6
19
1>
1C
b11 G
#340640000000
0!
0*
09
0>
0C
#340650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#340660000000
0!
0*
09
0>
0C
#340670000000
1!
1*
b101 6
19
1>
1C
b101 G
#340680000000
0!
0*
09
0>
0C
#340690000000
1!
1*
b110 6
19
1>
1C
b110 G
#340700000000
0!
0*
09
0>
0C
#340710000000
1!
1*
b111 6
19
1>
1C
b111 G
#340720000000
0!
1"
0*
1+
09
1:
0>
0C
#340730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#340740000000
0!
0*
09
0>
0C
#340750000000
1!
1*
b1 6
19
1>
1C
b1 G
#340760000000
0!
0*
09
0>
0C
#340770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#340780000000
0!
0*
09
0>
0C
#340790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#340800000000
0!
0*
09
0>
0C
#340810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#340820000000
0!
0*
09
0>
0C
#340830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#340840000000
0!
0#
0*
0,
09
0>
0?
0C
#340850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#340860000000
0!
0*
09
0>
0C
#340870000000
1!
1*
19
1>
1C
#340880000000
0!
0*
09
0>
0C
#340890000000
1!
1*
19
1>
1C
#340900000000
0!
0*
09
0>
0C
#340910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#340920000000
0!
0*
09
0>
0C
#340930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#340940000000
0!
0*
09
0>
0C
#340950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#340960000000
0!
0*
09
0>
0C
#340970000000
1!
1*
b10 6
19
1>
1C
b10 G
#340980000000
0!
0*
09
0>
0C
#340990000000
1!
1*
b11 6
19
1>
1C
b11 G
#341000000000
0!
0*
09
0>
0C
#341010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#341020000000
0!
0*
09
0>
0C
#341030000000
1!
1*
b101 6
19
1>
1C
b101 G
#341040000000
0!
0*
09
0>
0C
#341050000000
1!
1*
b110 6
19
1>
1C
b110 G
#341060000000
0!
0*
09
0>
0C
#341070000000
1!
1*
b111 6
19
1>
1C
b111 G
#341080000000
0!
0*
09
0>
0C
#341090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#341100000000
0!
0*
09
0>
0C
#341110000000
1!
1*
b1 6
19
1>
1C
b1 G
#341120000000
0!
0*
09
0>
0C
#341130000000
1!
1*
b10 6
19
1>
1C
b10 G
#341140000000
0!
0*
09
0>
0C
#341150000000
1!
1*
b11 6
19
1>
1C
b11 G
#341160000000
0!
0*
09
0>
0C
#341170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#341180000000
0!
0*
09
0>
0C
#341190000000
1!
1*
b101 6
19
1>
1C
b101 G
#341200000000
0!
0*
09
0>
0C
#341210000000
1!
1*
b110 6
19
1>
1C
b110 G
#341220000000
0!
0*
09
0>
0C
#341230000000
1!
1*
b111 6
19
1>
1C
b111 G
#341240000000
0!
0*
09
0>
0C
#341250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#341260000000
0!
0*
09
0>
0C
#341270000000
1!
1*
b1 6
19
1>
1C
b1 G
#341280000000
0!
0*
09
0>
0C
#341290000000
1!
1*
b10 6
19
1>
1C
b10 G
#341300000000
0!
0*
09
0>
0C
#341310000000
1!
1*
b11 6
19
1>
1C
b11 G
#341320000000
0!
0*
09
0>
0C
#341330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#341340000000
0!
0*
09
0>
0C
#341350000000
1!
1*
b101 6
19
1>
1C
b101 G
#341360000000
0!
0*
09
0>
0C
#341370000000
1!
1*
b110 6
19
1>
1C
b110 G
#341380000000
0!
0*
09
0>
0C
#341390000000
1!
1*
b111 6
19
1>
1C
b111 G
#341400000000
0!
1"
0*
1+
09
1:
0>
0C
#341410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#341420000000
0!
0*
09
0>
0C
#341430000000
1!
1*
b1 6
19
1>
1C
b1 G
#341440000000
0!
0*
09
0>
0C
#341450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#341460000000
0!
0*
09
0>
0C
#341470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#341480000000
0!
0*
09
0>
0C
#341490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#341500000000
0!
0*
09
0>
0C
#341510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#341520000000
0!
0#
0*
0,
09
0>
0?
0C
#341530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#341540000000
0!
0*
09
0>
0C
#341550000000
1!
1*
19
1>
1C
#341560000000
0!
0*
09
0>
0C
#341570000000
1!
1*
19
1>
1C
#341580000000
0!
0*
09
0>
0C
#341590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#341600000000
0!
0*
09
0>
0C
#341610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#341620000000
0!
0*
09
0>
0C
#341630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#341640000000
0!
0*
09
0>
0C
#341650000000
1!
1*
b10 6
19
1>
1C
b10 G
#341660000000
0!
0*
09
0>
0C
#341670000000
1!
1*
b11 6
19
1>
1C
b11 G
#341680000000
0!
0*
09
0>
0C
#341690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#341700000000
0!
0*
09
0>
0C
#341710000000
1!
1*
b101 6
19
1>
1C
b101 G
#341720000000
0!
0*
09
0>
0C
#341730000000
1!
1*
b110 6
19
1>
1C
b110 G
#341740000000
0!
0*
09
0>
0C
#341750000000
1!
1*
b111 6
19
1>
1C
b111 G
#341760000000
0!
0*
09
0>
0C
#341770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#341780000000
0!
0*
09
0>
0C
#341790000000
1!
1*
b1 6
19
1>
1C
b1 G
#341800000000
0!
0*
09
0>
0C
#341810000000
1!
1*
b10 6
19
1>
1C
b10 G
#341820000000
0!
0*
09
0>
0C
#341830000000
1!
1*
b11 6
19
1>
1C
b11 G
#341840000000
0!
0*
09
0>
0C
#341850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#341860000000
0!
0*
09
0>
0C
#341870000000
1!
1*
b101 6
19
1>
1C
b101 G
#341880000000
0!
0*
09
0>
0C
#341890000000
1!
1*
b110 6
19
1>
1C
b110 G
#341900000000
0!
0*
09
0>
0C
#341910000000
1!
1*
b111 6
19
1>
1C
b111 G
#341920000000
0!
0*
09
0>
0C
#341930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#341940000000
0!
0*
09
0>
0C
#341950000000
1!
1*
b1 6
19
1>
1C
b1 G
#341960000000
0!
0*
09
0>
0C
#341970000000
1!
1*
b10 6
19
1>
1C
b10 G
#341980000000
0!
0*
09
0>
0C
#341990000000
1!
1*
b11 6
19
1>
1C
b11 G
#342000000000
0!
0*
09
0>
0C
#342010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#342020000000
0!
0*
09
0>
0C
#342030000000
1!
1*
b101 6
19
1>
1C
b101 G
#342040000000
0!
0*
09
0>
0C
#342050000000
1!
1*
b110 6
19
1>
1C
b110 G
#342060000000
0!
0*
09
0>
0C
#342070000000
1!
1*
b111 6
19
1>
1C
b111 G
#342080000000
0!
1"
0*
1+
09
1:
0>
0C
#342090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#342100000000
0!
0*
09
0>
0C
#342110000000
1!
1*
b1 6
19
1>
1C
b1 G
#342120000000
0!
0*
09
0>
0C
#342130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#342140000000
0!
0*
09
0>
0C
#342150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#342160000000
0!
0*
09
0>
0C
#342170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#342180000000
0!
0*
09
0>
0C
#342190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#342200000000
0!
0#
0*
0,
09
0>
0?
0C
#342210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#342220000000
0!
0*
09
0>
0C
#342230000000
1!
1*
19
1>
1C
#342240000000
0!
0*
09
0>
0C
#342250000000
1!
1*
19
1>
1C
#342260000000
0!
0*
09
0>
0C
#342270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#342280000000
0!
0*
09
0>
0C
#342290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#342300000000
0!
0*
09
0>
0C
#342310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#342320000000
0!
0*
09
0>
0C
#342330000000
1!
1*
b10 6
19
1>
1C
b10 G
#342340000000
0!
0*
09
0>
0C
#342350000000
1!
1*
b11 6
19
1>
1C
b11 G
#342360000000
0!
0*
09
0>
0C
#342370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#342380000000
0!
0*
09
0>
0C
#342390000000
1!
1*
b101 6
19
1>
1C
b101 G
#342400000000
0!
0*
09
0>
0C
#342410000000
1!
1*
b110 6
19
1>
1C
b110 G
#342420000000
0!
0*
09
0>
0C
#342430000000
1!
1*
b111 6
19
1>
1C
b111 G
#342440000000
0!
0*
09
0>
0C
#342450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#342460000000
0!
0*
09
0>
0C
#342470000000
1!
1*
b1 6
19
1>
1C
b1 G
#342480000000
0!
0*
09
0>
0C
#342490000000
1!
1*
b10 6
19
1>
1C
b10 G
#342500000000
0!
0*
09
0>
0C
#342510000000
1!
1*
b11 6
19
1>
1C
b11 G
#342520000000
0!
0*
09
0>
0C
#342530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#342540000000
0!
0*
09
0>
0C
#342550000000
1!
1*
b101 6
19
1>
1C
b101 G
#342560000000
0!
0*
09
0>
0C
#342570000000
1!
1*
b110 6
19
1>
1C
b110 G
#342580000000
0!
0*
09
0>
0C
#342590000000
1!
1*
b111 6
19
1>
1C
b111 G
#342600000000
0!
0*
09
0>
0C
#342610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#342620000000
0!
0*
09
0>
0C
#342630000000
1!
1*
b1 6
19
1>
1C
b1 G
#342640000000
0!
0*
09
0>
0C
#342650000000
1!
1*
b10 6
19
1>
1C
b10 G
#342660000000
0!
0*
09
0>
0C
#342670000000
1!
1*
b11 6
19
1>
1C
b11 G
#342680000000
0!
0*
09
0>
0C
#342690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#342700000000
0!
0*
09
0>
0C
#342710000000
1!
1*
b101 6
19
1>
1C
b101 G
#342720000000
0!
0*
09
0>
0C
#342730000000
1!
1*
b110 6
19
1>
1C
b110 G
#342740000000
0!
0*
09
0>
0C
#342750000000
1!
1*
b111 6
19
1>
1C
b111 G
#342760000000
0!
1"
0*
1+
09
1:
0>
0C
#342770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#342780000000
0!
0*
09
0>
0C
#342790000000
1!
1*
b1 6
19
1>
1C
b1 G
#342800000000
0!
0*
09
0>
0C
#342810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#342820000000
0!
0*
09
0>
0C
#342830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#342840000000
0!
0*
09
0>
0C
#342850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#342860000000
0!
0*
09
0>
0C
#342870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#342880000000
0!
0#
0*
0,
09
0>
0?
0C
#342890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#342900000000
0!
0*
09
0>
0C
#342910000000
1!
1*
19
1>
1C
#342920000000
0!
0*
09
0>
0C
#342930000000
1!
1*
19
1>
1C
#342940000000
0!
0*
09
0>
0C
#342950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#342960000000
0!
0*
09
0>
0C
#342970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#342980000000
0!
0*
09
0>
0C
#342990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#343000000000
0!
0*
09
0>
0C
#343010000000
1!
1*
b10 6
19
1>
1C
b10 G
#343020000000
0!
0*
09
0>
0C
#343030000000
1!
1*
b11 6
19
1>
1C
b11 G
#343040000000
0!
0*
09
0>
0C
#343050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#343060000000
0!
0*
09
0>
0C
#343070000000
1!
1*
b101 6
19
1>
1C
b101 G
#343080000000
0!
0*
09
0>
0C
#343090000000
1!
1*
b110 6
19
1>
1C
b110 G
#343100000000
0!
0*
09
0>
0C
#343110000000
1!
1*
b111 6
19
1>
1C
b111 G
#343120000000
0!
0*
09
0>
0C
#343130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#343140000000
0!
0*
09
0>
0C
#343150000000
1!
1*
b1 6
19
1>
1C
b1 G
#343160000000
0!
0*
09
0>
0C
#343170000000
1!
1*
b10 6
19
1>
1C
b10 G
#343180000000
0!
0*
09
0>
0C
#343190000000
1!
1*
b11 6
19
1>
1C
b11 G
#343200000000
0!
0*
09
0>
0C
#343210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#343220000000
0!
0*
09
0>
0C
#343230000000
1!
1*
b101 6
19
1>
1C
b101 G
#343240000000
0!
0*
09
0>
0C
#343250000000
1!
1*
b110 6
19
1>
1C
b110 G
#343260000000
0!
0*
09
0>
0C
#343270000000
1!
1*
b111 6
19
1>
1C
b111 G
#343280000000
0!
0*
09
0>
0C
#343290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#343300000000
0!
0*
09
0>
0C
#343310000000
1!
1*
b1 6
19
1>
1C
b1 G
#343320000000
0!
0*
09
0>
0C
#343330000000
1!
1*
b10 6
19
1>
1C
b10 G
#343340000000
0!
0*
09
0>
0C
#343350000000
1!
1*
b11 6
19
1>
1C
b11 G
#343360000000
0!
0*
09
0>
0C
#343370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#343380000000
0!
0*
09
0>
0C
#343390000000
1!
1*
b101 6
19
1>
1C
b101 G
#343400000000
0!
0*
09
0>
0C
#343410000000
1!
1*
b110 6
19
1>
1C
b110 G
#343420000000
0!
0*
09
0>
0C
#343430000000
1!
1*
b111 6
19
1>
1C
b111 G
#343440000000
0!
1"
0*
1+
09
1:
0>
0C
#343450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#343460000000
0!
0*
09
0>
0C
#343470000000
1!
1*
b1 6
19
1>
1C
b1 G
#343480000000
0!
0*
09
0>
0C
#343490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#343500000000
0!
0*
09
0>
0C
#343510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#343520000000
0!
0*
09
0>
0C
#343530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#343540000000
0!
0*
09
0>
0C
#343550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#343560000000
0!
0#
0*
0,
09
0>
0?
0C
#343570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#343580000000
0!
0*
09
0>
0C
#343590000000
1!
1*
19
1>
1C
#343600000000
0!
0*
09
0>
0C
#343610000000
1!
1*
19
1>
1C
#343620000000
0!
0*
09
0>
0C
#343630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#343640000000
0!
0*
09
0>
0C
#343650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#343660000000
0!
0*
09
0>
0C
#343670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#343680000000
0!
0*
09
0>
0C
#343690000000
1!
1*
b10 6
19
1>
1C
b10 G
#343700000000
0!
0*
09
0>
0C
#343710000000
1!
1*
b11 6
19
1>
1C
b11 G
#343720000000
0!
0*
09
0>
0C
#343730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#343740000000
0!
0*
09
0>
0C
#343750000000
1!
1*
b101 6
19
1>
1C
b101 G
#343760000000
0!
0*
09
0>
0C
#343770000000
1!
1*
b110 6
19
1>
1C
b110 G
#343780000000
0!
0*
09
0>
0C
#343790000000
1!
1*
b111 6
19
1>
1C
b111 G
#343800000000
0!
0*
09
0>
0C
#343810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#343820000000
0!
0*
09
0>
0C
#343830000000
1!
1*
b1 6
19
1>
1C
b1 G
#343840000000
0!
0*
09
0>
0C
#343850000000
1!
1*
b10 6
19
1>
1C
b10 G
#343860000000
0!
0*
09
0>
0C
#343870000000
1!
1*
b11 6
19
1>
1C
b11 G
#343880000000
0!
0*
09
0>
0C
#343890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#343900000000
0!
0*
09
0>
0C
#343910000000
1!
1*
b101 6
19
1>
1C
b101 G
#343920000000
0!
0*
09
0>
0C
#343930000000
1!
1*
b110 6
19
1>
1C
b110 G
#343940000000
0!
0*
09
0>
0C
#343950000000
1!
1*
b111 6
19
1>
1C
b111 G
#343960000000
0!
0*
09
0>
0C
#343970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#343980000000
0!
0*
09
0>
0C
#343990000000
1!
1*
b1 6
19
1>
1C
b1 G
#344000000000
0!
0*
09
0>
0C
#344010000000
1!
1*
b10 6
19
1>
1C
b10 G
#344020000000
0!
0*
09
0>
0C
#344030000000
1!
1*
b11 6
19
1>
1C
b11 G
#344040000000
0!
0*
09
0>
0C
#344050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#344060000000
0!
0*
09
0>
0C
#344070000000
1!
1*
b101 6
19
1>
1C
b101 G
#344080000000
0!
0*
09
0>
0C
#344090000000
1!
1*
b110 6
19
1>
1C
b110 G
#344100000000
0!
0*
09
0>
0C
#344110000000
1!
1*
b111 6
19
1>
1C
b111 G
#344120000000
0!
1"
0*
1+
09
1:
0>
0C
#344130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#344140000000
0!
0*
09
0>
0C
#344150000000
1!
1*
b1 6
19
1>
1C
b1 G
#344160000000
0!
0*
09
0>
0C
#344170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#344180000000
0!
0*
09
0>
0C
#344190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#344200000000
0!
0*
09
0>
0C
#344210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#344220000000
0!
0*
09
0>
0C
#344230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#344240000000
0!
0#
0*
0,
09
0>
0?
0C
#344250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#344260000000
0!
0*
09
0>
0C
#344270000000
1!
1*
19
1>
1C
#344280000000
0!
0*
09
0>
0C
#344290000000
1!
1*
19
1>
1C
#344300000000
0!
0*
09
0>
0C
#344310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#344320000000
0!
0*
09
0>
0C
#344330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#344340000000
0!
0*
09
0>
0C
#344350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#344360000000
0!
0*
09
0>
0C
#344370000000
1!
1*
b10 6
19
1>
1C
b10 G
#344380000000
0!
0*
09
0>
0C
#344390000000
1!
1*
b11 6
19
1>
1C
b11 G
#344400000000
0!
0*
09
0>
0C
#344410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#344420000000
0!
0*
09
0>
0C
#344430000000
1!
1*
b101 6
19
1>
1C
b101 G
#344440000000
0!
0*
09
0>
0C
#344450000000
1!
1*
b110 6
19
1>
1C
b110 G
#344460000000
0!
0*
09
0>
0C
#344470000000
1!
1*
b111 6
19
1>
1C
b111 G
#344480000000
0!
0*
09
0>
0C
#344490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#344500000000
0!
0*
09
0>
0C
#344510000000
1!
1*
b1 6
19
1>
1C
b1 G
#344520000000
0!
0*
09
0>
0C
#344530000000
1!
1*
b10 6
19
1>
1C
b10 G
#344540000000
0!
0*
09
0>
0C
#344550000000
1!
1*
b11 6
19
1>
1C
b11 G
#344560000000
0!
0*
09
0>
0C
#344570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#344580000000
0!
0*
09
0>
0C
#344590000000
1!
1*
b101 6
19
1>
1C
b101 G
#344600000000
0!
0*
09
0>
0C
#344610000000
1!
1*
b110 6
19
1>
1C
b110 G
#344620000000
0!
0*
09
0>
0C
#344630000000
1!
1*
b111 6
19
1>
1C
b111 G
#344640000000
0!
0*
09
0>
0C
#344650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#344660000000
0!
0*
09
0>
0C
#344670000000
1!
1*
b1 6
19
1>
1C
b1 G
#344680000000
0!
0*
09
0>
0C
#344690000000
1!
1*
b10 6
19
1>
1C
b10 G
#344700000000
0!
0*
09
0>
0C
#344710000000
1!
1*
b11 6
19
1>
1C
b11 G
#344720000000
0!
0*
09
0>
0C
#344730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#344740000000
0!
0*
09
0>
0C
#344750000000
1!
1*
b101 6
19
1>
1C
b101 G
#344760000000
0!
0*
09
0>
0C
#344770000000
1!
1*
b110 6
19
1>
1C
b110 G
#344780000000
0!
0*
09
0>
0C
#344790000000
1!
1*
b111 6
19
1>
1C
b111 G
#344800000000
0!
1"
0*
1+
09
1:
0>
0C
#344810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#344820000000
0!
0*
09
0>
0C
#344830000000
1!
1*
b1 6
19
1>
1C
b1 G
#344840000000
0!
0*
09
0>
0C
#344850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#344860000000
0!
0*
09
0>
0C
#344870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#344880000000
0!
0*
09
0>
0C
#344890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#344900000000
0!
0*
09
0>
0C
#344910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#344920000000
0!
0#
0*
0,
09
0>
0?
0C
#344930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#344940000000
0!
0*
09
0>
0C
#344950000000
1!
1*
19
1>
1C
#344960000000
0!
0*
09
0>
0C
#344970000000
1!
1*
19
1>
1C
#344980000000
0!
0*
09
0>
0C
#344990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#345000000000
0!
0*
09
0>
0C
#345010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#345020000000
0!
0*
09
0>
0C
#345030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#345040000000
0!
0*
09
0>
0C
#345050000000
1!
1*
b10 6
19
1>
1C
b10 G
#345060000000
0!
0*
09
0>
0C
#345070000000
1!
1*
b11 6
19
1>
1C
b11 G
#345080000000
0!
0*
09
0>
0C
#345090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#345100000000
0!
0*
09
0>
0C
#345110000000
1!
1*
b101 6
19
1>
1C
b101 G
#345120000000
0!
0*
09
0>
0C
#345130000000
1!
1*
b110 6
19
1>
1C
b110 G
#345140000000
0!
0*
09
0>
0C
#345150000000
1!
1*
b111 6
19
1>
1C
b111 G
#345160000000
0!
0*
09
0>
0C
#345170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#345180000000
0!
0*
09
0>
0C
#345190000000
1!
1*
b1 6
19
1>
1C
b1 G
#345200000000
0!
0*
09
0>
0C
#345210000000
1!
1*
b10 6
19
1>
1C
b10 G
#345220000000
0!
0*
09
0>
0C
#345230000000
1!
1*
b11 6
19
1>
1C
b11 G
#345240000000
0!
0*
09
0>
0C
#345250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#345260000000
0!
0*
09
0>
0C
#345270000000
1!
1*
b101 6
19
1>
1C
b101 G
#345280000000
0!
0*
09
0>
0C
#345290000000
1!
1*
b110 6
19
1>
1C
b110 G
#345300000000
0!
0*
09
0>
0C
#345310000000
1!
1*
b111 6
19
1>
1C
b111 G
#345320000000
0!
0*
09
0>
0C
#345330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#345340000000
0!
0*
09
0>
0C
#345350000000
1!
1*
b1 6
19
1>
1C
b1 G
#345360000000
0!
0*
09
0>
0C
#345370000000
1!
1*
b10 6
19
1>
1C
b10 G
#345380000000
0!
0*
09
0>
0C
#345390000000
1!
1*
b11 6
19
1>
1C
b11 G
#345400000000
0!
0*
09
0>
0C
#345410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#345420000000
0!
0*
09
0>
0C
#345430000000
1!
1*
b101 6
19
1>
1C
b101 G
#345440000000
0!
0*
09
0>
0C
#345450000000
1!
1*
b110 6
19
1>
1C
b110 G
#345460000000
0!
0*
09
0>
0C
#345470000000
1!
1*
b111 6
19
1>
1C
b111 G
#345480000000
0!
1"
0*
1+
09
1:
0>
0C
#345490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#345500000000
0!
0*
09
0>
0C
#345510000000
1!
1*
b1 6
19
1>
1C
b1 G
#345520000000
0!
0*
09
0>
0C
#345530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#345540000000
0!
0*
09
0>
0C
#345550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#345560000000
0!
0*
09
0>
0C
#345570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#345580000000
0!
0*
09
0>
0C
#345590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#345600000000
0!
0#
0*
0,
09
0>
0?
0C
#345610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#345620000000
0!
0*
09
0>
0C
#345630000000
1!
1*
19
1>
1C
#345640000000
0!
0*
09
0>
0C
#345650000000
1!
1*
19
1>
1C
#345660000000
0!
0*
09
0>
0C
#345670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#345680000000
0!
0*
09
0>
0C
#345690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#345700000000
0!
0*
09
0>
0C
#345710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#345720000000
0!
0*
09
0>
0C
#345730000000
1!
1*
b10 6
19
1>
1C
b10 G
#345740000000
0!
0*
09
0>
0C
#345750000000
1!
1*
b11 6
19
1>
1C
b11 G
#345760000000
0!
0*
09
0>
0C
#345770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#345780000000
0!
0*
09
0>
0C
#345790000000
1!
1*
b101 6
19
1>
1C
b101 G
#345800000000
0!
0*
09
0>
0C
#345810000000
1!
1*
b110 6
19
1>
1C
b110 G
#345820000000
0!
0*
09
0>
0C
#345830000000
1!
1*
b111 6
19
1>
1C
b111 G
#345840000000
0!
0*
09
0>
0C
#345850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#345860000000
0!
0*
09
0>
0C
#345870000000
1!
1*
b1 6
19
1>
1C
b1 G
#345880000000
0!
0*
09
0>
0C
#345890000000
1!
1*
b10 6
19
1>
1C
b10 G
#345900000000
0!
0*
09
0>
0C
#345910000000
1!
1*
b11 6
19
1>
1C
b11 G
#345920000000
0!
0*
09
0>
0C
#345930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#345940000000
0!
0*
09
0>
0C
#345950000000
1!
1*
b101 6
19
1>
1C
b101 G
#345960000000
0!
0*
09
0>
0C
#345970000000
1!
1*
b110 6
19
1>
1C
b110 G
#345980000000
0!
0*
09
0>
0C
#345990000000
1!
1*
b111 6
19
1>
1C
b111 G
#346000000000
0!
0*
09
0>
0C
#346010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#346020000000
0!
0*
09
0>
0C
#346030000000
1!
1*
b1 6
19
1>
1C
b1 G
#346040000000
0!
0*
09
0>
0C
#346050000000
1!
1*
b10 6
19
1>
1C
b10 G
#346060000000
0!
0*
09
0>
0C
#346070000000
1!
1*
b11 6
19
1>
1C
b11 G
#346080000000
0!
0*
09
0>
0C
#346090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#346100000000
0!
0*
09
0>
0C
#346110000000
1!
1*
b101 6
19
1>
1C
b101 G
#346120000000
0!
0*
09
0>
0C
#346130000000
1!
1*
b110 6
19
1>
1C
b110 G
#346140000000
0!
0*
09
0>
0C
#346150000000
1!
1*
b111 6
19
1>
1C
b111 G
#346160000000
0!
1"
0*
1+
09
1:
0>
0C
#346170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#346180000000
0!
0*
09
0>
0C
#346190000000
1!
1*
b1 6
19
1>
1C
b1 G
#346200000000
0!
0*
09
0>
0C
#346210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#346220000000
0!
0*
09
0>
0C
#346230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#346240000000
0!
0*
09
0>
0C
#346250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#346260000000
0!
0*
09
0>
0C
#346270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#346280000000
0!
0#
0*
0,
09
0>
0?
0C
#346290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#346300000000
0!
0*
09
0>
0C
#346310000000
1!
1*
19
1>
1C
#346320000000
0!
0*
09
0>
0C
#346330000000
1!
1*
19
1>
1C
#346340000000
0!
0*
09
0>
0C
#346350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#346360000000
0!
0*
09
0>
0C
#346370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#346380000000
0!
0*
09
0>
0C
#346390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#346400000000
0!
0*
09
0>
0C
#346410000000
1!
1*
b10 6
19
1>
1C
b10 G
#346420000000
0!
0*
09
0>
0C
#346430000000
1!
1*
b11 6
19
1>
1C
b11 G
#346440000000
0!
0*
09
0>
0C
#346450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#346460000000
0!
0*
09
0>
0C
#346470000000
1!
1*
b101 6
19
1>
1C
b101 G
#346480000000
0!
0*
09
0>
0C
#346490000000
1!
1*
b110 6
19
1>
1C
b110 G
#346500000000
0!
0*
09
0>
0C
#346510000000
1!
1*
b111 6
19
1>
1C
b111 G
#346520000000
0!
0*
09
0>
0C
#346530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#346540000000
0!
0*
09
0>
0C
#346550000000
1!
1*
b1 6
19
1>
1C
b1 G
#346560000000
0!
0*
09
0>
0C
#346570000000
1!
1*
b10 6
19
1>
1C
b10 G
#346580000000
0!
0*
09
0>
0C
#346590000000
1!
1*
b11 6
19
1>
1C
b11 G
#346600000000
0!
0*
09
0>
0C
#346610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#346620000000
0!
0*
09
0>
0C
#346630000000
1!
1*
b101 6
19
1>
1C
b101 G
#346640000000
0!
0*
09
0>
0C
#346650000000
1!
1*
b110 6
19
1>
1C
b110 G
#346660000000
0!
0*
09
0>
0C
#346670000000
1!
1*
b111 6
19
1>
1C
b111 G
#346680000000
0!
0*
09
0>
0C
#346690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#346700000000
0!
0*
09
0>
0C
#346710000000
1!
1*
b1 6
19
1>
1C
b1 G
#346720000000
0!
0*
09
0>
0C
#346730000000
1!
1*
b10 6
19
1>
1C
b10 G
#346740000000
0!
0*
09
0>
0C
#346750000000
1!
1*
b11 6
19
1>
1C
b11 G
#346760000000
0!
0*
09
0>
0C
#346770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#346780000000
0!
0*
09
0>
0C
#346790000000
1!
1*
b101 6
19
1>
1C
b101 G
#346800000000
0!
0*
09
0>
0C
#346810000000
1!
1*
b110 6
19
1>
1C
b110 G
#346820000000
0!
0*
09
0>
0C
#346830000000
1!
1*
b111 6
19
1>
1C
b111 G
#346840000000
0!
1"
0*
1+
09
1:
0>
0C
#346850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#346860000000
0!
0*
09
0>
0C
#346870000000
1!
1*
b1 6
19
1>
1C
b1 G
#346880000000
0!
0*
09
0>
0C
#346890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#346900000000
0!
0*
09
0>
0C
#346910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#346920000000
0!
0*
09
0>
0C
#346930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#346940000000
0!
0*
09
0>
0C
#346950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#346960000000
0!
0#
0*
0,
09
0>
0?
0C
#346970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#346980000000
0!
0*
09
0>
0C
#346990000000
1!
1*
19
1>
1C
#347000000000
0!
0*
09
0>
0C
#347010000000
1!
1*
19
1>
1C
#347020000000
0!
0*
09
0>
0C
#347030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#347040000000
0!
0*
09
0>
0C
#347050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#347060000000
0!
0*
09
0>
0C
#347070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#347080000000
0!
0*
09
0>
0C
#347090000000
1!
1*
b10 6
19
1>
1C
b10 G
#347100000000
0!
0*
09
0>
0C
#347110000000
1!
1*
b11 6
19
1>
1C
b11 G
#347120000000
0!
0*
09
0>
0C
#347130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#347140000000
0!
0*
09
0>
0C
#347150000000
1!
1*
b101 6
19
1>
1C
b101 G
#347160000000
0!
0*
09
0>
0C
#347170000000
1!
1*
b110 6
19
1>
1C
b110 G
#347180000000
0!
0*
09
0>
0C
#347190000000
1!
1*
b111 6
19
1>
1C
b111 G
#347200000000
0!
0*
09
0>
0C
#347210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#347220000000
0!
0*
09
0>
0C
#347230000000
1!
1*
b1 6
19
1>
1C
b1 G
#347240000000
0!
0*
09
0>
0C
#347250000000
1!
1*
b10 6
19
1>
1C
b10 G
#347260000000
0!
0*
09
0>
0C
#347270000000
1!
1*
b11 6
19
1>
1C
b11 G
#347280000000
0!
0*
09
0>
0C
#347290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#347300000000
0!
0*
09
0>
0C
#347310000000
1!
1*
b101 6
19
1>
1C
b101 G
#347320000000
0!
0*
09
0>
0C
#347330000000
1!
1*
b110 6
19
1>
1C
b110 G
#347340000000
0!
0*
09
0>
0C
#347350000000
1!
1*
b111 6
19
1>
1C
b111 G
#347360000000
0!
0*
09
0>
0C
#347370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#347380000000
0!
0*
09
0>
0C
#347390000000
1!
1*
b1 6
19
1>
1C
b1 G
#347400000000
0!
0*
09
0>
0C
#347410000000
1!
1*
b10 6
19
1>
1C
b10 G
#347420000000
0!
0*
09
0>
0C
#347430000000
1!
1*
b11 6
19
1>
1C
b11 G
#347440000000
0!
0*
09
0>
0C
#347450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#347460000000
0!
0*
09
0>
0C
#347470000000
1!
1*
b101 6
19
1>
1C
b101 G
#347480000000
0!
0*
09
0>
0C
#347490000000
1!
1*
b110 6
19
1>
1C
b110 G
#347500000000
0!
0*
09
0>
0C
#347510000000
1!
1*
b111 6
19
1>
1C
b111 G
#347520000000
0!
1"
0*
1+
09
1:
0>
0C
#347530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#347540000000
0!
0*
09
0>
0C
#347550000000
1!
1*
b1 6
19
1>
1C
b1 G
#347560000000
0!
0*
09
0>
0C
#347570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#347580000000
0!
0*
09
0>
0C
#347590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#347600000000
0!
0*
09
0>
0C
#347610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#347620000000
0!
0*
09
0>
0C
#347630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#347640000000
0!
0#
0*
0,
09
0>
0?
0C
#347650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#347660000000
0!
0*
09
0>
0C
#347670000000
1!
1*
19
1>
1C
#347680000000
0!
0*
09
0>
0C
#347690000000
1!
1*
19
1>
1C
#347700000000
0!
0*
09
0>
0C
#347710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#347720000000
0!
0*
09
0>
0C
#347730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#347740000000
0!
0*
09
0>
0C
#347750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#347760000000
0!
0*
09
0>
0C
#347770000000
1!
1*
b10 6
19
1>
1C
b10 G
#347780000000
0!
0*
09
0>
0C
#347790000000
1!
1*
b11 6
19
1>
1C
b11 G
#347800000000
0!
0*
09
0>
0C
#347810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#347820000000
0!
0*
09
0>
0C
#347830000000
1!
1*
b101 6
19
1>
1C
b101 G
#347840000000
0!
0*
09
0>
0C
#347850000000
1!
1*
b110 6
19
1>
1C
b110 G
#347860000000
0!
0*
09
0>
0C
#347870000000
1!
1*
b111 6
19
1>
1C
b111 G
#347880000000
0!
0*
09
0>
0C
#347890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#347900000000
0!
0*
09
0>
0C
#347910000000
1!
1*
b1 6
19
1>
1C
b1 G
#347920000000
0!
0*
09
0>
0C
#347930000000
1!
1*
b10 6
19
1>
1C
b10 G
#347940000000
0!
0*
09
0>
0C
#347950000000
1!
1*
b11 6
19
1>
1C
b11 G
#347960000000
0!
0*
09
0>
0C
#347970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#347980000000
0!
0*
09
0>
0C
#347990000000
1!
1*
b101 6
19
1>
1C
b101 G
#348000000000
0!
0*
09
0>
0C
#348010000000
1!
1*
b110 6
19
1>
1C
b110 G
#348020000000
0!
0*
09
0>
0C
#348030000000
1!
1*
b111 6
19
1>
1C
b111 G
#348040000000
0!
0*
09
0>
0C
#348050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#348060000000
0!
0*
09
0>
0C
#348070000000
1!
1*
b1 6
19
1>
1C
b1 G
#348080000000
0!
0*
09
0>
0C
#348090000000
1!
1*
b10 6
19
1>
1C
b10 G
#348100000000
0!
0*
09
0>
0C
#348110000000
1!
1*
b11 6
19
1>
1C
b11 G
#348120000000
0!
0*
09
0>
0C
#348130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#348140000000
0!
0*
09
0>
0C
#348150000000
1!
1*
b101 6
19
1>
1C
b101 G
#348160000000
0!
0*
09
0>
0C
#348170000000
1!
1*
b110 6
19
1>
1C
b110 G
#348180000000
0!
0*
09
0>
0C
#348190000000
1!
1*
b111 6
19
1>
1C
b111 G
#348200000000
0!
1"
0*
1+
09
1:
0>
0C
#348210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#348220000000
0!
0*
09
0>
0C
#348230000000
1!
1*
b1 6
19
1>
1C
b1 G
#348240000000
0!
0*
09
0>
0C
#348250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#348260000000
0!
0*
09
0>
0C
#348270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#348280000000
0!
0*
09
0>
0C
#348290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#348300000000
0!
0*
09
0>
0C
#348310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#348320000000
0!
0#
0*
0,
09
0>
0?
0C
#348330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#348340000000
0!
0*
09
0>
0C
#348350000000
1!
1*
19
1>
1C
#348360000000
0!
0*
09
0>
0C
#348370000000
1!
1*
19
1>
1C
#348380000000
0!
0*
09
0>
0C
#348390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#348400000000
0!
0*
09
0>
0C
#348410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#348420000000
0!
0*
09
0>
0C
#348430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#348440000000
0!
0*
09
0>
0C
#348450000000
1!
1*
b10 6
19
1>
1C
b10 G
#348460000000
0!
0*
09
0>
0C
#348470000000
1!
1*
b11 6
19
1>
1C
b11 G
#348480000000
0!
0*
09
0>
0C
#348490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#348500000000
0!
0*
09
0>
0C
#348510000000
1!
1*
b101 6
19
1>
1C
b101 G
#348520000000
0!
0*
09
0>
0C
#348530000000
1!
1*
b110 6
19
1>
1C
b110 G
#348540000000
0!
0*
09
0>
0C
#348550000000
1!
1*
b111 6
19
1>
1C
b111 G
#348560000000
0!
0*
09
0>
0C
#348570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#348580000000
0!
0*
09
0>
0C
#348590000000
1!
1*
b1 6
19
1>
1C
b1 G
#348600000000
0!
0*
09
0>
0C
#348610000000
1!
1*
b10 6
19
1>
1C
b10 G
#348620000000
0!
0*
09
0>
0C
#348630000000
1!
1*
b11 6
19
1>
1C
b11 G
#348640000000
0!
0*
09
0>
0C
#348650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#348660000000
0!
0*
09
0>
0C
#348670000000
1!
1*
b101 6
19
1>
1C
b101 G
#348680000000
0!
0*
09
0>
0C
#348690000000
1!
1*
b110 6
19
1>
1C
b110 G
#348700000000
0!
0*
09
0>
0C
#348710000000
1!
1*
b111 6
19
1>
1C
b111 G
#348720000000
0!
0*
09
0>
0C
#348730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#348740000000
0!
0*
09
0>
0C
#348750000000
1!
1*
b1 6
19
1>
1C
b1 G
#348760000000
0!
0*
09
0>
0C
#348770000000
1!
1*
b10 6
19
1>
1C
b10 G
#348780000000
0!
0*
09
0>
0C
#348790000000
1!
1*
b11 6
19
1>
1C
b11 G
#348800000000
0!
0*
09
0>
0C
#348810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#348820000000
0!
0*
09
0>
0C
#348830000000
1!
1*
b101 6
19
1>
1C
b101 G
#348840000000
0!
0*
09
0>
0C
#348850000000
1!
1*
b110 6
19
1>
1C
b110 G
#348860000000
0!
0*
09
0>
0C
#348870000000
1!
1*
b111 6
19
1>
1C
b111 G
#348880000000
0!
1"
0*
1+
09
1:
0>
0C
#348890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#348900000000
0!
0*
09
0>
0C
#348910000000
1!
1*
b1 6
19
1>
1C
b1 G
#348920000000
0!
0*
09
0>
0C
#348930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#348940000000
0!
0*
09
0>
0C
#348950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#348960000000
0!
0*
09
0>
0C
#348970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#348980000000
0!
0*
09
0>
0C
#348990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#349000000000
0!
0#
0*
0,
09
0>
0?
0C
#349010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#349020000000
0!
0*
09
0>
0C
#349030000000
1!
1*
19
1>
1C
#349040000000
0!
0*
09
0>
0C
#349050000000
1!
1*
19
1>
1C
#349060000000
0!
0*
09
0>
0C
#349070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#349080000000
0!
0*
09
0>
0C
#349090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#349100000000
0!
0*
09
0>
0C
#349110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#349120000000
0!
0*
09
0>
0C
#349130000000
1!
1*
b10 6
19
1>
1C
b10 G
#349140000000
0!
0*
09
0>
0C
#349150000000
1!
1*
b11 6
19
1>
1C
b11 G
#349160000000
0!
0*
09
0>
0C
#349170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#349180000000
0!
0*
09
0>
0C
#349190000000
1!
1*
b101 6
19
1>
1C
b101 G
#349200000000
0!
0*
09
0>
0C
#349210000000
1!
1*
b110 6
19
1>
1C
b110 G
#349220000000
0!
0*
09
0>
0C
#349230000000
1!
1*
b111 6
19
1>
1C
b111 G
#349240000000
0!
0*
09
0>
0C
#349250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#349260000000
0!
0*
09
0>
0C
#349270000000
1!
1*
b1 6
19
1>
1C
b1 G
#349280000000
0!
0*
09
0>
0C
#349290000000
1!
1*
b10 6
19
1>
1C
b10 G
#349300000000
0!
0*
09
0>
0C
#349310000000
1!
1*
b11 6
19
1>
1C
b11 G
#349320000000
0!
0*
09
0>
0C
#349330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#349340000000
0!
0*
09
0>
0C
#349350000000
1!
1*
b101 6
19
1>
1C
b101 G
#349360000000
0!
0*
09
0>
0C
#349370000000
1!
1*
b110 6
19
1>
1C
b110 G
#349380000000
0!
0*
09
0>
0C
#349390000000
1!
1*
b111 6
19
1>
1C
b111 G
#349400000000
0!
0*
09
0>
0C
#349410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#349420000000
0!
0*
09
0>
0C
#349430000000
1!
1*
b1 6
19
1>
1C
b1 G
#349440000000
0!
0*
09
0>
0C
#349450000000
1!
1*
b10 6
19
1>
1C
b10 G
#349460000000
0!
0*
09
0>
0C
#349470000000
1!
1*
b11 6
19
1>
1C
b11 G
#349480000000
0!
0*
09
0>
0C
#349490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#349500000000
0!
0*
09
0>
0C
#349510000000
1!
1*
b101 6
19
1>
1C
b101 G
#349520000000
0!
0*
09
0>
0C
#349530000000
1!
1*
b110 6
19
1>
1C
b110 G
#349540000000
0!
0*
09
0>
0C
#349550000000
1!
1*
b111 6
19
1>
1C
b111 G
#349560000000
0!
1"
0*
1+
09
1:
0>
0C
#349570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#349580000000
0!
0*
09
0>
0C
#349590000000
1!
1*
b1 6
19
1>
1C
b1 G
#349600000000
0!
0*
09
0>
0C
#349610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#349620000000
0!
0*
09
0>
0C
#349630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#349640000000
0!
0*
09
0>
0C
#349650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#349660000000
0!
0*
09
0>
0C
#349670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#349680000000
0!
0#
0*
0,
09
0>
0?
0C
#349690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#349700000000
0!
0*
09
0>
0C
#349710000000
1!
1*
19
1>
1C
#349720000000
0!
0*
09
0>
0C
#349730000000
1!
1*
19
1>
1C
#349740000000
0!
0*
09
0>
0C
#349750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#349760000000
0!
0*
09
0>
0C
#349770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#349780000000
0!
0*
09
0>
0C
#349790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#349800000000
0!
0*
09
0>
0C
#349810000000
1!
1*
b10 6
19
1>
1C
b10 G
#349820000000
0!
0*
09
0>
0C
#349830000000
1!
1*
b11 6
19
1>
1C
b11 G
#349840000000
0!
0*
09
0>
0C
#349850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#349860000000
0!
0*
09
0>
0C
#349870000000
1!
1*
b101 6
19
1>
1C
b101 G
#349880000000
0!
0*
09
0>
0C
#349890000000
1!
1*
b110 6
19
1>
1C
b110 G
#349900000000
0!
0*
09
0>
0C
#349910000000
1!
1*
b111 6
19
1>
1C
b111 G
#349920000000
0!
0*
09
0>
0C
#349930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#349940000000
0!
0*
09
0>
0C
#349950000000
1!
1*
b1 6
19
1>
1C
b1 G
#349960000000
0!
0*
09
0>
0C
#349970000000
1!
1*
b10 6
19
1>
1C
b10 G
#349980000000
0!
0*
09
0>
0C
#349990000000
1!
1*
b11 6
19
1>
1C
b11 G
#350000000000
0!
0*
09
0>
0C
#350010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#350020000000
0!
0*
09
0>
0C
#350030000000
1!
1*
b101 6
19
1>
1C
b101 G
#350040000000
0!
0*
09
0>
0C
#350050000000
1!
1*
b110 6
19
1>
1C
b110 G
#350060000000
0!
0*
09
0>
0C
#350070000000
1!
1*
b111 6
19
1>
1C
b111 G
#350080000000
0!
0*
09
0>
0C
#350090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#350100000000
0!
0*
09
0>
0C
#350110000000
1!
1*
b1 6
19
1>
1C
b1 G
#350120000000
0!
0*
09
0>
0C
#350130000000
1!
1*
b10 6
19
1>
1C
b10 G
#350140000000
0!
0*
09
0>
0C
#350150000000
1!
1*
b11 6
19
1>
1C
b11 G
#350160000000
0!
0*
09
0>
0C
#350170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#350180000000
0!
0*
09
0>
0C
#350190000000
1!
1*
b101 6
19
1>
1C
b101 G
#350200000000
0!
0*
09
0>
0C
#350210000000
1!
1*
b110 6
19
1>
1C
b110 G
#350220000000
0!
0*
09
0>
0C
#350230000000
1!
1*
b111 6
19
1>
1C
b111 G
#350240000000
0!
1"
0*
1+
09
1:
0>
0C
#350250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#350260000000
0!
0*
09
0>
0C
#350270000000
1!
1*
b1 6
19
1>
1C
b1 G
#350280000000
0!
0*
09
0>
0C
#350290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#350300000000
0!
0*
09
0>
0C
#350310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#350320000000
0!
0*
09
0>
0C
#350330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#350340000000
0!
0*
09
0>
0C
#350350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#350360000000
0!
0#
0*
0,
09
0>
0?
0C
#350370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#350380000000
0!
0*
09
0>
0C
#350390000000
1!
1*
19
1>
1C
#350400000000
0!
0*
09
0>
0C
#350410000000
1!
1*
19
1>
1C
#350420000000
0!
0*
09
0>
0C
#350430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#350440000000
0!
0*
09
0>
0C
#350450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#350460000000
0!
0*
09
0>
0C
#350470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#350480000000
0!
0*
09
0>
0C
#350490000000
1!
1*
b10 6
19
1>
1C
b10 G
#350500000000
0!
0*
09
0>
0C
#350510000000
1!
1*
b11 6
19
1>
1C
b11 G
#350520000000
0!
0*
09
0>
0C
#350530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#350540000000
0!
0*
09
0>
0C
#350550000000
1!
1*
b101 6
19
1>
1C
b101 G
#350560000000
0!
0*
09
0>
0C
#350570000000
1!
1*
b110 6
19
1>
1C
b110 G
#350580000000
0!
0*
09
0>
0C
#350590000000
1!
1*
b111 6
19
1>
1C
b111 G
#350600000000
0!
0*
09
0>
0C
#350610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#350620000000
0!
0*
09
0>
0C
#350630000000
1!
1*
b1 6
19
1>
1C
b1 G
#350640000000
0!
0*
09
0>
0C
#350650000000
1!
1*
b10 6
19
1>
1C
b10 G
#350660000000
0!
0*
09
0>
0C
#350670000000
1!
1*
b11 6
19
1>
1C
b11 G
#350680000000
0!
0*
09
0>
0C
#350690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#350700000000
0!
0*
09
0>
0C
#350710000000
1!
1*
b101 6
19
1>
1C
b101 G
#350720000000
0!
0*
09
0>
0C
#350730000000
1!
1*
b110 6
19
1>
1C
b110 G
#350740000000
0!
0*
09
0>
0C
#350750000000
1!
1*
b111 6
19
1>
1C
b111 G
#350760000000
0!
0*
09
0>
0C
#350770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#350780000000
0!
0*
09
0>
0C
#350790000000
1!
1*
b1 6
19
1>
1C
b1 G
#350800000000
0!
0*
09
0>
0C
#350810000000
1!
1*
b10 6
19
1>
1C
b10 G
#350820000000
0!
0*
09
0>
0C
#350830000000
1!
1*
b11 6
19
1>
1C
b11 G
#350840000000
0!
0*
09
0>
0C
#350850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#350860000000
0!
0*
09
0>
0C
#350870000000
1!
1*
b101 6
19
1>
1C
b101 G
#350880000000
0!
0*
09
0>
0C
#350890000000
1!
1*
b110 6
19
1>
1C
b110 G
#350900000000
0!
0*
09
0>
0C
#350910000000
1!
1*
b111 6
19
1>
1C
b111 G
#350920000000
0!
1"
0*
1+
09
1:
0>
0C
#350930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#350940000000
0!
0*
09
0>
0C
#350950000000
1!
1*
b1 6
19
1>
1C
b1 G
#350960000000
0!
0*
09
0>
0C
#350970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#350980000000
0!
0*
09
0>
0C
#350990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#351000000000
0!
0*
09
0>
0C
#351010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#351020000000
0!
0*
09
0>
0C
#351030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#351040000000
0!
0#
0*
0,
09
0>
0?
0C
#351050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#351060000000
0!
0*
09
0>
0C
#351070000000
1!
1*
19
1>
1C
#351080000000
0!
0*
09
0>
0C
#351090000000
1!
1*
19
1>
1C
#351100000000
0!
0*
09
0>
0C
#351110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#351120000000
0!
0*
09
0>
0C
#351130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#351140000000
0!
0*
09
0>
0C
#351150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#351160000000
0!
0*
09
0>
0C
#351170000000
1!
1*
b10 6
19
1>
1C
b10 G
#351180000000
0!
0*
09
0>
0C
#351190000000
1!
1*
b11 6
19
1>
1C
b11 G
#351200000000
0!
0*
09
0>
0C
#351210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#351220000000
0!
0*
09
0>
0C
#351230000000
1!
1*
b101 6
19
1>
1C
b101 G
#351240000000
0!
0*
09
0>
0C
#351250000000
1!
1*
b110 6
19
1>
1C
b110 G
#351260000000
0!
0*
09
0>
0C
#351270000000
1!
1*
b111 6
19
1>
1C
b111 G
#351280000000
0!
0*
09
0>
0C
#351290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#351300000000
0!
0*
09
0>
0C
#351310000000
1!
1*
b1 6
19
1>
1C
b1 G
#351320000000
0!
0*
09
0>
0C
#351330000000
1!
1*
b10 6
19
1>
1C
b10 G
#351340000000
0!
0*
09
0>
0C
#351350000000
1!
1*
b11 6
19
1>
1C
b11 G
#351360000000
0!
0*
09
0>
0C
#351370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#351380000000
0!
0*
09
0>
0C
#351390000000
1!
1*
b101 6
19
1>
1C
b101 G
#351400000000
0!
0*
09
0>
0C
#351410000000
1!
1*
b110 6
19
1>
1C
b110 G
#351420000000
0!
0*
09
0>
0C
#351430000000
1!
1*
b111 6
19
1>
1C
b111 G
#351440000000
0!
0*
09
0>
0C
#351450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#351460000000
0!
0*
09
0>
0C
#351470000000
1!
1*
b1 6
19
1>
1C
b1 G
#351480000000
0!
0*
09
0>
0C
#351490000000
1!
1*
b10 6
19
1>
1C
b10 G
#351500000000
0!
0*
09
0>
0C
#351510000000
1!
1*
b11 6
19
1>
1C
b11 G
#351520000000
0!
0*
09
0>
0C
#351530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#351540000000
0!
0*
09
0>
0C
#351550000000
1!
1*
b101 6
19
1>
1C
b101 G
#351560000000
0!
0*
09
0>
0C
#351570000000
1!
1*
b110 6
19
1>
1C
b110 G
#351580000000
0!
0*
09
0>
0C
#351590000000
1!
1*
b111 6
19
1>
1C
b111 G
#351600000000
0!
1"
0*
1+
09
1:
0>
0C
#351610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#351620000000
0!
0*
09
0>
0C
#351630000000
1!
1*
b1 6
19
1>
1C
b1 G
#351640000000
0!
0*
09
0>
0C
#351650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#351660000000
0!
0*
09
0>
0C
#351670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#351680000000
0!
0*
09
0>
0C
#351690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#351700000000
0!
0*
09
0>
0C
#351710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#351720000000
0!
0#
0*
0,
09
0>
0?
0C
#351730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#351740000000
0!
0*
09
0>
0C
#351750000000
1!
1*
19
1>
1C
#351760000000
0!
0*
09
0>
0C
#351770000000
1!
1*
19
1>
1C
#351780000000
0!
0*
09
0>
0C
#351790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#351800000000
0!
0*
09
0>
0C
#351810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#351820000000
0!
0*
09
0>
0C
#351830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#351840000000
0!
0*
09
0>
0C
#351850000000
1!
1*
b10 6
19
1>
1C
b10 G
#351860000000
0!
0*
09
0>
0C
#351870000000
1!
1*
b11 6
19
1>
1C
b11 G
#351880000000
0!
0*
09
0>
0C
#351890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#351900000000
0!
0*
09
0>
0C
#351910000000
1!
1*
b101 6
19
1>
1C
b101 G
#351920000000
0!
0*
09
0>
0C
#351930000000
1!
1*
b110 6
19
1>
1C
b110 G
#351940000000
0!
0*
09
0>
0C
#351950000000
1!
1*
b111 6
19
1>
1C
b111 G
#351960000000
0!
0*
09
0>
0C
#351970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#351980000000
0!
0*
09
0>
0C
#351990000000
1!
1*
b1 6
19
1>
1C
b1 G
#352000000000
0!
0*
09
0>
0C
#352010000000
1!
1*
b10 6
19
1>
1C
b10 G
#352020000000
0!
0*
09
0>
0C
#352030000000
1!
1*
b11 6
19
1>
1C
b11 G
#352040000000
0!
0*
09
0>
0C
#352050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#352060000000
0!
0*
09
0>
0C
#352070000000
1!
1*
b101 6
19
1>
1C
b101 G
#352080000000
0!
0*
09
0>
0C
#352090000000
1!
1*
b110 6
19
1>
1C
b110 G
#352100000000
0!
0*
09
0>
0C
#352110000000
1!
1*
b111 6
19
1>
1C
b111 G
#352120000000
0!
0*
09
0>
0C
#352130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#352140000000
0!
0*
09
0>
0C
#352150000000
1!
1*
b1 6
19
1>
1C
b1 G
#352160000000
0!
0*
09
0>
0C
#352170000000
1!
1*
b10 6
19
1>
1C
b10 G
#352180000000
0!
0*
09
0>
0C
#352190000000
1!
1*
b11 6
19
1>
1C
b11 G
#352200000000
0!
0*
09
0>
0C
#352210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#352220000000
0!
0*
09
0>
0C
#352230000000
1!
1*
b101 6
19
1>
1C
b101 G
#352240000000
0!
0*
09
0>
0C
#352250000000
1!
1*
b110 6
19
1>
1C
b110 G
#352260000000
0!
0*
09
0>
0C
#352270000000
1!
1*
b111 6
19
1>
1C
b111 G
#352280000000
0!
1"
0*
1+
09
1:
0>
0C
#352290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#352300000000
0!
0*
09
0>
0C
#352310000000
1!
1*
b1 6
19
1>
1C
b1 G
#352320000000
0!
0*
09
0>
0C
#352330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#352340000000
0!
0*
09
0>
0C
#352350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#352360000000
0!
0*
09
0>
0C
#352370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#352380000000
0!
0*
09
0>
0C
#352390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#352400000000
0!
0#
0*
0,
09
0>
0?
0C
#352410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#352420000000
0!
0*
09
0>
0C
#352430000000
1!
1*
19
1>
1C
#352440000000
0!
0*
09
0>
0C
#352450000000
1!
1*
19
1>
1C
#352460000000
0!
0*
09
0>
0C
#352470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#352480000000
0!
0*
09
0>
0C
#352490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#352500000000
0!
0*
09
0>
0C
#352510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#352520000000
0!
0*
09
0>
0C
#352530000000
1!
1*
b10 6
19
1>
1C
b10 G
#352540000000
0!
0*
09
0>
0C
#352550000000
1!
1*
b11 6
19
1>
1C
b11 G
#352560000000
0!
0*
09
0>
0C
#352570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#352580000000
0!
0*
09
0>
0C
#352590000000
1!
1*
b101 6
19
1>
1C
b101 G
#352600000000
0!
0*
09
0>
0C
#352610000000
1!
1*
b110 6
19
1>
1C
b110 G
#352620000000
0!
0*
09
0>
0C
#352630000000
1!
1*
b111 6
19
1>
1C
b111 G
#352640000000
0!
0*
09
0>
0C
#352650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#352660000000
0!
0*
09
0>
0C
#352670000000
1!
1*
b1 6
19
1>
1C
b1 G
#352680000000
0!
0*
09
0>
0C
#352690000000
1!
1*
b10 6
19
1>
1C
b10 G
#352700000000
0!
0*
09
0>
0C
#352710000000
1!
1*
b11 6
19
1>
1C
b11 G
#352720000000
0!
0*
09
0>
0C
#352730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#352740000000
0!
0*
09
0>
0C
#352750000000
1!
1*
b101 6
19
1>
1C
b101 G
#352760000000
0!
0*
09
0>
0C
#352770000000
1!
1*
b110 6
19
1>
1C
b110 G
#352780000000
0!
0*
09
0>
0C
#352790000000
1!
1*
b111 6
19
1>
1C
b111 G
#352800000000
0!
0*
09
0>
0C
#352810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#352820000000
0!
0*
09
0>
0C
#352830000000
1!
1*
b1 6
19
1>
1C
b1 G
#352840000000
0!
0*
09
0>
0C
#352850000000
1!
1*
b10 6
19
1>
1C
b10 G
#352860000000
0!
0*
09
0>
0C
#352870000000
1!
1*
b11 6
19
1>
1C
b11 G
#352880000000
0!
0*
09
0>
0C
#352890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#352900000000
0!
0*
09
0>
0C
#352910000000
1!
1*
b101 6
19
1>
1C
b101 G
#352920000000
0!
0*
09
0>
0C
#352930000000
1!
1*
b110 6
19
1>
1C
b110 G
#352940000000
0!
0*
09
0>
0C
#352950000000
1!
1*
b111 6
19
1>
1C
b111 G
#352960000000
0!
1"
0*
1+
09
1:
0>
0C
#352970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#352980000000
0!
0*
09
0>
0C
#352990000000
1!
1*
b1 6
19
1>
1C
b1 G
#353000000000
0!
0*
09
0>
0C
#353010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#353020000000
0!
0*
09
0>
0C
#353030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#353040000000
0!
0*
09
0>
0C
#353050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#353060000000
0!
0*
09
0>
0C
#353070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#353080000000
0!
0#
0*
0,
09
0>
0?
0C
#353090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#353100000000
0!
0*
09
0>
0C
#353110000000
1!
1*
19
1>
1C
#353120000000
0!
0*
09
0>
0C
#353130000000
1!
1*
19
1>
1C
#353140000000
0!
0*
09
0>
0C
#353150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#353160000000
0!
0*
09
0>
0C
#353170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#353180000000
0!
0*
09
0>
0C
#353190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#353200000000
0!
0*
09
0>
0C
#353210000000
1!
1*
b10 6
19
1>
1C
b10 G
#353220000000
0!
0*
09
0>
0C
#353230000000
1!
1*
b11 6
19
1>
1C
b11 G
#353240000000
0!
0*
09
0>
0C
#353250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#353260000000
0!
0*
09
0>
0C
#353270000000
1!
1*
b101 6
19
1>
1C
b101 G
#353280000000
0!
0*
09
0>
0C
#353290000000
1!
1*
b110 6
19
1>
1C
b110 G
#353300000000
0!
0*
09
0>
0C
#353310000000
1!
1*
b111 6
19
1>
1C
b111 G
#353320000000
0!
0*
09
0>
0C
#353330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#353340000000
0!
0*
09
0>
0C
#353350000000
1!
1*
b1 6
19
1>
1C
b1 G
#353360000000
0!
0*
09
0>
0C
#353370000000
1!
1*
b10 6
19
1>
1C
b10 G
#353380000000
0!
0*
09
0>
0C
#353390000000
1!
1*
b11 6
19
1>
1C
b11 G
#353400000000
0!
0*
09
0>
0C
#353410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#353420000000
0!
0*
09
0>
0C
#353430000000
1!
1*
b101 6
19
1>
1C
b101 G
#353440000000
0!
0*
09
0>
0C
#353450000000
1!
1*
b110 6
19
1>
1C
b110 G
#353460000000
0!
0*
09
0>
0C
#353470000000
1!
1*
b111 6
19
1>
1C
b111 G
#353480000000
0!
0*
09
0>
0C
#353490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#353500000000
0!
0*
09
0>
0C
#353510000000
1!
1*
b1 6
19
1>
1C
b1 G
#353520000000
0!
0*
09
0>
0C
#353530000000
1!
1*
b10 6
19
1>
1C
b10 G
#353540000000
0!
0*
09
0>
0C
#353550000000
1!
1*
b11 6
19
1>
1C
b11 G
#353560000000
0!
0*
09
0>
0C
#353570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#353580000000
0!
0*
09
0>
0C
#353590000000
1!
1*
b101 6
19
1>
1C
b101 G
#353600000000
0!
0*
09
0>
0C
#353610000000
1!
1*
b110 6
19
1>
1C
b110 G
#353620000000
0!
0*
09
0>
0C
#353630000000
1!
1*
b111 6
19
1>
1C
b111 G
#353640000000
0!
1"
0*
1+
09
1:
0>
0C
#353650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#353660000000
0!
0*
09
0>
0C
#353670000000
1!
1*
b1 6
19
1>
1C
b1 G
#353680000000
0!
0*
09
0>
0C
#353690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#353700000000
0!
0*
09
0>
0C
#353710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#353720000000
0!
0*
09
0>
0C
#353730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#353740000000
0!
0*
09
0>
0C
#353750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#353760000000
0!
0#
0*
0,
09
0>
0?
0C
#353770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#353780000000
0!
0*
09
0>
0C
#353790000000
1!
1*
19
1>
1C
#353800000000
0!
0*
09
0>
0C
#353810000000
1!
1*
19
1>
1C
#353820000000
0!
0*
09
0>
0C
#353830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#353840000000
0!
0*
09
0>
0C
#353850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#353860000000
0!
0*
09
0>
0C
#353870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#353880000000
0!
0*
09
0>
0C
#353890000000
1!
1*
b10 6
19
1>
1C
b10 G
#353900000000
0!
0*
09
0>
0C
#353910000000
1!
1*
b11 6
19
1>
1C
b11 G
#353920000000
0!
0*
09
0>
0C
#353930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#353940000000
0!
0*
09
0>
0C
#353950000000
1!
1*
b101 6
19
1>
1C
b101 G
#353960000000
0!
0*
09
0>
0C
#353970000000
1!
1*
b110 6
19
1>
1C
b110 G
#353980000000
0!
0*
09
0>
0C
#353990000000
1!
1*
b111 6
19
1>
1C
b111 G
#354000000000
0!
0*
09
0>
0C
#354010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#354020000000
0!
0*
09
0>
0C
#354030000000
1!
1*
b1 6
19
1>
1C
b1 G
#354040000000
0!
0*
09
0>
0C
#354050000000
1!
1*
b10 6
19
1>
1C
b10 G
#354060000000
0!
0*
09
0>
0C
#354070000000
1!
1*
b11 6
19
1>
1C
b11 G
#354080000000
0!
0*
09
0>
0C
#354090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#354100000000
0!
0*
09
0>
0C
#354110000000
1!
1*
b101 6
19
1>
1C
b101 G
#354120000000
0!
0*
09
0>
0C
#354130000000
1!
1*
b110 6
19
1>
1C
b110 G
#354140000000
0!
0*
09
0>
0C
#354150000000
1!
1*
b111 6
19
1>
1C
b111 G
#354160000000
0!
0*
09
0>
0C
#354170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#354180000000
0!
0*
09
0>
0C
#354190000000
1!
1*
b1 6
19
1>
1C
b1 G
#354200000000
0!
0*
09
0>
0C
#354210000000
1!
1*
b10 6
19
1>
1C
b10 G
#354220000000
0!
0*
09
0>
0C
#354230000000
1!
1*
b11 6
19
1>
1C
b11 G
#354240000000
0!
0*
09
0>
0C
#354250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#354260000000
0!
0*
09
0>
0C
#354270000000
1!
1*
b101 6
19
1>
1C
b101 G
#354280000000
0!
0*
09
0>
0C
#354290000000
1!
1*
b110 6
19
1>
1C
b110 G
#354300000000
0!
0*
09
0>
0C
#354310000000
1!
1*
b111 6
19
1>
1C
b111 G
#354320000000
0!
1"
0*
1+
09
1:
0>
0C
#354330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#354340000000
0!
0*
09
0>
0C
#354350000000
1!
1*
b1 6
19
1>
1C
b1 G
#354360000000
0!
0*
09
0>
0C
#354370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#354380000000
0!
0*
09
0>
0C
#354390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#354400000000
0!
0*
09
0>
0C
#354410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#354420000000
0!
0*
09
0>
0C
#354430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#354440000000
0!
0#
0*
0,
09
0>
0?
0C
#354450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#354460000000
0!
0*
09
0>
0C
#354470000000
1!
1*
19
1>
1C
#354480000000
0!
0*
09
0>
0C
#354490000000
1!
1*
19
1>
1C
#354500000000
0!
0*
09
0>
0C
#354510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#354520000000
0!
0*
09
0>
0C
#354530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#354540000000
0!
0*
09
0>
0C
#354550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#354560000000
0!
0*
09
0>
0C
#354570000000
1!
1*
b10 6
19
1>
1C
b10 G
#354580000000
0!
0*
09
0>
0C
#354590000000
1!
1*
b11 6
19
1>
1C
b11 G
#354600000000
0!
0*
09
0>
0C
#354610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#354620000000
0!
0*
09
0>
0C
#354630000000
1!
1*
b101 6
19
1>
1C
b101 G
#354640000000
0!
0*
09
0>
0C
#354650000000
1!
1*
b110 6
19
1>
1C
b110 G
#354660000000
0!
0*
09
0>
0C
#354670000000
1!
1*
b111 6
19
1>
1C
b111 G
#354680000000
0!
0*
09
0>
0C
#354690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#354700000000
0!
0*
09
0>
0C
#354710000000
1!
1*
b1 6
19
1>
1C
b1 G
#354720000000
0!
0*
09
0>
0C
#354730000000
1!
1*
b10 6
19
1>
1C
b10 G
#354740000000
0!
0*
09
0>
0C
#354750000000
1!
1*
b11 6
19
1>
1C
b11 G
#354760000000
0!
0*
09
0>
0C
#354770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#354780000000
0!
0*
09
0>
0C
#354790000000
1!
1*
b101 6
19
1>
1C
b101 G
#354800000000
0!
0*
09
0>
0C
#354810000000
1!
1*
b110 6
19
1>
1C
b110 G
#354820000000
0!
0*
09
0>
0C
#354830000000
1!
1*
b111 6
19
1>
1C
b111 G
#354840000000
0!
0*
09
0>
0C
#354850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#354860000000
0!
0*
09
0>
0C
#354870000000
1!
1*
b1 6
19
1>
1C
b1 G
#354880000000
0!
0*
09
0>
0C
#354890000000
1!
1*
b10 6
19
1>
1C
b10 G
#354900000000
0!
0*
09
0>
0C
#354910000000
1!
1*
b11 6
19
1>
1C
b11 G
#354920000000
0!
0*
09
0>
0C
#354930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#354940000000
0!
0*
09
0>
0C
#354950000000
1!
1*
b101 6
19
1>
1C
b101 G
#354960000000
0!
0*
09
0>
0C
#354970000000
1!
1*
b110 6
19
1>
1C
b110 G
#354980000000
0!
0*
09
0>
0C
#354990000000
1!
1*
b111 6
19
1>
1C
b111 G
#355000000000
0!
1"
0*
1+
09
1:
0>
0C
#355010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#355020000000
0!
0*
09
0>
0C
#355030000000
1!
1*
b1 6
19
1>
1C
b1 G
#355040000000
0!
0*
09
0>
0C
#355050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#355060000000
0!
0*
09
0>
0C
#355070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#355080000000
0!
0*
09
0>
0C
#355090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#355100000000
0!
0*
09
0>
0C
#355110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#355120000000
0!
0#
0*
0,
09
0>
0?
0C
#355130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#355140000000
0!
0*
09
0>
0C
#355150000000
1!
1*
19
1>
1C
#355160000000
0!
0*
09
0>
0C
#355170000000
1!
1*
19
1>
1C
#355180000000
0!
0*
09
0>
0C
#355190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#355200000000
0!
0*
09
0>
0C
#355210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#355220000000
0!
0*
09
0>
0C
#355230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#355240000000
0!
0*
09
0>
0C
#355250000000
1!
1*
b10 6
19
1>
1C
b10 G
#355260000000
0!
0*
09
0>
0C
#355270000000
1!
1*
b11 6
19
1>
1C
b11 G
#355280000000
0!
0*
09
0>
0C
#355290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#355300000000
0!
0*
09
0>
0C
#355310000000
1!
1*
b101 6
19
1>
1C
b101 G
#355320000000
0!
0*
09
0>
0C
#355330000000
1!
1*
b110 6
19
1>
1C
b110 G
#355340000000
0!
0*
09
0>
0C
#355350000000
1!
1*
b111 6
19
1>
1C
b111 G
#355360000000
0!
0*
09
0>
0C
#355370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#355380000000
0!
0*
09
0>
0C
#355390000000
1!
1*
b1 6
19
1>
1C
b1 G
#355400000000
0!
0*
09
0>
0C
#355410000000
1!
1*
b10 6
19
1>
1C
b10 G
#355420000000
0!
0*
09
0>
0C
#355430000000
1!
1*
b11 6
19
1>
1C
b11 G
#355440000000
0!
0*
09
0>
0C
#355450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#355460000000
0!
0*
09
0>
0C
#355470000000
1!
1*
b101 6
19
1>
1C
b101 G
#355480000000
0!
0*
09
0>
0C
#355490000000
1!
1*
b110 6
19
1>
1C
b110 G
#355500000000
0!
0*
09
0>
0C
#355510000000
1!
1*
b111 6
19
1>
1C
b111 G
#355520000000
0!
0*
09
0>
0C
#355530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#355540000000
0!
0*
09
0>
0C
#355550000000
1!
1*
b1 6
19
1>
1C
b1 G
#355560000000
0!
0*
09
0>
0C
#355570000000
1!
1*
b10 6
19
1>
1C
b10 G
#355580000000
0!
0*
09
0>
0C
#355590000000
1!
1*
b11 6
19
1>
1C
b11 G
#355600000000
0!
0*
09
0>
0C
#355610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#355620000000
0!
0*
09
0>
0C
#355630000000
1!
1*
b101 6
19
1>
1C
b101 G
#355640000000
0!
0*
09
0>
0C
#355650000000
1!
1*
b110 6
19
1>
1C
b110 G
#355660000000
0!
0*
09
0>
0C
#355670000000
1!
1*
b111 6
19
1>
1C
b111 G
#355680000000
0!
1"
0*
1+
09
1:
0>
0C
#355690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#355700000000
0!
0*
09
0>
0C
#355710000000
1!
1*
b1 6
19
1>
1C
b1 G
#355720000000
0!
0*
09
0>
0C
#355730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#355740000000
0!
0*
09
0>
0C
#355750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#355760000000
0!
0*
09
0>
0C
#355770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#355780000000
0!
0*
09
0>
0C
#355790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#355800000000
0!
0#
0*
0,
09
0>
0?
0C
#355810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#355820000000
0!
0*
09
0>
0C
#355830000000
1!
1*
19
1>
1C
#355840000000
0!
0*
09
0>
0C
#355850000000
1!
1*
19
1>
1C
#355860000000
0!
0*
09
0>
0C
#355870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#355880000000
0!
0*
09
0>
0C
#355890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#355900000000
0!
0*
09
0>
0C
#355910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#355920000000
0!
0*
09
0>
0C
#355930000000
1!
1*
b10 6
19
1>
1C
b10 G
#355940000000
0!
0*
09
0>
0C
#355950000000
1!
1*
b11 6
19
1>
1C
b11 G
#355960000000
0!
0*
09
0>
0C
#355970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#355980000000
0!
0*
09
0>
0C
#355990000000
1!
1*
b101 6
19
1>
1C
b101 G
#356000000000
0!
0*
09
0>
0C
#356010000000
1!
1*
b110 6
19
1>
1C
b110 G
#356020000000
0!
0*
09
0>
0C
#356030000000
1!
1*
b111 6
19
1>
1C
b111 G
#356040000000
0!
0*
09
0>
0C
#356050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#356060000000
0!
0*
09
0>
0C
#356070000000
1!
1*
b1 6
19
1>
1C
b1 G
#356080000000
0!
0*
09
0>
0C
#356090000000
1!
1*
b10 6
19
1>
1C
b10 G
#356100000000
0!
0*
09
0>
0C
#356110000000
1!
1*
b11 6
19
1>
1C
b11 G
#356120000000
0!
0*
09
0>
0C
#356130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#356140000000
0!
0*
09
0>
0C
#356150000000
1!
1*
b101 6
19
1>
1C
b101 G
#356160000000
0!
0*
09
0>
0C
#356170000000
1!
1*
b110 6
19
1>
1C
b110 G
#356180000000
0!
0*
09
0>
0C
#356190000000
1!
1*
b111 6
19
1>
1C
b111 G
#356200000000
0!
0*
09
0>
0C
#356210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#356220000000
0!
0*
09
0>
0C
#356230000000
1!
1*
b1 6
19
1>
1C
b1 G
#356240000000
0!
0*
09
0>
0C
#356250000000
1!
1*
b10 6
19
1>
1C
b10 G
#356260000000
0!
0*
09
0>
0C
#356270000000
1!
1*
b11 6
19
1>
1C
b11 G
#356280000000
0!
0*
09
0>
0C
#356290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#356300000000
0!
0*
09
0>
0C
#356310000000
1!
1*
b101 6
19
1>
1C
b101 G
#356320000000
0!
0*
09
0>
0C
#356330000000
1!
1*
b110 6
19
1>
1C
b110 G
#356340000000
0!
0*
09
0>
0C
#356350000000
1!
1*
b111 6
19
1>
1C
b111 G
#356360000000
0!
1"
0*
1+
09
1:
0>
0C
#356370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#356380000000
0!
0*
09
0>
0C
#356390000000
1!
1*
b1 6
19
1>
1C
b1 G
#356400000000
0!
0*
09
0>
0C
#356410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#356420000000
0!
0*
09
0>
0C
#356430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#356440000000
0!
0*
09
0>
0C
#356450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#356460000000
0!
0*
09
0>
0C
#356470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#356480000000
0!
0#
0*
0,
09
0>
0?
0C
#356490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#356500000000
0!
0*
09
0>
0C
#356510000000
1!
1*
19
1>
1C
#356520000000
0!
0*
09
0>
0C
#356530000000
1!
1*
19
1>
1C
#356540000000
0!
0*
09
0>
0C
#356550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#356560000000
0!
0*
09
0>
0C
#356570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#356580000000
0!
0*
09
0>
0C
#356590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#356600000000
0!
0*
09
0>
0C
#356610000000
1!
1*
b10 6
19
1>
1C
b10 G
#356620000000
0!
0*
09
0>
0C
#356630000000
1!
1*
b11 6
19
1>
1C
b11 G
#356640000000
0!
0*
09
0>
0C
#356650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#356660000000
0!
0*
09
0>
0C
#356670000000
1!
1*
b101 6
19
1>
1C
b101 G
#356680000000
0!
0*
09
0>
0C
#356690000000
1!
1*
b110 6
19
1>
1C
b110 G
#356700000000
0!
0*
09
0>
0C
#356710000000
1!
1*
b111 6
19
1>
1C
b111 G
#356720000000
0!
0*
09
0>
0C
#356730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#356740000000
0!
0*
09
0>
0C
#356750000000
1!
1*
b1 6
19
1>
1C
b1 G
#356760000000
0!
0*
09
0>
0C
#356770000000
1!
1*
b10 6
19
1>
1C
b10 G
#356780000000
0!
0*
09
0>
0C
#356790000000
1!
1*
b11 6
19
1>
1C
b11 G
#356800000000
0!
0*
09
0>
0C
#356810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#356820000000
0!
0*
09
0>
0C
#356830000000
1!
1*
b101 6
19
1>
1C
b101 G
#356840000000
0!
0*
09
0>
0C
#356850000000
1!
1*
b110 6
19
1>
1C
b110 G
#356860000000
0!
0*
09
0>
0C
#356870000000
1!
1*
b111 6
19
1>
1C
b111 G
#356880000000
0!
0*
09
0>
0C
#356890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#356900000000
0!
0*
09
0>
0C
#356910000000
1!
1*
b1 6
19
1>
1C
b1 G
#356920000000
0!
0*
09
0>
0C
#356930000000
1!
1*
b10 6
19
1>
1C
b10 G
#356940000000
0!
0*
09
0>
0C
#356950000000
1!
1*
b11 6
19
1>
1C
b11 G
#356960000000
0!
0*
09
0>
0C
#356970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#356980000000
0!
0*
09
0>
0C
#356990000000
1!
1*
b101 6
19
1>
1C
b101 G
#357000000000
0!
0*
09
0>
0C
#357010000000
1!
1*
b110 6
19
1>
1C
b110 G
#357020000000
0!
0*
09
0>
0C
#357030000000
1!
1*
b111 6
19
1>
1C
b111 G
#357040000000
0!
1"
0*
1+
09
1:
0>
0C
#357050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#357060000000
0!
0*
09
0>
0C
#357070000000
1!
1*
b1 6
19
1>
1C
b1 G
#357080000000
0!
0*
09
0>
0C
#357090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#357100000000
0!
0*
09
0>
0C
#357110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#357120000000
0!
0*
09
0>
0C
#357130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#357140000000
0!
0*
09
0>
0C
#357150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#357160000000
0!
0#
0*
0,
09
0>
0?
0C
#357170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#357180000000
0!
0*
09
0>
0C
#357190000000
1!
1*
19
1>
1C
#357200000000
0!
0*
09
0>
0C
#357210000000
1!
1*
19
1>
1C
#357220000000
0!
0*
09
0>
0C
#357230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#357240000000
0!
0*
09
0>
0C
#357250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#357260000000
0!
0*
09
0>
0C
#357270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#357280000000
0!
0*
09
0>
0C
#357290000000
1!
1*
b10 6
19
1>
1C
b10 G
#357300000000
0!
0*
09
0>
0C
#357310000000
1!
1*
b11 6
19
1>
1C
b11 G
#357320000000
0!
0*
09
0>
0C
#357330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#357340000000
0!
0*
09
0>
0C
#357350000000
1!
1*
b101 6
19
1>
1C
b101 G
#357360000000
0!
0*
09
0>
0C
#357370000000
1!
1*
b110 6
19
1>
1C
b110 G
#357380000000
0!
0*
09
0>
0C
#357390000000
1!
1*
b111 6
19
1>
1C
b111 G
#357400000000
0!
0*
09
0>
0C
#357410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#357420000000
0!
0*
09
0>
0C
#357430000000
1!
1*
b1 6
19
1>
1C
b1 G
#357440000000
0!
0*
09
0>
0C
#357450000000
1!
1*
b10 6
19
1>
1C
b10 G
#357460000000
0!
0*
09
0>
0C
#357470000000
1!
1*
b11 6
19
1>
1C
b11 G
#357480000000
0!
0*
09
0>
0C
#357490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#357500000000
0!
0*
09
0>
0C
#357510000000
1!
1*
b101 6
19
1>
1C
b101 G
#357520000000
0!
0*
09
0>
0C
#357530000000
1!
1*
b110 6
19
1>
1C
b110 G
#357540000000
0!
0*
09
0>
0C
#357550000000
1!
1*
b111 6
19
1>
1C
b111 G
#357560000000
0!
0*
09
0>
0C
#357570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#357580000000
0!
0*
09
0>
0C
#357590000000
1!
1*
b1 6
19
1>
1C
b1 G
#357600000000
0!
0*
09
0>
0C
#357610000000
1!
1*
b10 6
19
1>
1C
b10 G
#357620000000
0!
0*
09
0>
0C
#357630000000
1!
1*
b11 6
19
1>
1C
b11 G
#357640000000
0!
0*
09
0>
0C
#357650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#357660000000
0!
0*
09
0>
0C
#357670000000
1!
1*
b101 6
19
1>
1C
b101 G
#357680000000
0!
0*
09
0>
0C
#357690000000
1!
1*
b110 6
19
1>
1C
b110 G
#357700000000
0!
0*
09
0>
0C
#357710000000
1!
1*
b111 6
19
1>
1C
b111 G
#357720000000
0!
1"
0*
1+
09
1:
0>
0C
#357730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#357740000000
0!
0*
09
0>
0C
#357750000000
1!
1*
b1 6
19
1>
1C
b1 G
#357760000000
0!
0*
09
0>
0C
#357770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#357780000000
0!
0*
09
0>
0C
#357790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#357800000000
0!
0*
09
0>
0C
#357810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#357820000000
0!
0*
09
0>
0C
#357830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#357840000000
0!
0#
0*
0,
09
0>
0?
0C
#357850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#357860000000
0!
0*
09
0>
0C
#357870000000
1!
1*
19
1>
1C
#357880000000
0!
0*
09
0>
0C
#357890000000
1!
1*
19
1>
1C
#357900000000
0!
0*
09
0>
0C
#357910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#357920000000
0!
0*
09
0>
0C
#357930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#357940000000
0!
0*
09
0>
0C
#357950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#357960000000
0!
0*
09
0>
0C
#357970000000
1!
1*
b10 6
19
1>
1C
b10 G
#357980000000
0!
0*
09
0>
0C
#357990000000
1!
1*
b11 6
19
1>
1C
b11 G
#358000000000
0!
0*
09
0>
0C
#358010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#358020000000
0!
0*
09
0>
0C
#358030000000
1!
1*
b101 6
19
1>
1C
b101 G
#358040000000
0!
0*
09
0>
0C
#358050000000
1!
1*
b110 6
19
1>
1C
b110 G
#358060000000
0!
0*
09
0>
0C
#358070000000
1!
1*
b111 6
19
1>
1C
b111 G
#358080000000
0!
0*
09
0>
0C
#358090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#358100000000
0!
0*
09
0>
0C
#358110000000
1!
1*
b1 6
19
1>
1C
b1 G
#358120000000
0!
0*
09
0>
0C
#358130000000
1!
1*
b10 6
19
1>
1C
b10 G
#358140000000
0!
0*
09
0>
0C
#358150000000
1!
1*
b11 6
19
1>
1C
b11 G
#358160000000
0!
0*
09
0>
0C
#358170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#358180000000
0!
0*
09
0>
0C
#358190000000
1!
1*
b101 6
19
1>
1C
b101 G
#358200000000
0!
0*
09
0>
0C
#358210000000
1!
1*
b110 6
19
1>
1C
b110 G
#358220000000
0!
0*
09
0>
0C
#358230000000
1!
1*
b111 6
19
1>
1C
b111 G
#358240000000
0!
0*
09
0>
0C
#358250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#358260000000
0!
0*
09
0>
0C
#358270000000
1!
1*
b1 6
19
1>
1C
b1 G
#358280000000
0!
0*
09
0>
0C
#358290000000
1!
1*
b10 6
19
1>
1C
b10 G
#358300000000
0!
0*
09
0>
0C
#358310000000
1!
1*
b11 6
19
1>
1C
b11 G
#358320000000
0!
0*
09
0>
0C
#358330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#358340000000
0!
0*
09
0>
0C
#358350000000
1!
1*
b101 6
19
1>
1C
b101 G
#358360000000
0!
0*
09
0>
0C
#358370000000
1!
1*
b110 6
19
1>
1C
b110 G
#358380000000
0!
0*
09
0>
0C
#358390000000
1!
1*
b111 6
19
1>
1C
b111 G
#358400000000
0!
1"
0*
1+
09
1:
0>
0C
#358410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#358420000000
0!
0*
09
0>
0C
#358430000000
1!
1*
b1 6
19
1>
1C
b1 G
#358440000000
0!
0*
09
0>
0C
#358450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#358460000000
0!
0*
09
0>
0C
#358470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#358480000000
0!
0*
09
0>
0C
#358490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#358500000000
0!
0*
09
0>
0C
#358510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#358520000000
0!
0#
0*
0,
09
0>
0?
0C
#358530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#358540000000
0!
0*
09
0>
0C
#358550000000
1!
1*
19
1>
1C
#358560000000
0!
0*
09
0>
0C
#358570000000
1!
1*
19
1>
1C
#358580000000
0!
0*
09
0>
0C
#358590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#358600000000
0!
0*
09
0>
0C
#358610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#358620000000
0!
0*
09
0>
0C
#358630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#358640000000
0!
0*
09
0>
0C
#358650000000
1!
1*
b10 6
19
1>
1C
b10 G
#358660000000
0!
0*
09
0>
0C
#358670000000
1!
1*
b11 6
19
1>
1C
b11 G
#358680000000
0!
0*
09
0>
0C
#358690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#358700000000
0!
0*
09
0>
0C
#358710000000
1!
1*
b101 6
19
1>
1C
b101 G
#358720000000
0!
0*
09
0>
0C
#358730000000
1!
1*
b110 6
19
1>
1C
b110 G
#358740000000
0!
0*
09
0>
0C
#358750000000
1!
1*
b111 6
19
1>
1C
b111 G
#358760000000
0!
0*
09
0>
0C
#358770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#358780000000
0!
0*
09
0>
0C
#358790000000
1!
1*
b1 6
19
1>
1C
b1 G
#358800000000
0!
0*
09
0>
0C
#358810000000
1!
1*
b10 6
19
1>
1C
b10 G
#358820000000
0!
0*
09
0>
0C
#358830000000
1!
1*
b11 6
19
1>
1C
b11 G
#358840000000
0!
0*
09
0>
0C
#358850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#358860000000
0!
0*
09
0>
0C
#358870000000
1!
1*
b101 6
19
1>
1C
b101 G
#358880000000
0!
0*
09
0>
0C
#358890000000
1!
1*
b110 6
19
1>
1C
b110 G
#358900000000
0!
0*
09
0>
0C
#358910000000
1!
1*
b111 6
19
1>
1C
b111 G
#358920000000
0!
0*
09
0>
0C
#358930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#358940000000
0!
0*
09
0>
0C
#358950000000
1!
1*
b1 6
19
1>
1C
b1 G
#358960000000
0!
0*
09
0>
0C
#358970000000
1!
1*
b10 6
19
1>
1C
b10 G
#358980000000
0!
0*
09
0>
0C
#358990000000
1!
1*
b11 6
19
1>
1C
b11 G
#359000000000
0!
0*
09
0>
0C
#359010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#359020000000
0!
0*
09
0>
0C
#359030000000
1!
1*
b101 6
19
1>
1C
b101 G
#359040000000
0!
0*
09
0>
0C
#359050000000
1!
1*
b110 6
19
1>
1C
b110 G
#359060000000
0!
0*
09
0>
0C
#359070000000
1!
1*
b111 6
19
1>
1C
b111 G
#359080000000
0!
1"
0*
1+
09
1:
0>
0C
#359090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#359100000000
0!
0*
09
0>
0C
#359110000000
1!
1*
b1 6
19
1>
1C
b1 G
#359120000000
0!
0*
09
0>
0C
#359130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#359140000000
0!
0*
09
0>
0C
#359150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#359160000000
0!
0*
09
0>
0C
#359170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#359180000000
0!
0*
09
0>
0C
#359190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#359200000000
0!
0#
0*
0,
09
0>
0?
0C
#359210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#359220000000
0!
0*
09
0>
0C
#359230000000
1!
1*
19
1>
1C
#359240000000
0!
0*
09
0>
0C
#359250000000
1!
1*
19
1>
1C
#359260000000
0!
0*
09
0>
0C
#359270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#359280000000
0!
0*
09
0>
0C
#359290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#359300000000
0!
0*
09
0>
0C
#359310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#359320000000
0!
0*
09
0>
0C
#359330000000
1!
1*
b10 6
19
1>
1C
b10 G
#359340000000
0!
0*
09
0>
0C
#359350000000
1!
1*
b11 6
19
1>
1C
b11 G
#359360000000
0!
0*
09
0>
0C
#359370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#359380000000
0!
0*
09
0>
0C
#359390000000
1!
1*
b101 6
19
1>
1C
b101 G
#359400000000
0!
0*
09
0>
0C
#359410000000
1!
1*
b110 6
19
1>
1C
b110 G
#359420000000
0!
0*
09
0>
0C
#359430000000
1!
1*
b111 6
19
1>
1C
b111 G
#359440000000
0!
0*
09
0>
0C
#359450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#359460000000
0!
0*
09
0>
0C
#359470000000
1!
1*
b1 6
19
1>
1C
b1 G
#359480000000
0!
0*
09
0>
0C
#359490000000
1!
1*
b10 6
19
1>
1C
b10 G
#359500000000
0!
0*
09
0>
0C
#359510000000
1!
1*
b11 6
19
1>
1C
b11 G
#359520000000
0!
0*
09
0>
0C
#359530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#359540000000
0!
0*
09
0>
0C
#359550000000
1!
1*
b101 6
19
1>
1C
b101 G
#359560000000
0!
0*
09
0>
0C
#359570000000
1!
1*
b110 6
19
1>
1C
b110 G
#359580000000
0!
0*
09
0>
0C
#359590000000
1!
1*
b111 6
19
1>
1C
b111 G
#359600000000
0!
0*
09
0>
0C
#359610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#359620000000
0!
0*
09
0>
0C
#359630000000
1!
1*
b1 6
19
1>
1C
b1 G
#359640000000
0!
0*
09
0>
0C
#359650000000
1!
1*
b10 6
19
1>
1C
b10 G
#359660000000
0!
0*
09
0>
0C
#359670000000
1!
1*
b11 6
19
1>
1C
b11 G
#359680000000
0!
0*
09
0>
0C
#359690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#359700000000
0!
0*
09
0>
0C
#359710000000
1!
1*
b101 6
19
1>
1C
b101 G
#359720000000
0!
0*
09
0>
0C
#359730000000
1!
1*
b110 6
19
1>
1C
b110 G
#359740000000
0!
0*
09
0>
0C
#359750000000
1!
1*
b111 6
19
1>
1C
b111 G
#359760000000
0!
1"
0*
1+
09
1:
0>
0C
#359770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#359780000000
0!
0*
09
0>
0C
#359790000000
1!
1*
b1 6
19
1>
1C
b1 G
#359800000000
0!
0*
09
0>
0C
#359810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#359820000000
0!
0*
09
0>
0C
#359830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#359840000000
0!
0*
09
0>
0C
#359850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#359860000000
0!
0*
09
0>
0C
#359870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#359880000000
0!
0#
0*
0,
09
0>
0?
0C
#359890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#359900000000
0!
0*
09
0>
0C
#359910000000
1!
1*
19
1>
1C
#359920000000
0!
0*
09
0>
0C
#359930000000
1!
1*
19
1>
1C
#359940000000
0!
0*
09
0>
0C
#359950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#359960000000
0!
0*
09
0>
0C
#359970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#359980000000
0!
0*
09
0>
0C
#359990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#360000000000
0!
0*
09
0>
0C
#360010000000
1!
1*
b10 6
19
1>
1C
b10 G
#360020000000
0!
0*
09
0>
0C
#360030000000
1!
1*
b11 6
19
1>
1C
b11 G
#360040000000
0!
0*
09
0>
0C
#360050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#360060000000
0!
0*
09
0>
0C
#360070000000
1!
1*
b101 6
19
1>
1C
b101 G
#360080000000
0!
0*
09
0>
0C
#360090000000
1!
1*
b110 6
19
1>
1C
b110 G
#360100000000
0!
0*
09
0>
0C
#360110000000
1!
1*
b111 6
19
1>
1C
b111 G
#360120000000
0!
0*
09
0>
0C
#360130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#360140000000
0!
0*
09
0>
0C
#360150000000
1!
1*
b1 6
19
1>
1C
b1 G
#360160000000
0!
0*
09
0>
0C
#360170000000
1!
1*
b10 6
19
1>
1C
b10 G
#360180000000
0!
0*
09
0>
0C
#360190000000
1!
1*
b11 6
19
1>
1C
b11 G
#360200000000
0!
0*
09
0>
0C
#360210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#360220000000
0!
0*
09
0>
0C
#360230000000
1!
1*
b101 6
19
1>
1C
b101 G
#360240000000
0!
0*
09
0>
0C
#360250000000
1!
1*
b110 6
19
1>
1C
b110 G
#360260000000
0!
0*
09
0>
0C
#360270000000
1!
1*
b111 6
19
1>
1C
b111 G
#360280000000
0!
0*
09
0>
0C
#360290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#360300000000
0!
0*
09
0>
0C
#360310000000
1!
1*
b1 6
19
1>
1C
b1 G
#360320000000
0!
0*
09
0>
0C
#360330000000
1!
1*
b10 6
19
1>
1C
b10 G
#360340000000
0!
0*
09
0>
0C
#360350000000
1!
1*
b11 6
19
1>
1C
b11 G
#360360000000
0!
0*
09
0>
0C
#360370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#360380000000
0!
0*
09
0>
0C
#360390000000
1!
1*
b101 6
19
1>
1C
b101 G
#360400000000
0!
0*
09
0>
0C
#360410000000
1!
1*
b110 6
19
1>
1C
b110 G
#360420000000
0!
0*
09
0>
0C
#360430000000
1!
1*
b111 6
19
1>
1C
b111 G
#360440000000
0!
1"
0*
1+
09
1:
0>
0C
#360450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#360460000000
0!
0*
09
0>
0C
#360470000000
1!
1*
b1 6
19
1>
1C
b1 G
#360480000000
0!
0*
09
0>
0C
#360490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#360500000000
0!
0*
09
0>
0C
#360510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#360520000000
0!
0*
09
0>
0C
#360530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#360540000000
0!
0*
09
0>
0C
#360550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#360560000000
0!
0#
0*
0,
09
0>
0?
0C
#360570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#360580000000
0!
0*
09
0>
0C
#360590000000
1!
1*
19
1>
1C
#360600000000
0!
0*
09
0>
0C
#360610000000
1!
1*
19
1>
1C
#360620000000
0!
0*
09
0>
0C
#360630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#360640000000
0!
0*
09
0>
0C
#360650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#360660000000
0!
0*
09
0>
0C
#360670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#360680000000
0!
0*
09
0>
0C
#360690000000
1!
1*
b10 6
19
1>
1C
b10 G
#360700000000
0!
0*
09
0>
0C
#360710000000
1!
1*
b11 6
19
1>
1C
b11 G
#360720000000
0!
0*
09
0>
0C
#360730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#360740000000
0!
0*
09
0>
0C
#360750000000
1!
1*
b101 6
19
1>
1C
b101 G
#360760000000
0!
0*
09
0>
0C
#360770000000
1!
1*
b110 6
19
1>
1C
b110 G
#360780000000
0!
0*
09
0>
0C
#360790000000
1!
1*
b111 6
19
1>
1C
b111 G
#360800000000
0!
0*
09
0>
0C
#360810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#360820000000
0!
0*
09
0>
0C
#360830000000
1!
1*
b1 6
19
1>
1C
b1 G
#360840000000
0!
0*
09
0>
0C
#360850000000
1!
1*
b10 6
19
1>
1C
b10 G
#360860000000
0!
0*
09
0>
0C
#360870000000
1!
1*
b11 6
19
1>
1C
b11 G
#360880000000
0!
0*
09
0>
0C
#360890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#360900000000
0!
0*
09
0>
0C
#360910000000
1!
1*
b101 6
19
1>
1C
b101 G
#360920000000
0!
0*
09
0>
0C
#360930000000
1!
1*
b110 6
19
1>
1C
b110 G
#360940000000
0!
0*
09
0>
0C
#360950000000
1!
1*
b111 6
19
1>
1C
b111 G
#360960000000
0!
0*
09
0>
0C
#360970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#360980000000
0!
0*
09
0>
0C
#360990000000
1!
1*
b1 6
19
1>
1C
b1 G
#361000000000
0!
0*
09
0>
0C
#361010000000
1!
1*
b10 6
19
1>
1C
b10 G
#361020000000
0!
0*
09
0>
0C
#361030000000
1!
1*
b11 6
19
1>
1C
b11 G
#361040000000
0!
0*
09
0>
0C
#361050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#361060000000
0!
0*
09
0>
0C
#361070000000
1!
1*
b101 6
19
1>
1C
b101 G
#361080000000
0!
0*
09
0>
0C
#361090000000
1!
1*
b110 6
19
1>
1C
b110 G
#361100000000
0!
0*
09
0>
0C
#361110000000
1!
1*
b111 6
19
1>
1C
b111 G
#361120000000
0!
1"
0*
1+
09
1:
0>
0C
#361130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#361140000000
0!
0*
09
0>
0C
#361150000000
1!
1*
b1 6
19
1>
1C
b1 G
#361160000000
0!
0*
09
0>
0C
#361170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#361180000000
0!
0*
09
0>
0C
#361190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#361200000000
0!
0*
09
0>
0C
#361210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#361220000000
0!
0*
09
0>
0C
#361230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#361240000000
0!
0#
0*
0,
09
0>
0?
0C
#361250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#361260000000
0!
0*
09
0>
0C
#361270000000
1!
1*
19
1>
1C
#361280000000
0!
0*
09
0>
0C
#361290000000
1!
1*
19
1>
1C
#361300000000
0!
0*
09
0>
0C
#361310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#361320000000
0!
0*
09
0>
0C
#361330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#361340000000
0!
0*
09
0>
0C
#361350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#361360000000
0!
0*
09
0>
0C
#361370000000
1!
1*
b10 6
19
1>
1C
b10 G
#361380000000
0!
0*
09
0>
0C
#361390000000
1!
1*
b11 6
19
1>
1C
b11 G
#361400000000
0!
0*
09
0>
0C
#361410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#361420000000
0!
0*
09
0>
0C
#361430000000
1!
1*
b101 6
19
1>
1C
b101 G
#361440000000
0!
0*
09
0>
0C
#361450000000
1!
1*
b110 6
19
1>
1C
b110 G
#361460000000
0!
0*
09
0>
0C
#361470000000
1!
1*
b111 6
19
1>
1C
b111 G
#361480000000
0!
0*
09
0>
0C
#361490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#361500000000
0!
0*
09
0>
0C
#361510000000
1!
1*
b1 6
19
1>
1C
b1 G
#361520000000
0!
0*
09
0>
0C
#361530000000
1!
1*
b10 6
19
1>
1C
b10 G
#361540000000
0!
0*
09
0>
0C
#361550000000
1!
1*
b11 6
19
1>
1C
b11 G
#361560000000
0!
0*
09
0>
0C
#361570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#361580000000
0!
0*
09
0>
0C
#361590000000
1!
1*
b101 6
19
1>
1C
b101 G
#361600000000
0!
0*
09
0>
0C
#361610000000
1!
1*
b110 6
19
1>
1C
b110 G
#361620000000
0!
0*
09
0>
0C
#361630000000
1!
1*
b111 6
19
1>
1C
b111 G
#361640000000
0!
0*
09
0>
0C
#361650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#361660000000
0!
0*
09
0>
0C
#361670000000
1!
1*
b1 6
19
1>
1C
b1 G
#361680000000
0!
0*
09
0>
0C
#361690000000
1!
1*
b10 6
19
1>
1C
b10 G
#361700000000
0!
0*
09
0>
0C
#361710000000
1!
1*
b11 6
19
1>
1C
b11 G
#361720000000
0!
0*
09
0>
0C
#361730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#361740000000
0!
0*
09
0>
0C
#361750000000
1!
1*
b101 6
19
1>
1C
b101 G
#361760000000
0!
0*
09
0>
0C
#361770000000
1!
1*
b110 6
19
1>
1C
b110 G
#361780000000
0!
0*
09
0>
0C
#361790000000
1!
1*
b111 6
19
1>
1C
b111 G
#361800000000
0!
1"
0*
1+
09
1:
0>
0C
#361810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#361820000000
0!
0*
09
0>
0C
#361830000000
1!
1*
b1 6
19
1>
1C
b1 G
#361840000000
0!
0*
09
0>
0C
#361850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#361860000000
0!
0*
09
0>
0C
#361870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#361880000000
0!
0*
09
0>
0C
#361890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#361900000000
0!
0*
09
0>
0C
#361910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#361920000000
0!
0#
0*
0,
09
0>
0?
0C
#361930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#361940000000
0!
0*
09
0>
0C
#361950000000
1!
1*
19
1>
1C
#361960000000
0!
0*
09
0>
0C
#361970000000
1!
1*
19
1>
1C
#361980000000
0!
0*
09
0>
0C
#361990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#362000000000
0!
0*
09
0>
0C
#362010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#362020000000
0!
0*
09
0>
0C
#362030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#362040000000
0!
0*
09
0>
0C
#362050000000
1!
1*
b10 6
19
1>
1C
b10 G
#362060000000
0!
0*
09
0>
0C
#362070000000
1!
1*
b11 6
19
1>
1C
b11 G
#362080000000
0!
0*
09
0>
0C
#362090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#362100000000
0!
0*
09
0>
0C
#362110000000
1!
1*
b101 6
19
1>
1C
b101 G
#362120000000
0!
0*
09
0>
0C
#362130000000
1!
1*
b110 6
19
1>
1C
b110 G
#362140000000
0!
0*
09
0>
0C
#362150000000
1!
1*
b111 6
19
1>
1C
b111 G
#362160000000
0!
0*
09
0>
0C
#362170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#362180000000
0!
0*
09
0>
0C
#362190000000
1!
1*
b1 6
19
1>
1C
b1 G
#362200000000
0!
0*
09
0>
0C
#362210000000
1!
1*
b10 6
19
1>
1C
b10 G
#362220000000
0!
0*
09
0>
0C
#362230000000
1!
1*
b11 6
19
1>
1C
b11 G
#362240000000
0!
0*
09
0>
0C
#362250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#362260000000
0!
0*
09
0>
0C
#362270000000
1!
1*
b101 6
19
1>
1C
b101 G
#362280000000
0!
0*
09
0>
0C
#362290000000
1!
1*
b110 6
19
1>
1C
b110 G
#362300000000
0!
0*
09
0>
0C
#362310000000
1!
1*
b111 6
19
1>
1C
b111 G
#362320000000
0!
0*
09
0>
0C
#362330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#362340000000
0!
0*
09
0>
0C
#362350000000
1!
1*
b1 6
19
1>
1C
b1 G
#362360000000
0!
0*
09
0>
0C
#362370000000
1!
1*
b10 6
19
1>
1C
b10 G
#362380000000
0!
0*
09
0>
0C
#362390000000
1!
1*
b11 6
19
1>
1C
b11 G
#362400000000
0!
0*
09
0>
0C
#362410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#362420000000
0!
0*
09
0>
0C
#362430000000
1!
1*
b101 6
19
1>
1C
b101 G
#362440000000
0!
0*
09
0>
0C
#362450000000
1!
1*
b110 6
19
1>
1C
b110 G
#362460000000
0!
0*
09
0>
0C
#362470000000
1!
1*
b111 6
19
1>
1C
b111 G
#362480000000
0!
1"
0*
1+
09
1:
0>
0C
#362490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#362500000000
0!
0*
09
0>
0C
#362510000000
1!
1*
b1 6
19
1>
1C
b1 G
#362520000000
0!
0*
09
0>
0C
#362530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#362540000000
0!
0*
09
0>
0C
#362550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#362560000000
0!
0*
09
0>
0C
#362570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#362580000000
0!
0*
09
0>
0C
#362590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#362600000000
0!
0#
0*
0,
09
0>
0?
0C
#362610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#362620000000
0!
0*
09
0>
0C
#362630000000
1!
1*
19
1>
1C
#362640000000
0!
0*
09
0>
0C
#362650000000
1!
1*
19
1>
1C
#362660000000
0!
0*
09
0>
0C
#362670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#362680000000
0!
0*
09
0>
0C
#362690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#362700000000
0!
0*
09
0>
0C
#362710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#362720000000
0!
0*
09
0>
0C
#362730000000
1!
1*
b10 6
19
1>
1C
b10 G
#362740000000
0!
0*
09
0>
0C
#362750000000
1!
1*
b11 6
19
1>
1C
b11 G
#362760000000
0!
0*
09
0>
0C
#362770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#362780000000
0!
0*
09
0>
0C
#362790000000
1!
1*
b101 6
19
1>
1C
b101 G
#362800000000
0!
0*
09
0>
0C
#362810000000
1!
1*
b110 6
19
1>
1C
b110 G
#362820000000
0!
0*
09
0>
0C
#362830000000
1!
1*
b111 6
19
1>
1C
b111 G
#362840000000
0!
0*
09
0>
0C
#362850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#362860000000
0!
0*
09
0>
0C
#362870000000
1!
1*
b1 6
19
1>
1C
b1 G
#362880000000
0!
0*
09
0>
0C
#362890000000
1!
1*
b10 6
19
1>
1C
b10 G
#362900000000
0!
0*
09
0>
0C
#362910000000
1!
1*
b11 6
19
1>
1C
b11 G
#362920000000
0!
0*
09
0>
0C
#362930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#362940000000
0!
0*
09
0>
0C
#362950000000
1!
1*
b101 6
19
1>
1C
b101 G
#362960000000
0!
0*
09
0>
0C
#362970000000
1!
1*
b110 6
19
1>
1C
b110 G
#362980000000
0!
0*
09
0>
0C
#362990000000
1!
1*
b111 6
19
1>
1C
b111 G
#363000000000
0!
0*
09
0>
0C
#363010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#363020000000
0!
0*
09
0>
0C
#363030000000
1!
1*
b1 6
19
1>
1C
b1 G
#363040000000
0!
0*
09
0>
0C
#363050000000
1!
1*
b10 6
19
1>
1C
b10 G
#363060000000
0!
0*
09
0>
0C
#363070000000
1!
1*
b11 6
19
1>
1C
b11 G
#363080000000
0!
0*
09
0>
0C
#363090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#363100000000
0!
0*
09
0>
0C
#363110000000
1!
1*
b101 6
19
1>
1C
b101 G
#363120000000
0!
0*
09
0>
0C
#363130000000
1!
1*
b110 6
19
1>
1C
b110 G
#363140000000
0!
0*
09
0>
0C
#363150000000
1!
1*
b111 6
19
1>
1C
b111 G
#363160000000
0!
1"
0*
1+
09
1:
0>
0C
#363170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#363180000000
0!
0*
09
0>
0C
#363190000000
1!
1*
b1 6
19
1>
1C
b1 G
#363200000000
0!
0*
09
0>
0C
#363210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#363220000000
0!
0*
09
0>
0C
#363230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#363240000000
0!
0*
09
0>
0C
#363250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#363260000000
0!
0*
09
0>
0C
#363270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#363280000000
0!
0#
0*
0,
09
0>
0?
0C
#363290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#363300000000
0!
0*
09
0>
0C
#363310000000
1!
1*
19
1>
1C
#363320000000
0!
0*
09
0>
0C
#363330000000
1!
1*
19
1>
1C
#363340000000
0!
0*
09
0>
0C
#363350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#363360000000
0!
0*
09
0>
0C
#363370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#363380000000
0!
0*
09
0>
0C
#363390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#363400000000
0!
0*
09
0>
0C
#363410000000
1!
1*
b10 6
19
1>
1C
b10 G
#363420000000
0!
0*
09
0>
0C
#363430000000
1!
1*
b11 6
19
1>
1C
b11 G
#363440000000
0!
0*
09
0>
0C
#363450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#363460000000
0!
0*
09
0>
0C
#363470000000
1!
1*
b101 6
19
1>
1C
b101 G
#363480000000
0!
0*
09
0>
0C
#363490000000
1!
1*
b110 6
19
1>
1C
b110 G
#363500000000
0!
0*
09
0>
0C
#363510000000
1!
1*
b111 6
19
1>
1C
b111 G
#363520000000
0!
0*
09
0>
0C
#363530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#363540000000
0!
0*
09
0>
0C
#363550000000
1!
1*
b1 6
19
1>
1C
b1 G
#363560000000
0!
0*
09
0>
0C
#363570000000
1!
1*
b10 6
19
1>
1C
b10 G
#363580000000
0!
0*
09
0>
0C
#363590000000
1!
1*
b11 6
19
1>
1C
b11 G
#363600000000
0!
0*
09
0>
0C
#363610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#363620000000
0!
0*
09
0>
0C
#363630000000
1!
1*
b101 6
19
1>
1C
b101 G
#363640000000
0!
0*
09
0>
0C
#363650000000
1!
1*
b110 6
19
1>
1C
b110 G
#363660000000
0!
0*
09
0>
0C
#363670000000
1!
1*
b111 6
19
1>
1C
b111 G
#363680000000
0!
0*
09
0>
0C
#363690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#363700000000
0!
0*
09
0>
0C
#363710000000
1!
1*
b1 6
19
1>
1C
b1 G
#363720000000
0!
0*
09
0>
0C
#363730000000
1!
1*
b10 6
19
1>
1C
b10 G
#363740000000
0!
0*
09
0>
0C
#363750000000
1!
1*
b11 6
19
1>
1C
b11 G
#363760000000
0!
0*
09
0>
0C
#363770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#363780000000
0!
0*
09
0>
0C
#363790000000
1!
1*
b101 6
19
1>
1C
b101 G
#363800000000
0!
0*
09
0>
0C
#363810000000
1!
1*
b110 6
19
1>
1C
b110 G
#363820000000
0!
0*
09
0>
0C
#363830000000
1!
1*
b111 6
19
1>
1C
b111 G
#363840000000
0!
1"
0*
1+
09
1:
0>
0C
#363850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#363860000000
0!
0*
09
0>
0C
#363870000000
1!
1*
b1 6
19
1>
1C
b1 G
#363880000000
0!
0*
09
0>
0C
#363890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#363900000000
0!
0*
09
0>
0C
#363910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#363920000000
0!
0*
09
0>
0C
#363930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#363940000000
0!
0*
09
0>
0C
#363950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#363960000000
0!
0#
0*
0,
09
0>
0?
0C
#363970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#363980000000
0!
0*
09
0>
0C
#363990000000
1!
1*
19
1>
1C
#364000000000
0!
0*
09
0>
0C
#364010000000
1!
1*
19
1>
1C
#364020000000
0!
0*
09
0>
0C
#364030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#364040000000
0!
0*
09
0>
0C
#364050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#364060000000
0!
0*
09
0>
0C
#364070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#364080000000
0!
0*
09
0>
0C
#364090000000
1!
1*
b10 6
19
1>
1C
b10 G
#364100000000
0!
0*
09
0>
0C
#364110000000
1!
1*
b11 6
19
1>
1C
b11 G
#364120000000
0!
0*
09
0>
0C
#364130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#364140000000
0!
0*
09
0>
0C
#364150000000
1!
1*
b101 6
19
1>
1C
b101 G
#364160000000
0!
0*
09
0>
0C
#364170000000
1!
1*
b110 6
19
1>
1C
b110 G
#364180000000
0!
0*
09
0>
0C
#364190000000
1!
1*
b111 6
19
1>
1C
b111 G
#364200000000
0!
0*
09
0>
0C
#364210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#364220000000
0!
0*
09
0>
0C
#364230000000
1!
1*
b1 6
19
1>
1C
b1 G
#364240000000
0!
0*
09
0>
0C
#364250000000
1!
1*
b10 6
19
1>
1C
b10 G
#364260000000
0!
0*
09
0>
0C
#364270000000
1!
1*
b11 6
19
1>
1C
b11 G
#364280000000
0!
0*
09
0>
0C
#364290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#364300000000
0!
0*
09
0>
0C
#364310000000
1!
1*
b101 6
19
1>
1C
b101 G
#364320000000
0!
0*
09
0>
0C
#364330000000
1!
1*
b110 6
19
1>
1C
b110 G
#364340000000
0!
0*
09
0>
0C
#364350000000
1!
1*
b111 6
19
1>
1C
b111 G
#364360000000
0!
0*
09
0>
0C
#364370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#364380000000
0!
0*
09
0>
0C
#364390000000
1!
1*
b1 6
19
1>
1C
b1 G
#364400000000
0!
0*
09
0>
0C
#364410000000
1!
1*
b10 6
19
1>
1C
b10 G
#364420000000
0!
0*
09
0>
0C
#364430000000
1!
1*
b11 6
19
1>
1C
b11 G
#364440000000
0!
0*
09
0>
0C
#364450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#364460000000
0!
0*
09
0>
0C
#364470000000
1!
1*
b101 6
19
1>
1C
b101 G
#364480000000
0!
0*
09
0>
0C
#364490000000
1!
1*
b110 6
19
1>
1C
b110 G
#364500000000
0!
0*
09
0>
0C
#364510000000
1!
1*
b111 6
19
1>
1C
b111 G
#364520000000
0!
1"
0*
1+
09
1:
0>
0C
#364530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#364540000000
0!
0*
09
0>
0C
#364550000000
1!
1*
b1 6
19
1>
1C
b1 G
#364560000000
0!
0*
09
0>
0C
#364570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#364580000000
0!
0*
09
0>
0C
#364590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#364600000000
0!
0*
09
0>
0C
#364610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#364620000000
0!
0*
09
0>
0C
#364630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#364640000000
0!
0#
0*
0,
09
0>
0?
0C
#364650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#364660000000
0!
0*
09
0>
0C
#364670000000
1!
1*
19
1>
1C
#364680000000
0!
0*
09
0>
0C
#364690000000
1!
1*
19
1>
1C
#364700000000
0!
0*
09
0>
0C
#364710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#364720000000
0!
0*
09
0>
0C
#364730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#364740000000
0!
0*
09
0>
0C
#364750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#364760000000
0!
0*
09
0>
0C
#364770000000
1!
1*
b10 6
19
1>
1C
b10 G
#364780000000
0!
0*
09
0>
0C
#364790000000
1!
1*
b11 6
19
1>
1C
b11 G
#364800000000
0!
0*
09
0>
0C
#364810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#364820000000
0!
0*
09
0>
0C
#364830000000
1!
1*
b101 6
19
1>
1C
b101 G
#364840000000
0!
0*
09
0>
0C
#364850000000
1!
1*
b110 6
19
1>
1C
b110 G
#364860000000
0!
0*
09
0>
0C
#364870000000
1!
1*
b111 6
19
1>
1C
b111 G
#364880000000
0!
0*
09
0>
0C
#364890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#364900000000
0!
0*
09
0>
0C
#364910000000
1!
1*
b1 6
19
1>
1C
b1 G
#364920000000
0!
0*
09
0>
0C
#364930000000
1!
1*
b10 6
19
1>
1C
b10 G
#364940000000
0!
0*
09
0>
0C
#364950000000
1!
1*
b11 6
19
1>
1C
b11 G
#364960000000
0!
0*
09
0>
0C
#364970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#364980000000
0!
0*
09
0>
0C
#364990000000
1!
1*
b101 6
19
1>
1C
b101 G
#365000000000
0!
0*
09
0>
0C
#365010000000
1!
1*
b110 6
19
1>
1C
b110 G
#365020000000
0!
0*
09
0>
0C
#365030000000
1!
1*
b111 6
19
1>
1C
b111 G
#365040000000
0!
0*
09
0>
0C
#365050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#365060000000
0!
0*
09
0>
0C
#365070000000
1!
1*
b1 6
19
1>
1C
b1 G
#365080000000
0!
0*
09
0>
0C
#365090000000
1!
1*
b10 6
19
1>
1C
b10 G
#365100000000
0!
0*
09
0>
0C
#365110000000
1!
1*
b11 6
19
1>
1C
b11 G
#365120000000
0!
0*
09
0>
0C
#365130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#365140000000
0!
0*
09
0>
0C
#365150000000
1!
1*
b101 6
19
1>
1C
b101 G
#365160000000
0!
0*
09
0>
0C
#365170000000
1!
1*
b110 6
19
1>
1C
b110 G
#365180000000
0!
0*
09
0>
0C
#365190000000
1!
1*
b111 6
19
1>
1C
b111 G
#365200000000
0!
1"
0*
1+
09
1:
0>
0C
#365210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#365220000000
0!
0*
09
0>
0C
#365230000000
1!
1*
b1 6
19
1>
1C
b1 G
#365240000000
0!
0*
09
0>
0C
#365250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#365260000000
0!
0*
09
0>
0C
#365270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#365280000000
0!
0*
09
0>
0C
#365290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#365300000000
0!
0*
09
0>
0C
#365310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#365320000000
0!
0#
0*
0,
09
0>
0?
0C
#365330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#365340000000
0!
0*
09
0>
0C
#365350000000
1!
1*
19
1>
1C
#365360000000
0!
0*
09
0>
0C
#365370000000
1!
1*
19
1>
1C
#365380000000
0!
0*
09
0>
0C
#365390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#365400000000
0!
0*
09
0>
0C
#365410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#365420000000
0!
0*
09
0>
0C
#365430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#365440000000
0!
0*
09
0>
0C
#365450000000
1!
1*
b10 6
19
1>
1C
b10 G
#365460000000
0!
0*
09
0>
0C
#365470000000
1!
1*
b11 6
19
1>
1C
b11 G
#365480000000
0!
0*
09
0>
0C
#365490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#365500000000
0!
0*
09
0>
0C
#365510000000
1!
1*
b101 6
19
1>
1C
b101 G
#365520000000
0!
0*
09
0>
0C
#365530000000
1!
1*
b110 6
19
1>
1C
b110 G
#365540000000
0!
0*
09
0>
0C
#365550000000
1!
1*
b111 6
19
1>
1C
b111 G
#365560000000
0!
0*
09
0>
0C
#365570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#365580000000
0!
0*
09
0>
0C
#365590000000
1!
1*
b1 6
19
1>
1C
b1 G
#365600000000
0!
0*
09
0>
0C
#365610000000
1!
1*
b10 6
19
1>
1C
b10 G
#365620000000
0!
0*
09
0>
0C
#365630000000
1!
1*
b11 6
19
1>
1C
b11 G
#365640000000
0!
0*
09
0>
0C
#365650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#365660000000
0!
0*
09
0>
0C
#365670000000
1!
1*
b101 6
19
1>
1C
b101 G
#365680000000
0!
0*
09
0>
0C
#365690000000
1!
1*
b110 6
19
1>
1C
b110 G
#365700000000
0!
0*
09
0>
0C
#365710000000
1!
1*
b111 6
19
1>
1C
b111 G
#365720000000
0!
0*
09
0>
0C
#365730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#365740000000
0!
0*
09
0>
0C
#365750000000
1!
1*
b1 6
19
1>
1C
b1 G
#365760000000
0!
0*
09
0>
0C
#365770000000
1!
1*
b10 6
19
1>
1C
b10 G
#365780000000
0!
0*
09
0>
0C
#365790000000
1!
1*
b11 6
19
1>
1C
b11 G
#365800000000
0!
0*
09
0>
0C
#365810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#365820000000
0!
0*
09
0>
0C
#365830000000
1!
1*
b101 6
19
1>
1C
b101 G
#365840000000
0!
0*
09
0>
0C
#365850000000
1!
1*
b110 6
19
1>
1C
b110 G
#365860000000
0!
0*
09
0>
0C
#365870000000
1!
1*
b111 6
19
1>
1C
b111 G
#365880000000
0!
1"
0*
1+
09
1:
0>
0C
#365890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#365900000000
0!
0*
09
0>
0C
#365910000000
1!
1*
b1 6
19
1>
1C
b1 G
#365920000000
0!
0*
09
0>
0C
#365930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#365940000000
0!
0*
09
0>
0C
#365950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#365960000000
0!
0*
09
0>
0C
#365970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#365980000000
0!
0*
09
0>
0C
#365990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#366000000000
0!
0#
0*
0,
09
0>
0?
0C
#366010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#366020000000
0!
0*
09
0>
0C
#366030000000
1!
1*
19
1>
1C
#366040000000
0!
0*
09
0>
0C
#366050000000
1!
1*
19
1>
1C
#366060000000
0!
0*
09
0>
0C
#366070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#366080000000
0!
0*
09
0>
0C
#366090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#366100000000
0!
0*
09
0>
0C
#366110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#366120000000
0!
0*
09
0>
0C
#366130000000
1!
1*
b10 6
19
1>
1C
b10 G
#366140000000
0!
0*
09
0>
0C
#366150000000
1!
1*
b11 6
19
1>
1C
b11 G
#366160000000
0!
0*
09
0>
0C
#366170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#366180000000
0!
0*
09
0>
0C
#366190000000
1!
1*
b101 6
19
1>
1C
b101 G
#366200000000
0!
0*
09
0>
0C
#366210000000
1!
1*
b110 6
19
1>
1C
b110 G
#366220000000
0!
0*
09
0>
0C
#366230000000
1!
1*
b111 6
19
1>
1C
b111 G
#366240000000
0!
0*
09
0>
0C
#366250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#366260000000
0!
0*
09
0>
0C
#366270000000
1!
1*
b1 6
19
1>
1C
b1 G
#366280000000
0!
0*
09
0>
0C
#366290000000
1!
1*
b10 6
19
1>
1C
b10 G
#366300000000
0!
0*
09
0>
0C
#366310000000
1!
1*
b11 6
19
1>
1C
b11 G
#366320000000
0!
0*
09
0>
0C
#366330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#366340000000
0!
0*
09
0>
0C
#366350000000
1!
1*
b101 6
19
1>
1C
b101 G
#366360000000
0!
0*
09
0>
0C
#366370000000
1!
1*
b110 6
19
1>
1C
b110 G
#366380000000
0!
0*
09
0>
0C
#366390000000
1!
1*
b111 6
19
1>
1C
b111 G
#366400000000
0!
0*
09
0>
0C
#366410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#366420000000
0!
0*
09
0>
0C
#366430000000
1!
1*
b1 6
19
1>
1C
b1 G
#366440000000
0!
0*
09
0>
0C
#366450000000
1!
1*
b10 6
19
1>
1C
b10 G
#366460000000
0!
0*
09
0>
0C
#366470000000
1!
1*
b11 6
19
1>
1C
b11 G
#366480000000
0!
0*
09
0>
0C
#366490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#366500000000
0!
0*
09
0>
0C
#366510000000
1!
1*
b101 6
19
1>
1C
b101 G
#366520000000
0!
0*
09
0>
0C
#366530000000
1!
1*
b110 6
19
1>
1C
b110 G
#366540000000
0!
0*
09
0>
0C
#366550000000
1!
1*
b111 6
19
1>
1C
b111 G
#366560000000
0!
1"
0*
1+
09
1:
0>
0C
#366570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#366580000000
0!
0*
09
0>
0C
#366590000000
1!
1*
b1 6
19
1>
1C
b1 G
#366600000000
0!
0*
09
0>
0C
#366610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#366620000000
0!
0*
09
0>
0C
#366630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#366640000000
0!
0*
09
0>
0C
#366650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#366660000000
0!
0*
09
0>
0C
#366670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#366680000000
0!
0#
0*
0,
09
0>
0?
0C
#366690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#366700000000
0!
0*
09
0>
0C
#366710000000
1!
1*
19
1>
1C
#366720000000
0!
0*
09
0>
0C
#366730000000
1!
1*
19
1>
1C
#366740000000
0!
0*
09
0>
0C
#366750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#366760000000
0!
0*
09
0>
0C
#366770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#366780000000
0!
0*
09
0>
0C
#366790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#366800000000
0!
0*
09
0>
0C
#366810000000
1!
1*
b10 6
19
1>
1C
b10 G
#366820000000
0!
0*
09
0>
0C
#366830000000
1!
1*
b11 6
19
1>
1C
b11 G
#366840000000
0!
0*
09
0>
0C
#366850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#366860000000
0!
0*
09
0>
0C
#366870000000
1!
1*
b101 6
19
1>
1C
b101 G
#366880000000
0!
0*
09
0>
0C
#366890000000
1!
1*
b110 6
19
1>
1C
b110 G
#366900000000
0!
0*
09
0>
0C
#366910000000
1!
1*
b111 6
19
1>
1C
b111 G
#366920000000
0!
0*
09
0>
0C
#366930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#366940000000
0!
0*
09
0>
0C
#366950000000
1!
1*
b1 6
19
1>
1C
b1 G
#366960000000
0!
0*
09
0>
0C
#366970000000
1!
1*
b10 6
19
1>
1C
b10 G
#366980000000
0!
0*
09
0>
0C
#366990000000
1!
1*
b11 6
19
1>
1C
b11 G
#367000000000
0!
0*
09
0>
0C
#367010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#367020000000
0!
0*
09
0>
0C
#367030000000
1!
1*
b101 6
19
1>
1C
b101 G
#367040000000
0!
0*
09
0>
0C
#367050000000
1!
1*
b110 6
19
1>
1C
b110 G
#367060000000
0!
0*
09
0>
0C
#367070000000
1!
1*
b111 6
19
1>
1C
b111 G
#367080000000
0!
0*
09
0>
0C
#367090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#367100000000
0!
0*
09
0>
0C
#367110000000
1!
1*
b1 6
19
1>
1C
b1 G
#367120000000
0!
0*
09
0>
0C
#367130000000
1!
1*
b10 6
19
1>
1C
b10 G
#367140000000
0!
0*
09
0>
0C
#367150000000
1!
1*
b11 6
19
1>
1C
b11 G
#367160000000
0!
0*
09
0>
0C
#367170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#367180000000
0!
0*
09
0>
0C
#367190000000
1!
1*
b101 6
19
1>
1C
b101 G
#367200000000
0!
0*
09
0>
0C
#367210000000
1!
1*
b110 6
19
1>
1C
b110 G
#367220000000
0!
0*
09
0>
0C
#367230000000
1!
1*
b111 6
19
1>
1C
b111 G
#367240000000
0!
1"
0*
1+
09
1:
0>
0C
#367250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#367260000000
0!
0*
09
0>
0C
#367270000000
1!
1*
b1 6
19
1>
1C
b1 G
#367280000000
0!
0*
09
0>
0C
#367290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#367300000000
0!
0*
09
0>
0C
#367310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#367320000000
0!
0*
09
0>
0C
#367330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#367340000000
0!
0*
09
0>
0C
#367350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#367360000000
0!
0#
0*
0,
09
0>
0?
0C
#367370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#367380000000
0!
0*
09
0>
0C
#367390000000
1!
1*
19
1>
1C
#367400000000
0!
0*
09
0>
0C
#367410000000
1!
1*
19
1>
1C
#367420000000
0!
0*
09
0>
0C
#367430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#367440000000
0!
0*
09
0>
0C
#367450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#367460000000
0!
0*
09
0>
0C
#367470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#367480000000
0!
0*
09
0>
0C
#367490000000
1!
1*
b10 6
19
1>
1C
b10 G
#367500000000
0!
0*
09
0>
0C
#367510000000
1!
1*
b11 6
19
1>
1C
b11 G
#367520000000
0!
0*
09
0>
0C
#367530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#367540000000
0!
0*
09
0>
0C
#367550000000
1!
1*
b101 6
19
1>
1C
b101 G
#367560000000
0!
0*
09
0>
0C
#367570000000
1!
1*
b110 6
19
1>
1C
b110 G
#367580000000
0!
0*
09
0>
0C
#367590000000
1!
1*
b111 6
19
1>
1C
b111 G
#367600000000
0!
0*
09
0>
0C
#367610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#367620000000
0!
0*
09
0>
0C
#367630000000
1!
1*
b1 6
19
1>
1C
b1 G
#367640000000
0!
0*
09
0>
0C
#367650000000
1!
1*
b10 6
19
1>
1C
b10 G
#367660000000
0!
0*
09
0>
0C
#367670000000
1!
1*
b11 6
19
1>
1C
b11 G
#367680000000
0!
0*
09
0>
0C
#367690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#367700000000
0!
0*
09
0>
0C
#367710000000
1!
1*
b101 6
19
1>
1C
b101 G
#367720000000
0!
0*
09
0>
0C
#367730000000
1!
1*
b110 6
19
1>
1C
b110 G
#367740000000
0!
0*
09
0>
0C
#367750000000
1!
1*
b111 6
19
1>
1C
b111 G
#367760000000
0!
0*
09
0>
0C
#367770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#367780000000
0!
0*
09
0>
0C
#367790000000
1!
1*
b1 6
19
1>
1C
b1 G
#367800000000
0!
0*
09
0>
0C
#367810000000
1!
1*
b10 6
19
1>
1C
b10 G
#367820000000
0!
0*
09
0>
0C
#367830000000
1!
1*
b11 6
19
1>
1C
b11 G
#367840000000
0!
0*
09
0>
0C
#367850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#367860000000
0!
0*
09
0>
0C
#367870000000
1!
1*
b101 6
19
1>
1C
b101 G
#367880000000
0!
0*
09
0>
0C
#367890000000
1!
1*
b110 6
19
1>
1C
b110 G
#367900000000
0!
0*
09
0>
0C
#367910000000
1!
1*
b111 6
19
1>
1C
b111 G
#367920000000
0!
1"
0*
1+
09
1:
0>
0C
#367930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#367940000000
0!
0*
09
0>
0C
#367950000000
1!
1*
b1 6
19
1>
1C
b1 G
#367960000000
0!
0*
09
0>
0C
#367970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#367980000000
0!
0*
09
0>
0C
#367990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#368000000000
0!
0*
09
0>
0C
#368010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#368020000000
0!
0*
09
0>
0C
#368030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#368040000000
0!
0#
0*
0,
09
0>
0?
0C
#368050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#368060000000
0!
0*
09
0>
0C
#368070000000
1!
1*
19
1>
1C
#368080000000
0!
0*
09
0>
0C
#368090000000
1!
1*
19
1>
1C
#368100000000
0!
0*
09
0>
0C
#368110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#368120000000
0!
0*
09
0>
0C
#368130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#368140000000
0!
0*
09
0>
0C
#368150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#368160000000
0!
0*
09
0>
0C
#368170000000
1!
1*
b10 6
19
1>
1C
b10 G
#368180000000
0!
0*
09
0>
0C
#368190000000
1!
1*
b11 6
19
1>
1C
b11 G
#368200000000
0!
0*
09
0>
0C
#368210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#368220000000
0!
0*
09
0>
0C
#368230000000
1!
1*
b101 6
19
1>
1C
b101 G
#368240000000
0!
0*
09
0>
0C
#368250000000
1!
1*
b110 6
19
1>
1C
b110 G
#368260000000
0!
0*
09
0>
0C
#368270000000
1!
1*
b111 6
19
1>
1C
b111 G
#368280000000
0!
0*
09
0>
0C
#368290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#368300000000
0!
0*
09
0>
0C
#368310000000
1!
1*
b1 6
19
1>
1C
b1 G
#368320000000
0!
0*
09
0>
0C
#368330000000
1!
1*
b10 6
19
1>
1C
b10 G
#368340000000
0!
0*
09
0>
0C
#368350000000
1!
1*
b11 6
19
1>
1C
b11 G
#368360000000
0!
0*
09
0>
0C
#368370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#368380000000
0!
0*
09
0>
0C
#368390000000
1!
1*
b101 6
19
1>
1C
b101 G
#368400000000
0!
0*
09
0>
0C
#368410000000
1!
1*
b110 6
19
1>
1C
b110 G
#368420000000
0!
0*
09
0>
0C
#368430000000
1!
1*
b111 6
19
1>
1C
b111 G
#368440000000
0!
0*
09
0>
0C
#368450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#368460000000
0!
0*
09
0>
0C
#368470000000
1!
1*
b1 6
19
1>
1C
b1 G
#368480000000
0!
0*
09
0>
0C
#368490000000
1!
1*
b10 6
19
1>
1C
b10 G
#368500000000
0!
0*
09
0>
0C
#368510000000
1!
1*
b11 6
19
1>
1C
b11 G
#368520000000
0!
0*
09
0>
0C
#368530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#368540000000
0!
0*
09
0>
0C
#368550000000
1!
1*
b101 6
19
1>
1C
b101 G
#368560000000
0!
0*
09
0>
0C
#368570000000
1!
1*
b110 6
19
1>
1C
b110 G
#368580000000
0!
0*
09
0>
0C
#368590000000
1!
1*
b111 6
19
1>
1C
b111 G
#368600000000
0!
1"
0*
1+
09
1:
0>
0C
#368610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#368620000000
0!
0*
09
0>
0C
#368630000000
1!
1*
b1 6
19
1>
1C
b1 G
#368640000000
0!
0*
09
0>
0C
#368650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#368660000000
0!
0*
09
0>
0C
#368670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#368680000000
0!
0*
09
0>
0C
#368690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#368700000000
0!
0*
09
0>
0C
#368710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#368720000000
0!
0#
0*
0,
09
0>
0?
0C
#368730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#368740000000
0!
0*
09
0>
0C
#368750000000
1!
1*
19
1>
1C
#368760000000
0!
0*
09
0>
0C
#368770000000
1!
1*
19
1>
1C
#368780000000
0!
0*
09
0>
0C
#368790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#368800000000
0!
0*
09
0>
0C
#368810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#368820000000
0!
0*
09
0>
0C
#368830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#368840000000
0!
0*
09
0>
0C
#368850000000
1!
1*
b10 6
19
1>
1C
b10 G
#368860000000
0!
0*
09
0>
0C
#368870000000
1!
1*
b11 6
19
1>
1C
b11 G
#368880000000
0!
0*
09
0>
0C
#368890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#368900000000
0!
0*
09
0>
0C
#368910000000
1!
1*
b101 6
19
1>
1C
b101 G
#368920000000
0!
0*
09
0>
0C
#368930000000
1!
1*
b110 6
19
1>
1C
b110 G
#368940000000
0!
0*
09
0>
0C
#368950000000
1!
1*
b111 6
19
1>
1C
b111 G
#368960000000
0!
0*
09
0>
0C
#368970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#368980000000
0!
0*
09
0>
0C
#368990000000
1!
1*
b1 6
19
1>
1C
b1 G
#369000000000
0!
0*
09
0>
0C
#369010000000
1!
1*
b10 6
19
1>
1C
b10 G
#369020000000
0!
0*
09
0>
0C
#369030000000
1!
1*
b11 6
19
1>
1C
b11 G
#369040000000
0!
0*
09
0>
0C
#369050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#369060000000
0!
0*
09
0>
0C
#369070000000
1!
1*
b101 6
19
1>
1C
b101 G
#369080000000
0!
0*
09
0>
0C
#369090000000
1!
1*
b110 6
19
1>
1C
b110 G
#369100000000
0!
0*
09
0>
0C
#369110000000
1!
1*
b111 6
19
1>
1C
b111 G
#369120000000
0!
0*
09
0>
0C
#369130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#369140000000
0!
0*
09
0>
0C
#369150000000
1!
1*
b1 6
19
1>
1C
b1 G
#369160000000
0!
0*
09
0>
0C
#369170000000
1!
1*
b10 6
19
1>
1C
b10 G
#369180000000
0!
0*
09
0>
0C
#369190000000
1!
1*
b11 6
19
1>
1C
b11 G
#369200000000
0!
0*
09
0>
0C
#369210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#369220000000
0!
0*
09
0>
0C
#369230000000
1!
1*
b101 6
19
1>
1C
b101 G
#369240000000
0!
0*
09
0>
0C
#369250000000
1!
1*
b110 6
19
1>
1C
b110 G
#369260000000
0!
0*
09
0>
0C
#369270000000
1!
1*
b111 6
19
1>
1C
b111 G
#369280000000
0!
1"
0*
1+
09
1:
0>
0C
#369290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#369300000000
0!
0*
09
0>
0C
#369310000000
1!
1*
b1 6
19
1>
1C
b1 G
#369320000000
0!
0*
09
0>
0C
#369330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#369340000000
0!
0*
09
0>
0C
#369350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#369360000000
0!
0*
09
0>
0C
#369370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#369380000000
0!
0*
09
0>
0C
#369390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#369400000000
0!
0#
0*
0,
09
0>
0?
0C
#369410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#369420000000
0!
0*
09
0>
0C
#369430000000
1!
1*
19
1>
1C
#369440000000
0!
0*
09
0>
0C
#369450000000
1!
1*
19
1>
1C
#369460000000
0!
0*
09
0>
0C
#369470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#369480000000
0!
0*
09
0>
0C
#369490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#369500000000
0!
0*
09
0>
0C
#369510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#369520000000
0!
0*
09
0>
0C
#369530000000
1!
1*
b10 6
19
1>
1C
b10 G
#369540000000
0!
0*
09
0>
0C
#369550000000
1!
1*
b11 6
19
1>
1C
b11 G
#369560000000
0!
0*
09
0>
0C
#369570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#369580000000
0!
0*
09
0>
0C
#369590000000
1!
1*
b101 6
19
1>
1C
b101 G
#369600000000
0!
0*
09
0>
0C
#369610000000
1!
1*
b110 6
19
1>
1C
b110 G
#369620000000
0!
0*
09
0>
0C
#369630000000
1!
1*
b111 6
19
1>
1C
b111 G
#369640000000
0!
0*
09
0>
0C
#369650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#369660000000
0!
0*
09
0>
0C
#369670000000
1!
1*
b1 6
19
1>
1C
b1 G
#369680000000
0!
0*
09
0>
0C
#369690000000
1!
1*
b10 6
19
1>
1C
b10 G
#369700000000
0!
0*
09
0>
0C
#369710000000
1!
1*
b11 6
19
1>
1C
b11 G
#369720000000
0!
0*
09
0>
0C
#369730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#369740000000
0!
0*
09
0>
0C
#369750000000
1!
1*
b101 6
19
1>
1C
b101 G
#369760000000
0!
0*
09
0>
0C
#369770000000
1!
1*
b110 6
19
1>
1C
b110 G
#369780000000
0!
0*
09
0>
0C
#369790000000
1!
1*
b111 6
19
1>
1C
b111 G
#369800000000
0!
0*
09
0>
0C
#369810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#369820000000
0!
0*
09
0>
0C
#369830000000
1!
1*
b1 6
19
1>
1C
b1 G
#369840000000
0!
0*
09
0>
0C
#369850000000
1!
1*
b10 6
19
1>
1C
b10 G
#369860000000
0!
0*
09
0>
0C
#369870000000
1!
1*
b11 6
19
1>
1C
b11 G
#369880000000
0!
0*
09
0>
0C
#369890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#369900000000
0!
0*
09
0>
0C
#369910000000
1!
1*
b101 6
19
1>
1C
b101 G
#369920000000
0!
0*
09
0>
0C
#369930000000
1!
1*
b110 6
19
1>
1C
b110 G
#369940000000
0!
0*
09
0>
0C
#369950000000
1!
1*
b111 6
19
1>
1C
b111 G
#369960000000
0!
1"
0*
1+
09
1:
0>
0C
#369970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#369980000000
0!
0*
09
0>
0C
#369990000000
1!
1*
b1 6
19
1>
1C
b1 G
#370000000000
0!
0*
09
0>
0C
#370010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#370020000000
0!
0*
09
0>
0C
#370030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#370040000000
0!
0*
09
0>
0C
#370050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#370060000000
0!
0*
09
0>
0C
#370070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#370080000000
0!
0#
0*
0,
09
0>
0?
0C
#370090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#370100000000
0!
0*
09
0>
0C
#370110000000
1!
1*
19
1>
1C
#370120000000
0!
0*
09
0>
0C
#370130000000
1!
1*
19
1>
1C
#370140000000
0!
0*
09
0>
0C
#370150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#370160000000
0!
0*
09
0>
0C
#370170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#370180000000
0!
0*
09
0>
0C
#370190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#370200000000
0!
0*
09
0>
0C
#370210000000
1!
1*
b10 6
19
1>
1C
b10 G
#370220000000
0!
0*
09
0>
0C
#370230000000
1!
1*
b11 6
19
1>
1C
b11 G
#370240000000
0!
0*
09
0>
0C
#370250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#370260000000
0!
0*
09
0>
0C
#370270000000
1!
1*
b101 6
19
1>
1C
b101 G
#370280000000
0!
0*
09
0>
0C
#370290000000
1!
1*
b110 6
19
1>
1C
b110 G
#370300000000
0!
0*
09
0>
0C
#370310000000
1!
1*
b111 6
19
1>
1C
b111 G
#370320000000
0!
0*
09
0>
0C
#370330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#370340000000
0!
0*
09
0>
0C
#370350000000
1!
1*
b1 6
19
1>
1C
b1 G
#370360000000
0!
0*
09
0>
0C
#370370000000
1!
1*
b10 6
19
1>
1C
b10 G
#370380000000
0!
0*
09
0>
0C
#370390000000
1!
1*
b11 6
19
1>
1C
b11 G
#370400000000
0!
0*
09
0>
0C
#370410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#370420000000
0!
0*
09
0>
0C
#370430000000
1!
1*
b101 6
19
1>
1C
b101 G
#370440000000
0!
0*
09
0>
0C
#370450000000
1!
1*
b110 6
19
1>
1C
b110 G
#370460000000
0!
0*
09
0>
0C
#370470000000
1!
1*
b111 6
19
1>
1C
b111 G
#370480000000
0!
0*
09
0>
0C
#370490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#370500000000
0!
0*
09
0>
0C
#370510000000
1!
1*
b1 6
19
1>
1C
b1 G
#370520000000
0!
0*
09
0>
0C
#370530000000
1!
1*
b10 6
19
1>
1C
b10 G
#370540000000
0!
0*
09
0>
0C
#370550000000
1!
1*
b11 6
19
1>
1C
b11 G
#370560000000
0!
0*
09
0>
0C
#370570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#370580000000
0!
0*
09
0>
0C
#370590000000
1!
1*
b101 6
19
1>
1C
b101 G
#370600000000
0!
0*
09
0>
0C
#370610000000
1!
1*
b110 6
19
1>
1C
b110 G
#370620000000
0!
0*
09
0>
0C
#370630000000
1!
1*
b111 6
19
1>
1C
b111 G
#370640000000
0!
1"
0*
1+
09
1:
0>
0C
#370650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#370660000000
0!
0*
09
0>
0C
#370670000000
1!
1*
b1 6
19
1>
1C
b1 G
#370680000000
0!
0*
09
0>
0C
#370690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#370700000000
0!
0*
09
0>
0C
#370710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#370720000000
0!
0*
09
0>
0C
#370730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#370740000000
0!
0*
09
0>
0C
#370750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#370760000000
0!
0#
0*
0,
09
0>
0?
0C
#370770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#370780000000
0!
0*
09
0>
0C
#370790000000
1!
1*
19
1>
1C
#370800000000
0!
0*
09
0>
0C
#370810000000
1!
1*
19
1>
1C
#370820000000
0!
0*
09
0>
0C
#370830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#370840000000
0!
0*
09
0>
0C
#370850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#370860000000
0!
0*
09
0>
0C
#370870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#370880000000
0!
0*
09
0>
0C
#370890000000
1!
1*
b10 6
19
1>
1C
b10 G
#370900000000
0!
0*
09
0>
0C
#370910000000
1!
1*
b11 6
19
1>
1C
b11 G
#370920000000
0!
0*
09
0>
0C
#370930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#370940000000
0!
0*
09
0>
0C
#370950000000
1!
1*
b101 6
19
1>
1C
b101 G
#370960000000
0!
0*
09
0>
0C
#370970000000
1!
1*
b110 6
19
1>
1C
b110 G
#370980000000
0!
0*
09
0>
0C
#370990000000
1!
1*
b111 6
19
1>
1C
b111 G
#371000000000
0!
0*
09
0>
0C
#371010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#371020000000
0!
0*
09
0>
0C
#371030000000
1!
1*
b1 6
19
1>
1C
b1 G
#371040000000
0!
0*
09
0>
0C
#371050000000
1!
1*
b10 6
19
1>
1C
b10 G
#371060000000
0!
0*
09
0>
0C
#371070000000
1!
1*
b11 6
19
1>
1C
b11 G
#371080000000
0!
0*
09
0>
0C
#371090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#371100000000
0!
0*
09
0>
0C
#371110000000
1!
1*
b101 6
19
1>
1C
b101 G
#371120000000
0!
0*
09
0>
0C
#371130000000
1!
1*
b110 6
19
1>
1C
b110 G
#371140000000
0!
0*
09
0>
0C
#371150000000
1!
1*
b111 6
19
1>
1C
b111 G
#371160000000
0!
0*
09
0>
0C
#371170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#371180000000
0!
0*
09
0>
0C
#371190000000
1!
1*
b1 6
19
1>
1C
b1 G
#371200000000
0!
0*
09
0>
0C
#371210000000
1!
1*
b10 6
19
1>
1C
b10 G
#371220000000
0!
0*
09
0>
0C
#371230000000
1!
1*
b11 6
19
1>
1C
b11 G
#371240000000
0!
0*
09
0>
0C
#371250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#371260000000
0!
0*
09
0>
0C
#371270000000
1!
1*
b101 6
19
1>
1C
b101 G
#371280000000
0!
0*
09
0>
0C
#371290000000
1!
1*
b110 6
19
1>
1C
b110 G
#371300000000
0!
0*
09
0>
0C
#371310000000
1!
1*
b111 6
19
1>
1C
b111 G
#371320000000
0!
1"
0*
1+
09
1:
0>
0C
#371330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#371340000000
0!
0*
09
0>
0C
#371350000000
1!
1*
b1 6
19
1>
1C
b1 G
#371360000000
0!
0*
09
0>
0C
#371370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#371380000000
0!
0*
09
0>
0C
#371390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#371400000000
0!
0*
09
0>
0C
#371410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#371420000000
0!
0*
09
0>
0C
#371430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#371440000000
0!
0#
0*
0,
09
0>
0?
0C
#371450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#371460000000
0!
0*
09
0>
0C
#371470000000
1!
1*
19
1>
1C
#371480000000
0!
0*
09
0>
0C
#371490000000
1!
1*
19
1>
1C
#371500000000
0!
0*
09
0>
0C
#371510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#371520000000
0!
0*
09
0>
0C
#371530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#371540000000
0!
0*
09
0>
0C
#371550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#371560000000
0!
0*
09
0>
0C
#371570000000
1!
1*
b10 6
19
1>
1C
b10 G
#371580000000
0!
0*
09
0>
0C
#371590000000
1!
1*
b11 6
19
1>
1C
b11 G
#371600000000
0!
0*
09
0>
0C
#371610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#371620000000
0!
0*
09
0>
0C
#371630000000
1!
1*
b101 6
19
1>
1C
b101 G
#371640000000
0!
0*
09
0>
0C
#371650000000
1!
1*
b110 6
19
1>
1C
b110 G
#371660000000
0!
0*
09
0>
0C
#371670000000
1!
1*
b111 6
19
1>
1C
b111 G
#371680000000
0!
0*
09
0>
0C
#371690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#371700000000
0!
0*
09
0>
0C
#371710000000
1!
1*
b1 6
19
1>
1C
b1 G
#371720000000
0!
0*
09
0>
0C
#371730000000
1!
1*
b10 6
19
1>
1C
b10 G
#371740000000
0!
0*
09
0>
0C
#371750000000
1!
1*
b11 6
19
1>
1C
b11 G
#371760000000
0!
0*
09
0>
0C
#371770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#371780000000
0!
0*
09
0>
0C
#371790000000
1!
1*
b101 6
19
1>
1C
b101 G
#371800000000
0!
0*
09
0>
0C
#371810000000
1!
1*
b110 6
19
1>
1C
b110 G
#371820000000
0!
0*
09
0>
0C
#371830000000
1!
1*
b111 6
19
1>
1C
b111 G
#371840000000
0!
0*
09
0>
0C
#371850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#371860000000
0!
0*
09
0>
0C
#371870000000
1!
1*
b1 6
19
1>
1C
b1 G
#371880000000
0!
0*
09
0>
0C
#371890000000
1!
1*
b10 6
19
1>
1C
b10 G
#371900000000
0!
0*
09
0>
0C
#371910000000
1!
1*
b11 6
19
1>
1C
b11 G
#371920000000
0!
0*
09
0>
0C
#371930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#371940000000
0!
0*
09
0>
0C
#371950000000
1!
1*
b101 6
19
1>
1C
b101 G
#371960000000
0!
0*
09
0>
0C
#371970000000
1!
1*
b110 6
19
1>
1C
b110 G
#371980000000
0!
0*
09
0>
0C
#371990000000
1!
1*
b111 6
19
1>
1C
b111 G
#372000000000
0!
1"
0*
1+
09
1:
0>
0C
#372010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#372020000000
0!
0*
09
0>
0C
#372030000000
1!
1*
b1 6
19
1>
1C
b1 G
#372040000000
0!
0*
09
0>
0C
#372050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#372060000000
0!
0*
09
0>
0C
#372070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#372080000000
0!
0*
09
0>
0C
#372090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#372100000000
0!
0*
09
0>
0C
#372110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#372120000000
0!
0#
0*
0,
09
0>
0?
0C
#372130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#372140000000
0!
0*
09
0>
0C
#372150000000
1!
1*
19
1>
1C
#372160000000
0!
0*
09
0>
0C
#372170000000
1!
1*
19
1>
1C
#372180000000
0!
0*
09
0>
0C
#372190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#372200000000
0!
0*
09
0>
0C
#372210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#372220000000
0!
0*
09
0>
0C
#372230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#372240000000
0!
0*
09
0>
0C
#372250000000
1!
1*
b10 6
19
1>
1C
b10 G
#372260000000
0!
0*
09
0>
0C
#372270000000
1!
1*
b11 6
19
1>
1C
b11 G
#372280000000
0!
0*
09
0>
0C
#372290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#372300000000
0!
0*
09
0>
0C
#372310000000
1!
1*
b101 6
19
1>
1C
b101 G
#372320000000
0!
0*
09
0>
0C
#372330000000
1!
1*
b110 6
19
1>
1C
b110 G
#372340000000
0!
0*
09
0>
0C
#372350000000
1!
1*
b111 6
19
1>
1C
b111 G
#372360000000
0!
0*
09
0>
0C
#372370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#372380000000
0!
0*
09
0>
0C
#372390000000
1!
1*
b1 6
19
1>
1C
b1 G
#372400000000
0!
0*
09
0>
0C
#372410000000
1!
1*
b10 6
19
1>
1C
b10 G
#372420000000
0!
0*
09
0>
0C
#372430000000
1!
1*
b11 6
19
1>
1C
b11 G
#372440000000
0!
0*
09
0>
0C
#372450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#372460000000
0!
0*
09
0>
0C
#372470000000
1!
1*
b101 6
19
1>
1C
b101 G
#372480000000
0!
0*
09
0>
0C
#372490000000
1!
1*
b110 6
19
1>
1C
b110 G
#372500000000
0!
0*
09
0>
0C
#372510000000
1!
1*
b111 6
19
1>
1C
b111 G
#372520000000
0!
0*
09
0>
0C
#372530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#372540000000
0!
0*
09
0>
0C
#372550000000
1!
1*
b1 6
19
1>
1C
b1 G
#372560000000
0!
0*
09
0>
0C
#372570000000
1!
1*
b10 6
19
1>
1C
b10 G
#372580000000
0!
0*
09
0>
0C
#372590000000
1!
1*
b11 6
19
1>
1C
b11 G
#372600000000
0!
0*
09
0>
0C
#372610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#372620000000
0!
0*
09
0>
0C
#372630000000
1!
1*
b101 6
19
1>
1C
b101 G
#372640000000
0!
0*
09
0>
0C
#372650000000
1!
1*
b110 6
19
1>
1C
b110 G
#372660000000
0!
0*
09
0>
0C
#372670000000
1!
1*
b111 6
19
1>
1C
b111 G
#372680000000
0!
1"
0*
1+
09
1:
0>
0C
#372690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#372700000000
0!
0*
09
0>
0C
#372710000000
1!
1*
b1 6
19
1>
1C
b1 G
#372720000000
0!
0*
09
0>
0C
#372730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#372740000000
0!
0*
09
0>
0C
#372750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#372760000000
0!
0*
09
0>
0C
#372770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#372780000000
0!
0*
09
0>
0C
#372790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#372800000000
0!
0#
0*
0,
09
0>
0?
0C
#372810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#372820000000
0!
0*
09
0>
0C
#372830000000
1!
1*
19
1>
1C
#372840000000
0!
0*
09
0>
0C
#372850000000
1!
1*
19
1>
1C
#372860000000
0!
0*
09
0>
0C
#372870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#372880000000
0!
0*
09
0>
0C
#372890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#372900000000
0!
0*
09
0>
0C
#372910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#372920000000
0!
0*
09
0>
0C
#372930000000
1!
1*
b10 6
19
1>
1C
b10 G
#372940000000
0!
0*
09
0>
0C
#372950000000
1!
1*
b11 6
19
1>
1C
b11 G
#372960000000
0!
0*
09
0>
0C
#372970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#372980000000
0!
0*
09
0>
0C
#372990000000
1!
1*
b101 6
19
1>
1C
b101 G
#373000000000
0!
0*
09
0>
0C
#373010000000
1!
1*
b110 6
19
1>
1C
b110 G
#373020000000
0!
0*
09
0>
0C
#373030000000
1!
1*
b111 6
19
1>
1C
b111 G
#373040000000
0!
0*
09
0>
0C
#373050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#373060000000
0!
0*
09
0>
0C
#373070000000
1!
1*
b1 6
19
1>
1C
b1 G
#373080000000
0!
0*
09
0>
0C
#373090000000
1!
1*
b10 6
19
1>
1C
b10 G
#373100000000
0!
0*
09
0>
0C
#373110000000
1!
1*
b11 6
19
1>
1C
b11 G
#373120000000
0!
0*
09
0>
0C
#373130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#373140000000
0!
0*
09
0>
0C
#373150000000
1!
1*
b101 6
19
1>
1C
b101 G
#373160000000
0!
0*
09
0>
0C
#373170000000
1!
1*
b110 6
19
1>
1C
b110 G
#373180000000
0!
0*
09
0>
0C
#373190000000
1!
1*
b111 6
19
1>
1C
b111 G
#373200000000
0!
0*
09
0>
0C
#373210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#373220000000
0!
0*
09
0>
0C
#373230000000
1!
1*
b1 6
19
1>
1C
b1 G
#373240000000
0!
0*
09
0>
0C
#373250000000
1!
1*
b10 6
19
1>
1C
b10 G
#373260000000
0!
0*
09
0>
0C
#373270000000
1!
1*
b11 6
19
1>
1C
b11 G
#373280000000
0!
0*
09
0>
0C
#373290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#373300000000
0!
0*
09
0>
0C
#373310000000
1!
1*
b101 6
19
1>
1C
b101 G
#373320000000
0!
0*
09
0>
0C
#373330000000
1!
1*
b110 6
19
1>
1C
b110 G
#373340000000
0!
0*
09
0>
0C
#373350000000
1!
1*
b111 6
19
1>
1C
b111 G
#373360000000
0!
1"
0*
1+
09
1:
0>
0C
#373370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#373380000000
0!
0*
09
0>
0C
#373390000000
1!
1*
b1 6
19
1>
1C
b1 G
#373400000000
0!
0*
09
0>
0C
#373410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#373420000000
0!
0*
09
0>
0C
#373430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#373440000000
0!
0*
09
0>
0C
#373450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#373460000000
0!
0*
09
0>
0C
#373470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#373480000000
0!
0#
0*
0,
09
0>
0?
0C
#373490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#373500000000
0!
0*
09
0>
0C
#373510000000
1!
1*
19
1>
1C
#373520000000
0!
0*
09
0>
0C
#373530000000
1!
1*
19
1>
1C
#373540000000
0!
0*
09
0>
0C
#373550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#373560000000
0!
0*
09
0>
0C
#373570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#373580000000
0!
0*
09
0>
0C
#373590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#373600000000
0!
0*
09
0>
0C
#373610000000
1!
1*
b10 6
19
1>
1C
b10 G
#373620000000
0!
0*
09
0>
0C
#373630000000
1!
1*
b11 6
19
1>
1C
b11 G
#373640000000
0!
0*
09
0>
0C
#373650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#373660000000
0!
0*
09
0>
0C
#373670000000
1!
1*
b101 6
19
1>
1C
b101 G
#373680000000
0!
0*
09
0>
0C
#373690000000
1!
1*
b110 6
19
1>
1C
b110 G
#373700000000
0!
0*
09
0>
0C
#373710000000
1!
1*
b111 6
19
1>
1C
b111 G
#373720000000
0!
0*
09
0>
0C
#373730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#373740000000
0!
0*
09
0>
0C
#373750000000
1!
1*
b1 6
19
1>
1C
b1 G
#373760000000
0!
0*
09
0>
0C
#373770000000
1!
1*
b10 6
19
1>
1C
b10 G
#373780000000
0!
0*
09
0>
0C
#373790000000
1!
1*
b11 6
19
1>
1C
b11 G
#373800000000
0!
0*
09
0>
0C
#373810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#373820000000
0!
0*
09
0>
0C
#373830000000
1!
1*
b101 6
19
1>
1C
b101 G
#373840000000
0!
0*
09
0>
0C
#373850000000
1!
1*
b110 6
19
1>
1C
b110 G
#373860000000
0!
0*
09
0>
0C
#373870000000
1!
1*
b111 6
19
1>
1C
b111 G
#373880000000
0!
0*
09
0>
0C
#373890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#373900000000
0!
0*
09
0>
0C
#373910000000
1!
1*
b1 6
19
1>
1C
b1 G
#373920000000
0!
0*
09
0>
0C
#373930000000
1!
1*
b10 6
19
1>
1C
b10 G
#373940000000
0!
0*
09
0>
0C
#373950000000
1!
1*
b11 6
19
1>
1C
b11 G
#373960000000
0!
0*
09
0>
0C
#373970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#373980000000
0!
0*
09
0>
0C
#373990000000
1!
1*
b101 6
19
1>
1C
b101 G
#374000000000
0!
0*
09
0>
0C
#374010000000
1!
1*
b110 6
19
1>
1C
b110 G
#374020000000
0!
0*
09
0>
0C
#374030000000
1!
1*
b111 6
19
1>
1C
b111 G
#374040000000
0!
1"
0*
1+
09
1:
0>
0C
#374050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#374060000000
0!
0*
09
0>
0C
#374070000000
1!
1*
b1 6
19
1>
1C
b1 G
#374080000000
0!
0*
09
0>
0C
#374090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#374100000000
0!
0*
09
0>
0C
#374110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#374120000000
0!
0*
09
0>
0C
#374130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#374140000000
0!
0*
09
0>
0C
#374150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#374160000000
0!
0#
0*
0,
09
0>
0?
0C
#374170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#374180000000
0!
0*
09
0>
0C
#374190000000
1!
1*
19
1>
1C
#374200000000
0!
0*
09
0>
0C
#374210000000
1!
1*
19
1>
1C
#374220000000
0!
0*
09
0>
0C
#374230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#374240000000
0!
0*
09
0>
0C
#374250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#374260000000
0!
0*
09
0>
0C
#374270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#374280000000
0!
0*
09
0>
0C
#374290000000
1!
1*
b10 6
19
1>
1C
b10 G
#374300000000
0!
0*
09
0>
0C
#374310000000
1!
1*
b11 6
19
1>
1C
b11 G
#374320000000
0!
0*
09
0>
0C
#374330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#374340000000
0!
0*
09
0>
0C
#374350000000
1!
1*
b101 6
19
1>
1C
b101 G
#374360000000
0!
0*
09
0>
0C
#374370000000
1!
1*
b110 6
19
1>
1C
b110 G
#374380000000
0!
0*
09
0>
0C
#374390000000
1!
1*
b111 6
19
1>
1C
b111 G
#374400000000
0!
0*
09
0>
0C
#374410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#374420000000
0!
0*
09
0>
0C
#374430000000
1!
1*
b1 6
19
1>
1C
b1 G
#374440000000
0!
0*
09
0>
0C
#374450000000
1!
1*
b10 6
19
1>
1C
b10 G
#374460000000
0!
0*
09
0>
0C
#374470000000
1!
1*
b11 6
19
1>
1C
b11 G
#374480000000
0!
0*
09
0>
0C
#374490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#374500000000
0!
0*
09
0>
0C
#374510000000
1!
1*
b101 6
19
1>
1C
b101 G
#374520000000
0!
0*
09
0>
0C
#374530000000
1!
1*
b110 6
19
1>
1C
b110 G
#374540000000
0!
0*
09
0>
0C
#374550000000
1!
1*
b111 6
19
1>
1C
b111 G
#374560000000
0!
0*
09
0>
0C
#374570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#374580000000
0!
0*
09
0>
0C
#374590000000
1!
1*
b1 6
19
1>
1C
b1 G
#374600000000
0!
0*
09
0>
0C
#374610000000
1!
1*
b10 6
19
1>
1C
b10 G
#374620000000
0!
0*
09
0>
0C
#374630000000
1!
1*
b11 6
19
1>
1C
b11 G
#374640000000
0!
0*
09
0>
0C
#374650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#374660000000
0!
0*
09
0>
0C
#374670000000
1!
1*
b101 6
19
1>
1C
b101 G
#374680000000
0!
0*
09
0>
0C
#374690000000
1!
1*
b110 6
19
1>
1C
b110 G
#374700000000
0!
0*
09
0>
0C
#374710000000
1!
1*
b111 6
19
1>
1C
b111 G
#374720000000
0!
1"
0*
1+
09
1:
0>
0C
#374730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#374740000000
0!
0*
09
0>
0C
#374750000000
1!
1*
b1 6
19
1>
1C
b1 G
#374760000000
0!
0*
09
0>
0C
#374770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#374780000000
0!
0*
09
0>
0C
#374790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#374800000000
0!
0*
09
0>
0C
#374810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#374820000000
0!
0*
09
0>
0C
#374830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#374840000000
0!
0#
0*
0,
09
0>
0?
0C
#374850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#374860000000
0!
0*
09
0>
0C
#374870000000
1!
1*
19
1>
1C
#374880000000
0!
0*
09
0>
0C
#374890000000
1!
1*
19
1>
1C
#374900000000
0!
0*
09
0>
0C
#374910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#374920000000
0!
0*
09
0>
0C
#374930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#374940000000
0!
0*
09
0>
0C
#374950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#374960000000
0!
0*
09
0>
0C
#374970000000
1!
1*
b10 6
19
1>
1C
b10 G
#374980000000
0!
0*
09
0>
0C
#374990000000
1!
1*
b11 6
19
1>
1C
b11 G
#375000000000
0!
0*
09
0>
0C
#375010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#375020000000
0!
0*
09
0>
0C
#375030000000
1!
1*
b101 6
19
1>
1C
b101 G
#375040000000
0!
0*
09
0>
0C
#375050000000
1!
1*
b110 6
19
1>
1C
b110 G
#375060000000
0!
0*
09
0>
0C
#375070000000
1!
1*
b111 6
19
1>
1C
b111 G
#375080000000
0!
0*
09
0>
0C
#375090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#375100000000
0!
0*
09
0>
0C
#375110000000
1!
1*
b1 6
19
1>
1C
b1 G
#375120000000
0!
0*
09
0>
0C
#375130000000
1!
1*
b10 6
19
1>
1C
b10 G
#375140000000
0!
0*
09
0>
0C
#375150000000
1!
1*
b11 6
19
1>
1C
b11 G
#375160000000
0!
0*
09
0>
0C
#375170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#375180000000
0!
0*
09
0>
0C
#375190000000
1!
1*
b101 6
19
1>
1C
b101 G
#375200000000
0!
0*
09
0>
0C
#375210000000
1!
1*
b110 6
19
1>
1C
b110 G
#375220000000
0!
0*
09
0>
0C
#375230000000
1!
1*
b111 6
19
1>
1C
b111 G
#375240000000
0!
0*
09
0>
0C
#375250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#375260000000
0!
0*
09
0>
0C
#375270000000
1!
1*
b1 6
19
1>
1C
b1 G
#375280000000
0!
0*
09
0>
0C
#375290000000
1!
1*
b10 6
19
1>
1C
b10 G
#375300000000
0!
0*
09
0>
0C
#375310000000
1!
1*
b11 6
19
1>
1C
b11 G
#375320000000
0!
0*
09
0>
0C
#375330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#375340000000
0!
0*
09
0>
0C
#375350000000
1!
1*
b101 6
19
1>
1C
b101 G
#375360000000
0!
0*
09
0>
0C
#375370000000
1!
1*
b110 6
19
1>
1C
b110 G
#375380000000
0!
0*
09
0>
0C
#375390000000
1!
1*
b111 6
19
1>
1C
b111 G
#375400000000
0!
1"
0*
1+
09
1:
0>
0C
#375410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#375420000000
0!
0*
09
0>
0C
#375430000000
1!
1*
b1 6
19
1>
1C
b1 G
#375440000000
0!
0*
09
0>
0C
#375450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#375460000000
0!
0*
09
0>
0C
#375470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#375480000000
0!
0*
09
0>
0C
#375490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#375500000000
0!
0*
09
0>
0C
#375510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#375520000000
0!
0#
0*
0,
09
0>
0?
0C
#375530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#375540000000
0!
0*
09
0>
0C
#375550000000
1!
1*
19
1>
1C
#375560000000
0!
0*
09
0>
0C
#375570000000
1!
1*
19
1>
1C
#375580000000
0!
0*
09
0>
0C
#375590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#375600000000
0!
0*
09
0>
0C
#375610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#375620000000
0!
0*
09
0>
0C
#375630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#375640000000
0!
0*
09
0>
0C
#375650000000
1!
1*
b10 6
19
1>
1C
b10 G
#375660000000
0!
0*
09
0>
0C
#375670000000
1!
1*
b11 6
19
1>
1C
b11 G
#375680000000
0!
0*
09
0>
0C
#375690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#375700000000
0!
0*
09
0>
0C
#375710000000
1!
1*
b101 6
19
1>
1C
b101 G
#375720000000
0!
0*
09
0>
0C
#375730000000
1!
1*
b110 6
19
1>
1C
b110 G
#375740000000
0!
0*
09
0>
0C
#375750000000
1!
1*
b111 6
19
1>
1C
b111 G
#375760000000
0!
0*
09
0>
0C
#375770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#375780000000
0!
0*
09
0>
0C
#375790000000
1!
1*
b1 6
19
1>
1C
b1 G
#375800000000
0!
0*
09
0>
0C
#375810000000
1!
1*
b10 6
19
1>
1C
b10 G
#375820000000
0!
0*
09
0>
0C
#375830000000
1!
1*
b11 6
19
1>
1C
b11 G
#375840000000
0!
0*
09
0>
0C
#375850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#375860000000
0!
0*
09
0>
0C
#375870000000
1!
1*
b101 6
19
1>
1C
b101 G
#375880000000
0!
0*
09
0>
0C
#375890000000
1!
1*
b110 6
19
1>
1C
b110 G
#375900000000
0!
0*
09
0>
0C
#375910000000
1!
1*
b111 6
19
1>
1C
b111 G
#375920000000
0!
0*
09
0>
0C
#375930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#375940000000
0!
0*
09
0>
0C
#375950000000
1!
1*
b1 6
19
1>
1C
b1 G
#375960000000
0!
0*
09
0>
0C
#375970000000
1!
1*
b10 6
19
1>
1C
b10 G
#375980000000
0!
0*
09
0>
0C
#375990000000
1!
1*
b11 6
19
1>
1C
b11 G
#376000000000
0!
0*
09
0>
0C
#376010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#376020000000
0!
0*
09
0>
0C
#376030000000
1!
1*
b101 6
19
1>
1C
b101 G
#376040000000
0!
0*
09
0>
0C
#376050000000
1!
1*
b110 6
19
1>
1C
b110 G
#376060000000
0!
0*
09
0>
0C
#376070000000
1!
1*
b111 6
19
1>
1C
b111 G
#376080000000
0!
1"
0*
1+
09
1:
0>
0C
#376090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#376100000000
0!
0*
09
0>
0C
#376110000000
1!
1*
b1 6
19
1>
1C
b1 G
#376120000000
0!
0*
09
0>
0C
#376130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#376140000000
0!
0*
09
0>
0C
#376150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#376160000000
0!
0*
09
0>
0C
#376170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#376180000000
0!
0*
09
0>
0C
#376190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#376200000000
0!
0#
0*
0,
09
0>
0?
0C
#376210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#376220000000
0!
0*
09
0>
0C
#376230000000
1!
1*
19
1>
1C
#376240000000
0!
0*
09
0>
0C
#376250000000
1!
1*
19
1>
1C
#376260000000
0!
0*
09
0>
0C
#376270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#376280000000
0!
0*
09
0>
0C
#376290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#376300000000
0!
0*
09
0>
0C
#376310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#376320000000
0!
0*
09
0>
0C
#376330000000
1!
1*
b10 6
19
1>
1C
b10 G
#376340000000
0!
0*
09
0>
0C
#376350000000
1!
1*
b11 6
19
1>
1C
b11 G
#376360000000
0!
0*
09
0>
0C
#376370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#376380000000
0!
0*
09
0>
0C
#376390000000
1!
1*
b101 6
19
1>
1C
b101 G
#376400000000
0!
0*
09
0>
0C
#376410000000
1!
1*
b110 6
19
1>
1C
b110 G
#376420000000
0!
0*
09
0>
0C
#376430000000
1!
1*
b111 6
19
1>
1C
b111 G
#376440000000
0!
0*
09
0>
0C
#376450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#376460000000
0!
0*
09
0>
0C
#376470000000
1!
1*
b1 6
19
1>
1C
b1 G
#376480000000
0!
0*
09
0>
0C
#376490000000
1!
1*
b10 6
19
1>
1C
b10 G
#376500000000
0!
0*
09
0>
0C
#376510000000
1!
1*
b11 6
19
1>
1C
b11 G
#376520000000
0!
0*
09
0>
0C
#376530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#376540000000
0!
0*
09
0>
0C
#376550000000
1!
1*
b101 6
19
1>
1C
b101 G
#376560000000
0!
0*
09
0>
0C
#376570000000
1!
1*
b110 6
19
1>
1C
b110 G
#376580000000
0!
0*
09
0>
0C
#376590000000
1!
1*
b111 6
19
1>
1C
b111 G
#376600000000
0!
0*
09
0>
0C
#376610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#376620000000
0!
0*
09
0>
0C
#376630000000
1!
1*
b1 6
19
1>
1C
b1 G
#376640000000
0!
0*
09
0>
0C
#376650000000
1!
1*
b10 6
19
1>
1C
b10 G
#376660000000
0!
0*
09
0>
0C
#376670000000
1!
1*
b11 6
19
1>
1C
b11 G
#376680000000
0!
0*
09
0>
0C
#376690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#376700000000
0!
0*
09
0>
0C
#376710000000
1!
1*
b101 6
19
1>
1C
b101 G
#376720000000
0!
0*
09
0>
0C
#376730000000
1!
1*
b110 6
19
1>
1C
b110 G
#376740000000
0!
0*
09
0>
0C
#376750000000
1!
1*
b111 6
19
1>
1C
b111 G
#376760000000
0!
1"
0*
1+
09
1:
0>
0C
#376770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#376780000000
0!
0*
09
0>
0C
#376790000000
1!
1*
b1 6
19
1>
1C
b1 G
#376800000000
0!
0*
09
0>
0C
#376810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#376820000000
0!
0*
09
0>
0C
#376830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#376840000000
0!
0*
09
0>
0C
#376850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#376860000000
0!
0*
09
0>
0C
#376870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#376880000000
0!
0#
0*
0,
09
0>
0?
0C
#376890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#376900000000
0!
0*
09
0>
0C
#376910000000
1!
1*
19
1>
1C
#376920000000
0!
0*
09
0>
0C
#376930000000
1!
1*
19
1>
1C
#376940000000
0!
0*
09
0>
0C
#376950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#376960000000
0!
0*
09
0>
0C
#376970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#376980000000
0!
0*
09
0>
0C
#376990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#377000000000
0!
0*
09
0>
0C
#377010000000
1!
1*
b10 6
19
1>
1C
b10 G
#377020000000
0!
0*
09
0>
0C
#377030000000
1!
1*
b11 6
19
1>
1C
b11 G
#377040000000
0!
0*
09
0>
0C
#377050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#377060000000
0!
0*
09
0>
0C
#377070000000
1!
1*
b101 6
19
1>
1C
b101 G
#377080000000
0!
0*
09
0>
0C
#377090000000
1!
1*
b110 6
19
1>
1C
b110 G
#377100000000
0!
0*
09
0>
0C
#377110000000
1!
1*
b111 6
19
1>
1C
b111 G
#377120000000
0!
0*
09
0>
0C
#377130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#377140000000
0!
0*
09
0>
0C
#377150000000
1!
1*
b1 6
19
1>
1C
b1 G
#377160000000
0!
0*
09
0>
0C
#377170000000
1!
1*
b10 6
19
1>
1C
b10 G
#377180000000
0!
0*
09
0>
0C
#377190000000
1!
1*
b11 6
19
1>
1C
b11 G
#377200000000
0!
0*
09
0>
0C
#377210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#377220000000
0!
0*
09
0>
0C
#377230000000
1!
1*
b101 6
19
1>
1C
b101 G
#377240000000
0!
0*
09
0>
0C
#377250000000
1!
1*
b110 6
19
1>
1C
b110 G
#377260000000
0!
0*
09
0>
0C
#377270000000
1!
1*
b111 6
19
1>
1C
b111 G
#377280000000
0!
0*
09
0>
0C
#377290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#377300000000
0!
0*
09
0>
0C
#377310000000
1!
1*
b1 6
19
1>
1C
b1 G
#377320000000
0!
0*
09
0>
0C
#377330000000
1!
1*
b10 6
19
1>
1C
b10 G
#377340000000
0!
0*
09
0>
0C
#377350000000
1!
1*
b11 6
19
1>
1C
b11 G
#377360000000
0!
0*
09
0>
0C
#377370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#377380000000
0!
0*
09
0>
0C
#377390000000
1!
1*
b101 6
19
1>
1C
b101 G
#377400000000
0!
0*
09
0>
0C
#377410000000
1!
1*
b110 6
19
1>
1C
b110 G
#377420000000
0!
0*
09
0>
0C
#377430000000
1!
1*
b111 6
19
1>
1C
b111 G
#377440000000
0!
1"
0*
1+
09
1:
0>
0C
#377450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#377460000000
0!
0*
09
0>
0C
#377470000000
1!
1*
b1 6
19
1>
1C
b1 G
#377480000000
0!
0*
09
0>
0C
#377490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#377500000000
0!
0*
09
0>
0C
#377510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#377520000000
0!
0*
09
0>
0C
#377530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#377540000000
0!
0*
09
0>
0C
#377550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#377560000000
0!
0#
0*
0,
09
0>
0?
0C
#377570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#377580000000
0!
0*
09
0>
0C
#377590000000
1!
1*
19
1>
1C
#377600000000
0!
0*
09
0>
0C
#377610000000
1!
1*
19
1>
1C
#377620000000
0!
0*
09
0>
0C
#377630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#377640000000
0!
0*
09
0>
0C
#377650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#377660000000
0!
0*
09
0>
0C
#377670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#377680000000
0!
0*
09
0>
0C
#377690000000
1!
1*
b10 6
19
1>
1C
b10 G
#377700000000
0!
0*
09
0>
0C
#377710000000
1!
1*
b11 6
19
1>
1C
b11 G
#377720000000
0!
0*
09
0>
0C
#377730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#377740000000
0!
0*
09
0>
0C
#377750000000
1!
1*
b101 6
19
1>
1C
b101 G
#377760000000
0!
0*
09
0>
0C
#377770000000
1!
1*
b110 6
19
1>
1C
b110 G
#377780000000
0!
0*
09
0>
0C
#377790000000
1!
1*
b111 6
19
1>
1C
b111 G
#377800000000
0!
0*
09
0>
0C
#377810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#377820000000
0!
0*
09
0>
0C
#377830000000
1!
1*
b1 6
19
1>
1C
b1 G
#377840000000
0!
0*
09
0>
0C
#377850000000
1!
1*
b10 6
19
1>
1C
b10 G
#377860000000
0!
0*
09
0>
0C
#377870000000
1!
1*
b11 6
19
1>
1C
b11 G
#377880000000
0!
0*
09
0>
0C
#377890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#377900000000
0!
0*
09
0>
0C
#377910000000
1!
1*
b101 6
19
1>
1C
b101 G
#377920000000
0!
0*
09
0>
0C
#377930000000
1!
1*
b110 6
19
1>
1C
b110 G
#377940000000
0!
0*
09
0>
0C
#377950000000
1!
1*
b111 6
19
1>
1C
b111 G
#377960000000
0!
0*
09
0>
0C
#377970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#377980000000
0!
0*
09
0>
0C
#377990000000
1!
1*
b1 6
19
1>
1C
b1 G
#378000000000
0!
0*
09
0>
0C
#378010000000
1!
1*
b10 6
19
1>
1C
b10 G
#378020000000
0!
0*
09
0>
0C
#378030000000
1!
1*
b11 6
19
1>
1C
b11 G
#378040000000
0!
0*
09
0>
0C
#378050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#378060000000
0!
0*
09
0>
0C
#378070000000
1!
1*
b101 6
19
1>
1C
b101 G
#378080000000
0!
0*
09
0>
0C
#378090000000
1!
1*
b110 6
19
1>
1C
b110 G
#378100000000
0!
0*
09
0>
0C
#378110000000
1!
1*
b111 6
19
1>
1C
b111 G
#378120000000
0!
1"
0*
1+
09
1:
0>
0C
#378130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#378140000000
0!
0*
09
0>
0C
#378150000000
1!
1*
b1 6
19
1>
1C
b1 G
#378160000000
0!
0*
09
0>
0C
#378170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#378180000000
0!
0*
09
0>
0C
#378190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#378200000000
0!
0*
09
0>
0C
#378210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#378220000000
0!
0*
09
0>
0C
#378230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#378240000000
0!
0#
0*
0,
09
0>
0?
0C
#378250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#378260000000
0!
0*
09
0>
0C
#378270000000
1!
1*
19
1>
1C
#378280000000
0!
0*
09
0>
0C
#378290000000
1!
1*
19
1>
1C
#378300000000
0!
0*
09
0>
0C
#378310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#378320000000
0!
0*
09
0>
0C
#378330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#378340000000
0!
0*
09
0>
0C
#378350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#378360000000
0!
0*
09
0>
0C
#378370000000
1!
1*
b10 6
19
1>
1C
b10 G
#378380000000
0!
0*
09
0>
0C
#378390000000
1!
1*
b11 6
19
1>
1C
b11 G
#378400000000
0!
0*
09
0>
0C
#378410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#378420000000
0!
0*
09
0>
0C
#378430000000
1!
1*
b101 6
19
1>
1C
b101 G
#378440000000
0!
0*
09
0>
0C
#378450000000
1!
1*
b110 6
19
1>
1C
b110 G
#378460000000
0!
0*
09
0>
0C
#378470000000
1!
1*
b111 6
19
1>
1C
b111 G
#378480000000
0!
0*
09
0>
0C
#378490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#378500000000
0!
0*
09
0>
0C
#378510000000
1!
1*
b1 6
19
1>
1C
b1 G
#378520000000
0!
0*
09
0>
0C
#378530000000
1!
1*
b10 6
19
1>
1C
b10 G
#378540000000
0!
0*
09
0>
0C
#378550000000
1!
1*
b11 6
19
1>
1C
b11 G
#378560000000
0!
0*
09
0>
0C
#378570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#378580000000
0!
0*
09
0>
0C
#378590000000
1!
1*
b101 6
19
1>
1C
b101 G
#378600000000
0!
0*
09
0>
0C
#378610000000
1!
1*
b110 6
19
1>
1C
b110 G
#378620000000
0!
0*
09
0>
0C
#378630000000
1!
1*
b111 6
19
1>
1C
b111 G
#378640000000
0!
0*
09
0>
0C
#378650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#378660000000
0!
0*
09
0>
0C
#378670000000
1!
1*
b1 6
19
1>
1C
b1 G
#378680000000
0!
0*
09
0>
0C
#378690000000
1!
1*
b10 6
19
1>
1C
b10 G
#378700000000
0!
0*
09
0>
0C
#378710000000
1!
1*
b11 6
19
1>
1C
b11 G
#378720000000
0!
0*
09
0>
0C
#378730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#378740000000
0!
0*
09
0>
0C
#378750000000
1!
1*
b101 6
19
1>
1C
b101 G
#378760000000
0!
0*
09
0>
0C
#378770000000
1!
1*
b110 6
19
1>
1C
b110 G
#378780000000
0!
0*
09
0>
0C
#378790000000
1!
1*
b111 6
19
1>
1C
b111 G
#378800000000
0!
1"
0*
1+
09
1:
0>
0C
#378810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#378820000000
0!
0*
09
0>
0C
#378830000000
1!
1*
b1 6
19
1>
1C
b1 G
#378840000000
0!
0*
09
0>
0C
#378850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#378860000000
0!
0*
09
0>
0C
#378870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#378880000000
0!
0*
09
0>
0C
#378890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#378900000000
0!
0*
09
0>
0C
#378910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#378920000000
0!
0#
0*
0,
09
0>
0?
0C
#378930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#378940000000
0!
0*
09
0>
0C
#378950000000
1!
1*
19
1>
1C
#378960000000
0!
0*
09
0>
0C
#378970000000
1!
1*
19
1>
1C
#378980000000
0!
0*
09
0>
0C
#378990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#379000000000
0!
0*
09
0>
0C
#379010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#379020000000
0!
0*
09
0>
0C
#379030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#379040000000
0!
0*
09
0>
0C
#379050000000
1!
1*
b10 6
19
1>
1C
b10 G
#379060000000
0!
0*
09
0>
0C
#379070000000
1!
1*
b11 6
19
1>
1C
b11 G
#379080000000
0!
0*
09
0>
0C
#379090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#379100000000
0!
0*
09
0>
0C
#379110000000
1!
1*
b101 6
19
1>
1C
b101 G
#379120000000
0!
0*
09
0>
0C
#379130000000
1!
1*
b110 6
19
1>
1C
b110 G
#379140000000
0!
0*
09
0>
0C
#379150000000
1!
1*
b111 6
19
1>
1C
b111 G
#379160000000
0!
0*
09
0>
0C
#379170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#379180000000
0!
0*
09
0>
0C
#379190000000
1!
1*
b1 6
19
1>
1C
b1 G
#379200000000
0!
0*
09
0>
0C
#379210000000
1!
1*
b10 6
19
1>
1C
b10 G
#379220000000
0!
0*
09
0>
0C
#379230000000
1!
1*
b11 6
19
1>
1C
b11 G
#379240000000
0!
0*
09
0>
0C
#379250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#379260000000
0!
0*
09
0>
0C
#379270000000
1!
1*
b101 6
19
1>
1C
b101 G
#379280000000
0!
0*
09
0>
0C
#379290000000
1!
1*
b110 6
19
1>
1C
b110 G
#379300000000
0!
0*
09
0>
0C
#379310000000
1!
1*
b111 6
19
1>
1C
b111 G
#379320000000
0!
0*
09
0>
0C
#379330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#379340000000
0!
0*
09
0>
0C
#379350000000
1!
1*
b1 6
19
1>
1C
b1 G
#379360000000
0!
0*
09
0>
0C
#379370000000
1!
1*
b10 6
19
1>
1C
b10 G
#379380000000
0!
0*
09
0>
0C
#379390000000
1!
1*
b11 6
19
1>
1C
b11 G
#379400000000
0!
0*
09
0>
0C
#379410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#379420000000
0!
0*
09
0>
0C
#379430000000
1!
1*
b101 6
19
1>
1C
b101 G
#379440000000
0!
0*
09
0>
0C
#379450000000
1!
1*
b110 6
19
1>
1C
b110 G
#379460000000
0!
0*
09
0>
0C
#379470000000
1!
1*
b111 6
19
1>
1C
b111 G
#379480000000
0!
1"
0*
1+
09
1:
0>
0C
#379490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#379500000000
0!
0*
09
0>
0C
#379510000000
1!
1*
b1 6
19
1>
1C
b1 G
#379520000000
0!
0*
09
0>
0C
#379530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#379540000000
0!
0*
09
0>
0C
#379550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#379560000000
0!
0*
09
0>
0C
#379570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#379580000000
0!
0*
09
0>
0C
#379590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#379600000000
0!
0#
0*
0,
09
0>
0?
0C
#379610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#379620000000
0!
0*
09
0>
0C
#379630000000
1!
1*
19
1>
1C
#379640000000
0!
0*
09
0>
0C
#379650000000
1!
1*
19
1>
1C
#379660000000
0!
0*
09
0>
0C
#379670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#379680000000
0!
0*
09
0>
0C
#379690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#379700000000
0!
0*
09
0>
0C
#379710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#379720000000
0!
0*
09
0>
0C
#379730000000
1!
1*
b10 6
19
1>
1C
b10 G
#379740000000
0!
0*
09
0>
0C
#379750000000
1!
1*
b11 6
19
1>
1C
b11 G
#379760000000
0!
0*
09
0>
0C
#379770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#379780000000
0!
0*
09
0>
0C
#379790000000
1!
1*
b101 6
19
1>
1C
b101 G
#379800000000
0!
0*
09
0>
0C
#379810000000
1!
1*
b110 6
19
1>
1C
b110 G
#379820000000
0!
0*
09
0>
0C
#379830000000
1!
1*
b111 6
19
1>
1C
b111 G
#379840000000
0!
0*
09
0>
0C
#379850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#379860000000
0!
0*
09
0>
0C
#379870000000
1!
1*
b1 6
19
1>
1C
b1 G
#379880000000
0!
0*
09
0>
0C
#379890000000
1!
1*
b10 6
19
1>
1C
b10 G
#379900000000
0!
0*
09
0>
0C
#379910000000
1!
1*
b11 6
19
1>
1C
b11 G
#379920000000
0!
0*
09
0>
0C
#379930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#379940000000
0!
0*
09
0>
0C
#379950000000
1!
1*
b101 6
19
1>
1C
b101 G
#379960000000
0!
0*
09
0>
0C
#379970000000
1!
1*
b110 6
19
1>
1C
b110 G
#379980000000
0!
0*
09
0>
0C
#379990000000
1!
1*
b111 6
19
1>
1C
b111 G
#380000000000
0!
0*
09
0>
0C
#380010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#380020000000
0!
0*
09
0>
0C
#380030000000
1!
1*
b1 6
19
1>
1C
b1 G
#380040000000
0!
0*
09
0>
0C
#380050000000
1!
1*
b10 6
19
1>
1C
b10 G
#380060000000
0!
0*
09
0>
0C
#380070000000
1!
1*
b11 6
19
1>
1C
b11 G
#380080000000
0!
0*
09
0>
0C
#380090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#380100000000
0!
0*
09
0>
0C
#380110000000
1!
1*
b101 6
19
1>
1C
b101 G
#380120000000
0!
0*
09
0>
0C
#380130000000
1!
1*
b110 6
19
1>
1C
b110 G
#380140000000
0!
0*
09
0>
0C
#380150000000
1!
1*
b111 6
19
1>
1C
b111 G
#380160000000
0!
1"
0*
1+
09
1:
0>
0C
#380170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#380180000000
0!
0*
09
0>
0C
#380190000000
1!
1*
b1 6
19
1>
1C
b1 G
#380200000000
0!
0*
09
0>
0C
#380210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#380220000000
0!
0*
09
0>
0C
#380230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#380240000000
0!
0*
09
0>
0C
#380250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#380260000000
0!
0*
09
0>
0C
#380270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#380280000000
0!
0#
0*
0,
09
0>
0?
0C
#380290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#380300000000
0!
0*
09
0>
0C
#380310000000
1!
1*
19
1>
1C
#380320000000
0!
0*
09
0>
0C
#380330000000
1!
1*
19
1>
1C
#380340000000
0!
0*
09
0>
0C
#380350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#380360000000
0!
0*
09
0>
0C
#380370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#380380000000
0!
0*
09
0>
0C
#380390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#380400000000
0!
0*
09
0>
0C
#380410000000
1!
1*
b10 6
19
1>
1C
b10 G
#380420000000
0!
0*
09
0>
0C
#380430000000
1!
1*
b11 6
19
1>
1C
b11 G
#380440000000
0!
0*
09
0>
0C
#380450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#380460000000
0!
0*
09
0>
0C
#380470000000
1!
1*
b101 6
19
1>
1C
b101 G
#380480000000
0!
0*
09
0>
0C
#380490000000
1!
1*
b110 6
19
1>
1C
b110 G
#380500000000
0!
0*
09
0>
0C
#380510000000
1!
1*
b111 6
19
1>
1C
b111 G
#380520000000
0!
0*
09
0>
0C
#380530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#380540000000
0!
0*
09
0>
0C
#380550000000
1!
1*
b1 6
19
1>
1C
b1 G
#380560000000
0!
0*
09
0>
0C
#380570000000
1!
1*
b10 6
19
1>
1C
b10 G
#380580000000
0!
0*
09
0>
0C
#380590000000
1!
1*
b11 6
19
1>
1C
b11 G
#380600000000
0!
0*
09
0>
0C
#380610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#380620000000
0!
0*
09
0>
0C
#380630000000
1!
1*
b101 6
19
1>
1C
b101 G
#380640000000
0!
0*
09
0>
0C
#380650000000
1!
1*
b110 6
19
1>
1C
b110 G
#380660000000
0!
0*
09
0>
0C
#380670000000
1!
1*
b111 6
19
1>
1C
b111 G
#380680000000
0!
0*
09
0>
0C
#380690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#380700000000
0!
0*
09
0>
0C
#380710000000
1!
1*
b1 6
19
1>
1C
b1 G
#380720000000
0!
0*
09
0>
0C
#380730000000
1!
1*
b10 6
19
1>
1C
b10 G
#380740000000
0!
0*
09
0>
0C
#380750000000
1!
1*
b11 6
19
1>
1C
b11 G
#380760000000
0!
0*
09
0>
0C
#380770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#380780000000
0!
0*
09
0>
0C
#380790000000
1!
1*
b101 6
19
1>
1C
b101 G
#380800000000
0!
0*
09
0>
0C
#380810000000
1!
1*
b110 6
19
1>
1C
b110 G
#380820000000
0!
0*
09
0>
0C
#380830000000
1!
1*
b111 6
19
1>
1C
b111 G
#380840000000
0!
1"
0*
1+
09
1:
0>
0C
#380850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#380860000000
0!
0*
09
0>
0C
#380870000000
1!
1*
b1 6
19
1>
1C
b1 G
#380880000000
0!
0*
09
0>
0C
#380890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#380900000000
0!
0*
09
0>
0C
#380910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#380920000000
0!
0*
09
0>
0C
#380930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#380940000000
0!
0*
09
0>
0C
#380950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#380960000000
0!
0#
0*
0,
09
0>
0?
0C
#380970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#380980000000
0!
0*
09
0>
0C
#380990000000
1!
1*
19
1>
1C
#381000000000
0!
0*
09
0>
0C
#381010000000
1!
1*
19
1>
1C
#381020000000
0!
0*
09
0>
0C
#381030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#381040000000
0!
0*
09
0>
0C
#381050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#381060000000
0!
0*
09
0>
0C
#381070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#381080000000
0!
0*
09
0>
0C
#381090000000
1!
1*
b10 6
19
1>
1C
b10 G
#381100000000
0!
0*
09
0>
0C
#381110000000
1!
1*
b11 6
19
1>
1C
b11 G
#381120000000
0!
0*
09
0>
0C
#381130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#381140000000
0!
0*
09
0>
0C
#381150000000
1!
1*
b101 6
19
1>
1C
b101 G
#381160000000
0!
0*
09
0>
0C
#381170000000
1!
1*
b110 6
19
1>
1C
b110 G
#381180000000
0!
0*
09
0>
0C
#381190000000
1!
1*
b111 6
19
1>
1C
b111 G
#381200000000
0!
0*
09
0>
0C
#381210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#381220000000
0!
0*
09
0>
0C
#381230000000
1!
1*
b1 6
19
1>
1C
b1 G
#381240000000
0!
0*
09
0>
0C
#381250000000
1!
1*
b10 6
19
1>
1C
b10 G
#381260000000
0!
0*
09
0>
0C
#381270000000
1!
1*
b11 6
19
1>
1C
b11 G
#381280000000
0!
0*
09
0>
0C
#381290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#381300000000
0!
0*
09
0>
0C
#381310000000
1!
1*
b101 6
19
1>
1C
b101 G
#381320000000
0!
0*
09
0>
0C
#381330000000
1!
1*
b110 6
19
1>
1C
b110 G
#381340000000
0!
0*
09
0>
0C
#381350000000
1!
1*
b111 6
19
1>
1C
b111 G
#381360000000
0!
0*
09
0>
0C
#381370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#381380000000
0!
0*
09
0>
0C
#381390000000
1!
1*
b1 6
19
1>
1C
b1 G
#381400000000
0!
0*
09
0>
0C
#381410000000
1!
1*
b10 6
19
1>
1C
b10 G
#381420000000
0!
0*
09
0>
0C
#381430000000
1!
1*
b11 6
19
1>
1C
b11 G
#381440000000
0!
0*
09
0>
0C
#381450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#381460000000
0!
0*
09
0>
0C
#381470000000
1!
1*
b101 6
19
1>
1C
b101 G
#381480000000
0!
0*
09
0>
0C
#381490000000
1!
1*
b110 6
19
1>
1C
b110 G
#381500000000
0!
0*
09
0>
0C
#381510000000
1!
1*
b111 6
19
1>
1C
b111 G
#381520000000
0!
1"
0*
1+
09
1:
0>
0C
#381530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#381540000000
0!
0*
09
0>
0C
#381550000000
1!
1*
b1 6
19
1>
1C
b1 G
#381560000000
0!
0*
09
0>
0C
#381570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#381580000000
0!
0*
09
0>
0C
#381590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#381600000000
0!
0*
09
0>
0C
#381610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#381620000000
0!
0*
09
0>
0C
#381630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#381640000000
0!
0#
0*
0,
09
0>
0?
0C
#381650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#381660000000
0!
0*
09
0>
0C
#381670000000
1!
1*
19
1>
1C
#381680000000
0!
0*
09
0>
0C
#381690000000
1!
1*
19
1>
1C
#381700000000
0!
0*
09
0>
0C
#381710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#381720000000
0!
0*
09
0>
0C
#381730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#381740000000
0!
0*
09
0>
0C
#381750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#381760000000
0!
0*
09
0>
0C
#381770000000
1!
1*
b10 6
19
1>
1C
b10 G
#381780000000
0!
0*
09
0>
0C
#381790000000
1!
1*
b11 6
19
1>
1C
b11 G
#381800000000
0!
0*
09
0>
0C
#381810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#381820000000
0!
0*
09
0>
0C
#381830000000
1!
1*
b101 6
19
1>
1C
b101 G
#381840000000
0!
0*
09
0>
0C
#381850000000
1!
1*
b110 6
19
1>
1C
b110 G
#381860000000
0!
0*
09
0>
0C
#381870000000
1!
1*
b111 6
19
1>
1C
b111 G
#381880000000
0!
0*
09
0>
0C
#381890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#381900000000
0!
0*
09
0>
0C
#381910000000
1!
1*
b1 6
19
1>
1C
b1 G
#381920000000
0!
0*
09
0>
0C
#381930000000
1!
1*
b10 6
19
1>
1C
b10 G
#381940000000
0!
0*
09
0>
0C
#381950000000
1!
1*
b11 6
19
1>
1C
b11 G
#381960000000
0!
0*
09
0>
0C
#381970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#381980000000
0!
0*
09
0>
0C
#381990000000
1!
1*
b101 6
19
1>
1C
b101 G
#382000000000
0!
0*
09
0>
0C
#382010000000
1!
1*
b110 6
19
1>
1C
b110 G
#382020000000
0!
0*
09
0>
0C
#382030000000
1!
1*
b111 6
19
1>
1C
b111 G
#382040000000
0!
0*
09
0>
0C
#382050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#382060000000
0!
0*
09
0>
0C
#382070000000
1!
1*
b1 6
19
1>
1C
b1 G
#382080000000
0!
0*
09
0>
0C
#382090000000
1!
1*
b10 6
19
1>
1C
b10 G
#382100000000
0!
0*
09
0>
0C
#382110000000
1!
1*
b11 6
19
1>
1C
b11 G
#382120000000
0!
0*
09
0>
0C
#382130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#382140000000
0!
0*
09
0>
0C
#382150000000
1!
1*
b101 6
19
1>
1C
b101 G
#382160000000
0!
0*
09
0>
0C
#382170000000
1!
1*
b110 6
19
1>
1C
b110 G
#382180000000
0!
0*
09
0>
0C
#382190000000
1!
1*
b111 6
19
1>
1C
b111 G
#382200000000
0!
1"
0*
1+
09
1:
0>
0C
#382210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#382220000000
0!
0*
09
0>
0C
#382230000000
1!
1*
b1 6
19
1>
1C
b1 G
#382240000000
0!
0*
09
0>
0C
#382250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#382260000000
0!
0*
09
0>
0C
#382270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#382280000000
0!
0*
09
0>
0C
#382290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#382300000000
0!
0*
09
0>
0C
#382310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#382320000000
0!
0#
0*
0,
09
0>
0?
0C
#382330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#382340000000
0!
0*
09
0>
0C
#382350000000
1!
1*
19
1>
1C
#382360000000
0!
0*
09
0>
0C
#382370000000
1!
1*
19
1>
1C
#382380000000
0!
0*
09
0>
0C
#382390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#382400000000
0!
0*
09
0>
0C
#382410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#382420000000
0!
0*
09
0>
0C
#382430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#382440000000
0!
0*
09
0>
0C
#382450000000
1!
1*
b10 6
19
1>
1C
b10 G
#382460000000
0!
0*
09
0>
0C
#382470000000
1!
1*
b11 6
19
1>
1C
b11 G
#382480000000
0!
0*
09
0>
0C
#382490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#382500000000
0!
0*
09
0>
0C
#382510000000
1!
1*
b101 6
19
1>
1C
b101 G
#382520000000
0!
0*
09
0>
0C
#382530000000
1!
1*
b110 6
19
1>
1C
b110 G
#382540000000
0!
0*
09
0>
0C
#382550000000
1!
1*
b111 6
19
1>
1C
b111 G
#382560000000
0!
0*
09
0>
0C
#382570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#382580000000
0!
0*
09
0>
0C
#382590000000
1!
1*
b1 6
19
1>
1C
b1 G
#382600000000
0!
0*
09
0>
0C
#382610000000
1!
1*
b10 6
19
1>
1C
b10 G
#382620000000
0!
0*
09
0>
0C
#382630000000
1!
1*
b11 6
19
1>
1C
b11 G
#382640000000
0!
0*
09
0>
0C
#382650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#382660000000
0!
0*
09
0>
0C
#382670000000
1!
1*
b101 6
19
1>
1C
b101 G
#382680000000
0!
0*
09
0>
0C
#382690000000
1!
1*
b110 6
19
1>
1C
b110 G
#382700000000
0!
0*
09
0>
0C
#382710000000
1!
1*
b111 6
19
1>
1C
b111 G
#382720000000
0!
0*
09
0>
0C
#382730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#382740000000
0!
0*
09
0>
0C
#382750000000
1!
1*
b1 6
19
1>
1C
b1 G
#382760000000
0!
0*
09
0>
0C
#382770000000
1!
1*
b10 6
19
1>
1C
b10 G
#382780000000
0!
0*
09
0>
0C
#382790000000
1!
1*
b11 6
19
1>
1C
b11 G
#382800000000
0!
0*
09
0>
0C
#382810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#382820000000
0!
0*
09
0>
0C
#382830000000
1!
1*
b101 6
19
1>
1C
b101 G
#382840000000
0!
0*
09
0>
0C
#382850000000
1!
1*
b110 6
19
1>
1C
b110 G
#382860000000
0!
0*
09
0>
0C
#382870000000
1!
1*
b111 6
19
1>
1C
b111 G
#382880000000
0!
1"
0*
1+
09
1:
0>
0C
#382890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#382900000000
0!
0*
09
0>
0C
#382910000000
1!
1*
b1 6
19
1>
1C
b1 G
#382920000000
0!
0*
09
0>
0C
#382930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#382940000000
0!
0*
09
0>
0C
#382950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#382960000000
0!
0*
09
0>
0C
#382970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#382980000000
0!
0*
09
0>
0C
#382990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#383000000000
0!
0#
0*
0,
09
0>
0?
0C
#383010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#383020000000
0!
0*
09
0>
0C
#383030000000
1!
1*
19
1>
1C
#383040000000
0!
0*
09
0>
0C
#383050000000
1!
1*
19
1>
1C
#383060000000
0!
0*
09
0>
0C
#383070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#383080000000
0!
0*
09
0>
0C
#383090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#383100000000
0!
0*
09
0>
0C
#383110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#383120000000
0!
0*
09
0>
0C
#383130000000
1!
1*
b10 6
19
1>
1C
b10 G
#383140000000
0!
0*
09
0>
0C
#383150000000
1!
1*
b11 6
19
1>
1C
b11 G
#383160000000
0!
0*
09
0>
0C
#383170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#383180000000
0!
0*
09
0>
0C
#383190000000
1!
1*
b101 6
19
1>
1C
b101 G
#383200000000
0!
0*
09
0>
0C
#383210000000
1!
1*
b110 6
19
1>
1C
b110 G
#383220000000
0!
0*
09
0>
0C
#383230000000
1!
1*
b111 6
19
1>
1C
b111 G
#383240000000
0!
0*
09
0>
0C
#383250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#383260000000
0!
0*
09
0>
0C
#383270000000
1!
1*
b1 6
19
1>
1C
b1 G
#383280000000
0!
0*
09
0>
0C
#383290000000
1!
1*
b10 6
19
1>
1C
b10 G
#383300000000
0!
0*
09
0>
0C
#383310000000
1!
1*
b11 6
19
1>
1C
b11 G
#383320000000
0!
0*
09
0>
0C
#383330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#383340000000
0!
0*
09
0>
0C
#383350000000
1!
1*
b101 6
19
1>
1C
b101 G
#383360000000
0!
0*
09
0>
0C
#383370000000
1!
1*
b110 6
19
1>
1C
b110 G
#383380000000
0!
0*
09
0>
0C
#383390000000
1!
1*
b111 6
19
1>
1C
b111 G
#383400000000
0!
0*
09
0>
0C
#383410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#383420000000
0!
0*
09
0>
0C
#383430000000
1!
1*
b1 6
19
1>
1C
b1 G
#383440000000
0!
0*
09
0>
0C
#383450000000
1!
1*
b10 6
19
1>
1C
b10 G
#383460000000
0!
0*
09
0>
0C
#383470000000
1!
1*
b11 6
19
1>
1C
b11 G
#383480000000
0!
0*
09
0>
0C
#383490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#383500000000
0!
0*
09
0>
0C
#383510000000
1!
1*
b101 6
19
1>
1C
b101 G
#383520000000
0!
0*
09
0>
0C
#383530000000
1!
1*
b110 6
19
1>
1C
b110 G
#383540000000
0!
0*
09
0>
0C
#383550000000
1!
1*
b111 6
19
1>
1C
b111 G
#383560000000
0!
1"
0*
1+
09
1:
0>
0C
#383570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#383580000000
0!
0*
09
0>
0C
#383590000000
1!
1*
b1 6
19
1>
1C
b1 G
#383600000000
0!
0*
09
0>
0C
#383610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#383620000000
0!
0*
09
0>
0C
#383630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#383640000000
0!
0*
09
0>
0C
#383650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#383660000000
0!
0*
09
0>
0C
#383670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#383680000000
0!
0#
0*
0,
09
0>
0?
0C
#383690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#383700000000
0!
0*
09
0>
0C
#383710000000
1!
1*
19
1>
1C
#383720000000
0!
0*
09
0>
0C
#383730000000
1!
1*
19
1>
1C
#383740000000
0!
0*
09
0>
0C
#383750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#383760000000
0!
0*
09
0>
0C
#383770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#383780000000
0!
0*
09
0>
0C
#383790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#383800000000
0!
0*
09
0>
0C
#383810000000
1!
1*
b10 6
19
1>
1C
b10 G
#383820000000
0!
0*
09
0>
0C
#383830000000
1!
1*
b11 6
19
1>
1C
b11 G
#383840000000
0!
0*
09
0>
0C
#383850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#383860000000
0!
0*
09
0>
0C
#383870000000
1!
1*
b101 6
19
1>
1C
b101 G
#383880000000
0!
0*
09
0>
0C
#383890000000
1!
1*
b110 6
19
1>
1C
b110 G
#383900000000
0!
0*
09
0>
0C
#383910000000
1!
1*
b111 6
19
1>
1C
b111 G
#383920000000
0!
0*
09
0>
0C
#383930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#383940000000
0!
0*
09
0>
0C
#383950000000
1!
1*
b1 6
19
1>
1C
b1 G
#383960000000
0!
0*
09
0>
0C
#383970000000
1!
1*
b10 6
19
1>
1C
b10 G
#383980000000
0!
0*
09
0>
0C
#383990000000
1!
1*
b11 6
19
1>
1C
b11 G
#384000000000
0!
0*
09
0>
0C
#384010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#384020000000
0!
0*
09
0>
0C
#384030000000
1!
1*
b101 6
19
1>
1C
b101 G
#384040000000
0!
0*
09
0>
0C
#384050000000
1!
1*
b110 6
19
1>
1C
b110 G
#384060000000
0!
0*
09
0>
0C
#384070000000
1!
1*
b111 6
19
1>
1C
b111 G
#384080000000
0!
0*
09
0>
0C
#384090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#384100000000
0!
0*
09
0>
0C
#384110000000
1!
1*
b1 6
19
1>
1C
b1 G
#384120000000
0!
0*
09
0>
0C
#384130000000
1!
1*
b10 6
19
1>
1C
b10 G
#384140000000
0!
0*
09
0>
0C
#384150000000
1!
1*
b11 6
19
1>
1C
b11 G
#384160000000
0!
0*
09
0>
0C
#384170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#384180000000
0!
0*
09
0>
0C
#384190000000
1!
1*
b101 6
19
1>
1C
b101 G
#384200000000
0!
0*
09
0>
0C
#384210000000
1!
1*
b110 6
19
1>
1C
b110 G
#384220000000
0!
0*
09
0>
0C
#384230000000
1!
1*
b111 6
19
1>
1C
b111 G
#384240000000
0!
1"
0*
1+
09
1:
0>
0C
#384250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#384260000000
0!
0*
09
0>
0C
#384270000000
1!
1*
b1 6
19
1>
1C
b1 G
#384280000000
0!
0*
09
0>
0C
#384290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#384300000000
0!
0*
09
0>
0C
#384310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#384320000000
0!
0*
09
0>
0C
#384330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#384340000000
0!
0*
09
0>
0C
#384350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#384360000000
0!
0#
0*
0,
09
0>
0?
0C
#384370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#384380000000
0!
0*
09
0>
0C
#384390000000
1!
1*
19
1>
1C
#384400000000
0!
0*
09
0>
0C
#384410000000
1!
1*
19
1>
1C
#384420000000
0!
0*
09
0>
0C
#384430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#384440000000
0!
0*
09
0>
0C
#384450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#384460000000
0!
0*
09
0>
0C
#384470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#384480000000
0!
0*
09
0>
0C
#384490000000
1!
1*
b10 6
19
1>
1C
b10 G
#384500000000
0!
0*
09
0>
0C
#384510000000
1!
1*
b11 6
19
1>
1C
b11 G
#384520000000
0!
0*
09
0>
0C
#384530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#384540000000
0!
0*
09
0>
0C
#384550000000
1!
1*
b101 6
19
1>
1C
b101 G
#384560000000
0!
0*
09
0>
0C
#384570000000
1!
1*
b110 6
19
1>
1C
b110 G
#384580000000
0!
0*
09
0>
0C
#384590000000
1!
1*
b111 6
19
1>
1C
b111 G
#384600000000
0!
0*
09
0>
0C
#384610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#384620000000
0!
0*
09
0>
0C
#384630000000
1!
1*
b1 6
19
1>
1C
b1 G
#384640000000
0!
0*
09
0>
0C
#384650000000
1!
1*
b10 6
19
1>
1C
b10 G
#384660000000
0!
0*
09
0>
0C
#384670000000
1!
1*
b11 6
19
1>
1C
b11 G
#384680000000
0!
0*
09
0>
0C
#384690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#384700000000
0!
0*
09
0>
0C
#384710000000
1!
1*
b101 6
19
1>
1C
b101 G
#384720000000
0!
0*
09
0>
0C
#384730000000
1!
1*
b110 6
19
1>
1C
b110 G
#384740000000
0!
0*
09
0>
0C
#384750000000
1!
1*
b111 6
19
1>
1C
b111 G
#384760000000
0!
0*
09
0>
0C
#384770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#384780000000
0!
0*
09
0>
0C
#384790000000
1!
1*
b1 6
19
1>
1C
b1 G
#384800000000
0!
0*
09
0>
0C
#384810000000
1!
1*
b10 6
19
1>
1C
b10 G
#384820000000
0!
0*
09
0>
0C
#384830000000
1!
1*
b11 6
19
1>
1C
b11 G
#384840000000
0!
0*
09
0>
0C
#384850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#384860000000
0!
0*
09
0>
0C
#384870000000
1!
1*
b101 6
19
1>
1C
b101 G
#384880000000
0!
0*
09
0>
0C
#384890000000
1!
1*
b110 6
19
1>
1C
b110 G
#384900000000
0!
0*
09
0>
0C
#384910000000
1!
1*
b111 6
19
1>
1C
b111 G
#384920000000
0!
1"
0*
1+
09
1:
0>
0C
#384930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#384940000000
0!
0*
09
0>
0C
#384950000000
1!
1*
b1 6
19
1>
1C
b1 G
#384960000000
0!
0*
09
0>
0C
#384970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#384980000000
0!
0*
09
0>
0C
#384990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#385000000000
0!
0*
09
0>
0C
#385010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#385020000000
0!
0*
09
0>
0C
#385030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#385040000000
0!
0#
0*
0,
09
0>
0?
0C
#385050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#385060000000
0!
0*
09
0>
0C
#385070000000
1!
1*
19
1>
1C
#385080000000
0!
0*
09
0>
0C
#385090000000
1!
1*
19
1>
1C
#385100000000
0!
0*
09
0>
0C
#385110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#385120000000
0!
0*
09
0>
0C
#385130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#385140000000
0!
0*
09
0>
0C
#385150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#385160000000
0!
0*
09
0>
0C
#385170000000
1!
1*
b10 6
19
1>
1C
b10 G
#385180000000
0!
0*
09
0>
0C
#385190000000
1!
1*
b11 6
19
1>
1C
b11 G
#385200000000
0!
0*
09
0>
0C
#385210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#385220000000
0!
0*
09
0>
0C
#385230000000
1!
1*
b101 6
19
1>
1C
b101 G
#385240000000
0!
0*
09
0>
0C
#385250000000
1!
1*
b110 6
19
1>
1C
b110 G
#385260000000
0!
0*
09
0>
0C
#385270000000
1!
1*
b111 6
19
1>
1C
b111 G
#385280000000
0!
0*
09
0>
0C
#385290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#385300000000
0!
0*
09
0>
0C
#385310000000
1!
1*
b1 6
19
1>
1C
b1 G
#385320000000
0!
0*
09
0>
0C
#385330000000
1!
1*
b10 6
19
1>
1C
b10 G
#385340000000
0!
0*
09
0>
0C
#385350000000
1!
1*
b11 6
19
1>
1C
b11 G
#385360000000
0!
0*
09
0>
0C
#385370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#385380000000
0!
0*
09
0>
0C
#385390000000
1!
1*
b101 6
19
1>
1C
b101 G
#385400000000
0!
0*
09
0>
0C
#385410000000
1!
1*
b110 6
19
1>
1C
b110 G
#385420000000
0!
0*
09
0>
0C
#385430000000
1!
1*
b111 6
19
1>
1C
b111 G
#385440000000
0!
0*
09
0>
0C
#385450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#385460000000
0!
0*
09
0>
0C
#385470000000
1!
1*
b1 6
19
1>
1C
b1 G
#385480000000
0!
0*
09
0>
0C
#385490000000
1!
1*
b10 6
19
1>
1C
b10 G
#385500000000
0!
0*
09
0>
0C
#385510000000
1!
1*
b11 6
19
1>
1C
b11 G
#385520000000
0!
0*
09
0>
0C
#385530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#385540000000
0!
0*
09
0>
0C
#385550000000
1!
1*
b101 6
19
1>
1C
b101 G
#385560000000
0!
0*
09
0>
0C
#385570000000
1!
1*
b110 6
19
1>
1C
b110 G
#385580000000
0!
0*
09
0>
0C
#385590000000
1!
1*
b111 6
19
1>
1C
b111 G
#385600000000
0!
1"
0*
1+
09
1:
0>
0C
#385610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#385620000000
0!
0*
09
0>
0C
#385630000000
1!
1*
b1 6
19
1>
1C
b1 G
#385640000000
0!
0*
09
0>
0C
#385650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#385660000000
0!
0*
09
0>
0C
#385670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#385680000000
0!
0*
09
0>
0C
#385690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#385700000000
0!
0*
09
0>
0C
#385710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#385720000000
0!
0#
0*
0,
09
0>
0?
0C
#385730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#385740000000
0!
0*
09
0>
0C
#385750000000
1!
1*
19
1>
1C
#385760000000
0!
0*
09
0>
0C
#385770000000
1!
1*
19
1>
1C
#385780000000
0!
0*
09
0>
0C
#385790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#385800000000
0!
0*
09
0>
0C
#385810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#385820000000
0!
0*
09
0>
0C
#385830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#385840000000
0!
0*
09
0>
0C
#385850000000
1!
1*
b10 6
19
1>
1C
b10 G
#385860000000
0!
0*
09
0>
0C
#385870000000
1!
1*
b11 6
19
1>
1C
b11 G
#385880000000
0!
0*
09
0>
0C
#385890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#385900000000
0!
0*
09
0>
0C
#385910000000
1!
1*
b101 6
19
1>
1C
b101 G
#385920000000
0!
0*
09
0>
0C
#385930000000
1!
1*
b110 6
19
1>
1C
b110 G
#385940000000
0!
0*
09
0>
0C
#385950000000
1!
1*
b111 6
19
1>
1C
b111 G
#385960000000
0!
0*
09
0>
0C
#385970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#385980000000
0!
0*
09
0>
0C
#385990000000
1!
1*
b1 6
19
1>
1C
b1 G
#386000000000
0!
0*
09
0>
0C
#386010000000
1!
1*
b10 6
19
1>
1C
b10 G
#386020000000
0!
0*
09
0>
0C
#386030000000
1!
1*
b11 6
19
1>
1C
b11 G
#386040000000
0!
0*
09
0>
0C
#386050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#386060000000
0!
0*
09
0>
0C
#386070000000
1!
1*
b101 6
19
1>
1C
b101 G
#386080000000
0!
0*
09
0>
0C
#386090000000
1!
1*
b110 6
19
1>
1C
b110 G
#386100000000
0!
0*
09
0>
0C
#386110000000
1!
1*
b111 6
19
1>
1C
b111 G
#386120000000
0!
0*
09
0>
0C
#386130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#386140000000
0!
0*
09
0>
0C
#386150000000
1!
1*
b1 6
19
1>
1C
b1 G
#386160000000
0!
0*
09
0>
0C
#386170000000
1!
1*
b10 6
19
1>
1C
b10 G
#386180000000
0!
0*
09
0>
0C
#386190000000
1!
1*
b11 6
19
1>
1C
b11 G
#386200000000
0!
0*
09
0>
0C
#386210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#386220000000
0!
0*
09
0>
0C
#386230000000
1!
1*
b101 6
19
1>
1C
b101 G
#386240000000
0!
0*
09
0>
0C
#386250000000
1!
1*
b110 6
19
1>
1C
b110 G
#386260000000
0!
0*
09
0>
0C
#386270000000
1!
1*
b111 6
19
1>
1C
b111 G
#386280000000
0!
1"
0*
1+
09
1:
0>
0C
#386290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#386300000000
0!
0*
09
0>
0C
#386310000000
1!
1*
b1 6
19
1>
1C
b1 G
#386320000000
0!
0*
09
0>
0C
#386330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#386340000000
0!
0*
09
0>
0C
#386350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#386360000000
0!
0*
09
0>
0C
#386370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#386380000000
0!
0*
09
0>
0C
#386390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#386400000000
0!
0#
0*
0,
09
0>
0?
0C
#386410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#386420000000
0!
0*
09
0>
0C
#386430000000
1!
1*
19
1>
1C
#386440000000
0!
0*
09
0>
0C
#386450000000
1!
1*
19
1>
1C
#386460000000
0!
0*
09
0>
0C
#386470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#386480000000
0!
0*
09
0>
0C
#386490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#386500000000
0!
0*
09
0>
0C
#386510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#386520000000
0!
0*
09
0>
0C
#386530000000
1!
1*
b10 6
19
1>
1C
b10 G
#386540000000
0!
0*
09
0>
0C
#386550000000
1!
1*
b11 6
19
1>
1C
b11 G
#386560000000
0!
0*
09
0>
0C
#386570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#386580000000
0!
0*
09
0>
0C
#386590000000
1!
1*
b101 6
19
1>
1C
b101 G
#386600000000
0!
0*
09
0>
0C
#386610000000
1!
1*
b110 6
19
1>
1C
b110 G
#386620000000
0!
0*
09
0>
0C
#386630000000
1!
1*
b111 6
19
1>
1C
b111 G
#386640000000
0!
0*
09
0>
0C
#386650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#386660000000
0!
0*
09
0>
0C
#386670000000
1!
1*
b1 6
19
1>
1C
b1 G
#386680000000
0!
0*
09
0>
0C
#386690000000
1!
1*
b10 6
19
1>
1C
b10 G
#386700000000
0!
0*
09
0>
0C
#386710000000
1!
1*
b11 6
19
1>
1C
b11 G
#386720000000
0!
0*
09
0>
0C
#386730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#386740000000
0!
0*
09
0>
0C
#386750000000
1!
1*
b101 6
19
1>
1C
b101 G
#386760000000
0!
0*
09
0>
0C
#386770000000
1!
1*
b110 6
19
1>
1C
b110 G
#386780000000
0!
0*
09
0>
0C
#386790000000
1!
1*
b111 6
19
1>
1C
b111 G
#386800000000
0!
0*
09
0>
0C
#386810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#386820000000
0!
0*
09
0>
0C
#386830000000
1!
1*
b1 6
19
1>
1C
b1 G
#386840000000
0!
0*
09
0>
0C
#386850000000
1!
1*
b10 6
19
1>
1C
b10 G
#386860000000
0!
0*
09
0>
0C
#386870000000
1!
1*
b11 6
19
1>
1C
b11 G
#386880000000
0!
0*
09
0>
0C
#386890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#386900000000
0!
0*
09
0>
0C
#386910000000
1!
1*
b101 6
19
1>
1C
b101 G
#386920000000
0!
0*
09
0>
0C
#386930000000
1!
1*
b110 6
19
1>
1C
b110 G
#386940000000
0!
0*
09
0>
0C
#386950000000
1!
1*
b111 6
19
1>
1C
b111 G
#386960000000
0!
1"
0*
1+
09
1:
0>
0C
#386970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#386980000000
0!
0*
09
0>
0C
#386990000000
1!
1*
b1 6
19
1>
1C
b1 G
#387000000000
0!
0*
09
0>
0C
#387010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#387020000000
0!
0*
09
0>
0C
#387030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#387040000000
0!
0*
09
0>
0C
#387050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#387060000000
0!
0*
09
0>
0C
#387070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#387080000000
0!
0#
0*
0,
09
0>
0?
0C
#387090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#387100000000
0!
0*
09
0>
0C
#387110000000
1!
1*
19
1>
1C
#387120000000
0!
0*
09
0>
0C
#387130000000
1!
1*
19
1>
1C
#387140000000
0!
0*
09
0>
0C
#387150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#387160000000
0!
0*
09
0>
0C
#387170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#387180000000
0!
0*
09
0>
0C
#387190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#387200000000
0!
0*
09
0>
0C
#387210000000
1!
1*
b10 6
19
1>
1C
b10 G
#387220000000
0!
0*
09
0>
0C
#387230000000
1!
1*
b11 6
19
1>
1C
b11 G
#387240000000
0!
0*
09
0>
0C
#387250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#387260000000
0!
0*
09
0>
0C
#387270000000
1!
1*
b101 6
19
1>
1C
b101 G
#387280000000
0!
0*
09
0>
0C
#387290000000
1!
1*
b110 6
19
1>
1C
b110 G
#387300000000
0!
0*
09
0>
0C
#387310000000
1!
1*
b111 6
19
1>
1C
b111 G
#387320000000
0!
0*
09
0>
0C
#387330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#387340000000
0!
0*
09
0>
0C
#387350000000
1!
1*
b1 6
19
1>
1C
b1 G
#387360000000
0!
0*
09
0>
0C
#387370000000
1!
1*
b10 6
19
1>
1C
b10 G
#387380000000
0!
0*
09
0>
0C
#387390000000
1!
1*
b11 6
19
1>
1C
b11 G
#387400000000
0!
0*
09
0>
0C
#387410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#387420000000
0!
0*
09
0>
0C
#387430000000
1!
1*
b101 6
19
1>
1C
b101 G
#387440000000
0!
0*
09
0>
0C
#387450000000
1!
1*
b110 6
19
1>
1C
b110 G
#387460000000
0!
0*
09
0>
0C
#387470000000
1!
1*
b111 6
19
1>
1C
b111 G
#387480000000
0!
0*
09
0>
0C
#387490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#387500000000
0!
0*
09
0>
0C
#387510000000
1!
1*
b1 6
19
1>
1C
b1 G
#387520000000
0!
0*
09
0>
0C
#387530000000
1!
1*
b10 6
19
1>
1C
b10 G
#387540000000
0!
0*
09
0>
0C
#387550000000
1!
1*
b11 6
19
1>
1C
b11 G
#387560000000
0!
0*
09
0>
0C
#387570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#387580000000
0!
0*
09
0>
0C
#387590000000
1!
1*
b101 6
19
1>
1C
b101 G
#387600000000
0!
0*
09
0>
0C
#387610000000
1!
1*
b110 6
19
1>
1C
b110 G
#387620000000
0!
0*
09
0>
0C
#387630000000
1!
1*
b111 6
19
1>
1C
b111 G
#387640000000
0!
1"
0*
1+
09
1:
0>
0C
#387650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#387660000000
0!
0*
09
0>
0C
#387670000000
1!
1*
b1 6
19
1>
1C
b1 G
#387680000000
0!
0*
09
0>
0C
#387690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#387700000000
0!
0*
09
0>
0C
#387710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#387720000000
0!
0*
09
0>
0C
#387730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#387740000000
0!
0*
09
0>
0C
#387750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#387760000000
0!
0#
0*
0,
09
0>
0?
0C
#387770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#387780000000
0!
0*
09
0>
0C
#387790000000
1!
1*
19
1>
1C
#387800000000
0!
0*
09
0>
0C
#387810000000
1!
1*
19
1>
1C
#387820000000
0!
0*
09
0>
0C
#387830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#387840000000
0!
0*
09
0>
0C
#387850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#387860000000
0!
0*
09
0>
0C
#387870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#387880000000
0!
0*
09
0>
0C
#387890000000
1!
1*
b10 6
19
1>
1C
b10 G
#387900000000
0!
0*
09
0>
0C
#387910000000
1!
1*
b11 6
19
1>
1C
b11 G
#387920000000
0!
0*
09
0>
0C
#387930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#387940000000
0!
0*
09
0>
0C
#387950000000
1!
1*
b101 6
19
1>
1C
b101 G
#387960000000
0!
0*
09
0>
0C
#387970000000
1!
1*
b110 6
19
1>
1C
b110 G
#387980000000
0!
0*
09
0>
0C
#387990000000
1!
1*
b111 6
19
1>
1C
b111 G
#388000000000
0!
0*
09
0>
0C
#388010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#388020000000
0!
0*
09
0>
0C
#388030000000
1!
1*
b1 6
19
1>
1C
b1 G
#388040000000
0!
0*
09
0>
0C
#388050000000
1!
1*
b10 6
19
1>
1C
b10 G
#388060000000
0!
0*
09
0>
0C
#388070000000
1!
1*
b11 6
19
1>
1C
b11 G
#388080000000
0!
0*
09
0>
0C
#388090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#388100000000
0!
0*
09
0>
0C
#388110000000
1!
1*
b101 6
19
1>
1C
b101 G
#388120000000
0!
0*
09
0>
0C
#388130000000
1!
1*
b110 6
19
1>
1C
b110 G
#388140000000
0!
0*
09
0>
0C
#388150000000
1!
1*
b111 6
19
1>
1C
b111 G
#388160000000
0!
0*
09
0>
0C
#388170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#388180000000
0!
0*
09
0>
0C
#388190000000
1!
1*
b1 6
19
1>
1C
b1 G
#388200000000
0!
0*
09
0>
0C
#388210000000
1!
1*
b10 6
19
1>
1C
b10 G
#388220000000
0!
0*
09
0>
0C
#388230000000
1!
1*
b11 6
19
1>
1C
b11 G
#388240000000
0!
0*
09
0>
0C
#388250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#388260000000
0!
0*
09
0>
0C
#388270000000
1!
1*
b101 6
19
1>
1C
b101 G
#388280000000
0!
0*
09
0>
0C
#388290000000
1!
1*
b110 6
19
1>
1C
b110 G
#388300000000
0!
0*
09
0>
0C
#388310000000
1!
1*
b111 6
19
1>
1C
b111 G
#388320000000
0!
1"
0*
1+
09
1:
0>
0C
#388330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#388340000000
0!
0*
09
0>
0C
#388350000000
1!
1*
b1 6
19
1>
1C
b1 G
#388360000000
0!
0*
09
0>
0C
#388370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#388380000000
0!
0*
09
0>
0C
#388390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#388400000000
0!
0*
09
0>
0C
#388410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#388420000000
0!
0*
09
0>
0C
#388430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#388440000000
0!
0#
0*
0,
09
0>
0?
0C
#388450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#388460000000
0!
0*
09
0>
0C
#388470000000
1!
1*
19
1>
1C
#388480000000
0!
0*
09
0>
0C
#388490000000
1!
1*
19
1>
1C
#388500000000
0!
0*
09
0>
0C
#388510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#388520000000
0!
0*
09
0>
0C
#388530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#388540000000
0!
0*
09
0>
0C
#388550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#388560000000
0!
0*
09
0>
0C
#388570000000
1!
1*
b10 6
19
1>
1C
b10 G
#388580000000
0!
0*
09
0>
0C
#388590000000
1!
1*
b11 6
19
1>
1C
b11 G
#388600000000
0!
0*
09
0>
0C
#388610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#388620000000
0!
0*
09
0>
0C
#388630000000
1!
1*
b101 6
19
1>
1C
b101 G
#388640000000
0!
0*
09
0>
0C
#388650000000
1!
1*
b110 6
19
1>
1C
b110 G
#388660000000
0!
0*
09
0>
0C
#388670000000
1!
1*
b111 6
19
1>
1C
b111 G
#388680000000
0!
0*
09
0>
0C
#388690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#388700000000
0!
0*
09
0>
0C
#388710000000
1!
1*
b1 6
19
1>
1C
b1 G
#388720000000
0!
0*
09
0>
0C
#388730000000
1!
1*
b10 6
19
1>
1C
b10 G
#388740000000
0!
0*
09
0>
0C
#388750000000
1!
1*
b11 6
19
1>
1C
b11 G
#388760000000
0!
0*
09
0>
0C
#388770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#388780000000
0!
0*
09
0>
0C
#388790000000
1!
1*
b101 6
19
1>
1C
b101 G
#388800000000
0!
0*
09
0>
0C
#388810000000
1!
1*
b110 6
19
1>
1C
b110 G
#388820000000
0!
0*
09
0>
0C
#388830000000
1!
1*
b111 6
19
1>
1C
b111 G
#388840000000
0!
0*
09
0>
0C
#388850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#388860000000
0!
0*
09
0>
0C
#388870000000
1!
1*
b1 6
19
1>
1C
b1 G
#388880000000
0!
0*
09
0>
0C
#388890000000
1!
1*
b10 6
19
1>
1C
b10 G
#388900000000
0!
0*
09
0>
0C
#388910000000
1!
1*
b11 6
19
1>
1C
b11 G
#388920000000
0!
0*
09
0>
0C
#388930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#388940000000
0!
0*
09
0>
0C
#388950000000
1!
1*
b101 6
19
1>
1C
b101 G
#388960000000
0!
0*
09
0>
0C
#388970000000
1!
1*
b110 6
19
1>
1C
b110 G
#388980000000
0!
0*
09
0>
0C
#388990000000
1!
1*
b111 6
19
1>
1C
b111 G
#389000000000
0!
1"
0*
1+
09
1:
0>
0C
#389010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#389020000000
0!
0*
09
0>
0C
#389030000000
1!
1*
b1 6
19
1>
1C
b1 G
#389040000000
0!
0*
09
0>
0C
#389050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#389060000000
0!
0*
09
0>
0C
#389070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#389080000000
0!
0*
09
0>
0C
#389090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#389100000000
0!
0*
09
0>
0C
#389110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#389120000000
0!
0#
0*
0,
09
0>
0?
0C
#389130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#389140000000
0!
0*
09
0>
0C
#389150000000
1!
1*
19
1>
1C
#389160000000
0!
0*
09
0>
0C
#389170000000
1!
1*
19
1>
1C
#389180000000
0!
0*
09
0>
0C
#389190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#389200000000
0!
0*
09
0>
0C
#389210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#389220000000
0!
0*
09
0>
0C
#389230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#389240000000
0!
0*
09
0>
0C
#389250000000
1!
1*
b10 6
19
1>
1C
b10 G
#389260000000
0!
0*
09
0>
0C
#389270000000
1!
1*
b11 6
19
1>
1C
b11 G
#389280000000
0!
0*
09
0>
0C
#389290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#389300000000
0!
0*
09
0>
0C
#389310000000
1!
1*
b101 6
19
1>
1C
b101 G
#389320000000
0!
0*
09
0>
0C
#389330000000
1!
1*
b110 6
19
1>
1C
b110 G
#389340000000
0!
0*
09
0>
0C
#389350000000
1!
1*
b111 6
19
1>
1C
b111 G
#389360000000
0!
0*
09
0>
0C
#389370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#389380000000
0!
0*
09
0>
0C
#389390000000
1!
1*
b1 6
19
1>
1C
b1 G
#389400000000
0!
0*
09
0>
0C
#389410000000
1!
1*
b10 6
19
1>
1C
b10 G
#389420000000
0!
0*
09
0>
0C
#389430000000
1!
1*
b11 6
19
1>
1C
b11 G
#389440000000
0!
0*
09
0>
0C
#389450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#389460000000
0!
0*
09
0>
0C
#389470000000
1!
1*
b101 6
19
1>
1C
b101 G
#389480000000
0!
0*
09
0>
0C
#389490000000
1!
1*
b110 6
19
1>
1C
b110 G
#389500000000
0!
0*
09
0>
0C
#389510000000
1!
1*
b111 6
19
1>
1C
b111 G
#389520000000
0!
0*
09
0>
0C
#389530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#389540000000
0!
0*
09
0>
0C
#389550000000
1!
1*
b1 6
19
1>
1C
b1 G
#389560000000
0!
0*
09
0>
0C
#389570000000
1!
1*
b10 6
19
1>
1C
b10 G
#389580000000
0!
0*
09
0>
0C
#389590000000
1!
1*
b11 6
19
1>
1C
b11 G
#389600000000
0!
0*
09
0>
0C
#389610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#389620000000
0!
0*
09
0>
0C
#389630000000
1!
1*
b101 6
19
1>
1C
b101 G
#389640000000
0!
0*
09
0>
0C
#389650000000
1!
1*
b110 6
19
1>
1C
b110 G
#389660000000
0!
0*
09
0>
0C
#389670000000
1!
1*
b111 6
19
1>
1C
b111 G
#389680000000
0!
1"
0*
1+
09
1:
0>
0C
#389690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#389700000000
0!
0*
09
0>
0C
#389710000000
1!
1*
b1 6
19
1>
1C
b1 G
#389720000000
0!
0*
09
0>
0C
#389730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#389740000000
0!
0*
09
0>
0C
#389750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#389760000000
0!
0*
09
0>
0C
#389770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#389780000000
0!
0*
09
0>
0C
#389790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#389800000000
0!
0#
0*
0,
09
0>
0?
0C
#389810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#389820000000
0!
0*
09
0>
0C
#389830000000
1!
1*
19
1>
1C
#389840000000
0!
0*
09
0>
0C
#389850000000
1!
1*
19
1>
1C
#389860000000
0!
0*
09
0>
0C
#389870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#389880000000
0!
0*
09
0>
0C
#389890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#389900000000
0!
0*
09
0>
0C
#389910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#389920000000
0!
0*
09
0>
0C
#389930000000
1!
1*
b10 6
19
1>
1C
b10 G
#389940000000
0!
0*
09
0>
0C
#389950000000
1!
1*
b11 6
19
1>
1C
b11 G
#389960000000
0!
0*
09
0>
0C
#389970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#389980000000
0!
0*
09
0>
0C
#389990000000
1!
1*
b101 6
19
1>
1C
b101 G
#390000000000
0!
0*
09
0>
0C
#390010000000
1!
1*
b110 6
19
1>
1C
b110 G
#390020000000
0!
0*
09
0>
0C
#390030000000
1!
1*
b111 6
19
1>
1C
b111 G
#390040000000
0!
0*
09
0>
0C
#390050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#390060000000
0!
0*
09
0>
0C
#390070000000
1!
1*
b1 6
19
1>
1C
b1 G
#390080000000
0!
0*
09
0>
0C
#390090000000
1!
1*
b10 6
19
1>
1C
b10 G
#390100000000
0!
0*
09
0>
0C
#390110000000
1!
1*
b11 6
19
1>
1C
b11 G
#390120000000
0!
0*
09
0>
0C
#390130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#390140000000
0!
0*
09
0>
0C
#390150000000
1!
1*
b101 6
19
1>
1C
b101 G
#390160000000
0!
0*
09
0>
0C
#390170000000
1!
1*
b110 6
19
1>
1C
b110 G
#390180000000
0!
0*
09
0>
0C
#390190000000
1!
1*
b111 6
19
1>
1C
b111 G
#390200000000
0!
0*
09
0>
0C
#390210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#390220000000
0!
0*
09
0>
0C
#390230000000
1!
1*
b1 6
19
1>
1C
b1 G
#390240000000
0!
0*
09
0>
0C
#390250000000
1!
1*
b10 6
19
1>
1C
b10 G
#390260000000
0!
0*
09
0>
0C
#390270000000
1!
1*
b11 6
19
1>
1C
b11 G
#390280000000
0!
0*
09
0>
0C
#390290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#390300000000
0!
0*
09
0>
0C
#390310000000
1!
1*
b101 6
19
1>
1C
b101 G
#390320000000
0!
0*
09
0>
0C
#390330000000
1!
1*
b110 6
19
1>
1C
b110 G
#390340000000
0!
0*
09
0>
0C
#390350000000
1!
1*
b111 6
19
1>
1C
b111 G
#390360000000
0!
1"
0*
1+
09
1:
0>
0C
#390370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#390380000000
0!
0*
09
0>
0C
#390390000000
1!
1*
b1 6
19
1>
1C
b1 G
#390400000000
0!
0*
09
0>
0C
#390410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#390420000000
0!
0*
09
0>
0C
#390430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#390440000000
0!
0*
09
0>
0C
#390450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#390460000000
0!
0*
09
0>
0C
#390470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#390480000000
0!
0#
0*
0,
09
0>
0?
0C
#390490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#390500000000
0!
0*
09
0>
0C
#390510000000
1!
1*
19
1>
1C
#390520000000
0!
0*
09
0>
0C
#390530000000
1!
1*
19
1>
1C
#390540000000
0!
0*
09
0>
0C
#390550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#390560000000
0!
0*
09
0>
0C
#390570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#390580000000
0!
0*
09
0>
0C
#390590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#390600000000
0!
0*
09
0>
0C
#390610000000
1!
1*
b10 6
19
1>
1C
b10 G
#390620000000
0!
0*
09
0>
0C
#390630000000
1!
1*
b11 6
19
1>
1C
b11 G
#390640000000
0!
0*
09
0>
0C
#390650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#390660000000
0!
0*
09
0>
0C
#390670000000
1!
1*
b101 6
19
1>
1C
b101 G
#390680000000
0!
0*
09
0>
0C
#390690000000
1!
1*
b110 6
19
1>
1C
b110 G
#390700000000
0!
0*
09
0>
0C
#390710000000
1!
1*
b111 6
19
1>
1C
b111 G
#390720000000
0!
0*
09
0>
0C
#390730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#390740000000
0!
0*
09
0>
0C
#390750000000
1!
1*
b1 6
19
1>
1C
b1 G
#390760000000
0!
0*
09
0>
0C
#390770000000
1!
1*
b10 6
19
1>
1C
b10 G
#390780000000
0!
0*
09
0>
0C
#390790000000
1!
1*
b11 6
19
1>
1C
b11 G
#390800000000
0!
0*
09
0>
0C
#390810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#390820000000
0!
0*
09
0>
0C
#390830000000
1!
1*
b101 6
19
1>
1C
b101 G
#390840000000
0!
0*
09
0>
0C
#390850000000
1!
1*
b110 6
19
1>
1C
b110 G
#390860000000
0!
0*
09
0>
0C
#390870000000
1!
1*
b111 6
19
1>
1C
b111 G
#390880000000
0!
0*
09
0>
0C
#390890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#390900000000
0!
0*
09
0>
0C
#390910000000
1!
1*
b1 6
19
1>
1C
b1 G
#390920000000
0!
0*
09
0>
0C
#390930000000
1!
1*
b10 6
19
1>
1C
b10 G
#390940000000
0!
0*
09
0>
0C
#390950000000
1!
1*
b11 6
19
1>
1C
b11 G
#390960000000
0!
0*
09
0>
0C
#390970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#390980000000
0!
0*
09
0>
0C
#390990000000
1!
1*
b101 6
19
1>
1C
b101 G
#391000000000
0!
0*
09
0>
0C
#391010000000
1!
1*
b110 6
19
1>
1C
b110 G
#391020000000
0!
0*
09
0>
0C
#391030000000
1!
1*
b111 6
19
1>
1C
b111 G
#391040000000
0!
1"
0*
1+
09
1:
0>
0C
#391050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#391060000000
0!
0*
09
0>
0C
#391070000000
1!
1*
b1 6
19
1>
1C
b1 G
#391080000000
0!
0*
09
0>
0C
#391090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#391100000000
0!
0*
09
0>
0C
#391110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#391120000000
0!
0*
09
0>
0C
#391130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#391140000000
0!
0*
09
0>
0C
#391150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#391160000000
0!
0#
0*
0,
09
0>
0?
0C
#391170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#391180000000
0!
0*
09
0>
0C
#391190000000
1!
1*
19
1>
1C
#391200000000
0!
0*
09
0>
0C
#391210000000
1!
1*
19
1>
1C
#391220000000
0!
0*
09
0>
0C
#391230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#391240000000
0!
0*
09
0>
0C
#391250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#391260000000
0!
0*
09
0>
0C
#391270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#391280000000
0!
0*
09
0>
0C
#391290000000
1!
1*
b10 6
19
1>
1C
b10 G
#391300000000
0!
0*
09
0>
0C
#391310000000
1!
1*
b11 6
19
1>
1C
b11 G
#391320000000
0!
0*
09
0>
0C
#391330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#391340000000
0!
0*
09
0>
0C
#391350000000
1!
1*
b101 6
19
1>
1C
b101 G
#391360000000
0!
0*
09
0>
0C
#391370000000
1!
1*
b110 6
19
1>
1C
b110 G
#391380000000
0!
0*
09
0>
0C
#391390000000
1!
1*
b111 6
19
1>
1C
b111 G
#391400000000
0!
0*
09
0>
0C
#391410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#391420000000
0!
0*
09
0>
0C
#391430000000
1!
1*
b1 6
19
1>
1C
b1 G
#391440000000
0!
0*
09
0>
0C
#391450000000
1!
1*
b10 6
19
1>
1C
b10 G
#391460000000
0!
0*
09
0>
0C
#391470000000
1!
1*
b11 6
19
1>
1C
b11 G
#391480000000
0!
0*
09
0>
0C
#391490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#391500000000
0!
0*
09
0>
0C
#391510000000
1!
1*
b101 6
19
1>
1C
b101 G
#391520000000
0!
0*
09
0>
0C
#391530000000
1!
1*
b110 6
19
1>
1C
b110 G
#391540000000
0!
0*
09
0>
0C
#391550000000
1!
1*
b111 6
19
1>
1C
b111 G
#391560000000
0!
0*
09
0>
0C
#391570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#391580000000
0!
0*
09
0>
0C
#391590000000
1!
1*
b1 6
19
1>
1C
b1 G
#391600000000
0!
0*
09
0>
0C
#391610000000
1!
1*
b10 6
19
1>
1C
b10 G
#391620000000
0!
0*
09
0>
0C
#391630000000
1!
1*
b11 6
19
1>
1C
b11 G
#391640000000
0!
0*
09
0>
0C
#391650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#391660000000
0!
0*
09
0>
0C
#391670000000
1!
1*
b101 6
19
1>
1C
b101 G
#391680000000
0!
0*
09
0>
0C
#391690000000
1!
1*
b110 6
19
1>
1C
b110 G
#391700000000
0!
0*
09
0>
0C
#391710000000
1!
1*
b111 6
19
1>
1C
b111 G
#391720000000
0!
1"
0*
1+
09
1:
0>
0C
#391730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#391740000000
0!
0*
09
0>
0C
#391750000000
1!
1*
b1 6
19
1>
1C
b1 G
#391760000000
0!
0*
09
0>
0C
#391770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#391780000000
0!
0*
09
0>
0C
#391790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#391800000000
0!
0*
09
0>
0C
#391810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#391820000000
0!
0*
09
0>
0C
#391830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#391840000000
0!
0#
0*
0,
09
0>
0?
0C
#391850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#391860000000
0!
0*
09
0>
0C
#391870000000
1!
1*
19
1>
1C
#391880000000
0!
0*
09
0>
0C
#391890000000
1!
1*
19
1>
1C
#391900000000
0!
0*
09
0>
0C
#391910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#391920000000
0!
0*
09
0>
0C
#391930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#391940000000
0!
0*
09
0>
0C
#391950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#391960000000
0!
0*
09
0>
0C
#391970000000
1!
1*
b10 6
19
1>
1C
b10 G
#391980000000
0!
0*
09
0>
0C
#391990000000
1!
1*
b11 6
19
1>
1C
b11 G
#392000000000
0!
0*
09
0>
0C
#392010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#392020000000
0!
0*
09
0>
0C
#392030000000
1!
1*
b101 6
19
1>
1C
b101 G
#392040000000
0!
0*
09
0>
0C
#392050000000
1!
1*
b110 6
19
1>
1C
b110 G
#392060000000
0!
0*
09
0>
0C
#392070000000
1!
1*
b111 6
19
1>
1C
b111 G
#392080000000
0!
0*
09
0>
0C
#392090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#392100000000
0!
0*
09
0>
0C
#392110000000
1!
1*
b1 6
19
1>
1C
b1 G
#392120000000
0!
0*
09
0>
0C
#392130000000
1!
1*
b10 6
19
1>
1C
b10 G
#392140000000
0!
0*
09
0>
0C
#392150000000
1!
1*
b11 6
19
1>
1C
b11 G
#392160000000
0!
0*
09
0>
0C
#392170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#392180000000
0!
0*
09
0>
0C
#392190000000
1!
1*
b101 6
19
1>
1C
b101 G
#392200000000
0!
0*
09
0>
0C
#392210000000
1!
1*
b110 6
19
1>
1C
b110 G
#392220000000
0!
0*
09
0>
0C
#392230000000
1!
1*
b111 6
19
1>
1C
b111 G
#392240000000
0!
0*
09
0>
0C
#392250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#392260000000
0!
0*
09
0>
0C
#392270000000
1!
1*
b1 6
19
1>
1C
b1 G
#392280000000
0!
0*
09
0>
0C
#392290000000
1!
1*
b10 6
19
1>
1C
b10 G
#392300000000
0!
0*
09
0>
0C
#392310000000
1!
1*
b11 6
19
1>
1C
b11 G
#392320000000
0!
0*
09
0>
0C
#392330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#392340000000
0!
0*
09
0>
0C
#392350000000
1!
1*
b101 6
19
1>
1C
b101 G
#392360000000
0!
0*
09
0>
0C
#392370000000
1!
1*
b110 6
19
1>
1C
b110 G
#392380000000
0!
0*
09
0>
0C
#392390000000
1!
1*
b111 6
19
1>
1C
b111 G
#392400000000
0!
1"
0*
1+
09
1:
0>
0C
#392410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#392420000000
0!
0*
09
0>
0C
#392430000000
1!
1*
b1 6
19
1>
1C
b1 G
#392440000000
0!
0*
09
0>
0C
#392450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#392460000000
0!
0*
09
0>
0C
#392470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#392480000000
0!
0*
09
0>
0C
#392490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#392500000000
0!
0*
09
0>
0C
#392510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#392520000000
0!
0#
0*
0,
09
0>
0?
0C
#392530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#392540000000
0!
0*
09
0>
0C
#392550000000
1!
1*
19
1>
1C
#392560000000
0!
0*
09
0>
0C
#392570000000
1!
1*
19
1>
1C
#392580000000
0!
0*
09
0>
0C
#392590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#392600000000
0!
0*
09
0>
0C
#392610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#392620000000
0!
0*
09
0>
0C
#392630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#392640000000
0!
0*
09
0>
0C
#392650000000
1!
1*
b10 6
19
1>
1C
b10 G
#392660000000
0!
0*
09
0>
0C
#392670000000
1!
1*
b11 6
19
1>
1C
b11 G
#392680000000
0!
0*
09
0>
0C
#392690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#392700000000
0!
0*
09
0>
0C
#392710000000
1!
1*
b101 6
19
1>
1C
b101 G
#392720000000
0!
0*
09
0>
0C
#392730000000
1!
1*
b110 6
19
1>
1C
b110 G
#392740000000
0!
0*
09
0>
0C
#392750000000
1!
1*
b111 6
19
1>
1C
b111 G
#392760000000
0!
0*
09
0>
0C
#392770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#392780000000
0!
0*
09
0>
0C
#392790000000
1!
1*
b1 6
19
1>
1C
b1 G
#392800000000
0!
0*
09
0>
0C
#392810000000
1!
1*
b10 6
19
1>
1C
b10 G
#392820000000
0!
0*
09
0>
0C
#392830000000
1!
1*
b11 6
19
1>
1C
b11 G
#392840000000
0!
0*
09
0>
0C
#392850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#392860000000
0!
0*
09
0>
0C
#392870000000
1!
1*
b101 6
19
1>
1C
b101 G
#392880000000
0!
0*
09
0>
0C
#392890000000
1!
1*
b110 6
19
1>
1C
b110 G
#392900000000
0!
0*
09
0>
0C
#392910000000
1!
1*
b111 6
19
1>
1C
b111 G
#392920000000
0!
0*
09
0>
0C
#392930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#392940000000
0!
0*
09
0>
0C
#392950000000
1!
1*
b1 6
19
1>
1C
b1 G
#392960000000
0!
0*
09
0>
0C
#392970000000
1!
1*
b10 6
19
1>
1C
b10 G
#392980000000
0!
0*
09
0>
0C
#392990000000
1!
1*
b11 6
19
1>
1C
b11 G
#393000000000
0!
0*
09
0>
0C
#393010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#393020000000
0!
0*
09
0>
0C
#393030000000
1!
1*
b101 6
19
1>
1C
b101 G
#393040000000
0!
0*
09
0>
0C
#393050000000
1!
1*
b110 6
19
1>
1C
b110 G
#393060000000
0!
0*
09
0>
0C
#393070000000
1!
1*
b111 6
19
1>
1C
b111 G
#393080000000
0!
1"
0*
1+
09
1:
0>
0C
#393090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#393100000000
0!
0*
09
0>
0C
#393110000000
1!
1*
b1 6
19
1>
1C
b1 G
#393120000000
0!
0*
09
0>
0C
#393130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#393140000000
0!
0*
09
0>
0C
#393150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#393160000000
0!
0*
09
0>
0C
#393170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#393180000000
0!
0*
09
0>
0C
#393190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#393200000000
0!
0#
0*
0,
09
0>
0?
0C
#393210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#393220000000
0!
0*
09
0>
0C
#393230000000
1!
1*
19
1>
1C
#393240000000
0!
0*
09
0>
0C
#393250000000
1!
1*
19
1>
1C
#393260000000
0!
0*
09
0>
0C
#393270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#393280000000
0!
0*
09
0>
0C
#393290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#393300000000
0!
0*
09
0>
0C
#393310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#393320000000
0!
0*
09
0>
0C
#393330000000
1!
1*
b10 6
19
1>
1C
b10 G
#393340000000
0!
0*
09
0>
0C
#393350000000
1!
1*
b11 6
19
1>
1C
b11 G
#393360000000
0!
0*
09
0>
0C
#393370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#393380000000
0!
0*
09
0>
0C
#393390000000
1!
1*
b101 6
19
1>
1C
b101 G
#393400000000
0!
0*
09
0>
0C
#393410000000
1!
1*
b110 6
19
1>
1C
b110 G
#393420000000
0!
0*
09
0>
0C
#393430000000
1!
1*
b111 6
19
1>
1C
b111 G
#393440000000
0!
0*
09
0>
0C
#393450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#393460000000
0!
0*
09
0>
0C
#393470000000
1!
1*
b1 6
19
1>
1C
b1 G
#393480000000
0!
0*
09
0>
0C
#393490000000
1!
1*
b10 6
19
1>
1C
b10 G
#393500000000
0!
0*
09
0>
0C
#393510000000
1!
1*
b11 6
19
1>
1C
b11 G
#393520000000
0!
0*
09
0>
0C
#393530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#393540000000
0!
0*
09
0>
0C
#393550000000
1!
1*
b101 6
19
1>
1C
b101 G
#393560000000
0!
0*
09
0>
0C
#393570000000
1!
1*
b110 6
19
1>
1C
b110 G
#393580000000
0!
0*
09
0>
0C
#393590000000
1!
1*
b111 6
19
1>
1C
b111 G
#393600000000
0!
0*
09
0>
0C
#393610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#393620000000
0!
0*
09
0>
0C
#393630000000
1!
1*
b1 6
19
1>
1C
b1 G
#393640000000
0!
0*
09
0>
0C
#393650000000
1!
1*
b10 6
19
1>
1C
b10 G
#393660000000
0!
0*
09
0>
0C
#393670000000
1!
1*
b11 6
19
1>
1C
b11 G
#393680000000
0!
0*
09
0>
0C
#393690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#393700000000
0!
0*
09
0>
0C
#393710000000
1!
1*
b101 6
19
1>
1C
b101 G
#393720000000
0!
0*
09
0>
0C
#393730000000
1!
1*
b110 6
19
1>
1C
b110 G
#393740000000
0!
0*
09
0>
0C
#393750000000
1!
1*
b111 6
19
1>
1C
b111 G
#393760000000
0!
1"
0*
1+
09
1:
0>
0C
#393770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#393780000000
0!
0*
09
0>
0C
#393790000000
1!
1*
b1 6
19
1>
1C
b1 G
#393800000000
0!
0*
09
0>
0C
#393810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#393820000000
0!
0*
09
0>
0C
#393830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#393840000000
0!
0*
09
0>
0C
#393850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#393860000000
0!
0*
09
0>
0C
#393870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#393880000000
0!
0#
0*
0,
09
0>
0?
0C
#393890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#393900000000
0!
0*
09
0>
0C
#393910000000
1!
1*
19
1>
1C
#393920000000
0!
0*
09
0>
0C
#393930000000
1!
1*
19
1>
1C
#393940000000
0!
0*
09
0>
0C
#393950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#393960000000
0!
0*
09
0>
0C
#393970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#393980000000
0!
0*
09
0>
0C
#393990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#394000000000
0!
0*
09
0>
0C
#394010000000
1!
1*
b10 6
19
1>
1C
b10 G
#394020000000
0!
0*
09
0>
0C
#394030000000
1!
1*
b11 6
19
1>
1C
b11 G
#394040000000
0!
0*
09
0>
0C
#394050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#394060000000
0!
0*
09
0>
0C
#394070000000
1!
1*
b101 6
19
1>
1C
b101 G
#394080000000
0!
0*
09
0>
0C
#394090000000
1!
1*
b110 6
19
1>
1C
b110 G
#394100000000
0!
0*
09
0>
0C
#394110000000
1!
1*
b111 6
19
1>
1C
b111 G
#394120000000
0!
0*
09
0>
0C
#394130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#394140000000
0!
0*
09
0>
0C
#394150000000
1!
1*
b1 6
19
1>
1C
b1 G
#394160000000
0!
0*
09
0>
0C
#394170000000
1!
1*
b10 6
19
1>
1C
b10 G
#394180000000
0!
0*
09
0>
0C
#394190000000
1!
1*
b11 6
19
1>
1C
b11 G
#394200000000
0!
0*
09
0>
0C
#394210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#394220000000
0!
0*
09
0>
0C
#394230000000
1!
1*
b101 6
19
1>
1C
b101 G
#394240000000
0!
0*
09
0>
0C
#394250000000
1!
1*
b110 6
19
1>
1C
b110 G
#394260000000
0!
0*
09
0>
0C
#394270000000
1!
1*
b111 6
19
1>
1C
b111 G
#394280000000
0!
0*
09
0>
0C
#394290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#394300000000
0!
0*
09
0>
0C
#394310000000
1!
1*
b1 6
19
1>
1C
b1 G
#394320000000
0!
0*
09
0>
0C
#394330000000
1!
1*
b10 6
19
1>
1C
b10 G
#394340000000
0!
0*
09
0>
0C
#394350000000
1!
1*
b11 6
19
1>
1C
b11 G
#394360000000
0!
0*
09
0>
0C
#394370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#394380000000
0!
0*
09
0>
0C
#394390000000
1!
1*
b101 6
19
1>
1C
b101 G
#394400000000
0!
0*
09
0>
0C
#394410000000
1!
1*
b110 6
19
1>
1C
b110 G
#394420000000
0!
0*
09
0>
0C
#394430000000
1!
1*
b111 6
19
1>
1C
b111 G
#394440000000
0!
1"
0*
1+
09
1:
0>
0C
#394450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#394460000000
0!
0*
09
0>
0C
#394470000000
1!
1*
b1 6
19
1>
1C
b1 G
#394480000000
0!
0*
09
0>
0C
#394490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#394500000000
0!
0*
09
0>
0C
#394510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#394520000000
0!
0*
09
0>
0C
#394530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#394540000000
0!
0*
09
0>
0C
#394550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#394560000000
0!
0#
0*
0,
09
0>
0?
0C
#394570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#394580000000
0!
0*
09
0>
0C
#394590000000
1!
1*
19
1>
1C
#394600000000
0!
0*
09
0>
0C
#394610000000
1!
1*
19
1>
1C
#394620000000
0!
0*
09
0>
0C
#394630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#394640000000
0!
0*
09
0>
0C
#394650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#394660000000
0!
0*
09
0>
0C
#394670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#394680000000
0!
0*
09
0>
0C
#394690000000
1!
1*
b10 6
19
1>
1C
b10 G
#394700000000
0!
0*
09
0>
0C
#394710000000
1!
1*
b11 6
19
1>
1C
b11 G
#394720000000
0!
0*
09
0>
0C
#394730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#394740000000
0!
0*
09
0>
0C
#394750000000
1!
1*
b101 6
19
1>
1C
b101 G
#394760000000
0!
0*
09
0>
0C
#394770000000
1!
1*
b110 6
19
1>
1C
b110 G
#394780000000
0!
0*
09
0>
0C
#394790000000
1!
1*
b111 6
19
1>
1C
b111 G
#394800000000
0!
0*
09
0>
0C
#394810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#394820000000
0!
0*
09
0>
0C
#394830000000
1!
1*
b1 6
19
1>
1C
b1 G
#394840000000
0!
0*
09
0>
0C
#394850000000
1!
1*
b10 6
19
1>
1C
b10 G
#394860000000
0!
0*
09
0>
0C
#394870000000
1!
1*
b11 6
19
1>
1C
b11 G
#394880000000
0!
0*
09
0>
0C
#394890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#394900000000
0!
0*
09
0>
0C
#394910000000
1!
1*
b101 6
19
1>
1C
b101 G
#394920000000
0!
0*
09
0>
0C
#394930000000
1!
1*
b110 6
19
1>
1C
b110 G
#394940000000
0!
0*
09
0>
0C
#394950000000
1!
1*
b111 6
19
1>
1C
b111 G
#394960000000
0!
0*
09
0>
0C
#394970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#394980000000
0!
0*
09
0>
0C
#394990000000
1!
1*
b1 6
19
1>
1C
b1 G
#395000000000
0!
0*
09
0>
0C
#395010000000
1!
1*
b10 6
19
1>
1C
b10 G
#395020000000
0!
0*
09
0>
0C
#395030000000
1!
1*
b11 6
19
1>
1C
b11 G
#395040000000
0!
0*
09
0>
0C
#395050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#395060000000
0!
0*
09
0>
0C
#395070000000
1!
1*
b101 6
19
1>
1C
b101 G
#395080000000
0!
0*
09
0>
0C
#395090000000
1!
1*
b110 6
19
1>
1C
b110 G
#395100000000
0!
0*
09
0>
0C
#395110000000
1!
1*
b111 6
19
1>
1C
b111 G
#395120000000
0!
1"
0*
1+
09
1:
0>
0C
#395130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#395140000000
0!
0*
09
0>
0C
#395150000000
1!
1*
b1 6
19
1>
1C
b1 G
#395160000000
0!
0*
09
0>
0C
#395170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#395180000000
0!
0*
09
0>
0C
#395190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#395200000000
0!
0*
09
0>
0C
#395210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#395220000000
0!
0*
09
0>
0C
#395230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#395240000000
0!
0#
0*
0,
09
0>
0?
0C
#395250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#395260000000
0!
0*
09
0>
0C
#395270000000
1!
1*
19
1>
1C
#395280000000
0!
0*
09
0>
0C
#395290000000
1!
1*
19
1>
1C
#395300000000
0!
0*
09
0>
0C
#395310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#395320000000
0!
0*
09
0>
0C
#395330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#395340000000
0!
0*
09
0>
0C
#395350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#395360000000
0!
0*
09
0>
0C
#395370000000
1!
1*
b10 6
19
1>
1C
b10 G
#395380000000
0!
0*
09
0>
0C
#395390000000
1!
1*
b11 6
19
1>
1C
b11 G
#395400000000
0!
0*
09
0>
0C
#395410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#395420000000
0!
0*
09
0>
0C
#395430000000
1!
1*
b101 6
19
1>
1C
b101 G
#395440000000
0!
0*
09
0>
0C
#395450000000
1!
1*
b110 6
19
1>
1C
b110 G
#395460000000
0!
0*
09
0>
0C
#395470000000
1!
1*
b111 6
19
1>
1C
b111 G
#395480000000
0!
0*
09
0>
0C
#395490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#395500000000
0!
0*
09
0>
0C
#395510000000
1!
1*
b1 6
19
1>
1C
b1 G
#395520000000
0!
0*
09
0>
0C
#395530000000
1!
1*
b10 6
19
1>
1C
b10 G
#395540000000
0!
0*
09
0>
0C
#395550000000
1!
1*
b11 6
19
1>
1C
b11 G
#395560000000
0!
0*
09
0>
0C
#395570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#395580000000
0!
0*
09
0>
0C
#395590000000
1!
1*
b101 6
19
1>
1C
b101 G
#395600000000
0!
0*
09
0>
0C
#395610000000
1!
1*
b110 6
19
1>
1C
b110 G
#395620000000
0!
0*
09
0>
0C
#395630000000
1!
1*
b111 6
19
1>
1C
b111 G
#395640000000
0!
0*
09
0>
0C
#395650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#395660000000
0!
0*
09
0>
0C
#395670000000
1!
1*
b1 6
19
1>
1C
b1 G
#395680000000
0!
0*
09
0>
0C
#395690000000
1!
1*
b10 6
19
1>
1C
b10 G
#395700000000
0!
0*
09
0>
0C
#395710000000
1!
1*
b11 6
19
1>
1C
b11 G
#395720000000
0!
0*
09
0>
0C
#395730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#395740000000
0!
0*
09
0>
0C
#395750000000
1!
1*
b101 6
19
1>
1C
b101 G
#395760000000
0!
0*
09
0>
0C
#395770000000
1!
1*
b110 6
19
1>
1C
b110 G
#395780000000
0!
0*
09
0>
0C
#395790000000
1!
1*
b111 6
19
1>
1C
b111 G
#395800000000
0!
1"
0*
1+
09
1:
0>
0C
#395810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#395820000000
0!
0*
09
0>
0C
#395830000000
1!
1*
b1 6
19
1>
1C
b1 G
#395840000000
0!
0*
09
0>
0C
#395850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#395860000000
0!
0*
09
0>
0C
#395870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#395880000000
0!
0*
09
0>
0C
#395890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#395900000000
0!
0*
09
0>
0C
#395910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#395920000000
0!
0#
0*
0,
09
0>
0?
0C
#395930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#395940000000
0!
0*
09
0>
0C
#395950000000
1!
1*
19
1>
1C
#395960000000
0!
0*
09
0>
0C
#395970000000
1!
1*
19
1>
1C
#395980000000
0!
0*
09
0>
0C
#395990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#396000000000
0!
0*
09
0>
0C
#396010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#396020000000
0!
0*
09
0>
0C
#396030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#396040000000
0!
0*
09
0>
0C
#396050000000
1!
1*
b10 6
19
1>
1C
b10 G
#396060000000
0!
0*
09
0>
0C
#396070000000
1!
1*
b11 6
19
1>
1C
b11 G
#396080000000
0!
0*
09
0>
0C
#396090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#396100000000
0!
0*
09
0>
0C
#396110000000
1!
1*
b101 6
19
1>
1C
b101 G
#396120000000
0!
0*
09
0>
0C
#396130000000
1!
1*
b110 6
19
1>
1C
b110 G
#396140000000
0!
0*
09
0>
0C
#396150000000
1!
1*
b111 6
19
1>
1C
b111 G
#396160000000
0!
0*
09
0>
0C
#396170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#396180000000
0!
0*
09
0>
0C
#396190000000
1!
1*
b1 6
19
1>
1C
b1 G
#396200000000
0!
0*
09
0>
0C
#396210000000
1!
1*
b10 6
19
1>
1C
b10 G
#396220000000
0!
0*
09
0>
0C
#396230000000
1!
1*
b11 6
19
1>
1C
b11 G
#396240000000
0!
0*
09
0>
0C
#396250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#396260000000
0!
0*
09
0>
0C
#396270000000
1!
1*
b101 6
19
1>
1C
b101 G
#396280000000
0!
0*
09
0>
0C
#396290000000
1!
1*
b110 6
19
1>
1C
b110 G
#396300000000
0!
0*
09
0>
0C
#396310000000
1!
1*
b111 6
19
1>
1C
b111 G
#396320000000
0!
0*
09
0>
0C
#396330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#396340000000
0!
0*
09
0>
0C
#396350000000
1!
1*
b1 6
19
1>
1C
b1 G
#396360000000
0!
0*
09
0>
0C
#396370000000
1!
1*
b10 6
19
1>
1C
b10 G
#396380000000
0!
0*
09
0>
0C
#396390000000
1!
1*
b11 6
19
1>
1C
b11 G
#396400000000
0!
0*
09
0>
0C
#396410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#396420000000
0!
0*
09
0>
0C
#396430000000
1!
1*
b101 6
19
1>
1C
b101 G
#396440000000
0!
0*
09
0>
0C
#396450000000
1!
1*
b110 6
19
1>
1C
b110 G
#396460000000
0!
0*
09
0>
0C
#396470000000
1!
1*
b111 6
19
1>
1C
b111 G
#396480000000
0!
1"
0*
1+
09
1:
0>
0C
#396490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#396500000000
0!
0*
09
0>
0C
#396510000000
1!
1*
b1 6
19
1>
1C
b1 G
#396520000000
0!
0*
09
0>
0C
#396530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#396540000000
0!
0*
09
0>
0C
#396550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#396560000000
0!
0*
09
0>
0C
#396570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#396580000000
0!
0*
09
0>
0C
#396590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#396600000000
0!
0#
0*
0,
09
0>
0?
0C
#396610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#396620000000
0!
0*
09
0>
0C
#396630000000
1!
1*
19
1>
1C
#396640000000
0!
0*
09
0>
0C
#396650000000
1!
1*
19
1>
1C
#396660000000
0!
0*
09
0>
0C
#396670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#396680000000
0!
0*
09
0>
0C
#396690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#396700000000
0!
0*
09
0>
0C
#396710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#396720000000
0!
0*
09
0>
0C
#396730000000
1!
1*
b10 6
19
1>
1C
b10 G
#396740000000
0!
0*
09
0>
0C
#396750000000
1!
1*
b11 6
19
1>
1C
b11 G
#396760000000
0!
0*
09
0>
0C
#396770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#396780000000
0!
0*
09
0>
0C
#396790000000
1!
1*
b101 6
19
1>
1C
b101 G
#396800000000
0!
0*
09
0>
0C
#396810000000
1!
1*
b110 6
19
1>
1C
b110 G
#396820000000
0!
0*
09
0>
0C
#396830000000
1!
1*
b111 6
19
1>
1C
b111 G
#396840000000
0!
0*
09
0>
0C
#396850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#396860000000
0!
0*
09
0>
0C
#396870000000
1!
1*
b1 6
19
1>
1C
b1 G
#396880000000
0!
0*
09
0>
0C
#396890000000
1!
1*
b10 6
19
1>
1C
b10 G
#396900000000
0!
0*
09
0>
0C
#396910000000
1!
1*
b11 6
19
1>
1C
b11 G
#396920000000
0!
0*
09
0>
0C
#396930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#396940000000
0!
0*
09
0>
0C
#396950000000
1!
1*
b101 6
19
1>
1C
b101 G
#396960000000
0!
0*
09
0>
0C
#396970000000
1!
1*
b110 6
19
1>
1C
b110 G
#396980000000
0!
0*
09
0>
0C
#396990000000
1!
1*
b111 6
19
1>
1C
b111 G
#397000000000
0!
0*
09
0>
0C
#397010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#397020000000
0!
0*
09
0>
0C
#397030000000
1!
1*
b1 6
19
1>
1C
b1 G
#397040000000
0!
0*
09
0>
0C
#397050000000
1!
1*
b10 6
19
1>
1C
b10 G
#397060000000
0!
0*
09
0>
0C
#397070000000
1!
1*
b11 6
19
1>
1C
b11 G
#397080000000
0!
0*
09
0>
0C
#397090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#397100000000
0!
0*
09
0>
0C
#397110000000
1!
1*
b101 6
19
1>
1C
b101 G
#397120000000
0!
0*
09
0>
0C
#397130000000
1!
1*
b110 6
19
1>
1C
b110 G
#397140000000
0!
0*
09
0>
0C
#397150000000
1!
1*
b111 6
19
1>
1C
b111 G
#397160000000
0!
1"
0*
1+
09
1:
0>
0C
#397170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#397180000000
0!
0*
09
0>
0C
#397190000000
1!
1*
b1 6
19
1>
1C
b1 G
#397200000000
0!
0*
09
0>
0C
#397210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#397220000000
0!
0*
09
0>
0C
#397230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#397240000000
0!
0*
09
0>
0C
#397250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#397260000000
0!
0*
09
0>
0C
#397270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#397280000000
0!
0#
0*
0,
09
0>
0?
0C
#397290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#397300000000
0!
0*
09
0>
0C
#397310000000
1!
1*
19
1>
1C
#397320000000
0!
0*
09
0>
0C
#397330000000
1!
1*
19
1>
1C
#397340000000
0!
0*
09
0>
0C
#397350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#397360000000
0!
0*
09
0>
0C
#397370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#397380000000
0!
0*
09
0>
0C
#397390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#397400000000
0!
0*
09
0>
0C
#397410000000
1!
1*
b10 6
19
1>
1C
b10 G
#397420000000
0!
0*
09
0>
0C
#397430000000
1!
1*
b11 6
19
1>
1C
b11 G
#397440000000
0!
0*
09
0>
0C
#397450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#397460000000
0!
0*
09
0>
0C
#397470000000
1!
1*
b101 6
19
1>
1C
b101 G
#397480000000
0!
0*
09
0>
0C
#397490000000
1!
1*
b110 6
19
1>
1C
b110 G
#397500000000
0!
0*
09
0>
0C
#397510000000
1!
1*
b111 6
19
1>
1C
b111 G
#397520000000
0!
0*
09
0>
0C
#397530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#397540000000
0!
0*
09
0>
0C
#397550000000
1!
1*
b1 6
19
1>
1C
b1 G
#397560000000
0!
0*
09
0>
0C
#397570000000
1!
1*
b10 6
19
1>
1C
b10 G
#397580000000
0!
0*
09
0>
0C
#397590000000
1!
1*
b11 6
19
1>
1C
b11 G
#397600000000
0!
0*
09
0>
0C
#397610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#397620000000
0!
0*
09
0>
0C
#397630000000
1!
1*
b101 6
19
1>
1C
b101 G
#397640000000
0!
0*
09
0>
0C
#397650000000
1!
1*
b110 6
19
1>
1C
b110 G
#397660000000
0!
0*
09
0>
0C
#397670000000
1!
1*
b111 6
19
1>
1C
b111 G
#397680000000
0!
0*
09
0>
0C
#397690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#397700000000
0!
0*
09
0>
0C
#397710000000
1!
1*
b1 6
19
1>
1C
b1 G
#397720000000
0!
0*
09
0>
0C
#397730000000
1!
1*
b10 6
19
1>
1C
b10 G
#397740000000
0!
0*
09
0>
0C
#397750000000
1!
1*
b11 6
19
1>
1C
b11 G
#397760000000
0!
0*
09
0>
0C
#397770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#397780000000
0!
0*
09
0>
0C
#397790000000
1!
1*
b101 6
19
1>
1C
b101 G
#397800000000
0!
0*
09
0>
0C
#397810000000
1!
1*
b110 6
19
1>
1C
b110 G
#397820000000
0!
0*
09
0>
0C
#397830000000
1!
1*
b111 6
19
1>
1C
b111 G
#397840000000
0!
1"
0*
1+
09
1:
0>
0C
#397850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#397860000000
0!
0*
09
0>
0C
#397870000000
1!
1*
b1 6
19
1>
1C
b1 G
#397880000000
0!
0*
09
0>
0C
#397890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#397900000000
0!
0*
09
0>
0C
#397910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#397920000000
0!
0*
09
0>
0C
#397930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#397940000000
0!
0*
09
0>
0C
#397950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#397960000000
0!
0#
0*
0,
09
0>
0?
0C
#397970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#397980000000
0!
0*
09
0>
0C
#397990000000
1!
1*
19
1>
1C
#398000000000
0!
0*
09
0>
0C
#398010000000
1!
1*
19
1>
1C
#398020000000
0!
0*
09
0>
0C
#398030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#398040000000
0!
0*
09
0>
0C
#398050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#398060000000
0!
0*
09
0>
0C
#398070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#398080000000
0!
0*
09
0>
0C
#398090000000
1!
1*
b10 6
19
1>
1C
b10 G
#398100000000
0!
0*
09
0>
0C
#398110000000
1!
1*
b11 6
19
1>
1C
b11 G
#398120000000
0!
0*
09
0>
0C
#398130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#398140000000
0!
0*
09
0>
0C
#398150000000
1!
1*
b101 6
19
1>
1C
b101 G
#398160000000
0!
0*
09
0>
0C
#398170000000
1!
1*
b110 6
19
1>
1C
b110 G
#398180000000
0!
0*
09
0>
0C
#398190000000
1!
1*
b111 6
19
1>
1C
b111 G
#398200000000
0!
0*
09
0>
0C
#398210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#398220000000
0!
0*
09
0>
0C
#398230000000
1!
1*
b1 6
19
1>
1C
b1 G
#398240000000
0!
0*
09
0>
0C
#398250000000
1!
1*
b10 6
19
1>
1C
b10 G
#398260000000
0!
0*
09
0>
0C
#398270000000
1!
1*
b11 6
19
1>
1C
b11 G
#398280000000
0!
0*
09
0>
0C
#398290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#398300000000
0!
0*
09
0>
0C
#398310000000
1!
1*
b101 6
19
1>
1C
b101 G
#398320000000
0!
0*
09
0>
0C
#398330000000
1!
1*
b110 6
19
1>
1C
b110 G
#398340000000
0!
0*
09
0>
0C
#398350000000
1!
1*
b111 6
19
1>
1C
b111 G
#398360000000
0!
0*
09
0>
0C
#398370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#398380000000
0!
0*
09
0>
0C
#398390000000
1!
1*
b1 6
19
1>
1C
b1 G
#398400000000
0!
0*
09
0>
0C
#398410000000
1!
1*
b10 6
19
1>
1C
b10 G
#398420000000
0!
0*
09
0>
0C
#398430000000
1!
1*
b11 6
19
1>
1C
b11 G
#398440000000
0!
0*
09
0>
0C
#398450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#398460000000
0!
0*
09
0>
0C
#398470000000
1!
1*
b101 6
19
1>
1C
b101 G
#398480000000
0!
0*
09
0>
0C
#398490000000
1!
1*
b110 6
19
1>
1C
b110 G
#398500000000
0!
0*
09
0>
0C
#398510000000
1!
1*
b111 6
19
1>
1C
b111 G
#398520000000
0!
1"
0*
1+
09
1:
0>
0C
#398530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#398540000000
0!
0*
09
0>
0C
#398550000000
1!
1*
b1 6
19
1>
1C
b1 G
#398560000000
0!
0*
09
0>
0C
#398570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#398580000000
0!
0*
09
0>
0C
#398590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#398600000000
0!
0*
09
0>
0C
#398610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#398620000000
0!
0*
09
0>
0C
#398630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#398640000000
0!
0#
0*
0,
09
0>
0?
0C
#398650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#398660000000
0!
0*
09
0>
0C
#398670000000
1!
1*
19
1>
1C
#398680000000
0!
0*
09
0>
0C
#398690000000
1!
1*
19
1>
1C
#398700000000
0!
0*
09
0>
0C
#398710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#398720000000
0!
0*
09
0>
0C
#398730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#398740000000
0!
0*
09
0>
0C
#398750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#398760000000
0!
0*
09
0>
0C
#398770000000
1!
1*
b10 6
19
1>
1C
b10 G
#398780000000
0!
0*
09
0>
0C
#398790000000
1!
1*
b11 6
19
1>
1C
b11 G
#398800000000
0!
0*
09
0>
0C
#398810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#398820000000
0!
0*
09
0>
0C
#398830000000
1!
1*
b101 6
19
1>
1C
b101 G
#398840000000
0!
0*
09
0>
0C
#398850000000
1!
1*
b110 6
19
1>
1C
b110 G
#398860000000
0!
0*
09
0>
0C
#398870000000
1!
1*
b111 6
19
1>
1C
b111 G
#398880000000
0!
0*
09
0>
0C
#398890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#398900000000
0!
0*
09
0>
0C
#398910000000
1!
1*
b1 6
19
1>
1C
b1 G
#398920000000
0!
0*
09
0>
0C
#398930000000
1!
1*
b10 6
19
1>
1C
b10 G
#398940000000
0!
0*
09
0>
0C
#398950000000
1!
1*
b11 6
19
1>
1C
b11 G
#398960000000
0!
0*
09
0>
0C
#398970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#398980000000
0!
0*
09
0>
0C
#398990000000
1!
1*
b101 6
19
1>
1C
b101 G
#399000000000
0!
0*
09
0>
0C
#399010000000
1!
1*
b110 6
19
1>
1C
b110 G
#399020000000
0!
0*
09
0>
0C
#399030000000
1!
1*
b111 6
19
1>
1C
b111 G
#399040000000
0!
0*
09
0>
0C
#399050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#399060000000
0!
0*
09
0>
0C
#399070000000
1!
1*
b1 6
19
1>
1C
b1 G
#399080000000
0!
0*
09
0>
0C
#399090000000
1!
1*
b10 6
19
1>
1C
b10 G
#399100000000
0!
0*
09
0>
0C
#399110000000
1!
1*
b11 6
19
1>
1C
b11 G
#399120000000
0!
0*
09
0>
0C
#399130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#399140000000
0!
0*
09
0>
0C
#399150000000
1!
1*
b101 6
19
1>
1C
b101 G
#399160000000
0!
0*
09
0>
0C
#399170000000
1!
1*
b110 6
19
1>
1C
b110 G
#399180000000
0!
0*
09
0>
0C
#399190000000
1!
1*
b111 6
19
1>
1C
b111 G
#399200000000
0!
1"
0*
1+
09
1:
0>
0C
#399210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#399220000000
0!
0*
09
0>
0C
#399230000000
1!
1*
b1 6
19
1>
1C
b1 G
#399240000000
0!
0*
09
0>
0C
#399250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#399260000000
0!
0*
09
0>
0C
#399270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#399280000000
0!
0*
09
0>
0C
#399290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#399300000000
0!
0*
09
0>
0C
#399310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#399320000000
0!
0#
0*
0,
09
0>
0?
0C
#399330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#399340000000
0!
0*
09
0>
0C
#399350000000
1!
1*
19
1>
1C
#399360000000
0!
0*
09
0>
0C
#399370000000
1!
1*
19
1>
1C
#399380000000
0!
0*
09
0>
0C
#399390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#399400000000
0!
0*
09
0>
0C
#399410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#399420000000
0!
0*
09
0>
0C
#399430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#399440000000
0!
0*
09
0>
0C
#399450000000
1!
1*
b10 6
19
1>
1C
b10 G
#399460000000
0!
0*
09
0>
0C
#399470000000
1!
1*
b11 6
19
1>
1C
b11 G
#399480000000
0!
0*
09
0>
0C
#399490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#399500000000
0!
0*
09
0>
0C
#399510000000
1!
1*
b101 6
19
1>
1C
b101 G
#399520000000
0!
0*
09
0>
0C
#399530000000
1!
1*
b110 6
19
1>
1C
b110 G
#399540000000
0!
0*
09
0>
0C
#399550000000
1!
1*
b111 6
19
1>
1C
b111 G
#399560000000
0!
0*
09
0>
0C
#399570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#399580000000
0!
0*
09
0>
0C
#399590000000
1!
1*
b1 6
19
1>
1C
b1 G
#399600000000
0!
0*
09
0>
0C
#399610000000
1!
1*
b10 6
19
1>
1C
b10 G
#399620000000
0!
0*
09
0>
0C
#399630000000
1!
1*
b11 6
19
1>
1C
b11 G
#399640000000
0!
0*
09
0>
0C
#399650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#399660000000
0!
0*
09
0>
0C
#399670000000
1!
1*
b101 6
19
1>
1C
b101 G
#399680000000
0!
0*
09
0>
0C
#399690000000
1!
1*
b110 6
19
1>
1C
b110 G
#399700000000
0!
0*
09
0>
0C
#399710000000
1!
1*
b111 6
19
1>
1C
b111 G
#399720000000
0!
0*
09
0>
0C
#399730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#399740000000
0!
0*
09
0>
0C
#399750000000
1!
1*
b1 6
19
1>
1C
b1 G
#399760000000
0!
0*
09
0>
0C
#399770000000
1!
1*
b10 6
19
1>
1C
b10 G
#399780000000
0!
0*
09
0>
0C
#399790000000
1!
1*
b11 6
19
1>
1C
b11 G
#399800000000
0!
0*
09
0>
0C
#399810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#399820000000
0!
0*
09
0>
0C
#399830000000
1!
1*
b101 6
19
1>
1C
b101 G
#399840000000
0!
0*
09
0>
0C
#399850000000
1!
1*
b110 6
19
1>
1C
b110 G
#399860000000
0!
0*
09
0>
0C
#399870000000
1!
1*
b111 6
19
1>
1C
b111 G
#399880000000
0!
1"
0*
1+
09
1:
0>
0C
#399890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#399900000000
0!
0*
09
0>
0C
#399910000000
1!
1*
b1 6
19
1>
1C
b1 G
#399920000000
0!
0*
09
0>
0C
#399930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#399940000000
0!
0*
09
0>
0C
#399950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#399960000000
0!
0*
09
0>
0C
#399970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#399980000000
0!
0*
09
0>
0C
#399990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#400000000000
0!
0#
0*
0,
09
0>
0?
0C
#400010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#400020000000
0!
0*
09
0>
0C
#400030000000
1!
1*
19
1>
1C
#400040000000
0!
0*
09
0>
0C
#400050000000
1!
1*
19
1>
1C
#400060000000
0!
0*
09
0>
0C
#400070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#400080000000
0!
0*
09
0>
0C
#400090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#400100000000
0!
0*
09
0>
0C
#400110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#400120000000
0!
0*
09
0>
0C
#400130000000
1!
1*
b10 6
19
1>
1C
b10 G
#400140000000
0!
0*
09
0>
0C
#400150000000
1!
1*
b11 6
19
1>
1C
b11 G
#400160000000
0!
0*
09
0>
0C
#400170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#400180000000
0!
0*
09
0>
0C
#400190000000
1!
1*
b101 6
19
1>
1C
b101 G
#400200000000
0!
0*
09
0>
0C
#400210000000
1!
1*
b110 6
19
1>
1C
b110 G
#400220000000
0!
0*
09
0>
0C
#400230000000
1!
1*
b111 6
19
1>
1C
b111 G
#400240000000
0!
0*
09
0>
0C
#400250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#400260000000
0!
0*
09
0>
0C
#400270000000
1!
1*
b1 6
19
1>
1C
b1 G
#400280000000
0!
0*
09
0>
0C
#400290000000
1!
1*
b10 6
19
1>
1C
b10 G
#400300000000
0!
0*
09
0>
0C
#400310000000
1!
1*
b11 6
19
1>
1C
b11 G
#400320000000
0!
0*
09
0>
0C
#400330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#400340000000
0!
0*
09
0>
0C
#400350000000
1!
1*
b101 6
19
1>
1C
b101 G
#400360000000
0!
0*
09
0>
0C
#400370000000
1!
1*
b110 6
19
1>
1C
b110 G
#400380000000
0!
0*
09
0>
0C
#400390000000
1!
1*
b111 6
19
1>
1C
b111 G
#400400000000
0!
0*
09
0>
0C
#400410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#400420000000
0!
0*
09
0>
0C
#400430000000
1!
1*
b1 6
19
1>
1C
b1 G
#400440000000
0!
0*
09
0>
0C
#400450000000
1!
1*
b10 6
19
1>
1C
b10 G
#400460000000
0!
0*
09
0>
0C
#400470000000
1!
1*
b11 6
19
1>
1C
b11 G
#400480000000
0!
0*
09
0>
0C
#400490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#400500000000
0!
0*
09
0>
0C
#400510000000
1!
1*
b101 6
19
1>
1C
b101 G
#400520000000
0!
0*
09
0>
0C
#400530000000
1!
1*
b110 6
19
1>
1C
b110 G
#400540000000
0!
0*
09
0>
0C
#400550000000
1!
1*
b111 6
19
1>
1C
b111 G
#400560000000
0!
1"
0*
1+
09
1:
0>
0C
#400570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#400580000000
0!
0*
09
0>
0C
#400590000000
1!
1*
b1 6
19
1>
1C
b1 G
#400600000000
0!
0*
09
0>
0C
#400610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#400620000000
0!
0*
09
0>
0C
#400630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#400640000000
0!
0*
09
0>
0C
#400650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#400660000000
0!
0*
09
0>
0C
#400670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#400680000000
0!
0#
0*
0,
09
0>
0?
0C
#400690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#400700000000
0!
0*
09
0>
0C
#400710000000
1!
1*
19
1>
1C
#400720000000
0!
0*
09
0>
0C
#400730000000
1!
1*
19
1>
1C
#400740000000
0!
0*
09
0>
0C
#400750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#400760000000
0!
0*
09
0>
0C
#400770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#400780000000
0!
0*
09
0>
0C
#400790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#400800000000
0!
0*
09
0>
0C
#400810000000
1!
1*
b10 6
19
1>
1C
b10 G
#400820000000
0!
0*
09
0>
0C
#400830000000
1!
1*
b11 6
19
1>
1C
b11 G
#400840000000
0!
0*
09
0>
0C
#400850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#400860000000
0!
0*
09
0>
0C
#400870000000
1!
1*
b101 6
19
1>
1C
b101 G
#400880000000
0!
0*
09
0>
0C
#400890000000
1!
1*
b110 6
19
1>
1C
b110 G
#400900000000
0!
0*
09
0>
0C
#400910000000
1!
1*
b111 6
19
1>
1C
b111 G
#400920000000
0!
0*
09
0>
0C
#400930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#400940000000
0!
0*
09
0>
0C
#400950000000
1!
1*
b1 6
19
1>
1C
b1 G
#400960000000
0!
0*
09
0>
0C
#400970000000
1!
1*
b10 6
19
1>
1C
b10 G
#400980000000
0!
0*
09
0>
0C
#400990000000
1!
1*
b11 6
19
1>
1C
b11 G
#401000000000
0!
0*
09
0>
0C
#401010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#401020000000
0!
0*
09
0>
0C
#401030000000
1!
1*
b101 6
19
1>
1C
b101 G
#401040000000
0!
0*
09
0>
0C
#401050000000
1!
1*
b110 6
19
1>
1C
b110 G
#401060000000
0!
0*
09
0>
0C
#401070000000
1!
1*
b111 6
19
1>
1C
b111 G
#401080000000
0!
0*
09
0>
0C
#401090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#401100000000
0!
0*
09
0>
0C
#401110000000
1!
1*
b1 6
19
1>
1C
b1 G
#401120000000
0!
0*
09
0>
0C
#401130000000
1!
1*
b10 6
19
1>
1C
b10 G
#401140000000
0!
0*
09
0>
0C
#401150000000
1!
1*
b11 6
19
1>
1C
b11 G
#401160000000
0!
0*
09
0>
0C
#401170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#401180000000
0!
0*
09
0>
0C
#401190000000
1!
1*
b101 6
19
1>
1C
b101 G
#401200000000
0!
0*
09
0>
0C
#401210000000
1!
1*
b110 6
19
1>
1C
b110 G
#401220000000
0!
0*
09
0>
0C
#401230000000
1!
1*
b111 6
19
1>
1C
b111 G
#401240000000
0!
1"
0*
1+
09
1:
0>
0C
#401250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#401260000000
0!
0*
09
0>
0C
#401270000000
1!
1*
b1 6
19
1>
1C
b1 G
#401280000000
0!
0*
09
0>
0C
#401290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#401300000000
0!
0*
09
0>
0C
#401310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#401320000000
0!
0*
09
0>
0C
#401330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#401340000000
0!
0*
09
0>
0C
#401350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#401360000000
0!
0#
0*
0,
09
0>
0?
0C
#401370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#401380000000
0!
0*
09
0>
0C
#401390000000
1!
1*
19
1>
1C
#401400000000
0!
0*
09
0>
0C
#401410000000
1!
1*
19
1>
1C
#401420000000
0!
0*
09
0>
0C
#401430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#401440000000
0!
0*
09
0>
0C
#401450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#401460000000
0!
0*
09
0>
0C
#401470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#401480000000
0!
0*
09
0>
0C
#401490000000
1!
1*
b10 6
19
1>
1C
b10 G
#401500000000
0!
0*
09
0>
0C
#401510000000
1!
1*
b11 6
19
1>
1C
b11 G
#401520000000
0!
0*
09
0>
0C
#401530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#401540000000
0!
0*
09
0>
0C
#401550000000
1!
1*
b101 6
19
1>
1C
b101 G
#401560000000
0!
0*
09
0>
0C
#401570000000
1!
1*
b110 6
19
1>
1C
b110 G
#401580000000
0!
0*
09
0>
0C
#401590000000
1!
1*
b111 6
19
1>
1C
b111 G
#401600000000
0!
0*
09
0>
0C
#401610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#401620000000
0!
0*
09
0>
0C
#401630000000
1!
1*
b1 6
19
1>
1C
b1 G
#401640000000
0!
0*
09
0>
0C
#401650000000
1!
1*
b10 6
19
1>
1C
b10 G
#401660000000
0!
0*
09
0>
0C
#401670000000
1!
1*
b11 6
19
1>
1C
b11 G
#401680000000
0!
0*
09
0>
0C
#401690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#401700000000
0!
0*
09
0>
0C
#401710000000
1!
1*
b101 6
19
1>
1C
b101 G
#401720000000
0!
0*
09
0>
0C
#401730000000
1!
1*
b110 6
19
1>
1C
b110 G
#401740000000
0!
0*
09
0>
0C
#401750000000
1!
1*
b111 6
19
1>
1C
b111 G
#401760000000
0!
0*
09
0>
0C
#401770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#401780000000
0!
0*
09
0>
0C
#401790000000
1!
1*
b1 6
19
1>
1C
b1 G
#401800000000
0!
0*
09
0>
0C
#401810000000
1!
1*
b10 6
19
1>
1C
b10 G
#401820000000
0!
0*
09
0>
0C
#401830000000
1!
1*
b11 6
19
1>
1C
b11 G
#401840000000
0!
0*
09
0>
0C
#401850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#401860000000
0!
0*
09
0>
0C
#401870000000
1!
1*
b101 6
19
1>
1C
b101 G
#401880000000
0!
0*
09
0>
0C
#401890000000
1!
1*
b110 6
19
1>
1C
b110 G
#401900000000
0!
0*
09
0>
0C
#401910000000
1!
1*
b111 6
19
1>
1C
b111 G
#401920000000
0!
1"
0*
1+
09
1:
0>
0C
#401930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#401940000000
0!
0*
09
0>
0C
#401950000000
1!
1*
b1 6
19
1>
1C
b1 G
#401960000000
0!
0*
09
0>
0C
#401970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#401980000000
0!
0*
09
0>
0C
#401990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#402000000000
0!
0*
09
0>
0C
#402010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#402020000000
0!
0*
09
0>
0C
#402030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#402040000000
0!
0#
0*
0,
09
0>
0?
0C
#402050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#402060000000
0!
0*
09
0>
0C
#402070000000
1!
1*
19
1>
1C
#402080000000
0!
0*
09
0>
0C
#402090000000
1!
1*
19
1>
1C
#402100000000
0!
0*
09
0>
0C
#402110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#402120000000
0!
0*
09
0>
0C
#402130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#402140000000
0!
0*
09
0>
0C
#402150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#402160000000
0!
0*
09
0>
0C
#402170000000
1!
1*
b10 6
19
1>
1C
b10 G
#402180000000
0!
0*
09
0>
0C
#402190000000
1!
1*
b11 6
19
1>
1C
b11 G
#402200000000
0!
0*
09
0>
0C
#402210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#402220000000
0!
0*
09
0>
0C
#402230000000
1!
1*
b101 6
19
1>
1C
b101 G
#402240000000
0!
0*
09
0>
0C
#402250000000
1!
1*
b110 6
19
1>
1C
b110 G
#402260000000
0!
0*
09
0>
0C
#402270000000
1!
1*
b111 6
19
1>
1C
b111 G
#402280000000
0!
0*
09
0>
0C
#402290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#402300000000
0!
0*
09
0>
0C
#402310000000
1!
1*
b1 6
19
1>
1C
b1 G
#402320000000
0!
0*
09
0>
0C
#402330000000
1!
1*
b10 6
19
1>
1C
b10 G
#402340000000
0!
0*
09
0>
0C
#402350000000
1!
1*
b11 6
19
1>
1C
b11 G
#402360000000
0!
0*
09
0>
0C
#402370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#402380000000
0!
0*
09
0>
0C
#402390000000
1!
1*
b101 6
19
1>
1C
b101 G
#402400000000
0!
0*
09
0>
0C
#402410000000
1!
1*
b110 6
19
1>
1C
b110 G
#402420000000
0!
0*
09
0>
0C
#402430000000
1!
1*
b111 6
19
1>
1C
b111 G
#402440000000
0!
0*
09
0>
0C
#402450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#402460000000
0!
0*
09
0>
0C
#402470000000
1!
1*
b1 6
19
1>
1C
b1 G
#402480000000
0!
0*
09
0>
0C
#402490000000
1!
1*
b10 6
19
1>
1C
b10 G
#402500000000
0!
0*
09
0>
0C
#402510000000
1!
1*
b11 6
19
1>
1C
b11 G
#402520000000
0!
0*
09
0>
0C
#402530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#402540000000
0!
0*
09
0>
0C
#402550000000
1!
1*
b101 6
19
1>
1C
b101 G
#402560000000
0!
0*
09
0>
0C
#402570000000
1!
1*
b110 6
19
1>
1C
b110 G
#402580000000
0!
0*
09
0>
0C
#402590000000
1!
1*
b111 6
19
1>
1C
b111 G
#402600000000
0!
1"
0*
1+
09
1:
0>
0C
#402610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#402620000000
0!
0*
09
0>
0C
#402630000000
1!
1*
b1 6
19
1>
1C
b1 G
#402640000000
0!
0*
09
0>
0C
#402650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#402660000000
0!
0*
09
0>
0C
#402670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#402680000000
0!
0*
09
0>
0C
#402690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#402700000000
0!
0*
09
0>
0C
#402710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#402720000000
0!
0#
0*
0,
09
0>
0?
0C
#402730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#402740000000
0!
0*
09
0>
0C
#402750000000
1!
1*
19
1>
1C
#402760000000
0!
0*
09
0>
0C
#402770000000
1!
1*
19
1>
1C
#402780000000
0!
0*
09
0>
0C
#402790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#402800000000
0!
0*
09
0>
0C
#402810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#402820000000
0!
0*
09
0>
0C
#402830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#402840000000
0!
0*
09
0>
0C
#402850000000
1!
1*
b10 6
19
1>
1C
b10 G
#402860000000
0!
0*
09
0>
0C
#402870000000
1!
1*
b11 6
19
1>
1C
b11 G
#402880000000
0!
0*
09
0>
0C
#402890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#402900000000
0!
0*
09
0>
0C
#402910000000
1!
1*
b101 6
19
1>
1C
b101 G
#402920000000
0!
0*
09
0>
0C
#402930000000
1!
1*
b110 6
19
1>
1C
b110 G
#402940000000
0!
0*
09
0>
0C
#402950000000
1!
1*
b111 6
19
1>
1C
b111 G
#402960000000
0!
0*
09
0>
0C
#402970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#402980000000
0!
0*
09
0>
0C
#402990000000
1!
1*
b1 6
19
1>
1C
b1 G
#403000000000
0!
0*
09
0>
0C
#403010000000
1!
1*
b10 6
19
1>
1C
b10 G
#403020000000
0!
0*
09
0>
0C
#403030000000
1!
1*
b11 6
19
1>
1C
b11 G
#403040000000
0!
0*
09
0>
0C
#403050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#403060000000
0!
0*
09
0>
0C
#403070000000
1!
1*
b101 6
19
1>
1C
b101 G
#403080000000
0!
0*
09
0>
0C
#403090000000
1!
1*
b110 6
19
1>
1C
b110 G
#403100000000
0!
0*
09
0>
0C
#403110000000
1!
1*
b111 6
19
1>
1C
b111 G
#403120000000
0!
0*
09
0>
0C
#403130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#403140000000
0!
0*
09
0>
0C
#403150000000
1!
1*
b1 6
19
1>
1C
b1 G
#403160000000
0!
0*
09
0>
0C
#403170000000
1!
1*
b10 6
19
1>
1C
b10 G
#403180000000
0!
0*
09
0>
0C
#403190000000
1!
1*
b11 6
19
1>
1C
b11 G
#403200000000
0!
0*
09
0>
0C
#403210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#403220000000
0!
0*
09
0>
0C
#403230000000
1!
1*
b101 6
19
1>
1C
b101 G
#403240000000
0!
0*
09
0>
0C
#403250000000
1!
1*
b110 6
19
1>
1C
b110 G
#403260000000
0!
0*
09
0>
0C
#403270000000
1!
1*
b111 6
19
1>
1C
b111 G
#403280000000
0!
1"
0*
1+
09
1:
0>
0C
#403290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#403300000000
0!
0*
09
0>
0C
#403310000000
1!
1*
b1 6
19
1>
1C
b1 G
#403320000000
0!
0*
09
0>
0C
#403330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#403340000000
0!
0*
09
0>
0C
#403350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#403360000000
0!
0*
09
0>
0C
#403370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#403380000000
0!
0*
09
0>
0C
#403390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#403400000000
0!
0#
0*
0,
09
0>
0?
0C
#403410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#403420000000
0!
0*
09
0>
0C
#403430000000
1!
1*
19
1>
1C
#403440000000
0!
0*
09
0>
0C
#403450000000
1!
1*
19
1>
1C
#403460000000
0!
0*
09
0>
0C
#403470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#403480000000
0!
0*
09
0>
0C
#403490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#403500000000
0!
0*
09
0>
0C
#403510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#403520000000
0!
0*
09
0>
0C
#403530000000
1!
1*
b10 6
19
1>
1C
b10 G
#403540000000
0!
0*
09
0>
0C
#403550000000
1!
1*
b11 6
19
1>
1C
b11 G
#403560000000
0!
0*
09
0>
0C
#403570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#403580000000
0!
0*
09
0>
0C
#403590000000
1!
1*
b101 6
19
1>
1C
b101 G
#403600000000
0!
0*
09
0>
0C
#403610000000
1!
1*
b110 6
19
1>
1C
b110 G
#403620000000
0!
0*
09
0>
0C
#403630000000
1!
1*
b111 6
19
1>
1C
b111 G
#403640000000
0!
0*
09
0>
0C
#403650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#403660000000
0!
0*
09
0>
0C
#403670000000
1!
1*
b1 6
19
1>
1C
b1 G
#403680000000
0!
0*
09
0>
0C
#403690000000
1!
1*
b10 6
19
1>
1C
b10 G
#403700000000
0!
0*
09
0>
0C
#403710000000
1!
1*
b11 6
19
1>
1C
b11 G
#403720000000
0!
0*
09
0>
0C
#403730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#403740000000
0!
0*
09
0>
0C
#403750000000
1!
1*
b101 6
19
1>
1C
b101 G
#403760000000
0!
0*
09
0>
0C
#403770000000
1!
1*
b110 6
19
1>
1C
b110 G
#403780000000
0!
0*
09
0>
0C
#403790000000
1!
1*
b111 6
19
1>
1C
b111 G
#403800000000
0!
0*
09
0>
0C
#403810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#403820000000
0!
0*
09
0>
0C
#403830000000
1!
1*
b1 6
19
1>
1C
b1 G
#403840000000
0!
0*
09
0>
0C
#403850000000
1!
1*
b10 6
19
1>
1C
b10 G
#403860000000
0!
0*
09
0>
0C
#403870000000
1!
1*
b11 6
19
1>
1C
b11 G
#403880000000
0!
0*
09
0>
0C
#403890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#403900000000
0!
0*
09
0>
0C
#403910000000
1!
1*
b101 6
19
1>
1C
b101 G
#403920000000
0!
0*
09
0>
0C
#403930000000
1!
1*
b110 6
19
1>
1C
b110 G
#403940000000
0!
0*
09
0>
0C
#403950000000
1!
1*
b111 6
19
1>
1C
b111 G
#403960000000
0!
1"
0*
1+
09
1:
0>
0C
#403970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#403980000000
0!
0*
09
0>
0C
#403990000000
1!
1*
b1 6
19
1>
1C
b1 G
#404000000000
0!
0*
09
0>
0C
#404010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#404020000000
0!
0*
09
0>
0C
#404030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#404040000000
0!
0*
09
0>
0C
#404050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#404060000000
0!
0*
09
0>
0C
#404070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#404080000000
0!
0#
0*
0,
09
0>
0?
0C
#404090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#404100000000
0!
0*
09
0>
0C
#404110000000
1!
1*
19
1>
1C
#404120000000
0!
0*
09
0>
0C
#404130000000
1!
1*
19
1>
1C
#404140000000
0!
0*
09
0>
0C
#404150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#404160000000
0!
0*
09
0>
0C
#404170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#404180000000
0!
0*
09
0>
0C
#404190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#404200000000
0!
0*
09
0>
0C
#404210000000
1!
1*
b10 6
19
1>
1C
b10 G
#404220000000
0!
0*
09
0>
0C
#404230000000
1!
1*
b11 6
19
1>
1C
b11 G
#404240000000
0!
0*
09
0>
0C
#404250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#404260000000
0!
0*
09
0>
0C
#404270000000
1!
1*
b101 6
19
1>
1C
b101 G
#404280000000
0!
0*
09
0>
0C
#404290000000
1!
1*
b110 6
19
1>
1C
b110 G
#404300000000
0!
0*
09
0>
0C
#404310000000
1!
1*
b111 6
19
1>
1C
b111 G
#404320000000
0!
0*
09
0>
0C
#404330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#404340000000
0!
0*
09
0>
0C
#404350000000
1!
1*
b1 6
19
1>
1C
b1 G
#404360000000
0!
0*
09
0>
0C
#404370000000
1!
1*
b10 6
19
1>
1C
b10 G
#404380000000
0!
0*
09
0>
0C
#404390000000
1!
1*
b11 6
19
1>
1C
b11 G
#404400000000
0!
0*
09
0>
0C
#404410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#404420000000
0!
0*
09
0>
0C
#404430000000
1!
1*
b101 6
19
1>
1C
b101 G
#404440000000
0!
0*
09
0>
0C
#404450000000
1!
1*
b110 6
19
1>
1C
b110 G
#404460000000
0!
0*
09
0>
0C
#404470000000
1!
1*
b111 6
19
1>
1C
b111 G
#404480000000
0!
0*
09
0>
0C
#404490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#404500000000
0!
0*
09
0>
0C
#404510000000
1!
1*
b1 6
19
1>
1C
b1 G
#404520000000
0!
0*
09
0>
0C
#404530000000
1!
1*
b10 6
19
1>
1C
b10 G
#404540000000
0!
0*
09
0>
0C
#404550000000
1!
1*
b11 6
19
1>
1C
b11 G
#404560000000
0!
0*
09
0>
0C
#404570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#404580000000
0!
0*
09
0>
0C
#404590000000
1!
1*
b101 6
19
1>
1C
b101 G
#404600000000
0!
0*
09
0>
0C
#404610000000
1!
1*
b110 6
19
1>
1C
b110 G
#404620000000
0!
0*
09
0>
0C
#404630000000
1!
1*
b111 6
19
1>
1C
b111 G
#404640000000
0!
1"
0*
1+
09
1:
0>
0C
#404650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#404660000000
0!
0*
09
0>
0C
#404670000000
1!
1*
b1 6
19
1>
1C
b1 G
#404680000000
0!
0*
09
0>
0C
#404690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#404700000000
0!
0*
09
0>
0C
#404710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#404720000000
0!
0*
09
0>
0C
#404730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#404740000000
0!
0*
09
0>
0C
#404750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#404760000000
0!
0#
0*
0,
09
0>
0?
0C
#404770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#404780000000
0!
0*
09
0>
0C
#404790000000
1!
1*
19
1>
1C
#404800000000
0!
0*
09
0>
0C
#404810000000
1!
1*
19
1>
1C
#404820000000
0!
0*
09
0>
0C
#404830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#404840000000
0!
0*
09
0>
0C
#404850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#404860000000
0!
0*
09
0>
0C
#404870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#404880000000
0!
0*
09
0>
0C
#404890000000
1!
1*
b10 6
19
1>
1C
b10 G
#404900000000
0!
0*
09
0>
0C
#404910000000
1!
1*
b11 6
19
1>
1C
b11 G
#404920000000
0!
0*
09
0>
0C
#404930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#404940000000
0!
0*
09
0>
0C
#404950000000
1!
1*
b101 6
19
1>
1C
b101 G
#404960000000
0!
0*
09
0>
0C
#404970000000
1!
1*
b110 6
19
1>
1C
b110 G
#404980000000
0!
0*
09
0>
0C
#404990000000
1!
1*
b111 6
19
1>
1C
b111 G
#405000000000
0!
0*
09
0>
0C
#405010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#405020000000
0!
0*
09
0>
0C
#405030000000
1!
1*
b1 6
19
1>
1C
b1 G
#405040000000
0!
0*
09
0>
0C
#405050000000
1!
1*
b10 6
19
1>
1C
b10 G
#405060000000
0!
0*
09
0>
0C
#405070000000
1!
1*
b11 6
19
1>
1C
b11 G
#405080000000
0!
0*
09
0>
0C
#405090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#405100000000
0!
0*
09
0>
0C
#405110000000
1!
1*
b101 6
19
1>
1C
b101 G
#405120000000
0!
0*
09
0>
0C
#405130000000
1!
1*
b110 6
19
1>
1C
b110 G
#405140000000
0!
0*
09
0>
0C
#405150000000
1!
1*
b111 6
19
1>
1C
b111 G
#405160000000
0!
0*
09
0>
0C
#405170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#405180000000
0!
0*
09
0>
0C
#405190000000
1!
1*
b1 6
19
1>
1C
b1 G
#405200000000
0!
0*
09
0>
0C
#405210000000
1!
1*
b10 6
19
1>
1C
b10 G
#405220000000
0!
0*
09
0>
0C
#405230000000
1!
1*
b11 6
19
1>
1C
b11 G
#405240000000
0!
0*
09
0>
0C
#405250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#405260000000
0!
0*
09
0>
0C
#405270000000
1!
1*
b101 6
19
1>
1C
b101 G
#405280000000
0!
0*
09
0>
0C
#405290000000
1!
1*
b110 6
19
1>
1C
b110 G
#405300000000
0!
0*
09
0>
0C
#405310000000
1!
1*
b111 6
19
1>
1C
b111 G
#405320000000
0!
1"
0*
1+
09
1:
0>
0C
#405330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#405340000000
0!
0*
09
0>
0C
#405350000000
1!
1*
b1 6
19
1>
1C
b1 G
#405360000000
0!
0*
09
0>
0C
#405370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#405380000000
0!
0*
09
0>
0C
#405390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#405400000000
0!
0*
09
0>
0C
#405410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#405420000000
0!
0*
09
0>
0C
#405430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#405440000000
0!
0#
0*
0,
09
0>
0?
0C
#405450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#405460000000
0!
0*
09
0>
0C
#405470000000
1!
1*
19
1>
1C
#405480000000
0!
0*
09
0>
0C
#405490000000
1!
1*
19
1>
1C
#405500000000
0!
0*
09
0>
0C
#405510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#405520000000
0!
0*
09
0>
0C
#405530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#405540000000
0!
0*
09
0>
0C
#405550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#405560000000
0!
0*
09
0>
0C
#405570000000
1!
1*
b10 6
19
1>
1C
b10 G
#405580000000
0!
0*
09
0>
0C
#405590000000
1!
1*
b11 6
19
1>
1C
b11 G
#405600000000
0!
0*
09
0>
0C
#405610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#405620000000
0!
0*
09
0>
0C
#405630000000
1!
1*
b101 6
19
1>
1C
b101 G
#405640000000
0!
0*
09
0>
0C
#405650000000
1!
1*
b110 6
19
1>
1C
b110 G
#405660000000
0!
0*
09
0>
0C
#405670000000
1!
1*
b111 6
19
1>
1C
b111 G
#405680000000
0!
0*
09
0>
0C
#405690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#405700000000
0!
0*
09
0>
0C
#405710000000
1!
1*
b1 6
19
1>
1C
b1 G
#405720000000
0!
0*
09
0>
0C
#405730000000
1!
1*
b10 6
19
1>
1C
b10 G
#405740000000
0!
0*
09
0>
0C
#405750000000
1!
1*
b11 6
19
1>
1C
b11 G
#405760000000
0!
0*
09
0>
0C
#405770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#405780000000
0!
0*
09
0>
0C
#405790000000
1!
1*
b101 6
19
1>
1C
b101 G
#405800000000
0!
0*
09
0>
0C
#405810000000
1!
1*
b110 6
19
1>
1C
b110 G
#405820000000
0!
0*
09
0>
0C
#405830000000
1!
1*
b111 6
19
1>
1C
b111 G
#405840000000
0!
0*
09
0>
0C
#405850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#405860000000
0!
0*
09
0>
0C
#405870000000
1!
1*
b1 6
19
1>
1C
b1 G
#405880000000
0!
0*
09
0>
0C
#405890000000
1!
1*
b10 6
19
1>
1C
b10 G
#405900000000
0!
0*
09
0>
0C
#405910000000
1!
1*
b11 6
19
1>
1C
b11 G
#405920000000
0!
0*
09
0>
0C
#405930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#405940000000
0!
0*
09
0>
0C
#405950000000
1!
1*
b101 6
19
1>
1C
b101 G
#405960000000
0!
0*
09
0>
0C
#405970000000
1!
1*
b110 6
19
1>
1C
b110 G
#405980000000
0!
0*
09
0>
0C
#405990000000
1!
1*
b111 6
19
1>
1C
b111 G
#406000000000
0!
1"
0*
1+
09
1:
0>
0C
#406010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#406020000000
0!
0*
09
0>
0C
#406030000000
1!
1*
b1 6
19
1>
1C
b1 G
#406040000000
0!
0*
09
0>
0C
#406050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#406060000000
0!
0*
09
0>
0C
#406070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#406080000000
0!
0*
09
0>
0C
#406090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#406100000000
0!
0*
09
0>
0C
#406110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#406120000000
0!
0#
0*
0,
09
0>
0?
0C
#406130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#406140000000
0!
0*
09
0>
0C
#406150000000
1!
1*
19
1>
1C
#406160000000
0!
0*
09
0>
0C
#406170000000
1!
1*
19
1>
1C
#406180000000
0!
0*
09
0>
0C
#406190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#406200000000
0!
0*
09
0>
0C
#406210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#406220000000
0!
0*
09
0>
0C
#406230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#406240000000
0!
0*
09
0>
0C
#406250000000
1!
1*
b10 6
19
1>
1C
b10 G
#406260000000
0!
0*
09
0>
0C
#406270000000
1!
1*
b11 6
19
1>
1C
b11 G
#406280000000
0!
0*
09
0>
0C
#406290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#406300000000
0!
0*
09
0>
0C
#406310000000
1!
1*
b101 6
19
1>
1C
b101 G
#406320000000
0!
0*
09
0>
0C
#406330000000
1!
1*
b110 6
19
1>
1C
b110 G
#406340000000
0!
0*
09
0>
0C
#406350000000
1!
1*
b111 6
19
1>
1C
b111 G
#406360000000
0!
0*
09
0>
0C
#406370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#406380000000
0!
0*
09
0>
0C
#406390000000
1!
1*
b1 6
19
1>
1C
b1 G
#406400000000
0!
0*
09
0>
0C
#406410000000
1!
1*
b10 6
19
1>
1C
b10 G
#406420000000
0!
0*
09
0>
0C
#406430000000
1!
1*
b11 6
19
1>
1C
b11 G
#406440000000
0!
0*
09
0>
0C
#406450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#406460000000
0!
0*
09
0>
0C
#406470000000
1!
1*
b101 6
19
1>
1C
b101 G
#406480000000
0!
0*
09
0>
0C
#406490000000
1!
1*
b110 6
19
1>
1C
b110 G
#406500000000
0!
0*
09
0>
0C
#406510000000
1!
1*
b111 6
19
1>
1C
b111 G
#406520000000
0!
0*
09
0>
0C
#406530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#406540000000
0!
0*
09
0>
0C
#406550000000
1!
1*
b1 6
19
1>
1C
b1 G
#406560000000
0!
0*
09
0>
0C
#406570000000
1!
1*
b10 6
19
1>
1C
b10 G
#406580000000
0!
0*
09
0>
0C
#406590000000
1!
1*
b11 6
19
1>
1C
b11 G
#406600000000
0!
0*
09
0>
0C
#406610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#406620000000
0!
0*
09
0>
0C
#406630000000
1!
1*
b101 6
19
1>
1C
b101 G
#406640000000
0!
0*
09
0>
0C
#406650000000
1!
1*
b110 6
19
1>
1C
b110 G
#406660000000
0!
0*
09
0>
0C
#406670000000
1!
1*
b111 6
19
1>
1C
b111 G
#406680000000
0!
1"
0*
1+
09
1:
0>
0C
#406690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#406700000000
0!
0*
09
0>
0C
#406710000000
1!
1*
b1 6
19
1>
1C
b1 G
#406720000000
0!
0*
09
0>
0C
#406730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#406740000000
0!
0*
09
0>
0C
#406750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#406760000000
0!
0*
09
0>
0C
#406770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#406780000000
0!
0*
09
0>
0C
#406790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#406800000000
0!
0#
0*
0,
09
0>
0?
0C
#406810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#406820000000
0!
0*
09
0>
0C
#406830000000
1!
1*
19
1>
1C
#406840000000
0!
0*
09
0>
0C
#406850000000
1!
1*
19
1>
1C
#406860000000
0!
0*
09
0>
0C
#406870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#406880000000
0!
0*
09
0>
0C
#406890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#406900000000
0!
0*
09
0>
0C
#406910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#406920000000
0!
0*
09
0>
0C
#406930000000
1!
1*
b10 6
19
1>
1C
b10 G
#406940000000
0!
0*
09
0>
0C
#406950000000
1!
1*
b11 6
19
1>
1C
b11 G
#406960000000
0!
0*
09
0>
0C
#406970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#406980000000
0!
0*
09
0>
0C
#406990000000
1!
1*
b101 6
19
1>
1C
b101 G
#407000000000
0!
0*
09
0>
0C
#407010000000
1!
1*
b110 6
19
1>
1C
b110 G
#407020000000
0!
0*
09
0>
0C
#407030000000
1!
1*
b111 6
19
1>
1C
b111 G
#407040000000
0!
0*
09
0>
0C
#407050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#407060000000
0!
0*
09
0>
0C
#407070000000
1!
1*
b1 6
19
1>
1C
b1 G
#407080000000
0!
0*
09
0>
0C
#407090000000
1!
1*
b10 6
19
1>
1C
b10 G
#407100000000
0!
0*
09
0>
0C
#407110000000
1!
1*
b11 6
19
1>
1C
b11 G
#407120000000
0!
0*
09
0>
0C
#407130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#407140000000
0!
0*
09
0>
0C
#407150000000
1!
1*
b101 6
19
1>
1C
b101 G
#407160000000
0!
0*
09
0>
0C
#407170000000
1!
1*
b110 6
19
1>
1C
b110 G
#407180000000
0!
0*
09
0>
0C
#407190000000
1!
1*
b111 6
19
1>
1C
b111 G
#407200000000
0!
0*
09
0>
0C
#407210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#407220000000
0!
0*
09
0>
0C
#407230000000
1!
1*
b1 6
19
1>
1C
b1 G
#407240000000
0!
0*
09
0>
0C
#407250000000
1!
1*
b10 6
19
1>
1C
b10 G
#407260000000
0!
0*
09
0>
0C
#407270000000
1!
1*
b11 6
19
1>
1C
b11 G
#407280000000
0!
0*
09
0>
0C
#407290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#407300000000
0!
0*
09
0>
0C
#407310000000
1!
1*
b101 6
19
1>
1C
b101 G
#407320000000
0!
0*
09
0>
0C
#407330000000
1!
1*
b110 6
19
1>
1C
b110 G
#407340000000
0!
0*
09
0>
0C
#407350000000
1!
1*
b111 6
19
1>
1C
b111 G
#407360000000
0!
1"
0*
1+
09
1:
0>
0C
#407370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#407380000000
0!
0*
09
0>
0C
#407390000000
1!
1*
b1 6
19
1>
1C
b1 G
#407400000000
0!
0*
09
0>
0C
#407410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#407420000000
0!
0*
09
0>
0C
#407430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#407440000000
0!
0*
09
0>
0C
#407450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#407460000000
0!
0*
09
0>
0C
#407470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#407480000000
0!
0#
0*
0,
09
0>
0?
0C
#407490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#407500000000
0!
0*
09
0>
0C
#407510000000
1!
1*
19
1>
1C
#407520000000
0!
0*
09
0>
0C
#407530000000
1!
1*
19
1>
1C
#407540000000
0!
0*
09
0>
0C
#407550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#407560000000
0!
0*
09
0>
0C
#407570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#407580000000
0!
0*
09
0>
0C
#407590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#407600000000
0!
0*
09
0>
0C
#407610000000
1!
1*
b10 6
19
1>
1C
b10 G
#407620000000
0!
0*
09
0>
0C
#407630000000
1!
1*
b11 6
19
1>
1C
b11 G
#407640000000
0!
0*
09
0>
0C
#407650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#407660000000
0!
0*
09
0>
0C
#407670000000
1!
1*
b101 6
19
1>
1C
b101 G
#407680000000
0!
0*
09
0>
0C
#407690000000
1!
1*
b110 6
19
1>
1C
b110 G
#407700000000
0!
0*
09
0>
0C
#407710000000
1!
1*
b111 6
19
1>
1C
b111 G
#407720000000
0!
0*
09
0>
0C
#407730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#407740000000
0!
0*
09
0>
0C
#407750000000
1!
1*
b1 6
19
1>
1C
b1 G
#407760000000
0!
0*
09
0>
0C
#407770000000
1!
1*
b10 6
19
1>
1C
b10 G
#407780000000
0!
0*
09
0>
0C
#407790000000
1!
1*
b11 6
19
1>
1C
b11 G
#407800000000
0!
0*
09
0>
0C
#407810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#407820000000
0!
0*
09
0>
0C
#407830000000
1!
1*
b101 6
19
1>
1C
b101 G
#407840000000
0!
0*
09
0>
0C
#407850000000
1!
1*
b110 6
19
1>
1C
b110 G
#407860000000
0!
0*
09
0>
0C
#407870000000
1!
1*
b111 6
19
1>
1C
b111 G
#407880000000
0!
0*
09
0>
0C
#407890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#407900000000
0!
0*
09
0>
0C
#407910000000
1!
1*
b1 6
19
1>
1C
b1 G
#407920000000
0!
0*
09
0>
0C
#407930000000
1!
1*
b10 6
19
1>
1C
b10 G
#407940000000
0!
0*
09
0>
0C
#407950000000
1!
1*
b11 6
19
1>
1C
b11 G
#407960000000
0!
0*
09
0>
0C
#407970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#407980000000
0!
0*
09
0>
0C
#407990000000
1!
1*
b101 6
19
1>
1C
b101 G
#408000000000
0!
0*
09
0>
0C
#408010000000
1!
1*
b110 6
19
1>
1C
b110 G
#408020000000
0!
0*
09
0>
0C
#408030000000
1!
1*
b111 6
19
1>
1C
b111 G
#408040000000
0!
1"
0*
1+
09
1:
0>
0C
#408050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#408060000000
0!
0*
09
0>
0C
#408070000000
1!
1*
b1 6
19
1>
1C
b1 G
#408080000000
0!
0*
09
0>
0C
#408090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#408100000000
0!
0*
09
0>
0C
#408110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#408120000000
0!
0*
09
0>
0C
#408130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#408140000000
0!
0*
09
0>
0C
#408150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#408160000000
0!
0#
0*
0,
09
0>
0?
0C
#408170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#408180000000
0!
0*
09
0>
0C
#408190000000
1!
1*
19
1>
1C
#408200000000
0!
0*
09
0>
0C
#408210000000
1!
1*
19
1>
1C
#408220000000
0!
0*
09
0>
0C
#408230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#408240000000
0!
0*
09
0>
0C
#408250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#408260000000
0!
0*
09
0>
0C
#408270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#408280000000
0!
0*
09
0>
0C
#408290000000
1!
1*
b10 6
19
1>
1C
b10 G
#408300000000
0!
0*
09
0>
0C
#408310000000
1!
1*
b11 6
19
1>
1C
b11 G
#408320000000
0!
0*
09
0>
0C
#408330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#408340000000
0!
0*
09
0>
0C
#408350000000
1!
1*
b101 6
19
1>
1C
b101 G
#408360000000
0!
0*
09
0>
0C
#408370000000
1!
1*
b110 6
19
1>
1C
b110 G
#408380000000
0!
0*
09
0>
0C
#408390000000
1!
1*
b111 6
19
1>
1C
b111 G
#408400000000
0!
0*
09
0>
0C
#408410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#408420000000
0!
0*
09
0>
0C
#408430000000
1!
1*
b1 6
19
1>
1C
b1 G
#408440000000
0!
0*
09
0>
0C
#408450000000
1!
1*
b10 6
19
1>
1C
b10 G
#408460000000
0!
0*
09
0>
0C
#408470000000
1!
1*
b11 6
19
1>
1C
b11 G
#408480000000
0!
0*
09
0>
0C
#408490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#408500000000
0!
0*
09
0>
0C
#408510000000
1!
1*
b101 6
19
1>
1C
b101 G
#408520000000
0!
0*
09
0>
0C
#408530000000
1!
1*
b110 6
19
1>
1C
b110 G
#408540000000
0!
0*
09
0>
0C
#408550000000
1!
1*
b111 6
19
1>
1C
b111 G
#408560000000
0!
0*
09
0>
0C
#408570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#408580000000
0!
0*
09
0>
0C
#408590000000
1!
1*
b1 6
19
1>
1C
b1 G
#408600000000
0!
0*
09
0>
0C
#408610000000
1!
1*
b10 6
19
1>
1C
b10 G
#408620000000
0!
0*
09
0>
0C
#408630000000
1!
1*
b11 6
19
1>
1C
b11 G
#408640000000
0!
0*
09
0>
0C
#408650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#408660000000
0!
0*
09
0>
0C
#408670000000
1!
1*
b101 6
19
1>
1C
b101 G
#408680000000
0!
0*
09
0>
0C
#408690000000
1!
1*
b110 6
19
1>
1C
b110 G
#408700000000
0!
0*
09
0>
0C
#408710000000
1!
1*
b111 6
19
1>
1C
b111 G
#408720000000
0!
1"
0*
1+
09
1:
0>
0C
#408730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#408740000000
0!
0*
09
0>
0C
#408750000000
1!
1*
b1 6
19
1>
1C
b1 G
#408760000000
0!
0*
09
0>
0C
#408770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#408780000000
0!
0*
09
0>
0C
#408790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#408800000000
0!
0*
09
0>
0C
#408810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#408820000000
0!
0*
09
0>
0C
#408830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#408840000000
0!
0#
0*
0,
09
0>
0?
0C
#408850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#408860000000
0!
0*
09
0>
0C
#408870000000
1!
1*
19
1>
1C
#408880000000
0!
0*
09
0>
0C
#408890000000
1!
1*
19
1>
1C
#408900000000
0!
0*
09
0>
0C
#408910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#408920000000
0!
0*
09
0>
0C
#408930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#408940000000
0!
0*
09
0>
0C
#408950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#408960000000
0!
0*
09
0>
0C
#408970000000
1!
1*
b10 6
19
1>
1C
b10 G
#408980000000
0!
0*
09
0>
0C
#408990000000
1!
1*
b11 6
19
1>
1C
b11 G
#409000000000
0!
0*
09
0>
0C
#409010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#409020000000
0!
0*
09
0>
0C
#409030000000
1!
1*
b101 6
19
1>
1C
b101 G
#409040000000
0!
0*
09
0>
0C
#409050000000
1!
1*
b110 6
19
1>
1C
b110 G
#409060000000
0!
0*
09
0>
0C
#409070000000
1!
1*
b111 6
19
1>
1C
b111 G
#409080000000
0!
0*
09
0>
0C
#409090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#409100000000
0!
0*
09
0>
0C
#409110000000
1!
1*
b1 6
19
1>
1C
b1 G
#409120000000
0!
0*
09
0>
0C
#409130000000
1!
1*
b10 6
19
1>
1C
b10 G
#409140000000
0!
0*
09
0>
0C
#409150000000
1!
1*
b11 6
19
1>
1C
b11 G
#409160000000
0!
0*
09
0>
0C
#409170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#409180000000
0!
0*
09
0>
0C
#409190000000
1!
1*
b101 6
19
1>
1C
b101 G
#409200000000
0!
0*
09
0>
0C
#409210000000
1!
1*
b110 6
19
1>
1C
b110 G
#409220000000
0!
0*
09
0>
0C
#409230000000
1!
1*
b111 6
19
1>
1C
b111 G
#409240000000
0!
0*
09
0>
0C
#409250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#409260000000
0!
0*
09
0>
0C
#409270000000
1!
1*
b1 6
19
1>
1C
b1 G
#409280000000
0!
0*
09
0>
0C
#409290000000
1!
1*
b10 6
19
1>
1C
b10 G
#409300000000
0!
0*
09
0>
0C
#409310000000
1!
1*
b11 6
19
1>
1C
b11 G
#409320000000
0!
0*
09
0>
0C
#409330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#409340000000
0!
0*
09
0>
0C
#409350000000
1!
1*
b101 6
19
1>
1C
b101 G
#409360000000
0!
0*
09
0>
0C
#409370000000
1!
1*
b110 6
19
1>
1C
b110 G
#409380000000
0!
0*
09
0>
0C
#409390000000
1!
1*
b111 6
19
1>
1C
b111 G
#409400000000
0!
1"
0*
1+
09
1:
0>
0C
#409410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#409420000000
0!
0*
09
0>
0C
#409430000000
1!
1*
b1 6
19
1>
1C
b1 G
#409440000000
0!
0*
09
0>
0C
#409450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#409460000000
0!
0*
09
0>
0C
#409470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#409480000000
0!
0*
09
0>
0C
#409490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#409500000000
0!
0*
09
0>
0C
#409510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#409520000000
0!
0#
0*
0,
09
0>
0?
0C
#409530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#409540000000
0!
0*
09
0>
0C
#409550000000
1!
1*
19
1>
1C
#409560000000
0!
0*
09
0>
0C
#409570000000
1!
1*
19
1>
1C
#409580000000
0!
0*
09
0>
0C
#409590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#409600000000
0!
0*
09
0>
0C
#409610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#409620000000
0!
0*
09
0>
0C
#409630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#409640000000
0!
0*
09
0>
0C
#409650000000
1!
1*
b10 6
19
1>
1C
b10 G
#409660000000
0!
0*
09
0>
0C
#409670000000
1!
1*
b11 6
19
1>
1C
b11 G
#409680000000
0!
0*
09
0>
0C
#409690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#409700000000
0!
0*
09
0>
0C
#409710000000
1!
1*
b101 6
19
1>
1C
b101 G
#409720000000
0!
0*
09
0>
0C
#409730000000
1!
1*
b110 6
19
1>
1C
b110 G
#409740000000
0!
0*
09
0>
0C
#409750000000
1!
1*
b111 6
19
1>
1C
b111 G
#409760000000
0!
0*
09
0>
0C
#409770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#409780000000
0!
0*
09
0>
0C
#409790000000
1!
1*
b1 6
19
1>
1C
b1 G
#409800000000
0!
0*
09
0>
0C
#409810000000
1!
1*
b10 6
19
1>
1C
b10 G
#409820000000
0!
0*
09
0>
0C
#409830000000
1!
1*
b11 6
19
1>
1C
b11 G
#409840000000
0!
0*
09
0>
0C
#409850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#409860000000
0!
0*
09
0>
0C
#409870000000
1!
1*
b101 6
19
1>
1C
b101 G
#409880000000
0!
0*
09
0>
0C
#409890000000
1!
1*
b110 6
19
1>
1C
b110 G
#409900000000
0!
0*
09
0>
0C
#409910000000
1!
1*
b111 6
19
1>
1C
b111 G
#409920000000
0!
0*
09
0>
0C
#409930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#409940000000
0!
0*
09
0>
0C
#409950000000
1!
1*
b1 6
19
1>
1C
b1 G
#409960000000
0!
0*
09
0>
0C
#409970000000
1!
1*
b10 6
19
1>
1C
b10 G
#409980000000
0!
0*
09
0>
0C
#409990000000
1!
1*
b11 6
19
1>
1C
b11 G
#410000000000
0!
0*
09
0>
0C
#410010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#410020000000
0!
0*
09
0>
0C
#410030000000
1!
1*
b101 6
19
1>
1C
b101 G
#410040000000
0!
0*
09
0>
0C
#410050000000
1!
1*
b110 6
19
1>
1C
b110 G
#410060000000
0!
0*
09
0>
0C
#410070000000
1!
1*
b111 6
19
1>
1C
b111 G
#410080000000
0!
1"
0*
1+
09
1:
0>
0C
#410090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#410100000000
0!
0*
09
0>
0C
#410110000000
1!
1*
b1 6
19
1>
1C
b1 G
#410120000000
0!
0*
09
0>
0C
#410130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#410140000000
0!
0*
09
0>
0C
#410150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#410160000000
0!
0*
09
0>
0C
#410170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#410180000000
0!
0*
09
0>
0C
#410190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#410200000000
0!
0#
0*
0,
09
0>
0?
0C
#410210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#410220000000
0!
0*
09
0>
0C
#410230000000
1!
1*
19
1>
1C
#410240000000
0!
0*
09
0>
0C
#410250000000
1!
1*
19
1>
1C
#410260000000
0!
0*
09
0>
0C
#410270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#410280000000
0!
0*
09
0>
0C
#410290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#410300000000
0!
0*
09
0>
0C
#410310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#410320000000
0!
0*
09
0>
0C
#410330000000
1!
1*
b10 6
19
1>
1C
b10 G
#410340000000
0!
0*
09
0>
0C
#410350000000
1!
1*
b11 6
19
1>
1C
b11 G
#410360000000
0!
0*
09
0>
0C
#410370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#410380000000
0!
0*
09
0>
0C
#410390000000
1!
1*
b101 6
19
1>
1C
b101 G
#410400000000
0!
0*
09
0>
0C
#410410000000
1!
1*
b110 6
19
1>
1C
b110 G
#410420000000
0!
0*
09
0>
0C
#410430000000
1!
1*
b111 6
19
1>
1C
b111 G
#410440000000
0!
0*
09
0>
0C
#410450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#410460000000
0!
0*
09
0>
0C
#410470000000
1!
1*
b1 6
19
1>
1C
b1 G
#410480000000
0!
0*
09
0>
0C
#410490000000
1!
1*
b10 6
19
1>
1C
b10 G
#410500000000
0!
0*
09
0>
0C
#410510000000
1!
1*
b11 6
19
1>
1C
b11 G
#410520000000
0!
0*
09
0>
0C
#410530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#410540000000
0!
0*
09
0>
0C
#410550000000
1!
1*
b101 6
19
1>
1C
b101 G
#410560000000
0!
0*
09
0>
0C
#410570000000
1!
1*
b110 6
19
1>
1C
b110 G
#410580000000
0!
0*
09
0>
0C
#410590000000
1!
1*
b111 6
19
1>
1C
b111 G
#410600000000
0!
0*
09
0>
0C
#410610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#410620000000
0!
0*
09
0>
0C
#410630000000
1!
1*
b1 6
19
1>
1C
b1 G
#410640000000
0!
0*
09
0>
0C
#410650000000
1!
1*
b10 6
19
1>
1C
b10 G
#410660000000
0!
0*
09
0>
0C
#410670000000
1!
1*
b11 6
19
1>
1C
b11 G
#410680000000
0!
0*
09
0>
0C
#410690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#410700000000
0!
0*
09
0>
0C
#410710000000
1!
1*
b101 6
19
1>
1C
b101 G
#410720000000
0!
0*
09
0>
0C
#410730000000
1!
1*
b110 6
19
1>
1C
b110 G
#410740000000
0!
0*
09
0>
0C
#410750000000
1!
1*
b111 6
19
1>
1C
b111 G
#410760000000
0!
1"
0*
1+
09
1:
0>
0C
#410770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#410780000000
0!
0*
09
0>
0C
#410790000000
1!
1*
b1 6
19
1>
1C
b1 G
#410800000000
0!
0*
09
0>
0C
#410810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#410820000000
0!
0*
09
0>
0C
#410830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#410840000000
0!
0*
09
0>
0C
#410850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#410860000000
0!
0*
09
0>
0C
#410870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#410880000000
0!
0#
0*
0,
09
0>
0?
0C
#410890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#410900000000
0!
0*
09
0>
0C
#410910000000
1!
1*
19
1>
1C
#410920000000
0!
0*
09
0>
0C
#410930000000
1!
1*
19
1>
1C
#410940000000
0!
0*
09
0>
0C
#410950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#410960000000
0!
0*
09
0>
0C
#410970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#410980000000
0!
0*
09
0>
0C
#410990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#411000000000
0!
0*
09
0>
0C
#411010000000
1!
1*
b10 6
19
1>
1C
b10 G
#411020000000
0!
0*
09
0>
0C
#411030000000
1!
1*
b11 6
19
1>
1C
b11 G
#411040000000
0!
0*
09
0>
0C
#411050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#411060000000
0!
0*
09
0>
0C
#411070000000
1!
1*
b101 6
19
1>
1C
b101 G
#411080000000
0!
0*
09
0>
0C
#411090000000
1!
1*
b110 6
19
1>
1C
b110 G
#411100000000
0!
0*
09
0>
0C
#411110000000
1!
1*
b111 6
19
1>
1C
b111 G
#411120000000
0!
0*
09
0>
0C
#411130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#411140000000
0!
0*
09
0>
0C
#411150000000
1!
1*
b1 6
19
1>
1C
b1 G
#411160000000
0!
0*
09
0>
0C
#411170000000
1!
1*
b10 6
19
1>
1C
b10 G
#411180000000
0!
0*
09
0>
0C
#411190000000
1!
1*
b11 6
19
1>
1C
b11 G
#411200000000
0!
0*
09
0>
0C
#411210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#411220000000
0!
0*
09
0>
0C
#411230000000
1!
1*
b101 6
19
1>
1C
b101 G
#411240000000
0!
0*
09
0>
0C
#411250000000
1!
1*
b110 6
19
1>
1C
b110 G
#411260000000
0!
0*
09
0>
0C
#411270000000
1!
1*
b111 6
19
1>
1C
b111 G
#411280000000
0!
0*
09
0>
0C
#411290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#411300000000
0!
0*
09
0>
0C
#411310000000
1!
1*
b1 6
19
1>
1C
b1 G
#411320000000
0!
0*
09
0>
0C
#411330000000
1!
1*
b10 6
19
1>
1C
b10 G
#411340000000
0!
0*
09
0>
0C
#411350000000
1!
1*
b11 6
19
1>
1C
b11 G
#411360000000
0!
0*
09
0>
0C
#411370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#411380000000
0!
0*
09
0>
0C
#411390000000
1!
1*
b101 6
19
1>
1C
b101 G
#411400000000
0!
0*
09
0>
0C
#411410000000
1!
1*
b110 6
19
1>
1C
b110 G
#411420000000
0!
0*
09
0>
0C
#411430000000
1!
1*
b111 6
19
1>
1C
b111 G
#411440000000
0!
1"
0*
1+
09
1:
0>
0C
#411450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#411460000000
0!
0*
09
0>
0C
#411470000000
1!
1*
b1 6
19
1>
1C
b1 G
#411480000000
0!
0*
09
0>
0C
#411490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#411500000000
0!
0*
09
0>
0C
#411510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#411520000000
0!
0*
09
0>
0C
#411530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#411540000000
0!
0*
09
0>
0C
#411550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#411560000000
0!
0#
0*
0,
09
0>
0?
0C
#411570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#411580000000
0!
0*
09
0>
0C
#411590000000
1!
1*
19
1>
1C
#411600000000
0!
0*
09
0>
0C
#411610000000
1!
1*
19
1>
1C
#411620000000
0!
0*
09
0>
0C
#411630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#411640000000
0!
0*
09
0>
0C
#411650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#411660000000
0!
0*
09
0>
0C
#411670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#411680000000
0!
0*
09
0>
0C
#411690000000
1!
1*
b10 6
19
1>
1C
b10 G
#411700000000
0!
0*
09
0>
0C
#411710000000
1!
1*
b11 6
19
1>
1C
b11 G
#411720000000
0!
0*
09
0>
0C
#411730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#411740000000
0!
0*
09
0>
0C
#411750000000
1!
1*
b101 6
19
1>
1C
b101 G
#411760000000
0!
0*
09
0>
0C
#411770000000
1!
1*
b110 6
19
1>
1C
b110 G
#411780000000
0!
0*
09
0>
0C
#411790000000
1!
1*
b111 6
19
1>
1C
b111 G
#411800000000
0!
0*
09
0>
0C
#411810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#411820000000
0!
0*
09
0>
0C
#411830000000
1!
1*
b1 6
19
1>
1C
b1 G
#411840000000
0!
0*
09
0>
0C
#411850000000
1!
1*
b10 6
19
1>
1C
b10 G
#411860000000
0!
0*
09
0>
0C
#411870000000
1!
1*
b11 6
19
1>
1C
b11 G
#411880000000
0!
0*
09
0>
0C
#411890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#411900000000
0!
0*
09
0>
0C
#411910000000
1!
1*
b101 6
19
1>
1C
b101 G
#411920000000
0!
0*
09
0>
0C
#411930000000
1!
1*
b110 6
19
1>
1C
b110 G
#411940000000
0!
0*
09
0>
0C
#411950000000
1!
1*
b111 6
19
1>
1C
b111 G
#411960000000
0!
0*
09
0>
0C
#411970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#411980000000
0!
0*
09
0>
0C
#411990000000
1!
1*
b1 6
19
1>
1C
b1 G
#412000000000
0!
0*
09
0>
0C
#412010000000
1!
1*
b10 6
19
1>
1C
b10 G
#412020000000
0!
0*
09
0>
0C
#412030000000
1!
1*
b11 6
19
1>
1C
b11 G
#412040000000
0!
0*
09
0>
0C
#412050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#412060000000
0!
0*
09
0>
0C
#412070000000
1!
1*
b101 6
19
1>
1C
b101 G
#412080000000
0!
0*
09
0>
0C
#412090000000
1!
1*
b110 6
19
1>
1C
b110 G
#412100000000
0!
0*
09
0>
0C
#412110000000
1!
1*
b111 6
19
1>
1C
b111 G
#412120000000
0!
1"
0*
1+
09
1:
0>
0C
#412130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#412140000000
0!
0*
09
0>
0C
#412150000000
1!
1*
b1 6
19
1>
1C
b1 G
#412160000000
0!
0*
09
0>
0C
#412170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#412180000000
0!
0*
09
0>
0C
#412190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#412200000000
0!
0*
09
0>
0C
#412210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#412220000000
0!
0*
09
0>
0C
#412230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#412240000000
0!
0#
0*
0,
09
0>
0?
0C
#412250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#412260000000
0!
0*
09
0>
0C
#412270000000
1!
1*
19
1>
1C
#412280000000
0!
0*
09
0>
0C
#412290000000
1!
1*
19
1>
1C
#412300000000
0!
0*
09
0>
0C
#412310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#412320000000
0!
0*
09
0>
0C
#412330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#412340000000
0!
0*
09
0>
0C
#412350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#412360000000
0!
0*
09
0>
0C
#412370000000
1!
1*
b10 6
19
1>
1C
b10 G
#412380000000
0!
0*
09
0>
0C
#412390000000
1!
1*
b11 6
19
1>
1C
b11 G
#412400000000
0!
0*
09
0>
0C
#412410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#412420000000
0!
0*
09
0>
0C
#412430000000
1!
1*
b101 6
19
1>
1C
b101 G
#412440000000
0!
0*
09
0>
0C
#412450000000
1!
1*
b110 6
19
1>
1C
b110 G
#412460000000
0!
0*
09
0>
0C
#412470000000
1!
1*
b111 6
19
1>
1C
b111 G
#412480000000
0!
0*
09
0>
0C
#412490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#412500000000
0!
0*
09
0>
0C
#412510000000
1!
1*
b1 6
19
1>
1C
b1 G
#412520000000
0!
0*
09
0>
0C
#412530000000
1!
1*
b10 6
19
1>
1C
b10 G
#412540000000
0!
0*
09
0>
0C
#412550000000
1!
1*
b11 6
19
1>
1C
b11 G
#412560000000
0!
0*
09
0>
0C
#412570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#412580000000
0!
0*
09
0>
0C
#412590000000
1!
1*
b101 6
19
1>
1C
b101 G
#412600000000
0!
0*
09
0>
0C
#412610000000
1!
1*
b110 6
19
1>
1C
b110 G
#412620000000
0!
0*
09
0>
0C
#412630000000
1!
1*
b111 6
19
1>
1C
b111 G
#412640000000
0!
0*
09
0>
0C
#412650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#412660000000
0!
0*
09
0>
0C
#412670000000
1!
1*
b1 6
19
1>
1C
b1 G
#412680000000
0!
0*
09
0>
0C
#412690000000
1!
1*
b10 6
19
1>
1C
b10 G
#412700000000
0!
0*
09
0>
0C
#412710000000
1!
1*
b11 6
19
1>
1C
b11 G
#412720000000
0!
0*
09
0>
0C
#412730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#412740000000
0!
0*
09
0>
0C
#412750000000
1!
1*
b101 6
19
1>
1C
b101 G
#412760000000
0!
0*
09
0>
0C
#412770000000
1!
1*
b110 6
19
1>
1C
b110 G
#412780000000
0!
0*
09
0>
0C
#412790000000
1!
1*
b111 6
19
1>
1C
b111 G
#412800000000
0!
1"
0*
1+
09
1:
0>
0C
#412810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#412820000000
0!
0*
09
0>
0C
#412830000000
1!
1*
b1 6
19
1>
1C
b1 G
#412840000000
0!
0*
09
0>
0C
#412850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#412860000000
0!
0*
09
0>
0C
#412870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#412880000000
0!
0*
09
0>
0C
#412890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#412900000000
0!
0*
09
0>
0C
#412910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#412920000000
0!
0#
0*
0,
09
0>
0?
0C
#412930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#412940000000
0!
0*
09
0>
0C
#412950000000
1!
1*
19
1>
1C
#412960000000
0!
0*
09
0>
0C
#412970000000
1!
1*
19
1>
1C
#412980000000
0!
0*
09
0>
0C
#412990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#413000000000
0!
0*
09
0>
0C
#413010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#413020000000
0!
0*
09
0>
0C
#413030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#413040000000
0!
0*
09
0>
0C
#413050000000
1!
1*
b10 6
19
1>
1C
b10 G
#413060000000
0!
0*
09
0>
0C
#413070000000
1!
1*
b11 6
19
1>
1C
b11 G
#413080000000
0!
0*
09
0>
0C
#413090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#413100000000
0!
0*
09
0>
0C
#413110000000
1!
1*
b101 6
19
1>
1C
b101 G
#413120000000
0!
0*
09
0>
0C
#413130000000
1!
1*
b110 6
19
1>
1C
b110 G
#413140000000
0!
0*
09
0>
0C
#413150000000
1!
1*
b111 6
19
1>
1C
b111 G
#413160000000
0!
0*
09
0>
0C
#413170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#413180000000
0!
0*
09
0>
0C
#413190000000
1!
1*
b1 6
19
1>
1C
b1 G
#413200000000
0!
0*
09
0>
0C
#413210000000
1!
1*
b10 6
19
1>
1C
b10 G
#413220000000
0!
0*
09
0>
0C
#413230000000
1!
1*
b11 6
19
1>
1C
b11 G
#413240000000
0!
0*
09
0>
0C
#413250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#413260000000
0!
0*
09
0>
0C
#413270000000
1!
1*
b101 6
19
1>
1C
b101 G
#413280000000
0!
0*
09
0>
0C
#413290000000
1!
1*
b110 6
19
1>
1C
b110 G
#413300000000
0!
0*
09
0>
0C
#413310000000
1!
1*
b111 6
19
1>
1C
b111 G
#413320000000
0!
0*
09
0>
0C
#413330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#413340000000
0!
0*
09
0>
0C
#413350000000
1!
1*
b1 6
19
1>
1C
b1 G
#413360000000
0!
0*
09
0>
0C
#413370000000
1!
1*
b10 6
19
1>
1C
b10 G
#413380000000
0!
0*
09
0>
0C
#413390000000
1!
1*
b11 6
19
1>
1C
b11 G
#413400000000
0!
0*
09
0>
0C
#413410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#413420000000
0!
0*
09
0>
0C
#413430000000
1!
1*
b101 6
19
1>
1C
b101 G
#413440000000
0!
0*
09
0>
0C
#413450000000
1!
1*
b110 6
19
1>
1C
b110 G
#413460000000
0!
0*
09
0>
0C
#413470000000
1!
1*
b111 6
19
1>
1C
b111 G
#413480000000
0!
1"
0*
1+
09
1:
0>
0C
#413490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#413500000000
0!
0*
09
0>
0C
#413510000000
1!
1*
b1 6
19
1>
1C
b1 G
#413520000000
0!
0*
09
0>
0C
#413530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#413540000000
0!
0*
09
0>
0C
#413550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#413560000000
0!
0*
09
0>
0C
#413570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#413580000000
0!
0*
09
0>
0C
#413590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#413600000000
0!
0#
0*
0,
09
0>
0?
0C
#413610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#413620000000
0!
0*
09
0>
0C
#413630000000
1!
1*
19
1>
1C
#413640000000
0!
0*
09
0>
0C
#413650000000
1!
1*
19
1>
1C
#413660000000
0!
0*
09
0>
0C
#413670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#413680000000
0!
0*
09
0>
0C
#413690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#413700000000
0!
0*
09
0>
0C
#413710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#413720000000
0!
0*
09
0>
0C
#413730000000
1!
1*
b10 6
19
1>
1C
b10 G
#413740000000
0!
0*
09
0>
0C
#413750000000
1!
1*
b11 6
19
1>
1C
b11 G
#413760000000
0!
0*
09
0>
0C
#413770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#413780000000
0!
0*
09
0>
0C
#413790000000
1!
1*
b101 6
19
1>
1C
b101 G
#413800000000
0!
0*
09
0>
0C
#413810000000
1!
1*
b110 6
19
1>
1C
b110 G
#413820000000
0!
0*
09
0>
0C
#413830000000
1!
1*
b111 6
19
1>
1C
b111 G
#413840000000
0!
0*
09
0>
0C
#413850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#413860000000
0!
0*
09
0>
0C
#413870000000
1!
1*
b1 6
19
1>
1C
b1 G
#413880000000
0!
0*
09
0>
0C
#413890000000
1!
1*
b10 6
19
1>
1C
b10 G
#413900000000
0!
0*
09
0>
0C
#413910000000
1!
1*
b11 6
19
1>
1C
b11 G
#413920000000
0!
0*
09
0>
0C
#413930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#413940000000
0!
0*
09
0>
0C
#413950000000
1!
1*
b101 6
19
1>
1C
b101 G
#413960000000
0!
0*
09
0>
0C
#413970000000
1!
1*
b110 6
19
1>
1C
b110 G
#413980000000
0!
0*
09
0>
0C
#413990000000
1!
1*
b111 6
19
1>
1C
b111 G
#414000000000
0!
0*
09
0>
0C
#414010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#414020000000
0!
0*
09
0>
0C
#414030000000
1!
1*
b1 6
19
1>
1C
b1 G
#414040000000
0!
0*
09
0>
0C
#414050000000
1!
1*
b10 6
19
1>
1C
b10 G
#414060000000
0!
0*
09
0>
0C
#414070000000
1!
1*
b11 6
19
1>
1C
b11 G
#414080000000
0!
0*
09
0>
0C
#414090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#414100000000
0!
0*
09
0>
0C
#414110000000
1!
1*
b101 6
19
1>
1C
b101 G
#414120000000
0!
0*
09
0>
0C
#414130000000
1!
1*
b110 6
19
1>
1C
b110 G
#414140000000
0!
0*
09
0>
0C
#414150000000
1!
1*
b111 6
19
1>
1C
b111 G
#414160000000
0!
1"
0*
1+
09
1:
0>
0C
#414170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#414180000000
0!
0*
09
0>
0C
#414190000000
1!
1*
b1 6
19
1>
1C
b1 G
#414200000000
0!
0*
09
0>
0C
#414210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#414220000000
0!
0*
09
0>
0C
#414230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#414240000000
0!
0*
09
0>
0C
#414250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#414260000000
0!
0*
09
0>
0C
#414270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#414280000000
0!
0#
0*
0,
09
0>
0?
0C
#414290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#414300000000
0!
0*
09
0>
0C
#414310000000
1!
1*
19
1>
1C
#414320000000
0!
0*
09
0>
0C
#414330000000
1!
1*
19
1>
1C
#414340000000
0!
0*
09
0>
0C
#414350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#414360000000
0!
0*
09
0>
0C
#414370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#414380000000
0!
0*
09
0>
0C
#414390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#414400000000
0!
0*
09
0>
0C
#414410000000
1!
1*
b10 6
19
1>
1C
b10 G
#414420000000
0!
0*
09
0>
0C
#414430000000
1!
1*
b11 6
19
1>
1C
b11 G
#414440000000
0!
0*
09
0>
0C
#414450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#414460000000
0!
0*
09
0>
0C
#414470000000
1!
1*
b101 6
19
1>
1C
b101 G
#414480000000
0!
0*
09
0>
0C
#414490000000
1!
1*
b110 6
19
1>
1C
b110 G
#414500000000
0!
0*
09
0>
0C
#414510000000
1!
1*
b111 6
19
1>
1C
b111 G
#414520000000
0!
0*
09
0>
0C
#414530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#414540000000
0!
0*
09
0>
0C
#414550000000
1!
1*
b1 6
19
1>
1C
b1 G
#414560000000
0!
0*
09
0>
0C
#414570000000
1!
1*
b10 6
19
1>
1C
b10 G
#414580000000
0!
0*
09
0>
0C
#414590000000
1!
1*
b11 6
19
1>
1C
b11 G
#414600000000
0!
0*
09
0>
0C
#414610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#414620000000
0!
0*
09
0>
0C
#414630000000
1!
1*
b101 6
19
1>
1C
b101 G
#414640000000
0!
0*
09
0>
0C
#414650000000
1!
1*
b110 6
19
1>
1C
b110 G
#414660000000
0!
0*
09
0>
0C
#414670000000
1!
1*
b111 6
19
1>
1C
b111 G
#414680000000
0!
0*
09
0>
0C
#414690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#414700000000
0!
0*
09
0>
0C
#414710000000
1!
1*
b1 6
19
1>
1C
b1 G
#414720000000
0!
0*
09
0>
0C
#414730000000
1!
1*
b10 6
19
1>
1C
b10 G
#414740000000
0!
0*
09
0>
0C
#414750000000
1!
1*
b11 6
19
1>
1C
b11 G
#414760000000
0!
0*
09
0>
0C
#414770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#414780000000
0!
0*
09
0>
0C
#414790000000
1!
1*
b101 6
19
1>
1C
b101 G
#414800000000
0!
0*
09
0>
0C
#414810000000
1!
1*
b110 6
19
1>
1C
b110 G
#414820000000
0!
0*
09
0>
0C
#414830000000
1!
1*
b111 6
19
1>
1C
b111 G
#414840000000
0!
1"
0*
1+
09
1:
0>
0C
#414850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#414860000000
0!
0*
09
0>
0C
#414870000000
1!
1*
b1 6
19
1>
1C
b1 G
#414880000000
0!
0*
09
0>
0C
#414890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#414900000000
0!
0*
09
0>
0C
#414910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#414920000000
0!
0*
09
0>
0C
#414930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#414940000000
0!
0*
09
0>
0C
#414950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#414960000000
0!
0#
0*
0,
09
0>
0?
0C
#414970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#414980000000
0!
0*
09
0>
0C
#414990000000
1!
1*
19
1>
1C
#415000000000
0!
0*
09
0>
0C
#415010000000
1!
1*
19
1>
1C
#415020000000
0!
0*
09
0>
0C
#415030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#415040000000
0!
0*
09
0>
0C
#415050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#415060000000
0!
0*
09
0>
0C
#415070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#415080000000
0!
0*
09
0>
0C
#415090000000
1!
1*
b10 6
19
1>
1C
b10 G
#415100000000
0!
0*
09
0>
0C
#415110000000
1!
1*
b11 6
19
1>
1C
b11 G
#415120000000
0!
0*
09
0>
0C
#415130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#415140000000
0!
0*
09
0>
0C
#415150000000
1!
1*
b101 6
19
1>
1C
b101 G
#415160000000
0!
0*
09
0>
0C
#415170000000
1!
1*
b110 6
19
1>
1C
b110 G
#415180000000
0!
0*
09
0>
0C
#415190000000
1!
1*
b111 6
19
1>
1C
b111 G
#415200000000
0!
0*
09
0>
0C
#415210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#415220000000
0!
0*
09
0>
0C
#415230000000
1!
1*
b1 6
19
1>
1C
b1 G
#415240000000
0!
0*
09
0>
0C
#415250000000
1!
1*
b10 6
19
1>
1C
b10 G
#415260000000
0!
0*
09
0>
0C
#415270000000
1!
1*
b11 6
19
1>
1C
b11 G
#415280000000
0!
0*
09
0>
0C
#415290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#415300000000
0!
0*
09
0>
0C
#415310000000
1!
1*
b101 6
19
1>
1C
b101 G
#415320000000
0!
0*
09
0>
0C
#415330000000
1!
1*
b110 6
19
1>
1C
b110 G
#415340000000
0!
0*
09
0>
0C
#415350000000
1!
1*
b111 6
19
1>
1C
b111 G
#415360000000
0!
0*
09
0>
0C
#415370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#415380000000
0!
0*
09
0>
0C
#415390000000
1!
1*
b1 6
19
1>
1C
b1 G
#415400000000
0!
0*
09
0>
0C
#415410000000
1!
1*
b10 6
19
1>
1C
b10 G
#415420000000
0!
0*
09
0>
0C
#415430000000
1!
1*
b11 6
19
1>
1C
b11 G
#415440000000
0!
0*
09
0>
0C
#415450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#415460000000
0!
0*
09
0>
0C
#415470000000
1!
1*
b101 6
19
1>
1C
b101 G
#415480000000
0!
0*
09
0>
0C
#415490000000
1!
1*
b110 6
19
1>
1C
b110 G
#415500000000
0!
0*
09
0>
0C
#415510000000
1!
1*
b111 6
19
1>
1C
b111 G
#415520000000
0!
1"
0*
1+
09
1:
0>
0C
#415530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#415540000000
0!
0*
09
0>
0C
#415550000000
1!
1*
b1 6
19
1>
1C
b1 G
#415560000000
0!
0*
09
0>
0C
#415570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#415580000000
0!
0*
09
0>
0C
#415590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#415600000000
0!
0*
09
0>
0C
#415610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#415620000000
0!
0*
09
0>
0C
#415630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#415640000000
0!
0#
0*
0,
09
0>
0?
0C
#415650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#415660000000
0!
0*
09
0>
0C
#415670000000
1!
1*
19
1>
1C
#415680000000
0!
0*
09
0>
0C
#415690000000
1!
1*
19
1>
1C
#415700000000
0!
0*
09
0>
0C
#415710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#415720000000
0!
0*
09
0>
0C
#415730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#415740000000
0!
0*
09
0>
0C
#415750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#415760000000
0!
0*
09
0>
0C
#415770000000
1!
1*
b10 6
19
1>
1C
b10 G
#415780000000
0!
0*
09
0>
0C
#415790000000
1!
1*
b11 6
19
1>
1C
b11 G
#415800000000
0!
0*
09
0>
0C
#415810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#415820000000
0!
0*
09
0>
0C
#415830000000
1!
1*
b101 6
19
1>
1C
b101 G
#415840000000
0!
0*
09
0>
0C
#415850000000
1!
1*
b110 6
19
1>
1C
b110 G
#415860000000
0!
0*
09
0>
0C
#415870000000
1!
1*
b111 6
19
1>
1C
b111 G
#415880000000
0!
0*
09
0>
0C
#415890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#415900000000
0!
0*
09
0>
0C
#415910000000
1!
1*
b1 6
19
1>
1C
b1 G
#415920000000
0!
0*
09
0>
0C
#415930000000
1!
1*
b10 6
19
1>
1C
b10 G
#415940000000
0!
0*
09
0>
0C
#415950000000
1!
1*
b11 6
19
1>
1C
b11 G
#415960000000
0!
0*
09
0>
0C
#415970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#415980000000
0!
0*
09
0>
0C
#415990000000
1!
1*
b101 6
19
1>
1C
b101 G
#416000000000
0!
0*
09
0>
0C
#416010000000
1!
1*
b110 6
19
1>
1C
b110 G
#416020000000
0!
0*
09
0>
0C
#416030000000
1!
1*
b111 6
19
1>
1C
b111 G
#416040000000
0!
0*
09
0>
0C
#416050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#416060000000
0!
0*
09
0>
0C
#416070000000
1!
1*
b1 6
19
1>
1C
b1 G
#416080000000
0!
0*
09
0>
0C
#416090000000
1!
1*
b10 6
19
1>
1C
b10 G
#416100000000
0!
0*
09
0>
0C
#416110000000
1!
1*
b11 6
19
1>
1C
b11 G
#416120000000
0!
0*
09
0>
0C
#416130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#416140000000
0!
0*
09
0>
0C
#416150000000
1!
1*
b101 6
19
1>
1C
b101 G
#416160000000
0!
0*
09
0>
0C
#416170000000
1!
1*
b110 6
19
1>
1C
b110 G
#416180000000
0!
0*
09
0>
0C
#416190000000
1!
1*
b111 6
19
1>
1C
b111 G
#416200000000
0!
1"
0*
1+
09
1:
0>
0C
#416210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#416220000000
0!
0*
09
0>
0C
#416230000000
1!
1*
b1 6
19
1>
1C
b1 G
#416240000000
0!
0*
09
0>
0C
#416250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#416260000000
0!
0*
09
0>
0C
#416270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#416280000000
0!
0*
09
0>
0C
#416290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#416300000000
0!
0*
09
0>
0C
#416310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#416320000000
0!
0#
0*
0,
09
0>
0?
0C
#416330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#416340000000
0!
0*
09
0>
0C
#416350000000
1!
1*
19
1>
1C
#416360000000
0!
0*
09
0>
0C
#416370000000
1!
1*
19
1>
1C
#416380000000
0!
0*
09
0>
0C
#416390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#416400000000
0!
0*
09
0>
0C
#416410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#416420000000
0!
0*
09
0>
0C
#416430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#416440000000
0!
0*
09
0>
0C
#416450000000
1!
1*
b10 6
19
1>
1C
b10 G
#416460000000
0!
0*
09
0>
0C
#416470000000
1!
1*
b11 6
19
1>
1C
b11 G
#416480000000
0!
0*
09
0>
0C
#416490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#416500000000
0!
0*
09
0>
0C
#416510000000
1!
1*
b101 6
19
1>
1C
b101 G
#416520000000
0!
0*
09
0>
0C
#416530000000
1!
1*
b110 6
19
1>
1C
b110 G
#416540000000
0!
0*
09
0>
0C
#416550000000
1!
1*
b111 6
19
1>
1C
b111 G
#416560000000
0!
0*
09
0>
0C
#416570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#416580000000
0!
0*
09
0>
0C
#416590000000
1!
1*
b1 6
19
1>
1C
b1 G
#416600000000
0!
0*
09
0>
0C
#416610000000
1!
1*
b10 6
19
1>
1C
b10 G
#416620000000
0!
0*
09
0>
0C
#416630000000
1!
1*
b11 6
19
1>
1C
b11 G
#416640000000
0!
0*
09
0>
0C
#416650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#416660000000
0!
0*
09
0>
0C
#416670000000
1!
1*
b101 6
19
1>
1C
b101 G
#416680000000
0!
0*
09
0>
0C
#416690000000
1!
1*
b110 6
19
1>
1C
b110 G
#416700000000
0!
0*
09
0>
0C
#416710000000
1!
1*
b111 6
19
1>
1C
b111 G
#416720000000
0!
0*
09
0>
0C
#416730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#416740000000
0!
0*
09
0>
0C
#416750000000
1!
1*
b1 6
19
1>
1C
b1 G
#416760000000
0!
0*
09
0>
0C
#416770000000
1!
1*
b10 6
19
1>
1C
b10 G
#416780000000
0!
0*
09
0>
0C
#416790000000
1!
1*
b11 6
19
1>
1C
b11 G
#416800000000
0!
0*
09
0>
0C
#416810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#416820000000
0!
0*
09
0>
0C
#416830000000
1!
1*
b101 6
19
1>
1C
b101 G
#416840000000
0!
0*
09
0>
0C
#416850000000
1!
1*
b110 6
19
1>
1C
b110 G
#416860000000
0!
0*
09
0>
0C
#416870000000
1!
1*
b111 6
19
1>
1C
b111 G
#416880000000
0!
1"
0*
1+
09
1:
0>
0C
#416890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#416900000000
0!
0*
09
0>
0C
#416910000000
1!
1*
b1 6
19
1>
1C
b1 G
#416920000000
0!
0*
09
0>
0C
#416930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#416940000000
0!
0*
09
0>
0C
#416950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#416960000000
0!
0*
09
0>
0C
#416970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#416980000000
0!
0*
09
0>
0C
#416990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#417000000000
0!
0#
0*
0,
09
0>
0?
0C
#417010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#417020000000
0!
0*
09
0>
0C
#417030000000
1!
1*
19
1>
1C
#417040000000
0!
0*
09
0>
0C
#417050000000
1!
1*
19
1>
1C
#417060000000
0!
0*
09
0>
0C
#417070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#417080000000
0!
0*
09
0>
0C
#417090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#417100000000
0!
0*
09
0>
0C
#417110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#417120000000
0!
0*
09
0>
0C
#417130000000
1!
1*
b10 6
19
1>
1C
b10 G
#417140000000
0!
0*
09
0>
0C
#417150000000
1!
1*
b11 6
19
1>
1C
b11 G
#417160000000
0!
0*
09
0>
0C
#417170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#417180000000
0!
0*
09
0>
0C
#417190000000
1!
1*
b101 6
19
1>
1C
b101 G
#417200000000
0!
0*
09
0>
0C
#417210000000
1!
1*
b110 6
19
1>
1C
b110 G
#417220000000
0!
0*
09
0>
0C
#417230000000
1!
1*
b111 6
19
1>
1C
b111 G
#417240000000
0!
0*
09
0>
0C
#417250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#417260000000
0!
0*
09
0>
0C
#417270000000
1!
1*
b1 6
19
1>
1C
b1 G
#417280000000
0!
0*
09
0>
0C
#417290000000
1!
1*
b10 6
19
1>
1C
b10 G
#417300000000
0!
0*
09
0>
0C
#417310000000
1!
1*
b11 6
19
1>
1C
b11 G
#417320000000
0!
0*
09
0>
0C
#417330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#417340000000
0!
0*
09
0>
0C
#417350000000
1!
1*
b101 6
19
1>
1C
b101 G
#417360000000
0!
0*
09
0>
0C
#417370000000
1!
1*
b110 6
19
1>
1C
b110 G
#417380000000
0!
0*
09
0>
0C
#417390000000
1!
1*
b111 6
19
1>
1C
b111 G
#417400000000
0!
0*
09
0>
0C
#417410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#417420000000
0!
0*
09
0>
0C
#417430000000
1!
1*
b1 6
19
1>
1C
b1 G
#417440000000
0!
0*
09
0>
0C
#417450000000
1!
1*
b10 6
19
1>
1C
b10 G
#417460000000
0!
0*
09
0>
0C
#417470000000
1!
1*
b11 6
19
1>
1C
b11 G
#417480000000
0!
0*
09
0>
0C
#417490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#417500000000
0!
0*
09
0>
0C
#417510000000
1!
1*
b101 6
19
1>
1C
b101 G
#417520000000
0!
0*
09
0>
0C
#417530000000
1!
1*
b110 6
19
1>
1C
b110 G
#417540000000
0!
0*
09
0>
0C
#417550000000
1!
1*
b111 6
19
1>
1C
b111 G
#417560000000
0!
1"
0*
1+
09
1:
0>
0C
#417570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#417580000000
0!
0*
09
0>
0C
#417590000000
1!
1*
b1 6
19
1>
1C
b1 G
#417600000000
0!
0*
09
0>
0C
#417610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#417620000000
0!
0*
09
0>
0C
#417630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#417640000000
0!
0*
09
0>
0C
#417650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#417660000000
0!
0*
09
0>
0C
#417670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#417680000000
0!
0#
0*
0,
09
0>
0?
0C
#417690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#417700000000
0!
0*
09
0>
0C
#417710000000
1!
1*
19
1>
1C
#417720000000
0!
0*
09
0>
0C
#417730000000
1!
1*
19
1>
1C
#417740000000
0!
0*
09
0>
0C
#417750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#417760000000
0!
0*
09
0>
0C
#417770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#417780000000
0!
0*
09
0>
0C
#417790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#417800000000
0!
0*
09
0>
0C
#417810000000
1!
1*
b10 6
19
1>
1C
b10 G
#417820000000
0!
0*
09
0>
0C
#417830000000
1!
1*
b11 6
19
1>
1C
b11 G
#417840000000
0!
0*
09
0>
0C
#417850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#417860000000
0!
0*
09
0>
0C
#417870000000
1!
1*
b101 6
19
1>
1C
b101 G
#417880000000
0!
0*
09
0>
0C
#417890000000
1!
1*
b110 6
19
1>
1C
b110 G
#417900000000
0!
0*
09
0>
0C
#417910000000
1!
1*
b111 6
19
1>
1C
b111 G
#417920000000
0!
0*
09
0>
0C
#417930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#417940000000
0!
0*
09
0>
0C
#417950000000
1!
1*
b1 6
19
1>
1C
b1 G
#417960000000
0!
0*
09
0>
0C
#417970000000
1!
1*
b10 6
19
1>
1C
b10 G
#417980000000
0!
0*
09
0>
0C
#417990000000
1!
1*
b11 6
19
1>
1C
b11 G
#418000000000
0!
0*
09
0>
0C
#418010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#418020000000
0!
0*
09
0>
0C
#418030000000
1!
1*
b101 6
19
1>
1C
b101 G
#418040000000
0!
0*
09
0>
0C
#418050000000
1!
1*
b110 6
19
1>
1C
b110 G
#418060000000
0!
0*
09
0>
0C
#418070000000
1!
1*
b111 6
19
1>
1C
b111 G
#418080000000
0!
0*
09
0>
0C
#418090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#418100000000
0!
0*
09
0>
0C
#418110000000
1!
1*
b1 6
19
1>
1C
b1 G
#418120000000
0!
0*
09
0>
0C
#418130000000
1!
1*
b10 6
19
1>
1C
b10 G
#418140000000
0!
0*
09
0>
0C
#418150000000
1!
1*
b11 6
19
1>
1C
b11 G
#418160000000
0!
0*
09
0>
0C
#418170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#418180000000
0!
0*
09
0>
0C
#418190000000
1!
1*
b101 6
19
1>
1C
b101 G
#418200000000
0!
0*
09
0>
0C
#418210000000
1!
1*
b110 6
19
1>
1C
b110 G
#418220000000
0!
0*
09
0>
0C
#418230000000
1!
1*
b111 6
19
1>
1C
b111 G
#418240000000
0!
1"
0*
1+
09
1:
0>
0C
#418250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#418260000000
0!
0*
09
0>
0C
#418270000000
1!
1*
b1 6
19
1>
1C
b1 G
#418280000000
0!
0*
09
0>
0C
#418290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#418300000000
0!
0*
09
0>
0C
#418310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#418320000000
0!
0*
09
0>
0C
#418330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#418340000000
0!
0*
09
0>
0C
#418350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#418360000000
0!
0#
0*
0,
09
0>
0?
0C
#418370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#418380000000
0!
0*
09
0>
0C
#418390000000
1!
1*
19
1>
1C
#418400000000
0!
0*
09
0>
0C
#418410000000
1!
1*
19
1>
1C
#418420000000
0!
0*
09
0>
0C
#418430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#418440000000
0!
0*
09
0>
0C
#418450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#418460000000
0!
0*
09
0>
0C
#418470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#418480000000
0!
0*
09
0>
0C
#418490000000
1!
1*
b10 6
19
1>
1C
b10 G
#418500000000
0!
0*
09
0>
0C
#418510000000
1!
1*
b11 6
19
1>
1C
b11 G
#418520000000
0!
0*
09
0>
0C
#418530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#418540000000
0!
0*
09
0>
0C
#418550000000
1!
1*
b101 6
19
1>
1C
b101 G
#418560000000
0!
0*
09
0>
0C
#418570000000
1!
1*
b110 6
19
1>
1C
b110 G
#418580000000
0!
0*
09
0>
0C
#418590000000
1!
1*
b111 6
19
1>
1C
b111 G
#418600000000
0!
0*
09
0>
0C
#418610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#418620000000
0!
0*
09
0>
0C
#418630000000
1!
1*
b1 6
19
1>
1C
b1 G
#418640000000
0!
0*
09
0>
0C
#418650000000
1!
1*
b10 6
19
1>
1C
b10 G
#418660000000
0!
0*
09
0>
0C
#418670000000
1!
1*
b11 6
19
1>
1C
b11 G
#418680000000
0!
0*
09
0>
0C
#418690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#418700000000
0!
0*
09
0>
0C
#418710000000
1!
1*
b101 6
19
1>
1C
b101 G
#418720000000
0!
0*
09
0>
0C
#418730000000
1!
1*
b110 6
19
1>
1C
b110 G
#418740000000
0!
0*
09
0>
0C
#418750000000
1!
1*
b111 6
19
1>
1C
b111 G
#418760000000
0!
0*
09
0>
0C
#418770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#418780000000
0!
0*
09
0>
0C
#418790000000
1!
1*
b1 6
19
1>
1C
b1 G
#418800000000
0!
0*
09
0>
0C
#418810000000
1!
1*
b10 6
19
1>
1C
b10 G
#418820000000
0!
0*
09
0>
0C
#418830000000
1!
1*
b11 6
19
1>
1C
b11 G
#418840000000
0!
0*
09
0>
0C
#418850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#418860000000
0!
0*
09
0>
0C
#418870000000
1!
1*
b101 6
19
1>
1C
b101 G
#418880000000
0!
0*
09
0>
0C
#418890000000
1!
1*
b110 6
19
1>
1C
b110 G
#418900000000
0!
0*
09
0>
0C
#418910000000
1!
1*
b111 6
19
1>
1C
b111 G
#418920000000
0!
1"
0*
1+
09
1:
0>
0C
#418930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#418940000000
0!
0*
09
0>
0C
#418950000000
1!
1*
b1 6
19
1>
1C
b1 G
#418960000000
0!
0*
09
0>
0C
#418970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#418980000000
0!
0*
09
0>
0C
#418990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#419000000000
0!
0*
09
0>
0C
#419010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#419020000000
0!
0*
09
0>
0C
#419030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#419040000000
0!
0#
0*
0,
09
0>
0?
0C
#419050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#419060000000
0!
0*
09
0>
0C
#419070000000
1!
1*
19
1>
1C
#419080000000
0!
0*
09
0>
0C
#419090000000
1!
1*
19
1>
1C
#419100000000
0!
0*
09
0>
0C
#419110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#419120000000
0!
0*
09
0>
0C
#419130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#419140000000
0!
0*
09
0>
0C
#419150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#419160000000
0!
0*
09
0>
0C
#419170000000
1!
1*
b10 6
19
1>
1C
b10 G
#419180000000
0!
0*
09
0>
0C
#419190000000
1!
1*
b11 6
19
1>
1C
b11 G
#419200000000
0!
0*
09
0>
0C
#419210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#419220000000
0!
0*
09
0>
0C
#419230000000
1!
1*
b101 6
19
1>
1C
b101 G
#419240000000
0!
0*
09
0>
0C
#419250000000
1!
1*
b110 6
19
1>
1C
b110 G
#419260000000
0!
0*
09
0>
0C
#419270000000
1!
1*
b111 6
19
1>
1C
b111 G
#419280000000
0!
0*
09
0>
0C
#419290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#419300000000
0!
0*
09
0>
0C
#419310000000
1!
1*
b1 6
19
1>
1C
b1 G
#419320000000
0!
0*
09
0>
0C
#419330000000
1!
1*
b10 6
19
1>
1C
b10 G
#419340000000
0!
0*
09
0>
0C
#419350000000
1!
1*
b11 6
19
1>
1C
b11 G
#419360000000
0!
0*
09
0>
0C
#419370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#419380000000
0!
0*
09
0>
0C
#419390000000
1!
1*
b101 6
19
1>
1C
b101 G
#419400000000
0!
0*
09
0>
0C
#419410000000
1!
1*
b110 6
19
1>
1C
b110 G
#419420000000
0!
0*
09
0>
0C
#419430000000
1!
1*
b111 6
19
1>
1C
b111 G
#419440000000
0!
0*
09
0>
0C
#419450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#419460000000
0!
0*
09
0>
0C
#419470000000
1!
1*
b1 6
19
1>
1C
b1 G
#419480000000
0!
0*
09
0>
0C
#419490000000
1!
1*
b10 6
19
1>
1C
b10 G
#419500000000
0!
0*
09
0>
0C
#419510000000
1!
1*
b11 6
19
1>
1C
b11 G
#419520000000
0!
0*
09
0>
0C
#419530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#419540000000
0!
0*
09
0>
0C
#419550000000
1!
1*
b101 6
19
1>
1C
b101 G
#419560000000
0!
0*
09
0>
0C
#419570000000
1!
1*
b110 6
19
1>
1C
b110 G
#419580000000
0!
0*
09
0>
0C
#419590000000
1!
1*
b111 6
19
1>
1C
b111 G
#419600000000
0!
1"
0*
1+
09
1:
0>
0C
#419610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#419620000000
0!
0*
09
0>
0C
#419630000000
1!
1*
b1 6
19
1>
1C
b1 G
#419640000000
0!
0*
09
0>
0C
#419650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#419660000000
0!
0*
09
0>
0C
#419670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#419680000000
0!
0*
09
0>
0C
#419690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#419700000000
0!
0*
09
0>
0C
#419710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#419720000000
0!
0#
0*
0,
09
0>
0?
0C
#419730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#419740000000
0!
0*
09
0>
0C
#419750000000
1!
1*
19
1>
1C
#419760000000
0!
0*
09
0>
0C
#419770000000
1!
1*
19
1>
1C
#419780000000
0!
0*
09
0>
0C
#419790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#419800000000
0!
0*
09
0>
0C
#419810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#419820000000
0!
0*
09
0>
0C
#419830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#419840000000
0!
0*
09
0>
0C
#419850000000
1!
1*
b10 6
19
1>
1C
b10 G
#419860000000
0!
0*
09
0>
0C
#419870000000
1!
1*
b11 6
19
1>
1C
b11 G
#419880000000
0!
0*
09
0>
0C
#419890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#419900000000
0!
0*
09
0>
0C
#419910000000
1!
1*
b101 6
19
1>
1C
b101 G
#419920000000
0!
0*
09
0>
0C
#419930000000
1!
1*
b110 6
19
1>
1C
b110 G
#419940000000
0!
0*
09
0>
0C
#419950000000
1!
1*
b111 6
19
1>
1C
b111 G
#419960000000
0!
0*
09
0>
0C
#419970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#419980000000
0!
0*
09
0>
0C
#419990000000
1!
1*
b1 6
19
1>
1C
b1 G
#420000000000
0!
0*
09
0>
0C
#420010000000
1!
1*
b10 6
19
1>
1C
b10 G
#420020000000
0!
0*
09
0>
0C
#420030000000
1!
1*
b11 6
19
1>
1C
b11 G
#420040000000
0!
0*
09
0>
0C
#420050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#420060000000
0!
0*
09
0>
0C
#420070000000
1!
1*
b101 6
19
1>
1C
b101 G
#420080000000
0!
0*
09
0>
0C
#420090000000
1!
1*
b110 6
19
1>
1C
b110 G
#420100000000
0!
0*
09
0>
0C
#420110000000
1!
1*
b111 6
19
1>
1C
b111 G
#420120000000
0!
0*
09
0>
0C
#420130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#420140000000
0!
0*
09
0>
0C
#420150000000
1!
1*
b1 6
19
1>
1C
b1 G
#420160000000
0!
0*
09
0>
0C
#420170000000
1!
1*
b10 6
19
1>
1C
b10 G
#420180000000
0!
0*
09
0>
0C
#420190000000
1!
1*
b11 6
19
1>
1C
b11 G
#420200000000
0!
0*
09
0>
0C
#420210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#420220000000
0!
0*
09
0>
0C
#420230000000
1!
1*
b101 6
19
1>
1C
b101 G
#420240000000
0!
0*
09
0>
0C
#420250000000
1!
1*
b110 6
19
1>
1C
b110 G
#420260000000
0!
0*
09
0>
0C
#420270000000
1!
1*
b111 6
19
1>
1C
b111 G
#420280000000
0!
1"
0*
1+
09
1:
0>
0C
#420290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#420300000000
0!
0*
09
0>
0C
#420310000000
1!
1*
b1 6
19
1>
1C
b1 G
#420320000000
0!
0*
09
0>
0C
#420330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#420340000000
0!
0*
09
0>
0C
#420350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#420360000000
0!
0*
09
0>
0C
#420370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#420380000000
0!
0*
09
0>
0C
#420390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#420400000000
0!
0#
0*
0,
09
0>
0?
0C
#420410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#420420000000
0!
0*
09
0>
0C
#420430000000
1!
1*
19
1>
1C
#420440000000
0!
0*
09
0>
0C
#420450000000
1!
1*
19
1>
1C
#420460000000
0!
0*
09
0>
0C
#420470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#420480000000
0!
0*
09
0>
0C
#420490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#420500000000
0!
0*
09
0>
0C
#420510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#420520000000
0!
0*
09
0>
0C
#420530000000
1!
1*
b10 6
19
1>
1C
b10 G
#420540000000
0!
0*
09
0>
0C
#420550000000
1!
1*
b11 6
19
1>
1C
b11 G
#420560000000
0!
0*
09
0>
0C
#420570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#420580000000
0!
0*
09
0>
0C
#420590000000
1!
1*
b101 6
19
1>
1C
b101 G
#420600000000
0!
0*
09
0>
0C
#420610000000
1!
1*
b110 6
19
1>
1C
b110 G
#420620000000
0!
0*
09
0>
0C
#420630000000
1!
1*
b111 6
19
1>
1C
b111 G
#420640000000
0!
0*
09
0>
0C
#420650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#420660000000
0!
0*
09
0>
0C
#420670000000
1!
1*
b1 6
19
1>
1C
b1 G
#420680000000
0!
0*
09
0>
0C
#420690000000
1!
1*
b10 6
19
1>
1C
b10 G
#420700000000
0!
0*
09
0>
0C
#420710000000
1!
1*
b11 6
19
1>
1C
b11 G
#420720000000
0!
0*
09
0>
0C
#420730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#420740000000
0!
0*
09
0>
0C
#420750000000
1!
1*
b101 6
19
1>
1C
b101 G
#420760000000
0!
0*
09
0>
0C
#420770000000
1!
1*
b110 6
19
1>
1C
b110 G
#420780000000
0!
0*
09
0>
0C
#420790000000
1!
1*
b111 6
19
1>
1C
b111 G
#420800000000
0!
0*
09
0>
0C
#420810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#420820000000
0!
0*
09
0>
0C
#420830000000
1!
1*
b1 6
19
1>
1C
b1 G
#420840000000
0!
0*
09
0>
0C
#420850000000
1!
1*
b10 6
19
1>
1C
b10 G
#420860000000
0!
0*
09
0>
0C
#420870000000
1!
1*
b11 6
19
1>
1C
b11 G
#420880000000
0!
0*
09
0>
0C
#420890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#420900000000
0!
0*
09
0>
0C
#420910000000
1!
1*
b101 6
19
1>
1C
b101 G
#420920000000
0!
0*
09
0>
0C
#420930000000
1!
1*
b110 6
19
1>
1C
b110 G
#420940000000
0!
0*
09
0>
0C
#420950000000
1!
1*
b111 6
19
1>
1C
b111 G
#420960000000
0!
1"
0*
1+
09
1:
0>
0C
#420970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#420980000000
0!
0*
09
0>
0C
#420990000000
1!
1*
b1 6
19
1>
1C
b1 G
#421000000000
0!
0*
09
0>
0C
#421010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#421020000000
0!
0*
09
0>
0C
#421030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#421040000000
0!
0*
09
0>
0C
#421050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#421060000000
0!
0*
09
0>
0C
#421070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#421080000000
0!
0#
0*
0,
09
0>
0?
0C
#421090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#421100000000
0!
0*
09
0>
0C
#421110000000
1!
1*
19
1>
1C
#421120000000
0!
0*
09
0>
0C
#421130000000
1!
1*
19
1>
1C
#421140000000
0!
0*
09
0>
0C
#421150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#421160000000
0!
0*
09
0>
0C
#421170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#421180000000
0!
0*
09
0>
0C
#421190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#421200000000
0!
0*
09
0>
0C
#421210000000
1!
1*
b10 6
19
1>
1C
b10 G
#421220000000
0!
0*
09
0>
0C
#421230000000
1!
1*
b11 6
19
1>
1C
b11 G
#421240000000
0!
0*
09
0>
0C
#421250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#421260000000
0!
0*
09
0>
0C
#421270000000
1!
1*
b101 6
19
1>
1C
b101 G
#421280000000
0!
0*
09
0>
0C
#421290000000
1!
1*
b110 6
19
1>
1C
b110 G
#421300000000
0!
0*
09
0>
0C
#421310000000
1!
1*
b111 6
19
1>
1C
b111 G
#421320000000
0!
0*
09
0>
0C
#421330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#421340000000
0!
0*
09
0>
0C
#421350000000
1!
1*
b1 6
19
1>
1C
b1 G
#421360000000
0!
0*
09
0>
0C
#421370000000
1!
1*
b10 6
19
1>
1C
b10 G
#421380000000
0!
0*
09
0>
0C
#421390000000
1!
1*
b11 6
19
1>
1C
b11 G
#421400000000
0!
0*
09
0>
0C
#421410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#421420000000
0!
0*
09
0>
0C
#421430000000
1!
1*
b101 6
19
1>
1C
b101 G
#421440000000
0!
0*
09
0>
0C
#421450000000
1!
1*
b110 6
19
1>
1C
b110 G
#421460000000
0!
0*
09
0>
0C
#421470000000
1!
1*
b111 6
19
1>
1C
b111 G
#421480000000
0!
0*
09
0>
0C
#421490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#421500000000
0!
0*
09
0>
0C
#421510000000
1!
1*
b1 6
19
1>
1C
b1 G
#421520000000
0!
0*
09
0>
0C
#421530000000
1!
1*
b10 6
19
1>
1C
b10 G
#421540000000
0!
0*
09
0>
0C
#421550000000
1!
1*
b11 6
19
1>
1C
b11 G
#421560000000
0!
0*
09
0>
0C
#421570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#421580000000
0!
0*
09
0>
0C
#421590000000
1!
1*
b101 6
19
1>
1C
b101 G
#421600000000
0!
0*
09
0>
0C
#421610000000
1!
1*
b110 6
19
1>
1C
b110 G
#421620000000
0!
0*
09
0>
0C
#421630000000
1!
1*
b111 6
19
1>
1C
b111 G
#421640000000
0!
1"
0*
1+
09
1:
0>
0C
#421650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#421660000000
0!
0*
09
0>
0C
#421670000000
1!
1*
b1 6
19
1>
1C
b1 G
#421680000000
0!
0*
09
0>
0C
#421690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#421700000000
0!
0*
09
0>
0C
#421710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#421720000000
0!
0*
09
0>
0C
#421730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#421740000000
0!
0*
09
0>
0C
#421750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#421760000000
0!
0#
0*
0,
09
0>
0?
0C
#421770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#421780000000
0!
0*
09
0>
0C
#421790000000
1!
1*
19
1>
1C
#421800000000
0!
0*
09
0>
0C
#421810000000
1!
1*
19
1>
1C
#421820000000
0!
0*
09
0>
0C
#421830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#421840000000
0!
0*
09
0>
0C
#421850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#421860000000
0!
0*
09
0>
0C
#421870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#421880000000
0!
0*
09
0>
0C
#421890000000
1!
1*
b10 6
19
1>
1C
b10 G
#421900000000
0!
0*
09
0>
0C
#421910000000
1!
1*
b11 6
19
1>
1C
b11 G
#421920000000
0!
0*
09
0>
0C
#421930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#421940000000
0!
0*
09
0>
0C
#421950000000
1!
1*
b101 6
19
1>
1C
b101 G
#421960000000
0!
0*
09
0>
0C
#421970000000
1!
1*
b110 6
19
1>
1C
b110 G
#421980000000
0!
0*
09
0>
0C
#421990000000
1!
1*
b111 6
19
1>
1C
b111 G
#422000000000
0!
0*
09
0>
0C
#422010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#422020000000
0!
0*
09
0>
0C
#422030000000
1!
1*
b1 6
19
1>
1C
b1 G
#422040000000
0!
0*
09
0>
0C
#422050000000
1!
1*
b10 6
19
1>
1C
b10 G
#422060000000
0!
0*
09
0>
0C
#422070000000
1!
1*
b11 6
19
1>
1C
b11 G
#422080000000
0!
0*
09
0>
0C
#422090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#422100000000
0!
0*
09
0>
0C
#422110000000
1!
1*
b101 6
19
1>
1C
b101 G
#422120000000
0!
0*
09
0>
0C
#422130000000
1!
1*
b110 6
19
1>
1C
b110 G
#422140000000
0!
0*
09
0>
0C
#422150000000
1!
1*
b111 6
19
1>
1C
b111 G
#422160000000
0!
0*
09
0>
0C
#422170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#422180000000
0!
0*
09
0>
0C
#422190000000
1!
1*
b1 6
19
1>
1C
b1 G
#422200000000
0!
0*
09
0>
0C
#422210000000
1!
1*
b10 6
19
1>
1C
b10 G
#422220000000
0!
0*
09
0>
0C
#422230000000
1!
1*
b11 6
19
1>
1C
b11 G
#422240000000
0!
0*
09
0>
0C
#422250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#422260000000
0!
0*
09
0>
0C
#422270000000
1!
1*
b101 6
19
1>
1C
b101 G
#422280000000
0!
0*
09
0>
0C
#422290000000
1!
1*
b110 6
19
1>
1C
b110 G
#422300000000
0!
0*
09
0>
0C
#422310000000
1!
1*
b111 6
19
1>
1C
b111 G
#422320000000
0!
1"
0*
1+
09
1:
0>
0C
#422330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#422340000000
0!
0*
09
0>
0C
#422350000000
1!
1*
b1 6
19
1>
1C
b1 G
#422360000000
0!
0*
09
0>
0C
#422370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#422380000000
0!
0*
09
0>
0C
#422390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#422400000000
0!
0*
09
0>
0C
#422410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#422420000000
0!
0*
09
0>
0C
#422430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#422440000000
0!
0#
0*
0,
09
0>
0?
0C
#422450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#422460000000
0!
0*
09
0>
0C
#422470000000
1!
1*
19
1>
1C
#422480000000
0!
0*
09
0>
0C
#422490000000
1!
1*
19
1>
1C
#422500000000
0!
0*
09
0>
0C
#422510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#422520000000
0!
0*
09
0>
0C
#422530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#422540000000
0!
0*
09
0>
0C
#422550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#422560000000
0!
0*
09
0>
0C
#422570000000
1!
1*
b10 6
19
1>
1C
b10 G
#422580000000
0!
0*
09
0>
0C
#422590000000
1!
1*
b11 6
19
1>
1C
b11 G
#422600000000
0!
0*
09
0>
0C
#422610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#422620000000
0!
0*
09
0>
0C
#422630000000
1!
1*
b101 6
19
1>
1C
b101 G
#422640000000
0!
0*
09
0>
0C
#422650000000
1!
1*
b110 6
19
1>
1C
b110 G
#422660000000
0!
0*
09
0>
0C
#422670000000
1!
1*
b111 6
19
1>
1C
b111 G
#422680000000
0!
0*
09
0>
0C
#422690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#422700000000
0!
0*
09
0>
0C
#422710000000
1!
1*
b1 6
19
1>
1C
b1 G
#422720000000
0!
0*
09
0>
0C
#422730000000
1!
1*
b10 6
19
1>
1C
b10 G
#422740000000
0!
0*
09
0>
0C
#422750000000
1!
1*
b11 6
19
1>
1C
b11 G
#422760000000
0!
0*
09
0>
0C
#422770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#422780000000
0!
0*
09
0>
0C
#422790000000
1!
1*
b101 6
19
1>
1C
b101 G
#422800000000
0!
0*
09
0>
0C
#422810000000
1!
1*
b110 6
19
1>
1C
b110 G
#422820000000
0!
0*
09
0>
0C
#422830000000
1!
1*
b111 6
19
1>
1C
b111 G
#422840000000
0!
0*
09
0>
0C
#422850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#422860000000
0!
0*
09
0>
0C
#422870000000
1!
1*
b1 6
19
1>
1C
b1 G
#422880000000
0!
0*
09
0>
0C
#422890000000
1!
1*
b10 6
19
1>
1C
b10 G
#422900000000
0!
0*
09
0>
0C
#422910000000
1!
1*
b11 6
19
1>
1C
b11 G
#422920000000
0!
0*
09
0>
0C
#422930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#422940000000
0!
0*
09
0>
0C
#422950000000
1!
1*
b101 6
19
1>
1C
b101 G
#422960000000
0!
0*
09
0>
0C
#422970000000
1!
1*
b110 6
19
1>
1C
b110 G
#422980000000
0!
0*
09
0>
0C
#422990000000
1!
1*
b111 6
19
1>
1C
b111 G
#423000000000
0!
1"
0*
1+
09
1:
0>
0C
#423010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#423020000000
0!
0*
09
0>
0C
#423030000000
1!
1*
b1 6
19
1>
1C
b1 G
#423040000000
0!
0*
09
0>
0C
#423050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#423060000000
0!
0*
09
0>
0C
#423070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#423080000000
0!
0*
09
0>
0C
#423090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#423100000000
0!
0*
09
0>
0C
#423110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#423120000000
0!
0#
0*
0,
09
0>
0?
0C
#423130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#423140000000
0!
0*
09
0>
0C
#423150000000
1!
1*
19
1>
1C
#423160000000
0!
0*
09
0>
0C
#423170000000
1!
1*
19
1>
1C
#423180000000
0!
0*
09
0>
0C
#423190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#423200000000
0!
0*
09
0>
0C
#423210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#423220000000
0!
0*
09
0>
0C
#423230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#423240000000
0!
0*
09
0>
0C
#423250000000
1!
1*
b10 6
19
1>
1C
b10 G
#423260000000
0!
0*
09
0>
0C
#423270000000
1!
1*
b11 6
19
1>
1C
b11 G
#423280000000
0!
0*
09
0>
0C
#423290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#423300000000
0!
0*
09
0>
0C
#423310000000
1!
1*
b101 6
19
1>
1C
b101 G
#423320000000
0!
0*
09
0>
0C
#423330000000
1!
1*
b110 6
19
1>
1C
b110 G
#423340000000
0!
0*
09
0>
0C
#423350000000
1!
1*
b111 6
19
1>
1C
b111 G
#423360000000
0!
0*
09
0>
0C
#423370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#423380000000
0!
0*
09
0>
0C
#423390000000
1!
1*
b1 6
19
1>
1C
b1 G
#423400000000
0!
0*
09
0>
0C
#423410000000
1!
1*
b10 6
19
1>
1C
b10 G
#423420000000
0!
0*
09
0>
0C
#423430000000
1!
1*
b11 6
19
1>
1C
b11 G
#423440000000
0!
0*
09
0>
0C
#423450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#423460000000
0!
0*
09
0>
0C
#423470000000
1!
1*
b101 6
19
1>
1C
b101 G
#423480000000
0!
0*
09
0>
0C
#423490000000
1!
1*
b110 6
19
1>
1C
b110 G
#423500000000
0!
0*
09
0>
0C
#423510000000
1!
1*
b111 6
19
1>
1C
b111 G
#423520000000
0!
0*
09
0>
0C
#423530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#423540000000
0!
0*
09
0>
0C
#423550000000
1!
1*
b1 6
19
1>
1C
b1 G
#423560000000
0!
0*
09
0>
0C
#423570000000
1!
1*
b10 6
19
1>
1C
b10 G
#423580000000
0!
0*
09
0>
0C
#423590000000
1!
1*
b11 6
19
1>
1C
b11 G
#423600000000
0!
0*
09
0>
0C
#423610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#423620000000
0!
0*
09
0>
0C
#423630000000
1!
1*
b101 6
19
1>
1C
b101 G
#423640000000
0!
0*
09
0>
0C
#423650000000
1!
1*
b110 6
19
1>
1C
b110 G
#423660000000
0!
0*
09
0>
0C
#423670000000
1!
1*
b111 6
19
1>
1C
b111 G
#423680000000
0!
1"
0*
1+
09
1:
0>
0C
#423690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#423700000000
0!
0*
09
0>
0C
#423710000000
1!
1*
b1 6
19
1>
1C
b1 G
#423720000000
0!
0*
09
0>
0C
#423730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#423740000000
0!
0*
09
0>
0C
#423750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#423760000000
0!
0*
09
0>
0C
#423770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#423780000000
0!
0*
09
0>
0C
#423790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#423800000000
0!
0#
0*
0,
09
0>
0?
0C
#423810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#423820000000
0!
0*
09
0>
0C
#423830000000
1!
1*
19
1>
1C
#423840000000
0!
0*
09
0>
0C
#423850000000
1!
1*
19
1>
1C
#423860000000
0!
0*
09
0>
0C
#423870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#423880000000
0!
0*
09
0>
0C
#423890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#423900000000
0!
0*
09
0>
0C
#423910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#423920000000
0!
0*
09
0>
0C
#423930000000
1!
1*
b10 6
19
1>
1C
b10 G
#423940000000
0!
0*
09
0>
0C
#423950000000
1!
1*
b11 6
19
1>
1C
b11 G
#423960000000
0!
0*
09
0>
0C
#423970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#423980000000
0!
0*
09
0>
0C
#423990000000
1!
1*
b101 6
19
1>
1C
b101 G
#424000000000
0!
0*
09
0>
0C
#424010000000
1!
1*
b110 6
19
1>
1C
b110 G
#424020000000
0!
0*
09
0>
0C
#424030000000
1!
1*
b111 6
19
1>
1C
b111 G
#424040000000
0!
0*
09
0>
0C
#424050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#424060000000
0!
0*
09
0>
0C
#424070000000
1!
1*
b1 6
19
1>
1C
b1 G
#424080000000
0!
0*
09
0>
0C
#424090000000
1!
1*
b10 6
19
1>
1C
b10 G
#424100000000
0!
0*
09
0>
0C
#424110000000
1!
1*
b11 6
19
1>
1C
b11 G
#424120000000
0!
0*
09
0>
0C
#424130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#424140000000
0!
0*
09
0>
0C
#424150000000
1!
1*
b101 6
19
1>
1C
b101 G
#424160000000
0!
0*
09
0>
0C
#424170000000
1!
1*
b110 6
19
1>
1C
b110 G
#424180000000
0!
0*
09
0>
0C
#424190000000
1!
1*
b111 6
19
1>
1C
b111 G
#424200000000
0!
0*
09
0>
0C
#424210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#424220000000
0!
0*
09
0>
0C
#424230000000
1!
1*
b1 6
19
1>
1C
b1 G
#424240000000
0!
0*
09
0>
0C
#424250000000
1!
1*
b10 6
19
1>
1C
b10 G
#424260000000
0!
0*
09
0>
0C
#424270000000
1!
1*
b11 6
19
1>
1C
b11 G
#424280000000
0!
0*
09
0>
0C
#424290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#424300000000
0!
0*
09
0>
0C
#424310000000
1!
1*
b101 6
19
1>
1C
b101 G
#424320000000
0!
0*
09
0>
0C
#424330000000
1!
1*
b110 6
19
1>
1C
b110 G
#424340000000
0!
0*
09
0>
0C
#424350000000
1!
1*
b111 6
19
1>
1C
b111 G
#424360000000
0!
1"
0*
1+
09
1:
0>
0C
#424370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#424380000000
0!
0*
09
0>
0C
#424390000000
1!
1*
b1 6
19
1>
1C
b1 G
#424400000000
0!
0*
09
0>
0C
#424410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#424420000000
0!
0*
09
0>
0C
#424430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#424440000000
0!
0*
09
0>
0C
#424450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#424460000000
0!
0*
09
0>
0C
#424470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#424480000000
0!
0#
0*
0,
09
0>
0?
0C
#424490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#424500000000
0!
0*
09
0>
0C
#424510000000
1!
1*
19
1>
1C
#424520000000
0!
0*
09
0>
0C
#424530000000
1!
1*
19
1>
1C
#424540000000
0!
0*
09
0>
0C
#424550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#424560000000
0!
0*
09
0>
0C
#424570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#424580000000
0!
0*
09
0>
0C
#424590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#424600000000
0!
0*
09
0>
0C
#424610000000
1!
1*
b10 6
19
1>
1C
b10 G
#424620000000
0!
0*
09
0>
0C
#424630000000
1!
1*
b11 6
19
1>
1C
b11 G
#424640000000
0!
0*
09
0>
0C
#424650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#424660000000
0!
0*
09
0>
0C
#424670000000
1!
1*
b101 6
19
1>
1C
b101 G
#424680000000
0!
0*
09
0>
0C
#424690000000
1!
1*
b110 6
19
1>
1C
b110 G
#424700000000
0!
0*
09
0>
0C
#424710000000
1!
1*
b111 6
19
1>
1C
b111 G
#424720000000
0!
0*
09
0>
0C
#424730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#424740000000
0!
0*
09
0>
0C
#424750000000
1!
1*
b1 6
19
1>
1C
b1 G
#424760000000
0!
0*
09
0>
0C
#424770000000
1!
1*
b10 6
19
1>
1C
b10 G
#424780000000
0!
0*
09
0>
0C
#424790000000
1!
1*
b11 6
19
1>
1C
b11 G
#424800000000
0!
0*
09
0>
0C
#424810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#424820000000
0!
0*
09
0>
0C
#424830000000
1!
1*
b101 6
19
1>
1C
b101 G
#424840000000
0!
0*
09
0>
0C
#424850000000
1!
1*
b110 6
19
1>
1C
b110 G
#424860000000
0!
0*
09
0>
0C
#424870000000
1!
1*
b111 6
19
1>
1C
b111 G
#424880000000
0!
0*
09
0>
0C
#424890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#424900000000
0!
0*
09
0>
0C
#424910000000
1!
1*
b1 6
19
1>
1C
b1 G
#424920000000
0!
0*
09
0>
0C
#424930000000
1!
1*
b10 6
19
1>
1C
b10 G
#424940000000
0!
0*
09
0>
0C
#424950000000
1!
1*
b11 6
19
1>
1C
b11 G
#424960000000
0!
0*
09
0>
0C
#424970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#424980000000
0!
0*
09
0>
0C
#424990000000
1!
1*
b101 6
19
1>
1C
b101 G
#425000000000
0!
0*
09
0>
0C
#425010000000
1!
1*
b110 6
19
1>
1C
b110 G
#425020000000
0!
0*
09
0>
0C
#425030000000
1!
1*
b111 6
19
1>
1C
b111 G
#425040000000
0!
1"
0*
1+
09
1:
0>
0C
#425050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#425060000000
0!
0*
09
0>
0C
#425070000000
1!
1*
b1 6
19
1>
1C
b1 G
#425080000000
0!
0*
09
0>
0C
#425090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#425100000000
0!
0*
09
0>
0C
#425110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#425120000000
0!
0*
09
0>
0C
#425130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#425140000000
0!
0*
09
0>
0C
#425150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#425160000000
0!
0#
0*
0,
09
0>
0?
0C
#425170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#425180000000
0!
0*
09
0>
0C
#425190000000
1!
1*
19
1>
1C
#425200000000
0!
0*
09
0>
0C
#425210000000
1!
1*
19
1>
1C
#425220000000
0!
0*
09
0>
0C
#425230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#425240000000
0!
0*
09
0>
0C
#425250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#425260000000
0!
0*
09
0>
0C
#425270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#425280000000
0!
0*
09
0>
0C
#425290000000
1!
1*
b10 6
19
1>
1C
b10 G
#425300000000
0!
0*
09
0>
0C
#425310000000
1!
1*
b11 6
19
1>
1C
b11 G
#425320000000
0!
0*
09
0>
0C
#425330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#425340000000
0!
0*
09
0>
0C
#425350000000
1!
1*
b101 6
19
1>
1C
b101 G
#425360000000
0!
0*
09
0>
0C
#425370000000
1!
1*
b110 6
19
1>
1C
b110 G
#425380000000
0!
0*
09
0>
0C
#425390000000
1!
1*
b111 6
19
1>
1C
b111 G
#425400000000
0!
0*
09
0>
0C
#425410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#425420000000
0!
0*
09
0>
0C
#425430000000
1!
1*
b1 6
19
1>
1C
b1 G
#425440000000
0!
0*
09
0>
0C
#425450000000
1!
1*
b10 6
19
1>
1C
b10 G
#425460000000
0!
0*
09
0>
0C
#425470000000
1!
1*
b11 6
19
1>
1C
b11 G
#425480000000
0!
0*
09
0>
0C
#425490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#425500000000
0!
0*
09
0>
0C
#425510000000
1!
1*
b101 6
19
1>
1C
b101 G
#425520000000
0!
0*
09
0>
0C
#425530000000
1!
1*
b110 6
19
1>
1C
b110 G
#425540000000
0!
0*
09
0>
0C
#425550000000
1!
1*
b111 6
19
1>
1C
b111 G
#425560000000
0!
0*
09
0>
0C
#425570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#425580000000
0!
0*
09
0>
0C
#425590000000
1!
1*
b1 6
19
1>
1C
b1 G
#425600000000
0!
0*
09
0>
0C
#425610000000
1!
1*
b10 6
19
1>
1C
b10 G
#425620000000
0!
0*
09
0>
0C
#425630000000
1!
1*
b11 6
19
1>
1C
b11 G
#425640000000
0!
0*
09
0>
0C
#425650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#425660000000
0!
0*
09
0>
0C
#425670000000
1!
1*
b101 6
19
1>
1C
b101 G
#425680000000
0!
0*
09
0>
0C
#425690000000
1!
1*
b110 6
19
1>
1C
b110 G
#425700000000
0!
0*
09
0>
0C
#425710000000
1!
1*
b111 6
19
1>
1C
b111 G
#425720000000
0!
1"
0*
1+
09
1:
0>
0C
#425730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#425740000000
0!
0*
09
0>
0C
#425750000000
1!
1*
b1 6
19
1>
1C
b1 G
#425760000000
0!
0*
09
0>
0C
#425770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#425780000000
0!
0*
09
0>
0C
#425790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#425800000000
0!
0*
09
0>
0C
#425810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#425820000000
0!
0*
09
0>
0C
#425830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#425840000000
0!
0#
0*
0,
09
0>
0?
0C
#425850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#425860000000
0!
0*
09
0>
0C
#425870000000
1!
1*
19
1>
1C
#425880000000
0!
0*
09
0>
0C
#425890000000
1!
1*
19
1>
1C
#425900000000
0!
0*
09
0>
0C
#425910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#425920000000
0!
0*
09
0>
0C
#425930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#425940000000
0!
0*
09
0>
0C
#425950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#425960000000
0!
0*
09
0>
0C
#425970000000
1!
1*
b10 6
19
1>
1C
b10 G
#425980000000
0!
0*
09
0>
0C
#425990000000
1!
1*
b11 6
19
1>
1C
b11 G
#426000000000
0!
0*
09
0>
0C
#426010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#426020000000
0!
0*
09
0>
0C
#426030000000
1!
1*
b101 6
19
1>
1C
b101 G
#426040000000
0!
0*
09
0>
0C
#426050000000
1!
1*
b110 6
19
1>
1C
b110 G
#426060000000
0!
0*
09
0>
0C
#426070000000
1!
1*
b111 6
19
1>
1C
b111 G
#426080000000
0!
0*
09
0>
0C
#426090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#426100000000
0!
0*
09
0>
0C
#426110000000
1!
1*
b1 6
19
1>
1C
b1 G
#426120000000
0!
0*
09
0>
0C
#426130000000
1!
1*
b10 6
19
1>
1C
b10 G
#426140000000
0!
0*
09
0>
0C
#426150000000
1!
1*
b11 6
19
1>
1C
b11 G
#426160000000
0!
0*
09
0>
0C
#426170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#426180000000
0!
0*
09
0>
0C
#426190000000
1!
1*
b101 6
19
1>
1C
b101 G
#426200000000
0!
0*
09
0>
0C
#426210000000
1!
1*
b110 6
19
1>
1C
b110 G
#426220000000
0!
0*
09
0>
0C
#426230000000
1!
1*
b111 6
19
1>
1C
b111 G
#426240000000
0!
0*
09
0>
0C
#426250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#426260000000
0!
0*
09
0>
0C
#426270000000
1!
1*
b1 6
19
1>
1C
b1 G
#426280000000
0!
0*
09
0>
0C
#426290000000
1!
1*
b10 6
19
1>
1C
b10 G
#426300000000
0!
0*
09
0>
0C
#426310000000
1!
1*
b11 6
19
1>
1C
b11 G
#426320000000
0!
0*
09
0>
0C
#426330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#426340000000
0!
0*
09
0>
0C
#426350000000
1!
1*
b101 6
19
1>
1C
b101 G
#426360000000
0!
0*
09
0>
0C
#426370000000
1!
1*
b110 6
19
1>
1C
b110 G
#426380000000
0!
0*
09
0>
0C
#426390000000
1!
1*
b111 6
19
1>
1C
b111 G
#426400000000
0!
1"
0*
1+
09
1:
0>
0C
#426410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#426420000000
0!
0*
09
0>
0C
#426430000000
1!
1*
b1 6
19
1>
1C
b1 G
#426440000000
0!
0*
09
0>
0C
#426450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#426460000000
0!
0*
09
0>
0C
#426470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#426480000000
0!
0*
09
0>
0C
#426490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#426500000000
0!
0*
09
0>
0C
#426510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#426520000000
0!
0#
0*
0,
09
0>
0?
0C
#426530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#426540000000
0!
0*
09
0>
0C
#426550000000
1!
1*
19
1>
1C
#426560000000
0!
0*
09
0>
0C
#426570000000
1!
1*
19
1>
1C
#426580000000
0!
0*
09
0>
0C
#426590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#426600000000
0!
0*
09
0>
0C
#426610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#426620000000
0!
0*
09
0>
0C
#426630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#426640000000
0!
0*
09
0>
0C
#426650000000
1!
1*
b10 6
19
1>
1C
b10 G
#426660000000
0!
0*
09
0>
0C
#426670000000
1!
1*
b11 6
19
1>
1C
b11 G
#426680000000
0!
0*
09
0>
0C
#426690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#426700000000
0!
0*
09
0>
0C
#426710000000
1!
1*
b101 6
19
1>
1C
b101 G
#426720000000
0!
0*
09
0>
0C
#426730000000
1!
1*
b110 6
19
1>
1C
b110 G
#426740000000
0!
0*
09
0>
0C
#426750000000
1!
1*
b111 6
19
1>
1C
b111 G
#426760000000
0!
0*
09
0>
0C
#426770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#426780000000
0!
0*
09
0>
0C
#426790000000
1!
1*
b1 6
19
1>
1C
b1 G
#426800000000
0!
0*
09
0>
0C
#426810000000
1!
1*
b10 6
19
1>
1C
b10 G
#426820000000
0!
0*
09
0>
0C
#426830000000
1!
1*
b11 6
19
1>
1C
b11 G
#426840000000
0!
0*
09
0>
0C
#426850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#426860000000
0!
0*
09
0>
0C
#426870000000
1!
1*
b101 6
19
1>
1C
b101 G
#426880000000
0!
0*
09
0>
0C
#426890000000
1!
1*
b110 6
19
1>
1C
b110 G
#426900000000
0!
0*
09
0>
0C
#426910000000
1!
1*
b111 6
19
1>
1C
b111 G
#426920000000
0!
0*
09
0>
0C
#426930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#426940000000
0!
0*
09
0>
0C
#426950000000
1!
1*
b1 6
19
1>
1C
b1 G
#426960000000
0!
0*
09
0>
0C
#426970000000
1!
1*
b10 6
19
1>
1C
b10 G
#426980000000
0!
0*
09
0>
0C
#426990000000
1!
1*
b11 6
19
1>
1C
b11 G
#427000000000
0!
0*
09
0>
0C
#427010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#427020000000
0!
0*
09
0>
0C
#427030000000
1!
1*
b101 6
19
1>
1C
b101 G
#427040000000
0!
0*
09
0>
0C
#427050000000
1!
1*
b110 6
19
1>
1C
b110 G
#427060000000
0!
0*
09
0>
0C
#427070000000
1!
1*
b111 6
19
1>
1C
b111 G
#427080000000
0!
1"
0*
1+
09
1:
0>
0C
#427090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#427100000000
0!
0*
09
0>
0C
#427110000000
1!
1*
b1 6
19
1>
1C
b1 G
#427120000000
0!
0*
09
0>
0C
#427130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#427140000000
0!
0*
09
0>
0C
#427150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#427160000000
0!
0*
09
0>
0C
#427170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#427180000000
0!
0*
09
0>
0C
#427190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#427200000000
0!
0#
0*
0,
09
0>
0?
0C
#427210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#427220000000
0!
0*
09
0>
0C
#427230000000
1!
1*
19
1>
1C
#427240000000
0!
0*
09
0>
0C
#427250000000
1!
1*
19
1>
1C
#427260000000
0!
0*
09
0>
0C
#427270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#427280000000
0!
0*
09
0>
0C
#427290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#427300000000
0!
0*
09
0>
0C
#427310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#427320000000
0!
0*
09
0>
0C
#427330000000
1!
1*
b10 6
19
1>
1C
b10 G
#427340000000
0!
0*
09
0>
0C
#427350000000
1!
1*
b11 6
19
1>
1C
b11 G
#427360000000
0!
0*
09
0>
0C
#427370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#427380000000
0!
0*
09
0>
0C
#427390000000
1!
1*
b101 6
19
1>
1C
b101 G
#427400000000
0!
0*
09
0>
0C
#427410000000
1!
1*
b110 6
19
1>
1C
b110 G
#427420000000
0!
0*
09
0>
0C
#427430000000
1!
1*
b111 6
19
1>
1C
b111 G
#427440000000
0!
0*
09
0>
0C
#427450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#427460000000
0!
0*
09
0>
0C
#427470000000
1!
1*
b1 6
19
1>
1C
b1 G
#427480000000
0!
0*
09
0>
0C
#427490000000
1!
1*
b10 6
19
1>
1C
b10 G
#427500000000
0!
0*
09
0>
0C
#427510000000
1!
1*
b11 6
19
1>
1C
b11 G
#427520000000
0!
0*
09
0>
0C
#427530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#427540000000
0!
0*
09
0>
0C
#427550000000
1!
1*
b101 6
19
1>
1C
b101 G
#427560000000
0!
0*
09
0>
0C
#427570000000
1!
1*
b110 6
19
1>
1C
b110 G
#427580000000
0!
0*
09
0>
0C
#427590000000
1!
1*
b111 6
19
1>
1C
b111 G
#427600000000
0!
0*
09
0>
0C
#427610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#427620000000
0!
0*
09
0>
0C
#427630000000
1!
1*
b1 6
19
1>
1C
b1 G
#427640000000
0!
0*
09
0>
0C
#427650000000
1!
1*
b10 6
19
1>
1C
b10 G
#427660000000
0!
0*
09
0>
0C
#427670000000
1!
1*
b11 6
19
1>
1C
b11 G
#427680000000
0!
0*
09
0>
0C
#427690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#427700000000
0!
0*
09
0>
0C
#427710000000
1!
1*
b101 6
19
1>
1C
b101 G
#427720000000
0!
0*
09
0>
0C
#427730000000
1!
1*
b110 6
19
1>
1C
b110 G
#427740000000
0!
0*
09
0>
0C
#427750000000
1!
1*
b111 6
19
1>
1C
b111 G
#427760000000
0!
1"
0*
1+
09
1:
0>
0C
#427770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#427780000000
0!
0*
09
0>
0C
#427790000000
1!
1*
b1 6
19
1>
1C
b1 G
#427800000000
0!
0*
09
0>
0C
#427810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#427820000000
0!
0*
09
0>
0C
#427830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#427840000000
0!
0*
09
0>
0C
#427850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#427860000000
0!
0*
09
0>
0C
#427870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#427880000000
0!
0#
0*
0,
09
0>
0?
0C
#427890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#427900000000
0!
0*
09
0>
0C
#427910000000
1!
1*
19
1>
1C
#427920000000
0!
0*
09
0>
0C
#427930000000
1!
1*
19
1>
1C
#427940000000
0!
0*
09
0>
0C
#427950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#427960000000
0!
0*
09
0>
0C
#427970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#427980000000
0!
0*
09
0>
0C
#427990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#428000000000
0!
0*
09
0>
0C
#428010000000
1!
1*
b10 6
19
1>
1C
b10 G
#428020000000
0!
0*
09
0>
0C
#428030000000
1!
1*
b11 6
19
1>
1C
b11 G
#428040000000
0!
0*
09
0>
0C
#428050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#428060000000
0!
0*
09
0>
0C
#428070000000
1!
1*
b101 6
19
1>
1C
b101 G
#428080000000
0!
0*
09
0>
0C
#428090000000
1!
1*
b110 6
19
1>
1C
b110 G
#428100000000
0!
0*
09
0>
0C
#428110000000
1!
1*
b111 6
19
1>
1C
b111 G
#428120000000
0!
0*
09
0>
0C
#428130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#428140000000
0!
0*
09
0>
0C
#428150000000
1!
1*
b1 6
19
1>
1C
b1 G
#428160000000
0!
0*
09
0>
0C
#428170000000
1!
1*
b10 6
19
1>
1C
b10 G
#428180000000
0!
0*
09
0>
0C
#428190000000
1!
1*
b11 6
19
1>
1C
b11 G
#428200000000
0!
0*
09
0>
0C
#428210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#428220000000
0!
0*
09
0>
0C
#428230000000
1!
1*
b101 6
19
1>
1C
b101 G
#428240000000
0!
0*
09
0>
0C
#428250000000
1!
1*
b110 6
19
1>
1C
b110 G
#428260000000
0!
0*
09
0>
0C
#428270000000
1!
1*
b111 6
19
1>
1C
b111 G
#428280000000
0!
0*
09
0>
0C
#428290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#428300000000
0!
0*
09
0>
0C
#428310000000
1!
1*
b1 6
19
1>
1C
b1 G
#428320000000
0!
0*
09
0>
0C
#428330000000
1!
1*
b10 6
19
1>
1C
b10 G
#428340000000
0!
0*
09
0>
0C
#428350000000
1!
1*
b11 6
19
1>
1C
b11 G
#428360000000
0!
0*
09
0>
0C
#428370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#428380000000
0!
0*
09
0>
0C
#428390000000
1!
1*
b101 6
19
1>
1C
b101 G
#428400000000
0!
0*
09
0>
0C
#428410000000
1!
1*
b110 6
19
1>
1C
b110 G
#428420000000
0!
0*
09
0>
0C
#428430000000
1!
1*
b111 6
19
1>
1C
b111 G
#428440000000
0!
1"
0*
1+
09
1:
0>
0C
#428450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#428460000000
0!
0*
09
0>
0C
#428470000000
1!
1*
b1 6
19
1>
1C
b1 G
#428480000000
0!
0*
09
0>
0C
#428490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#428500000000
0!
0*
09
0>
0C
#428510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#428520000000
0!
0*
09
0>
0C
#428530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#428540000000
0!
0*
09
0>
0C
#428550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#428560000000
0!
0#
0*
0,
09
0>
0?
0C
#428570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#428580000000
0!
0*
09
0>
0C
#428590000000
1!
1*
19
1>
1C
#428600000000
0!
0*
09
0>
0C
#428610000000
1!
1*
19
1>
1C
#428620000000
0!
0*
09
0>
0C
#428630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#428640000000
0!
0*
09
0>
0C
#428650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#428660000000
0!
0*
09
0>
0C
#428670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#428680000000
0!
0*
09
0>
0C
#428690000000
1!
1*
b10 6
19
1>
1C
b10 G
#428700000000
0!
0*
09
0>
0C
#428710000000
1!
1*
b11 6
19
1>
1C
b11 G
#428720000000
0!
0*
09
0>
0C
#428730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#428740000000
0!
0*
09
0>
0C
#428750000000
1!
1*
b101 6
19
1>
1C
b101 G
#428760000000
0!
0*
09
0>
0C
#428770000000
1!
1*
b110 6
19
1>
1C
b110 G
#428780000000
0!
0*
09
0>
0C
#428790000000
1!
1*
b111 6
19
1>
1C
b111 G
#428800000000
0!
0*
09
0>
0C
#428810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#428820000000
0!
0*
09
0>
0C
#428830000000
1!
1*
b1 6
19
1>
1C
b1 G
#428840000000
0!
0*
09
0>
0C
#428850000000
1!
1*
b10 6
19
1>
1C
b10 G
#428860000000
0!
0*
09
0>
0C
#428870000000
1!
1*
b11 6
19
1>
1C
b11 G
#428880000000
0!
0*
09
0>
0C
#428890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#428900000000
0!
0*
09
0>
0C
#428910000000
1!
1*
b101 6
19
1>
1C
b101 G
#428920000000
0!
0*
09
0>
0C
#428930000000
1!
1*
b110 6
19
1>
1C
b110 G
#428940000000
0!
0*
09
0>
0C
#428950000000
1!
1*
b111 6
19
1>
1C
b111 G
#428960000000
0!
0*
09
0>
0C
#428970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#428980000000
0!
0*
09
0>
0C
#428990000000
1!
1*
b1 6
19
1>
1C
b1 G
#429000000000
0!
0*
09
0>
0C
#429010000000
1!
1*
b10 6
19
1>
1C
b10 G
#429020000000
0!
0*
09
0>
0C
#429030000000
1!
1*
b11 6
19
1>
1C
b11 G
#429040000000
0!
0*
09
0>
0C
#429050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#429060000000
0!
0*
09
0>
0C
#429070000000
1!
1*
b101 6
19
1>
1C
b101 G
#429080000000
0!
0*
09
0>
0C
#429090000000
1!
1*
b110 6
19
1>
1C
b110 G
#429100000000
0!
0*
09
0>
0C
#429110000000
1!
1*
b111 6
19
1>
1C
b111 G
#429120000000
0!
1"
0*
1+
09
1:
0>
0C
#429130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#429140000000
0!
0*
09
0>
0C
#429150000000
1!
1*
b1 6
19
1>
1C
b1 G
#429160000000
0!
0*
09
0>
0C
#429170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#429180000000
0!
0*
09
0>
0C
#429190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#429200000000
0!
0*
09
0>
0C
#429210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#429220000000
0!
0*
09
0>
0C
#429230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#429240000000
0!
0#
0*
0,
09
0>
0?
0C
#429250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#429260000000
0!
0*
09
0>
0C
#429270000000
1!
1*
19
1>
1C
#429280000000
0!
0*
09
0>
0C
#429290000000
1!
1*
19
1>
1C
#429300000000
0!
0*
09
0>
0C
#429310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#429320000000
0!
0*
09
0>
0C
#429330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#429340000000
0!
0*
09
0>
0C
#429350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#429360000000
0!
0*
09
0>
0C
#429370000000
1!
1*
b10 6
19
1>
1C
b10 G
#429380000000
0!
0*
09
0>
0C
#429390000000
1!
1*
b11 6
19
1>
1C
b11 G
#429400000000
0!
0*
09
0>
0C
#429410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#429420000000
0!
0*
09
0>
0C
#429430000000
1!
1*
b101 6
19
1>
1C
b101 G
#429440000000
0!
0*
09
0>
0C
#429450000000
1!
1*
b110 6
19
1>
1C
b110 G
#429460000000
0!
0*
09
0>
0C
#429470000000
1!
1*
b111 6
19
1>
1C
b111 G
#429480000000
0!
0*
09
0>
0C
#429490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#429500000000
0!
0*
09
0>
0C
#429510000000
1!
1*
b1 6
19
1>
1C
b1 G
#429520000000
0!
0*
09
0>
0C
#429530000000
1!
1*
b10 6
19
1>
1C
b10 G
#429540000000
0!
0*
09
0>
0C
#429550000000
1!
1*
b11 6
19
1>
1C
b11 G
#429560000000
0!
0*
09
0>
0C
#429570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#429580000000
0!
0*
09
0>
0C
#429590000000
1!
1*
b101 6
19
1>
1C
b101 G
#429600000000
0!
0*
09
0>
0C
#429610000000
1!
1*
b110 6
19
1>
1C
b110 G
#429620000000
0!
0*
09
0>
0C
#429630000000
1!
1*
b111 6
19
1>
1C
b111 G
#429640000000
0!
0*
09
0>
0C
#429650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#429660000000
0!
0*
09
0>
0C
#429670000000
1!
1*
b1 6
19
1>
1C
b1 G
#429680000000
0!
0*
09
0>
0C
#429690000000
1!
1*
b10 6
19
1>
1C
b10 G
#429700000000
0!
0*
09
0>
0C
#429710000000
1!
1*
b11 6
19
1>
1C
b11 G
#429720000000
0!
0*
09
0>
0C
#429730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#429740000000
0!
0*
09
0>
0C
#429750000000
1!
1*
b101 6
19
1>
1C
b101 G
#429760000000
0!
0*
09
0>
0C
#429770000000
1!
1*
b110 6
19
1>
1C
b110 G
#429780000000
0!
0*
09
0>
0C
#429790000000
1!
1*
b111 6
19
1>
1C
b111 G
#429800000000
0!
1"
0*
1+
09
1:
0>
0C
#429810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#429820000000
0!
0*
09
0>
0C
#429830000000
1!
1*
b1 6
19
1>
1C
b1 G
#429840000000
0!
0*
09
0>
0C
#429850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#429860000000
0!
0*
09
0>
0C
#429870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#429880000000
0!
0*
09
0>
0C
#429890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#429900000000
0!
0*
09
0>
0C
#429910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#429920000000
0!
0#
0*
0,
09
0>
0?
0C
#429930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#429940000000
0!
0*
09
0>
0C
#429950000000
1!
1*
19
1>
1C
#429960000000
0!
0*
09
0>
0C
#429970000000
1!
1*
19
1>
1C
#429980000000
0!
0*
09
0>
0C
#429990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#430000000000
0!
0*
09
0>
0C
#430010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#430020000000
0!
0*
09
0>
0C
#430030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#430040000000
0!
0*
09
0>
0C
#430050000000
1!
1*
b10 6
19
1>
1C
b10 G
#430060000000
0!
0*
09
0>
0C
#430070000000
1!
1*
b11 6
19
1>
1C
b11 G
#430080000000
0!
0*
09
0>
0C
#430090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#430100000000
0!
0*
09
0>
0C
#430110000000
1!
1*
b101 6
19
1>
1C
b101 G
#430120000000
0!
0*
09
0>
0C
#430130000000
1!
1*
b110 6
19
1>
1C
b110 G
#430140000000
0!
0*
09
0>
0C
#430150000000
1!
1*
b111 6
19
1>
1C
b111 G
#430160000000
0!
0*
09
0>
0C
#430170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#430180000000
0!
0*
09
0>
0C
#430190000000
1!
1*
b1 6
19
1>
1C
b1 G
#430200000000
0!
0*
09
0>
0C
#430210000000
1!
1*
b10 6
19
1>
1C
b10 G
#430220000000
0!
0*
09
0>
0C
#430230000000
1!
1*
b11 6
19
1>
1C
b11 G
#430240000000
0!
0*
09
0>
0C
#430250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#430260000000
0!
0*
09
0>
0C
#430270000000
1!
1*
b101 6
19
1>
1C
b101 G
#430280000000
0!
0*
09
0>
0C
#430290000000
1!
1*
b110 6
19
1>
1C
b110 G
#430300000000
0!
0*
09
0>
0C
#430310000000
1!
1*
b111 6
19
1>
1C
b111 G
#430320000000
0!
0*
09
0>
0C
#430330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#430340000000
0!
0*
09
0>
0C
#430350000000
1!
1*
b1 6
19
1>
1C
b1 G
#430360000000
0!
0*
09
0>
0C
#430370000000
1!
1*
b10 6
19
1>
1C
b10 G
#430380000000
0!
0*
09
0>
0C
#430390000000
1!
1*
b11 6
19
1>
1C
b11 G
#430400000000
0!
0*
09
0>
0C
#430410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#430420000000
0!
0*
09
0>
0C
#430430000000
1!
1*
b101 6
19
1>
1C
b101 G
#430440000000
0!
0*
09
0>
0C
#430450000000
1!
1*
b110 6
19
1>
1C
b110 G
#430460000000
0!
0*
09
0>
0C
#430470000000
1!
1*
b111 6
19
1>
1C
b111 G
#430480000000
0!
1"
0*
1+
09
1:
0>
0C
#430490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#430500000000
0!
0*
09
0>
0C
#430510000000
1!
1*
b1 6
19
1>
1C
b1 G
#430520000000
0!
0*
09
0>
0C
#430530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#430540000000
0!
0*
09
0>
0C
#430550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#430560000000
0!
0*
09
0>
0C
#430570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#430580000000
0!
0*
09
0>
0C
#430590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#430600000000
0!
0#
0*
0,
09
0>
0?
0C
#430610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#430620000000
0!
0*
09
0>
0C
#430630000000
1!
1*
19
1>
1C
#430640000000
0!
0*
09
0>
0C
#430650000000
1!
1*
19
1>
1C
#430660000000
0!
0*
09
0>
0C
#430670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#430680000000
0!
0*
09
0>
0C
#430690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#430700000000
0!
0*
09
0>
0C
#430710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#430720000000
0!
0*
09
0>
0C
#430730000000
1!
1*
b10 6
19
1>
1C
b10 G
#430740000000
0!
0*
09
0>
0C
#430750000000
1!
1*
b11 6
19
1>
1C
b11 G
#430760000000
0!
0*
09
0>
0C
#430770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#430780000000
0!
0*
09
0>
0C
#430790000000
1!
1*
b101 6
19
1>
1C
b101 G
#430800000000
0!
0*
09
0>
0C
#430810000000
1!
1*
b110 6
19
1>
1C
b110 G
#430820000000
0!
0*
09
0>
0C
#430830000000
1!
1*
b111 6
19
1>
1C
b111 G
#430840000000
0!
0*
09
0>
0C
#430850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#430860000000
0!
0*
09
0>
0C
#430870000000
1!
1*
b1 6
19
1>
1C
b1 G
#430880000000
0!
0*
09
0>
0C
#430890000000
1!
1*
b10 6
19
1>
1C
b10 G
#430900000000
0!
0*
09
0>
0C
#430910000000
1!
1*
b11 6
19
1>
1C
b11 G
#430920000000
0!
0*
09
0>
0C
#430930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#430940000000
0!
0*
09
0>
0C
#430950000000
1!
1*
b101 6
19
1>
1C
b101 G
#430960000000
0!
0*
09
0>
0C
#430970000000
1!
1*
b110 6
19
1>
1C
b110 G
#430980000000
0!
0*
09
0>
0C
#430990000000
1!
1*
b111 6
19
1>
1C
b111 G
#431000000000
0!
0*
09
0>
0C
#431010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#431020000000
0!
0*
09
0>
0C
#431030000000
1!
1*
b1 6
19
1>
1C
b1 G
#431040000000
0!
0*
09
0>
0C
#431050000000
1!
1*
b10 6
19
1>
1C
b10 G
#431060000000
0!
0*
09
0>
0C
#431070000000
1!
1*
b11 6
19
1>
1C
b11 G
#431080000000
0!
0*
09
0>
0C
#431090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#431100000000
0!
0*
09
0>
0C
#431110000000
1!
1*
b101 6
19
1>
1C
b101 G
#431120000000
0!
0*
09
0>
0C
#431130000000
1!
1*
b110 6
19
1>
1C
b110 G
#431140000000
0!
0*
09
0>
0C
#431150000000
1!
1*
b111 6
19
1>
1C
b111 G
#431160000000
0!
1"
0*
1+
09
1:
0>
0C
#431170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#431180000000
0!
0*
09
0>
0C
#431190000000
1!
1*
b1 6
19
1>
1C
b1 G
#431200000000
0!
0*
09
0>
0C
#431210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#431220000000
0!
0*
09
0>
0C
#431230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#431240000000
0!
0*
09
0>
0C
#431250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#431260000000
0!
0*
09
0>
0C
#431270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#431280000000
0!
0#
0*
0,
09
0>
0?
0C
#431290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#431300000000
0!
0*
09
0>
0C
#431310000000
1!
1*
19
1>
1C
#431320000000
0!
0*
09
0>
0C
#431330000000
1!
1*
19
1>
1C
#431340000000
0!
0*
09
0>
0C
#431350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#431360000000
0!
0*
09
0>
0C
#431370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#431380000000
0!
0*
09
0>
0C
#431390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#431400000000
0!
0*
09
0>
0C
#431410000000
1!
1*
b10 6
19
1>
1C
b10 G
#431420000000
0!
0*
09
0>
0C
#431430000000
1!
1*
b11 6
19
1>
1C
b11 G
#431440000000
0!
0*
09
0>
0C
#431450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#431460000000
0!
0*
09
0>
0C
#431470000000
1!
1*
b101 6
19
1>
1C
b101 G
#431480000000
0!
0*
09
0>
0C
#431490000000
1!
1*
b110 6
19
1>
1C
b110 G
#431500000000
0!
0*
09
0>
0C
#431510000000
1!
1*
b111 6
19
1>
1C
b111 G
#431520000000
0!
0*
09
0>
0C
#431530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#431540000000
0!
0*
09
0>
0C
#431550000000
1!
1*
b1 6
19
1>
1C
b1 G
#431560000000
0!
0*
09
0>
0C
#431570000000
1!
1*
b10 6
19
1>
1C
b10 G
#431580000000
0!
0*
09
0>
0C
#431590000000
1!
1*
b11 6
19
1>
1C
b11 G
#431600000000
0!
0*
09
0>
0C
#431610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#431620000000
0!
0*
09
0>
0C
#431630000000
1!
1*
b101 6
19
1>
1C
b101 G
#431640000000
0!
0*
09
0>
0C
#431650000000
1!
1*
b110 6
19
1>
1C
b110 G
#431660000000
0!
0*
09
0>
0C
#431670000000
1!
1*
b111 6
19
1>
1C
b111 G
#431680000000
0!
0*
09
0>
0C
#431690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#431700000000
0!
0*
09
0>
0C
#431710000000
1!
1*
b1 6
19
1>
1C
b1 G
#431720000000
0!
0*
09
0>
0C
#431730000000
1!
1*
b10 6
19
1>
1C
b10 G
#431740000000
0!
0*
09
0>
0C
#431750000000
1!
1*
b11 6
19
1>
1C
b11 G
#431760000000
0!
0*
09
0>
0C
#431770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#431780000000
0!
0*
09
0>
0C
#431790000000
1!
1*
b101 6
19
1>
1C
b101 G
#431800000000
0!
0*
09
0>
0C
#431810000000
1!
1*
b110 6
19
1>
1C
b110 G
#431820000000
0!
0*
09
0>
0C
#431830000000
1!
1*
b111 6
19
1>
1C
b111 G
#431840000000
0!
1"
0*
1+
09
1:
0>
0C
#431850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#431860000000
0!
0*
09
0>
0C
#431870000000
1!
1*
b1 6
19
1>
1C
b1 G
#431880000000
0!
0*
09
0>
0C
#431890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#431900000000
0!
0*
09
0>
0C
#431910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#431920000000
0!
0*
09
0>
0C
#431930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#431940000000
0!
0*
09
0>
0C
#431950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#431960000000
0!
0#
0*
0,
09
0>
0?
0C
#431970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#431980000000
0!
0*
09
0>
0C
#431990000000
1!
1*
19
1>
1C
#432000000000
0!
0*
09
0>
0C
#432010000000
1!
1*
19
1>
1C
#432020000000
0!
0*
09
0>
0C
#432030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#432040000000
0!
0*
09
0>
0C
#432050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#432060000000
0!
0*
09
0>
0C
#432070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#432080000000
0!
0*
09
0>
0C
#432090000000
1!
1*
b10 6
19
1>
1C
b10 G
#432100000000
0!
0*
09
0>
0C
#432110000000
1!
1*
b11 6
19
1>
1C
b11 G
#432120000000
0!
0*
09
0>
0C
#432130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#432140000000
0!
0*
09
0>
0C
#432150000000
1!
1*
b101 6
19
1>
1C
b101 G
#432160000000
0!
0*
09
0>
0C
#432170000000
1!
1*
b110 6
19
1>
1C
b110 G
#432180000000
0!
0*
09
0>
0C
#432190000000
1!
1*
b111 6
19
1>
1C
b111 G
#432200000000
0!
0*
09
0>
0C
#432210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#432220000000
0!
0*
09
0>
0C
#432230000000
1!
1*
b1 6
19
1>
1C
b1 G
#432240000000
0!
0*
09
0>
0C
#432250000000
1!
1*
b10 6
19
1>
1C
b10 G
#432260000000
0!
0*
09
0>
0C
#432270000000
1!
1*
b11 6
19
1>
1C
b11 G
#432280000000
0!
0*
09
0>
0C
#432290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#432300000000
0!
0*
09
0>
0C
#432310000000
1!
1*
b101 6
19
1>
1C
b101 G
#432320000000
0!
0*
09
0>
0C
#432330000000
1!
1*
b110 6
19
1>
1C
b110 G
#432340000000
0!
0*
09
0>
0C
#432350000000
1!
1*
b111 6
19
1>
1C
b111 G
#432360000000
0!
0*
09
0>
0C
#432370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#432380000000
0!
0*
09
0>
0C
#432390000000
1!
1*
b1 6
19
1>
1C
b1 G
#432400000000
0!
0*
09
0>
0C
#432410000000
1!
1*
b10 6
19
1>
1C
b10 G
#432420000000
0!
0*
09
0>
0C
#432430000000
1!
1*
b11 6
19
1>
1C
b11 G
#432440000000
0!
0*
09
0>
0C
#432450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#432460000000
0!
0*
09
0>
0C
#432470000000
1!
1*
b101 6
19
1>
1C
b101 G
#432480000000
0!
0*
09
0>
0C
#432490000000
1!
1*
b110 6
19
1>
1C
b110 G
#432500000000
0!
0*
09
0>
0C
#432510000000
1!
1*
b111 6
19
1>
1C
b111 G
#432520000000
0!
1"
0*
1+
09
1:
0>
0C
#432530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#432540000000
0!
0*
09
0>
0C
#432550000000
1!
1*
b1 6
19
1>
1C
b1 G
#432560000000
0!
0*
09
0>
0C
#432570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#432580000000
0!
0*
09
0>
0C
#432590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#432600000000
0!
0*
09
0>
0C
#432610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#432620000000
0!
0*
09
0>
0C
#432630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#432640000000
0!
0#
0*
0,
09
0>
0?
0C
#432650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#432660000000
0!
0*
09
0>
0C
#432670000000
1!
1*
19
1>
1C
#432680000000
0!
0*
09
0>
0C
#432690000000
1!
1*
19
1>
1C
#432700000000
0!
0*
09
0>
0C
#432710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#432720000000
0!
0*
09
0>
0C
#432730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#432740000000
0!
0*
09
0>
0C
#432750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#432760000000
0!
0*
09
0>
0C
#432770000000
1!
1*
b10 6
19
1>
1C
b10 G
#432780000000
0!
0*
09
0>
0C
#432790000000
1!
1*
b11 6
19
1>
1C
b11 G
#432800000000
0!
0*
09
0>
0C
#432810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#432820000000
0!
0*
09
0>
0C
#432830000000
1!
1*
b101 6
19
1>
1C
b101 G
#432840000000
0!
0*
09
0>
0C
#432850000000
1!
1*
b110 6
19
1>
1C
b110 G
#432860000000
0!
0*
09
0>
0C
#432870000000
1!
1*
b111 6
19
1>
1C
b111 G
#432880000000
0!
0*
09
0>
0C
#432890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#432900000000
0!
0*
09
0>
0C
#432910000000
1!
1*
b1 6
19
1>
1C
b1 G
#432920000000
0!
0*
09
0>
0C
#432930000000
1!
1*
b10 6
19
1>
1C
b10 G
#432940000000
0!
0*
09
0>
0C
#432950000000
1!
1*
b11 6
19
1>
1C
b11 G
#432960000000
0!
0*
09
0>
0C
#432970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#432980000000
0!
0*
09
0>
0C
#432990000000
1!
1*
b101 6
19
1>
1C
b101 G
#433000000000
0!
0*
09
0>
0C
#433010000000
1!
1*
b110 6
19
1>
1C
b110 G
#433020000000
0!
0*
09
0>
0C
#433030000000
1!
1*
b111 6
19
1>
1C
b111 G
#433040000000
0!
0*
09
0>
0C
#433050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#433060000000
0!
0*
09
0>
0C
#433070000000
1!
1*
b1 6
19
1>
1C
b1 G
#433080000000
0!
0*
09
0>
0C
#433090000000
1!
1*
b10 6
19
1>
1C
b10 G
#433100000000
0!
0*
09
0>
0C
#433110000000
1!
1*
b11 6
19
1>
1C
b11 G
#433120000000
0!
0*
09
0>
0C
#433130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#433140000000
0!
0*
09
0>
0C
#433150000000
1!
1*
b101 6
19
1>
1C
b101 G
#433160000000
0!
0*
09
0>
0C
#433170000000
1!
1*
b110 6
19
1>
1C
b110 G
#433180000000
0!
0*
09
0>
0C
#433190000000
1!
1*
b111 6
19
1>
1C
b111 G
#433200000000
0!
1"
0*
1+
09
1:
0>
0C
#433210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#433220000000
0!
0*
09
0>
0C
#433230000000
1!
1*
b1 6
19
1>
1C
b1 G
#433240000000
0!
0*
09
0>
0C
#433250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#433260000000
0!
0*
09
0>
0C
#433270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#433280000000
0!
0*
09
0>
0C
#433290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#433300000000
0!
0*
09
0>
0C
#433310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#433320000000
0!
0#
0*
0,
09
0>
0?
0C
#433330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#433340000000
0!
0*
09
0>
0C
#433350000000
1!
1*
19
1>
1C
#433360000000
0!
0*
09
0>
0C
#433370000000
1!
1*
19
1>
1C
#433380000000
0!
0*
09
0>
0C
#433390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#433400000000
0!
0*
09
0>
0C
#433410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#433420000000
0!
0*
09
0>
0C
#433430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#433440000000
0!
0*
09
0>
0C
#433450000000
1!
1*
b10 6
19
1>
1C
b10 G
#433460000000
0!
0*
09
0>
0C
#433470000000
1!
1*
b11 6
19
1>
1C
b11 G
#433480000000
0!
0*
09
0>
0C
#433490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#433500000000
0!
0*
09
0>
0C
#433510000000
1!
1*
b101 6
19
1>
1C
b101 G
#433520000000
0!
0*
09
0>
0C
#433530000000
1!
1*
b110 6
19
1>
1C
b110 G
#433540000000
0!
0*
09
0>
0C
#433550000000
1!
1*
b111 6
19
1>
1C
b111 G
#433560000000
0!
0*
09
0>
0C
#433570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#433580000000
0!
0*
09
0>
0C
#433590000000
1!
1*
b1 6
19
1>
1C
b1 G
#433600000000
0!
0*
09
0>
0C
#433610000000
1!
1*
b10 6
19
1>
1C
b10 G
#433620000000
0!
0*
09
0>
0C
#433630000000
1!
1*
b11 6
19
1>
1C
b11 G
#433640000000
0!
0*
09
0>
0C
#433650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#433660000000
0!
0*
09
0>
0C
#433670000000
1!
1*
b101 6
19
1>
1C
b101 G
#433680000000
0!
0*
09
0>
0C
#433690000000
1!
1*
b110 6
19
1>
1C
b110 G
#433700000000
0!
0*
09
0>
0C
#433710000000
1!
1*
b111 6
19
1>
1C
b111 G
#433720000000
0!
0*
09
0>
0C
#433730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#433740000000
0!
0*
09
0>
0C
#433750000000
1!
1*
b1 6
19
1>
1C
b1 G
#433760000000
0!
0*
09
0>
0C
#433770000000
1!
1*
b10 6
19
1>
1C
b10 G
#433780000000
0!
0*
09
0>
0C
#433790000000
1!
1*
b11 6
19
1>
1C
b11 G
#433800000000
0!
0*
09
0>
0C
#433810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#433820000000
0!
0*
09
0>
0C
#433830000000
1!
1*
b101 6
19
1>
1C
b101 G
#433840000000
0!
0*
09
0>
0C
#433850000000
1!
1*
b110 6
19
1>
1C
b110 G
#433860000000
0!
0*
09
0>
0C
#433870000000
1!
1*
b111 6
19
1>
1C
b111 G
#433880000000
0!
1"
0*
1+
09
1:
0>
0C
#433890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#433900000000
0!
0*
09
0>
0C
#433910000000
1!
1*
b1 6
19
1>
1C
b1 G
#433920000000
0!
0*
09
0>
0C
#433930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#433940000000
0!
0*
09
0>
0C
#433950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#433960000000
0!
0*
09
0>
0C
#433970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#433980000000
0!
0*
09
0>
0C
#433990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#434000000000
0!
0#
0*
0,
09
0>
0?
0C
#434010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#434020000000
0!
0*
09
0>
0C
#434030000000
1!
1*
19
1>
1C
#434040000000
0!
0*
09
0>
0C
#434050000000
1!
1*
19
1>
1C
#434060000000
0!
0*
09
0>
0C
#434070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#434080000000
0!
0*
09
0>
0C
#434090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#434100000000
0!
0*
09
0>
0C
#434110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#434120000000
0!
0*
09
0>
0C
#434130000000
1!
1*
b10 6
19
1>
1C
b10 G
#434140000000
0!
0*
09
0>
0C
#434150000000
1!
1*
b11 6
19
1>
1C
b11 G
#434160000000
0!
0*
09
0>
0C
#434170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#434180000000
0!
0*
09
0>
0C
#434190000000
1!
1*
b101 6
19
1>
1C
b101 G
#434200000000
0!
0*
09
0>
0C
#434210000000
1!
1*
b110 6
19
1>
1C
b110 G
#434220000000
0!
0*
09
0>
0C
#434230000000
1!
1*
b111 6
19
1>
1C
b111 G
#434240000000
0!
0*
09
0>
0C
#434250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#434260000000
0!
0*
09
0>
0C
#434270000000
1!
1*
b1 6
19
1>
1C
b1 G
#434280000000
0!
0*
09
0>
0C
#434290000000
1!
1*
b10 6
19
1>
1C
b10 G
#434300000000
0!
0*
09
0>
0C
#434310000000
1!
1*
b11 6
19
1>
1C
b11 G
#434320000000
0!
0*
09
0>
0C
#434330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#434340000000
0!
0*
09
0>
0C
#434350000000
1!
1*
b101 6
19
1>
1C
b101 G
#434360000000
0!
0*
09
0>
0C
#434370000000
1!
1*
b110 6
19
1>
1C
b110 G
#434380000000
0!
0*
09
0>
0C
#434390000000
1!
1*
b111 6
19
1>
1C
b111 G
#434400000000
0!
0*
09
0>
0C
#434410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#434420000000
0!
0*
09
0>
0C
#434430000000
1!
1*
b1 6
19
1>
1C
b1 G
#434440000000
0!
0*
09
0>
0C
#434450000000
1!
1*
b10 6
19
1>
1C
b10 G
#434460000000
0!
0*
09
0>
0C
#434470000000
1!
1*
b11 6
19
1>
1C
b11 G
#434480000000
0!
0*
09
0>
0C
#434490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#434500000000
0!
0*
09
0>
0C
#434510000000
1!
1*
b101 6
19
1>
1C
b101 G
#434520000000
0!
0*
09
0>
0C
#434530000000
1!
1*
b110 6
19
1>
1C
b110 G
#434540000000
0!
0*
09
0>
0C
#434550000000
1!
1*
b111 6
19
1>
1C
b111 G
#434560000000
0!
1"
0*
1+
09
1:
0>
0C
#434570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#434580000000
0!
0*
09
0>
0C
#434590000000
1!
1*
b1 6
19
1>
1C
b1 G
#434600000000
0!
0*
09
0>
0C
#434610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#434620000000
0!
0*
09
0>
0C
#434630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#434640000000
0!
0*
09
0>
0C
#434650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#434660000000
0!
0*
09
0>
0C
#434670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#434680000000
0!
0#
0*
0,
09
0>
0?
0C
#434690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#434700000000
0!
0*
09
0>
0C
#434710000000
1!
1*
19
1>
1C
#434720000000
0!
0*
09
0>
0C
#434730000000
1!
1*
19
1>
1C
#434740000000
0!
0*
09
0>
0C
#434750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#434760000000
0!
0*
09
0>
0C
#434770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#434780000000
0!
0*
09
0>
0C
#434790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#434800000000
0!
0*
09
0>
0C
#434810000000
1!
1*
b10 6
19
1>
1C
b10 G
#434820000000
0!
0*
09
0>
0C
#434830000000
1!
1*
b11 6
19
1>
1C
b11 G
#434840000000
0!
0*
09
0>
0C
#434850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#434860000000
0!
0*
09
0>
0C
#434870000000
1!
1*
b101 6
19
1>
1C
b101 G
#434880000000
0!
0*
09
0>
0C
#434890000000
1!
1*
b110 6
19
1>
1C
b110 G
#434900000000
0!
0*
09
0>
0C
#434910000000
1!
1*
b111 6
19
1>
1C
b111 G
#434920000000
0!
0*
09
0>
0C
#434930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#434940000000
0!
0*
09
0>
0C
#434950000000
1!
1*
b1 6
19
1>
1C
b1 G
#434960000000
0!
0*
09
0>
0C
#434970000000
1!
1*
b10 6
19
1>
1C
b10 G
#434980000000
0!
0*
09
0>
0C
#434990000000
1!
1*
b11 6
19
1>
1C
b11 G
#435000000000
0!
0*
09
0>
0C
#435010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#435020000000
0!
0*
09
0>
0C
#435030000000
1!
1*
b101 6
19
1>
1C
b101 G
#435040000000
0!
0*
09
0>
0C
#435050000000
1!
1*
b110 6
19
1>
1C
b110 G
#435060000000
0!
0*
09
0>
0C
#435070000000
1!
1*
b111 6
19
1>
1C
b111 G
#435080000000
0!
0*
09
0>
0C
#435090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#435100000000
0!
0*
09
0>
0C
#435110000000
1!
1*
b1 6
19
1>
1C
b1 G
#435120000000
0!
0*
09
0>
0C
#435130000000
1!
1*
b10 6
19
1>
1C
b10 G
#435140000000
0!
0*
09
0>
0C
#435150000000
1!
1*
b11 6
19
1>
1C
b11 G
#435160000000
0!
0*
09
0>
0C
#435170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#435180000000
0!
0*
09
0>
0C
#435190000000
1!
1*
b101 6
19
1>
1C
b101 G
#435200000000
0!
0*
09
0>
0C
#435210000000
1!
1*
b110 6
19
1>
1C
b110 G
#435220000000
0!
0*
09
0>
0C
#435230000000
1!
1*
b111 6
19
1>
1C
b111 G
#435240000000
0!
1"
0*
1+
09
1:
0>
0C
#435250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#435260000000
0!
0*
09
0>
0C
#435270000000
1!
1*
b1 6
19
1>
1C
b1 G
#435280000000
0!
0*
09
0>
0C
#435290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#435300000000
0!
0*
09
0>
0C
#435310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#435320000000
0!
0*
09
0>
0C
#435330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#435340000000
0!
0*
09
0>
0C
#435350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#435360000000
0!
0#
0*
0,
09
0>
0?
0C
#435370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#435380000000
0!
0*
09
0>
0C
#435390000000
1!
1*
19
1>
1C
#435400000000
0!
0*
09
0>
0C
#435410000000
1!
1*
19
1>
1C
#435420000000
0!
0*
09
0>
0C
#435430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#435440000000
0!
0*
09
0>
0C
#435450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#435460000000
0!
0*
09
0>
0C
#435470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#435480000000
0!
0*
09
0>
0C
#435490000000
1!
1*
b10 6
19
1>
1C
b10 G
#435500000000
0!
0*
09
0>
0C
#435510000000
1!
1*
b11 6
19
1>
1C
b11 G
#435520000000
0!
0*
09
0>
0C
#435530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#435540000000
0!
0*
09
0>
0C
#435550000000
1!
1*
b101 6
19
1>
1C
b101 G
#435560000000
0!
0*
09
0>
0C
#435570000000
1!
1*
b110 6
19
1>
1C
b110 G
#435580000000
0!
0*
09
0>
0C
#435590000000
1!
1*
b111 6
19
1>
1C
b111 G
#435600000000
0!
0*
09
0>
0C
#435610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#435620000000
0!
0*
09
0>
0C
#435630000000
1!
1*
b1 6
19
1>
1C
b1 G
#435640000000
0!
0*
09
0>
0C
#435650000000
1!
1*
b10 6
19
1>
1C
b10 G
#435660000000
0!
0*
09
0>
0C
#435670000000
1!
1*
b11 6
19
1>
1C
b11 G
#435680000000
0!
0*
09
0>
0C
#435690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#435700000000
0!
0*
09
0>
0C
#435710000000
1!
1*
b101 6
19
1>
1C
b101 G
#435720000000
0!
0*
09
0>
0C
#435730000000
1!
1*
b110 6
19
1>
1C
b110 G
#435740000000
0!
0*
09
0>
0C
#435750000000
1!
1*
b111 6
19
1>
1C
b111 G
#435760000000
0!
0*
09
0>
0C
#435770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#435780000000
0!
0*
09
0>
0C
#435790000000
1!
1*
b1 6
19
1>
1C
b1 G
#435800000000
0!
0*
09
0>
0C
#435810000000
1!
1*
b10 6
19
1>
1C
b10 G
#435820000000
0!
0*
09
0>
0C
#435830000000
1!
1*
b11 6
19
1>
1C
b11 G
#435840000000
0!
0*
09
0>
0C
#435850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#435860000000
0!
0*
09
0>
0C
#435870000000
1!
1*
b101 6
19
1>
1C
b101 G
#435880000000
0!
0*
09
0>
0C
#435890000000
1!
1*
b110 6
19
1>
1C
b110 G
#435900000000
0!
0*
09
0>
0C
#435910000000
1!
1*
b111 6
19
1>
1C
b111 G
#435920000000
0!
1"
0*
1+
09
1:
0>
0C
#435930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#435940000000
0!
0*
09
0>
0C
#435950000000
1!
1*
b1 6
19
1>
1C
b1 G
#435960000000
0!
0*
09
0>
0C
#435970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#435980000000
0!
0*
09
0>
0C
#435990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#436000000000
0!
0*
09
0>
0C
#436010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#436020000000
0!
0*
09
0>
0C
#436030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#436040000000
0!
0#
0*
0,
09
0>
0?
0C
#436050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#436060000000
0!
0*
09
0>
0C
#436070000000
1!
1*
19
1>
1C
#436080000000
0!
0*
09
0>
0C
#436090000000
1!
1*
19
1>
1C
#436100000000
0!
0*
09
0>
0C
#436110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#436120000000
0!
0*
09
0>
0C
#436130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#436140000000
0!
0*
09
0>
0C
#436150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#436160000000
0!
0*
09
0>
0C
#436170000000
1!
1*
b10 6
19
1>
1C
b10 G
#436180000000
0!
0*
09
0>
0C
#436190000000
1!
1*
b11 6
19
1>
1C
b11 G
#436200000000
0!
0*
09
0>
0C
#436210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#436220000000
0!
0*
09
0>
0C
#436230000000
1!
1*
b101 6
19
1>
1C
b101 G
#436240000000
0!
0*
09
0>
0C
#436250000000
1!
1*
b110 6
19
1>
1C
b110 G
#436260000000
0!
0*
09
0>
0C
#436270000000
1!
1*
b111 6
19
1>
1C
b111 G
#436280000000
0!
0*
09
0>
0C
#436290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#436300000000
0!
0*
09
0>
0C
#436310000000
1!
1*
b1 6
19
1>
1C
b1 G
#436320000000
0!
0*
09
0>
0C
#436330000000
1!
1*
b10 6
19
1>
1C
b10 G
#436340000000
0!
0*
09
0>
0C
#436350000000
1!
1*
b11 6
19
1>
1C
b11 G
#436360000000
0!
0*
09
0>
0C
#436370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#436380000000
0!
0*
09
0>
0C
#436390000000
1!
1*
b101 6
19
1>
1C
b101 G
#436400000000
0!
0*
09
0>
0C
#436410000000
1!
1*
b110 6
19
1>
1C
b110 G
#436420000000
0!
0*
09
0>
0C
#436430000000
1!
1*
b111 6
19
1>
1C
b111 G
#436440000000
0!
0*
09
0>
0C
#436450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#436460000000
0!
0*
09
0>
0C
#436470000000
1!
1*
b1 6
19
1>
1C
b1 G
#436480000000
0!
0*
09
0>
0C
#436490000000
1!
1*
b10 6
19
1>
1C
b10 G
#436500000000
0!
0*
09
0>
0C
#436510000000
1!
1*
b11 6
19
1>
1C
b11 G
#436520000000
0!
0*
09
0>
0C
#436530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#436540000000
0!
0*
09
0>
0C
#436550000000
1!
1*
b101 6
19
1>
1C
b101 G
#436560000000
0!
0*
09
0>
0C
#436570000000
1!
1*
b110 6
19
1>
1C
b110 G
#436580000000
0!
0*
09
0>
0C
#436590000000
1!
1*
b111 6
19
1>
1C
b111 G
#436600000000
0!
1"
0*
1+
09
1:
0>
0C
#436610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#436620000000
0!
0*
09
0>
0C
#436630000000
1!
1*
b1 6
19
1>
1C
b1 G
#436640000000
0!
0*
09
0>
0C
#436650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#436660000000
0!
0*
09
0>
0C
#436670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#436680000000
0!
0*
09
0>
0C
#436690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#436700000000
0!
0*
09
0>
0C
#436710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#436720000000
0!
0#
0*
0,
09
0>
0?
0C
#436730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#436740000000
0!
0*
09
0>
0C
#436750000000
1!
1*
19
1>
1C
#436760000000
0!
0*
09
0>
0C
#436770000000
1!
1*
19
1>
1C
#436780000000
0!
0*
09
0>
0C
#436790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#436800000000
0!
0*
09
0>
0C
#436810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#436820000000
0!
0*
09
0>
0C
#436830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#436840000000
0!
0*
09
0>
0C
#436850000000
1!
1*
b10 6
19
1>
1C
b10 G
#436860000000
0!
0*
09
0>
0C
#436870000000
1!
1*
b11 6
19
1>
1C
b11 G
#436880000000
0!
0*
09
0>
0C
#436890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#436900000000
0!
0*
09
0>
0C
#436910000000
1!
1*
b101 6
19
1>
1C
b101 G
#436920000000
0!
0*
09
0>
0C
#436930000000
1!
1*
b110 6
19
1>
1C
b110 G
#436940000000
0!
0*
09
0>
0C
#436950000000
1!
1*
b111 6
19
1>
1C
b111 G
#436960000000
0!
0*
09
0>
0C
#436970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#436980000000
0!
0*
09
0>
0C
#436990000000
1!
1*
b1 6
19
1>
1C
b1 G
#437000000000
0!
0*
09
0>
0C
#437010000000
1!
1*
b10 6
19
1>
1C
b10 G
#437020000000
0!
0*
09
0>
0C
#437030000000
1!
1*
b11 6
19
1>
1C
b11 G
#437040000000
0!
0*
09
0>
0C
#437050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#437060000000
0!
0*
09
0>
0C
#437070000000
1!
1*
b101 6
19
1>
1C
b101 G
#437080000000
0!
0*
09
0>
0C
#437090000000
1!
1*
b110 6
19
1>
1C
b110 G
#437100000000
0!
0*
09
0>
0C
#437110000000
1!
1*
b111 6
19
1>
1C
b111 G
#437120000000
0!
0*
09
0>
0C
#437130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#437140000000
0!
0*
09
0>
0C
#437150000000
1!
1*
b1 6
19
1>
1C
b1 G
#437160000000
0!
0*
09
0>
0C
#437170000000
1!
1*
b10 6
19
1>
1C
b10 G
#437180000000
0!
0*
09
0>
0C
#437190000000
1!
1*
b11 6
19
1>
1C
b11 G
#437200000000
0!
0*
09
0>
0C
#437210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#437220000000
0!
0*
09
0>
0C
#437230000000
1!
1*
b101 6
19
1>
1C
b101 G
#437240000000
0!
0*
09
0>
0C
#437250000000
1!
1*
b110 6
19
1>
1C
b110 G
#437260000000
0!
0*
09
0>
0C
#437270000000
1!
1*
b111 6
19
1>
1C
b111 G
#437280000000
0!
1"
0*
1+
09
1:
0>
0C
#437290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#437300000000
0!
0*
09
0>
0C
#437310000000
1!
1*
b1 6
19
1>
1C
b1 G
#437320000000
0!
0*
09
0>
0C
#437330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#437340000000
0!
0*
09
0>
0C
#437350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#437360000000
0!
0*
09
0>
0C
#437370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#437380000000
0!
0*
09
0>
0C
#437390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#437400000000
0!
0#
0*
0,
09
0>
0?
0C
#437410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#437420000000
0!
0*
09
0>
0C
#437430000000
1!
1*
19
1>
1C
#437440000000
0!
0*
09
0>
0C
#437450000000
1!
1*
19
1>
1C
#437460000000
0!
0*
09
0>
0C
#437470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#437480000000
0!
0*
09
0>
0C
#437490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#437500000000
0!
0*
09
0>
0C
#437510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#437520000000
0!
0*
09
0>
0C
#437530000000
1!
1*
b10 6
19
1>
1C
b10 G
#437540000000
0!
0*
09
0>
0C
#437550000000
1!
1*
b11 6
19
1>
1C
b11 G
#437560000000
0!
0*
09
0>
0C
#437570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#437580000000
0!
0*
09
0>
0C
#437590000000
1!
1*
b101 6
19
1>
1C
b101 G
#437600000000
0!
0*
09
0>
0C
#437610000000
1!
1*
b110 6
19
1>
1C
b110 G
#437620000000
0!
0*
09
0>
0C
#437630000000
1!
1*
b111 6
19
1>
1C
b111 G
#437640000000
0!
0*
09
0>
0C
#437650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#437660000000
0!
0*
09
0>
0C
#437670000000
1!
1*
b1 6
19
1>
1C
b1 G
#437680000000
0!
0*
09
0>
0C
#437690000000
1!
1*
b10 6
19
1>
1C
b10 G
#437700000000
0!
0*
09
0>
0C
#437710000000
1!
1*
b11 6
19
1>
1C
b11 G
#437720000000
0!
0*
09
0>
0C
#437730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#437740000000
0!
0*
09
0>
0C
#437750000000
1!
1*
b101 6
19
1>
1C
b101 G
#437760000000
0!
0*
09
0>
0C
#437770000000
1!
1*
b110 6
19
1>
1C
b110 G
#437780000000
0!
0*
09
0>
0C
#437790000000
1!
1*
b111 6
19
1>
1C
b111 G
#437800000000
0!
0*
09
0>
0C
#437810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#437820000000
0!
0*
09
0>
0C
#437830000000
1!
1*
b1 6
19
1>
1C
b1 G
#437840000000
0!
0*
09
0>
0C
#437850000000
1!
1*
b10 6
19
1>
1C
b10 G
#437860000000
0!
0*
09
0>
0C
#437870000000
1!
1*
b11 6
19
1>
1C
b11 G
#437880000000
0!
0*
09
0>
0C
#437890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#437900000000
0!
0*
09
0>
0C
#437910000000
1!
1*
b101 6
19
1>
1C
b101 G
#437920000000
0!
0*
09
0>
0C
#437930000000
1!
1*
b110 6
19
1>
1C
b110 G
#437940000000
0!
0*
09
0>
0C
#437950000000
1!
1*
b111 6
19
1>
1C
b111 G
#437960000000
0!
1"
0*
1+
09
1:
0>
0C
#437970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#437980000000
0!
0*
09
0>
0C
#437990000000
1!
1*
b1 6
19
1>
1C
b1 G
#438000000000
0!
0*
09
0>
0C
#438010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#438020000000
0!
0*
09
0>
0C
#438030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#438040000000
0!
0*
09
0>
0C
#438050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#438060000000
0!
0*
09
0>
0C
#438070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#438080000000
0!
0#
0*
0,
09
0>
0?
0C
#438090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#438100000000
0!
0*
09
0>
0C
#438110000000
1!
1*
19
1>
1C
#438120000000
0!
0*
09
0>
0C
#438130000000
1!
1*
19
1>
1C
#438140000000
0!
0*
09
0>
0C
#438150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#438160000000
0!
0*
09
0>
0C
#438170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#438180000000
0!
0*
09
0>
0C
#438190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#438200000000
0!
0*
09
0>
0C
#438210000000
1!
1*
b10 6
19
1>
1C
b10 G
#438220000000
0!
0*
09
0>
0C
#438230000000
1!
1*
b11 6
19
1>
1C
b11 G
#438240000000
0!
0*
09
0>
0C
#438250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#438260000000
0!
0*
09
0>
0C
#438270000000
1!
1*
b101 6
19
1>
1C
b101 G
#438280000000
0!
0*
09
0>
0C
#438290000000
1!
1*
b110 6
19
1>
1C
b110 G
#438300000000
0!
0*
09
0>
0C
#438310000000
1!
1*
b111 6
19
1>
1C
b111 G
#438320000000
0!
0*
09
0>
0C
#438330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#438340000000
0!
0*
09
0>
0C
#438350000000
1!
1*
b1 6
19
1>
1C
b1 G
#438360000000
0!
0*
09
0>
0C
#438370000000
1!
1*
b10 6
19
1>
1C
b10 G
#438380000000
0!
0*
09
0>
0C
#438390000000
1!
1*
b11 6
19
1>
1C
b11 G
#438400000000
0!
0*
09
0>
0C
#438410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#438420000000
0!
0*
09
0>
0C
#438430000000
1!
1*
b101 6
19
1>
1C
b101 G
#438440000000
0!
0*
09
0>
0C
#438450000000
1!
1*
b110 6
19
1>
1C
b110 G
#438460000000
0!
0*
09
0>
0C
#438470000000
1!
1*
b111 6
19
1>
1C
b111 G
#438480000000
0!
0*
09
0>
0C
#438490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#438500000000
0!
0*
09
0>
0C
#438510000000
1!
1*
b1 6
19
1>
1C
b1 G
#438520000000
0!
0*
09
0>
0C
#438530000000
1!
1*
b10 6
19
1>
1C
b10 G
#438540000000
0!
0*
09
0>
0C
#438550000000
1!
1*
b11 6
19
1>
1C
b11 G
#438560000000
0!
0*
09
0>
0C
#438570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#438580000000
0!
0*
09
0>
0C
#438590000000
1!
1*
b101 6
19
1>
1C
b101 G
#438600000000
0!
0*
09
0>
0C
#438610000000
1!
1*
b110 6
19
1>
1C
b110 G
#438620000000
0!
0*
09
0>
0C
#438630000000
1!
1*
b111 6
19
1>
1C
b111 G
#438640000000
0!
1"
0*
1+
09
1:
0>
0C
#438650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#438660000000
0!
0*
09
0>
0C
#438670000000
1!
1*
b1 6
19
1>
1C
b1 G
#438680000000
0!
0*
09
0>
0C
#438690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#438700000000
0!
0*
09
0>
0C
#438710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#438720000000
0!
0*
09
0>
0C
#438730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#438740000000
0!
0*
09
0>
0C
#438750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#438760000000
0!
0#
0*
0,
09
0>
0?
0C
#438770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#438780000000
0!
0*
09
0>
0C
#438790000000
1!
1*
19
1>
1C
#438800000000
0!
0*
09
0>
0C
#438810000000
1!
1*
19
1>
1C
#438820000000
0!
0*
09
0>
0C
#438830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#438840000000
0!
0*
09
0>
0C
#438850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#438860000000
0!
0*
09
0>
0C
#438870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#438880000000
0!
0*
09
0>
0C
#438890000000
1!
1*
b10 6
19
1>
1C
b10 G
#438900000000
0!
0*
09
0>
0C
#438910000000
1!
1*
b11 6
19
1>
1C
b11 G
#438920000000
0!
0*
09
0>
0C
#438930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#438940000000
0!
0*
09
0>
0C
#438950000000
1!
1*
b101 6
19
1>
1C
b101 G
#438960000000
0!
0*
09
0>
0C
#438970000000
1!
1*
b110 6
19
1>
1C
b110 G
#438980000000
0!
0*
09
0>
0C
#438990000000
1!
1*
b111 6
19
1>
1C
b111 G
#439000000000
0!
0*
09
0>
0C
#439010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#439020000000
0!
0*
09
0>
0C
#439030000000
1!
1*
b1 6
19
1>
1C
b1 G
#439040000000
0!
0*
09
0>
0C
#439050000000
1!
1*
b10 6
19
1>
1C
b10 G
#439060000000
0!
0*
09
0>
0C
#439070000000
1!
1*
b11 6
19
1>
1C
b11 G
#439080000000
0!
0*
09
0>
0C
#439090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#439100000000
0!
0*
09
0>
0C
#439110000000
1!
1*
b101 6
19
1>
1C
b101 G
#439120000000
0!
0*
09
0>
0C
#439130000000
1!
1*
b110 6
19
1>
1C
b110 G
#439140000000
0!
0*
09
0>
0C
#439150000000
1!
1*
b111 6
19
1>
1C
b111 G
#439160000000
0!
0*
09
0>
0C
#439170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#439180000000
0!
0*
09
0>
0C
#439190000000
1!
1*
b1 6
19
1>
1C
b1 G
#439200000000
0!
0*
09
0>
0C
#439210000000
1!
1*
b10 6
19
1>
1C
b10 G
#439220000000
0!
0*
09
0>
0C
#439230000000
1!
1*
b11 6
19
1>
1C
b11 G
#439240000000
0!
0*
09
0>
0C
#439250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#439260000000
0!
0*
09
0>
0C
#439270000000
1!
1*
b101 6
19
1>
1C
b101 G
#439280000000
0!
0*
09
0>
0C
#439290000000
1!
1*
b110 6
19
1>
1C
b110 G
#439300000000
0!
0*
09
0>
0C
#439310000000
1!
1*
b111 6
19
1>
1C
b111 G
#439320000000
0!
1"
0*
1+
09
1:
0>
0C
#439330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#439340000000
0!
0*
09
0>
0C
#439350000000
1!
1*
b1 6
19
1>
1C
b1 G
#439360000000
0!
0*
09
0>
0C
#439370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#439380000000
0!
0*
09
0>
0C
#439390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#439400000000
0!
0*
09
0>
0C
#439410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#439420000000
0!
0*
09
0>
0C
#439430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#439440000000
0!
0#
0*
0,
09
0>
0?
0C
#439450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#439460000000
0!
0*
09
0>
0C
#439470000000
1!
1*
19
1>
1C
#439480000000
0!
0*
09
0>
0C
#439490000000
1!
1*
19
1>
1C
#439500000000
0!
0*
09
0>
0C
#439510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#439520000000
0!
0*
09
0>
0C
#439530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#439540000000
0!
0*
09
0>
0C
#439550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#439560000000
0!
0*
09
0>
0C
#439570000000
1!
1*
b10 6
19
1>
1C
b10 G
#439580000000
0!
0*
09
0>
0C
#439590000000
1!
1*
b11 6
19
1>
1C
b11 G
#439600000000
0!
0*
09
0>
0C
#439610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#439620000000
0!
0*
09
0>
0C
#439630000000
1!
1*
b101 6
19
1>
1C
b101 G
#439640000000
0!
0*
09
0>
0C
#439650000000
1!
1*
b110 6
19
1>
1C
b110 G
#439660000000
0!
0*
09
0>
0C
#439670000000
1!
1*
b111 6
19
1>
1C
b111 G
#439680000000
0!
0*
09
0>
0C
#439690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#439700000000
0!
0*
09
0>
0C
#439710000000
1!
1*
b1 6
19
1>
1C
b1 G
#439720000000
0!
0*
09
0>
0C
#439730000000
1!
1*
b10 6
19
1>
1C
b10 G
#439740000000
0!
0*
09
0>
0C
#439750000000
1!
1*
b11 6
19
1>
1C
b11 G
#439760000000
0!
0*
09
0>
0C
#439770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#439780000000
0!
0*
09
0>
0C
#439790000000
1!
1*
b101 6
19
1>
1C
b101 G
#439800000000
0!
0*
09
0>
0C
#439810000000
1!
1*
b110 6
19
1>
1C
b110 G
#439820000000
0!
0*
09
0>
0C
#439830000000
1!
1*
b111 6
19
1>
1C
b111 G
#439840000000
0!
0*
09
0>
0C
#439850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#439860000000
0!
0*
09
0>
0C
#439870000000
1!
1*
b1 6
19
1>
1C
b1 G
#439880000000
0!
0*
09
0>
0C
#439890000000
1!
1*
b10 6
19
1>
1C
b10 G
#439900000000
0!
0*
09
0>
0C
#439910000000
1!
1*
b11 6
19
1>
1C
b11 G
#439920000000
0!
0*
09
0>
0C
#439930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#439940000000
0!
0*
09
0>
0C
#439950000000
1!
1*
b101 6
19
1>
1C
b101 G
#439960000000
0!
0*
09
0>
0C
#439970000000
1!
1*
b110 6
19
1>
1C
b110 G
#439980000000
0!
0*
09
0>
0C
#439990000000
1!
1*
b111 6
19
1>
1C
b111 G
#440000000000
0!
1"
0*
1+
09
1:
0>
0C
#440010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#440020000000
0!
0*
09
0>
0C
#440030000000
1!
1*
b1 6
19
1>
1C
b1 G
#440040000000
0!
0*
09
0>
0C
#440050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#440060000000
0!
0*
09
0>
0C
#440070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#440080000000
0!
0*
09
0>
0C
#440090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#440100000000
0!
0*
09
0>
0C
#440110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#440120000000
0!
0#
0*
0,
09
0>
0?
0C
#440130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#440140000000
0!
0*
09
0>
0C
#440150000000
1!
1*
19
1>
1C
#440160000000
0!
0*
09
0>
0C
#440170000000
1!
1*
19
1>
1C
#440180000000
0!
0*
09
0>
0C
#440190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#440200000000
0!
0*
09
0>
0C
#440210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#440220000000
0!
0*
09
0>
0C
#440230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#440240000000
0!
0*
09
0>
0C
#440250000000
1!
1*
b10 6
19
1>
1C
b10 G
#440260000000
0!
0*
09
0>
0C
#440270000000
1!
1*
b11 6
19
1>
1C
b11 G
#440280000000
0!
0*
09
0>
0C
#440290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#440300000000
0!
0*
09
0>
0C
#440310000000
1!
1*
b101 6
19
1>
1C
b101 G
#440320000000
0!
0*
09
0>
0C
#440330000000
1!
1*
b110 6
19
1>
1C
b110 G
#440340000000
0!
0*
09
0>
0C
#440350000000
1!
1*
b111 6
19
1>
1C
b111 G
#440360000000
0!
0*
09
0>
0C
#440370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#440380000000
0!
0*
09
0>
0C
#440390000000
1!
1*
b1 6
19
1>
1C
b1 G
#440400000000
0!
0*
09
0>
0C
#440410000000
1!
1*
b10 6
19
1>
1C
b10 G
#440420000000
0!
0*
09
0>
0C
#440430000000
1!
1*
b11 6
19
1>
1C
b11 G
#440440000000
0!
0*
09
0>
0C
#440450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#440460000000
0!
0*
09
0>
0C
#440470000000
1!
1*
b101 6
19
1>
1C
b101 G
#440480000000
0!
0*
09
0>
0C
#440490000000
1!
1*
b110 6
19
1>
1C
b110 G
#440500000000
0!
0*
09
0>
0C
#440510000000
1!
1*
b111 6
19
1>
1C
b111 G
#440520000000
0!
0*
09
0>
0C
#440530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#440540000000
0!
0*
09
0>
0C
#440550000000
1!
1*
b1 6
19
1>
1C
b1 G
#440560000000
0!
0*
09
0>
0C
#440570000000
1!
1*
b10 6
19
1>
1C
b10 G
#440580000000
0!
0*
09
0>
0C
#440590000000
1!
1*
b11 6
19
1>
1C
b11 G
#440600000000
0!
0*
09
0>
0C
#440610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#440620000000
0!
0*
09
0>
0C
#440630000000
1!
1*
b101 6
19
1>
1C
b101 G
#440640000000
0!
0*
09
0>
0C
#440650000000
1!
1*
b110 6
19
1>
1C
b110 G
#440660000000
0!
0*
09
0>
0C
#440670000000
1!
1*
b111 6
19
1>
1C
b111 G
#440680000000
0!
1"
0*
1+
09
1:
0>
0C
#440690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#440700000000
0!
0*
09
0>
0C
#440710000000
1!
1*
b1 6
19
1>
1C
b1 G
#440720000000
0!
0*
09
0>
0C
#440730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#440740000000
0!
0*
09
0>
0C
#440750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#440760000000
0!
0*
09
0>
0C
#440770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#440780000000
0!
0*
09
0>
0C
#440790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#440800000000
0!
0#
0*
0,
09
0>
0?
0C
#440810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#440820000000
0!
0*
09
0>
0C
#440830000000
1!
1*
19
1>
1C
#440840000000
0!
0*
09
0>
0C
#440850000000
1!
1*
19
1>
1C
#440860000000
0!
0*
09
0>
0C
#440870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#440880000000
0!
0*
09
0>
0C
#440890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#440900000000
0!
0*
09
0>
0C
#440910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#440920000000
0!
0*
09
0>
0C
#440930000000
1!
1*
b10 6
19
1>
1C
b10 G
#440940000000
0!
0*
09
0>
0C
#440950000000
1!
1*
b11 6
19
1>
1C
b11 G
#440960000000
0!
0*
09
0>
0C
#440970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#440980000000
0!
0*
09
0>
0C
#440990000000
1!
1*
b101 6
19
1>
1C
b101 G
#441000000000
0!
0*
09
0>
0C
#441010000000
1!
1*
b110 6
19
1>
1C
b110 G
#441020000000
0!
0*
09
0>
0C
#441030000000
1!
1*
b111 6
19
1>
1C
b111 G
#441040000000
0!
0*
09
0>
0C
#441050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#441060000000
0!
0*
09
0>
0C
#441070000000
1!
1*
b1 6
19
1>
1C
b1 G
#441080000000
0!
0*
09
0>
0C
#441090000000
1!
1*
b10 6
19
1>
1C
b10 G
#441100000000
0!
0*
09
0>
0C
#441110000000
1!
1*
b11 6
19
1>
1C
b11 G
#441120000000
0!
0*
09
0>
0C
#441130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#441140000000
0!
0*
09
0>
0C
#441150000000
1!
1*
b101 6
19
1>
1C
b101 G
#441160000000
0!
0*
09
0>
0C
#441170000000
1!
1*
b110 6
19
1>
1C
b110 G
#441180000000
0!
0*
09
0>
0C
#441190000000
1!
1*
b111 6
19
1>
1C
b111 G
#441200000000
0!
0*
09
0>
0C
#441210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#441220000000
0!
0*
09
0>
0C
#441230000000
1!
1*
b1 6
19
1>
1C
b1 G
#441240000000
0!
0*
09
0>
0C
#441250000000
1!
1*
b10 6
19
1>
1C
b10 G
#441260000000
0!
0*
09
0>
0C
#441270000000
1!
1*
b11 6
19
1>
1C
b11 G
#441280000000
0!
0*
09
0>
0C
#441290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#441300000000
0!
0*
09
0>
0C
#441310000000
1!
1*
b101 6
19
1>
1C
b101 G
#441320000000
0!
0*
09
0>
0C
#441330000000
1!
1*
b110 6
19
1>
1C
b110 G
#441340000000
0!
0*
09
0>
0C
#441350000000
1!
1*
b111 6
19
1>
1C
b111 G
#441360000000
0!
1"
0*
1+
09
1:
0>
0C
#441370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#441380000000
0!
0*
09
0>
0C
#441390000000
1!
1*
b1 6
19
1>
1C
b1 G
#441400000000
0!
0*
09
0>
0C
#441410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#441420000000
0!
0*
09
0>
0C
#441430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#441440000000
0!
0*
09
0>
0C
#441450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#441460000000
0!
0*
09
0>
0C
#441470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#441480000000
0!
0#
0*
0,
09
0>
0?
0C
#441490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#441500000000
0!
0*
09
0>
0C
#441510000000
1!
1*
19
1>
1C
#441520000000
0!
0*
09
0>
0C
#441530000000
1!
1*
19
1>
1C
#441540000000
0!
0*
09
0>
0C
#441550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#441560000000
0!
0*
09
0>
0C
#441570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#441580000000
0!
0*
09
0>
0C
#441590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#441600000000
0!
0*
09
0>
0C
#441610000000
1!
1*
b10 6
19
1>
1C
b10 G
#441620000000
0!
0*
09
0>
0C
#441630000000
1!
1*
b11 6
19
1>
1C
b11 G
#441640000000
0!
0*
09
0>
0C
#441650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#441660000000
0!
0*
09
0>
0C
#441670000000
1!
1*
b101 6
19
1>
1C
b101 G
#441680000000
0!
0*
09
0>
0C
#441690000000
1!
1*
b110 6
19
1>
1C
b110 G
#441700000000
0!
0*
09
0>
0C
#441710000000
1!
1*
b111 6
19
1>
1C
b111 G
#441720000000
0!
0*
09
0>
0C
#441730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#441740000000
0!
0*
09
0>
0C
#441750000000
1!
1*
b1 6
19
1>
1C
b1 G
#441760000000
0!
0*
09
0>
0C
#441770000000
1!
1*
b10 6
19
1>
1C
b10 G
#441780000000
0!
0*
09
0>
0C
#441790000000
1!
1*
b11 6
19
1>
1C
b11 G
#441800000000
0!
0*
09
0>
0C
#441810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#441820000000
0!
0*
09
0>
0C
#441830000000
1!
1*
b101 6
19
1>
1C
b101 G
#441840000000
0!
0*
09
0>
0C
#441850000000
1!
1*
b110 6
19
1>
1C
b110 G
#441860000000
0!
0*
09
0>
0C
#441870000000
1!
1*
b111 6
19
1>
1C
b111 G
#441880000000
0!
0*
09
0>
0C
#441890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#441900000000
0!
0*
09
0>
0C
#441910000000
1!
1*
b1 6
19
1>
1C
b1 G
#441920000000
0!
0*
09
0>
0C
#441930000000
1!
1*
b10 6
19
1>
1C
b10 G
#441940000000
0!
0*
09
0>
0C
#441950000000
1!
1*
b11 6
19
1>
1C
b11 G
#441960000000
0!
0*
09
0>
0C
#441970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#441980000000
0!
0*
09
0>
0C
#441990000000
1!
1*
b101 6
19
1>
1C
b101 G
#442000000000
0!
0*
09
0>
0C
#442010000000
1!
1*
b110 6
19
1>
1C
b110 G
#442020000000
0!
0*
09
0>
0C
#442030000000
1!
1*
b111 6
19
1>
1C
b111 G
#442040000000
0!
1"
0*
1+
09
1:
0>
0C
#442050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#442060000000
0!
0*
09
0>
0C
#442070000000
1!
1*
b1 6
19
1>
1C
b1 G
#442080000000
0!
0*
09
0>
0C
#442090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#442100000000
0!
0*
09
0>
0C
#442110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#442120000000
0!
0*
09
0>
0C
#442130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#442140000000
0!
0*
09
0>
0C
#442150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#442160000000
0!
0#
0*
0,
09
0>
0?
0C
#442170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#442180000000
0!
0*
09
0>
0C
#442190000000
1!
1*
19
1>
1C
#442200000000
0!
0*
09
0>
0C
#442210000000
1!
1*
19
1>
1C
#442220000000
0!
0*
09
0>
0C
#442230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#442240000000
0!
0*
09
0>
0C
#442250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#442260000000
0!
0*
09
0>
0C
#442270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#442280000000
0!
0*
09
0>
0C
#442290000000
1!
1*
b10 6
19
1>
1C
b10 G
#442300000000
0!
0*
09
0>
0C
#442310000000
1!
1*
b11 6
19
1>
1C
b11 G
#442320000000
0!
0*
09
0>
0C
#442330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#442340000000
0!
0*
09
0>
0C
#442350000000
1!
1*
b101 6
19
1>
1C
b101 G
#442360000000
0!
0*
09
0>
0C
#442370000000
1!
1*
b110 6
19
1>
1C
b110 G
#442380000000
0!
0*
09
0>
0C
#442390000000
1!
1*
b111 6
19
1>
1C
b111 G
#442400000000
0!
0*
09
0>
0C
#442410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#442420000000
0!
0*
09
0>
0C
#442430000000
1!
1*
b1 6
19
1>
1C
b1 G
#442440000000
0!
0*
09
0>
0C
#442450000000
1!
1*
b10 6
19
1>
1C
b10 G
#442460000000
0!
0*
09
0>
0C
#442470000000
1!
1*
b11 6
19
1>
1C
b11 G
#442480000000
0!
0*
09
0>
0C
#442490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#442500000000
0!
0*
09
0>
0C
#442510000000
1!
1*
b101 6
19
1>
1C
b101 G
#442520000000
0!
0*
09
0>
0C
#442530000000
1!
1*
b110 6
19
1>
1C
b110 G
#442540000000
0!
0*
09
0>
0C
#442550000000
1!
1*
b111 6
19
1>
1C
b111 G
#442560000000
0!
0*
09
0>
0C
#442570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#442580000000
0!
0*
09
0>
0C
#442590000000
1!
1*
b1 6
19
1>
1C
b1 G
#442600000000
0!
0*
09
0>
0C
#442610000000
1!
1*
b10 6
19
1>
1C
b10 G
#442620000000
0!
0*
09
0>
0C
#442630000000
1!
1*
b11 6
19
1>
1C
b11 G
#442640000000
0!
0*
09
0>
0C
#442650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#442660000000
0!
0*
09
0>
0C
#442670000000
1!
1*
b101 6
19
1>
1C
b101 G
#442680000000
0!
0*
09
0>
0C
#442690000000
1!
1*
b110 6
19
1>
1C
b110 G
#442700000000
0!
0*
09
0>
0C
#442710000000
1!
1*
b111 6
19
1>
1C
b111 G
#442720000000
0!
1"
0*
1+
09
1:
0>
0C
#442730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#442740000000
0!
0*
09
0>
0C
#442750000000
1!
1*
b1 6
19
1>
1C
b1 G
#442760000000
0!
0*
09
0>
0C
#442770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#442780000000
0!
0*
09
0>
0C
#442790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#442800000000
0!
0*
09
0>
0C
#442810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#442820000000
0!
0*
09
0>
0C
#442830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#442840000000
0!
0#
0*
0,
09
0>
0?
0C
#442850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#442860000000
0!
0*
09
0>
0C
#442870000000
1!
1*
19
1>
1C
#442880000000
0!
0*
09
0>
0C
#442890000000
1!
1*
19
1>
1C
#442900000000
0!
0*
09
0>
0C
#442910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#442920000000
0!
0*
09
0>
0C
#442930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#442940000000
0!
0*
09
0>
0C
#442950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#442960000000
0!
0*
09
0>
0C
#442970000000
1!
1*
b10 6
19
1>
1C
b10 G
#442980000000
0!
0*
09
0>
0C
#442990000000
1!
1*
b11 6
19
1>
1C
b11 G
#443000000000
0!
0*
09
0>
0C
#443010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#443020000000
0!
0*
09
0>
0C
#443030000000
1!
1*
b101 6
19
1>
1C
b101 G
#443040000000
0!
0*
09
0>
0C
#443050000000
1!
1*
b110 6
19
1>
1C
b110 G
#443060000000
0!
0*
09
0>
0C
#443070000000
1!
1*
b111 6
19
1>
1C
b111 G
#443080000000
0!
0*
09
0>
0C
#443090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#443100000000
0!
0*
09
0>
0C
#443110000000
1!
1*
b1 6
19
1>
1C
b1 G
#443120000000
0!
0*
09
0>
0C
#443130000000
1!
1*
b10 6
19
1>
1C
b10 G
#443140000000
0!
0*
09
0>
0C
#443150000000
1!
1*
b11 6
19
1>
1C
b11 G
#443160000000
0!
0*
09
0>
0C
#443170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#443180000000
0!
0*
09
0>
0C
#443190000000
1!
1*
b101 6
19
1>
1C
b101 G
#443200000000
0!
0*
09
0>
0C
#443210000000
1!
1*
b110 6
19
1>
1C
b110 G
#443220000000
0!
0*
09
0>
0C
#443230000000
1!
1*
b111 6
19
1>
1C
b111 G
#443240000000
0!
0*
09
0>
0C
#443250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#443260000000
0!
0*
09
0>
0C
#443270000000
1!
1*
b1 6
19
1>
1C
b1 G
#443280000000
0!
0*
09
0>
0C
#443290000000
1!
1*
b10 6
19
1>
1C
b10 G
#443300000000
0!
0*
09
0>
0C
#443310000000
1!
1*
b11 6
19
1>
1C
b11 G
#443320000000
0!
0*
09
0>
0C
#443330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#443340000000
0!
0*
09
0>
0C
#443350000000
1!
1*
b101 6
19
1>
1C
b101 G
#443360000000
0!
0*
09
0>
0C
#443370000000
1!
1*
b110 6
19
1>
1C
b110 G
#443380000000
0!
0*
09
0>
0C
#443390000000
1!
1*
b111 6
19
1>
1C
b111 G
#443400000000
0!
1"
0*
1+
09
1:
0>
0C
#443410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#443420000000
0!
0*
09
0>
0C
#443430000000
1!
1*
b1 6
19
1>
1C
b1 G
#443440000000
0!
0*
09
0>
0C
#443450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#443460000000
0!
0*
09
0>
0C
#443470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#443480000000
0!
0*
09
0>
0C
#443490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#443500000000
0!
0*
09
0>
0C
#443510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#443520000000
0!
0#
0*
0,
09
0>
0?
0C
#443530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#443540000000
0!
0*
09
0>
0C
#443550000000
1!
1*
19
1>
1C
#443560000000
0!
0*
09
0>
0C
#443570000000
1!
1*
19
1>
1C
#443580000000
0!
0*
09
0>
0C
#443590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#443600000000
0!
0*
09
0>
0C
#443610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#443620000000
0!
0*
09
0>
0C
#443630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#443640000000
0!
0*
09
0>
0C
#443650000000
1!
1*
b10 6
19
1>
1C
b10 G
#443660000000
0!
0*
09
0>
0C
#443670000000
1!
1*
b11 6
19
1>
1C
b11 G
#443680000000
0!
0*
09
0>
0C
#443690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#443700000000
0!
0*
09
0>
0C
#443710000000
1!
1*
b101 6
19
1>
1C
b101 G
#443720000000
0!
0*
09
0>
0C
#443730000000
1!
1*
b110 6
19
1>
1C
b110 G
#443740000000
0!
0*
09
0>
0C
#443750000000
1!
1*
b111 6
19
1>
1C
b111 G
#443760000000
0!
0*
09
0>
0C
#443770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#443780000000
0!
0*
09
0>
0C
#443790000000
1!
1*
b1 6
19
1>
1C
b1 G
#443800000000
0!
0*
09
0>
0C
#443810000000
1!
1*
b10 6
19
1>
1C
b10 G
#443820000000
0!
0*
09
0>
0C
#443830000000
1!
1*
b11 6
19
1>
1C
b11 G
#443840000000
0!
0*
09
0>
0C
#443850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#443860000000
0!
0*
09
0>
0C
#443870000000
1!
1*
b101 6
19
1>
1C
b101 G
#443880000000
0!
0*
09
0>
0C
#443890000000
1!
1*
b110 6
19
1>
1C
b110 G
#443900000000
0!
0*
09
0>
0C
#443910000000
1!
1*
b111 6
19
1>
1C
b111 G
#443920000000
0!
0*
09
0>
0C
#443930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#443940000000
0!
0*
09
0>
0C
#443950000000
1!
1*
b1 6
19
1>
1C
b1 G
#443960000000
0!
0*
09
0>
0C
#443970000000
1!
1*
b10 6
19
1>
1C
b10 G
#443980000000
0!
0*
09
0>
0C
#443990000000
1!
1*
b11 6
19
1>
1C
b11 G
#444000000000
0!
0*
09
0>
0C
#444010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#444020000000
0!
0*
09
0>
0C
#444030000000
1!
1*
b101 6
19
1>
1C
b101 G
#444040000000
0!
0*
09
0>
0C
#444050000000
1!
1*
b110 6
19
1>
1C
b110 G
#444060000000
0!
0*
09
0>
0C
#444070000000
1!
1*
b111 6
19
1>
1C
b111 G
#444080000000
0!
1"
0*
1+
09
1:
0>
0C
#444090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#444100000000
0!
0*
09
0>
0C
#444110000000
1!
1*
b1 6
19
1>
1C
b1 G
#444120000000
0!
0*
09
0>
0C
#444130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#444140000000
0!
0*
09
0>
0C
#444150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#444160000000
0!
0*
09
0>
0C
#444170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#444180000000
0!
0*
09
0>
0C
#444190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#444200000000
0!
0#
0*
0,
09
0>
0?
0C
#444210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#444220000000
0!
0*
09
0>
0C
#444230000000
1!
1*
19
1>
1C
#444240000000
0!
0*
09
0>
0C
#444250000000
1!
1*
19
1>
1C
#444260000000
0!
0*
09
0>
0C
#444270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#444280000000
0!
0*
09
0>
0C
#444290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#444300000000
0!
0*
09
0>
0C
#444310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#444320000000
0!
0*
09
0>
0C
#444330000000
1!
1*
b10 6
19
1>
1C
b10 G
#444340000000
0!
0*
09
0>
0C
#444350000000
1!
1*
b11 6
19
1>
1C
b11 G
#444360000000
0!
0*
09
0>
0C
#444370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#444380000000
0!
0*
09
0>
0C
#444390000000
1!
1*
b101 6
19
1>
1C
b101 G
#444400000000
0!
0*
09
0>
0C
#444410000000
1!
1*
b110 6
19
1>
1C
b110 G
#444420000000
0!
0*
09
0>
0C
#444430000000
1!
1*
b111 6
19
1>
1C
b111 G
#444440000000
0!
0*
09
0>
0C
#444450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#444460000000
0!
0*
09
0>
0C
#444470000000
1!
1*
b1 6
19
1>
1C
b1 G
#444480000000
0!
0*
09
0>
0C
#444490000000
1!
1*
b10 6
19
1>
1C
b10 G
#444500000000
0!
0*
09
0>
0C
#444510000000
1!
1*
b11 6
19
1>
1C
b11 G
#444520000000
0!
0*
09
0>
0C
#444530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#444540000000
0!
0*
09
0>
0C
#444550000000
1!
1*
b101 6
19
1>
1C
b101 G
#444560000000
0!
0*
09
0>
0C
#444570000000
1!
1*
b110 6
19
1>
1C
b110 G
#444580000000
0!
0*
09
0>
0C
#444590000000
1!
1*
b111 6
19
1>
1C
b111 G
#444600000000
0!
0*
09
0>
0C
#444610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#444620000000
0!
0*
09
0>
0C
#444630000000
1!
1*
b1 6
19
1>
1C
b1 G
#444640000000
0!
0*
09
0>
0C
#444650000000
1!
1*
b10 6
19
1>
1C
b10 G
#444660000000
0!
0*
09
0>
0C
#444670000000
1!
1*
b11 6
19
1>
1C
b11 G
#444680000000
0!
0*
09
0>
0C
#444690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#444700000000
0!
0*
09
0>
0C
#444710000000
1!
1*
b101 6
19
1>
1C
b101 G
#444720000000
0!
0*
09
0>
0C
#444730000000
1!
1*
b110 6
19
1>
1C
b110 G
#444740000000
0!
0*
09
0>
0C
#444750000000
1!
1*
b111 6
19
1>
1C
b111 G
#444760000000
0!
1"
0*
1+
09
1:
0>
0C
#444770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#444780000000
0!
0*
09
0>
0C
#444790000000
1!
1*
b1 6
19
1>
1C
b1 G
#444800000000
0!
0*
09
0>
0C
#444810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#444820000000
0!
0*
09
0>
0C
#444830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#444840000000
0!
0*
09
0>
0C
#444850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#444860000000
0!
0*
09
0>
0C
#444870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#444880000000
0!
0#
0*
0,
09
0>
0?
0C
#444890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#444900000000
0!
0*
09
0>
0C
#444910000000
1!
1*
19
1>
1C
#444920000000
0!
0*
09
0>
0C
#444930000000
1!
1*
19
1>
1C
#444940000000
0!
0*
09
0>
0C
#444950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#444960000000
0!
0*
09
0>
0C
#444970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#444980000000
0!
0*
09
0>
0C
#444990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#445000000000
0!
0*
09
0>
0C
#445010000000
1!
1*
b10 6
19
1>
1C
b10 G
#445020000000
0!
0*
09
0>
0C
#445030000000
1!
1*
b11 6
19
1>
1C
b11 G
#445040000000
0!
0*
09
0>
0C
#445050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#445060000000
0!
0*
09
0>
0C
#445070000000
1!
1*
b101 6
19
1>
1C
b101 G
#445080000000
0!
0*
09
0>
0C
#445090000000
1!
1*
b110 6
19
1>
1C
b110 G
#445100000000
0!
0*
09
0>
0C
#445110000000
1!
1*
b111 6
19
1>
1C
b111 G
#445120000000
0!
0*
09
0>
0C
#445130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#445140000000
0!
0*
09
0>
0C
#445150000000
1!
1*
b1 6
19
1>
1C
b1 G
#445160000000
0!
0*
09
0>
0C
#445170000000
1!
1*
b10 6
19
1>
1C
b10 G
#445180000000
0!
0*
09
0>
0C
#445190000000
1!
1*
b11 6
19
1>
1C
b11 G
#445200000000
0!
0*
09
0>
0C
#445210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#445220000000
0!
0*
09
0>
0C
#445230000000
1!
1*
b101 6
19
1>
1C
b101 G
#445240000000
0!
0*
09
0>
0C
#445250000000
1!
1*
b110 6
19
1>
1C
b110 G
#445260000000
0!
0*
09
0>
0C
#445270000000
1!
1*
b111 6
19
1>
1C
b111 G
#445280000000
0!
0*
09
0>
0C
#445290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#445300000000
0!
0*
09
0>
0C
#445310000000
1!
1*
b1 6
19
1>
1C
b1 G
#445320000000
0!
0*
09
0>
0C
#445330000000
1!
1*
b10 6
19
1>
1C
b10 G
#445340000000
0!
0*
09
0>
0C
#445350000000
1!
1*
b11 6
19
1>
1C
b11 G
#445360000000
0!
0*
09
0>
0C
#445370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#445380000000
0!
0*
09
0>
0C
#445390000000
1!
1*
b101 6
19
1>
1C
b101 G
#445400000000
0!
0*
09
0>
0C
#445410000000
1!
1*
b110 6
19
1>
1C
b110 G
#445420000000
0!
0*
09
0>
0C
#445430000000
1!
1*
b111 6
19
1>
1C
b111 G
#445440000000
0!
1"
0*
1+
09
1:
0>
0C
#445450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#445460000000
0!
0*
09
0>
0C
#445470000000
1!
1*
b1 6
19
1>
1C
b1 G
#445480000000
0!
0*
09
0>
0C
#445490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#445500000000
0!
0*
09
0>
0C
#445510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#445520000000
0!
0*
09
0>
0C
#445530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#445540000000
0!
0*
09
0>
0C
#445550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#445560000000
0!
0#
0*
0,
09
0>
0?
0C
#445570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#445580000000
0!
0*
09
0>
0C
#445590000000
1!
1*
19
1>
1C
#445600000000
0!
0*
09
0>
0C
#445610000000
1!
1*
19
1>
1C
#445620000000
0!
0*
09
0>
0C
#445630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#445640000000
0!
0*
09
0>
0C
#445650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#445660000000
0!
0*
09
0>
0C
#445670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#445680000000
0!
0*
09
0>
0C
#445690000000
1!
1*
b10 6
19
1>
1C
b10 G
#445700000000
0!
0*
09
0>
0C
#445710000000
1!
1*
b11 6
19
1>
1C
b11 G
#445720000000
0!
0*
09
0>
0C
#445730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#445740000000
0!
0*
09
0>
0C
#445750000000
1!
1*
b101 6
19
1>
1C
b101 G
#445760000000
0!
0*
09
0>
0C
#445770000000
1!
1*
b110 6
19
1>
1C
b110 G
#445780000000
0!
0*
09
0>
0C
#445790000000
1!
1*
b111 6
19
1>
1C
b111 G
#445800000000
0!
0*
09
0>
0C
#445810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#445820000000
0!
0*
09
0>
0C
#445830000000
1!
1*
b1 6
19
1>
1C
b1 G
#445840000000
0!
0*
09
0>
0C
#445850000000
1!
1*
b10 6
19
1>
1C
b10 G
#445860000000
0!
0*
09
0>
0C
#445870000000
1!
1*
b11 6
19
1>
1C
b11 G
#445880000000
0!
0*
09
0>
0C
#445890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#445900000000
0!
0*
09
0>
0C
#445910000000
1!
1*
b101 6
19
1>
1C
b101 G
#445920000000
0!
0*
09
0>
0C
#445930000000
1!
1*
b110 6
19
1>
1C
b110 G
#445940000000
0!
0*
09
0>
0C
#445950000000
1!
1*
b111 6
19
1>
1C
b111 G
#445960000000
0!
0*
09
0>
0C
#445970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#445980000000
0!
0*
09
0>
0C
#445990000000
1!
1*
b1 6
19
1>
1C
b1 G
#446000000000
0!
0*
09
0>
0C
#446010000000
1!
1*
b10 6
19
1>
1C
b10 G
#446020000000
0!
0*
09
0>
0C
#446030000000
1!
1*
b11 6
19
1>
1C
b11 G
#446040000000
0!
0*
09
0>
0C
#446050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#446060000000
0!
0*
09
0>
0C
#446070000000
1!
1*
b101 6
19
1>
1C
b101 G
#446080000000
0!
0*
09
0>
0C
#446090000000
1!
1*
b110 6
19
1>
1C
b110 G
#446100000000
0!
0*
09
0>
0C
#446110000000
1!
1*
b111 6
19
1>
1C
b111 G
#446120000000
0!
1"
0*
1+
09
1:
0>
0C
#446130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#446140000000
0!
0*
09
0>
0C
#446150000000
1!
1*
b1 6
19
1>
1C
b1 G
#446160000000
0!
0*
09
0>
0C
#446170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#446180000000
0!
0*
09
0>
0C
#446190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#446200000000
0!
0*
09
0>
0C
#446210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#446220000000
0!
0*
09
0>
0C
#446230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#446240000000
0!
0#
0*
0,
09
0>
0?
0C
#446250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#446260000000
0!
0*
09
0>
0C
#446270000000
1!
1*
19
1>
1C
#446280000000
0!
0*
09
0>
0C
#446290000000
1!
1*
19
1>
1C
#446300000000
0!
0*
09
0>
0C
#446310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#446320000000
0!
0*
09
0>
0C
#446330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#446340000000
0!
0*
09
0>
0C
#446350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#446360000000
0!
0*
09
0>
0C
#446370000000
1!
1*
b10 6
19
1>
1C
b10 G
#446380000000
0!
0*
09
0>
0C
#446390000000
1!
1*
b11 6
19
1>
1C
b11 G
#446400000000
0!
0*
09
0>
0C
#446410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#446420000000
0!
0*
09
0>
0C
#446430000000
1!
1*
b101 6
19
1>
1C
b101 G
#446440000000
0!
0*
09
0>
0C
#446450000000
1!
1*
b110 6
19
1>
1C
b110 G
#446460000000
0!
0*
09
0>
0C
#446470000000
1!
1*
b111 6
19
1>
1C
b111 G
#446480000000
0!
0*
09
0>
0C
#446490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#446500000000
0!
0*
09
0>
0C
#446510000000
1!
1*
b1 6
19
1>
1C
b1 G
#446520000000
0!
0*
09
0>
0C
#446530000000
1!
1*
b10 6
19
1>
1C
b10 G
#446540000000
0!
0*
09
0>
0C
#446550000000
1!
1*
b11 6
19
1>
1C
b11 G
#446560000000
0!
0*
09
0>
0C
#446570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#446580000000
0!
0*
09
0>
0C
#446590000000
1!
1*
b101 6
19
1>
1C
b101 G
#446600000000
0!
0*
09
0>
0C
#446610000000
1!
1*
b110 6
19
1>
1C
b110 G
#446620000000
0!
0*
09
0>
0C
#446630000000
1!
1*
b111 6
19
1>
1C
b111 G
#446640000000
0!
0*
09
0>
0C
#446650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#446660000000
0!
0*
09
0>
0C
#446670000000
1!
1*
b1 6
19
1>
1C
b1 G
#446680000000
0!
0*
09
0>
0C
#446690000000
1!
1*
b10 6
19
1>
1C
b10 G
#446700000000
0!
0*
09
0>
0C
#446710000000
1!
1*
b11 6
19
1>
1C
b11 G
#446720000000
0!
0*
09
0>
0C
#446730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#446740000000
0!
0*
09
0>
0C
#446750000000
1!
1*
b101 6
19
1>
1C
b101 G
#446760000000
0!
0*
09
0>
0C
#446770000000
1!
1*
b110 6
19
1>
1C
b110 G
#446780000000
0!
0*
09
0>
0C
#446790000000
1!
1*
b111 6
19
1>
1C
b111 G
#446800000000
0!
1"
0*
1+
09
1:
0>
0C
#446810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#446820000000
0!
0*
09
0>
0C
#446830000000
1!
1*
b1 6
19
1>
1C
b1 G
#446840000000
0!
0*
09
0>
0C
#446850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#446860000000
0!
0*
09
0>
0C
#446870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#446880000000
0!
0*
09
0>
0C
#446890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#446900000000
0!
0*
09
0>
0C
#446910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#446920000000
0!
0#
0*
0,
09
0>
0?
0C
#446930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#446940000000
0!
0*
09
0>
0C
#446950000000
1!
1*
19
1>
1C
#446960000000
0!
0*
09
0>
0C
#446970000000
1!
1*
19
1>
1C
#446980000000
0!
0*
09
0>
0C
#446990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#447000000000
0!
0*
09
0>
0C
#447010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#447020000000
0!
0*
09
0>
0C
#447030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#447040000000
0!
0*
09
0>
0C
#447050000000
1!
1*
b10 6
19
1>
1C
b10 G
#447060000000
0!
0*
09
0>
0C
#447070000000
1!
1*
b11 6
19
1>
1C
b11 G
#447080000000
0!
0*
09
0>
0C
#447090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#447100000000
0!
0*
09
0>
0C
#447110000000
1!
1*
b101 6
19
1>
1C
b101 G
#447120000000
0!
0*
09
0>
0C
#447130000000
1!
1*
b110 6
19
1>
1C
b110 G
#447140000000
0!
0*
09
0>
0C
#447150000000
1!
1*
b111 6
19
1>
1C
b111 G
#447160000000
0!
0*
09
0>
0C
#447170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#447180000000
0!
0*
09
0>
0C
#447190000000
1!
1*
b1 6
19
1>
1C
b1 G
#447200000000
0!
0*
09
0>
0C
#447210000000
1!
1*
b10 6
19
1>
1C
b10 G
#447220000000
0!
0*
09
0>
0C
#447230000000
1!
1*
b11 6
19
1>
1C
b11 G
#447240000000
0!
0*
09
0>
0C
#447250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#447260000000
0!
0*
09
0>
0C
#447270000000
1!
1*
b101 6
19
1>
1C
b101 G
#447280000000
0!
0*
09
0>
0C
#447290000000
1!
1*
b110 6
19
1>
1C
b110 G
#447300000000
0!
0*
09
0>
0C
#447310000000
1!
1*
b111 6
19
1>
1C
b111 G
#447320000000
0!
0*
09
0>
0C
#447330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#447340000000
0!
0*
09
0>
0C
#447350000000
1!
1*
b1 6
19
1>
1C
b1 G
#447360000000
0!
0*
09
0>
0C
#447370000000
1!
1*
b10 6
19
1>
1C
b10 G
#447380000000
0!
0*
09
0>
0C
#447390000000
1!
1*
b11 6
19
1>
1C
b11 G
#447400000000
0!
0*
09
0>
0C
#447410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#447420000000
0!
0*
09
0>
0C
#447430000000
1!
1*
b101 6
19
1>
1C
b101 G
#447440000000
0!
0*
09
0>
0C
#447450000000
1!
1*
b110 6
19
1>
1C
b110 G
#447460000000
0!
0*
09
0>
0C
#447470000000
1!
1*
b111 6
19
1>
1C
b111 G
#447480000000
0!
1"
0*
1+
09
1:
0>
0C
#447490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#447500000000
0!
0*
09
0>
0C
#447510000000
1!
1*
b1 6
19
1>
1C
b1 G
#447520000000
0!
0*
09
0>
0C
#447530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#447540000000
0!
0*
09
0>
0C
#447550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#447560000000
0!
0*
09
0>
0C
#447570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#447580000000
0!
0*
09
0>
0C
#447590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#447600000000
0!
0#
0*
0,
09
0>
0?
0C
#447610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#447620000000
0!
0*
09
0>
0C
#447630000000
1!
1*
19
1>
1C
#447640000000
0!
0*
09
0>
0C
#447650000000
1!
1*
19
1>
1C
#447660000000
0!
0*
09
0>
0C
#447670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#447680000000
0!
0*
09
0>
0C
#447690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#447700000000
0!
0*
09
0>
0C
#447710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#447720000000
0!
0*
09
0>
0C
#447730000000
1!
1*
b10 6
19
1>
1C
b10 G
#447740000000
0!
0*
09
0>
0C
#447750000000
1!
1*
b11 6
19
1>
1C
b11 G
#447760000000
0!
0*
09
0>
0C
#447770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#447780000000
0!
0*
09
0>
0C
#447790000000
1!
1*
b101 6
19
1>
1C
b101 G
#447800000000
0!
0*
09
0>
0C
#447810000000
1!
1*
b110 6
19
1>
1C
b110 G
#447820000000
0!
0*
09
0>
0C
#447830000000
1!
1*
b111 6
19
1>
1C
b111 G
#447840000000
0!
0*
09
0>
0C
#447850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#447860000000
0!
0*
09
0>
0C
#447870000000
1!
1*
b1 6
19
1>
1C
b1 G
#447880000000
0!
0*
09
0>
0C
#447890000000
1!
1*
b10 6
19
1>
1C
b10 G
#447900000000
0!
0*
09
0>
0C
#447910000000
1!
1*
b11 6
19
1>
1C
b11 G
#447920000000
0!
0*
09
0>
0C
#447930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#447940000000
0!
0*
09
0>
0C
#447950000000
1!
1*
b101 6
19
1>
1C
b101 G
#447960000000
0!
0*
09
0>
0C
#447970000000
1!
1*
b110 6
19
1>
1C
b110 G
#447980000000
0!
0*
09
0>
0C
#447990000000
1!
1*
b111 6
19
1>
1C
b111 G
#448000000000
0!
0*
09
0>
0C
#448010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#448020000000
0!
0*
09
0>
0C
#448030000000
1!
1*
b1 6
19
1>
1C
b1 G
#448040000000
0!
0*
09
0>
0C
#448050000000
1!
1*
b10 6
19
1>
1C
b10 G
#448060000000
0!
0*
09
0>
0C
#448070000000
1!
1*
b11 6
19
1>
1C
b11 G
#448080000000
0!
0*
09
0>
0C
#448090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#448100000000
0!
0*
09
0>
0C
#448110000000
1!
1*
b101 6
19
1>
1C
b101 G
#448120000000
0!
0*
09
0>
0C
#448130000000
1!
1*
b110 6
19
1>
1C
b110 G
#448140000000
0!
0*
09
0>
0C
#448150000000
1!
1*
b111 6
19
1>
1C
b111 G
#448160000000
0!
1"
0*
1+
09
1:
0>
0C
#448170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#448180000000
0!
0*
09
0>
0C
#448190000000
1!
1*
b1 6
19
1>
1C
b1 G
#448200000000
0!
0*
09
0>
0C
#448210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#448220000000
0!
0*
09
0>
0C
#448230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#448240000000
0!
0*
09
0>
0C
#448250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#448260000000
0!
0*
09
0>
0C
#448270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#448280000000
0!
0#
0*
0,
09
0>
0?
0C
#448290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#448300000000
0!
0*
09
0>
0C
#448310000000
1!
1*
19
1>
1C
#448320000000
0!
0*
09
0>
0C
#448330000000
1!
1*
19
1>
1C
#448340000000
0!
0*
09
0>
0C
#448350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#448360000000
0!
0*
09
0>
0C
#448370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#448380000000
0!
0*
09
0>
0C
#448390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#448400000000
0!
0*
09
0>
0C
#448410000000
1!
1*
b10 6
19
1>
1C
b10 G
#448420000000
0!
0*
09
0>
0C
#448430000000
1!
1*
b11 6
19
1>
1C
b11 G
#448440000000
0!
0*
09
0>
0C
#448450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#448460000000
0!
0*
09
0>
0C
#448470000000
1!
1*
b101 6
19
1>
1C
b101 G
#448480000000
0!
0*
09
0>
0C
#448490000000
1!
1*
b110 6
19
1>
1C
b110 G
#448500000000
0!
0*
09
0>
0C
#448510000000
1!
1*
b111 6
19
1>
1C
b111 G
#448520000000
0!
0*
09
0>
0C
#448530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#448540000000
0!
0*
09
0>
0C
#448550000000
1!
1*
b1 6
19
1>
1C
b1 G
#448560000000
0!
0*
09
0>
0C
#448570000000
1!
1*
b10 6
19
1>
1C
b10 G
#448580000000
0!
0*
09
0>
0C
#448590000000
1!
1*
b11 6
19
1>
1C
b11 G
#448600000000
0!
0*
09
0>
0C
#448610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#448620000000
0!
0*
09
0>
0C
#448630000000
1!
1*
b101 6
19
1>
1C
b101 G
#448640000000
0!
0*
09
0>
0C
#448650000000
1!
1*
b110 6
19
1>
1C
b110 G
#448660000000
0!
0*
09
0>
0C
#448670000000
1!
1*
b111 6
19
1>
1C
b111 G
#448680000000
0!
0*
09
0>
0C
#448690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#448700000000
0!
0*
09
0>
0C
#448710000000
1!
1*
b1 6
19
1>
1C
b1 G
#448720000000
0!
0*
09
0>
0C
#448730000000
1!
1*
b10 6
19
1>
1C
b10 G
#448740000000
0!
0*
09
0>
0C
#448750000000
1!
1*
b11 6
19
1>
1C
b11 G
#448760000000
0!
0*
09
0>
0C
#448770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#448780000000
0!
0*
09
0>
0C
#448790000000
1!
1*
b101 6
19
1>
1C
b101 G
#448800000000
0!
0*
09
0>
0C
#448810000000
1!
1*
b110 6
19
1>
1C
b110 G
#448820000000
0!
0*
09
0>
0C
#448830000000
1!
1*
b111 6
19
1>
1C
b111 G
#448840000000
0!
1"
0*
1+
09
1:
0>
0C
#448850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#448860000000
0!
0*
09
0>
0C
#448870000000
1!
1*
b1 6
19
1>
1C
b1 G
#448880000000
0!
0*
09
0>
0C
#448890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#448900000000
0!
0*
09
0>
0C
#448910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#448920000000
0!
0*
09
0>
0C
#448930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#448940000000
0!
0*
09
0>
0C
#448950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#448960000000
0!
0#
0*
0,
09
0>
0?
0C
#448970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#448980000000
0!
0*
09
0>
0C
#448990000000
1!
1*
19
1>
1C
#449000000000
0!
0*
09
0>
0C
#449010000000
1!
1*
19
1>
1C
#449020000000
0!
0*
09
0>
0C
#449030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#449040000000
0!
0*
09
0>
0C
#449050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#449060000000
0!
0*
09
0>
0C
#449070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#449080000000
0!
0*
09
0>
0C
#449090000000
1!
1*
b10 6
19
1>
1C
b10 G
#449100000000
0!
0*
09
0>
0C
#449110000000
1!
1*
b11 6
19
1>
1C
b11 G
#449120000000
0!
0*
09
0>
0C
#449130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#449140000000
0!
0*
09
0>
0C
#449150000000
1!
1*
b101 6
19
1>
1C
b101 G
#449160000000
0!
0*
09
0>
0C
#449170000000
1!
1*
b110 6
19
1>
1C
b110 G
#449180000000
0!
0*
09
0>
0C
#449190000000
1!
1*
b111 6
19
1>
1C
b111 G
#449200000000
0!
0*
09
0>
0C
#449210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#449220000000
0!
0*
09
0>
0C
#449230000000
1!
1*
b1 6
19
1>
1C
b1 G
#449240000000
0!
0*
09
0>
0C
#449250000000
1!
1*
b10 6
19
1>
1C
b10 G
#449260000000
0!
0*
09
0>
0C
#449270000000
1!
1*
b11 6
19
1>
1C
b11 G
#449280000000
0!
0*
09
0>
0C
#449290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#449300000000
0!
0*
09
0>
0C
#449310000000
1!
1*
b101 6
19
1>
1C
b101 G
#449320000000
0!
0*
09
0>
0C
#449330000000
1!
1*
b110 6
19
1>
1C
b110 G
#449340000000
0!
0*
09
0>
0C
#449350000000
1!
1*
b111 6
19
1>
1C
b111 G
#449360000000
0!
0*
09
0>
0C
#449370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#449380000000
0!
0*
09
0>
0C
#449390000000
1!
1*
b1 6
19
1>
1C
b1 G
#449400000000
0!
0*
09
0>
0C
#449410000000
1!
1*
b10 6
19
1>
1C
b10 G
#449420000000
0!
0*
09
0>
0C
#449430000000
1!
1*
b11 6
19
1>
1C
b11 G
#449440000000
0!
0*
09
0>
0C
#449450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#449460000000
0!
0*
09
0>
0C
#449470000000
1!
1*
b101 6
19
1>
1C
b101 G
#449480000000
0!
0*
09
0>
0C
#449490000000
1!
1*
b110 6
19
1>
1C
b110 G
#449500000000
0!
0*
09
0>
0C
#449510000000
1!
1*
b111 6
19
1>
1C
b111 G
#449520000000
0!
1"
0*
1+
09
1:
0>
0C
#449530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#449540000000
0!
0*
09
0>
0C
#449550000000
1!
1*
b1 6
19
1>
1C
b1 G
#449560000000
0!
0*
09
0>
0C
#449570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#449580000000
0!
0*
09
0>
0C
#449590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#449600000000
0!
0*
09
0>
0C
#449610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#449620000000
0!
0*
09
0>
0C
#449630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#449640000000
0!
0#
0*
0,
09
0>
0?
0C
#449650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#449660000000
0!
0*
09
0>
0C
#449670000000
1!
1*
19
1>
1C
#449680000000
0!
0*
09
0>
0C
#449690000000
1!
1*
19
1>
1C
#449700000000
0!
0*
09
0>
0C
#449710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#449720000000
0!
0*
09
0>
0C
#449730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#449740000000
0!
0*
09
0>
0C
#449750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#449760000000
0!
0*
09
0>
0C
#449770000000
1!
1*
b10 6
19
1>
1C
b10 G
#449780000000
0!
0*
09
0>
0C
#449790000000
1!
1*
b11 6
19
1>
1C
b11 G
#449800000000
0!
0*
09
0>
0C
#449810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#449820000000
0!
0*
09
0>
0C
#449830000000
1!
1*
b101 6
19
1>
1C
b101 G
#449840000000
0!
0*
09
0>
0C
#449850000000
1!
1*
b110 6
19
1>
1C
b110 G
#449860000000
0!
0*
09
0>
0C
#449870000000
1!
1*
b111 6
19
1>
1C
b111 G
#449880000000
0!
0*
09
0>
0C
#449890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#449900000000
0!
0*
09
0>
0C
#449910000000
1!
1*
b1 6
19
1>
1C
b1 G
#449920000000
0!
0*
09
0>
0C
#449930000000
1!
1*
b10 6
19
1>
1C
b10 G
#449940000000
0!
0*
09
0>
0C
#449950000000
1!
1*
b11 6
19
1>
1C
b11 G
#449960000000
0!
0*
09
0>
0C
#449970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#449980000000
0!
0*
09
0>
0C
#449990000000
1!
1*
b101 6
19
1>
1C
b101 G
#450000000000
0!
0*
09
0>
0C
#450010000000
1!
1*
b110 6
19
1>
1C
b110 G
#450020000000
0!
0*
09
0>
0C
#450030000000
1!
1*
b111 6
19
1>
1C
b111 G
#450040000000
0!
0*
09
0>
0C
#450050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#450060000000
0!
0*
09
0>
0C
#450070000000
1!
1*
b1 6
19
1>
1C
b1 G
#450080000000
0!
0*
09
0>
0C
#450090000000
1!
1*
b10 6
19
1>
1C
b10 G
#450100000000
0!
0*
09
0>
0C
#450110000000
1!
1*
b11 6
19
1>
1C
b11 G
#450120000000
0!
0*
09
0>
0C
#450130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#450140000000
0!
0*
09
0>
0C
#450150000000
1!
1*
b101 6
19
1>
1C
b101 G
#450160000000
0!
0*
09
0>
0C
#450170000000
1!
1*
b110 6
19
1>
1C
b110 G
#450180000000
0!
0*
09
0>
0C
#450190000000
1!
1*
b111 6
19
1>
1C
b111 G
#450200000000
0!
1"
0*
1+
09
1:
0>
0C
#450210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#450220000000
0!
0*
09
0>
0C
#450230000000
1!
1*
b1 6
19
1>
1C
b1 G
#450240000000
0!
0*
09
0>
0C
#450250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#450260000000
0!
0*
09
0>
0C
#450270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#450280000000
0!
0*
09
0>
0C
#450290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#450300000000
0!
0*
09
0>
0C
#450310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#450320000000
0!
0#
0*
0,
09
0>
0?
0C
#450330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#450340000000
0!
0*
09
0>
0C
#450350000000
1!
1*
19
1>
1C
#450360000000
0!
0*
09
0>
0C
#450370000000
1!
1*
19
1>
1C
#450380000000
0!
0*
09
0>
0C
#450390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#450400000000
0!
0*
09
0>
0C
#450410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#450420000000
0!
0*
09
0>
0C
#450430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#450440000000
0!
0*
09
0>
0C
#450450000000
1!
1*
b10 6
19
1>
1C
b10 G
#450460000000
0!
0*
09
0>
0C
#450470000000
1!
1*
b11 6
19
1>
1C
b11 G
#450480000000
0!
0*
09
0>
0C
#450490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#450500000000
0!
0*
09
0>
0C
#450510000000
1!
1*
b101 6
19
1>
1C
b101 G
#450520000000
0!
0*
09
0>
0C
#450530000000
1!
1*
b110 6
19
1>
1C
b110 G
#450540000000
0!
0*
09
0>
0C
#450550000000
1!
1*
b111 6
19
1>
1C
b111 G
#450560000000
0!
0*
09
0>
0C
#450570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#450580000000
0!
0*
09
0>
0C
#450590000000
1!
1*
b1 6
19
1>
1C
b1 G
#450600000000
0!
0*
09
0>
0C
#450610000000
1!
1*
b10 6
19
1>
1C
b10 G
#450620000000
0!
0*
09
0>
0C
#450630000000
1!
1*
b11 6
19
1>
1C
b11 G
#450640000000
0!
0*
09
0>
0C
#450650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#450660000000
0!
0*
09
0>
0C
#450670000000
1!
1*
b101 6
19
1>
1C
b101 G
#450680000000
0!
0*
09
0>
0C
#450690000000
1!
1*
b110 6
19
1>
1C
b110 G
#450700000000
0!
0*
09
0>
0C
#450710000000
1!
1*
b111 6
19
1>
1C
b111 G
#450720000000
0!
0*
09
0>
0C
#450730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#450740000000
0!
0*
09
0>
0C
#450750000000
1!
1*
b1 6
19
1>
1C
b1 G
#450760000000
0!
0*
09
0>
0C
#450770000000
1!
1*
b10 6
19
1>
1C
b10 G
#450780000000
0!
0*
09
0>
0C
#450790000000
1!
1*
b11 6
19
1>
1C
b11 G
#450800000000
0!
0*
09
0>
0C
#450810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#450820000000
0!
0*
09
0>
0C
#450830000000
1!
1*
b101 6
19
1>
1C
b101 G
#450840000000
0!
0*
09
0>
0C
#450850000000
1!
1*
b110 6
19
1>
1C
b110 G
#450860000000
0!
0*
09
0>
0C
#450870000000
1!
1*
b111 6
19
1>
1C
b111 G
#450880000000
0!
1"
0*
1+
09
1:
0>
0C
#450890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#450900000000
0!
0*
09
0>
0C
#450910000000
1!
1*
b1 6
19
1>
1C
b1 G
#450920000000
0!
0*
09
0>
0C
#450930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#450940000000
0!
0*
09
0>
0C
#450950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#450960000000
0!
0*
09
0>
0C
#450970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#450980000000
0!
0*
09
0>
0C
#450990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#451000000000
0!
0#
0*
0,
09
0>
0?
0C
#451010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#451020000000
0!
0*
09
0>
0C
#451030000000
1!
1*
19
1>
1C
#451040000000
0!
0*
09
0>
0C
#451050000000
1!
1*
19
1>
1C
#451060000000
0!
0*
09
0>
0C
#451070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#451080000000
0!
0*
09
0>
0C
#451090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#451100000000
0!
0*
09
0>
0C
#451110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#451120000000
0!
0*
09
0>
0C
#451130000000
1!
1*
b10 6
19
1>
1C
b10 G
#451140000000
0!
0*
09
0>
0C
#451150000000
1!
1*
b11 6
19
1>
1C
b11 G
#451160000000
0!
0*
09
0>
0C
#451170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#451180000000
0!
0*
09
0>
0C
#451190000000
1!
1*
b101 6
19
1>
1C
b101 G
#451200000000
0!
0*
09
0>
0C
#451210000000
1!
1*
b110 6
19
1>
1C
b110 G
#451220000000
0!
0*
09
0>
0C
#451230000000
1!
1*
b111 6
19
1>
1C
b111 G
#451240000000
0!
0*
09
0>
0C
#451250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#451260000000
0!
0*
09
0>
0C
#451270000000
1!
1*
b1 6
19
1>
1C
b1 G
#451280000000
0!
0*
09
0>
0C
#451290000000
1!
1*
b10 6
19
1>
1C
b10 G
#451300000000
0!
0*
09
0>
0C
#451310000000
1!
1*
b11 6
19
1>
1C
b11 G
#451320000000
0!
0*
09
0>
0C
#451330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#451340000000
0!
0*
09
0>
0C
#451350000000
1!
1*
b101 6
19
1>
1C
b101 G
#451360000000
0!
0*
09
0>
0C
#451370000000
1!
1*
b110 6
19
1>
1C
b110 G
#451380000000
0!
0*
09
0>
0C
#451390000000
1!
1*
b111 6
19
1>
1C
b111 G
#451400000000
0!
0*
09
0>
0C
#451410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#451420000000
0!
0*
09
0>
0C
#451430000000
1!
1*
b1 6
19
1>
1C
b1 G
#451440000000
0!
0*
09
0>
0C
#451450000000
1!
1*
b10 6
19
1>
1C
b10 G
#451460000000
0!
0*
09
0>
0C
#451470000000
1!
1*
b11 6
19
1>
1C
b11 G
#451480000000
0!
0*
09
0>
0C
#451490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#451500000000
0!
0*
09
0>
0C
#451510000000
1!
1*
b101 6
19
1>
1C
b101 G
#451520000000
0!
0*
09
0>
0C
#451530000000
1!
1*
b110 6
19
1>
1C
b110 G
#451540000000
0!
0*
09
0>
0C
#451550000000
1!
1*
b111 6
19
1>
1C
b111 G
#451560000000
0!
1"
0*
1+
09
1:
0>
0C
#451570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#451580000000
0!
0*
09
0>
0C
#451590000000
1!
1*
b1 6
19
1>
1C
b1 G
#451600000000
0!
0*
09
0>
0C
#451610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#451620000000
0!
0*
09
0>
0C
#451630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#451640000000
0!
0*
09
0>
0C
#451650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#451660000000
0!
0*
09
0>
0C
#451670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#451680000000
0!
0#
0*
0,
09
0>
0?
0C
#451690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#451700000000
0!
0*
09
0>
0C
#451710000000
1!
1*
19
1>
1C
#451720000000
0!
0*
09
0>
0C
#451730000000
1!
1*
19
1>
1C
#451740000000
0!
0*
09
0>
0C
#451750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#451760000000
0!
0*
09
0>
0C
#451770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#451780000000
0!
0*
09
0>
0C
#451790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#451800000000
0!
0*
09
0>
0C
#451810000000
1!
1*
b10 6
19
1>
1C
b10 G
#451820000000
0!
0*
09
0>
0C
#451830000000
1!
1*
b11 6
19
1>
1C
b11 G
#451840000000
0!
0*
09
0>
0C
#451850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#451860000000
0!
0*
09
0>
0C
#451870000000
1!
1*
b101 6
19
1>
1C
b101 G
#451880000000
0!
0*
09
0>
0C
#451890000000
1!
1*
b110 6
19
1>
1C
b110 G
#451900000000
0!
0*
09
0>
0C
#451910000000
1!
1*
b111 6
19
1>
1C
b111 G
#451920000000
0!
0*
09
0>
0C
#451930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#451940000000
0!
0*
09
0>
0C
#451950000000
1!
1*
b1 6
19
1>
1C
b1 G
#451960000000
0!
0*
09
0>
0C
#451970000000
1!
1*
b10 6
19
1>
1C
b10 G
#451980000000
0!
0*
09
0>
0C
#451990000000
1!
1*
b11 6
19
1>
1C
b11 G
#452000000000
0!
0*
09
0>
0C
#452010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#452020000000
0!
0*
09
0>
0C
#452030000000
1!
1*
b101 6
19
1>
1C
b101 G
#452040000000
0!
0*
09
0>
0C
#452050000000
1!
1*
b110 6
19
1>
1C
b110 G
#452060000000
0!
0*
09
0>
0C
#452070000000
1!
1*
b111 6
19
1>
1C
b111 G
#452080000000
0!
0*
09
0>
0C
#452090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#452100000000
0!
0*
09
0>
0C
#452110000000
1!
1*
b1 6
19
1>
1C
b1 G
#452120000000
0!
0*
09
0>
0C
#452130000000
1!
1*
b10 6
19
1>
1C
b10 G
#452140000000
0!
0*
09
0>
0C
#452150000000
1!
1*
b11 6
19
1>
1C
b11 G
#452160000000
0!
0*
09
0>
0C
#452170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#452180000000
0!
0*
09
0>
0C
#452190000000
1!
1*
b101 6
19
1>
1C
b101 G
#452200000000
0!
0*
09
0>
0C
#452210000000
1!
1*
b110 6
19
1>
1C
b110 G
#452220000000
0!
0*
09
0>
0C
#452230000000
1!
1*
b111 6
19
1>
1C
b111 G
#452240000000
0!
1"
0*
1+
09
1:
0>
0C
#452250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#452260000000
0!
0*
09
0>
0C
#452270000000
1!
1*
b1 6
19
1>
1C
b1 G
#452280000000
0!
0*
09
0>
0C
#452290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#452300000000
0!
0*
09
0>
0C
#452310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#452320000000
0!
0*
09
0>
0C
#452330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#452340000000
0!
0*
09
0>
0C
#452350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#452360000000
0!
0#
0*
0,
09
0>
0?
0C
#452370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#452380000000
0!
0*
09
0>
0C
#452390000000
1!
1*
19
1>
1C
#452400000000
0!
0*
09
0>
0C
#452410000000
1!
1*
19
1>
1C
#452420000000
0!
0*
09
0>
0C
#452430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#452440000000
0!
0*
09
0>
0C
#452450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#452460000000
0!
0*
09
0>
0C
#452470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#452480000000
0!
0*
09
0>
0C
#452490000000
1!
1*
b10 6
19
1>
1C
b10 G
#452500000000
0!
0*
09
0>
0C
#452510000000
1!
1*
b11 6
19
1>
1C
b11 G
#452520000000
0!
0*
09
0>
0C
#452530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#452540000000
0!
0*
09
0>
0C
#452550000000
1!
1*
b101 6
19
1>
1C
b101 G
#452560000000
0!
0*
09
0>
0C
#452570000000
1!
1*
b110 6
19
1>
1C
b110 G
#452580000000
0!
0*
09
0>
0C
#452590000000
1!
1*
b111 6
19
1>
1C
b111 G
#452600000000
0!
0*
09
0>
0C
#452610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#452620000000
0!
0*
09
0>
0C
#452630000000
1!
1*
b1 6
19
1>
1C
b1 G
#452640000000
0!
0*
09
0>
0C
#452650000000
1!
1*
b10 6
19
1>
1C
b10 G
#452660000000
0!
0*
09
0>
0C
#452670000000
1!
1*
b11 6
19
1>
1C
b11 G
#452680000000
0!
0*
09
0>
0C
#452690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#452700000000
0!
0*
09
0>
0C
#452710000000
1!
1*
b101 6
19
1>
1C
b101 G
#452720000000
0!
0*
09
0>
0C
#452730000000
1!
1*
b110 6
19
1>
1C
b110 G
#452740000000
0!
0*
09
0>
0C
#452750000000
1!
1*
b111 6
19
1>
1C
b111 G
#452760000000
0!
0*
09
0>
0C
#452770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#452780000000
0!
0*
09
0>
0C
#452790000000
1!
1*
b1 6
19
1>
1C
b1 G
#452800000000
0!
0*
09
0>
0C
#452810000000
1!
1*
b10 6
19
1>
1C
b10 G
#452820000000
0!
0*
09
0>
0C
#452830000000
1!
1*
b11 6
19
1>
1C
b11 G
#452840000000
0!
0*
09
0>
0C
#452850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#452860000000
0!
0*
09
0>
0C
#452870000000
1!
1*
b101 6
19
1>
1C
b101 G
#452880000000
0!
0*
09
0>
0C
#452890000000
1!
1*
b110 6
19
1>
1C
b110 G
#452900000000
0!
0*
09
0>
0C
#452910000000
1!
1*
b111 6
19
1>
1C
b111 G
#452920000000
0!
1"
0*
1+
09
1:
0>
0C
#452930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#452940000000
0!
0*
09
0>
0C
#452950000000
1!
1*
b1 6
19
1>
1C
b1 G
#452960000000
0!
0*
09
0>
0C
#452970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#452980000000
0!
0*
09
0>
0C
#452990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#453000000000
0!
0*
09
0>
0C
#453010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#453020000000
0!
0*
09
0>
0C
#453030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#453040000000
0!
0#
0*
0,
09
0>
0?
0C
#453050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#453060000000
0!
0*
09
0>
0C
#453070000000
1!
1*
19
1>
1C
#453080000000
0!
0*
09
0>
0C
#453090000000
1!
1*
19
1>
1C
#453100000000
0!
0*
09
0>
0C
#453110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#453120000000
0!
0*
09
0>
0C
#453130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#453140000000
0!
0*
09
0>
0C
#453150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#453160000000
0!
0*
09
0>
0C
#453170000000
1!
1*
b10 6
19
1>
1C
b10 G
#453180000000
0!
0*
09
0>
0C
#453190000000
1!
1*
b11 6
19
1>
1C
b11 G
#453200000000
0!
0*
09
0>
0C
#453210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#453220000000
0!
0*
09
0>
0C
#453230000000
1!
1*
b101 6
19
1>
1C
b101 G
#453240000000
0!
0*
09
0>
0C
#453250000000
1!
1*
b110 6
19
1>
1C
b110 G
#453260000000
0!
0*
09
0>
0C
#453270000000
1!
1*
b111 6
19
1>
1C
b111 G
#453280000000
0!
0*
09
0>
0C
#453290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#453300000000
0!
0*
09
0>
0C
#453310000000
1!
1*
b1 6
19
1>
1C
b1 G
#453320000000
0!
0*
09
0>
0C
#453330000000
1!
1*
b10 6
19
1>
1C
b10 G
#453340000000
0!
0*
09
0>
0C
#453350000000
1!
1*
b11 6
19
1>
1C
b11 G
#453360000000
0!
0*
09
0>
0C
#453370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#453380000000
0!
0*
09
0>
0C
#453390000000
1!
1*
b101 6
19
1>
1C
b101 G
#453400000000
0!
0*
09
0>
0C
#453410000000
1!
1*
b110 6
19
1>
1C
b110 G
#453420000000
0!
0*
09
0>
0C
#453430000000
1!
1*
b111 6
19
1>
1C
b111 G
#453440000000
0!
0*
09
0>
0C
#453450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#453460000000
0!
0*
09
0>
0C
#453470000000
1!
1*
b1 6
19
1>
1C
b1 G
#453480000000
0!
0*
09
0>
0C
#453490000000
1!
1*
b10 6
19
1>
1C
b10 G
#453500000000
0!
0*
09
0>
0C
#453510000000
1!
1*
b11 6
19
1>
1C
b11 G
#453520000000
0!
0*
09
0>
0C
#453530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#453540000000
0!
0*
09
0>
0C
#453550000000
1!
1*
b101 6
19
1>
1C
b101 G
#453560000000
0!
0*
09
0>
0C
#453570000000
1!
1*
b110 6
19
1>
1C
b110 G
#453580000000
0!
0*
09
0>
0C
#453590000000
1!
1*
b111 6
19
1>
1C
b111 G
#453600000000
0!
1"
0*
1+
09
1:
0>
0C
#453610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#453620000000
0!
0*
09
0>
0C
#453630000000
1!
1*
b1 6
19
1>
1C
b1 G
#453640000000
0!
0*
09
0>
0C
#453650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#453660000000
0!
0*
09
0>
0C
#453670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#453680000000
0!
0*
09
0>
0C
#453690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#453700000000
0!
0*
09
0>
0C
#453710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#453720000000
0!
0#
0*
0,
09
0>
0?
0C
#453730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#453740000000
0!
0*
09
0>
0C
#453750000000
1!
1*
19
1>
1C
#453760000000
0!
0*
09
0>
0C
#453770000000
1!
1*
19
1>
1C
#453780000000
0!
0*
09
0>
0C
#453790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#453800000000
0!
0*
09
0>
0C
#453810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#453820000000
0!
0*
09
0>
0C
#453830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#453840000000
0!
0*
09
0>
0C
#453850000000
1!
1*
b10 6
19
1>
1C
b10 G
#453860000000
0!
0*
09
0>
0C
#453870000000
1!
1*
b11 6
19
1>
1C
b11 G
#453880000000
0!
0*
09
0>
0C
#453890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#453900000000
0!
0*
09
0>
0C
#453910000000
1!
1*
b101 6
19
1>
1C
b101 G
#453920000000
0!
0*
09
0>
0C
#453930000000
1!
1*
b110 6
19
1>
1C
b110 G
#453940000000
0!
0*
09
0>
0C
#453950000000
1!
1*
b111 6
19
1>
1C
b111 G
#453960000000
0!
0*
09
0>
0C
#453970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#453980000000
0!
0*
09
0>
0C
#453990000000
1!
1*
b1 6
19
1>
1C
b1 G
#454000000000
0!
0*
09
0>
0C
#454010000000
1!
1*
b10 6
19
1>
1C
b10 G
#454020000000
0!
0*
09
0>
0C
#454030000000
1!
1*
b11 6
19
1>
1C
b11 G
#454040000000
0!
0*
09
0>
0C
#454050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#454060000000
0!
0*
09
0>
0C
#454070000000
1!
1*
b101 6
19
1>
1C
b101 G
#454080000000
0!
0*
09
0>
0C
#454090000000
1!
1*
b110 6
19
1>
1C
b110 G
#454100000000
0!
0*
09
0>
0C
#454110000000
1!
1*
b111 6
19
1>
1C
b111 G
#454120000000
0!
0*
09
0>
0C
#454130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#454140000000
0!
0*
09
0>
0C
#454150000000
1!
1*
b1 6
19
1>
1C
b1 G
#454160000000
0!
0*
09
0>
0C
#454170000000
1!
1*
b10 6
19
1>
1C
b10 G
#454180000000
0!
0*
09
0>
0C
#454190000000
1!
1*
b11 6
19
1>
1C
b11 G
#454200000000
0!
0*
09
0>
0C
#454210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#454220000000
0!
0*
09
0>
0C
#454230000000
1!
1*
b101 6
19
1>
1C
b101 G
#454240000000
0!
0*
09
0>
0C
#454250000000
1!
1*
b110 6
19
1>
1C
b110 G
#454260000000
0!
0*
09
0>
0C
#454270000000
1!
1*
b111 6
19
1>
1C
b111 G
#454280000000
0!
1"
0*
1+
09
1:
0>
0C
#454290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#454300000000
0!
0*
09
0>
0C
#454310000000
1!
1*
b1 6
19
1>
1C
b1 G
#454320000000
0!
0*
09
0>
0C
#454330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#454340000000
0!
0*
09
0>
0C
#454350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#454360000000
0!
0*
09
0>
0C
#454370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#454380000000
0!
0*
09
0>
0C
#454390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#454400000000
0!
0#
0*
0,
09
0>
0?
0C
#454410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#454420000000
0!
0*
09
0>
0C
#454430000000
1!
1*
19
1>
1C
#454440000000
0!
0*
09
0>
0C
#454450000000
1!
1*
19
1>
1C
#454460000000
0!
0*
09
0>
0C
#454470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#454480000000
0!
0*
09
0>
0C
#454490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#454500000000
0!
0*
09
0>
0C
#454510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#454520000000
0!
0*
09
0>
0C
#454530000000
1!
1*
b10 6
19
1>
1C
b10 G
#454540000000
0!
0*
09
0>
0C
#454550000000
1!
1*
b11 6
19
1>
1C
b11 G
#454560000000
0!
0*
09
0>
0C
#454570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#454580000000
0!
0*
09
0>
0C
#454590000000
1!
1*
b101 6
19
1>
1C
b101 G
#454600000000
0!
0*
09
0>
0C
#454610000000
1!
1*
b110 6
19
1>
1C
b110 G
#454620000000
0!
0*
09
0>
0C
#454630000000
1!
1*
b111 6
19
1>
1C
b111 G
#454640000000
0!
0*
09
0>
0C
#454650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#454660000000
0!
0*
09
0>
0C
#454670000000
1!
1*
b1 6
19
1>
1C
b1 G
#454680000000
0!
0*
09
0>
0C
#454690000000
1!
1*
b10 6
19
1>
1C
b10 G
#454700000000
0!
0*
09
0>
0C
#454710000000
1!
1*
b11 6
19
1>
1C
b11 G
#454720000000
0!
0*
09
0>
0C
#454730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#454740000000
0!
0*
09
0>
0C
#454750000000
1!
1*
b101 6
19
1>
1C
b101 G
#454760000000
0!
0*
09
0>
0C
#454770000000
1!
1*
b110 6
19
1>
1C
b110 G
#454780000000
0!
0*
09
0>
0C
#454790000000
1!
1*
b111 6
19
1>
1C
b111 G
#454800000000
0!
0*
09
0>
0C
#454810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#454820000000
0!
0*
09
0>
0C
#454830000000
1!
1*
b1 6
19
1>
1C
b1 G
#454840000000
0!
0*
09
0>
0C
#454850000000
1!
1*
b10 6
19
1>
1C
b10 G
#454860000000
0!
0*
09
0>
0C
#454870000000
1!
1*
b11 6
19
1>
1C
b11 G
#454880000000
0!
0*
09
0>
0C
#454890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#454900000000
0!
0*
09
0>
0C
#454910000000
1!
1*
b101 6
19
1>
1C
b101 G
#454920000000
0!
0*
09
0>
0C
#454930000000
1!
1*
b110 6
19
1>
1C
b110 G
#454940000000
0!
0*
09
0>
0C
#454950000000
1!
1*
b111 6
19
1>
1C
b111 G
#454960000000
0!
1"
0*
1+
09
1:
0>
0C
#454970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#454980000000
0!
0*
09
0>
0C
#454990000000
1!
1*
b1 6
19
1>
1C
b1 G
#455000000000
0!
0*
09
0>
0C
#455010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#455020000000
0!
0*
09
0>
0C
#455030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#455040000000
0!
0*
09
0>
0C
#455050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#455060000000
0!
0*
09
0>
0C
#455070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#455080000000
0!
0#
0*
0,
09
0>
0?
0C
#455090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#455100000000
0!
0*
09
0>
0C
#455110000000
1!
1*
19
1>
1C
#455120000000
0!
0*
09
0>
0C
#455130000000
1!
1*
19
1>
1C
#455140000000
0!
0*
09
0>
0C
#455150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#455160000000
0!
0*
09
0>
0C
#455170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#455180000000
0!
0*
09
0>
0C
#455190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#455200000000
0!
0*
09
0>
0C
#455210000000
1!
1*
b10 6
19
1>
1C
b10 G
#455220000000
0!
0*
09
0>
0C
#455230000000
1!
1*
b11 6
19
1>
1C
b11 G
#455240000000
0!
0*
09
0>
0C
#455250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#455260000000
0!
0*
09
0>
0C
#455270000000
1!
1*
b101 6
19
1>
1C
b101 G
#455280000000
0!
0*
09
0>
0C
#455290000000
1!
1*
b110 6
19
1>
1C
b110 G
#455300000000
0!
0*
09
0>
0C
#455310000000
1!
1*
b111 6
19
1>
1C
b111 G
#455320000000
0!
0*
09
0>
0C
#455330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#455340000000
0!
0*
09
0>
0C
#455350000000
1!
1*
b1 6
19
1>
1C
b1 G
#455360000000
0!
0*
09
0>
0C
#455370000000
1!
1*
b10 6
19
1>
1C
b10 G
#455380000000
0!
0*
09
0>
0C
#455390000000
1!
1*
b11 6
19
1>
1C
b11 G
#455400000000
0!
0*
09
0>
0C
#455410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#455420000000
0!
0*
09
0>
0C
#455430000000
1!
1*
b101 6
19
1>
1C
b101 G
#455440000000
0!
0*
09
0>
0C
#455450000000
1!
1*
b110 6
19
1>
1C
b110 G
#455460000000
0!
0*
09
0>
0C
#455470000000
1!
1*
b111 6
19
1>
1C
b111 G
#455480000000
0!
0*
09
0>
0C
#455490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#455500000000
0!
0*
09
0>
0C
#455510000000
1!
1*
b1 6
19
1>
1C
b1 G
#455520000000
0!
0*
09
0>
0C
#455530000000
1!
1*
b10 6
19
1>
1C
b10 G
#455540000000
0!
0*
09
0>
0C
#455550000000
1!
1*
b11 6
19
1>
1C
b11 G
#455560000000
0!
0*
09
0>
0C
#455570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#455580000000
0!
0*
09
0>
0C
#455590000000
1!
1*
b101 6
19
1>
1C
b101 G
#455600000000
0!
0*
09
0>
0C
#455610000000
1!
1*
b110 6
19
1>
1C
b110 G
#455620000000
0!
0*
09
0>
0C
#455630000000
1!
1*
b111 6
19
1>
1C
b111 G
#455640000000
0!
1"
0*
1+
09
1:
0>
0C
#455650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#455660000000
0!
0*
09
0>
0C
#455670000000
1!
1*
b1 6
19
1>
1C
b1 G
#455680000000
0!
0*
09
0>
0C
#455690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#455700000000
0!
0*
09
0>
0C
#455710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#455720000000
0!
0*
09
0>
0C
#455730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#455740000000
0!
0*
09
0>
0C
#455750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#455760000000
0!
0#
0*
0,
09
0>
0?
0C
#455770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#455780000000
0!
0*
09
0>
0C
#455790000000
1!
1*
19
1>
1C
#455800000000
0!
0*
09
0>
0C
#455810000000
1!
1*
19
1>
1C
#455820000000
0!
0*
09
0>
0C
#455830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#455840000000
0!
0*
09
0>
0C
#455850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#455860000000
0!
0*
09
0>
0C
#455870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#455880000000
0!
0*
09
0>
0C
#455890000000
1!
1*
b10 6
19
1>
1C
b10 G
#455900000000
0!
0*
09
0>
0C
#455910000000
1!
1*
b11 6
19
1>
1C
b11 G
#455920000000
0!
0*
09
0>
0C
#455930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#455940000000
0!
0*
09
0>
0C
#455950000000
1!
1*
b101 6
19
1>
1C
b101 G
#455960000000
0!
0*
09
0>
0C
#455970000000
1!
1*
b110 6
19
1>
1C
b110 G
#455980000000
0!
0*
09
0>
0C
#455990000000
1!
1*
b111 6
19
1>
1C
b111 G
#456000000000
0!
0*
09
0>
0C
#456010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#456020000000
0!
0*
09
0>
0C
#456030000000
1!
1*
b1 6
19
1>
1C
b1 G
#456040000000
0!
0*
09
0>
0C
#456050000000
1!
1*
b10 6
19
1>
1C
b10 G
#456060000000
0!
0*
09
0>
0C
#456070000000
1!
1*
b11 6
19
1>
1C
b11 G
#456080000000
0!
0*
09
0>
0C
#456090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#456100000000
0!
0*
09
0>
0C
#456110000000
1!
1*
b101 6
19
1>
1C
b101 G
#456120000000
0!
0*
09
0>
0C
#456130000000
1!
1*
b110 6
19
1>
1C
b110 G
#456140000000
0!
0*
09
0>
0C
#456150000000
1!
1*
b111 6
19
1>
1C
b111 G
#456160000000
0!
0*
09
0>
0C
#456170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#456180000000
0!
0*
09
0>
0C
#456190000000
1!
1*
b1 6
19
1>
1C
b1 G
#456200000000
0!
0*
09
0>
0C
#456210000000
1!
1*
b10 6
19
1>
1C
b10 G
#456220000000
0!
0*
09
0>
0C
#456230000000
1!
1*
b11 6
19
1>
1C
b11 G
#456240000000
0!
0*
09
0>
0C
#456250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#456260000000
0!
0*
09
0>
0C
#456270000000
1!
1*
b101 6
19
1>
1C
b101 G
#456280000000
0!
0*
09
0>
0C
#456290000000
1!
1*
b110 6
19
1>
1C
b110 G
#456300000000
0!
0*
09
0>
0C
#456310000000
1!
1*
b111 6
19
1>
1C
b111 G
#456320000000
0!
1"
0*
1+
09
1:
0>
0C
#456330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#456340000000
0!
0*
09
0>
0C
#456350000000
1!
1*
b1 6
19
1>
1C
b1 G
#456360000000
0!
0*
09
0>
0C
#456370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#456380000000
0!
0*
09
0>
0C
#456390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#456400000000
0!
0*
09
0>
0C
#456410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#456420000000
0!
0*
09
0>
0C
#456430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#456440000000
0!
0#
0*
0,
09
0>
0?
0C
#456450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#456460000000
0!
0*
09
0>
0C
#456470000000
1!
1*
19
1>
1C
#456480000000
0!
0*
09
0>
0C
#456490000000
1!
1*
19
1>
1C
#456500000000
0!
0*
09
0>
0C
#456510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#456520000000
0!
0*
09
0>
0C
#456530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#456540000000
0!
0*
09
0>
0C
#456550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#456560000000
0!
0*
09
0>
0C
#456570000000
1!
1*
b10 6
19
1>
1C
b10 G
#456580000000
0!
0*
09
0>
0C
#456590000000
1!
1*
b11 6
19
1>
1C
b11 G
#456600000000
0!
0*
09
0>
0C
#456610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#456620000000
0!
0*
09
0>
0C
#456630000000
1!
1*
b101 6
19
1>
1C
b101 G
#456640000000
0!
0*
09
0>
0C
#456650000000
1!
1*
b110 6
19
1>
1C
b110 G
#456660000000
0!
0*
09
0>
0C
#456670000000
1!
1*
b111 6
19
1>
1C
b111 G
#456680000000
0!
0*
09
0>
0C
#456690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#456700000000
0!
0*
09
0>
0C
#456710000000
1!
1*
b1 6
19
1>
1C
b1 G
#456720000000
0!
0*
09
0>
0C
#456730000000
1!
1*
b10 6
19
1>
1C
b10 G
#456740000000
0!
0*
09
0>
0C
#456750000000
1!
1*
b11 6
19
1>
1C
b11 G
#456760000000
0!
0*
09
0>
0C
#456770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#456780000000
0!
0*
09
0>
0C
#456790000000
1!
1*
b101 6
19
1>
1C
b101 G
#456800000000
0!
0*
09
0>
0C
#456810000000
1!
1*
b110 6
19
1>
1C
b110 G
#456820000000
0!
0*
09
0>
0C
#456830000000
1!
1*
b111 6
19
1>
1C
b111 G
#456840000000
0!
0*
09
0>
0C
#456850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#456860000000
0!
0*
09
0>
0C
#456870000000
1!
1*
b1 6
19
1>
1C
b1 G
#456880000000
0!
0*
09
0>
0C
#456890000000
1!
1*
b10 6
19
1>
1C
b10 G
#456900000000
0!
0*
09
0>
0C
#456910000000
1!
1*
b11 6
19
1>
1C
b11 G
#456920000000
0!
0*
09
0>
0C
#456930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#456940000000
0!
0*
09
0>
0C
#456950000000
1!
1*
b101 6
19
1>
1C
b101 G
#456960000000
0!
0*
09
0>
0C
#456970000000
1!
1*
b110 6
19
1>
1C
b110 G
#456980000000
0!
0*
09
0>
0C
#456990000000
1!
1*
b111 6
19
1>
1C
b111 G
#457000000000
0!
1"
0*
1+
09
1:
0>
0C
#457010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#457020000000
0!
0*
09
0>
0C
#457030000000
1!
1*
b1 6
19
1>
1C
b1 G
#457040000000
0!
0*
09
0>
0C
#457050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#457060000000
0!
0*
09
0>
0C
#457070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#457080000000
0!
0*
09
0>
0C
#457090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#457100000000
0!
0*
09
0>
0C
#457110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#457120000000
0!
0#
0*
0,
09
0>
0?
0C
#457130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#457140000000
0!
0*
09
0>
0C
#457150000000
1!
1*
19
1>
1C
#457160000000
0!
0*
09
0>
0C
#457170000000
1!
1*
19
1>
1C
#457180000000
0!
0*
09
0>
0C
#457190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#457200000000
0!
0*
09
0>
0C
#457210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#457220000000
0!
0*
09
0>
0C
#457230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#457240000000
0!
0*
09
0>
0C
#457250000000
1!
1*
b10 6
19
1>
1C
b10 G
#457260000000
0!
0*
09
0>
0C
#457270000000
1!
1*
b11 6
19
1>
1C
b11 G
#457280000000
0!
0*
09
0>
0C
#457290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#457300000000
0!
0*
09
0>
0C
#457310000000
1!
1*
b101 6
19
1>
1C
b101 G
#457320000000
0!
0*
09
0>
0C
#457330000000
1!
1*
b110 6
19
1>
1C
b110 G
#457340000000
0!
0*
09
0>
0C
#457350000000
1!
1*
b111 6
19
1>
1C
b111 G
#457360000000
0!
0*
09
0>
0C
#457370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#457380000000
0!
0*
09
0>
0C
#457390000000
1!
1*
b1 6
19
1>
1C
b1 G
#457400000000
0!
0*
09
0>
0C
#457410000000
1!
1*
b10 6
19
1>
1C
b10 G
#457420000000
0!
0*
09
0>
0C
#457430000000
1!
1*
b11 6
19
1>
1C
b11 G
#457440000000
0!
0*
09
0>
0C
#457450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#457460000000
0!
0*
09
0>
0C
#457470000000
1!
1*
b101 6
19
1>
1C
b101 G
#457480000000
0!
0*
09
0>
0C
#457490000000
1!
1*
b110 6
19
1>
1C
b110 G
#457500000000
0!
0*
09
0>
0C
#457510000000
1!
1*
b111 6
19
1>
1C
b111 G
#457520000000
0!
0*
09
0>
0C
#457530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#457540000000
0!
0*
09
0>
0C
#457550000000
1!
1*
b1 6
19
1>
1C
b1 G
#457560000000
0!
0*
09
0>
0C
#457570000000
1!
1*
b10 6
19
1>
1C
b10 G
#457580000000
0!
0*
09
0>
0C
#457590000000
1!
1*
b11 6
19
1>
1C
b11 G
#457600000000
0!
0*
09
0>
0C
#457610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#457620000000
0!
0*
09
0>
0C
#457630000000
1!
1*
b101 6
19
1>
1C
b101 G
#457640000000
0!
0*
09
0>
0C
#457650000000
1!
1*
b110 6
19
1>
1C
b110 G
#457660000000
0!
0*
09
0>
0C
#457670000000
1!
1*
b111 6
19
1>
1C
b111 G
#457680000000
0!
1"
0*
1+
09
1:
0>
0C
#457690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#457700000000
0!
0*
09
0>
0C
#457710000000
1!
1*
b1 6
19
1>
1C
b1 G
#457720000000
0!
0*
09
0>
0C
#457730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#457740000000
0!
0*
09
0>
0C
#457750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#457760000000
0!
0*
09
0>
0C
#457770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#457780000000
0!
0*
09
0>
0C
#457790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#457800000000
0!
0#
0*
0,
09
0>
0?
0C
#457810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#457820000000
0!
0*
09
0>
0C
#457830000000
1!
1*
19
1>
1C
#457840000000
0!
0*
09
0>
0C
#457850000000
1!
1*
19
1>
1C
#457860000000
0!
0*
09
0>
0C
#457870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#457880000000
0!
0*
09
0>
0C
#457890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#457900000000
0!
0*
09
0>
0C
#457910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#457920000000
0!
0*
09
0>
0C
#457930000000
1!
1*
b10 6
19
1>
1C
b10 G
#457940000000
0!
0*
09
0>
0C
#457950000000
1!
1*
b11 6
19
1>
1C
b11 G
#457960000000
0!
0*
09
0>
0C
#457970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#457980000000
0!
0*
09
0>
0C
#457990000000
1!
1*
b101 6
19
1>
1C
b101 G
#458000000000
0!
0*
09
0>
0C
#458010000000
1!
1*
b110 6
19
1>
1C
b110 G
#458020000000
0!
0*
09
0>
0C
#458030000000
1!
1*
b111 6
19
1>
1C
b111 G
#458040000000
0!
0*
09
0>
0C
#458050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#458060000000
0!
0*
09
0>
0C
#458070000000
1!
1*
b1 6
19
1>
1C
b1 G
#458080000000
0!
0*
09
0>
0C
#458090000000
1!
1*
b10 6
19
1>
1C
b10 G
#458100000000
0!
0*
09
0>
0C
#458110000000
1!
1*
b11 6
19
1>
1C
b11 G
#458120000000
0!
0*
09
0>
0C
#458130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#458140000000
0!
0*
09
0>
0C
#458150000000
1!
1*
b101 6
19
1>
1C
b101 G
#458160000000
0!
0*
09
0>
0C
#458170000000
1!
1*
b110 6
19
1>
1C
b110 G
#458180000000
0!
0*
09
0>
0C
#458190000000
1!
1*
b111 6
19
1>
1C
b111 G
#458200000000
0!
0*
09
0>
0C
#458210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#458220000000
0!
0*
09
0>
0C
#458230000000
1!
1*
b1 6
19
1>
1C
b1 G
#458240000000
0!
0*
09
0>
0C
#458250000000
1!
1*
b10 6
19
1>
1C
b10 G
#458260000000
0!
0*
09
0>
0C
#458270000000
1!
1*
b11 6
19
1>
1C
b11 G
#458280000000
0!
0*
09
0>
0C
#458290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#458300000000
0!
0*
09
0>
0C
#458310000000
1!
1*
b101 6
19
1>
1C
b101 G
#458320000000
0!
0*
09
0>
0C
#458330000000
1!
1*
b110 6
19
1>
1C
b110 G
#458340000000
0!
0*
09
0>
0C
#458350000000
1!
1*
b111 6
19
1>
1C
b111 G
#458360000000
0!
1"
0*
1+
09
1:
0>
0C
#458370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#458380000000
0!
0*
09
0>
0C
#458390000000
1!
1*
b1 6
19
1>
1C
b1 G
#458400000000
0!
0*
09
0>
0C
#458410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#458420000000
0!
0*
09
0>
0C
#458430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#458440000000
0!
0*
09
0>
0C
#458450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#458460000000
0!
0*
09
0>
0C
#458470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#458480000000
0!
0#
0*
0,
09
0>
0?
0C
#458490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#458500000000
0!
0*
09
0>
0C
#458510000000
1!
1*
19
1>
1C
#458520000000
0!
0*
09
0>
0C
#458530000000
1!
1*
19
1>
1C
#458540000000
0!
0*
09
0>
0C
#458550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#458560000000
0!
0*
09
0>
0C
#458570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#458580000000
0!
0*
09
0>
0C
#458590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#458600000000
0!
0*
09
0>
0C
#458610000000
1!
1*
b10 6
19
1>
1C
b10 G
#458620000000
0!
0*
09
0>
0C
#458630000000
1!
1*
b11 6
19
1>
1C
b11 G
#458640000000
0!
0*
09
0>
0C
#458650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#458660000000
0!
0*
09
0>
0C
#458670000000
1!
1*
b101 6
19
1>
1C
b101 G
#458680000000
0!
0*
09
0>
0C
#458690000000
1!
1*
b110 6
19
1>
1C
b110 G
#458700000000
0!
0*
09
0>
0C
#458710000000
1!
1*
b111 6
19
1>
1C
b111 G
#458720000000
0!
0*
09
0>
0C
#458730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#458740000000
0!
0*
09
0>
0C
#458750000000
1!
1*
b1 6
19
1>
1C
b1 G
#458760000000
0!
0*
09
0>
0C
#458770000000
1!
1*
b10 6
19
1>
1C
b10 G
#458780000000
0!
0*
09
0>
0C
#458790000000
1!
1*
b11 6
19
1>
1C
b11 G
#458800000000
0!
0*
09
0>
0C
#458810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#458820000000
0!
0*
09
0>
0C
#458830000000
1!
1*
b101 6
19
1>
1C
b101 G
#458840000000
0!
0*
09
0>
0C
#458850000000
1!
1*
b110 6
19
1>
1C
b110 G
#458860000000
0!
0*
09
0>
0C
#458870000000
1!
1*
b111 6
19
1>
1C
b111 G
#458880000000
0!
0*
09
0>
0C
#458890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#458900000000
0!
0*
09
0>
0C
#458910000000
1!
1*
b1 6
19
1>
1C
b1 G
#458920000000
0!
0*
09
0>
0C
#458930000000
1!
1*
b10 6
19
1>
1C
b10 G
#458940000000
0!
0*
09
0>
0C
#458950000000
1!
1*
b11 6
19
1>
1C
b11 G
#458960000000
0!
0*
09
0>
0C
#458970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#458980000000
0!
0*
09
0>
0C
#458990000000
1!
1*
b101 6
19
1>
1C
b101 G
#459000000000
0!
0*
09
0>
0C
#459010000000
1!
1*
b110 6
19
1>
1C
b110 G
#459020000000
0!
0*
09
0>
0C
#459030000000
1!
1*
b111 6
19
1>
1C
b111 G
#459040000000
0!
1"
0*
1+
09
1:
0>
0C
#459050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#459060000000
0!
0*
09
0>
0C
#459070000000
1!
1*
b1 6
19
1>
1C
b1 G
#459080000000
0!
0*
09
0>
0C
#459090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#459100000000
0!
0*
09
0>
0C
#459110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#459120000000
0!
0*
09
0>
0C
#459130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#459140000000
0!
0*
09
0>
0C
#459150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#459160000000
0!
0#
0*
0,
09
0>
0?
0C
#459170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#459180000000
0!
0*
09
0>
0C
#459190000000
1!
1*
19
1>
1C
#459200000000
0!
0*
09
0>
0C
#459210000000
1!
1*
19
1>
1C
#459220000000
0!
0*
09
0>
0C
#459230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#459240000000
0!
0*
09
0>
0C
#459250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#459260000000
0!
0*
09
0>
0C
#459270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#459280000000
0!
0*
09
0>
0C
#459290000000
1!
1*
b10 6
19
1>
1C
b10 G
#459300000000
0!
0*
09
0>
0C
#459310000000
1!
1*
b11 6
19
1>
1C
b11 G
#459320000000
0!
0*
09
0>
0C
#459330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#459340000000
0!
0*
09
0>
0C
#459350000000
1!
1*
b101 6
19
1>
1C
b101 G
#459360000000
0!
0*
09
0>
0C
#459370000000
1!
1*
b110 6
19
1>
1C
b110 G
#459380000000
0!
0*
09
0>
0C
#459390000000
1!
1*
b111 6
19
1>
1C
b111 G
#459400000000
0!
0*
09
0>
0C
#459410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#459420000000
0!
0*
09
0>
0C
#459430000000
1!
1*
b1 6
19
1>
1C
b1 G
#459440000000
0!
0*
09
0>
0C
#459450000000
1!
1*
b10 6
19
1>
1C
b10 G
#459460000000
0!
0*
09
0>
0C
#459470000000
1!
1*
b11 6
19
1>
1C
b11 G
#459480000000
0!
0*
09
0>
0C
#459490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#459500000000
0!
0*
09
0>
0C
#459510000000
1!
1*
b101 6
19
1>
1C
b101 G
#459520000000
0!
0*
09
0>
0C
#459530000000
1!
1*
b110 6
19
1>
1C
b110 G
#459540000000
0!
0*
09
0>
0C
#459550000000
1!
1*
b111 6
19
1>
1C
b111 G
#459560000000
0!
0*
09
0>
0C
#459570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#459580000000
0!
0*
09
0>
0C
#459590000000
1!
1*
b1 6
19
1>
1C
b1 G
#459600000000
0!
0*
09
0>
0C
#459610000000
1!
1*
b10 6
19
1>
1C
b10 G
#459620000000
0!
0*
09
0>
0C
#459630000000
1!
1*
b11 6
19
1>
1C
b11 G
#459640000000
0!
0*
09
0>
0C
#459650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#459660000000
0!
0*
09
0>
0C
#459670000000
1!
1*
b101 6
19
1>
1C
b101 G
#459680000000
0!
0*
09
0>
0C
#459690000000
1!
1*
b110 6
19
1>
1C
b110 G
#459700000000
0!
0*
09
0>
0C
#459710000000
1!
1*
b111 6
19
1>
1C
b111 G
#459720000000
0!
1"
0*
1+
09
1:
0>
0C
#459730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#459740000000
0!
0*
09
0>
0C
#459750000000
1!
1*
b1 6
19
1>
1C
b1 G
#459760000000
0!
0*
09
0>
0C
#459770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#459780000000
0!
0*
09
0>
0C
#459790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#459800000000
0!
0*
09
0>
0C
#459810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#459820000000
0!
0*
09
0>
0C
#459830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#459840000000
0!
0#
0*
0,
09
0>
0?
0C
#459850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#459860000000
0!
0*
09
0>
0C
#459870000000
1!
1*
19
1>
1C
#459880000000
0!
0*
09
0>
0C
#459890000000
1!
1*
19
1>
1C
#459900000000
0!
0*
09
0>
0C
#459910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#459920000000
0!
0*
09
0>
0C
#459930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#459940000000
0!
0*
09
0>
0C
#459950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#459960000000
0!
0*
09
0>
0C
#459970000000
1!
1*
b10 6
19
1>
1C
b10 G
#459980000000
0!
0*
09
0>
0C
#459990000000
1!
1*
b11 6
19
1>
1C
b11 G
#460000000000
0!
0*
09
0>
0C
#460010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#460020000000
0!
0*
09
0>
0C
#460030000000
1!
1*
b101 6
19
1>
1C
b101 G
#460040000000
0!
0*
09
0>
0C
#460050000000
1!
1*
b110 6
19
1>
1C
b110 G
#460060000000
0!
0*
09
0>
0C
#460070000000
1!
1*
b111 6
19
1>
1C
b111 G
#460080000000
0!
0*
09
0>
0C
#460090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#460100000000
0!
0*
09
0>
0C
#460110000000
1!
1*
b1 6
19
1>
1C
b1 G
#460120000000
0!
0*
09
0>
0C
#460130000000
1!
1*
b10 6
19
1>
1C
b10 G
#460140000000
0!
0*
09
0>
0C
#460150000000
1!
1*
b11 6
19
1>
1C
b11 G
#460160000000
0!
0*
09
0>
0C
#460170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#460180000000
0!
0*
09
0>
0C
#460190000000
1!
1*
b101 6
19
1>
1C
b101 G
#460200000000
0!
0*
09
0>
0C
#460210000000
1!
1*
b110 6
19
1>
1C
b110 G
#460220000000
0!
0*
09
0>
0C
#460230000000
1!
1*
b111 6
19
1>
1C
b111 G
#460240000000
0!
0*
09
0>
0C
#460250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#460260000000
0!
0*
09
0>
0C
#460270000000
1!
1*
b1 6
19
1>
1C
b1 G
#460280000000
0!
0*
09
0>
0C
#460290000000
1!
1*
b10 6
19
1>
1C
b10 G
#460300000000
0!
0*
09
0>
0C
#460310000000
1!
1*
b11 6
19
1>
1C
b11 G
#460320000000
0!
0*
09
0>
0C
#460330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#460340000000
0!
0*
09
0>
0C
#460350000000
1!
1*
b101 6
19
1>
1C
b101 G
#460360000000
0!
0*
09
0>
0C
#460370000000
1!
1*
b110 6
19
1>
1C
b110 G
#460380000000
0!
0*
09
0>
0C
#460390000000
1!
1*
b111 6
19
1>
1C
b111 G
#460400000000
0!
1"
0*
1+
09
1:
0>
0C
#460410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#460420000000
0!
0*
09
0>
0C
#460430000000
1!
1*
b1 6
19
1>
1C
b1 G
#460440000000
0!
0*
09
0>
0C
#460450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#460460000000
0!
0*
09
0>
0C
#460470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#460480000000
0!
0*
09
0>
0C
#460490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#460500000000
0!
0*
09
0>
0C
#460510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#460520000000
0!
0#
0*
0,
09
0>
0?
0C
#460530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#460540000000
0!
0*
09
0>
0C
#460550000000
1!
1*
19
1>
1C
#460560000000
0!
0*
09
0>
0C
#460570000000
1!
1*
19
1>
1C
#460580000000
0!
0*
09
0>
0C
#460590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#460600000000
0!
0*
09
0>
0C
#460610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#460620000000
0!
0*
09
0>
0C
#460630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#460640000000
0!
0*
09
0>
0C
#460650000000
1!
1*
b10 6
19
1>
1C
b10 G
#460660000000
0!
0*
09
0>
0C
#460670000000
1!
1*
b11 6
19
1>
1C
b11 G
#460680000000
0!
0*
09
0>
0C
#460690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#460700000000
0!
0*
09
0>
0C
#460710000000
1!
1*
b101 6
19
1>
1C
b101 G
#460720000000
0!
0*
09
0>
0C
#460730000000
1!
1*
b110 6
19
1>
1C
b110 G
#460740000000
0!
0*
09
0>
0C
#460750000000
1!
1*
b111 6
19
1>
1C
b111 G
#460760000000
0!
0*
09
0>
0C
#460770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#460780000000
0!
0*
09
0>
0C
#460790000000
1!
1*
b1 6
19
1>
1C
b1 G
#460800000000
0!
0*
09
0>
0C
#460810000000
1!
1*
b10 6
19
1>
1C
b10 G
#460820000000
0!
0*
09
0>
0C
#460830000000
1!
1*
b11 6
19
1>
1C
b11 G
#460840000000
0!
0*
09
0>
0C
#460850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#460860000000
0!
0*
09
0>
0C
#460870000000
1!
1*
b101 6
19
1>
1C
b101 G
#460880000000
0!
0*
09
0>
0C
#460890000000
1!
1*
b110 6
19
1>
1C
b110 G
#460900000000
0!
0*
09
0>
0C
#460910000000
1!
1*
b111 6
19
1>
1C
b111 G
#460920000000
0!
0*
09
0>
0C
#460930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#460940000000
0!
0*
09
0>
0C
#460950000000
1!
1*
b1 6
19
1>
1C
b1 G
#460960000000
0!
0*
09
0>
0C
#460970000000
1!
1*
b10 6
19
1>
1C
b10 G
#460980000000
0!
0*
09
0>
0C
#460990000000
1!
1*
b11 6
19
1>
1C
b11 G
#461000000000
0!
0*
09
0>
0C
#461010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#461020000000
0!
0*
09
0>
0C
#461030000000
1!
1*
b101 6
19
1>
1C
b101 G
#461040000000
0!
0*
09
0>
0C
#461050000000
1!
1*
b110 6
19
1>
1C
b110 G
#461060000000
0!
0*
09
0>
0C
#461070000000
1!
1*
b111 6
19
1>
1C
b111 G
#461080000000
0!
1"
0*
1+
09
1:
0>
0C
#461090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#461100000000
0!
0*
09
0>
0C
#461110000000
1!
1*
b1 6
19
1>
1C
b1 G
#461120000000
0!
0*
09
0>
0C
#461130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#461140000000
0!
0*
09
0>
0C
#461150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#461160000000
0!
0*
09
0>
0C
#461170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#461180000000
0!
0*
09
0>
0C
#461190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#461200000000
0!
0#
0*
0,
09
0>
0?
0C
#461210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#461220000000
0!
0*
09
0>
0C
#461230000000
1!
1*
19
1>
1C
#461240000000
0!
0*
09
0>
0C
#461250000000
1!
1*
19
1>
1C
#461260000000
0!
0*
09
0>
0C
#461270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#461280000000
0!
0*
09
0>
0C
#461290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#461300000000
0!
0*
09
0>
0C
#461310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#461320000000
0!
0*
09
0>
0C
#461330000000
1!
1*
b10 6
19
1>
1C
b10 G
#461340000000
0!
0*
09
0>
0C
#461350000000
1!
1*
b11 6
19
1>
1C
b11 G
#461360000000
0!
0*
09
0>
0C
#461370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#461380000000
0!
0*
09
0>
0C
#461390000000
1!
1*
b101 6
19
1>
1C
b101 G
#461400000000
0!
0*
09
0>
0C
#461410000000
1!
1*
b110 6
19
1>
1C
b110 G
#461420000000
0!
0*
09
0>
0C
#461430000000
1!
1*
b111 6
19
1>
1C
b111 G
#461440000000
0!
0*
09
0>
0C
#461450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#461460000000
0!
0*
09
0>
0C
#461470000000
1!
1*
b1 6
19
1>
1C
b1 G
#461480000000
0!
0*
09
0>
0C
#461490000000
1!
1*
b10 6
19
1>
1C
b10 G
#461500000000
0!
0*
09
0>
0C
#461510000000
1!
1*
b11 6
19
1>
1C
b11 G
#461520000000
0!
0*
09
0>
0C
#461530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#461540000000
0!
0*
09
0>
0C
#461550000000
1!
1*
b101 6
19
1>
1C
b101 G
#461560000000
0!
0*
09
0>
0C
#461570000000
1!
1*
b110 6
19
1>
1C
b110 G
#461580000000
0!
0*
09
0>
0C
#461590000000
1!
1*
b111 6
19
1>
1C
b111 G
#461600000000
0!
0*
09
0>
0C
#461610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#461620000000
0!
0*
09
0>
0C
#461630000000
1!
1*
b1 6
19
1>
1C
b1 G
#461640000000
0!
0*
09
0>
0C
#461650000000
1!
1*
b10 6
19
1>
1C
b10 G
#461660000000
0!
0*
09
0>
0C
#461670000000
1!
1*
b11 6
19
1>
1C
b11 G
#461680000000
0!
0*
09
0>
0C
#461690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#461700000000
0!
0*
09
0>
0C
#461710000000
1!
1*
b101 6
19
1>
1C
b101 G
#461720000000
0!
0*
09
0>
0C
#461730000000
1!
1*
b110 6
19
1>
1C
b110 G
#461740000000
0!
0*
09
0>
0C
#461750000000
1!
1*
b111 6
19
1>
1C
b111 G
#461760000000
0!
1"
0*
1+
09
1:
0>
0C
#461770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#461780000000
0!
0*
09
0>
0C
#461790000000
1!
1*
b1 6
19
1>
1C
b1 G
#461800000000
0!
0*
09
0>
0C
#461810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#461820000000
0!
0*
09
0>
0C
#461830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#461840000000
0!
0*
09
0>
0C
#461850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#461860000000
0!
0*
09
0>
0C
#461870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#461880000000
0!
0#
0*
0,
09
0>
0?
0C
#461890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#461900000000
0!
0*
09
0>
0C
#461910000000
1!
1*
19
1>
1C
#461920000000
0!
0*
09
0>
0C
#461930000000
1!
1*
19
1>
1C
#461940000000
0!
0*
09
0>
0C
#461950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#461960000000
0!
0*
09
0>
0C
#461970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#461980000000
0!
0*
09
0>
0C
#461990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#462000000000
0!
0*
09
0>
0C
#462010000000
1!
1*
b10 6
19
1>
1C
b10 G
#462020000000
0!
0*
09
0>
0C
#462030000000
1!
1*
b11 6
19
1>
1C
b11 G
#462040000000
0!
0*
09
0>
0C
#462050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#462060000000
0!
0*
09
0>
0C
#462070000000
1!
1*
b101 6
19
1>
1C
b101 G
#462080000000
0!
0*
09
0>
0C
#462090000000
1!
1*
b110 6
19
1>
1C
b110 G
#462100000000
0!
0*
09
0>
0C
#462110000000
1!
1*
b111 6
19
1>
1C
b111 G
#462120000000
0!
0*
09
0>
0C
#462130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#462140000000
0!
0*
09
0>
0C
#462150000000
1!
1*
b1 6
19
1>
1C
b1 G
#462160000000
0!
0*
09
0>
0C
#462170000000
1!
1*
b10 6
19
1>
1C
b10 G
#462180000000
0!
0*
09
0>
0C
#462190000000
1!
1*
b11 6
19
1>
1C
b11 G
#462200000000
0!
0*
09
0>
0C
#462210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#462220000000
0!
0*
09
0>
0C
#462230000000
1!
1*
b101 6
19
1>
1C
b101 G
#462240000000
0!
0*
09
0>
0C
#462250000000
1!
1*
b110 6
19
1>
1C
b110 G
#462260000000
0!
0*
09
0>
0C
#462270000000
1!
1*
b111 6
19
1>
1C
b111 G
#462280000000
0!
0*
09
0>
0C
#462290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#462300000000
0!
0*
09
0>
0C
#462310000000
1!
1*
b1 6
19
1>
1C
b1 G
#462320000000
0!
0*
09
0>
0C
#462330000000
1!
1*
b10 6
19
1>
1C
b10 G
#462340000000
0!
0*
09
0>
0C
#462350000000
1!
1*
b11 6
19
1>
1C
b11 G
#462360000000
0!
0*
09
0>
0C
#462370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#462380000000
0!
0*
09
0>
0C
#462390000000
1!
1*
b101 6
19
1>
1C
b101 G
#462400000000
0!
0*
09
0>
0C
#462410000000
1!
1*
b110 6
19
1>
1C
b110 G
#462420000000
0!
0*
09
0>
0C
#462430000000
1!
1*
b111 6
19
1>
1C
b111 G
#462440000000
0!
1"
0*
1+
09
1:
0>
0C
#462450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#462460000000
0!
0*
09
0>
0C
#462470000000
1!
1*
b1 6
19
1>
1C
b1 G
#462480000000
0!
0*
09
0>
0C
#462490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#462500000000
0!
0*
09
0>
0C
#462510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#462520000000
0!
0*
09
0>
0C
#462530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#462540000000
0!
0*
09
0>
0C
#462550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#462560000000
0!
0#
0*
0,
09
0>
0?
0C
#462570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#462580000000
0!
0*
09
0>
0C
#462590000000
1!
1*
19
1>
1C
#462600000000
0!
0*
09
0>
0C
#462610000000
1!
1*
19
1>
1C
#462620000000
0!
0*
09
0>
0C
#462630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#462640000000
0!
0*
09
0>
0C
#462650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#462660000000
0!
0*
09
0>
0C
#462670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#462680000000
0!
0*
09
0>
0C
#462690000000
1!
1*
b10 6
19
1>
1C
b10 G
#462700000000
0!
0*
09
0>
0C
#462710000000
1!
1*
b11 6
19
1>
1C
b11 G
#462720000000
0!
0*
09
0>
0C
#462730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#462740000000
0!
0*
09
0>
0C
#462750000000
1!
1*
b101 6
19
1>
1C
b101 G
#462760000000
0!
0*
09
0>
0C
#462770000000
1!
1*
b110 6
19
1>
1C
b110 G
#462780000000
0!
0*
09
0>
0C
#462790000000
1!
1*
b111 6
19
1>
1C
b111 G
#462800000000
0!
0*
09
0>
0C
#462810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#462820000000
0!
0*
09
0>
0C
#462830000000
1!
1*
b1 6
19
1>
1C
b1 G
#462840000000
0!
0*
09
0>
0C
#462850000000
1!
1*
b10 6
19
1>
1C
b10 G
#462860000000
0!
0*
09
0>
0C
#462870000000
1!
1*
b11 6
19
1>
1C
b11 G
#462880000000
0!
0*
09
0>
0C
#462890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#462900000000
0!
0*
09
0>
0C
#462910000000
1!
1*
b101 6
19
1>
1C
b101 G
#462920000000
0!
0*
09
0>
0C
#462930000000
1!
1*
b110 6
19
1>
1C
b110 G
#462940000000
0!
0*
09
0>
0C
#462950000000
1!
1*
b111 6
19
1>
1C
b111 G
#462960000000
0!
0*
09
0>
0C
#462970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#462980000000
0!
0*
09
0>
0C
#462990000000
1!
1*
b1 6
19
1>
1C
b1 G
#463000000000
0!
0*
09
0>
0C
#463010000000
1!
1*
b10 6
19
1>
1C
b10 G
#463020000000
0!
0*
09
0>
0C
#463030000000
1!
1*
b11 6
19
1>
1C
b11 G
#463040000000
0!
0*
09
0>
0C
#463050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#463060000000
0!
0*
09
0>
0C
#463070000000
1!
1*
b101 6
19
1>
1C
b101 G
#463080000000
0!
0*
09
0>
0C
#463090000000
1!
1*
b110 6
19
1>
1C
b110 G
#463100000000
0!
0*
09
0>
0C
#463110000000
1!
1*
b111 6
19
1>
1C
b111 G
#463120000000
0!
1"
0*
1+
09
1:
0>
0C
#463130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#463140000000
0!
0*
09
0>
0C
#463150000000
1!
1*
b1 6
19
1>
1C
b1 G
#463160000000
0!
0*
09
0>
0C
#463170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#463180000000
0!
0*
09
0>
0C
#463190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#463200000000
0!
0*
09
0>
0C
#463210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#463220000000
0!
0*
09
0>
0C
#463230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#463240000000
0!
0#
0*
0,
09
0>
0?
0C
#463250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#463260000000
0!
0*
09
0>
0C
#463270000000
1!
1*
19
1>
1C
#463280000000
0!
0*
09
0>
0C
#463290000000
1!
1*
19
1>
1C
#463300000000
0!
0*
09
0>
0C
#463310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#463320000000
0!
0*
09
0>
0C
#463330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#463340000000
0!
0*
09
0>
0C
#463350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#463360000000
0!
0*
09
0>
0C
#463370000000
1!
1*
b10 6
19
1>
1C
b10 G
#463380000000
0!
0*
09
0>
0C
#463390000000
1!
1*
b11 6
19
1>
1C
b11 G
#463400000000
0!
0*
09
0>
0C
#463410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#463420000000
0!
0*
09
0>
0C
#463430000000
1!
1*
b101 6
19
1>
1C
b101 G
#463440000000
0!
0*
09
0>
0C
#463450000000
1!
1*
b110 6
19
1>
1C
b110 G
#463460000000
0!
0*
09
0>
0C
#463470000000
1!
1*
b111 6
19
1>
1C
b111 G
#463480000000
0!
0*
09
0>
0C
#463490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#463500000000
0!
0*
09
0>
0C
#463510000000
1!
1*
b1 6
19
1>
1C
b1 G
#463520000000
0!
0*
09
0>
0C
#463530000000
1!
1*
b10 6
19
1>
1C
b10 G
#463540000000
0!
0*
09
0>
0C
#463550000000
1!
1*
b11 6
19
1>
1C
b11 G
#463560000000
0!
0*
09
0>
0C
#463570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#463580000000
0!
0*
09
0>
0C
#463590000000
1!
1*
b101 6
19
1>
1C
b101 G
#463600000000
0!
0*
09
0>
0C
#463610000000
1!
1*
b110 6
19
1>
1C
b110 G
#463620000000
0!
0*
09
0>
0C
#463630000000
1!
1*
b111 6
19
1>
1C
b111 G
#463640000000
0!
0*
09
0>
0C
#463650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#463660000000
0!
0*
09
0>
0C
#463670000000
1!
1*
b1 6
19
1>
1C
b1 G
#463680000000
0!
0*
09
0>
0C
#463690000000
1!
1*
b10 6
19
1>
1C
b10 G
#463700000000
0!
0*
09
0>
0C
#463710000000
1!
1*
b11 6
19
1>
1C
b11 G
#463720000000
0!
0*
09
0>
0C
#463730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#463740000000
0!
0*
09
0>
0C
#463750000000
1!
1*
b101 6
19
1>
1C
b101 G
#463760000000
0!
0*
09
0>
0C
#463770000000
1!
1*
b110 6
19
1>
1C
b110 G
#463780000000
0!
0*
09
0>
0C
#463790000000
1!
1*
b111 6
19
1>
1C
b111 G
#463800000000
0!
1"
0*
1+
09
1:
0>
0C
#463810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#463820000000
0!
0*
09
0>
0C
#463830000000
1!
1*
b1 6
19
1>
1C
b1 G
#463840000000
0!
0*
09
0>
0C
#463850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#463860000000
0!
0*
09
0>
0C
#463870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#463880000000
0!
0*
09
0>
0C
#463890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#463900000000
0!
0*
09
0>
0C
#463910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#463920000000
0!
0#
0*
0,
09
0>
0?
0C
#463930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#463940000000
0!
0*
09
0>
0C
#463950000000
1!
1*
19
1>
1C
#463960000000
0!
0*
09
0>
0C
#463970000000
1!
1*
19
1>
1C
#463980000000
0!
0*
09
0>
0C
#463990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#464000000000
0!
0*
09
0>
0C
#464010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#464020000000
0!
0*
09
0>
0C
#464030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#464040000000
0!
0*
09
0>
0C
#464050000000
1!
1*
b10 6
19
1>
1C
b10 G
#464060000000
0!
0*
09
0>
0C
#464070000000
1!
1*
b11 6
19
1>
1C
b11 G
#464080000000
0!
0*
09
0>
0C
#464090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#464100000000
0!
0*
09
0>
0C
#464110000000
1!
1*
b101 6
19
1>
1C
b101 G
#464120000000
0!
0*
09
0>
0C
#464130000000
1!
1*
b110 6
19
1>
1C
b110 G
#464140000000
0!
0*
09
0>
0C
#464150000000
1!
1*
b111 6
19
1>
1C
b111 G
#464160000000
0!
0*
09
0>
0C
#464170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#464180000000
0!
0*
09
0>
0C
#464190000000
1!
1*
b1 6
19
1>
1C
b1 G
#464200000000
0!
0*
09
0>
0C
#464210000000
1!
1*
b10 6
19
1>
1C
b10 G
#464220000000
0!
0*
09
0>
0C
#464230000000
1!
1*
b11 6
19
1>
1C
b11 G
#464240000000
0!
0*
09
0>
0C
#464250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#464260000000
0!
0*
09
0>
0C
#464270000000
1!
1*
b101 6
19
1>
1C
b101 G
#464280000000
0!
0*
09
0>
0C
#464290000000
1!
1*
b110 6
19
1>
1C
b110 G
#464300000000
0!
0*
09
0>
0C
#464310000000
1!
1*
b111 6
19
1>
1C
b111 G
#464320000000
0!
0*
09
0>
0C
#464330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#464340000000
0!
0*
09
0>
0C
#464350000000
1!
1*
b1 6
19
1>
1C
b1 G
#464360000000
0!
0*
09
0>
0C
#464370000000
1!
1*
b10 6
19
1>
1C
b10 G
#464380000000
0!
0*
09
0>
0C
#464390000000
1!
1*
b11 6
19
1>
1C
b11 G
#464400000000
0!
0*
09
0>
0C
#464410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#464420000000
0!
0*
09
0>
0C
#464430000000
1!
1*
b101 6
19
1>
1C
b101 G
#464440000000
0!
0*
09
0>
0C
#464450000000
1!
1*
b110 6
19
1>
1C
b110 G
#464460000000
0!
0*
09
0>
0C
#464470000000
1!
1*
b111 6
19
1>
1C
b111 G
#464480000000
0!
1"
0*
1+
09
1:
0>
0C
#464490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#464500000000
0!
0*
09
0>
0C
#464510000000
1!
1*
b1 6
19
1>
1C
b1 G
#464520000000
0!
0*
09
0>
0C
#464530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#464540000000
0!
0*
09
0>
0C
#464550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#464560000000
0!
0*
09
0>
0C
#464570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#464580000000
0!
0*
09
0>
0C
#464590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#464600000000
0!
0#
0*
0,
09
0>
0?
0C
#464610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#464620000000
0!
0*
09
0>
0C
#464630000000
1!
1*
19
1>
1C
#464640000000
0!
0*
09
0>
0C
#464650000000
1!
1*
19
1>
1C
#464660000000
0!
0*
09
0>
0C
#464670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#464680000000
0!
0*
09
0>
0C
#464690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#464700000000
0!
0*
09
0>
0C
#464710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#464720000000
0!
0*
09
0>
0C
#464730000000
1!
1*
b10 6
19
1>
1C
b10 G
#464740000000
0!
0*
09
0>
0C
#464750000000
1!
1*
b11 6
19
1>
1C
b11 G
#464760000000
0!
0*
09
0>
0C
#464770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#464780000000
0!
0*
09
0>
0C
#464790000000
1!
1*
b101 6
19
1>
1C
b101 G
#464800000000
0!
0*
09
0>
0C
#464810000000
1!
1*
b110 6
19
1>
1C
b110 G
#464820000000
0!
0*
09
0>
0C
#464830000000
1!
1*
b111 6
19
1>
1C
b111 G
#464840000000
0!
0*
09
0>
0C
#464850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#464860000000
0!
0*
09
0>
0C
#464870000000
1!
1*
b1 6
19
1>
1C
b1 G
#464880000000
0!
0*
09
0>
0C
#464890000000
1!
1*
b10 6
19
1>
1C
b10 G
#464900000000
0!
0*
09
0>
0C
#464910000000
1!
1*
b11 6
19
1>
1C
b11 G
#464920000000
0!
0*
09
0>
0C
#464930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#464940000000
0!
0*
09
0>
0C
#464950000000
1!
1*
b101 6
19
1>
1C
b101 G
#464960000000
0!
0*
09
0>
0C
#464970000000
1!
1*
b110 6
19
1>
1C
b110 G
#464980000000
0!
0*
09
0>
0C
#464990000000
1!
1*
b111 6
19
1>
1C
b111 G
#465000000000
0!
0*
09
0>
0C
#465010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#465020000000
0!
0*
09
0>
0C
#465030000000
1!
1*
b1 6
19
1>
1C
b1 G
#465040000000
0!
0*
09
0>
0C
#465050000000
1!
1*
b10 6
19
1>
1C
b10 G
#465060000000
0!
0*
09
0>
0C
#465070000000
1!
1*
b11 6
19
1>
1C
b11 G
#465080000000
0!
0*
09
0>
0C
#465090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#465100000000
0!
0*
09
0>
0C
#465110000000
1!
1*
b101 6
19
1>
1C
b101 G
#465120000000
0!
0*
09
0>
0C
#465130000000
1!
1*
b110 6
19
1>
1C
b110 G
#465140000000
0!
0*
09
0>
0C
#465150000000
1!
1*
b111 6
19
1>
1C
b111 G
#465160000000
0!
1"
0*
1+
09
1:
0>
0C
#465170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#465180000000
0!
0*
09
0>
0C
#465190000000
1!
1*
b1 6
19
1>
1C
b1 G
#465200000000
0!
0*
09
0>
0C
#465210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#465220000000
0!
0*
09
0>
0C
#465230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#465240000000
0!
0*
09
0>
0C
#465250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#465260000000
0!
0*
09
0>
0C
#465270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#465280000000
0!
0#
0*
0,
09
0>
0?
0C
#465290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#465300000000
0!
0*
09
0>
0C
#465310000000
1!
1*
19
1>
1C
#465320000000
0!
0*
09
0>
0C
#465330000000
1!
1*
19
1>
1C
#465340000000
0!
0*
09
0>
0C
#465350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#465360000000
0!
0*
09
0>
0C
#465370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#465380000000
0!
0*
09
0>
0C
#465390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#465400000000
0!
0*
09
0>
0C
#465410000000
1!
1*
b10 6
19
1>
1C
b10 G
#465420000000
0!
0*
09
0>
0C
#465430000000
1!
1*
b11 6
19
1>
1C
b11 G
#465440000000
0!
0*
09
0>
0C
#465450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#465460000000
0!
0*
09
0>
0C
#465470000000
1!
1*
b101 6
19
1>
1C
b101 G
#465480000000
0!
0*
09
0>
0C
#465490000000
1!
1*
b110 6
19
1>
1C
b110 G
#465500000000
0!
0*
09
0>
0C
#465510000000
1!
1*
b111 6
19
1>
1C
b111 G
#465520000000
0!
0*
09
0>
0C
#465530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#465540000000
0!
0*
09
0>
0C
#465550000000
1!
1*
b1 6
19
1>
1C
b1 G
#465560000000
0!
0*
09
0>
0C
#465570000000
1!
1*
b10 6
19
1>
1C
b10 G
#465580000000
0!
0*
09
0>
0C
#465590000000
1!
1*
b11 6
19
1>
1C
b11 G
#465600000000
0!
0*
09
0>
0C
#465610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#465620000000
0!
0*
09
0>
0C
#465630000000
1!
1*
b101 6
19
1>
1C
b101 G
#465640000000
0!
0*
09
0>
0C
#465650000000
1!
1*
b110 6
19
1>
1C
b110 G
#465660000000
0!
0*
09
0>
0C
#465670000000
1!
1*
b111 6
19
1>
1C
b111 G
#465680000000
0!
0*
09
0>
0C
#465690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#465700000000
0!
0*
09
0>
0C
#465710000000
1!
1*
b1 6
19
1>
1C
b1 G
#465720000000
0!
0*
09
0>
0C
#465730000000
1!
1*
b10 6
19
1>
1C
b10 G
#465740000000
0!
0*
09
0>
0C
#465750000000
1!
1*
b11 6
19
1>
1C
b11 G
#465760000000
0!
0*
09
0>
0C
#465770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#465780000000
0!
0*
09
0>
0C
#465790000000
1!
1*
b101 6
19
1>
1C
b101 G
#465800000000
0!
0*
09
0>
0C
#465810000000
1!
1*
b110 6
19
1>
1C
b110 G
#465820000000
0!
0*
09
0>
0C
#465830000000
1!
1*
b111 6
19
1>
1C
b111 G
#465840000000
0!
1"
0*
1+
09
1:
0>
0C
#465850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#465860000000
0!
0*
09
0>
0C
#465870000000
1!
1*
b1 6
19
1>
1C
b1 G
#465880000000
0!
0*
09
0>
0C
#465890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#465900000000
0!
0*
09
0>
0C
#465910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#465920000000
0!
0*
09
0>
0C
#465930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#465940000000
0!
0*
09
0>
0C
#465950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#465960000000
0!
0#
0*
0,
09
0>
0?
0C
#465970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#465980000000
0!
0*
09
0>
0C
#465990000000
1!
1*
19
1>
1C
#466000000000
0!
0*
09
0>
0C
#466010000000
1!
1*
19
1>
1C
#466020000000
0!
0*
09
0>
0C
#466030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#466040000000
0!
0*
09
0>
0C
#466050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#466060000000
0!
0*
09
0>
0C
#466070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#466080000000
0!
0*
09
0>
0C
#466090000000
1!
1*
b10 6
19
1>
1C
b10 G
#466100000000
0!
0*
09
0>
0C
#466110000000
1!
1*
b11 6
19
1>
1C
b11 G
#466120000000
0!
0*
09
0>
0C
#466130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#466140000000
0!
0*
09
0>
0C
#466150000000
1!
1*
b101 6
19
1>
1C
b101 G
#466160000000
0!
0*
09
0>
0C
#466170000000
1!
1*
b110 6
19
1>
1C
b110 G
#466180000000
0!
0*
09
0>
0C
#466190000000
1!
1*
b111 6
19
1>
1C
b111 G
#466200000000
0!
0*
09
0>
0C
#466210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#466220000000
0!
0*
09
0>
0C
#466230000000
1!
1*
b1 6
19
1>
1C
b1 G
#466240000000
0!
0*
09
0>
0C
#466250000000
1!
1*
b10 6
19
1>
1C
b10 G
#466260000000
0!
0*
09
0>
0C
#466270000000
1!
1*
b11 6
19
1>
1C
b11 G
#466280000000
0!
0*
09
0>
0C
#466290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#466300000000
0!
0*
09
0>
0C
#466310000000
1!
1*
b101 6
19
1>
1C
b101 G
#466320000000
0!
0*
09
0>
0C
#466330000000
1!
1*
b110 6
19
1>
1C
b110 G
#466340000000
0!
0*
09
0>
0C
#466350000000
1!
1*
b111 6
19
1>
1C
b111 G
#466360000000
0!
0*
09
0>
0C
#466370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#466380000000
0!
0*
09
0>
0C
#466390000000
1!
1*
b1 6
19
1>
1C
b1 G
#466400000000
0!
0*
09
0>
0C
#466410000000
1!
1*
b10 6
19
1>
1C
b10 G
#466420000000
0!
0*
09
0>
0C
#466430000000
1!
1*
b11 6
19
1>
1C
b11 G
#466440000000
0!
0*
09
0>
0C
#466450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#466460000000
0!
0*
09
0>
0C
#466470000000
1!
1*
b101 6
19
1>
1C
b101 G
#466480000000
0!
0*
09
0>
0C
#466490000000
1!
1*
b110 6
19
1>
1C
b110 G
#466500000000
0!
0*
09
0>
0C
#466510000000
1!
1*
b111 6
19
1>
1C
b111 G
#466520000000
0!
1"
0*
1+
09
1:
0>
0C
#466530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#466540000000
0!
0*
09
0>
0C
#466550000000
1!
1*
b1 6
19
1>
1C
b1 G
#466560000000
0!
0*
09
0>
0C
#466570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#466580000000
0!
0*
09
0>
0C
#466590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#466600000000
0!
0*
09
0>
0C
#466610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#466620000000
0!
0*
09
0>
0C
#466630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#466640000000
0!
0#
0*
0,
09
0>
0?
0C
#466650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#466660000000
0!
0*
09
0>
0C
#466670000000
1!
1*
19
1>
1C
#466680000000
0!
0*
09
0>
0C
#466690000000
1!
1*
19
1>
1C
#466700000000
0!
0*
09
0>
0C
#466710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#466720000000
0!
0*
09
0>
0C
#466730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#466740000000
0!
0*
09
0>
0C
#466750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#466760000000
0!
0*
09
0>
0C
#466770000000
1!
1*
b10 6
19
1>
1C
b10 G
#466780000000
0!
0*
09
0>
0C
#466790000000
1!
1*
b11 6
19
1>
1C
b11 G
#466800000000
0!
0*
09
0>
0C
#466810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#466820000000
0!
0*
09
0>
0C
#466830000000
1!
1*
b101 6
19
1>
1C
b101 G
#466840000000
0!
0*
09
0>
0C
#466850000000
1!
1*
b110 6
19
1>
1C
b110 G
#466860000000
0!
0*
09
0>
0C
#466870000000
1!
1*
b111 6
19
1>
1C
b111 G
#466880000000
0!
0*
09
0>
0C
#466890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#466900000000
0!
0*
09
0>
0C
#466910000000
1!
1*
b1 6
19
1>
1C
b1 G
#466920000000
0!
0*
09
0>
0C
#466930000000
1!
1*
b10 6
19
1>
1C
b10 G
#466940000000
0!
0*
09
0>
0C
#466950000000
1!
1*
b11 6
19
1>
1C
b11 G
#466960000000
0!
0*
09
0>
0C
#466970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#466980000000
0!
0*
09
0>
0C
#466990000000
1!
1*
b101 6
19
1>
1C
b101 G
#467000000000
0!
0*
09
0>
0C
#467010000000
1!
1*
b110 6
19
1>
1C
b110 G
#467020000000
0!
0*
09
0>
0C
#467030000000
1!
1*
b111 6
19
1>
1C
b111 G
#467040000000
0!
0*
09
0>
0C
#467050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#467060000000
0!
0*
09
0>
0C
#467070000000
1!
1*
b1 6
19
1>
1C
b1 G
#467080000000
0!
0*
09
0>
0C
#467090000000
1!
1*
b10 6
19
1>
1C
b10 G
#467100000000
0!
0*
09
0>
0C
#467110000000
1!
1*
b11 6
19
1>
1C
b11 G
#467120000000
0!
0*
09
0>
0C
#467130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#467140000000
0!
0*
09
0>
0C
#467150000000
1!
1*
b101 6
19
1>
1C
b101 G
#467160000000
0!
0*
09
0>
0C
#467170000000
1!
1*
b110 6
19
1>
1C
b110 G
#467180000000
0!
0*
09
0>
0C
#467190000000
1!
1*
b111 6
19
1>
1C
b111 G
#467200000000
0!
1"
0*
1+
09
1:
0>
0C
#467210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#467220000000
0!
0*
09
0>
0C
#467230000000
1!
1*
b1 6
19
1>
1C
b1 G
#467240000000
0!
0*
09
0>
0C
#467250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#467260000000
0!
0*
09
0>
0C
#467270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#467280000000
0!
0*
09
0>
0C
#467290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#467300000000
0!
0*
09
0>
0C
#467310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#467320000000
0!
0#
0*
0,
09
0>
0?
0C
#467330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#467340000000
0!
0*
09
0>
0C
#467350000000
1!
1*
19
1>
1C
#467360000000
0!
0*
09
0>
0C
#467370000000
1!
1*
19
1>
1C
#467380000000
0!
0*
09
0>
0C
#467390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#467400000000
0!
0*
09
0>
0C
#467410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#467420000000
0!
0*
09
0>
0C
#467430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#467440000000
0!
0*
09
0>
0C
#467450000000
1!
1*
b10 6
19
1>
1C
b10 G
#467460000000
0!
0*
09
0>
0C
#467470000000
1!
1*
b11 6
19
1>
1C
b11 G
#467480000000
0!
0*
09
0>
0C
#467490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#467500000000
0!
0*
09
0>
0C
#467510000000
1!
1*
b101 6
19
1>
1C
b101 G
#467520000000
0!
0*
09
0>
0C
#467530000000
1!
1*
b110 6
19
1>
1C
b110 G
#467540000000
0!
0*
09
0>
0C
#467550000000
1!
1*
b111 6
19
1>
1C
b111 G
#467560000000
0!
0*
09
0>
0C
#467570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#467580000000
0!
0*
09
0>
0C
#467590000000
1!
1*
b1 6
19
1>
1C
b1 G
#467600000000
0!
0*
09
0>
0C
#467610000000
1!
1*
b10 6
19
1>
1C
b10 G
#467620000000
0!
0*
09
0>
0C
#467630000000
1!
1*
b11 6
19
1>
1C
b11 G
#467640000000
0!
0*
09
0>
0C
#467650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#467660000000
0!
0*
09
0>
0C
#467670000000
1!
1*
b101 6
19
1>
1C
b101 G
#467680000000
0!
0*
09
0>
0C
#467690000000
1!
1*
b110 6
19
1>
1C
b110 G
#467700000000
0!
0*
09
0>
0C
#467710000000
1!
1*
b111 6
19
1>
1C
b111 G
#467720000000
0!
0*
09
0>
0C
#467730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#467740000000
0!
0*
09
0>
0C
#467750000000
1!
1*
b1 6
19
1>
1C
b1 G
#467760000000
0!
0*
09
0>
0C
#467770000000
1!
1*
b10 6
19
1>
1C
b10 G
#467780000000
0!
0*
09
0>
0C
#467790000000
1!
1*
b11 6
19
1>
1C
b11 G
#467800000000
0!
0*
09
0>
0C
#467810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#467820000000
0!
0*
09
0>
0C
#467830000000
1!
1*
b101 6
19
1>
1C
b101 G
#467840000000
0!
0*
09
0>
0C
#467850000000
1!
1*
b110 6
19
1>
1C
b110 G
#467860000000
0!
0*
09
0>
0C
#467870000000
1!
1*
b111 6
19
1>
1C
b111 G
#467880000000
0!
1"
0*
1+
09
1:
0>
0C
#467890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#467900000000
0!
0*
09
0>
0C
#467910000000
1!
1*
b1 6
19
1>
1C
b1 G
#467920000000
0!
0*
09
0>
0C
#467930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#467940000000
0!
0*
09
0>
0C
#467950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#467960000000
0!
0*
09
0>
0C
#467970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#467980000000
0!
0*
09
0>
0C
#467990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#468000000000
0!
0#
0*
0,
09
0>
0?
0C
#468010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#468020000000
0!
0*
09
0>
0C
#468030000000
1!
1*
19
1>
1C
#468040000000
0!
0*
09
0>
0C
#468050000000
1!
1*
19
1>
1C
#468060000000
0!
0*
09
0>
0C
#468070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#468080000000
0!
0*
09
0>
0C
#468090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#468100000000
0!
0*
09
0>
0C
#468110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#468120000000
0!
0*
09
0>
0C
#468130000000
1!
1*
b10 6
19
1>
1C
b10 G
#468140000000
0!
0*
09
0>
0C
#468150000000
1!
1*
b11 6
19
1>
1C
b11 G
#468160000000
0!
0*
09
0>
0C
#468170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#468180000000
0!
0*
09
0>
0C
#468190000000
1!
1*
b101 6
19
1>
1C
b101 G
#468200000000
0!
0*
09
0>
0C
#468210000000
1!
1*
b110 6
19
1>
1C
b110 G
#468220000000
0!
0*
09
0>
0C
#468230000000
1!
1*
b111 6
19
1>
1C
b111 G
#468240000000
0!
0*
09
0>
0C
#468250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#468260000000
0!
0*
09
0>
0C
#468270000000
1!
1*
b1 6
19
1>
1C
b1 G
#468280000000
0!
0*
09
0>
0C
#468290000000
1!
1*
b10 6
19
1>
1C
b10 G
#468300000000
0!
0*
09
0>
0C
#468310000000
1!
1*
b11 6
19
1>
1C
b11 G
#468320000000
0!
0*
09
0>
0C
#468330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#468340000000
0!
0*
09
0>
0C
#468350000000
1!
1*
b101 6
19
1>
1C
b101 G
#468360000000
0!
0*
09
0>
0C
#468370000000
1!
1*
b110 6
19
1>
1C
b110 G
#468380000000
0!
0*
09
0>
0C
#468390000000
1!
1*
b111 6
19
1>
1C
b111 G
#468400000000
0!
0*
09
0>
0C
#468410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#468420000000
0!
0*
09
0>
0C
#468430000000
1!
1*
b1 6
19
1>
1C
b1 G
#468440000000
0!
0*
09
0>
0C
#468450000000
1!
1*
b10 6
19
1>
1C
b10 G
#468460000000
0!
0*
09
0>
0C
#468470000000
1!
1*
b11 6
19
1>
1C
b11 G
#468480000000
0!
0*
09
0>
0C
#468490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#468500000000
0!
0*
09
0>
0C
#468510000000
1!
1*
b101 6
19
1>
1C
b101 G
#468520000000
0!
0*
09
0>
0C
#468530000000
1!
1*
b110 6
19
1>
1C
b110 G
#468540000000
0!
0*
09
0>
0C
#468550000000
1!
1*
b111 6
19
1>
1C
b111 G
#468560000000
0!
1"
0*
1+
09
1:
0>
0C
#468570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#468580000000
0!
0*
09
0>
0C
#468590000000
1!
1*
b1 6
19
1>
1C
b1 G
#468600000000
0!
0*
09
0>
0C
#468610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#468620000000
0!
0*
09
0>
0C
#468630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#468640000000
0!
0*
09
0>
0C
#468650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#468660000000
0!
0*
09
0>
0C
#468670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#468680000000
0!
0#
0*
0,
09
0>
0?
0C
#468690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#468700000000
0!
0*
09
0>
0C
#468710000000
1!
1*
19
1>
1C
#468720000000
0!
0*
09
0>
0C
#468730000000
1!
1*
19
1>
1C
#468740000000
0!
0*
09
0>
0C
#468750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#468760000000
0!
0*
09
0>
0C
#468770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#468780000000
0!
0*
09
0>
0C
#468790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#468800000000
0!
0*
09
0>
0C
#468810000000
1!
1*
b10 6
19
1>
1C
b10 G
#468820000000
0!
0*
09
0>
0C
#468830000000
1!
1*
b11 6
19
1>
1C
b11 G
#468840000000
0!
0*
09
0>
0C
#468850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#468860000000
0!
0*
09
0>
0C
#468870000000
1!
1*
b101 6
19
1>
1C
b101 G
#468880000000
0!
0*
09
0>
0C
#468890000000
1!
1*
b110 6
19
1>
1C
b110 G
#468900000000
0!
0*
09
0>
0C
#468910000000
1!
1*
b111 6
19
1>
1C
b111 G
#468920000000
0!
0*
09
0>
0C
#468930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#468940000000
0!
0*
09
0>
0C
#468950000000
1!
1*
b1 6
19
1>
1C
b1 G
#468960000000
0!
0*
09
0>
0C
#468970000000
1!
1*
b10 6
19
1>
1C
b10 G
#468980000000
0!
0*
09
0>
0C
#468990000000
1!
1*
b11 6
19
1>
1C
b11 G
#469000000000
0!
0*
09
0>
0C
#469010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#469020000000
0!
0*
09
0>
0C
#469030000000
1!
1*
b101 6
19
1>
1C
b101 G
#469040000000
0!
0*
09
0>
0C
#469050000000
1!
1*
b110 6
19
1>
1C
b110 G
#469060000000
0!
0*
09
0>
0C
#469070000000
1!
1*
b111 6
19
1>
1C
b111 G
#469080000000
0!
0*
09
0>
0C
#469090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#469100000000
0!
0*
09
0>
0C
#469110000000
1!
1*
b1 6
19
1>
1C
b1 G
#469120000000
0!
0*
09
0>
0C
#469130000000
1!
1*
b10 6
19
1>
1C
b10 G
#469140000000
0!
0*
09
0>
0C
#469150000000
1!
1*
b11 6
19
1>
1C
b11 G
#469160000000
0!
0*
09
0>
0C
#469170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#469180000000
0!
0*
09
0>
0C
#469190000000
1!
1*
b101 6
19
1>
1C
b101 G
#469200000000
0!
0*
09
0>
0C
#469210000000
1!
1*
b110 6
19
1>
1C
b110 G
#469220000000
0!
0*
09
0>
0C
#469230000000
1!
1*
b111 6
19
1>
1C
b111 G
#469240000000
0!
1"
0*
1+
09
1:
0>
0C
#469250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#469260000000
0!
0*
09
0>
0C
#469270000000
1!
1*
b1 6
19
1>
1C
b1 G
#469280000000
0!
0*
09
0>
0C
#469290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#469300000000
0!
0*
09
0>
0C
#469310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#469320000000
0!
0*
09
0>
0C
#469330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#469340000000
0!
0*
09
0>
0C
#469350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#469360000000
0!
0#
0*
0,
09
0>
0?
0C
#469370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#469380000000
0!
0*
09
0>
0C
#469390000000
1!
1*
19
1>
1C
#469400000000
0!
0*
09
0>
0C
#469410000000
1!
1*
19
1>
1C
#469420000000
0!
0*
09
0>
0C
#469430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#469440000000
0!
0*
09
0>
0C
#469450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#469460000000
0!
0*
09
0>
0C
#469470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#469480000000
0!
0*
09
0>
0C
#469490000000
1!
1*
b10 6
19
1>
1C
b10 G
#469500000000
0!
0*
09
0>
0C
#469510000000
1!
1*
b11 6
19
1>
1C
b11 G
#469520000000
0!
0*
09
0>
0C
#469530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#469540000000
0!
0*
09
0>
0C
#469550000000
1!
1*
b101 6
19
1>
1C
b101 G
#469560000000
0!
0*
09
0>
0C
#469570000000
1!
1*
b110 6
19
1>
1C
b110 G
#469580000000
0!
0*
09
0>
0C
#469590000000
1!
1*
b111 6
19
1>
1C
b111 G
#469600000000
0!
0*
09
0>
0C
#469610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#469620000000
0!
0*
09
0>
0C
#469630000000
1!
1*
b1 6
19
1>
1C
b1 G
#469640000000
0!
0*
09
0>
0C
#469650000000
1!
1*
b10 6
19
1>
1C
b10 G
#469660000000
0!
0*
09
0>
0C
#469670000000
1!
1*
b11 6
19
1>
1C
b11 G
#469680000000
0!
0*
09
0>
0C
#469690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#469700000000
0!
0*
09
0>
0C
#469710000000
1!
1*
b101 6
19
1>
1C
b101 G
#469720000000
0!
0*
09
0>
0C
#469730000000
1!
1*
b110 6
19
1>
1C
b110 G
#469740000000
0!
0*
09
0>
0C
#469750000000
1!
1*
b111 6
19
1>
1C
b111 G
#469760000000
0!
0*
09
0>
0C
#469770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#469780000000
0!
0*
09
0>
0C
#469790000000
1!
1*
b1 6
19
1>
1C
b1 G
#469800000000
0!
0*
09
0>
0C
#469810000000
1!
1*
b10 6
19
1>
1C
b10 G
#469820000000
0!
0*
09
0>
0C
#469830000000
1!
1*
b11 6
19
1>
1C
b11 G
#469840000000
0!
0*
09
0>
0C
#469850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#469860000000
0!
0*
09
0>
0C
#469870000000
1!
1*
b101 6
19
1>
1C
b101 G
#469880000000
0!
0*
09
0>
0C
#469890000000
1!
1*
b110 6
19
1>
1C
b110 G
#469900000000
0!
0*
09
0>
0C
#469910000000
1!
1*
b111 6
19
1>
1C
b111 G
#469920000000
0!
1"
0*
1+
09
1:
0>
0C
#469930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#469940000000
0!
0*
09
0>
0C
#469950000000
1!
1*
b1 6
19
1>
1C
b1 G
#469960000000
0!
0*
09
0>
0C
#469970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#469980000000
0!
0*
09
0>
0C
#469990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#470000000000
0!
0*
09
0>
0C
#470010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#470020000000
0!
0*
09
0>
0C
#470030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#470040000000
0!
0#
0*
0,
09
0>
0?
0C
#470050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#470060000000
0!
0*
09
0>
0C
#470070000000
1!
1*
19
1>
1C
#470080000000
0!
0*
09
0>
0C
#470090000000
1!
1*
19
1>
1C
#470100000000
0!
0*
09
0>
0C
#470110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#470120000000
0!
0*
09
0>
0C
#470130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#470140000000
0!
0*
09
0>
0C
#470150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#470160000000
0!
0*
09
0>
0C
#470170000000
1!
1*
b10 6
19
1>
1C
b10 G
#470180000000
0!
0*
09
0>
0C
#470190000000
1!
1*
b11 6
19
1>
1C
b11 G
#470200000000
0!
0*
09
0>
0C
#470210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#470220000000
0!
0*
09
0>
0C
#470230000000
1!
1*
b101 6
19
1>
1C
b101 G
#470240000000
0!
0*
09
0>
0C
#470250000000
1!
1*
b110 6
19
1>
1C
b110 G
#470260000000
0!
0*
09
0>
0C
#470270000000
1!
1*
b111 6
19
1>
1C
b111 G
#470280000000
0!
0*
09
0>
0C
#470290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#470300000000
0!
0*
09
0>
0C
#470310000000
1!
1*
b1 6
19
1>
1C
b1 G
#470320000000
0!
0*
09
0>
0C
#470330000000
1!
1*
b10 6
19
1>
1C
b10 G
#470340000000
0!
0*
09
0>
0C
#470350000000
1!
1*
b11 6
19
1>
1C
b11 G
#470360000000
0!
0*
09
0>
0C
#470370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#470380000000
0!
0*
09
0>
0C
#470390000000
1!
1*
b101 6
19
1>
1C
b101 G
#470400000000
0!
0*
09
0>
0C
#470410000000
1!
1*
b110 6
19
1>
1C
b110 G
#470420000000
0!
0*
09
0>
0C
#470430000000
1!
1*
b111 6
19
1>
1C
b111 G
#470440000000
0!
0*
09
0>
0C
#470450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#470460000000
0!
0*
09
0>
0C
#470470000000
1!
1*
b1 6
19
1>
1C
b1 G
#470480000000
0!
0*
09
0>
0C
#470490000000
1!
1*
b10 6
19
1>
1C
b10 G
#470500000000
0!
0*
09
0>
0C
#470510000000
1!
1*
b11 6
19
1>
1C
b11 G
#470520000000
0!
0*
09
0>
0C
#470530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#470540000000
0!
0*
09
0>
0C
#470550000000
1!
1*
b101 6
19
1>
1C
b101 G
#470560000000
0!
0*
09
0>
0C
#470570000000
1!
1*
b110 6
19
1>
1C
b110 G
#470580000000
0!
0*
09
0>
0C
#470590000000
1!
1*
b111 6
19
1>
1C
b111 G
#470600000000
0!
1"
0*
1+
09
1:
0>
0C
#470610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#470620000000
0!
0*
09
0>
0C
#470630000000
1!
1*
b1 6
19
1>
1C
b1 G
#470640000000
0!
0*
09
0>
0C
#470650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#470660000000
0!
0*
09
0>
0C
#470670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#470680000000
0!
0*
09
0>
0C
#470690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#470700000000
0!
0*
09
0>
0C
#470710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#470720000000
0!
0#
0*
0,
09
0>
0?
0C
#470730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#470740000000
0!
0*
09
0>
0C
#470750000000
1!
1*
19
1>
1C
#470760000000
0!
0*
09
0>
0C
#470770000000
1!
1*
19
1>
1C
#470780000000
0!
0*
09
0>
0C
#470790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#470800000000
0!
0*
09
0>
0C
#470810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#470820000000
0!
0*
09
0>
0C
#470830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#470840000000
0!
0*
09
0>
0C
#470850000000
1!
1*
b10 6
19
1>
1C
b10 G
#470860000000
0!
0*
09
0>
0C
#470870000000
1!
1*
b11 6
19
1>
1C
b11 G
#470880000000
0!
0*
09
0>
0C
#470890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#470900000000
0!
0*
09
0>
0C
#470910000000
1!
1*
b101 6
19
1>
1C
b101 G
#470920000000
0!
0*
09
0>
0C
#470930000000
1!
1*
b110 6
19
1>
1C
b110 G
#470940000000
0!
0*
09
0>
0C
#470950000000
1!
1*
b111 6
19
1>
1C
b111 G
#470960000000
0!
0*
09
0>
0C
#470970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#470980000000
0!
0*
09
0>
0C
#470990000000
1!
1*
b1 6
19
1>
1C
b1 G
#471000000000
0!
0*
09
0>
0C
#471010000000
1!
1*
b10 6
19
1>
1C
b10 G
#471020000000
0!
0*
09
0>
0C
#471030000000
1!
1*
b11 6
19
1>
1C
b11 G
#471040000000
0!
0*
09
0>
0C
#471050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#471060000000
0!
0*
09
0>
0C
#471070000000
1!
1*
b101 6
19
1>
1C
b101 G
#471080000000
0!
0*
09
0>
0C
#471090000000
1!
1*
b110 6
19
1>
1C
b110 G
#471100000000
0!
0*
09
0>
0C
#471110000000
1!
1*
b111 6
19
1>
1C
b111 G
#471120000000
0!
0*
09
0>
0C
#471130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#471140000000
0!
0*
09
0>
0C
#471150000000
1!
1*
b1 6
19
1>
1C
b1 G
#471160000000
0!
0*
09
0>
0C
#471170000000
1!
1*
b10 6
19
1>
1C
b10 G
#471180000000
0!
0*
09
0>
0C
#471190000000
1!
1*
b11 6
19
1>
1C
b11 G
#471200000000
0!
0*
09
0>
0C
#471210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#471220000000
0!
0*
09
0>
0C
#471230000000
1!
1*
b101 6
19
1>
1C
b101 G
#471240000000
0!
0*
09
0>
0C
#471250000000
1!
1*
b110 6
19
1>
1C
b110 G
#471260000000
0!
0*
09
0>
0C
#471270000000
1!
1*
b111 6
19
1>
1C
b111 G
#471280000000
0!
1"
0*
1+
09
1:
0>
0C
#471290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#471300000000
0!
0*
09
0>
0C
#471310000000
1!
1*
b1 6
19
1>
1C
b1 G
#471320000000
0!
0*
09
0>
0C
#471330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#471340000000
0!
0*
09
0>
0C
#471350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#471360000000
0!
0*
09
0>
0C
#471370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#471380000000
0!
0*
09
0>
0C
#471390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#471400000000
0!
0#
0*
0,
09
0>
0?
0C
#471410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#471420000000
0!
0*
09
0>
0C
#471430000000
1!
1*
19
1>
1C
#471440000000
0!
0*
09
0>
0C
#471450000000
1!
1*
19
1>
1C
#471460000000
0!
0*
09
0>
0C
#471470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#471480000000
0!
0*
09
0>
0C
#471490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#471500000000
0!
0*
09
0>
0C
#471510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#471520000000
0!
0*
09
0>
0C
#471530000000
1!
1*
b10 6
19
1>
1C
b10 G
#471540000000
0!
0*
09
0>
0C
#471550000000
1!
1*
b11 6
19
1>
1C
b11 G
#471560000000
0!
0*
09
0>
0C
#471570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#471580000000
0!
0*
09
0>
0C
#471590000000
1!
1*
b101 6
19
1>
1C
b101 G
#471600000000
0!
0*
09
0>
0C
#471610000000
1!
1*
b110 6
19
1>
1C
b110 G
#471620000000
0!
0*
09
0>
0C
#471630000000
1!
1*
b111 6
19
1>
1C
b111 G
#471640000000
0!
0*
09
0>
0C
#471650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#471660000000
0!
0*
09
0>
0C
#471670000000
1!
1*
b1 6
19
1>
1C
b1 G
#471680000000
0!
0*
09
0>
0C
#471690000000
1!
1*
b10 6
19
1>
1C
b10 G
#471700000000
0!
0*
09
0>
0C
#471710000000
1!
1*
b11 6
19
1>
1C
b11 G
#471720000000
0!
0*
09
0>
0C
#471730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#471740000000
0!
0*
09
0>
0C
#471750000000
1!
1*
b101 6
19
1>
1C
b101 G
#471760000000
0!
0*
09
0>
0C
#471770000000
1!
1*
b110 6
19
1>
1C
b110 G
#471780000000
0!
0*
09
0>
0C
#471790000000
1!
1*
b111 6
19
1>
1C
b111 G
#471800000000
0!
0*
09
0>
0C
#471810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#471820000000
0!
0*
09
0>
0C
#471830000000
1!
1*
b1 6
19
1>
1C
b1 G
#471840000000
0!
0*
09
0>
0C
#471850000000
1!
1*
b10 6
19
1>
1C
b10 G
#471860000000
0!
0*
09
0>
0C
#471870000000
1!
1*
b11 6
19
1>
1C
b11 G
#471880000000
0!
0*
09
0>
0C
#471890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#471900000000
0!
0*
09
0>
0C
#471910000000
1!
1*
b101 6
19
1>
1C
b101 G
#471920000000
0!
0*
09
0>
0C
#471930000000
1!
1*
b110 6
19
1>
1C
b110 G
#471940000000
0!
0*
09
0>
0C
#471950000000
1!
1*
b111 6
19
1>
1C
b111 G
#471960000000
0!
1"
0*
1+
09
1:
0>
0C
#471970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#471980000000
0!
0*
09
0>
0C
#471990000000
1!
1*
b1 6
19
1>
1C
b1 G
#472000000000
0!
0*
09
0>
0C
#472010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#472020000000
0!
0*
09
0>
0C
#472030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#472040000000
0!
0*
09
0>
0C
#472050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#472060000000
0!
0*
09
0>
0C
#472070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#472080000000
0!
0#
0*
0,
09
0>
0?
0C
#472090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#472100000000
0!
0*
09
0>
0C
#472110000000
1!
1*
19
1>
1C
#472120000000
0!
0*
09
0>
0C
#472130000000
1!
1*
19
1>
1C
#472140000000
0!
0*
09
0>
0C
#472150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#472160000000
0!
0*
09
0>
0C
#472170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#472180000000
0!
0*
09
0>
0C
#472190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#472200000000
0!
0*
09
0>
0C
#472210000000
1!
1*
b10 6
19
1>
1C
b10 G
#472220000000
0!
0*
09
0>
0C
#472230000000
1!
1*
b11 6
19
1>
1C
b11 G
#472240000000
0!
0*
09
0>
0C
#472250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#472260000000
0!
0*
09
0>
0C
#472270000000
1!
1*
b101 6
19
1>
1C
b101 G
#472280000000
0!
0*
09
0>
0C
#472290000000
1!
1*
b110 6
19
1>
1C
b110 G
#472300000000
0!
0*
09
0>
0C
#472310000000
1!
1*
b111 6
19
1>
1C
b111 G
#472320000000
0!
0*
09
0>
0C
#472330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#472340000000
0!
0*
09
0>
0C
#472350000000
1!
1*
b1 6
19
1>
1C
b1 G
#472360000000
0!
0*
09
0>
0C
#472370000000
1!
1*
b10 6
19
1>
1C
b10 G
#472380000000
0!
0*
09
0>
0C
#472390000000
1!
1*
b11 6
19
1>
1C
b11 G
#472400000000
0!
0*
09
0>
0C
#472410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#472420000000
0!
0*
09
0>
0C
#472430000000
1!
1*
b101 6
19
1>
1C
b101 G
#472440000000
0!
0*
09
0>
0C
#472450000000
1!
1*
b110 6
19
1>
1C
b110 G
#472460000000
0!
0*
09
0>
0C
#472470000000
1!
1*
b111 6
19
1>
1C
b111 G
#472480000000
0!
0*
09
0>
0C
#472490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#472500000000
0!
0*
09
0>
0C
#472510000000
1!
1*
b1 6
19
1>
1C
b1 G
#472520000000
0!
0*
09
0>
0C
#472530000000
1!
1*
b10 6
19
1>
1C
b10 G
#472540000000
0!
0*
09
0>
0C
#472550000000
1!
1*
b11 6
19
1>
1C
b11 G
#472560000000
0!
0*
09
0>
0C
#472570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#472580000000
0!
0*
09
0>
0C
#472590000000
1!
1*
b101 6
19
1>
1C
b101 G
#472600000000
0!
0*
09
0>
0C
#472610000000
1!
1*
b110 6
19
1>
1C
b110 G
#472620000000
0!
0*
09
0>
0C
#472630000000
1!
1*
b111 6
19
1>
1C
b111 G
#472640000000
0!
1"
0*
1+
09
1:
0>
0C
#472650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#472660000000
0!
0*
09
0>
0C
#472670000000
1!
1*
b1 6
19
1>
1C
b1 G
#472680000000
0!
0*
09
0>
0C
#472690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#472700000000
0!
0*
09
0>
0C
#472710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#472720000000
0!
0*
09
0>
0C
#472730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#472740000000
0!
0*
09
0>
0C
#472750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#472760000000
0!
0#
0*
0,
09
0>
0?
0C
#472770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#472780000000
0!
0*
09
0>
0C
#472790000000
1!
1*
19
1>
1C
#472800000000
0!
0*
09
0>
0C
#472810000000
1!
1*
19
1>
1C
#472820000000
0!
0*
09
0>
0C
#472830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#472840000000
0!
0*
09
0>
0C
#472850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#472860000000
0!
0*
09
0>
0C
#472870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#472880000000
0!
0*
09
0>
0C
#472890000000
1!
1*
b10 6
19
1>
1C
b10 G
#472900000000
0!
0*
09
0>
0C
#472910000000
1!
1*
b11 6
19
1>
1C
b11 G
#472920000000
0!
0*
09
0>
0C
#472930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#472940000000
0!
0*
09
0>
0C
#472950000000
1!
1*
b101 6
19
1>
1C
b101 G
#472960000000
0!
0*
09
0>
0C
#472970000000
1!
1*
b110 6
19
1>
1C
b110 G
#472980000000
0!
0*
09
0>
0C
#472990000000
1!
1*
b111 6
19
1>
1C
b111 G
#473000000000
0!
0*
09
0>
0C
#473010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#473020000000
0!
0*
09
0>
0C
#473030000000
1!
1*
b1 6
19
1>
1C
b1 G
#473040000000
0!
0*
09
0>
0C
#473050000000
1!
1*
b10 6
19
1>
1C
b10 G
#473060000000
0!
0*
09
0>
0C
#473070000000
1!
1*
b11 6
19
1>
1C
b11 G
#473080000000
0!
0*
09
0>
0C
#473090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#473100000000
0!
0*
09
0>
0C
#473110000000
1!
1*
b101 6
19
1>
1C
b101 G
#473120000000
0!
0*
09
0>
0C
#473130000000
1!
1*
b110 6
19
1>
1C
b110 G
#473140000000
0!
0*
09
0>
0C
#473150000000
1!
1*
b111 6
19
1>
1C
b111 G
#473160000000
0!
0*
09
0>
0C
#473170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#473180000000
0!
0*
09
0>
0C
#473190000000
1!
1*
b1 6
19
1>
1C
b1 G
#473200000000
0!
0*
09
0>
0C
#473210000000
1!
1*
b10 6
19
1>
1C
b10 G
#473220000000
0!
0*
09
0>
0C
#473230000000
1!
1*
b11 6
19
1>
1C
b11 G
#473240000000
0!
0*
09
0>
0C
#473250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#473260000000
0!
0*
09
0>
0C
#473270000000
1!
1*
b101 6
19
1>
1C
b101 G
#473280000000
0!
0*
09
0>
0C
#473290000000
1!
1*
b110 6
19
1>
1C
b110 G
#473300000000
0!
0*
09
0>
0C
#473310000000
1!
1*
b111 6
19
1>
1C
b111 G
#473320000000
0!
1"
0*
1+
09
1:
0>
0C
#473330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#473340000000
0!
0*
09
0>
0C
#473350000000
1!
1*
b1 6
19
1>
1C
b1 G
#473360000000
0!
0*
09
0>
0C
#473370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#473380000000
0!
0*
09
0>
0C
#473390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#473400000000
0!
0*
09
0>
0C
#473410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#473420000000
0!
0*
09
0>
0C
#473430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#473440000000
0!
0#
0*
0,
09
0>
0?
0C
#473450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#473460000000
0!
0*
09
0>
0C
#473470000000
1!
1*
19
1>
1C
#473480000000
0!
0*
09
0>
0C
#473490000000
1!
1*
19
1>
1C
#473500000000
0!
0*
09
0>
0C
#473510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#473520000000
0!
0*
09
0>
0C
#473530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#473540000000
0!
0*
09
0>
0C
#473550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#473560000000
0!
0*
09
0>
0C
#473570000000
1!
1*
b10 6
19
1>
1C
b10 G
#473580000000
0!
0*
09
0>
0C
#473590000000
1!
1*
b11 6
19
1>
1C
b11 G
#473600000000
0!
0*
09
0>
0C
#473610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#473620000000
0!
0*
09
0>
0C
#473630000000
1!
1*
b101 6
19
1>
1C
b101 G
#473640000000
0!
0*
09
0>
0C
#473650000000
1!
1*
b110 6
19
1>
1C
b110 G
#473660000000
0!
0*
09
0>
0C
#473670000000
1!
1*
b111 6
19
1>
1C
b111 G
#473680000000
0!
0*
09
0>
0C
#473690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#473700000000
0!
0*
09
0>
0C
#473710000000
1!
1*
b1 6
19
1>
1C
b1 G
#473720000000
0!
0*
09
0>
0C
#473730000000
1!
1*
b10 6
19
1>
1C
b10 G
#473740000000
0!
0*
09
0>
0C
#473750000000
1!
1*
b11 6
19
1>
1C
b11 G
#473760000000
0!
0*
09
0>
0C
#473770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#473780000000
0!
0*
09
0>
0C
#473790000000
1!
1*
b101 6
19
1>
1C
b101 G
#473800000000
0!
0*
09
0>
0C
#473810000000
1!
1*
b110 6
19
1>
1C
b110 G
#473820000000
0!
0*
09
0>
0C
#473830000000
1!
1*
b111 6
19
1>
1C
b111 G
#473840000000
0!
0*
09
0>
0C
#473850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#473860000000
0!
0*
09
0>
0C
#473870000000
1!
1*
b1 6
19
1>
1C
b1 G
#473880000000
0!
0*
09
0>
0C
#473890000000
1!
1*
b10 6
19
1>
1C
b10 G
#473900000000
0!
0*
09
0>
0C
#473910000000
1!
1*
b11 6
19
1>
1C
b11 G
#473920000000
0!
0*
09
0>
0C
#473930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#473940000000
0!
0*
09
0>
0C
#473950000000
1!
1*
b101 6
19
1>
1C
b101 G
#473960000000
0!
0*
09
0>
0C
#473970000000
1!
1*
b110 6
19
1>
1C
b110 G
#473980000000
0!
0*
09
0>
0C
#473990000000
1!
1*
b111 6
19
1>
1C
b111 G
#474000000000
0!
1"
0*
1+
09
1:
0>
0C
#474010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#474020000000
0!
0*
09
0>
0C
#474030000000
1!
1*
b1 6
19
1>
1C
b1 G
#474040000000
0!
0*
09
0>
0C
#474050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#474060000000
0!
0*
09
0>
0C
#474070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#474080000000
0!
0*
09
0>
0C
#474090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#474100000000
0!
0*
09
0>
0C
#474110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#474120000000
0!
0#
0*
0,
09
0>
0?
0C
#474130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#474140000000
0!
0*
09
0>
0C
#474150000000
1!
1*
19
1>
1C
#474160000000
0!
0*
09
0>
0C
#474170000000
1!
1*
19
1>
1C
#474180000000
0!
0*
09
0>
0C
#474190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#474200000000
0!
0*
09
0>
0C
#474210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#474220000000
0!
0*
09
0>
0C
#474230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#474240000000
0!
0*
09
0>
0C
#474250000000
1!
1*
b10 6
19
1>
1C
b10 G
#474260000000
0!
0*
09
0>
0C
#474270000000
1!
1*
b11 6
19
1>
1C
b11 G
#474280000000
0!
0*
09
0>
0C
#474290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#474300000000
0!
0*
09
0>
0C
#474310000000
1!
1*
b101 6
19
1>
1C
b101 G
#474320000000
0!
0*
09
0>
0C
#474330000000
1!
1*
b110 6
19
1>
1C
b110 G
#474340000000
0!
0*
09
0>
0C
#474350000000
1!
1*
b111 6
19
1>
1C
b111 G
#474360000000
0!
0*
09
0>
0C
#474370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#474380000000
0!
0*
09
0>
0C
#474390000000
1!
1*
b1 6
19
1>
1C
b1 G
#474400000000
0!
0*
09
0>
0C
#474410000000
1!
1*
b10 6
19
1>
1C
b10 G
#474420000000
0!
0*
09
0>
0C
#474430000000
1!
1*
b11 6
19
1>
1C
b11 G
#474440000000
0!
0*
09
0>
0C
#474450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#474460000000
0!
0*
09
0>
0C
#474470000000
1!
1*
b101 6
19
1>
1C
b101 G
#474480000000
0!
0*
09
0>
0C
#474490000000
1!
1*
b110 6
19
1>
1C
b110 G
#474500000000
0!
0*
09
0>
0C
#474510000000
1!
1*
b111 6
19
1>
1C
b111 G
#474520000000
0!
0*
09
0>
0C
#474530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#474540000000
0!
0*
09
0>
0C
#474550000000
1!
1*
b1 6
19
1>
1C
b1 G
#474560000000
0!
0*
09
0>
0C
#474570000000
1!
1*
b10 6
19
1>
1C
b10 G
#474580000000
0!
0*
09
0>
0C
#474590000000
1!
1*
b11 6
19
1>
1C
b11 G
#474600000000
0!
0*
09
0>
0C
#474610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#474620000000
0!
0*
09
0>
0C
#474630000000
1!
1*
b101 6
19
1>
1C
b101 G
#474640000000
0!
0*
09
0>
0C
#474650000000
1!
1*
b110 6
19
1>
1C
b110 G
#474660000000
0!
0*
09
0>
0C
#474670000000
1!
1*
b111 6
19
1>
1C
b111 G
#474680000000
0!
1"
0*
1+
09
1:
0>
0C
#474690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#474700000000
0!
0*
09
0>
0C
#474710000000
1!
1*
b1 6
19
1>
1C
b1 G
#474720000000
0!
0*
09
0>
0C
#474730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#474740000000
0!
0*
09
0>
0C
#474750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#474760000000
0!
0*
09
0>
0C
#474770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#474780000000
0!
0*
09
0>
0C
#474790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#474800000000
0!
0#
0*
0,
09
0>
0?
0C
#474810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#474820000000
0!
0*
09
0>
0C
#474830000000
1!
1*
19
1>
1C
#474840000000
0!
0*
09
0>
0C
#474850000000
1!
1*
19
1>
1C
#474860000000
0!
0*
09
0>
0C
#474870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#474880000000
0!
0*
09
0>
0C
#474890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#474900000000
0!
0*
09
0>
0C
#474910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#474920000000
0!
0*
09
0>
0C
#474930000000
1!
1*
b10 6
19
1>
1C
b10 G
#474940000000
0!
0*
09
0>
0C
#474950000000
1!
1*
b11 6
19
1>
1C
b11 G
#474960000000
0!
0*
09
0>
0C
#474970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#474980000000
0!
0*
09
0>
0C
#474990000000
1!
1*
b101 6
19
1>
1C
b101 G
#475000000000
0!
0*
09
0>
0C
#475010000000
1!
1*
b110 6
19
1>
1C
b110 G
#475020000000
0!
0*
09
0>
0C
#475030000000
1!
1*
b111 6
19
1>
1C
b111 G
#475040000000
0!
0*
09
0>
0C
#475050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#475060000000
0!
0*
09
0>
0C
#475070000000
1!
1*
b1 6
19
1>
1C
b1 G
#475080000000
0!
0*
09
0>
0C
#475090000000
1!
1*
b10 6
19
1>
1C
b10 G
#475100000000
0!
0*
09
0>
0C
#475110000000
1!
1*
b11 6
19
1>
1C
b11 G
#475120000000
0!
0*
09
0>
0C
#475130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#475140000000
0!
0*
09
0>
0C
#475150000000
1!
1*
b101 6
19
1>
1C
b101 G
#475160000000
0!
0*
09
0>
0C
#475170000000
1!
1*
b110 6
19
1>
1C
b110 G
#475180000000
0!
0*
09
0>
0C
#475190000000
1!
1*
b111 6
19
1>
1C
b111 G
#475200000000
0!
0*
09
0>
0C
#475210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#475220000000
0!
0*
09
0>
0C
#475230000000
1!
1*
b1 6
19
1>
1C
b1 G
#475240000000
0!
0*
09
0>
0C
#475250000000
1!
1*
b10 6
19
1>
1C
b10 G
#475260000000
0!
0*
09
0>
0C
#475270000000
1!
1*
b11 6
19
1>
1C
b11 G
#475280000000
0!
0*
09
0>
0C
#475290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#475300000000
0!
0*
09
0>
0C
#475310000000
1!
1*
b101 6
19
1>
1C
b101 G
#475320000000
0!
0*
09
0>
0C
#475330000000
1!
1*
b110 6
19
1>
1C
b110 G
#475340000000
0!
0*
09
0>
0C
#475350000000
1!
1*
b111 6
19
1>
1C
b111 G
#475360000000
0!
1"
0*
1+
09
1:
0>
0C
#475370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#475380000000
0!
0*
09
0>
0C
#475390000000
1!
1*
b1 6
19
1>
1C
b1 G
#475400000000
0!
0*
09
0>
0C
#475410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#475420000000
0!
0*
09
0>
0C
#475430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#475440000000
0!
0*
09
0>
0C
#475450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#475460000000
0!
0*
09
0>
0C
#475470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#475480000000
0!
0#
0*
0,
09
0>
0?
0C
#475490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#475500000000
0!
0*
09
0>
0C
#475510000000
1!
1*
19
1>
1C
#475520000000
0!
0*
09
0>
0C
#475530000000
1!
1*
19
1>
1C
#475540000000
0!
0*
09
0>
0C
#475550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#475560000000
0!
0*
09
0>
0C
#475570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#475580000000
0!
0*
09
0>
0C
#475590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#475600000000
0!
0*
09
0>
0C
#475610000000
1!
1*
b10 6
19
1>
1C
b10 G
#475620000000
0!
0*
09
0>
0C
#475630000000
1!
1*
b11 6
19
1>
1C
b11 G
#475640000000
0!
0*
09
0>
0C
#475650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#475660000000
0!
0*
09
0>
0C
#475670000000
1!
1*
b101 6
19
1>
1C
b101 G
#475680000000
0!
0*
09
0>
0C
#475690000000
1!
1*
b110 6
19
1>
1C
b110 G
#475700000000
0!
0*
09
0>
0C
#475710000000
1!
1*
b111 6
19
1>
1C
b111 G
#475720000000
0!
0*
09
0>
0C
#475730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#475740000000
0!
0*
09
0>
0C
#475750000000
1!
1*
b1 6
19
1>
1C
b1 G
#475760000000
0!
0*
09
0>
0C
#475770000000
1!
1*
b10 6
19
1>
1C
b10 G
#475780000000
0!
0*
09
0>
0C
#475790000000
1!
1*
b11 6
19
1>
1C
b11 G
#475800000000
0!
0*
09
0>
0C
#475810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#475820000000
0!
0*
09
0>
0C
#475830000000
1!
1*
b101 6
19
1>
1C
b101 G
#475840000000
0!
0*
09
0>
0C
#475850000000
1!
1*
b110 6
19
1>
1C
b110 G
#475860000000
0!
0*
09
0>
0C
#475870000000
1!
1*
b111 6
19
1>
1C
b111 G
#475880000000
0!
0*
09
0>
0C
#475890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#475900000000
0!
0*
09
0>
0C
#475910000000
1!
1*
b1 6
19
1>
1C
b1 G
#475920000000
0!
0*
09
0>
0C
#475930000000
1!
1*
b10 6
19
1>
1C
b10 G
#475940000000
0!
0*
09
0>
0C
#475950000000
1!
1*
b11 6
19
1>
1C
b11 G
#475960000000
0!
0*
09
0>
0C
#475970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#475980000000
0!
0*
09
0>
0C
#475990000000
1!
1*
b101 6
19
1>
1C
b101 G
#476000000000
0!
0*
09
0>
0C
#476010000000
1!
1*
b110 6
19
1>
1C
b110 G
#476020000000
0!
0*
09
0>
0C
#476030000000
1!
1*
b111 6
19
1>
1C
b111 G
#476040000000
0!
1"
0*
1+
09
1:
0>
0C
#476050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#476060000000
0!
0*
09
0>
0C
#476070000000
1!
1*
b1 6
19
1>
1C
b1 G
#476080000000
0!
0*
09
0>
0C
#476090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#476100000000
0!
0*
09
0>
0C
#476110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#476120000000
0!
0*
09
0>
0C
#476130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#476140000000
0!
0*
09
0>
0C
#476150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#476160000000
0!
0#
0*
0,
09
0>
0?
0C
#476170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#476180000000
0!
0*
09
0>
0C
#476190000000
1!
1*
19
1>
1C
#476200000000
0!
0*
09
0>
0C
#476210000000
1!
1*
19
1>
1C
#476220000000
0!
0*
09
0>
0C
#476230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#476240000000
0!
0*
09
0>
0C
#476250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#476260000000
0!
0*
09
0>
0C
#476270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#476280000000
0!
0*
09
0>
0C
#476290000000
1!
1*
b10 6
19
1>
1C
b10 G
#476300000000
0!
0*
09
0>
0C
#476310000000
1!
1*
b11 6
19
1>
1C
b11 G
#476320000000
0!
0*
09
0>
0C
#476330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#476340000000
0!
0*
09
0>
0C
#476350000000
1!
1*
b101 6
19
1>
1C
b101 G
#476360000000
0!
0*
09
0>
0C
#476370000000
1!
1*
b110 6
19
1>
1C
b110 G
#476380000000
0!
0*
09
0>
0C
#476390000000
1!
1*
b111 6
19
1>
1C
b111 G
#476400000000
0!
0*
09
0>
0C
#476410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#476420000000
0!
0*
09
0>
0C
#476430000000
1!
1*
b1 6
19
1>
1C
b1 G
#476440000000
0!
0*
09
0>
0C
#476450000000
1!
1*
b10 6
19
1>
1C
b10 G
#476460000000
0!
0*
09
0>
0C
#476470000000
1!
1*
b11 6
19
1>
1C
b11 G
#476480000000
0!
0*
09
0>
0C
#476490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#476500000000
0!
0*
09
0>
0C
#476510000000
1!
1*
b101 6
19
1>
1C
b101 G
#476520000000
0!
0*
09
0>
0C
#476530000000
1!
1*
b110 6
19
1>
1C
b110 G
#476540000000
0!
0*
09
0>
0C
#476550000000
1!
1*
b111 6
19
1>
1C
b111 G
#476560000000
0!
0*
09
0>
0C
#476570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#476580000000
0!
0*
09
0>
0C
#476590000000
1!
1*
b1 6
19
1>
1C
b1 G
#476600000000
0!
0*
09
0>
0C
#476610000000
1!
1*
b10 6
19
1>
1C
b10 G
#476620000000
0!
0*
09
0>
0C
#476630000000
1!
1*
b11 6
19
1>
1C
b11 G
#476640000000
0!
0*
09
0>
0C
#476650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#476660000000
0!
0*
09
0>
0C
#476670000000
1!
1*
b101 6
19
1>
1C
b101 G
#476680000000
0!
0*
09
0>
0C
#476690000000
1!
1*
b110 6
19
1>
1C
b110 G
#476700000000
0!
0*
09
0>
0C
#476710000000
1!
1*
b111 6
19
1>
1C
b111 G
#476720000000
0!
1"
0*
1+
09
1:
0>
0C
#476730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#476740000000
0!
0*
09
0>
0C
#476750000000
1!
1*
b1 6
19
1>
1C
b1 G
#476760000000
0!
0*
09
0>
0C
#476770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#476780000000
0!
0*
09
0>
0C
#476790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#476800000000
0!
0*
09
0>
0C
#476810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#476820000000
0!
0*
09
0>
0C
#476830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#476840000000
0!
0#
0*
0,
09
0>
0?
0C
#476850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#476860000000
0!
0*
09
0>
0C
#476870000000
1!
1*
19
1>
1C
#476880000000
0!
0*
09
0>
0C
#476890000000
1!
1*
19
1>
1C
#476900000000
0!
0*
09
0>
0C
#476910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#476920000000
0!
0*
09
0>
0C
#476930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#476940000000
0!
0*
09
0>
0C
#476950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#476960000000
0!
0*
09
0>
0C
#476970000000
1!
1*
b10 6
19
1>
1C
b10 G
#476980000000
0!
0*
09
0>
0C
#476990000000
1!
1*
b11 6
19
1>
1C
b11 G
#477000000000
0!
0*
09
0>
0C
#477010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#477020000000
0!
0*
09
0>
0C
#477030000000
1!
1*
b101 6
19
1>
1C
b101 G
#477040000000
0!
0*
09
0>
0C
#477050000000
1!
1*
b110 6
19
1>
1C
b110 G
#477060000000
0!
0*
09
0>
0C
#477070000000
1!
1*
b111 6
19
1>
1C
b111 G
#477080000000
0!
0*
09
0>
0C
#477090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#477100000000
0!
0*
09
0>
0C
#477110000000
1!
1*
b1 6
19
1>
1C
b1 G
#477120000000
0!
0*
09
0>
0C
#477130000000
1!
1*
b10 6
19
1>
1C
b10 G
#477140000000
0!
0*
09
0>
0C
#477150000000
1!
1*
b11 6
19
1>
1C
b11 G
#477160000000
0!
0*
09
0>
0C
#477170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#477180000000
0!
0*
09
0>
0C
#477190000000
1!
1*
b101 6
19
1>
1C
b101 G
#477200000000
0!
0*
09
0>
0C
#477210000000
1!
1*
b110 6
19
1>
1C
b110 G
#477220000000
0!
0*
09
0>
0C
#477230000000
1!
1*
b111 6
19
1>
1C
b111 G
#477240000000
0!
0*
09
0>
0C
#477250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#477260000000
0!
0*
09
0>
0C
#477270000000
1!
1*
b1 6
19
1>
1C
b1 G
#477280000000
0!
0*
09
0>
0C
#477290000000
1!
1*
b10 6
19
1>
1C
b10 G
#477300000000
0!
0*
09
0>
0C
#477310000000
1!
1*
b11 6
19
1>
1C
b11 G
#477320000000
0!
0*
09
0>
0C
#477330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#477340000000
0!
0*
09
0>
0C
#477350000000
1!
1*
b101 6
19
1>
1C
b101 G
#477360000000
0!
0*
09
0>
0C
#477370000000
1!
1*
b110 6
19
1>
1C
b110 G
#477380000000
0!
0*
09
0>
0C
#477390000000
1!
1*
b111 6
19
1>
1C
b111 G
#477400000000
0!
1"
0*
1+
09
1:
0>
0C
#477410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#477420000000
0!
0*
09
0>
0C
#477430000000
1!
1*
b1 6
19
1>
1C
b1 G
#477440000000
0!
0*
09
0>
0C
#477450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#477460000000
0!
0*
09
0>
0C
#477470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#477480000000
0!
0*
09
0>
0C
#477490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#477500000000
0!
0*
09
0>
0C
#477510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#477520000000
0!
0#
0*
0,
09
0>
0?
0C
#477530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#477540000000
0!
0*
09
0>
0C
#477550000000
1!
1*
19
1>
1C
#477560000000
0!
0*
09
0>
0C
#477570000000
1!
1*
19
1>
1C
#477580000000
0!
0*
09
0>
0C
#477590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#477600000000
0!
0*
09
0>
0C
#477610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#477620000000
0!
0*
09
0>
0C
#477630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#477640000000
0!
0*
09
0>
0C
#477650000000
1!
1*
b10 6
19
1>
1C
b10 G
#477660000000
0!
0*
09
0>
0C
#477670000000
1!
1*
b11 6
19
1>
1C
b11 G
#477680000000
0!
0*
09
0>
0C
#477690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#477700000000
0!
0*
09
0>
0C
#477710000000
1!
1*
b101 6
19
1>
1C
b101 G
#477720000000
0!
0*
09
0>
0C
#477730000000
1!
1*
b110 6
19
1>
1C
b110 G
#477740000000
0!
0*
09
0>
0C
#477750000000
1!
1*
b111 6
19
1>
1C
b111 G
#477760000000
0!
0*
09
0>
0C
#477770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#477780000000
0!
0*
09
0>
0C
#477790000000
1!
1*
b1 6
19
1>
1C
b1 G
#477800000000
0!
0*
09
0>
0C
#477810000000
1!
1*
b10 6
19
1>
1C
b10 G
#477820000000
0!
0*
09
0>
0C
#477830000000
1!
1*
b11 6
19
1>
1C
b11 G
#477840000000
0!
0*
09
0>
0C
#477850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#477860000000
0!
0*
09
0>
0C
#477870000000
1!
1*
b101 6
19
1>
1C
b101 G
#477880000000
0!
0*
09
0>
0C
#477890000000
1!
1*
b110 6
19
1>
1C
b110 G
#477900000000
0!
0*
09
0>
0C
#477910000000
1!
1*
b111 6
19
1>
1C
b111 G
#477920000000
0!
0*
09
0>
0C
#477930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#477940000000
0!
0*
09
0>
0C
#477950000000
1!
1*
b1 6
19
1>
1C
b1 G
#477960000000
0!
0*
09
0>
0C
#477970000000
1!
1*
b10 6
19
1>
1C
b10 G
#477980000000
0!
0*
09
0>
0C
#477990000000
1!
1*
b11 6
19
1>
1C
b11 G
#478000000000
0!
0*
09
0>
0C
#478010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#478020000000
0!
0*
09
0>
0C
#478030000000
1!
1*
b101 6
19
1>
1C
b101 G
#478040000000
0!
0*
09
0>
0C
#478050000000
1!
1*
b110 6
19
1>
1C
b110 G
#478060000000
0!
0*
09
0>
0C
#478070000000
1!
1*
b111 6
19
1>
1C
b111 G
#478080000000
0!
1"
0*
1+
09
1:
0>
0C
#478090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#478100000000
0!
0*
09
0>
0C
#478110000000
1!
1*
b1 6
19
1>
1C
b1 G
#478120000000
0!
0*
09
0>
0C
#478130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#478140000000
0!
0*
09
0>
0C
#478150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#478160000000
0!
0*
09
0>
0C
#478170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#478180000000
0!
0*
09
0>
0C
#478190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#478200000000
0!
0#
0*
0,
09
0>
0?
0C
#478210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#478220000000
0!
0*
09
0>
0C
#478230000000
1!
1*
19
1>
1C
#478240000000
0!
0*
09
0>
0C
#478250000000
1!
1*
19
1>
1C
#478260000000
0!
0*
09
0>
0C
#478270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#478280000000
0!
0*
09
0>
0C
#478290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#478300000000
0!
0*
09
0>
0C
#478310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#478320000000
0!
0*
09
0>
0C
#478330000000
1!
1*
b10 6
19
1>
1C
b10 G
#478340000000
0!
0*
09
0>
0C
#478350000000
1!
1*
b11 6
19
1>
1C
b11 G
#478360000000
0!
0*
09
0>
0C
#478370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#478380000000
0!
0*
09
0>
0C
#478390000000
1!
1*
b101 6
19
1>
1C
b101 G
#478400000000
0!
0*
09
0>
0C
#478410000000
1!
1*
b110 6
19
1>
1C
b110 G
#478420000000
0!
0*
09
0>
0C
#478430000000
1!
1*
b111 6
19
1>
1C
b111 G
#478440000000
0!
0*
09
0>
0C
#478450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#478460000000
0!
0*
09
0>
0C
#478470000000
1!
1*
b1 6
19
1>
1C
b1 G
#478480000000
0!
0*
09
0>
0C
#478490000000
1!
1*
b10 6
19
1>
1C
b10 G
#478500000000
0!
0*
09
0>
0C
#478510000000
1!
1*
b11 6
19
1>
1C
b11 G
#478520000000
0!
0*
09
0>
0C
#478530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#478540000000
0!
0*
09
0>
0C
#478550000000
1!
1*
b101 6
19
1>
1C
b101 G
#478560000000
0!
0*
09
0>
0C
#478570000000
1!
1*
b110 6
19
1>
1C
b110 G
#478580000000
0!
0*
09
0>
0C
#478590000000
1!
1*
b111 6
19
1>
1C
b111 G
#478600000000
0!
0*
09
0>
0C
#478610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#478620000000
0!
0*
09
0>
0C
#478630000000
1!
1*
b1 6
19
1>
1C
b1 G
#478640000000
0!
0*
09
0>
0C
#478650000000
1!
1*
b10 6
19
1>
1C
b10 G
#478660000000
0!
0*
09
0>
0C
#478670000000
1!
1*
b11 6
19
1>
1C
b11 G
#478680000000
0!
0*
09
0>
0C
#478690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#478700000000
0!
0*
09
0>
0C
#478710000000
1!
1*
b101 6
19
1>
1C
b101 G
#478720000000
0!
0*
09
0>
0C
#478730000000
1!
1*
b110 6
19
1>
1C
b110 G
#478740000000
0!
0*
09
0>
0C
#478750000000
1!
1*
b111 6
19
1>
1C
b111 G
#478760000000
0!
1"
0*
1+
09
1:
0>
0C
#478770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#478780000000
0!
0*
09
0>
0C
#478790000000
1!
1*
b1 6
19
1>
1C
b1 G
#478800000000
0!
0*
09
0>
0C
#478810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#478820000000
0!
0*
09
0>
0C
#478830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#478840000000
0!
0*
09
0>
0C
#478850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#478860000000
0!
0*
09
0>
0C
#478870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#478880000000
0!
0#
0*
0,
09
0>
0?
0C
#478890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#478900000000
0!
0*
09
0>
0C
#478910000000
1!
1*
19
1>
1C
#478920000000
0!
0*
09
0>
0C
#478930000000
1!
1*
19
1>
1C
#478940000000
0!
0*
09
0>
0C
#478950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#478960000000
0!
0*
09
0>
0C
#478970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#478980000000
0!
0*
09
0>
0C
#478990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#479000000000
0!
0*
09
0>
0C
#479010000000
1!
1*
b10 6
19
1>
1C
b10 G
#479020000000
0!
0*
09
0>
0C
#479030000000
1!
1*
b11 6
19
1>
1C
b11 G
#479040000000
0!
0*
09
0>
0C
#479050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#479060000000
0!
0*
09
0>
0C
#479070000000
1!
1*
b101 6
19
1>
1C
b101 G
#479080000000
0!
0*
09
0>
0C
#479090000000
1!
1*
b110 6
19
1>
1C
b110 G
#479100000000
0!
0*
09
0>
0C
#479110000000
1!
1*
b111 6
19
1>
1C
b111 G
#479120000000
0!
0*
09
0>
0C
#479130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#479140000000
0!
0*
09
0>
0C
#479150000000
1!
1*
b1 6
19
1>
1C
b1 G
#479160000000
0!
0*
09
0>
0C
#479170000000
1!
1*
b10 6
19
1>
1C
b10 G
#479180000000
0!
0*
09
0>
0C
#479190000000
1!
1*
b11 6
19
1>
1C
b11 G
#479200000000
0!
0*
09
0>
0C
#479210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#479220000000
0!
0*
09
0>
0C
#479230000000
1!
1*
b101 6
19
1>
1C
b101 G
#479240000000
0!
0*
09
0>
0C
#479250000000
1!
1*
b110 6
19
1>
1C
b110 G
#479260000000
0!
0*
09
0>
0C
#479270000000
1!
1*
b111 6
19
1>
1C
b111 G
#479280000000
0!
0*
09
0>
0C
#479290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#479300000000
0!
0*
09
0>
0C
#479310000000
1!
1*
b1 6
19
1>
1C
b1 G
#479320000000
0!
0*
09
0>
0C
#479330000000
1!
1*
b10 6
19
1>
1C
b10 G
#479340000000
0!
0*
09
0>
0C
#479350000000
1!
1*
b11 6
19
1>
1C
b11 G
#479360000000
0!
0*
09
0>
0C
#479370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#479380000000
0!
0*
09
0>
0C
#479390000000
1!
1*
b101 6
19
1>
1C
b101 G
#479400000000
0!
0*
09
0>
0C
#479410000000
1!
1*
b110 6
19
1>
1C
b110 G
#479420000000
0!
0*
09
0>
0C
#479430000000
1!
1*
b111 6
19
1>
1C
b111 G
#479440000000
0!
1"
0*
1+
09
1:
0>
0C
#479450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#479460000000
0!
0*
09
0>
0C
#479470000000
1!
1*
b1 6
19
1>
1C
b1 G
#479480000000
0!
0*
09
0>
0C
#479490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#479500000000
0!
0*
09
0>
0C
#479510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#479520000000
0!
0*
09
0>
0C
#479530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#479540000000
0!
0*
09
0>
0C
#479550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#479560000000
0!
0#
0*
0,
09
0>
0?
0C
#479570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#479580000000
0!
0*
09
0>
0C
#479590000000
1!
1*
19
1>
1C
#479600000000
0!
0*
09
0>
0C
#479610000000
1!
1*
19
1>
1C
#479620000000
0!
0*
09
0>
0C
#479630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#479640000000
0!
0*
09
0>
0C
#479650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#479660000000
0!
0*
09
0>
0C
#479670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#479680000000
0!
0*
09
0>
0C
#479690000000
1!
1*
b10 6
19
1>
1C
b10 G
#479700000000
0!
0*
09
0>
0C
#479710000000
1!
1*
b11 6
19
1>
1C
b11 G
#479720000000
0!
0*
09
0>
0C
#479730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#479740000000
0!
0*
09
0>
0C
#479750000000
1!
1*
b101 6
19
1>
1C
b101 G
#479760000000
0!
0*
09
0>
0C
#479770000000
1!
1*
b110 6
19
1>
1C
b110 G
#479780000000
0!
0*
09
0>
0C
#479790000000
1!
1*
b111 6
19
1>
1C
b111 G
#479800000000
0!
0*
09
0>
0C
#479810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#479820000000
0!
0*
09
0>
0C
#479830000000
1!
1*
b1 6
19
1>
1C
b1 G
#479840000000
0!
0*
09
0>
0C
#479850000000
1!
1*
b10 6
19
1>
1C
b10 G
#479860000000
0!
0*
09
0>
0C
#479870000000
1!
1*
b11 6
19
1>
1C
b11 G
#479880000000
0!
0*
09
0>
0C
#479890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#479900000000
0!
0*
09
0>
0C
#479910000000
1!
1*
b101 6
19
1>
1C
b101 G
#479920000000
0!
0*
09
0>
0C
#479930000000
1!
1*
b110 6
19
1>
1C
b110 G
#479940000000
0!
0*
09
0>
0C
#479950000000
1!
1*
b111 6
19
1>
1C
b111 G
#479960000000
0!
0*
09
0>
0C
#479970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#479980000000
0!
0*
09
0>
0C
#479990000000
1!
1*
b1 6
19
1>
1C
b1 G
#480000000000
0!
0*
09
0>
0C
#480010000000
1!
1*
b10 6
19
1>
1C
b10 G
#480020000000
0!
0*
09
0>
0C
#480030000000
1!
1*
b11 6
19
1>
1C
b11 G
#480040000000
0!
0*
09
0>
0C
#480050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#480060000000
0!
0*
09
0>
0C
#480070000000
1!
1*
b101 6
19
1>
1C
b101 G
#480080000000
0!
0*
09
0>
0C
#480090000000
1!
1*
b110 6
19
1>
1C
b110 G
#480100000000
0!
0*
09
0>
0C
#480110000000
1!
1*
b111 6
19
1>
1C
b111 G
#480120000000
0!
1"
0*
1+
09
1:
0>
0C
#480130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#480140000000
0!
0*
09
0>
0C
#480150000000
1!
1*
b1 6
19
1>
1C
b1 G
#480160000000
0!
0*
09
0>
0C
#480170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#480180000000
0!
0*
09
0>
0C
#480190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#480200000000
0!
0*
09
0>
0C
#480210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#480220000000
0!
0*
09
0>
0C
#480230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#480240000000
0!
0#
0*
0,
09
0>
0?
0C
#480250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#480260000000
0!
0*
09
0>
0C
#480270000000
1!
1*
19
1>
1C
#480280000000
0!
0*
09
0>
0C
#480290000000
1!
1*
19
1>
1C
#480300000000
0!
0*
09
0>
0C
#480310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#480320000000
0!
0*
09
0>
0C
#480330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#480340000000
0!
0*
09
0>
0C
#480350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#480360000000
0!
0*
09
0>
0C
#480370000000
1!
1*
b10 6
19
1>
1C
b10 G
#480380000000
0!
0*
09
0>
0C
#480390000000
1!
1*
b11 6
19
1>
1C
b11 G
#480400000000
0!
0*
09
0>
0C
#480410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#480420000000
0!
0*
09
0>
0C
#480430000000
1!
1*
b101 6
19
1>
1C
b101 G
#480440000000
0!
0*
09
0>
0C
#480450000000
1!
1*
b110 6
19
1>
1C
b110 G
#480460000000
0!
0*
09
0>
0C
#480470000000
1!
1*
b111 6
19
1>
1C
b111 G
#480480000000
0!
0*
09
0>
0C
#480490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#480500000000
0!
0*
09
0>
0C
#480510000000
1!
1*
b1 6
19
1>
1C
b1 G
#480520000000
0!
0*
09
0>
0C
#480530000000
1!
1*
b10 6
19
1>
1C
b10 G
#480540000000
0!
0*
09
0>
0C
#480550000000
1!
1*
b11 6
19
1>
1C
b11 G
#480560000000
0!
0*
09
0>
0C
#480570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#480580000000
0!
0*
09
0>
0C
#480590000000
1!
1*
b101 6
19
1>
1C
b101 G
#480600000000
0!
0*
09
0>
0C
#480610000000
1!
1*
b110 6
19
1>
1C
b110 G
#480620000000
0!
0*
09
0>
0C
#480630000000
1!
1*
b111 6
19
1>
1C
b111 G
#480640000000
0!
0*
09
0>
0C
#480650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#480660000000
0!
0*
09
0>
0C
#480670000000
1!
1*
b1 6
19
1>
1C
b1 G
#480680000000
0!
0*
09
0>
0C
#480690000000
1!
1*
b10 6
19
1>
1C
b10 G
#480700000000
0!
0*
09
0>
0C
#480710000000
1!
1*
b11 6
19
1>
1C
b11 G
#480720000000
0!
0*
09
0>
0C
#480730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#480740000000
0!
0*
09
0>
0C
#480750000000
1!
1*
b101 6
19
1>
1C
b101 G
#480760000000
0!
0*
09
0>
0C
#480770000000
1!
1*
b110 6
19
1>
1C
b110 G
#480780000000
0!
0*
09
0>
0C
#480790000000
1!
1*
b111 6
19
1>
1C
b111 G
#480800000000
0!
1"
0*
1+
09
1:
0>
0C
#480810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#480820000000
0!
0*
09
0>
0C
#480830000000
1!
1*
b1 6
19
1>
1C
b1 G
#480840000000
0!
0*
09
0>
0C
#480850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#480860000000
0!
0*
09
0>
0C
#480870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#480880000000
0!
0*
09
0>
0C
#480890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#480900000000
0!
0*
09
0>
0C
#480910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#480920000000
0!
0#
0*
0,
09
0>
0?
0C
#480930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#480940000000
0!
0*
09
0>
0C
#480950000000
1!
1*
19
1>
1C
#480960000000
0!
0*
09
0>
0C
#480970000000
1!
1*
19
1>
1C
#480980000000
0!
0*
09
0>
0C
#480990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#481000000000
0!
0*
09
0>
0C
#481010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#481020000000
0!
0*
09
0>
0C
#481030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#481040000000
0!
0*
09
0>
0C
#481050000000
1!
1*
b10 6
19
1>
1C
b10 G
#481060000000
0!
0*
09
0>
0C
#481070000000
1!
1*
b11 6
19
1>
1C
b11 G
#481080000000
0!
0*
09
0>
0C
#481090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#481100000000
0!
0*
09
0>
0C
#481110000000
1!
1*
b101 6
19
1>
1C
b101 G
#481120000000
0!
0*
09
0>
0C
#481130000000
1!
1*
b110 6
19
1>
1C
b110 G
#481140000000
0!
0*
09
0>
0C
#481150000000
1!
1*
b111 6
19
1>
1C
b111 G
#481160000000
0!
0*
09
0>
0C
#481170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#481180000000
0!
0*
09
0>
0C
#481190000000
1!
1*
b1 6
19
1>
1C
b1 G
#481200000000
0!
0*
09
0>
0C
#481210000000
1!
1*
b10 6
19
1>
1C
b10 G
#481220000000
0!
0*
09
0>
0C
#481230000000
1!
1*
b11 6
19
1>
1C
b11 G
#481240000000
0!
0*
09
0>
0C
#481250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#481260000000
0!
0*
09
0>
0C
#481270000000
1!
1*
b101 6
19
1>
1C
b101 G
#481280000000
0!
0*
09
0>
0C
#481290000000
1!
1*
b110 6
19
1>
1C
b110 G
#481300000000
0!
0*
09
0>
0C
#481310000000
1!
1*
b111 6
19
1>
1C
b111 G
#481320000000
0!
0*
09
0>
0C
#481330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#481340000000
0!
0*
09
0>
0C
#481350000000
1!
1*
b1 6
19
1>
1C
b1 G
#481360000000
0!
0*
09
0>
0C
#481370000000
1!
1*
b10 6
19
1>
1C
b10 G
#481380000000
0!
0*
09
0>
0C
#481390000000
1!
1*
b11 6
19
1>
1C
b11 G
#481400000000
0!
0*
09
0>
0C
#481410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#481420000000
0!
0*
09
0>
0C
#481430000000
1!
1*
b101 6
19
1>
1C
b101 G
#481440000000
0!
0*
09
0>
0C
#481450000000
1!
1*
b110 6
19
1>
1C
b110 G
#481460000000
0!
0*
09
0>
0C
#481470000000
1!
1*
b111 6
19
1>
1C
b111 G
#481480000000
0!
1"
0*
1+
09
1:
0>
0C
#481490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#481500000000
0!
0*
09
0>
0C
#481510000000
1!
1*
b1 6
19
1>
1C
b1 G
#481520000000
0!
0*
09
0>
0C
#481530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#481540000000
0!
0*
09
0>
0C
#481550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#481560000000
0!
0*
09
0>
0C
#481570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#481580000000
0!
0*
09
0>
0C
#481590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#481600000000
0!
0#
0*
0,
09
0>
0?
0C
#481610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#481620000000
0!
0*
09
0>
0C
#481630000000
1!
1*
19
1>
1C
#481640000000
0!
0*
09
0>
0C
#481650000000
1!
1*
19
1>
1C
#481660000000
0!
0*
09
0>
0C
#481670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#481680000000
0!
0*
09
0>
0C
#481690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#481700000000
0!
0*
09
0>
0C
#481710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#481720000000
0!
0*
09
0>
0C
#481730000000
1!
1*
b10 6
19
1>
1C
b10 G
#481740000000
0!
0*
09
0>
0C
#481750000000
1!
1*
b11 6
19
1>
1C
b11 G
#481760000000
0!
0*
09
0>
0C
#481770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#481780000000
0!
0*
09
0>
0C
#481790000000
1!
1*
b101 6
19
1>
1C
b101 G
#481800000000
0!
0*
09
0>
0C
#481810000000
1!
1*
b110 6
19
1>
1C
b110 G
#481820000000
0!
0*
09
0>
0C
#481830000000
1!
1*
b111 6
19
1>
1C
b111 G
#481840000000
0!
0*
09
0>
0C
#481850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#481860000000
0!
0*
09
0>
0C
#481870000000
1!
1*
b1 6
19
1>
1C
b1 G
#481880000000
0!
0*
09
0>
0C
#481890000000
1!
1*
b10 6
19
1>
1C
b10 G
#481900000000
0!
0*
09
0>
0C
#481910000000
1!
1*
b11 6
19
1>
1C
b11 G
#481920000000
0!
0*
09
0>
0C
#481930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#481940000000
0!
0*
09
0>
0C
#481950000000
1!
1*
b101 6
19
1>
1C
b101 G
#481960000000
0!
0*
09
0>
0C
#481970000000
1!
1*
b110 6
19
1>
1C
b110 G
#481980000000
0!
0*
09
0>
0C
#481990000000
1!
1*
b111 6
19
1>
1C
b111 G
#482000000000
0!
0*
09
0>
0C
#482010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#482020000000
0!
0*
09
0>
0C
#482030000000
1!
1*
b1 6
19
1>
1C
b1 G
#482040000000
0!
0*
09
0>
0C
#482050000000
1!
1*
b10 6
19
1>
1C
b10 G
#482060000000
0!
0*
09
0>
0C
#482070000000
1!
1*
b11 6
19
1>
1C
b11 G
#482080000000
0!
0*
09
0>
0C
#482090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#482100000000
0!
0*
09
0>
0C
#482110000000
1!
1*
b101 6
19
1>
1C
b101 G
#482120000000
0!
0*
09
0>
0C
#482130000000
1!
1*
b110 6
19
1>
1C
b110 G
#482140000000
0!
0*
09
0>
0C
#482150000000
1!
1*
b111 6
19
1>
1C
b111 G
#482160000000
0!
1"
0*
1+
09
1:
0>
0C
#482170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#482180000000
0!
0*
09
0>
0C
#482190000000
1!
1*
b1 6
19
1>
1C
b1 G
#482200000000
0!
0*
09
0>
0C
#482210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#482220000000
0!
0*
09
0>
0C
#482230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#482240000000
0!
0*
09
0>
0C
#482250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#482260000000
0!
0*
09
0>
0C
#482270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#482280000000
0!
0#
0*
0,
09
0>
0?
0C
#482290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#482300000000
0!
0*
09
0>
0C
#482310000000
1!
1*
19
1>
1C
#482320000000
0!
0*
09
0>
0C
#482330000000
1!
1*
19
1>
1C
#482340000000
0!
0*
09
0>
0C
#482350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#482360000000
0!
0*
09
0>
0C
#482370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#482380000000
0!
0*
09
0>
0C
#482390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#482400000000
0!
0*
09
0>
0C
#482410000000
1!
1*
b10 6
19
1>
1C
b10 G
#482420000000
0!
0*
09
0>
0C
#482430000000
1!
1*
b11 6
19
1>
1C
b11 G
#482440000000
0!
0*
09
0>
0C
#482450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#482460000000
0!
0*
09
0>
0C
#482470000000
1!
1*
b101 6
19
1>
1C
b101 G
#482480000000
0!
0*
09
0>
0C
#482490000000
1!
1*
b110 6
19
1>
1C
b110 G
#482500000000
0!
0*
09
0>
0C
#482510000000
1!
1*
b111 6
19
1>
1C
b111 G
#482520000000
0!
0*
09
0>
0C
#482530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#482540000000
0!
0*
09
0>
0C
#482550000000
1!
1*
b1 6
19
1>
1C
b1 G
#482560000000
0!
0*
09
0>
0C
#482570000000
1!
1*
b10 6
19
1>
1C
b10 G
#482580000000
0!
0*
09
0>
0C
#482590000000
1!
1*
b11 6
19
1>
1C
b11 G
#482600000000
0!
0*
09
0>
0C
#482610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#482620000000
0!
0*
09
0>
0C
#482630000000
1!
1*
b101 6
19
1>
1C
b101 G
#482640000000
0!
0*
09
0>
0C
#482650000000
1!
1*
b110 6
19
1>
1C
b110 G
#482660000000
0!
0*
09
0>
0C
#482670000000
1!
1*
b111 6
19
1>
1C
b111 G
#482680000000
0!
0*
09
0>
0C
#482690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#482700000000
0!
0*
09
0>
0C
#482710000000
1!
1*
b1 6
19
1>
1C
b1 G
#482720000000
0!
0*
09
0>
0C
#482730000000
1!
1*
b10 6
19
1>
1C
b10 G
#482740000000
0!
0*
09
0>
0C
#482750000000
1!
1*
b11 6
19
1>
1C
b11 G
#482760000000
0!
0*
09
0>
0C
#482770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#482780000000
0!
0*
09
0>
0C
#482790000000
1!
1*
b101 6
19
1>
1C
b101 G
#482800000000
0!
0*
09
0>
0C
#482810000000
1!
1*
b110 6
19
1>
1C
b110 G
#482820000000
0!
0*
09
0>
0C
#482830000000
1!
1*
b111 6
19
1>
1C
b111 G
#482840000000
0!
1"
0*
1+
09
1:
0>
0C
#482850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#482860000000
0!
0*
09
0>
0C
#482870000000
1!
1*
b1 6
19
1>
1C
b1 G
#482880000000
0!
0*
09
0>
0C
#482890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#482900000000
0!
0*
09
0>
0C
#482910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#482920000000
0!
0*
09
0>
0C
#482930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#482940000000
0!
0*
09
0>
0C
#482950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#482960000000
0!
0#
0*
0,
09
0>
0?
0C
#482970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#482980000000
0!
0*
09
0>
0C
#482990000000
1!
1*
19
1>
1C
#483000000000
0!
0*
09
0>
0C
#483010000000
1!
1*
19
1>
1C
#483020000000
0!
0*
09
0>
0C
#483030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#483040000000
0!
0*
09
0>
0C
#483050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#483060000000
0!
0*
09
0>
0C
#483070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#483080000000
0!
0*
09
0>
0C
#483090000000
1!
1*
b10 6
19
1>
1C
b10 G
#483100000000
0!
0*
09
0>
0C
#483110000000
1!
1*
b11 6
19
1>
1C
b11 G
#483120000000
0!
0*
09
0>
0C
#483130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#483140000000
0!
0*
09
0>
0C
#483150000000
1!
1*
b101 6
19
1>
1C
b101 G
#483160000000
0!
0*
09
0>
0C
#483170000000
1!
1*
b110 6
19
1>
1C
b110 G
#483180000000
0!
0*
09
0>
0C
#483190000000
1!
1*
b111 6
19
1>
1C
b111 G
#483200000000
0!
0*
09
0>
0C
#483210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#483220000000
0!
0*
09
0>
0C
#483230000000
1!
1*
b1 6
19
1>
1C
b1 G
#483240000000
0!
0*
09
0>
0C
#483250000000
1!
1*
b10 6
19
1>
1C
b10 G
#483260000000
0!
0*
09
0>
0C
#483270000000
1!
1*
b11 6
19
1>
1C
b11 G
#483280000000
0!
0*
09
0>
0C
#483290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#483300000000
0!
0*
09
0>
0C
#483310000000
1!
1*
b101 6
19
1>
1C
b101 G
#483320000000
0!
0*
09
0>
0C
#483330000000
1!
1*
b110 6
19
1>
1C
b110 G
#483340000000
0!
0*
09
0>
0C
#483350000000
1!
1*
b111 6
19
1>
1C
b111 G
#483360000000
0!
0*
09
0>
0C
#483370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#483380000000
0!
0*
09
0>
0C
#483390000000
1!
1*
b1 6
19
1>
1C
b1 G
#483400000000
0!
0*
09
0>
0C
#483410000000
1!
1*
b10 6
19
1>
1C
b10 G
#483420000000
0!
0*
09
0>
0C
#483430000000
1!
1*
b11 6
19
1>
1C
b11 G
#483440000000
0!
0*
09
0>
0C
#483450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#483460000000
0!
0*
09
0>
0C
#483470000000
1!
1*
b101 6
19
1>
1C
b101 G
#483480000000
0!
0*
09
0>
0C
#483490000000
1!
1*
b110 6
19
1>
1C
b110 G
#483500000000
0!
0*
09
0>
0C
#483510000000
1!
1*
b111 6
19
1>
1C
b111 G
#483520000000
0!
1"
0*
1+
09
1:
0>
0C
#483530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#483540000000
0!
0*
09
0>
0C
#483550000000
1!
1*
b1 6
19
1>
1C
b1 G
#483560000000
0!
0*
09
0>
0C
#483570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#483580000000
0!
0*
09
0>
0C
#483590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#483600000000
0!
0*
09
0>
0C
#483610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#483620000000
0!
0*
09
0>
0C
#483630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#483640000000
0!
0#
0*
0,
09
0>
0?
0C
#483650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#483660000000
0!
0*
09
0>
0C
#483670000000
1!
1*
19
1>
1C
#483680000000
0!
0*
09
0>
0C
#483690000000
1!
1*
19
1>
1C
#483700000000
0!
0*
09
0>
0C
#483710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#483720000000
0!
0*
09
0>
0C
#483730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#483740000000
0!
0*
09
0>
0C
#483750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#483760000000
0!
0*
09
0>
0C
#483770000000
1!
1*
b10 6
19
1>
1C
b10 G
#483780000000
0!
0*
09
0>
0C
#483790000000
1!
1*
b11 6
19
1>
1C
b11 G
#483800000000
0!
0*
09
0>
0C
#483810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#483820000000
0!
0*
09
0>
0C
#483830000000
1!
1*
b101 6
19
1>
1C
b101 G
#483840000000
0!
0*
09
0>
0C
#483850000000
1!
1*
b110 6
19
1>
1C
b110 G
#483860000000
0!
0*
09
0>
0C
#483870000000
1!
1*
b111 6
19
1>
1C
b111 G
#483880000000
0!
0*
09
0>
0C
#483890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#483900000000
0!
0*
09
0>
0C
#483910000000
1!
1*
b1 6
19
1>
1C
b1 G
#483920000000
0!
0*
09
0>
0C
#483930000000
1!
1*
b10 6
19
1>
1C
b10 G
#483940000000
0!
0*
09
0>
0C
#483950000000
1!
1*
b11 6
19
1>
1C
b11 G
#483960000000
0!
0*
09
0>
0C
#483970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#483980000000
0!
0*
09
0>
0C
#483990000000
1!
1*
b101 6
19
1>
1C
b101 G
#484000000000
0!
0*
09
0>
0C
#484010000000
1!
1*
b110 6
19
1>
1C
b110 G
#484020000000
0!
0*
09
0>
0C
#484030000000
1!
1*
b111 6
19
1>
1C
b111 G
#484040000000
0!
0*
09
0>
0C
#484050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#484060000000
0!
0*
09
0>
0C
#484070000000
1!
1*
b1 6
19
1>
1C
b1 G
#484080000000
0!
0*
09
0>
0C
#484090000000
1!
1*
b10 6
19
1>
1C
b10 G
#484100000000
0!
0*
09
0>
0C
#484110000000
1!
1*
b11 6
19
1>
1C
b11 G
#484120000000
0!
0*
09
0>
0C
#484130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#484140000000
0!
0*
09
0>
0C
#484150000000
1!
1*
b101 6
19
1>
1C
b101 G
#484160000000
0!
0*
09
0>
0C
#484170000000
1!
1*
b110 6
19
1>
1C
b110 G
#484180000000
0!
0*
09
0>
0C
#484190000000
1!
1*
b111 6
19
1>
1C
b111 G
#484200000000
0!
1"
0*
1+
09
1:
0>
0C
#484210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#484220000000
0!
0*
09
0>
0C
#484230000000
1!
1*
b1 6
19
1>
1C
b1 G
#484240000000
0!
0*
09
0>
0C
#484250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#484260000000
0!
0*
09
0>
0C
#484270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#484280000000
0!
0*
09
0>
0C
#484290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#484300000000
0!
0*
09
0>
0C
#484310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#484320000000
0!
0#
0*
0,
09
0>
0?
0C
#484330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#484340000000
0!
0*
09
0>
0C
#484350000000
1!
1*
19
1>
1C
#484360000000
0!
0*
09
0>
0C
#484370000000
1!
1*
19
1>
1C
#484380000000
0!
0*
09
0>
0C
#484390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#484400000000
0!
0*
09
0>
0C
#484410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#484420000000
0!
0*
09
0>
0C
#484430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#484440000000
0!
0*
09
0>
0C
#484450000000
1!
1*
b10 6
19
1>
1C
b10 G
#484460000000
0!
0*
09
0>
0C
#484470000000
1!
1*
b11 6
19
1>
1C
b11 G
#484480000000
0!
0*
09
0>
0C
#484490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#484500000000
0!
0*
09
0>
0C
#484510000000
1!
1*
b101 6
19
1>
1C
b101 G
#484520000000
0!
0*
09
0>
0C
#484530000000
1!
1*
b110 6
19
1>
1C
b110 G
#484540000000
0!
0*
09
0>
0C
#484550000000
1!
1*
b111 6
19
1>
1C
b111 G
#484560000000
0!
0*
09
0>
0C
#484570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#484580000000
0!
0*
09
0>
0C
#484590000000
1!
1*
b1 6
19
1>
1C
b1 G
#484600000000
0!
0*
09
0>
0C
#484610000000
1!
1*
b10 6
19
1>
1C
b10 G
#484620000000
0!
0*
09
0>
0C
#484630000000
1!
1*
b11 6
19
1>
1C
b11 G
#484640000000
0!
0*
09
0>
0C
#484650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#484660000000
0!
0*
09
0>
0C
#484670000000
1!
1*
b101 6
19
1>
1C
b101 G
#484680000000
0!
0*
09
0>
0C
#484690000000
1!
1*
b110 6
19
1>
1C
b110 G
#484700000000
0!
0*
09
0>
0C
#484710000000
1!
1*
b111 6
19
1>
1C
b111 G
#484720000000
0!
0*
09
0>
0C
#484730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#484740000000
0!
0*
09
0>
0C
#484750000000
1!
1*
b1 6
19
1>
1C
b1 G
#484760000000
0!
0*
09
0>
0C
#484770000000
1!
1*
b10 6
19
1>
1C
b10 G
#484780000000
0!
0*
09
0>
0C
#484790000000
1!
1*
b11 6
19
1>
1C
b11 G
#484800000000
0!
0*
09
0>
0C
#484810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#484820000000
0!
0*
09
0>
0C
#484830000000
1!
1*
b101 6
19
1>
1C
b101 G
#484840000000
0!
0*
09
0>
0C
#484850000000
1!
1*
b110 6
19
1>
1C
b110 G
#484860000000
0!
0*
09
0>
0C
#484870000000
1!
1*
b111 6
19
1>
1C
b111 G
#484880000000
0!
1"
0*
1+
09
1:
0>
0C
#484890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#484900000000
0!
0*
09
0>
0C
#484910000000
1!
1*
b1 6
19
1>
1C
b1 G
#484920000000
0!
0*
09
0>
0C
#484930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#484940000000
0!
0*
09
0>
0C
#484950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#484960000000
0!
0*
09
0>
0C
#484970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#484980000000
0!
0*
09
0>
0C
#484990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#485000000000
0!
0#
0*
0,
09
0>
0?
0C
#485010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#485020000000
0!
0*
09
0>
0C
#485030000000
1!
1*
19
1>
1C
#485040000000
0!
0*
09
0>
0C
#485050000000
1!
1*
19
1>
1C
#485060000000
0!
0*
09
0>
0C
#485070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#485080000000
0!
0*
09
0>
0C
#485090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#485100000000
0!
0*
09
0>
0C
#485110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#485120000000
0!
0*
09
0>
0C
#485130000000
1!
1*
b10 6
19
1>
1C
b10 G
#485140000000
0!
0*
09
0>
0C
#485150000000
1!
1*
b11 6
19
1>
1C
b11 G
#485160000000
0!
0*
09
0>
0C
#485170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#485180000000
0!
0*
09
0>
0C
#485190000000
1!
1*
b101 6
19
1>
1C
b101 G
#485200000000
0!
0*
09
0>
0C
#485210000000
1!
1*
b110 6
19
1>
1C
b110 G
#485220000000
0!
0*
09
0>
0C
#485230000000
1!
1*
b111 6
19
1>
1C
b111 G
#485240000000
0!
0*
09
0>
0C
#485250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#485260000000
0!
0*
09
0>
0C
#485270000000
1!
1*
b1 6
19
1>
1C
b1 G
#485280000000
0!
0*
09
0>
0C
#485290000000
1!
1*
b10 6
19
1>
1C
b10 G
#485300000000
0!
0*
09
0>
0C
#485310000000
1!
1*
b11 6
19
1>
1C
b11 G
#485320000000
0!
0*
09
0>
0C
#485330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#485340000000
0!
0*
09
0>
0C
#485350000000
1!
1*
b101 6
19
1>
1C
b101 G
#485360000000
0!
0*
09
0>
0C
#485370000000
1!
1*
b110 6
19
1>
1C
b110 G
#485380000000
0!
0*
09
0>
0C
#485390000000
1!
1*
b111 6
19
1>
1C
b111 G
#485400000000
0!
0*
09
0>
0C
#485410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#485420000000
0!
0*
09
0>
0C
#485430000000
1!
1*
b1 6
19
1>
1C
b1 G
#485440000000
0!
0*
09
0>
0C
#485450000000
1!
1*
b10 6
19
1>
1C
b10 G
#485460000000
0!
0*
09
0>
0C
#485470000000
1!
1*
b11 6
19
1>
1C
b11 G
#485480000000
0!
0*
09
0>
0C
#485490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#485500000000
0!
0*
09
0>
0C
#485510000000
1!
1*
b101 6
19
1>
1C
b101 G
#485520000000
0!
0*
09
0>
0C
#485530000000
1!
1*
b110 6
19
1>
1C
b110 G
#485540000000
0!
0*
09
0>
0C
#485550000000
1!
1*
b111 6
19
1>
1C
b111 G
#485560000000
0!
1"
0*
1+
09
1:
0>
0C
#485570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#485580000000
0!
0*
09
0>
0C
#485590000000
1!
1*
b1 6
19
1>
1C
b1 G
#485600000000
0!
0*
09
0>
0C
#485610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#485620000000
0!
0*
09
0>
0C
#485630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#485640000000
0!
0*
09
0>
0C
#485650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#485660000000
0!
0*
09
0>
0C
#485670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#485680000000
0!
0#
0*
0,
09
0>
0?
0C
#485690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#485700000000
0!
0*
09
0>
0C
#485710000000
1!
1*
19
1>
1C
#485720000000
0!
0*
09
0>
0C
#485730000000
1!
1*
19
1>
1C
#485740000000
0!
0*
09
0>
0C
#485750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#485760000000
0!
0*
09
0>
0C
#485770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#485780000000
0!
0*
09
0>
0C
#485790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#485800000000
0!
0*
09
0>
0C
#485810000000
1!
1*
b10 6
19
1>
1C
b10 G
#485820000000
0!
0*
09
0>
0C
#485830000000
1!
1*
b11 6
19
1>
1C
b11 G
#485840000000
0!
0*
09
0>
0C
#485850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#485860000000
0!
0*
09
0>
0C
#485870000000
1!
1*
b101 6
19
1>
1C
b101 G
#485880000000
0!
0*
09
0>
0C
#485890000000
1!
1*
b110 6
19
1>
1C
b110 G
#485900000000
0!
0*
09
0>
0C
#485910000000
1!
1*
b111 6
19
1>
1C
b111 G
#485920000000
0!
0*
09
0>
0C
#485930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#485940000000
0!
0*
09
0>
0C
#485950000000
1!
1*
b1 6
19
1>
1C
b1 G
#485960000000
0!
0*
09
0>
0C
#485970000000
1!
1*
b10 6
19
1>
1C
b10 G
#485980000000
0!
0*
09
0>
0C
#485990000000
1!
1*
b11 6
19
1>
1C
b11 G
#486000000000
0!
0*
09
0>
0C
#486010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#486020000000
0!
0*
09
0>
0C
#486030000000
1!
1*
b101 6
19
1>
1C
b101 G
#486040000000
0!
0*
09
0>
0C
#486050000000
1!
1*
b110 6
19
1>
1C
b110 G
#486060000000
0!
0*
09
0>
0C
#486070000000
1!
1*
b111 6
19
1>
1C
b111 G
#486080000000
0!
0*
09
0>
0C
#486090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#486100000000
0!
0*
09
0>
0C
#486110000000
1!
1*
b1 6
19
1>
1C
b1 G
#486120000000
0!
0*
09
0>
0C
#486130000000
1!
1*
b10 6
19
1>
1C
b10 G
#486140000000
0!
0*
09
0>
0C
#486150000000
1!
1*
b11 6
19
1>
1C
b11 G
#486160000000
0!
0*
09
0>
0C
#486170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#486180000000
0!
0*
09
0>
0C
#486190000000
1!
1*
b101 6
19
1>
1C
b101 G
#486200000000
0!
0*
09
0>
0C
#486210000000
1!
1*
b110 6
19
1>
1C
b110 G
#486220000000
0!
0*
09
0>
0C
#486230000000
1!
1*
b111 6
19
1>
1C
b111 G
#486240000000
0!
1"
0*
1+
09
1:
0>
0C
#486250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#486260000000
0!
0*
09
0>
0C
#486270000000
1!
1*
b1 6
19
1>
1C
b1 G
#486280000000
0!
0*
09
0>
0C
#486290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#486300000000
0!
0*
09
0>
0C
#486310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#486320000000
0!
0*
09
0>
0C
#486330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#486340000000
0!
0*
09
0>
0C
#486350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#486360000000
0!
0#
0*
0,
09
0>
0?
0C
#486370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#486380000000
0!
0*
09
0>
0C
#486390000000
1!
1*
19
1>
1C
#486400000000
0!
0*
09
0>
0C
#486410000000
1!
1*
19
1>
1C
#486420000000
0!
0*
09
0>
0C
#486430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#486440000000
0!
0*
09
0>
0C
#486450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#486460000000
0!
0*
09
0>
0C
#486470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#486480000000
0!
0*
09
0>
0C
#486490000000
1!
1*
b10 6
19
1>
1C
b10 G
#486500000000
0!
0*
09
0>
0C
#486510000000
1!
1*
b11 6
19
1>
1C
b11 G
#486520000000
0!
0*
09
0>
0C
#486530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#486540000000
0!
0*
09
0>
0C
#486550000000
1!
1*
b101 6
19
1>
1C
b101 G
#486560000000
0!
0*
09
0>
0C
#486570000000
1!
1*
b110 6
19
1>
1C
b110 G
#486580000000
0!
0*
09
0>
0C
#486590000000
1!
1*
b111 6
19
1>
1C
b111 G
#486600000000
0!
0*
09
0>
0C
#486610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#486620000000
0!
0*
09
0>
0C
#486630000000
1!
1*
b1 6
19
1>
1C
b1 G
#486640000000
0!
0*
09
0>
0C
#486650000000
1!
1*
b10 6
19
1>
1C
b10 G
#486660000000
0!
0*
09
0>
0C
#486670000000
1!
1*
b11 6
19
1>
1C
b11 G
#486680000000
0!
0*
09
0>
0C
#486690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#486700000000
0!
0*
09
0>
0C
#486710000000
1!
1*
b101 6
19
1>
1C
b101 G
#486720000000
0!
0*
09
0>
0C
#486730000000
1!
1*
b110 6
19
1>
1C
b110 G
#486740000000
0!
0*
09
0>
0C
#486750000000
1!
1*
b111 6
19
1>
1C
b111 G
#486760000000
0!
0*
09
0>
0C
#486770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#486780000000
0!
0*
09
0>
0C
#486790000000
1!
1*
b1 6
19
1>
1C
b1 G
#486800000000
0!
0*
09
0>
0C
#486810000000
1!
1*
b10 6
19
1>
1C
b10 G
#486820000000
0!
0*
09
0>
0C
#486830000000
1!
1*
b11 6
19
1>
1C
b11 G
#486840000000
0!
0*
09
0>
0C
#486850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#486860000000
0!
0*
09
0>
0C
#486870000000
1!
1*
b101 6
19
1>
1C
b101 G
#486880000000
0!
0*
09
0>
0C
#486890000000
1!
1*
b110 6
19
1>
1C
b110 G
#486900000000
0!
0*
09
0>
0C
#486910000000
1!
1*
b111 6
19
1>
1C
b111 G
#486920000000
0!
1"
0*
1+
09
1:
0>
0C
#486930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#486940000000
0!
0*
09
0>
0C
#486950000000
1!
1*
b1 6
19
1>
1C
b1 G
#486960000000
0!
0*
09
0>
0C
#486970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#486980000000
0!
0*
09
0>
0C
#486990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#487000000000
0!
0*
09
0>
0C
#487010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#487020000000
0!
0*
09
0>
0C
#487030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#487040000000
0!
0#
0*
0,
09
0>
0?
0C
#487050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#487060000000
0!
0*
09
0>
0C
#487070000000
1!
1*
19
1>
1C
#487080000000
0!
0*
09
0>
0C
#487090000000
1!
1*
19
1>
1C
#487100000000
0!
0*
09
0>
0C
#487110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#487120000000
0!
0*
09
0>
0C
#487130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#487140000000
0!
0*
09
0>
0C
#487150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#487160000000
0!
0*
09
0>
0C
#487170000000
1!
1*
b10 6
19
1>
1C
b10 G
#487180000000
0!
0*
09
0>
0C
#487190000000
1!
1*
b11 6
19
1>
1C
b11 G
#487200000000
0!
0*
09
0>
0C
#487210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#487220000000
0!
0*
09
0>
0C
#487230000000
1!
1*
b101 6
19
1>
1C
b101 G
#487240000000
0!
0*
09
0>
0C
#487250000000
1!
1*
b110 6
19
1>
1C
b110 G
#487260000000
0!
0*
09
0>
0C
#487270000000
1!
1*
b111 6
19
1>
1C
b111 G
#487280000000
0!
0*
09
0>
0C
#487290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#487300000000
0!
0*
09
0>
0C
#487310000000
1!
1*
b1 6
19
1>
1C
b1 G
#487320000000
0!
0*
09
0>
0C
#487330000000
1!
1*
b10 6
19
1>
1C
b10 G
#487340000000
0!
0*
09
0>
0C
#487350000000
1!
1*
b11 6
19
1>
1C
b11 G
#487360000000
0!
0*
09
0>
0C
#487370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#487380000000
0!
0*
09
0>
0C
#487390000000
1!
1*
b101 6
19
1>
1C
b101 G
#487400000000
0!
0*
09
0>
0C
#487410000000
1!
1*
b110 6
19
1>
1C
b110 G
#487420000000
0!
0*
09
0>
0C
#487430000000
1!
1*
b111 6
19
1>
1C
b111 G
#487440000000
0!
0*
09
0>
0C
#487450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#487460000000
0!
0*
09
0>
0C
#487470000000
1!
1*
b1 6
19
1>
1C
b1 G
#487480000000
0!
0*
09
0>
0C
#487490000000
1!
1*
b10 6
19
1>
1C
b10 G
#487500000000
0!
0*
09
0>
0C
#487510000000
1!
1*
b11 6
19
1>
1C
b11 G
#487520000000
0!
0*
09
0>
0C
#487530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#487540000000
0!
0*
09
0>
0C
#487550000000
1!
1*
b101 6
19
1>
1C
b101 G
#487560000000
0!
0*
09
0>
0C
#487570000000
1!
1*
b110 6
19
1>
1C
b110 G
#487580000000
0!
0*
09
0>
0C
#487590000000
1!
1*
b111 6
19
1>
1C
b111 G
#487600000000
0!
1"
0*
1+
09
1:
0>
0C
#487610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#487620000000
0!
0*
09
0>
0C
#487630000000
1!
1*
b1 6
19
1>
1C
b1 G
#487640000000
0!
0*
09
0>
0C
#487650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#487660000000
0!
0*
09
0>
0C
#487670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#487680000000
0!
0*
09
0>
0C
#487690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#487700000000
0!
0*
09
0>
0C
#487710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#487720000000
0!
0#
0*
0,
09
0>
0?
0C
#487730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#487740000000
0!
0*
09
0>
0C
#487750000000
1!
1*
19
1>
1C
#487760000000
0!
0*
09
0>
0C
#487770000000
1!
1*
19
1>
1C
#487780000000
0!
0*
09
0>
0C
#487790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#487800000000
0!
0*
09
0>
0C
#487810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#487820000000
0!
0*
09
0>
0C
#487830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#487840000000
0!
0*
09
0>
0C
#487850000000
1!
1*
b10 6
19
1>
1C
b10 G
#487860000000
0!
0*
09
0>
0C
#487870000000
1!
1*
b11 6
19
1>
1C
b11 G
#487880000000
0!
0*
09
0>
0C
#487890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#487900000000
0!
0*
09
0>
0C
#487910000000
1!
1*
b101 6
19
1>
1C
b101 G
#487920000000
0!
0*
09
0>
0C
#487930000000
1!
1*
b110 6
19
1>
1C
b110 G
#487940000000
0!
0*
09
0>
0C
#487950000000
1!
1*
b111 6
19
1>
1C
b111 G
#487960000000
0!
0*
09
0>
0C
#487970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#487980000000
0!
0*
09
0>
0C
#487990000000
1!
1*
b1 6
19
1>
1C
b1 G
#488000000000
0!
0*
09
0>
0C
#488010000000
1!
1*
b10 6
19
1>
1C
b10 G
#488020000000
0!
0*
09
0>
0C
#488030000000
1!
1*
b11 6
19
1>
1C
b11 G
#488040000000
0!
0*
09
0>
0C
#488050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#488060000000
0!
0*
09
0>
0C
#488070000000
1!
1*
b101 6
19
1>
1C
b101 G
#488080000000
0!
0*
09
0>
0C
#488090000000
1!
1*
b110 6
19
1>
1C
b110 G
#488100000000
0!
0*
09
0>
0C
#488110000000
1!
1*
b111 6
19
1>
1C
b111 G
#488120000000
0!
0*
09
0>
0C
#488130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#488140000000
0!
0*
09
0>
0C
#488150000000
1!
1*
b1 6
19
1>
1C
b1 G
#488160000000
0!
0*
09
0>
0C
#488170000000
1!
1*
b10 6
19
1>
1C
b10 G
#488180000000
0!
0*
09
0>
0C
#488190000000
1!
1*
b11 6
19
1>
1C
b11 G
#488200000000
0!
0*
09
0>
0C
#488210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#488220000000
0!
0*
09
0>
0C
#488230000000
1!
1*
b101 6
19
1>
1C
b101 G
#488240000000
0!
0*
09
0>
0C
#488250000000
1!
1*
b110 6
19
1>
1C
b110 G
#488260000000
0!
0*
09
0>
0C
#488270000000
1!
1*
b111 6
19
1>
1C
b111 G
#488280000000
0!
1"
0*
1+
09
1:
0>
0C
#488290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#488300000000
0!
0*
09
0>
0C
#488310000000
1!
1*
b1 6
19
1>
1C
b1 G
#488320000000
0!
0*
09
0>
0C
#488330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#488340000000
0!
0*
09
0>
0C
#488350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#488360000000
0!
0*
09
0>
0C
#488370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#488380000000
0!
0*
09
0>
0C
#488390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#488400000000
0!
0#
0*
0,
09
0>
0?
0C
#488410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#488420000000
0!
0*
09
0>
0C
#488430000000
1!
1*
19
1>
1C
#488440000000
0!
0*
09
0>
0C
#488450000000
1!
1*
19
1>
1C
#488460000000
0!
0*
09
0>
0C
#488470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#488480000000
0!
0*
09
0>
0C
#488490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#488500000000
0!
0*
09
0>
0C
#488510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#488520000000
0!
0*
09
0>
0C
#488530000000
1!
1*
b10 6
19
1>
1C
b10 G
#488540000000
0!
0*
09
0>
0C
#488550000000
1!
1*
b11 6
19
1>
1C
b11 G
#488560000000
0!
0*
09
0>
0C
#488570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#488580000000
0!
0*
09
0>
0C
#488590000000
1!
1*
b101 6
19
1>
1C
b101 G
#488600000000
0!
0*
09
0>
0C
#488610000000
1!
1*
b110 6
19
1>
1C
b110 G
#488620000000
0!
0*
09
0>
0C
#488630000000
1!
1*
b111 6
19
1>
1C
b111 G
#488640000000
0!
0*
09
0>
0C
#488650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#488660000000
0!
0*
09
0>
0C
#488670000000
1!
1*
b1 6
19
1>
1C
b1 G
#488680000000
0!
0*
09
0>
0C
#488690000000
1!
1*
b10 6
19
1>
1C
b10 G
#488700000000
0!
0*
09
0>
0C
#488710000000
1!
1*
b11 6
19
1>
1C
b11 G
#488720000000
0!
0*
09
0>
0C
#488730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#488740000000
0!
0*
09
0>
0C
#488750000000
1!
1*
b101 6
19
1>
1C
b101 G
#488760000000
0!
0*
09
0>
0C
#488770000000
1!
1*
b110 6
19
1>
1C
b110 G
#488780000000
0!
0*
09
0>
0C
#488790000000
1!
1*
b111 6
19
1>
1C
b111 G
#488800000000
0!
0*
09
0>
0C
#488810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#488820000000
0!
0*
09
0>
0C
#488830000000
1!
1*
b1 6
19
1>
1C
b1 G
#488840000000
0!
0*
09
0>
0C
#488850000000
1!
1*
b10 6
19
1>
1C
b10 G
#488860000000
0!
0*
09
0>
0C
#488870000000
1!
1*
b11 6
19
1>
1C
b11 G
#488880000000
0!
0*
09
0>
0C
#488890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#488900000000
0!
0*
09
0>
0C
#488910000000
1!
1*
b101 6
19
1>
1C
b101 G
#488920000000
0!
0*
09
0>
0C
#488930000000
1!
1*
b110 6
19
1>
1C
b110 G
#488940000000
0!
0*
09
0>
0C
#488950000000
1!
1*
b111 6
19
1>
1C
b111 G
#488960000000
0!
1"
0*
1+
09
1:
0>
0C
#488970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#488980000000
0!
0*
09
0>
0C
#488990000000
1!
1*
b1 6
19
1>
1C
b1 G
#489000000000
0!
0*
09
0>
0C
#489010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#489020000000
0!
0*
09
0>
0C
#489030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#489040000000
0!
0*
09
0>
0C
#489050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#489060000000
0!
0*
09
0>
0C
#489070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#489080000000
0!
0#
0*
0,
09
0>
0?
0C
#489090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#489100000000
0!
0*
09
0>
0C
#489110000000
1!
1*
19
1>
1C
#489120000000
0!
0*
09
0>
0C
#489130000000
1!
1*
19
1>
1C
#489140000000
0!
0*
09
0>
0C
#489150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#489160000000
0!
0*
09
0>
0C
#489170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#489180000000
0!
0*
09
0>
0C
#489190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#489200000000
0!
0*
09
0>
0C
#489210000000
1!
1*
b10 6
19
1>
1C
b10 G
#489220000000
0!
0*
09
0>
0C
#489230000000
1!
1*
b11 6
19
1>
1C
b11 G
#489240000000
0!
0*
09
0>
0C
#489250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#489260000000
0!
0*
09
0>
0C
#489270000000
1!
1*
b101 6
19
1>
1C
b101 G
#489280000000
0!
0*
09
0>
0C
#489290000000
1!
1*
b110 6
19
1>
1C
b110 G
#489300000000
0!
0*
09
0>
0C
#489310000000
1!
1*
b111 6
19
1>
1C
b111 G
#489320000000
0!
0*
09
0>
0C
#489330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#489340000000
0!
0*
09
0>
0C
#489350000000
1!
1*
b1 6
19
1>
1C
b1 G
#489360000000
0!
0*
09
0>
0C
#489370000000
1!
1*
b10 6
19
1>
1C
b10 G
#489380000000
0!
0*
09
0>
0C
#489390000000
1!
1*
b11 6
19
1>
1C
b11 G
#489400000000
0!
0*
09
0>
0C
#489410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#489420000000
0!
0*
09
0>
0C
#489430000000
1!
1*
b101 6
19
1>
1C
b101 G
#489440000000
0!
0*
09
0>
0C
#489450000000
1!
1*
b110 6
19
1>
1C
b110 G
#489460000000
0!
0*
09
0>
0C
#489470000000
1!
1*
b111 6
19
1>
1C
b111 G
#489480000000
0!
0*
09
0>
0C
#489490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#489500000000
0!
0*
09
0>
0C
#489510000000
1!
1*
b1 6
19
1>
1C
b1 G
#489520000000
0!
0*
09
0>
0C
#489530000000
1!
1*
b10 6
19
1>
1C
b10 G
#489540000000
0!
0*
09
0>
0C
#489550000000
1!
1*
b11 6
19
1>
1C
b11 G
#489560000000
0!
0*
09
0>
0C
#489570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#489580000000
0!
0*
09
0>
0C
#489590000000
1!
1*
b101 6
19
1>
1C
b101 G
#489600000000
0!
0*
09
0>
0C
#489610000000
1!
1*
b110 6
19
1>
1C
b110 G
#489620000000
0!
0*
09
0>
0C
#489630000000
1!
1*
b111 6
19
1>
1C
b111 G
#489640000000
0!
1"
0*
1+
09
1:
0>
0C
#489650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#489660000000
0!
0*
09
0>
0C
#489670000000
1!
1*
b1 6
19
1>
1C
b1 G
#489680000000
0!
0*
09
0>
0C
#489690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#489700000000
0!
0*
09
0>
0C
#489710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#489720000000
0!
0*
09
0>
0C
#489730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#489740000000
0!
0*
09
0>
0C
#489750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#489760000000
0!
0#
0*
0,
09
0>
0?
0C
#489770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#489780000000
0!
0*
09
0>
0C
#489790000000
1!
1*
19
1>
1C
#489800000000
0!
0*
09
0>
0C
#489810000000
1!
1*
19
1>
1C
#489820000000
0!
0*
09
0>
0C
#489830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#489840000000
0!
0*
09
0>
0C
#489850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#489860000000
0!
0*
09
0>
0C
#489870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#489880000000
0!
0*
09
0>
0C
#489890000000
1!
1*
b10 6
19
1>
1C
b10 G
#489900000000
0!
0*
09
0>
0C
#489910000000
1!
1*
b11 6
19
1>
1C
b11 G
#489920000000
0!
0*
09
0>
0C
#489930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#489940000000
0!
0*
09
0>
0C
#489950000000
1!
1*
b101 6
19
1>
1C
b101 G
#489960000000
0!
0*
09
0>
0C
#489970000000
1!
1*
b110 6
19
1>
1C
b110 G
#489980000000
0!
0*
09
0>
0C
#489990000000
1!
1*
b111 6
19
1>
1C
b111 G
#490000000000
0!
0*
09
0>
0C
#490010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#490020000000
0!
0*
09
0>
0C
#490030000000
1!
1*
b1 6
19
1>
1C
b1 G
#490040000000
0!
0*
09
0>
0C
#490050000000
1!
1*
b10 6
19
1>
1C
b10 G
#490060000000
0!
0*
09
0>
0C
#490070000000
1!
1*
b11 6
19
1>
1C
b11 G
#490080000000
0!
0*
09
0>
0C
#490090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#490100000000
0!
0*
09
0>
0C
#490110000000
1!
1*
b101 6
19
1>
1C
b101 G
#490120000000
0!
0*
09
0>
0C
#490130000000
1!
1*
b110 6
19
1>
1C
b110 G
#490140000000
0!
0*
09
0>
0C
#490150000000
1!
1*
b111 6
19
1>
1C
b111 G
#490160000000
0!
0*
09
0>
0C
#490170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#490180000000
0!
0*
09
0>
0C
#490190000000
1!
1*
b1 6
19
1>
1C
b1 G
#490200000000
0!
0*
09
0>
0C
#490210000000
1!
1*
b10 6
19
1>
1C
b10 G
#490220000000
0!
0*
09
0>
0C
#490230000000
1!
1*
b11 6
19
1>
1C
b11 G
#490240000000
0!
0*
09
0>
0C
#490250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#490260000000
0!
0*
09
0>
0C
#490270000000
1!
1*
b101 6
19
1>
1C
b101 G
#490280000000
0!
0*
09
0>
0C
#490290000000
1!
1*
b110 6
19
1>
1C
b110 G
#490300000000
0!
0*
09
0>
0C
#490310000000
1!
1*
b111 6
19
1>
1C
b111 G
#490320000000
0!
1"
0*
1+
09
1:
0>
0C
#490330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#490340000000
0!
0*
09
0>
0C
#490350000000
1!
1*
b1 6
19
1>
1C
b1 G
#490360000000
0!
0*
09
0>
0C
#490370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#490380000000
0!
0*
09
0>
0C
#490390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#490400000000
0!
0*
09
0>
0C
#490410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#490420000000
0!
0*
09
0>
0C
#490430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#490440000000
0!
0#
0*
0,
09
0>
0?
0C
#490450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#490460000000
0!
0*
09
0>
0C
#490470000000
1!
1*
19
1>
1C
#490480000000
0!
0*
09
0>
0C
#490490000000
1!
1*
19
1>
1C
#490500000000
0!
0*
09
0>
0C
#490510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#490520000000
0!
0*
09
0>
0C
#490530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#490540000000
0!
0*
09
0>
0C
#490550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#490560000000
0!
0*
09
0>
0C
#490570000000
1!
1*
b10 6
19
1>
1C
b10 G
#490580000000
0!
0*
09
0>
0C
#490590000000
1!
1*
b11 6
19
1>
1C
b11 G
#490600000000
0!
0*
09
0>
0C
#490610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#490620000000
0!
0*
09
0>
0C
#490630000000
1!
1*
b101 6
19
1>
1C
b101 G
#490640000000
0!
0*
09
0>
0C
#490650000000
1!
1*
b110 6
19
1>
1C
b110 G
#490660000000
0!
0*
09
0>
0C
#490670000000
1!
1*
b111 6
19
1>
1C
b111 G
#490680000000
0!
0*
09
0>
0C
#490690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#490700000000
0!
0*
09
0>
0C
#490710000000
1!
1*
b1 6
19
1>
1C
b1 G
#490720000000
0!
0*
09
0>
0C
#490730000000
1!
1*
b10 6
19
1>
1C
b10 G
#490740000000
0!
0*
09
0>
0C
#490750000000
1!
1*
b11 6
19
1>
1C
b11 G
#490760000000
0!
0*
09
0>
0C
#490770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#490780000000
0!
0*
09
0>
0C
#490790000000
1!
1*
b101 6
19
1>
1C
b101 G
#490800000000
0!
0*
09
0>
0C
#490810000000
1!
1*
b110 6
19
1>
1C
b110 G
#490820000000
0!
0*
09
0>
0C
#490830000000
1!
1*
b111 6
19
1>
1C
b111 G
#490840000000
0!
0*
09
0>
0C
#490850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#490860000000
0!
0*
09
0>
0C
#490870000000
1!
1*
b1 6
19
1>
1C
b1 G
#490880000000
0!
0*
09
0>
0C
#490890000000
1!
1*
b10 6
19
1>
1C
b10 G
#490900000000
0!
0*
09
0>
0C
#490910000000
1!
1*
b11 6
19
1>
1C
b11 G
#490920000000
0!
0*
09
0>
0C
#490930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#490940000000
0!
0*
09
0>
0C
#490950000000
1!
1*
b101 6
19
1>
1C
b101 G
#490960000000
0!
0*
09
0>
0C
#490970000000
1!
1*
b110 6
19
1>
1C
b110 G
#490980000000
0!
0*
09
0>
0C
#490990000000
1!
1*
b111 6
19
1>
1C
b111 G
#491000000000
0!
1"
0*
1+
09
1:
0>
0C
#491010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#491020000000
0!
0*
09
0>
0C
#491030000000
1!
1*
b1 6
19
1>
1C
b1 G
#491040000000
0!
0*
09
0>
0C
#491050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#491060000000
0!
0*
09
0>
0C
#491070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#491080000000
0!
0*
09
0>
0C
#491090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#491100000000
0!
0*
09
0>
0C
#491110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#491120000000
0!
0#
0*
0,
09
0>
0?
0C
#491130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#491140000000
0!
0*
09
0>
0C
#491150000000
1!
1*
19
1>
1C
#491160000000
0!
0*
09
0>
0C
#491170000000
1!
1*
19
1>
1C
#491180000000
0!
0*
09
0>
0C
#491190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#491200000000
0!
0*
09
0>
0C
#491210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#491220000000
0!
0*
09
0>
0C
#491230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#491240000000
0!
0*
09
0>
0C
#491250000000
1!
1*
b10 6
19
1>
1C
b10 G
#491260000000
0!
0*
09
0>
0C
#491270000000
1!
1*
b11 6
19
1>
1C
b11 G
#491280000000
0!
0*
09
0>
0C
#491290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#491300000000
0!
0*
09
0>
0C
#491310000000
1!
1*
b101 6
19
1>
1C
b101 G
#491320000000
0!
0*
09
0>
0C
#491330000000
1!
1*
b110 6
19
1>
1C
b110 G
#491340000000
0!
0*
09
0>
0C
#491350000000
1!
1*
b111 6
19
1>
1C
b111 G
#491360000000
0!
0*
09
0>
0C
#491370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#491380000000
0!
0*
09
0>
0C
#491390000000
1!
1*
b1 6
19
1>
1C
b1 G
#491400000000
0!
0*
09
0>
0C
#491410000000
1!
1*
b10 6
19
1>
1C
b10 G
#491420000000
0!
0*
09
0>
0C
#491430000000
1!
1*
b11 6
19
1>
1C
b11 G
#491440000000
0!
0*
09
0>
0C
#491450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#491460000000
0!
0*
09
0>
0C
#491470000000
1!
1*
b101 6
19
1>
1C
b101 G
#491480000000
0!
0*
09
0>
0C
#491490000000
1!
1*
b110 6
19
1>
1C
b110 G
#491500000000
0!
0*
09
0>
0C
#491510000000
1!
1*
b111 6
19
1>
1C
b111 G
#491520000000
0!
0*
09
0>
0C
#491530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#491540000000
0!
0*
09
0>
0C
#491550000000
1!
1*
b1 6
19
1>
1C
b1 G
#491560000000
0!
0*
09
0>
0C
#491570000000
1!
1*
b10 6
19
1>
1C
b10 G
#491580000000
0!
0*
09
0>
0C
#491590000000
1!
1*
b11 6
19
1>
1C
b11 G
#491600000000
0!
0*
09
0>
0C
#491610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#491620000000
0!
0*
09
0>
0C
#491630000000
1!
1*
b101 6
19
1>
1C
b101 G
#491640000000
0!
0*
09
0>
0C
#491650000000
1!
1*
b110 6
19
1>
1C
b110 G
#491660000000
0!
0*
09
0>
0C
#491670000000
1!
1*
b111 6
19
1>
1C
b111 G
#491680000000
0!
1"
0*
1+
09
1:
0>
0C
#491690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#491700000000
0!
0*
09
0>
0C
#491710000000
1!
1*
b1 6
19
1>
1C
b1 G
#491720000000
0!
0*
09
0>
0C
#491730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#491740000000
0!
0*
09
0>
0C
#491750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#491760000000
0!
0*
09
0>
0C
#491770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#491780000000
0!
0*
09
0>
0C
#491790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#491800000000
0!
0#
0*
0,
09
0>
0?
0C
#491810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#491820000000
0!
0*
09
0>
0C
#491830000000
1!
1*
19
1>
1C
#491840000000
0!
0*
09
0>
0C
#491850000000
1!
1*
19
1>
1C
#491860000000
0!
0*
09
0>
0C
#491870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#491880000000
0!
0*
09
0>
0C
#491890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#491900000000
0!
0*
09
0>
0C
#491910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#491920000000
0!
0*
09
0>
0C
#491930000000
1!
1*
b10 6
19
1>
1C
b10 G
#491940000000
0!
0*
09
0>
0C
#491950000000
1!
1*
b11 6
19
1>
1C
b11 G
#491960000000
0!
0*
09
0>
0C
#491970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#491980000000
0!
0*
09
0>
0C
#491990000000
1!
1*
b101 6
19
1>
1C
b101 G
#492000000000
0!
0*
09
0>
0C
#492010000000
1!
1*
b110 6
19
1>
1C
b110 G
#492020000000
0!
0*
09
0>
0C
#492030000000
1!
1*
b111 6
19
1>
1C
b111 G
#492040000000
0!
0*
09
0>
0C
#492050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#492060000000
0!
0*
09
0>
0C
#492070000000
1!
1*
b1 6
19
1>
1C
b1 G
#492080000000
0!
0*
09
0>
0C
#492090000000
1!
1*
b10 6
19
1>
1C
b10 G
#492100000000
0!
0*
09
0>
0C
#492110000000
1!
1*
b11 6
19
1>
1C
b11 G
#492120000000
0!
0*
09
0>
0C
#492130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#492140000000
0!
0*
09
0>
0C
#492150000000
1!
1*
b101 6
19
1>
1C
b101 G
#492160000000
0!
0*
09
0>
0C
#492170000000
1!
1*
b110 6
19
1>
1C
b110 G
#492180000000
0!
0*
09
0>
0C
#492190000000
1!
1*
b111 6
19
1>
1C
b111 G
#492200000000
0!
0*
09
0>
0C
#492210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#492220000000
0!
0*
09
0>
0C
#492230000000
1!
1*
b1 6
19
1>
1C
b1 G
#492240000000
0!
0*
09
0>
0C
#492250000000
1!
1*
b10 6
19
1>
1C
b10 G
#492260000000
0!
0*
09
0>
0C
#492270000000
1!
1*
b11 6
19
1>
1C
b11 G
#492280000000
0!
0*
09
0>
0C
#492290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#492300000000
0!
0*
09
0>
0C
#492310000000
1!
1*
b101 6
19
1>
1C
b101 G
#492320000000
0!
0*
09
0>
0C
#492330000000
1!
1*
b110 6
19
1>
1C
b110 G
#492340000000
0!
0*
09
0>
0C
#492350000000
1!
1*
b111 6
19
1>
1C
b111 G
#492360000000
0!
1"
0*
1+
09
1:
0>
0C
#492370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#492380000000
0!
0*
09
0>
0C
#492390000000
1!
1*
b1 6
19
1>
1C
b1 G
#492400000000
0!
0*
09
0>
0C
#492410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#492420000000
0!
0*
09
0>
0C
#492430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#492440000000
0!
0*
09
0>
0C
#492450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#492460000000
0!
0*
09
0>
0C
#492470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#492480000000
0!
0#
0*
0,
09
0>
0?
0C
#492490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#492500000000
0!
0*
09
0>
0C
#492510000000
1!
1*
19
1>
1C
#492520000000
0!
0*
09
0>
0C
#492530000000
1!
1*
19
1>
1C
#492540000000
0!
0*
09
0>
0C
#492550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#492560000000
0!
0*
09
0>
0C
#492570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#492580000000
0!
0*
09
0>
0C
#492590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#492600000000
0!
0*
09
0>
0C
#492610000000
1!
1*
b10 6
19
1>
1C
b10 G
#492620000000
0!
0*
09
0>
0C
#492630000000
1!
1*
b11 6
19
1>
1C
b11 G
#492640000000
0!
0*
09
0>
0C
#492650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#492660000000
0!
0*
09
0>
0C
#492670000000
1!
1*
b101 6
19
1>
1C
b101 G
#492680000000
0!
0*
09
0>
0C
#492690000000
1!
1*
b110 6
19
1>
1C
b110 G
#492700000000
0!
0*
09
0>
0C
#492710000000
1!
1*
b111 6
19
1>
1C
b111 G
#492720000000
0!
0*
09
0>
0C
#492730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#492740000000
0!
0*
09
0>
0C
#492750000000
1!
1*
b1 6
19
1>
1C
b1 G
#492760000000
0!
0*
09
0>
0C
#492770000000
1!
1*
b10 6
19
1>
1C
b10 G
#492780000000
0!
0*
09
0>
0C
#492790000000
1!
1*
b11 6
19
1>
1C
b11 G
#492800000000
0!
0*
09
0>
0C
#492810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#492820000000
0!
0*
09
0>
0C
#492830000000
1!
1*
b101 6
19
1>
1C
b101 G
#492840000000
0!
0*
09
0>
0C
#492850000000
1!
1*
b110 6
19
1>
1C
b110 G
#492860000000
0!
0*
09
0>
0C
#492870000000
1!
1*
b111 6
19
1>
1C
b111 G
#492880000000
0!
0*
09
0>
0C
#492890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#492900000000
0!
0*
09
0>
0C
#492910000000
1!
1*
b1 6
19
1>
1C
b1 G
#492920000000
0!
0*
09
0>
0C
#492930000000
1!
1*
b10 6
19
1>
1C
b10 G
#492940000000
0!
0*
09
0>
0C
#492950000000
1!
1*
b11 6
19
1>
1C
b11 G
#492960000000
0!
0*
09
0>
0C
#492970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#492980000000
0!
0*
09
0>
0C
#492990000000
1!
1*
b101 6
19
1>
1C
b101 G
#493000000000
0!
0*
09
0>
0C
#493010000000
1!
1*
b110 6
19
1>
1C
b110 G
#493020000000
0!
0*
09
0>
0C
#493030000000
1!
1*
b111 6
19
1>
1C
b111 G
#493040000000
0!
1"
0*
1+
09
1:
0>
0C
#493050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#493060000000
0!
0*
09
0>
0C
#493070000000
1!
1*
b1 6
19
1>
1C
b1 G
#493080000000
0!
0*
09
0>
0C
#493090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#493100000000
0!
0*
09
0>
0C
#493110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#493120000000
0!
0*
09
0>
0C
#493130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#493140000000
0!
0*
09
0>
0C
#493150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#493160000000
0!
0#
0*
0,
09
0>
0?
0C
#493170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#493180000000
0!
0*
09
0>
0C
#493190000000
1!
1*
19
1>
1C
#493200000000
0!
0*
09
0>
0C
#493210000000
1!
1*
19
1>
1C
#493220000000
0!
0*
09
0>
0C
#493230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#493240000000
0!
0*
09
0>
0C
#493250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#493260000000
0!
0*
09
0>
0C
#493270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#493280000000
0!
0*
09
0>
0C
#493290000000
1!
1*
b10 6
19
1>
1C
b10 G
#493300000000
0!
0*
09
0>
0C
#493310000000
1!
1*
b11 6
19
1>
1C
b11 G
#493320000000
0!
0*
09
0>
0C
#493330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#493340000000
0!
0*
09
0>
0C
#493350000000
1!
1*
b101 6
19
1>
1C
b101 G
#493360000000
0!
0*
09
0>
0C
#493370000000
1!
1*
b110 6
19
1>
1C
b110 G
#493380000000
0!
0*
09
0>
0C
#493390000000
1!
1*
b111 6
19
1>
1C
b111 G
#493400000000
0!
0*
09
0>
0C
#493410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#493420000000
0!
0*
09
0>
0C
#493430000000
1!
1*
b1 6
19
1>
1C
b1 G
#493440000000
0!
0*
09
0>
0C
#493450000000
1!
1*
b10 6
19
1>
1C
b10 G
#493460000000
0!
0*
09
0>
0C
#493470000000
1!
1*
b11 6
19
1>
1C
b11 G
#493480000000
0!
0*
09
0>
0C
#493490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#493500000000
0!
0*
09
0>
0C
#493510000000
1!
1*
b101 6
19
1>
1C
b101 G
#493520000000
0!
0*
09
0>
0C
#493530000000
1!
1*
b110 6
19
1>
1C
b110 G
#493540000000
0!
0*
09
0>
0C
#493550000000
1!
1*
b111 6
19
1>
1C
b111 G
#493560000000
0!
0*
09
0>
0C
#493570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#493580000000
0!
0*
09
0>
0C
#493590000000
1!
1*
b1 6
19
1>
1C
b1 G
#493600000000
0!
0*
09
0>
0C
#493610000000
1!
1*
b10 6
19
1>
1C
b10 G
#493620000000
0!
0*
09
0>
0C
#493630000000
1!
1*
b11 6
19
1>
1C
b11 G
#493640000000
0!
0*
09
0>
0C
#493650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#493660000000
0!
0*
09
0>
0C
#493670000000
1!
1*
b101 6
19
1>
1C
b101 G
#493680000000
0!
0*
09
0>
0C
#493690000000
1!
1*
b110 6
19
1>
1C
b110 G
#493700000000
0!
0*
09
0>
0C
#493710000000
1!
1*
b111 6
19
1>
1C
b111 G
#493720000000
0!
1"
0*
1+
09
1:
0>
0C
#493730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#493740000000
0!
0*
09
0>
0C
#493750000000
1!
1*
b1 6
19
1>
1C
b1 G
#493760000000
0!
0*
09
0>
0C
#493770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#493780000000
0!
0*
09
0>
0C
#493790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#493800000000
0!
0*
09
0>
0C
#493810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#493820000000
0!
0*
09
0>
0C
#493830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#493840000000
0!
0#
0*
0,
09
0>
0?
0C
#493850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#493860000000
0!
0*
09
0>
0C
#493870000000
1!
1*
19
1>
1C
#493880000000
0!
0*
09
0>
0C
#493890000000
1!
1*
19
1>
1C
#493900000000
0!
0*
09
0>
0C
#493910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#493920000000
0!
0*
09
0>
0C
#493930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#493940000000
0!
0*
09
0>
0C
#493950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#493960000000
0!
0*
09
0>
0C
#493970000000
1!
1*
b10 6
19
1>
1C
b10 G
#493980000000
0!
0*
09
0>
0C
#493990000000
1!
1*
b11 6
19
1>
1C
b11 G
#494000000000
0!
0*
09
0>
0C
#494010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#494020000000
0!
0*
09
0>
0C
#494030000000
1!
1*
b101 6
19
1>
1C
b101 G
#494040000000
0!
0*
09
0>
0C
#494050000000
1!
1*
b110 6
19
1>
1C
b110 G
#494060000000
0!
0*
09
0>
0C
#494070000000
1!
1*
b111 6
19
1>
1C
b111 G
#494080000000
0!
0*
09
0>
0C
#494090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#494100000000
0!
0*
09
0>
0C
#494110000000
1!
1*
b1 6
19
1>
1C
b1 G
#494120000000
0!
0*
09
0>
0C
#494130000000
1!
1*
b10 6
19
1>
1C
b10 G
#494140000000
0!
0*
09
0>
0C
#494150000000
1!
1*
b11 6
19
1>
1C
b11 G
#494160000000
0!
0*
09
0>
0C
#494170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#494180000000
0!
0*
09
0>
0C
#494190000000
1!
1*
b101 6
19
1>
1C
b101 G
#494200000000
0!
0*
09
0>
0C
#494210000000
1!
1*
b110 6
19
1>
1C
b110 G
#494220000000
0!
0*
09
0>
0C
#494230000000
1!
1*
b111 6
19
1>
1C
b111 G
#494240000000
0!
0*
09
0>
0C
#494250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#494260000000
0!
0*
09
0>
0C
#494270000000
1!
1*
b1 6
19
1>
1C
b1 G
#494280000000
0!
0*
09
0>
0C
#494290000000
1!
1*
b10 6
19
1>
1C
b10 G
#494300000000
0!
0*
09
0>
0C
#494310000000
1!
1*
b11 6
19
1>
1C
b11 G
#494320000000
0!
0*
09
0>
0C
#494330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#494340000000
0!
0*
09
0>
0C
#494350000000
1!
1*
b101 6
19
1>
1C
b101 G
#494360000000
0!
0*
09
0>
0C
#494370000000
1!
1*
b110 6
19
1>
1C
b110 G
#494380000000
0!
0*
09
0>
0C
#494390000000
1!
1*
b111 6
19
1>
1C
b111 G
#494400000000
0!
1"
0*
1+
09
1:
0>
0C
#494410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#494420000000
0!
0*
09
0>
0C
#494430000000
1!
1*
b1 6
19
1>
1C
b1 G
#494440000000
0!
0*
09
0>
0C
#494450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#494460000000
0!
0*
09
0>
0C
#494470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#494480000000
0!
0*
09
0>
0C
#494490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#494500000000
0!
0*
09
0>
0C
#494510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#494520000000
0!
0#
0*
0,
09
0>
0?
0C
#494530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#494540000000
0!
0*
09
0>
0C
#494550000000
1!
1*
19
1>
1C
#494560000000
0!
0*
09
0>
0C
#494570000000
1!
1*
19
1>
1C
#494580000000
0!
0*
09
0>
0C
#494590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#494600000000
0!
0*
09
0>
0C
#494610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#494620000000
0!
0*
09
0>
0C
#494630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#494640000000
0!
0*
09
0>
0C
#494650000000
1!
1*
b10 6
19
1>
1C
b10 G
#494660000000
0!
0*
09
0>
0C
#494670000000
1!
1*
b11 6
19
1>
1C
b11 G
#494680000000
0!
0*
09
0>
0C
#494690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#494700000000
0!
0*
09
0>
0C
#494710000000
1!
1*
b101 6
19
1>
1C
b101 G
#494720000000
0!
0*
09
0>
0C
#494730000000
1!
1*
b110 6
19
1>
1C
b110 G
#494740000000
0!
0*
09
0>
0C
#494750000000
1!
1*
b111 6
19
1>
1C
b111 G
#494760000000
0!
0*
09
0>
0C
#494770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#494780000000
0!
0*
09
0>
0C
#494790000000
1!
1*
b1 6
19
1>
1C
b1 G
#494800000000
0!
0*
09
0>
0C
#494810000000
1!
1*
b10 6
19
1>
1C
b10 G
#494820000000
0!
0*
09
0>
0C
#494830000000
1!
1*
b11 6
19
1>
1C
b11 G
#494840000000
0!
0*
09
0>
0C
#494850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#494860000000
0!
0*
09
0>
0C
#494870000000
1!
1*
b101 6
19
1>
1C
b101 G
#494880000000
0!
0*
09
0>
0C
#494890000000
1!
1*
b110 6
19
1>
1C
b110 G
#494900000000
0!
0*
09
0>
0C
#494910000000
1!
1*
b111 6
19
1>
1C
b111 G
#494920000000
0!
0*
09
0>
0C
#494930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#494940000000
0!
0*
09
0>
0C
#494950000000
1!
1*
b1 6
19
1>
1C
b1 G
#494960000000
0!
0*
09
0>
0C
#494970000000
1!
1*
b10 6
19
1>
1C
b10 G
#494980000000
0!
0*
09
0>
0C
#494990000000
1!
1*
b11 6
19
1>
1C
b11 G
#495000000000
0!
0*
09
0>
0C
#495010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#495020000000
0!
0*
09
0>
0C
#495030000000
1!
1*
b101 6
19
1>
1C
b101 G
#495040000000
0!
0*
09
0>
0C
#495050000000
1!
1*
b110 6
19
1>
1C
b110 G
#495060000000
0!
0*
09
0>
0C
#495070000000
1!
1*
b111 6
19
1>
1C
b111 G
#495080000000
0!
1"
0*
1+
09
1:
0>
0C
#495090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#495100000000
0!
0*
09
0>
0C
#495110000000
1!
1*
b1 6
19
1>
1C
b1 G
#495120000000
0!
0*
09
0>
0C
#495130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#495140000000
0!
0*
09
0>
0C
#495150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#495160000000
0!
0*
09
0>
0C
#495170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#495180000000
0!
0*
09
0>
0C
#495190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#495200000000
0!
0#
0*
0,
09
0>
0?
0C
#495210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#495220000000
0!
0*
09
0>
0C
#495230000000
1!
1*
19
1>
1C
#495240000000
0!
0*
09
0>
0C
#495250000000
1!
1*
19
1>
1C
#495260000000
0!
0*
09
0>
0C
#495270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#495280000000
0!
0*
09
0>
0C
#495290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#495300000000
0!
0*
09
0>
0C
#495310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#495320000000
0!
0*
09
0>
0C
#495330000000
1!
1*
b10 6
19
1>
1C
b10 G
#495340000000
0!
0*
09
0>
0C
#495350000000
1!
1*
b11 6
19
1>
1C
b11 G
#495360000000
0!
0*
09
0>
0C
#495370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#495380000000
0!
0*
09
0>
0C
#495390000000
1!
1*
b101 6
19
1>
1C
b101 G
#495400000000
0!
0*
09
0>
0C
#495410000000
1!
1*
b110 6
19
1>
1C
b110 G
#495420000000
0!
0*
09
0>
0C
#495430000000
1!
1*
b111 6
19
1>
1C
b111 G
#495440000000
0!
0*
09
0>
0C
#495450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#495460000000
0!
0*
09
0>
0C
#495470000000
1!
1*
b1 6
19
1>
1C
b1 G
#495480000000
0!
0*
09
0>
0C
#495490000000
1!
1*
b10 6
19
1>
1C
b10 G
#495500000000
0!
0*
09
0>
0C
#495510000000
1!
1*
b11 6
19
1>
1C
b11 G
#495520000000
0!
0*
09
0>
0C
#495530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#495540000000
0!
0*
09
0>
0C
#495550000000
1!
1*
b101 6
19
1>
1C
b101 G
#495560000000
0!
0*
09
0>
0C
#495570000000
1!
1*
b110 6
19
1>
1C
b110 G
#495580000000
0!
0*
09
0>
0C
#495590000000
1!
1*
b111 6
19
1>
1C
b111 G
#495600000000
0!
0*
09
0>
0C
#495610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#495620000000
0!
0*
09
0>
0C
#495630000000
1!
1*
b1 6
19
1>
1C
b1 G
#495640000000
0!
0*
09
0>
0C
#495650000000
1!
1*
b10 6
19
1>
1C
b10 G
#495660000000
0!
0*
09
0>
0C
#495670000000
1!
1*
b11 6
19
1>
1C
b11 G
#495680000000
0!
0*
09
0>
0C
#495690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#495700000000
0!
0*
09
0>
0C
#495710000000
1!
1*
b101 6
19
1>
1C
b101 G
#495720000000
0!
0*
09
0>
0C
#495730000000
1!
1*
b110 6
19
1>
1C
b110 G
#495740000000
0!
0*
09
0>
0C
#495750000000
1!
1*
b111 6
19
1>
1C
b111 G
#495760000000
0!
1"
0*
1+
09
1:
0>
0C
#495770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#495780000000
0!
0*
09
0>
0C
#495790000000
1!
1*
b1 6
19
1>
1C
b1 G
#495800000000
0!
0*
09
0>
0C
#495810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#495820000000
0!
0*
09
0>
0C
#495830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#495840000000
0!
0*
09
0>
0C
#495850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#495860000000
0!
0*
09
0>
0C
#495870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#495880000000
0!
0#
0*
0,
09
0>
0?
0C
#495890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#495900000000
0!
0*
09
0>
0C
#495910000000
1!
1*
19
1>
1C
#495920000000
0!
0*
09
0>
0C
#495930000000
1!
1*
19
1>
1C
#495940000000
0!
0*
09
0>
0C
#495950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#495960000000
0!
0*
09
0>
0C
#495970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#495980000000
0!
0*
09
0>
0C
#495990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#496000000000
0!
0*
09
0>
0C
#496010000000
1!
1*
b10 6
19
1>
1C
b10 G
#496020000000
0!
0*
09
0>
0C
#496030000000
1!
1*
b11 6
19
1>
1C
b11 G
#496040000000
0!
0*
09
0>
0C
#496050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#496060000000
0!
0*
09
0>
0C
#496070000000
1!
1*
b101 6
19
1>
1C
b101 G
#496080000000
0!
0*
09
0>
0C
#496090000000
1!
1*
b110 6
19
1>
1C
b110 G
#496100000000
0!
0*
09
0>
0C
#496110000000
1!
1*
b111 6
19
1>
1C
b111 G
#496120000000
0!
0*
09
0>
0C
#496130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#496140000000
0!
0*
09
0>
0C
#496150000000
1!
1*
b1 6
19
1>
1C
b1 G
#496160000000
0!
0*
09
0>
0C
#496170000000
1!
1*
b10 6
19
1>
1C
b10 G
#496180000000
0!
0*
09
0>
0C
#496190000000
1!
1*
b11 6
19
1>
1C
b11 G
#496200000000
0!
0*
09
0>
0C
#496210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#496220000000
0!
0*
09
0>
0C
#496230000000
1!
1*
b101 6
19
1>
1C
b101 G
#496240000000
0!
0*
09
0>
0C
#496250000000
1!
1*
b110 6
19
1>
1C
b110 G
#496260000000
0!
0*
09
0>
0C
#496270000000
1!
1*
b111 6
19
1>
1C
b111 G
#496280000000
0!
0*
09
0>
0C
#496290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#496300000000
0!
0*
09
0>
0C
#496310000000
1!
1*
b1 6
19
1>
1C
b1 G
#496320000000
0!
0*
09
0>
0C
#496330000000
1!
1*
b10 6
19
1>
1C
b10 G
#496340000000
0!
0*
09
0>
0C
#496350000000
1!
1*
b11 6
19
1>
1C
b11 G
#496360000000
0!
0*
09
0>
0C
#496370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#496380000000
0!
0*
09
0>
0C
#496390000000
1!
1*
b101 6
19
1>
1C
b101 G
#496400000000
0!
0*
09
0>
0C
#496410000000
1!
1*
b110 6
19
1>
1C
b110 G
#496420000000
0!
0*
09
0>
0C
#496430000000
1!
1*
b111 6
19
1>
1C
b111 G
#496440000000
0!
1"
0*
1+
09
1:
0>
0C
#496450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#496460000000
0!
0*
09
0>
0C
#496470000000
1!
1*
b1 6
19
1>
1C
b1 G
#496480000000
0!
0*
09
0>
0C
#496490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#496500000000
0!
0*
09
0>
0C
#496510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#496520000000
0!
0*
09
0>
0C
#496530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#496540000000
0!
0*
09
0>
0C
#496550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#496560000000
0!
0#
0*
0,
09
0>
0?
0C
#496570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#496580000000
0!
0*
09
0>
0C
#496590000000
1!
1*
19
1>
1C
#496600000000
0!
0*
09
0>
0C
#496610000000
1!
1*
19
1>
1C
#496620000000
0!
0*
09
0>
0C
#496630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#496640000000
0!
0*
09
0>
0C
#496650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#496660000000
0!
0*
09
0>
0C
#496670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#496680000000
0!
0*
09
0>
0C
#496690000000
1!
1*
b10 6
19
1>
1C
b10 G
#496700000000
0!
0*
09
0>
0C
#496710000000
1!
1*
b11 6
19
1>
1C
b11 G
#496720000000
0!
0*
09
0>
0C
#496730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#496740000000
0!
0*
09
0>
0C
#496750000000
1!
1*
b101 6
19
1>
1C
b101 G
#496760000000
0!
0*
09
0>
0C
#496770000000
1!
1*
b110 6
19
1>
1C
b110 G
#496780000000
0!
0*
09
0>
0C
#496790000000
1!
1*
b111 6
19
1>
1C
b111 G
#496800000000
0!
0*
09
0>
0C
#496810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#496820000000
0!
0*
09
0>
0C
#496830000000
1!
1*
b1 6
19
1>
1C
b1 G
#496840000000
0!
0*
09
0>
0C
#496850000000
1!
1*
b10 6
19
1>
1C
b10 G
#496860000000
0!
0*
09
0>
0C
#496870000000
1!
1*
b11 6
19
1>
1C
b11 G
#496880000000
0!
0*
09
0>
0C
#496890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#496900000000
0!
0*
09
0>
0C
#496910000000
1!
1*
b101 6
19
1>
1C
b101 G
#496920000000
0!
0*
09
0>
0C
#496930000000
1!
1*
b110 6
19
1>
1C
b110 G
#496940000000
0!
0*
09
0>
0C
#496950000000
1!
1*
b111 6
19
1>
1C
b111 G
#496960000000
0!
0*
09
0>
0C
#496970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#496980000000
0!
0*
09
0>
0C
#496990000000
1!
1*
b1 6
19
1>
1C
b1 G
#497000000000
0!
0*
09
0>
0C
#497010000000
1!
1*
b10 6
19
1>
1C
b10 G
#497020000000
0!
0*
09
0>
0C
#497030000000
1!
1*
b11 6
19
1>
1C
b11 G
#497040000000
0!
0*
09
0>
0C
#497050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#497060000000
0!
0*
09
0>
0C
#497070000000
1!
1*
b101 6
19
1>
1C
b101 G
#497080000000
0!
0*
09
0>
0C
#497090000000
1!
1*
b110 6
19
1>
1C
b110 G
#497100000000
0!
0*
09
0>
0C
#497110000000
1!
1*
b111 6
19
1>
1C
b111 G
#497120000000
0!
1"
0*
1+
09
1:
0>
0C
#497130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#497140000000
0!
0*
09
0>
0C
#497150000000
1!
1*
b1 6
19
1>
1C
b1 G
#497160000000
0!
0*
09
0>
0C
#497170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#497180000000
0!
0*
09
0>
0C
#497190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#497200000000
0!
0*
09
0>
0C
#497210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#497220000000
0!
0*
09
0>
0C
#497230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#497240000000
0!
0#
0*
0,
09
0>
0?
0C
#497250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#497260000000
0!
0*
09
0>
0C
#497270000000
1!
1*
19
1>
1C
#497280000000
0!
0*
09
0>
0C
#497290000000
1!
1*
19
1>
1C
#497300000000
0!
0*
09
0>
0C
#497310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#497320000000
0!
0*
09
0>
0C
#497330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#497340000000
0!
0*
09
0>
0C
#497350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#497360000000
0!
0*
09
0>
0C
#497370000000
1!
1*
b10 6
19
1>
1C
b10 G
#497380000000
0!
0*
09
0>
0C
#497390000000
1!
1*
b11 6
19
1>
1C
b11 G
#497400000000
0!
0*
09
0>
0C
#497410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#497420000000
0!
0*
09
0>
0C
#497430000000
1!
1*
b101 6
19
1>
1C
b101 G
#497440000000
0!
0*
09
0>
0C
#497450000000
1!
1*
b110 6
19
1>
1C
b110 G
#497460000000
0!
0*
09
0>
0C
#497470000000
1!
1*
b111 6
19
1>
1C
b111 G
#497480000000
0!
0*
09
0>
0C
#497490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#497500000000
0!
0*
09
0>
0C
#497510000000
1!
1*
b1 6
19
1>
1C
b1 G
#497520000000
0!
0*
09
0>
0C
#497530000000
1!
1*
b10 6
19
1>
1C
b10 G
#497540000000
0!
0*
09
0>
0C
#497550000000
1!
1*
b11 6
19
1>
1C
b11 G
#497560000000
0!
0*
09
0>
0C
#497570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#497580000000
0!
0*
09
0>
0C
#497590000000
1!
1*
b101 6
19
1>
1C
b101 G
#497600000000
0!
0*
09
0>
0C
#497610000000
1!
1*
b110 6
19
1>
1C
b110 G
#497620000000
0!
0*
09
0>
0C
#497630000000
1!
1*
b111 6
19
1>
1C
b111 G
#497640000000
0!
0*
09
0>
0C
#497650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#497660000000
0!
0*
09
0>
0C
#497670000000
1!
1*
b1 6
19
1>
1C
b1 G
#497680000000
0!
0*
09
0>
0C
#497690000000
1!
1*
b10 6
19
1>
1C
b10 G
#497700000000
0!
0*
09
0>
0C
#497710000000
1!
1*
b11 6
19
1>
1C
b11 G
#497720000000
0!
0*
09
0>
0C
#497730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#497740000000
0!
0*
09
0>
0C
#497750000000
1!
1*
b101 6
19
1>
1C
b101 G
#497760000000
0!
0*
09
0>
0C
#497770000000
1!
1*
b110 6
19
1>
1C
b110 G
#497780000000
0!
0*
09
0>
0C
#497790000000
1!
1*
b111 6
19
1>
1C
b111 G
#497800000000
0!
1"
0*
1+
09
1:
0>
0C
#497810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#497820000000
0!
0*
09
0>
0C
#497830000000
1!
1*
b1 6
19
1>
1C
b1 G
#497840000000
0!
0*
09
0>
0C
#497850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#497860000000
0!
0*
09
0>
0C
#497870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#497880000000
0!
0*
09
0>
0C
#497890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#497900000000
0!
0*
09
0>
0C
#497910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#497920000000
0!
0#
0*
0,
09
0>
0?
0C
#497930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#497940000000
0!
0*
09
0>
0C
#497950000000
1!
1*
19
1>
1C
#497960000000
0!
0*
09
0>
0C
#497970000000
1!
1*
19
1>
1C
#497980000000
0!
0*
09
0>
0C
#497990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#498000000000
0!
0*
09
0>
0C
#498010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#498020000000
0!
0*
09
0>
0C
#498030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#498040000000
0!
0*
09
0>
0C
#498050000000
1!
1*
b10 6
19
1>
1C
b10 G
#498060000000
0!
0*
09
0>
0C
#498070000000
1!
1*
b11 6
19
1>
1C
b11 G
#498080000000
0!
0*
09
0>
0C
#498090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#498100000000
0!
0*
09
0>
0C
#498110000000
1!
1*
b101 6
19
1>
1C
b101 G
#498120000000
0!
0*
09
0>
0C
#498130000000
1!
1*
b110 6
19
1>
1C
b110 G
#498140000000
0!
0*
09
0>
0C
#498150000000
1!
1*
b111 6
19
1>
1C
b111 G
#498160000000
0!
0*
09
0>
0C
#498170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#498180000000
0!
0*
09
0>
0C
#498190000000
1!
1*
b1 6
19
1>
1C
b1 G
#498200000000
0!
0*
09
0>
0C
#498210000000
1!
1*
b10 6
19
1>
1C
b10 G
#498220000000
0!
0*
09
0>
0C
#498230000000
1!
1*
b11 6
19
1>
1C
b11 G
#498240000000
0!
0*
09
0>
0C
#498250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#498260000000
0!
0*
09
0>
0C
#498270000000
1!
1*
b101 6
19
1>
1C
b101 G
#498280000000
0!
0*
09
0>
0C
#498290000000
1!
1*
b110 6
19
1>
1C
b110 G
#498300000000
0!
0*
09
0>
0C
#498310000000
1!
1*
b111 6
19
1>
1C
b111 G
#498320000000
0!
0*
09
0>
0C
#498330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#498340000000
0!
0*
09
0>
0C
#498350000000
1!
1*
b1 6
19
1>
1C
b1 G
#498360000000
0!
0*
09
0>
0C
#498370000000
1!
1*
b10 6
19
1>
1C
b10 G
#498380000000
0!
0*
09
0>
0C
#498390000000
1!
1*
b11 6
19
1>
1C
b11 G
#498400000000
0!
0*
09
0>
0C
#498410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#498420000000
0!
0*
09
0>
0C
#498430000000
1!
1*
b101 6
19
1>
1C
b101 G
#498440000000
0!
0*
09
0>
0C
#498450000000
1!
1*
b110 6
19
1>
1C
b110 G
#498460000000
0!
0*
09
0>
0C
#498470000000
1!
1*
b111 6
19
1>
1C
b111 G
#498480000000
0!
1"
0*
1+
09
1:
0>
0C
#498490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#498500000000
0!
0*
09
0>
0C
#498510000000
1!
1*
b1 6
19
1>
1C
b1 G
#498520000000
0!
0*
09
0>
0C
#498530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#498540000000
0!
0*
09
0>
0C
#498550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#498560000000
0!
0*
09
0>
0C
#498570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#498580000000
0!
0*
09
0>
0C
#498590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#498600000000
0!
0#
0*
0,
09
0>
0?
0C
#498610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#498620000000
0!
0*
09
0>
0C
#498630000000
1!
1*
19
1>
1C
#498640000000
0!
0*
09
0>
0C
#498650000000
1!
1*
19
1>
1C
#498660000000
0!
0*
09
0>
0C
#498670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#498680000000
0!
0*
09
0>
0C
#498690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#498700000000
0!
0*
09
0>
0C
#498710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#498720000000
0!
0*
09
0>
0C
#498730000000
1!
1*
b10 6
19
1>
1C
b10 G
#498740000000
0!
0*
09
0>
0C
#498750000000
1!
1*
b11 6
19
1>
1C
b11 G
#498760000000
0!
0*
09
0>
0C
#498770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#498780000000
0!
0*
09
0>
0C
#498790000000
1!
1*
b101 6
19
1>
1C
b101 G
#498800000000
0!
0*
09
0>
0C
#498810000000
1!
1*
b110 6
19
1>
1C
b110 G
#498820000000
0!
0*
09
0>
0C
#498830000000
1!
1*
b111 6
19
1>
1C
b111 G
#498840000000
0!
0*
09
0>
0C
#498850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#498860000000
0!
0*
09
0>
0C
#498870000000
1!
1*
b1 6
19
1>
1C
b1 G
#498880000000
0!
0*
09
0>
0C
#498890000000
1!
1*
b10 6
19
1>
1C
b10 G
#498900000000
0!
0*
09
0>
0C
#498910000000
1!
1*
b11 6
19
1>
1C
b11 G
#498920000000
0!
0*
09
0>
0C
#498930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#498940000000
0!
0*
09
0>
0C
#498950000000
1!
1*
b101 6
19
1>
1C
b101 G
#498960000000
0!
0*
09
0>
0C
#498970000000
1!
1*
b110 6
19
1>
1C
b110 G
#498980000000
0!
0*
09
0>
0C
#498990000000
1!
1*
b111 6
19
1>
1C
b111 G
#499000000000
0!
0*
09
0>
0C
#499010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#499020000000
0!
0*
09
0>
0C
#499030000000
1!
1*
b1 6
19
1>
1C
b1 G
#499040000000
0!
0*
09
0>
0C
#499050000000
1!
1*
b10 6
19
1>
1C
b10 G
#499060000000
0!
0*
09
0>
0C
#499070000000
1!
1*
b11 6
19
1>
1C
b11 G
#499080000000
0!
0*
09
0>
0C
#499090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#499100000000
0!
0*
09
0>
0C
#499110000000
1!
1*
b101 6
19
1>
1C
b101 G
#499120000000
0!
0*
09
0>
0C
#499130000000
1!
1*
b110 6
19
1>
1C
b110 G
#499140000000
0!
0*
09
0>
0C
#499150000000
1!
1*
b111 6
19
1>
1C
b111 G
#499160000000
0!
1"
0*
1+
09
1:
0>
0C
#499170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#499180000000
0!
0*
09
0>
0C
#499190000000
1!
1*
b1 6
19
1>
1C
b1 G
#499200000000
0!
0*
09
0>
0C
#499210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#499220000000
0!
0*
09
0>
0C
#499230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#499240000000
0!
0*
09
0>
0C
#499250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#499260000000
0!
0*
09
0>
0C
#499270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#499280000000
0!
0#
0*
0,
09
0>
0?
0C
#499290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#499300000000
0!
0*
09
0>
0C
#499310000000
1!
1*
19
1>
1C
#499320000000
0!
0*
09
0>
0C
#499330000000
1!
1*
19
1>
1C
#499340000000
0!
0*
09
0>
0C
#499350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#499360000000
0!
0*
09
0>
0C
#499370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#499380000000
0!
0*
09
0>
0C
#499390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#499400000000
0!
0*
09
0>
0C
#499410000000
1!
1*
b10 6
19
1>
1C
b10 G
#499420000000
0!
0*
09
0>
0C
#499430000000
1!
1*
b11 6
19
1>
1C
b11 G
#499440000000
0!
0*
09
0>
0C
#499450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#499460000000
0!
0*
09
0>
0C
#499470000000
1!
1*
b101 6
19
1>
1C
b101 G
#499480000000
0!
0*
09
0>
0C
#499490000000
1!
1*
b110 6
19
1>
1C
b110 G
#499500000000
0!
0*
09
0>
0C
#499510000000
1!
1*
b111 6
19
1>
1C
b111 G
#499520000000
0!
0*
09
0>
0C
#499530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#499540000000
0!
0*
09
0>
0C
#499550000000
1!
1*
b1 6
19
1>
1C
b1 G
#499560000000
0!
0*
09
0>
0C
#499570000000
1!
1*
b10 6
19
1>
1C
b10 G
#499580000000
0!
0*
09
0>
0C
#499590000000
1!
1*
b11 6
19
1>
1C
b11 G
#499600000000
0!
0*
09
0>
0C
#499610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#499620000000
0!
0*
09
0>
0C
#499630000000
1!
1*
b101 6
19
1>
1C
b101 G
#499640000000
0!
0*
09
0>
0C
#499650000000
1!
1*
b110 6
19
1>
1C
b110 G
#499660000000
0!
0*
09
0>
0C
#499670000000
1!
1*
b111 6
19
1>
1C
b111 G
#499680000000
0!
0*
09
0>
0C
#499690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#499700000000
0!
0*
09
0>
0C
#499710000000
1!
1*
b1 6
19
1>
1C
b1 G
#499720000000
0!
0*
09
0>
0C
#499730000000
1!
1*
b10 6
19
1>
1C
b10 G
#499740000000
0!
0*
09
0>
0C
#499750000000
1!
1*
b11 6
19
1>
1C
b11 G
#499760000000
0!
0*
09
0>
0C
#499770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#499780000000
0!
0*
09
0>
0C
#499790000000
1!
1*
b101 6
19
1>
1C
b101 G
#499800000000
0!
0*
09
0>
0C
#499810000000
1!
1*
b110 6
19
1>
1C
b110 G
#499820000000
0!
0*
09
0>
0C
#499830000000
1!
1*
b111 6
19
1>
1C
b111 G
#499840000000
0!
1"
0*
1+
09
1:
0>
0C
#499850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#499860000000
0!
0*
09
0>
0C
#499870000000
1!
1*
b1 6
19
1>
1C
b1 G
#499880000000
0!
0*
09
0>
0C
#499890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#499900000000
0!
0*
09
0>
0C
#499910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#499920000000
0!
0*
09
0>
0C
#499930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#499940000000
0!
0*
09
0>
0C
#499950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#499960000000
0!
0#
0*
0,
09
0>
0?
0C
#499970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#499980000000
0!
0*
09
0>
0C
#499990000000
1!
1*
19
1>
1C
#500000000000
0!
0*
09
0>
0C
#500010000000
1!
1*
19
1>
1C
#500020000000
0!
0*
09
0>
0C
#500030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#500040000000
0!
0*
09
0>
0C
#500050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#500060000000
0!
0*
09
0>
0C
#500070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#500080000000
0!
0*
09
0>
0C
#500090000000
1!
1*
b10 6
19
1>
1C
b10 G
#500100000000
0!
0*
09
0>
0C
#500110000000
1!
1*
b11 6
19
1>
1C
b11 G
#500120000000
0!
0*
09
0>
0C
#500130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#500140000000
0!
0*
09
0>
0C
#500150000000
1!
1*
b101 6
19
1>
1C
b101 G
#500160000000
0!
0*
09
0>
0C
#500170000000
1!
1*
b110 6
19
1>
1C
b110 G
#500180000000
0!
0*
09
0>
0C
#500190000000
1!
1*
b111 6
19
1>
1C
b111 G
#500200000000
0!
0*
09
0>
0C
#500210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#500220000000
0!
0*
09
0>
0C
#500230000000
1!
1*
b1 6
19
1>
1C
b1 G
#500240000000
0!
0*
09
0>
0C
#500250000000
1!
1*
b10 6
19
1>
1C
b10 G
#500260000000
0!
0*
09
0>
0C
#500270000000
1!
1*
b11 6
19
1>
1C
b11 G
#500280000000
0!
0*
09
0>
0C
#500290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#500300000000
0!
0*
09
0>
0C
#500310000000
1!
1*
b101 6
19
1>
1C
b101 G
#500320000000
0!
0*
09
0>
0C
#500330000000
1!
1*
b110 6
19
1>
1C
b110 G
#500340000000
0!
0*
09
0>
0C
#500350000000
1!
1*
b111 6
19
1>
1C
b111 G
#500360000000
0!
0*
09
0>
0C
#500370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#500380000000
0!
0*
09
0>
0C
#500390000000
1!
1*
b1 6
19
1>
1C
b1 G
#500400000000
0!
0*
09
0>
0C
#500410000000
1!
1*
b10 6
19
1>
1C
b10 G
#500420000000
0!
0*
09
0>
0C
#500430000000
1!
1*
b11 6
19
1>
1C
b11 G
#500440000000
0!
0*
09
0>
0C
#500450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#500460000000
0!
0*
09
0>
0C
#500470000000
1!
1*
b101 6
19
1>
1C
b101 G
#500480000000
0!
0*
09
0>
0C
#500490000000
1!
1*
b110 6
19
1>
1C
b110 G
#500500000000
0!
0*
09
0>
0C
#500510000000
1!
1*
b111 6
19
1>
1C
b111 G
#500520000000
0!
1"
0*
1+
09
1:
0>
0C
#500530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#500540000000
0!
0*
09
0>
0C
#500550000000
1!
1*
b1 6
19
1>
1C
b1 G
#500560000000
0!
0*
09
0>
0C
#500570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#500580000000
0!
0*
09
0>
0C
#500590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#500600000000
0!
0*
09
0>
0C
#500610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#500620000000
0!
0*
09
0>
0C
#500630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#500640000000
0!
0#
0*
0,
09
0>
0?
0C
#500650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#500660000000
0!
0*
09
0>
0C
#500670000000
1!
1*
19
1>
1C
#500680000000
0!
0*
09
0>
0C
#500690000000
1!
1*
19
1>
1C
#500700000000
0!
0*
09
0>
0C
#500710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#500720000000
0!
0*
09
0>
0C
#500730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#500740000000
0!
0*
09
0>
0C
#500750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#500760000000
0!
0*
09
0>
0C
#500770000000
1!
1*
b10 6
19
1>
1C
b10 G
#500780000000
0!
0*
09
0>
0C
#500790000000
1!
1*
b11 6
19
1>
1C
b11 G
#500800000000
0!
0*
09
0>
0C
#500810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#500820000000
0!
0*
09
0>
0C
#500830000000
1!
1*
b101 6
19
1>
1C
b101 G
#500840000000
0!
0*
09
0>
0C
#500850000000
1!
1*
b110 6
19
1>
1C
b110 G
#500860000000
0!
0*
09
0>
0C
#500870000000
1!
1*
b111 6
19
1>
1C
b111 G
#500880000000
0!
0*
09
0>
0C
#500890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#500900000000
0!
0*
09
0>
0C
#500910000000
1!
1*
b1 6
19
1>
1C
b1 G
#500920000000
0!
0*
09
0>
0C
#500930000000
1!
1*
b10 6
19
1>
1C
b10 G
#500940000000
0!
0*
09
0>
0C
#500950000000
1!
1*
b11 6
19
1>
1C
b11 G
#500960000000
0!
0*
09
0>
0C
#500970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#500980000000
0!
0*
09
0>
0C
#500990000000
1!
1*
b101 6
19
1>
1C
b101 G
#501000000000
0!
0*
09
0>
0C
#501010000000
1!
1*
b110 6
19
1>
1C
b110 G
#501020000000
0!
0*
09
0>
0C
#501030000000
1!
1*
b111 6
19
1>
1C
b111 G
#501040000000
0!
0*
09
0>
0C
#501050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#501060000000
0!
0*
09
0>
0C
#501070000000
1!
1*
b1 6
19
1>
1C
b1 G
#501080000000
0!
0*
09
0>
0C
#501090000000
1!
1*
b10 6
19
1>
1C
b10 G
#501100000000
0!
0*
09
0>
0C
#501110000000
1!
1*
b11 6
19
1>
1C
b11 G
#501120000000
0!
0*
09
0>
0C
#501130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#501140000000
0!
0*
09
0>
0C
#501150000000
1!
1*
b101 6
19
1>
1C
b101 G
#501160000000
0!
0*
09
0>
0C
#501170000000
1!
1*
b110 6
19
1>
1C
b110 G
#501180000000
0!
0*
09
0>
0C
#501190000000
1!
1*
b111 6
19
1>
1C
b111 G
#501200000000
0!
1"
0*
1+
09
1:
0>
0C
#501210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#501220000000
0!
0*
09
0>
0C
#501230000000
1!
1*
b1 6
19
1>
1C
b1 G
#501240000000
0!
0*
09
0>
0C
#501250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#501260000000
0!
0*
09
0>
0C
#501270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#501280000000
0!
0*
09
0>
0C
#501290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#501300000000
0!
0*
09
0>
0C
#501310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#501320000000
0!
0#
0*
0,
09
0>
0?
0C
#501330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#501340000000
0!
0*
09
0>
0C
#501350000000
1!
1*
19
1>
1C
#501360000000
0!
0*
09
0>
0C
#501370000000
1!
1*
19
1>
1C
#501380000000
0!
0*
09
0>
0C
#501390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#501400000000
0!
0*
09
0>
0C
#501410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#501420000000
0!
0*
09
0>
0C
#501430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#501440000000
0!
0*
09
0>
0C
#501450000000
1!
1*
b10 6
19
1>
1C
b10 G
#501460000000
0!
0*
09
0>
0C
#501470000000
1!
1*
b11 6
19
1>
1C
b11 G
#501480000000
0!
0*
09
0>
0C
#501490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#501500000000
0!
0*
09
0>
0C
#501510000000
1!
1*
b101 6
19
1>
1C
b101 G
#501520000000
0!
0*
09
0>
0C
#501530000000
1!
1*
b110 6
19
1>
1C
b110 G
#501540000000
0!
0*
09
0>
0C
#501550000000
1!
1*
b111 6
19
1>
1C
b111 G
#501560000000
0!
0*
09
0>
0C
#501570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#501580000000
0!
0*
09
0>
0C
#501590000000
1!
1*
b1 6
19
1>
1C
b1 G
#501600000000
0!
0*
09
0>
0C
#501610000000
1!
1*
b10 6
19
1>
1C
b10 G
#501620000000
0!
0*
09
0>
0C
#501630000000
1!
1*
b11 6
19
1>
1C
b11 G
#501640000000
0!
0*
09
0>
0C
#501650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#501660000000
0!
0*
09
0>
0C
#501670000000
1!
1*
b101 6
19
1>
1C
b101 G
#501680000000
0!
0*
09
0>
0C
#501690000000
1!
1*
b110 6
19
1>
1C
b110 G
#501700000000
0!
0*
09
0>
0C
#501710000000
1!
1*
b111 6
19
1>
1C
b111 G
#501720000000
0!
0*
09
0>
0C
#501730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#501740000000
0!
0*
09
0>
0C
#501750000000
1!
1*
b1 6
19
1>
1C
b1 G
#501760000000
0!
0*
09
0>
0C
#501770000000
1!
1*
b10 6
19
1>
1C
b10 G
#501780000000
0!
0*
09
0>
0C
#501790000000
1!
1*
b11 6
19
1>
1C
b11 G
#501800000000
0!
0*
09
0>
0C
#501810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#501820000000
0!
0*
09
0>
0C
#501830000000
1!
1*
b101 6
19
1>
1C
b101 G
#501840000000
0!
0*
09
0>
0C
#501850000000
1!
1*
b110 6
19
1>
1C
b110 G
#501860000000
0!
0*
09
0>
0C
#501870000000
1!
1*
b111 6
19
1>
1C
b111 G
#501880000000
0!
1"
0*
1+
09
1:
0>
0C
#501890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#501900000000
0!
0*
09
0>
0C
#501910000000
1!
1*
b1 6
19
1>
1C
b1 G
#501920000000
0!
0*
09
0>
0C
#501930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#501940000000
0!
0*
09
0>
0C
#501950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#501960000000
0!
0*
09
0>
0C
#501970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#501980000000
0!
0*
09
0>
0C
#501990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#502000000000
0!
0#
0*
0,
09
0>
0?
0C
#502010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#502020000000
0!
0*
09
0>
0C
#502030000000
1!
1*
19
1>
1C
#502040000000
0!
0*
09
0>
0C
#502050000000
1!
1*
19
1>
1C
#502060000000
0!
0*
09
0>
0C
#502070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#502080000000
0!
0*
09
0>
0C
#502090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#502100000000
0!
0*
09
0>
0C
#502110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#502120000000
0!
0*
09
0>
0C
#502130000000
1!
1*
b10 6
19
1>
1C
b10 G
#502140000000
0!
0*
09
0>
0C
#502150000000
1!
1*
b11 6
19
1>
1C
b11 G
#502160000000
0!
0*
09
0>
0C
#502170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#502180000000
0!
0*
09
0>
0C
#502190000000
1!
1*
b101 6
19
1>
1C
b101 G
#502200000000
0!
0*
09
0>
0C
#502210000000
1!
1*
b110 6
19
1>
1C
b110 G
#502220000000
0!
0*
09
0>
0C
#502230000000
1!
1*
b111 6
19
1>
1C
b111 G
#502240000000
0!
0*
09
0>
0C
#502250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#502260000000
0!
0*
09
0>
0C
#502270000000
1!
1*
b1 6
19
1>
1C
b1 G
#502280000000
0!
0*
09
0>
0C
#502290000000
1!
1*
b10 6
19
1>
1C
b10 G
#502300000000
0!
0*
09
0>
0C
#502310000000
1!
1*
b11 6
19
1>
1C
b11 G
#502320000000
0!
0*
09
0>
0C
#502330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#502340000000
0!
0*
09
0>
0C
#502350000000
1!
1*
b101 6
19
1>
1C
b101 G
#502360000000
0!
0*
09
0>
0C
#502370000000
1!
1*
b110 6
19
1>
1C
b110 G
#502380000000
0!
0*
09
0>
0C
#502390000000
1!
1*
b111 6
19
1>
1C
b111 G
#502400000000
0!
0*
09
0>
0C
#502410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#502420000000
0!
0*
09
0>
0C
#502430000000
1!
1*
b1 6
19
1>
1C
b1 G
#502440000000
0!
0*
09
0>
0C
#502450000000
1!
1*
b10 6
19
1>
1C
b10 G
#502460000000
0!
0*
09
0>
0C
#502470000000
1!
1*
b11 6
19
1>
1C
b11 G
#502480000000
0!
0*
09
0>
0C
#502490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#502500000000
0!
0*
09
0>
0C
#502510000000
1!
1*
b101 6
19
1>
1C
b101 G
#502520000000
0!
0*
09
0>
0C
#502530000000
1!
1*
b110 6
19
1>
1C
b110 G
#502540000000
0!
0*
09
0>
0C
#502550000000
1!
1*
b111 6
19
1>
1C
b111 G
#502560000000
0!
1"
0*
1+
09
1:
0>
0C
#502570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#502580000000
0!
0*
09
0>
0C
#502590000000
1!
1*
b1 6
19
1>
1C
b1 G
#502600000000
0!
0*
09
0>
0C
#502610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#502620000000
0!
0*
09
0>
0C
#502630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#502640000000
0!
0*
09
0>
0C
#502650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#502660000000
0!
0*
09
0>
0C
#502670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#502680000000
0!
0#
0*
0,
09
0>
0?
0C
#502690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#502700000000
0!
0*
09
0>
0C
#502710000000
1!
1*
19
1>
1C
#502720000000
0!
0*
09
0>
0C
#502730000000
1!
1*
19
1>
1C
#502740000000
0!
0*
09
0>
0C
#502750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#502760000000
0!
0*
09
0>
0C
#502770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#502780000000
0!
0*
09
0>
0C
#502790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#502800000000
0!
0*
09
0>
0C
#502810000000
1!
1*
b10 6
19
1>
1C
b10 G
#502820000000
0!
0*
09
0>
0C
#502830000000
1!
1*
b11 6
19
1>
1C
b11 G
#502840000000
0!
0*
09
0>
0C
#502850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#502860000000
0!
0*
09
0>
0C
#502870000000
1!
1*
b101 6
19
1>
1C
b101 G
#502880000000
0!
0*
09
0>
0C
#502890000000
1!
1*
b110 6
19
1>
1C
b110 G
#502900000000
0!
0*
09
0>
0C
#502910000000
1!
1*
b111 6
19
1>
1C
b111 G
#502920000000
0!
0*
09
0>
0C
#502930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#502940000000
0!
0*
09
0>
0C
#502950000000
1!
1*
b1 6
19
1>
1C
b1 G
#502960000000
0!
0*
09
0>
0C
#502970000000
1!
1*
b10 6
19
1>
1C
b10 G
#502980000000
0!
0*
09
0>
0C
#502990000000
1!
1*
b11 6
19
1>
1C
b11 G
#503000000000
0!
0*
09
0>
0C
#503010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#503020000000
0!
0*
09
0>
0C
#503030000000
1!
1*
b101 6
19
1>
1C
b101 G
#503040000000
0!
0*
09
0>
0C
#503050000000
1!
1*
b110 6
19
1>
1C
b110 G
#503060000000
0!
0*
09
0>
0C
#503070000000
1!
1*
b111 6
19
1>
1C
b111 G
#503080000000
0!
0*
09
0>
0C
#503090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#503100000000
0!
0*
09
0>
0C
#503110000000
1!
1*
b1 6
19
1>
1C
b1 G
#503120000000
0!
0*
09
0>
0C
#503130000000
1!
1*
b10 6
19
1>
1C
b10 G
#503140000000
0!
0*
09
0>
0C
#503150000000
1!
1*
b11 6
19
1>
1C
b11 G
#503160000000
0!
0*
09
0>
0C
#503170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#503180000000
0!
0*
09
0>
0C
#503190000000
1!
1*
b101 6
19
1>
1C
b101 G
#503200000000
0!
0*
09
0>
0C
#503210000000
1!
1*
b110 6
19
1>
1C
b110 G
#503220000000
0!
0*
09
0>
0C
#503230000000
1!
1*
b111 6
19
1>
1C
b111 G
#503240000000
0!
1"
0*
1+
09
1:
0>
0C
#503250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#503260000000
0!
0*
09
0>
0C
#503270000000
1!
1*
b1 6
19
1>
1C
b1 G
#503280000000
0!
0*
09
0>
0C
#503290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#503300000000
0!
0*
09
0>
0C
#503310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#503320000000
0!
0*
09
0>
0C
#503330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#503340000000
0!
0*
09
0>
0C
#503350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#503360000000
0!
0#
0*
0,
09
0>
0?
0C
#503370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#503380000000
0!
0*
09
0>
0C
#503390000000
1!
1*
19
1>
1C
#503400000000
0!
0*
09
0>
0C
#503410000000
1!
1*
19
1>
1C
#503420000000
0!
0*
09
0>
0C
#503430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#503440000000
0!
0*
09
0>
0C
#503450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#503460000000
0!
0*
09
0>
0C
#503470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#503480000000
0!
0*
09
0>
0C
#503490000000
1!
1*
b10 6
19
1>
1C
b10 G
#503500000000
0!
0*
09
0>
0C
#503510000000
1!
1*
b11 6
19
1>
1C
b11 G
#503520000000
0!
0*
09
0>
0C
#503530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#503540000000
0!
0*
09
0>
0C
#503550000000
1!
1*
b101 6
19
1>
1C
b101 G
#503560000000
0!
0*
09
0>
0C
#503570000000
1!
1*
b110 6
19
1>
1C
b110 G
#503580000000
0!
0*
09
0>
0C
#503590000000
1!
1*
b111 6
19
1>
1C
b111 G
#503600000000
0!
0*
09
0>
0C
#503610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#503620000000
0!
0*
09
0>
0C
#503630000000
1!
1*
b1 6
19
1>
1C
b1 G
#503640000000
0!
0*
09
0>
0C
#503650000000
1!
1*
b10 6
19
1>
1C
b10 G
#503660000000
0!
0*
09
0>
0C
#503670000000
1!
1*
b11 6
19
1>
1C
b11 G
#503680000000
0!
0*
09
0>
0C
#503690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#503700000000
0!
0*
09
0>
0C
#503710000000
1!
1*
b101 6
19
1>
1C
b101 G
#503720000000
0!
0*
09
0>
0C
#503730000000
1!
1*
b110 6
19
1>
1C
b110 G
#503740000000
0!
0*
09
0>
0C
#503750000000
1!
1*
b111 6
19
1>
1C
b111 G
#503760000000
0!
0*
09
0>
0C
#503770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#503780000000
0!
0*
09
0>
0C
#503790000000
1!
1*
b1 6
19
1>
1C
b1 G
#503800000000
0!
0*
09
0>
0C
#503810000000
1!
1*
b10 6
19
1>
1C
b10 G
#503820000000
0!
0*
09
0>
0C
#503830000000
1!
1*
b11 6
19
1>
1C
b11 G
#503840000000
0!
0*
09
0>
0C
#503850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#503860000000
0!
0*
09
0>
0C
#503870000000
1!
1*
b101 6
19
1>
1C
b101 G
#503880000000
0!
0*
09
0>
0C
#503890000000
1!
1*
b110 6
19
1>
1C
b110 G
#503900000000
0!
0*
09
0>
0C
#503910000000
1!
1*
b111 6
19
1>
1C
b111 G
#503920000000
0!
1"
0*
1+
09
1:
0>
0C
#503930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#503940000000
0!
0*
09
0>
0C
#503950000000
1!
1*
b1 6
19
1>
1C
b1 G
#503960000000
0!
0*
09
0>
0C
#503970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#503980000000
0!
0*
09
0>
0C
#503990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#504000000000
0!
0*
09
0>
0C
#504010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#504020000000
0!
0*
09
0>
0C
#504030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#504040000000
0!
0#
0*
0,
09
0>
0?
0C
#504050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#504060000000
0!
0*
09
0>
0C
#504070000000
1!
1*
19
1>
1C
#504080000000
0!
0*
09
0>
0C
#504090000000
1!
1*
19
1>
1C
#504100000000
0!
0*
09
0>
0C
#504110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#504120000000
0!
0*
09
0>
0C
#504130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#504140000000
0!
0*
09
0>
0C
#504150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#504160000000
0!
0*
09
0>
0C
#504170000000
1!
1*
b10 6
19
1>
1C
b10 G
#504180000000
0!
0*
09
0>
0C
#504190000000
1!
1*
b11 6
19
1>
1C
b11 G
#504200000000
0!
0*
09
0>
0C
#504210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#504220000000
0!
0*
09
0>
0C
#504230000000
1!
1*
b101 6
19
1>
1C
b101 G
#504240000000
0!
0*
09
0>
0C
#504250000000
1!
1*
b110 6
19
1>
1C
b110 G
#504260000000
0!
0*
09
0>
0C
#504270000000
1!
1*
b111 6
19
1>
1C
b111 G
#504280000000
0!
0*
09
0>
0C
#504290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#504300000000
0!
0*
09
0>
0C
#504310000000
1!
1*
b1 6
19
1>
1C
b1 G
#504320000000
0!
0*
09
0>
0C
#504330000000
1!
1*
b10 6
19
1>
1C
b10 G
#504340000000
0!
0*
09
0>
0C
#504350000000
1!
1*
b11 6
19
1>
1C
b11 G
#504360000000
0!
0*
09
0>
0C
#504370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#504380000000
0!
0*
09
0>
0C
#504390000000
1!
1*
b101 6
19
1>
1C
b101 G
#504400000000
0!
0*
09
0>
0C
#504410000000
1!
1*
b110 6
19
1>
1C
b110 G
#504420000000
0!
0*
09
0>
0C
#504430000000
1!
1*
b111 6
19
1>
1C
b111 G
#504440000000
0!
0*
09
0>
0C
#504450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#504460000000
0!
0*
09
0>
0C
#504470000000
1!
1*
b1 6
19
1>
1C
b1 G
#504480000000
0!
0*
09
0>
0C
#504490000000
1!
1*
b10 6
19
1>
1C
b10 G
#504500000000
0!
0*
09
0>
0C
#504510000000
1!
1*
b11 6
19
1>
1C
b11 G
#504520000000
0!
0*
09
0>
0C
#504530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#504540000000
0!
0*
09
0>
0C
#504550000000
1!
1*
b101 6
19
1>
1C
b101 G
#504560000000
0!
0*
09
0>
0C
#504570000000
1!
1*
b110 6
19
1>
1C
b110 G
#504580000000
0!
0*
09
0>
0C
#504590000000
1!
1*
b111 6
19
1>
1C
b111 G
#504600000000
0!
1"
0*
1+
09
1:
0>
0C
#504610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#504620000000
0!
0*
09
0>
0C
#504630000000
1!
1*
b1 6
19
1>
1C
b1 G
#504640000000
0!
0*
09
0>
0C
#504650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#504660000000
0!
0*
09
0>
0C
#504670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#504680000000
0!
0*
09
0>
0C
#504690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#504700000000
0!
0*
09
0>
0C
#504710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#504720000000
0!
0#
0*
0,
09
0>
0?
0C
#504730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#504740000000
0!
0*
09
0>
0C
#504750000000
1!
1*
19
1>
1C
#504760000000
0!
0*
09
0>
0C
#504770000000
1!
1*
19
1>
1C
#504780000000
0!
0*
09
0>
0C
#504790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#504800000000
0!
0*
09
0>
0C
#504810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#504820000000
0!
0*
09
0>
0C
#504830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#504840000000
0!
0*
09
0>
0C
#504850000000
1!
1*
b10 6
19
1>
1C
b10 G
#504860000000
0!
0*
09
0>
0C
#504870000000
1!
1*
b11 6
19
1>
1C
b11 G
#504880000000
0!
0*
09
0>
0C
#504890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#504900000000
0!
0*
09
0>
0C
#504910000000
1!
1*
b101 6
19
1>
1C
b101 G
#504920000000
0!
0*
09
0>
0C
#504930000000
1!
1*
b110 6
19
1>
1C
b110 G
#504940000000
0!
0*
09
0>
0C
#504950000000
1!
1*
b111 6
19
1>
1C
b111 G
#504960000000
0!
0*
09
0>
0C
#504970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#504980000000
0!
0*
09
0>
0C
#504990000000
1!
1*
b1 6
19
1>
1C
b1 G
#505000000000
0!
0*
09
0>
0C
#505010000000
1!
1*
b10 6
19
1>
1C
b10 G
#505020000000
0!
0*
09
0>
0C
#505030000000
1!
1*
b11 6
19
1>
1C
b11 G
#505040000000
0!
0*
09
0>
0C
#505050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#505060000000
0!
0*
09
0>
0C
#505070000000
1!
1*
b101 6
19
1>
1C
b101 G
#505080000000
0!
0*
09
0>
0C
#505090000000
1!
1*
b110 6
19
1>
1C
b110 G
#505100000000
0!
0*
09
0>
0C
#505110000000
1!
1*
b111 6
19
1>
1C
b111 G
#505120000000
0!
0*
09
0>
0C
#505130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#505140000000
0!
0*
09
0>
0C
#505150000000
1!
1*
b1 6
19
1>
1C
b1 G
#505160000000
0!
0*
09
0>
0C
#505170000000
1!
1*
b10 6
19
1>
1C
b10 G
#505180000000
0!
0*
09
0>
0C
#505190000000
1!
1*
b11 6
19
1>
1C
b11 G
#505200000000
0!
0*
09
0>
0C
#505210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#505220000000
0!
0*
09
0>
0C
#505230000000
1!
1*
b101 6
19
1>
1C
b101 G
#505240000000
0!
0*
09
0>
0C
#505250000000
1!
1*
b110 6
19
1>
1C
b110 G
#505260000000
0!
0*
09
0>
0C
#505270000000
1!
1*
b111 6
19
1>
1C
b111 G
#505280000000
0!
1"
0*
1+
09
1:
0>
0C
#505290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#505300000000
0!
0*
09
0>
0C
#505310000000
1!
1*
b1 6
19
1>
1C
b1 G
#505320000000
0!
0*
09
0>
0C
#505330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#505340000000
0!
0*
09
0>
0C
#505350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#505360000000
0!
0*
09
0>
0C
#505370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#505380000000
0!
0*
09
0>
0C
#505390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#505400000000
0!
0#
0*
0,
09
0>
0?
0C
#505410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#505420000000
0!
0*
09
0>
0C
#505430000000
1!
1*
19
1>
1C
#505440000000
0!
0*
09
0>
0C
#505450000000
1!
1*
19
1>
1C
#505460000000
0!
0*
09
0>
0C
#505470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#505480000000
0!
0*
09
0>
0C
#505490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#505500000000
0!
0*
09
0>
0C
#505510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#505520000000
0!
0*
09
0>
0C
#505530000000
1!
1*
b10 6
19
1>
1C
b10 G
#505540000000
0!
0*
09
0>
0C
#505550000000
1!
1*
b11 6
19
1>
1C
b11 G
#505560000000
0!
0*
09
0>
0C
#505570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#505580000000
0!
0*
09
0>
0C
#505590000000
1!
1*
b101 6
19
1>
1C
b101 G
#505600000000
0!
0*
09
0>
0C
#505610000000
1!
1*
b110 6
19
1>
1C
b110 G
#505620000000
0!
0*
09
0>
0C
#505630000000
1!
1*
b111 6
19
1>
1C
b111 G
#505640000000
0!
0*
09
0>
0C
#505650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#505660000000
0!
0*
09
0>
0C
#505670000000
1!
1*
b1 6
19
1>
1C
b1 G
#505680000000
0!
0*
09
0>
0C
#505690000000
1!
1*
b10 6
19
1>
1C
b10 G
#505700000000
0!
0*
09
0>
0C
#505710000000
1!
1*
b11 6
19
1>
1C
b11 G
#505720000000
0!
0*
09
0>
0C
#505730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#505740000000
0!
0*
09
0>
0C
#505750000000
1!
1*
b101 6
19
1>
1C
b101 G
#505760000000
0!
0*
09
0>
0C
#505770000000
1!
1*
b110 6
19
1>
1C
b110 G
#505780000000
0!
0*
09
0>
0C
#505790000000
1!
1*
b111 6
19
1>
1C
b111 G
#505800000000
0!
0*
09
0>
0C
#505810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#505820000000
0!
0*
09
0>
0C
#505830000000
1!
1*
b1 6
19
1>
1C
b1 G
#505840000000
0!
0*
09
0>
0C
#505850000000
1!
1*
b10 6
19
1>
1C
b10 G
#505860000000
0!
0*
09
0>
0C
#505870000000
1!
1*
b11 6
19
1>
1C
b11 G
#505880000000
0!
0*
09
0>
0C
#505890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#505900000000
0!
0*
09
0>
0C
#505910000000
1!
1*
b101 6
19
1>
1C
b101 G
#505920000000
0!
0*
09
0>
0C
#505930000000
1!
1*
b110 6
19
1>
1C
b110 G
#505940000000
0!
0*
09
0>
0C
#505950000000
1!
1*
b111 6
19
1>
1C
b111 G
#505960000000
0!
1"
0*
1+
09
1:
0>
0C
#505970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#505980000000
0!
0*
09
0>
0C
#505990000000
1!
1*
b1 6
19
1>
1C
b1 G
#506000000000
0!
0*
09
0>
0C
#506010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#506020000000
0!
0*
09
0>
0C
#506030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#506040000000
0!
0*
09
0>
0C
#506050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#506060000000
0!
0*
09
0>
0C
#506070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#506080000000
0!
0#
0*
0,
09
0>
0?
0C
#506090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#506100000000
0!
0*
09
0>
0C
#506110000000
1!
1*
19
1>
1C
#506120000000
0!
0*
09
0>
0C
#506130000000
1!
1*
19
1>
1C
#506140000000
0!
0*
09
0>
0C
#506150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#506160000000
0!
0*
09
0>
0C
#506170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#506180000000
0!
0*
09
0>
0C
#506190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#506200000000
0!
0*
09
0>
0C
#506210000000
1!
1*
b10 6
19
1>
1C
b10 G
#506220000000
0!
0*
09
0>
0C
#506230000000
1!
1*
b11 6
19
1>
1C
b11 G
#506240000000
0!
0*
09
0>
0C
#506250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#506260000000
0!
0*
09
0>
0C
#506270000000
1!
1*
b101 6
19
1>
1C
b101 G
#506280000000
0!
0*
09
0>
0C
#506290000000
1!
1*
b110 6
19
1>
1C
b110 G
#506300000000
0!
0*
09
0>
0C
#506310000000
1!
1*
b111 6
19
1>
1C
b111 G
#506320000000
0!
0*
09
0>
0C
#506330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#506340000000
0!
0*
09
0>
0C
#506350000000
1!
1*
b1 6
19
1>
1C
b1 G
#506360000000
0!
0*
09
0>
0C
#506370000000
1!
1*
b10 6
19
1>
1C
b10 G
#506380000000
0!
0*
09
0>
0C
#506390000000
1!
1*
b11 6
19
1>
1C
b11 G
#506400000000
0!
0*
09
0>
0C
#506410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#506420000000
0!
0*
09
0>
0C
#506430000000
1!
1*
b101 6
19
1>
1C
b101 G
#506440000000
0!
0*
09
0>
0C
#506450000000
1!
1*
b110 6
19
1>
1C
b110 G
#506460000000
0!
0*
09
0>
0C
#506470000000
1!
1*
b111 6
19
1>
1C
b111 G
#506480000000
0!
0*
09
0>
0C
#506490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#506500000000
0!
0*
09
0>
0C
#506510000000
1!
1*
b1 6
19
1>
1C
b1 G
#506520000000
0!
0*
09
0>
0C
#506530000000
1!
1*
b10 6
19
1>
1C
b10 G
#506540000000
0!
0*
09
0>
0C
#506550000000
1!
1*
b11 6
19
1>
1C
b11 G
#506560000000
0!
0*
09
0>
0C
#506570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#506580000000
0!
0*
09
0>
0C
#506590000000
1!
1*
b101 6
19
1>
1C
b101 G
#506600000000
0!
0*
09
0>
0C
#506610000000
1!
1*
b110 6
19
1>
1C
b110 G
#506620000000
0!
0*
09
0>
0C
#506630000000
1!
1*
b111 6
19
1>
1C
b111 G
#506640000000
0!
1"
0*
1+
09
1:
0>
0C
#506650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#506660000000
0!
0*
09
0>
0C
#506670000000
1!
1*
b1 6
19
1>
1C
b1 G
#506680000000
0!
0*
09
0>
0C
#506690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#506700000000
0!
0*
09
0>
0C
#506710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#506720000000
0!
0*
09
0>
0C
#506730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#506740000000
0!
0*
09
0>
0C
#506750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#506760000000
0!
0#
0*
0,
09
0>
0?
0C
#506770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#506780000000
0!
0*
09
0>
0C
#506790000000
1!
1*
19
1>
1C
#506800000000
0!
0*
09
0>
0C
#506810000000
1!
1*
19
1>
1C
#506820000000
0!
0*
09
0>
0C
#506830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#506840000000
0!
0*
09
0>
0C
#506850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#506860000000
0!
0*
09
0>
0C
#506870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#506880000000
0!
0*
09
0>
0C
#506890000000
1!
1*
b10 6
19
1>
1C
b10 G
#506900000000
0!
0*
09
0>
0C
#506910000000
1!
1*
b11 6
19
1>
1C
b11 G
#506920000000
0!
0*
09
0>
0C
#506930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#506940000000
0!
0*
09
0>
0C
#506950000000
1!
1*
b101 6
19
1>
1C
b101 G
#506960000000
0!
0*
09
0>
0C
#506970000000
1!
1*
b110 6
19
1>
1C
b110 G
#506980000000
0!
0*
09
0>
0C
#506990000000
1!
1*
b111 6
19
1>
1C
b111 G
#507000000000
0!
0*
09
0>
0C
#507010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#507020000000
0!
0*
09
0>
0C
#507030000000
1!
1*
b1 6
19
1>
1C
b1 G
#507040000000
0!
0*
09
0>
0C
#507050000000
1!
1*
b10 6
19
1>
1C
b10 G
#507060000000
0!
0*
09
0>
0C
#507070000000
1!
1*
b11 6
19
1>
1C
b11 G
#507080000000
0!
0*
09
0>
0C
#507090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#507100000000
0!
0*
09
0>
0C
#507110000000
1!
1*
b101 6
19
1>
1C
b101 G
#507120000000
0!
0*
09
0>
0C
#507130000000
1!
1*
b110 6
19
1>
1C
b110 G
#507140000000
0!
0*
09
0>
0C
#507150000000
1!
1*
b111 6
19
1>
1C
b111 G
#507160000000
0!
0*
09
0>
0C
#507170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#507180000000
0!
0*
09
0>
0C
#507190000000
1!
1*
b1 6
19
1>
1C
b1 G
#507200000000
0!
0*
09
0>
0C
#507210000000
1!
1*
b10 6
19
1>
1C
b10 G
#507220000000
0!
0*
09
0>
0C
#507230000000
1!
1*
b11 6
19
1>
1C
b11 G
#507240000000
0!
0*
09
0>
0C
#507250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#507260000000
0!
0*
09
0>
0C
#507270000000
1!
1*
b101 6
19
1>
1C
b101 G
#507280000000
0!
0*
09
0>
0C
#507290000000
1!
1*
b110 6
19
1>
1C
b110 G
#507300000000
0!
0*
09
0>
0C
#507310000000
1!
1*
b111 6
19
1>
1C
b111 G
#507320000000
0!
1"
0*
1+
09
1:
0>
0C
#507330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#507340000000
0!
0*
09
0>
0C
#507350000000
1!
1*
b1 6
19
1>
1C
b1 G
#507360000000
0!
0*
09
0>
0C
#507370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#507380000000
0!
0*
09
0>
0C
#507390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#507400000000
0!
0*
09
0>
0C
#507410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#507420000000
0!
0*
09
0>
0C
#507430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#507440000000
0!
0#
0*
0,
09
0>
0?
0C
#507450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#507460000000
0!
0*
09
0>
0C
#507470000000
1!
1*
19
1>
1C
#507480000000
0!
0*
09
0>
0C
#507490000000
1!
1*
19
1>
1C
#507500000000
0!
0*
09
0>
0C
#507510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#507520000000
0!
0*
09
0>
0C
#507530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#507540000000
0!
0*
09
0>
0C
#507550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#507560000000
0!
0*
09
0>
0C
#507570000000
1!
1*
b10 6
19
1>
1C
b10 G
#507580000000
0!
0*
09
0>
0C
#507590000000
1!
1*
b11 6
19
1>
1C
b11 G
#507600000000
0!
0*
09
0>
0C
#507610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#507620000000
0!
0*
09
0>
0C
#507630000000
1!
1*
b101 6
19
1>
1C
b101 G
#507640000000
0!
0*
09
0>
0C
#507650000000
1!
1*
b110 6
19
1>
1C
b110 G
#507660000000
0!
0*
09
0>
0C
#507670000000
1!
1*
b111 6
19
1>
1C
b111 G
#507680000000
0!
0*
09
0>
0C
#507690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#507700000000
0!
0*
09
0>
0C
#507710000000
1!
1*
b1 6
19
1>
1C
b1 G
#507720000000
0!
0*
09
0>
0C
#507730000000
1!
1*
b10 6
19
1>
1C
b10 G
#507740000000
0!
0*
09
0>
0C
#507750000000
1!
1*
b11 6
19
1>
1C
b11 G
#507760000000
0!
0*
09
0>
0C
#507770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#507780000000
0!
0*
09
0>
0C
#507790000000
1!
1*
b101 6
19
1>
1C
b101 G
#507800000000
0!
0*
09
0>
0C
#507810000000
1!
1*
b110 6
19
1>
1C
b110 G
#507820000000
0!
0*
09
0>
0C
#507830000000
1!
1*
b111 6
19
1>
1C
b111 G
#507840000000
0!
0*
09
0>
0C
#507850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#507860000000
0!
0*
09
0>
0C
#507870000000
1!
1*
b1 6
19
1>
1C
b1 G
#507880000000
0!
0*
09
0>
0C
#507890000000
1!
1*
b10 6
19
1>
1C
b10 G
#507900000000
0!
0*
09
0>
0C
#507910000000
1!
1*
b11 6
19
1>
1C
b11 G
#507920000000
0!
0*
09
0>
0C
#507930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#507940000000
0!
0*
09
0>
0C
#507950000000
1!
1*
b101 6
19
1>
1C
b101 G
#507960000000
0!
0*
09
0>
0C
#507970000000
1!
1*
b110 6
19
1>
1C
b110 G
#507980000000
0!
0*
09
0>
0C
#507990000000
1!
1*
b111 6
19
1>
1C
b111 G
#508000000000
0!
1"
0*
1+
09
1:
0>
0C
#508010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#508020000000
0!
0*
09
0>
0C
#508030000000
1!
1*
b1 6
19
1>
1C
b1 G
#508040000000
0!
0*
09
0>
0C
#508050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#508060000000
0!
0*
09
0>
0C
#508070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#508080000000
0!
0*
09
0>
0C
#508090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#508100000000
0!
0*
09
0>
0C
#508110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#508120000000
0!
0#
0*
0,
09
0>
0?
0C
#508130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#508140000000
0!
0*
09
0>
0C
#508150000000
1!
1*
19
1>
1C
#508160000000
0!
0*
09
0>
0C
#508170000000
1!
1*
19
1>
1C
#508180000000
0!
0*
09
0>
0C
#508190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#508200000000
0!
0*
09
0>
0C
#508210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#508220000000
0!
0*
09
0>
0C
#508230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#508240000000
0!
0*
09
0>
0C
#508250000000
1!
1*
b10 6
19
1>
1C
b10 G
#508260000000
0!
0*
09
0>
0C
#508270000000
1!
1*
b11 6
19
1>
1C
b11 G
#508280000000
0!
0*
09
0>
0C
#508290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#508300000000
0!
0*
09
0>
0C
#508310000000
1!
1*
b101 6
19
1>
1C
b101 G
#508320000000
0!
0*
09
0>
0C
#508330000000
1!
1*
b110 6
19
1>
1C
b110 G
#508340000000
0!
0*
09
0>
0C
#508350000000
1!
1*
b111 6
19
1>
1C
b111 G
#508360000000
0!
0*
09
0>
0C
#508370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#508380000000
0!
0*
09
0>
0C
#508390000000
1!
1*
b1 6
19
1>
1C
b1 G
#508400000000
0!
0*
09
0>
0C
#508410000000
1!
1*
b10 6
19
1>
1C
b10 G
#508420000000
0!
0*
09
0>
0C
#508430000000
1!
1*
b11 6
19
1>
1C
b11 G
#508440000000
0!
0*
09
0>
0C
#508450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#508460000000
0!
0*
09
0>
0C
#508470000000
1!
1*
b101 6
19
1>
1C
b101 G
#508480000000
0!
0*
09
0>
0C
#508490000000
1!
1*
b110 6
19
1>
1C
b110 G
#508500000000
0!
0*
09
0>
0C
#508510000000
1!
1*
b111 6
19
1>
1C
b111 G
#508520000000
0!
0*
09
0>
0C
#508530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#508540000000
0!
0*
09
0>
0C
#508550000000
1!
1*
b1 6
19
1>
1C
b1 G
#508560000000
0!
0*
09
0>
0C
#508570000000
1!
1*
b10 6
19
1>
1C
b10 G
#508580000000
0!
0*
09
0>
0C
#508590000000
1!
1*
b11 6
19
1>
1C
b11 G
#508600000000
0!
0*
09
0>
0C
#508610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#508620000000
0!
0*
09
0>
0C
#508630000000
1!
1*
b101 6
19
1>
1C
b101 G
#508640000000
0!
0*
09
0>
0C
#508650000000
1!
1*
b110 6
19
1>
1C
b110 G
#508660000000
0!
0*
09
0>
0C
#508670000000
1!
1*
b111 6
19
1>
1C
b111 G
#508680000000
0!
1"
0*
1+
09
1:
0>
0C
#508690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#508700000000
0!
0*
09
0>
0C
#508710000000
1!
1*
b1 6
19
1>
1C
b1 G
#508720000000
0!
0*
09
0>
0C
#508730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#508740000000
0!
0*
09
0>
0C
#508750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#508760000000
0!
0*
09
0>
0C
#508770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#508780000000
0!
0*
09
0>
0C
#508790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#508800000000
0!
0#
0*
0,
09
0>
0?
0C
#508810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#508820000000
0!
0*
09
0>
0C
#508830000000
1!
1*
19
1>
1C
#508840000000
0!
0*
09
0>
0C
#508850000000
1!
1*
19
1>
1C
#508860000000
0!
0*
09
0>
0C
#508870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#508880000000
0!
0*
09
0>
0C
#508890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#508900000000
0!
0*
09
0>
0C
#508910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#508920000000
0!
0*
09
0>
0C
#508930000000
1!
1*
b10 6
19
1>
1C
b10 G
#508940000000
0!
0*
09
0>
0C
#508950000000
1!
1*
b11 6
19
1>
1C
b11 G
#508960000000
0!
0*
09
0>
0C
#508970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#508980000000
0!
0*
09
0>
0C
#508990000000
1!
1*
b101 6
19
1>
1C
b101 G
#509000000000
0!
0*
09
0>
0C
#509010000000
1!
1*
b110 6
19
1>
1C
b110 G
#509020000000
0!
0*
09
0>
0C
#509030000000
1!
1*
b111 6
19
1>
1C
b111 G
#509040000000
0!
0*
09
0>
0C
#509050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#509060000000
0!
0*
09
0>
0C
#509070000000
1!
1*
b1 6
19
1>
1C
b1 G
#509080000000
0!
0*
09
0>
0C
#509090000000
1!
1*
b10 6
19
1>
1C
b10 G
#509100000000
0!
0*
09
0>
0C
#509110000000
1!
1*
b11 6
19
1>
1C
b11 G
#509120000000
0!
0*
09
0>
0C
#509130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#509140000000
0!
0*
09
0>
0C
#509150000000
1!
1*
b101 6
19
1>
1C
b101 G
#509160000000
0!
0*
09
0>
0C
#509170000000
1!
1*
b110 6
19
1>
1C
b110 G
#509180000000
0!
0*
09
0>
0C
#509190000000
1!
1*
b111 6
19
1>
1C
b111 G
#509200000000
0!
0*
09
0>
0C
#509210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#509220000000
0!
0*
09
0>
0C
#509230000000
1!
1*
b1 6
19
1>
1C
b1 G
#509240000000
0!
0*
09
0>
0C
#509250000000
1!
1*
b10 6
19
1>
1C
b10 G
#509260000000
0!
0*
09
0>
0C
#509270000000
1!
1*
b11 6
19
1>
1C
b11 G
#509280000000
0!
0*
09
0>
0C
#509290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#509300000000
0!
0*
09
0>
0C
#509310000000
1!
1*
b101 6
19
1>
1C
b101 G
#509320000000
0!
0*
09
0>
0C
#509330000000
1!
1*
b110 6
19
1>
1C
b110 G
#509340000000
0!
0*
09
0>
0C
#509350000000
1!
1*
b111 6
19
1>
1C
b111 G
#509360000000
0!
1"
0*
1+
09
1:
0>
0C
#509370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#509380000000
0!
0*
09
0>
0C
#509390000000
1!
1*
b1 6
19
1>
1C
b1 G
#509400000000
0!
0*
09
0>
0C
#509410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#509420000000
0!
0*
09
0>
0C
#509430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#509440000000
0!
0*
09
0>
0C
#509450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#509460000000
0!
0*
09
0>
0C
#509470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#509480000000
0!
0#
0*
0,
09
0>
0?
0C
#509490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#509500000000
0!
0*
09
0>
0C
#509510000000
1!
1*
19
1>
1C
#509520000000
0!
0*
09
0>
0C
#509530000000
1!
1*
19
1>
1C
#509540000000
0!
0*
09
0>
0C
#509550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#509560000000
0!
0*
09
0>
0C
#509570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#509580000000
0!
0*
09
0>
0C
#509590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#509600000000
0!
0*
09
0>
0C
#509610000000
1!
1*
b10 6
19
1>
1C
b10 G
#509620000000
0!
0*
09
0>
0C
#509630000000
1!
1*
b11 6
19
1>
1C
b11 G
#509640000000
0!
0*
09
0>
0C
#509650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#509660000000
0!
0*
09
0>
0C
#509670000000
1!
1*
b101 6
19
1>
1C
b101 G
#509680000000
0!
0*
09
0>
0C
#509690000000
1!
1*
b110 6
19
1>
1C
b110 G
#509700000000
0!
0*
09
0>
0C
#509710000000
1!
1*
b111 6
19
1>
1C
b111 G
#509720000000
0!
0*
09
0>
0C
#509730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#509740000000
0!
0*
09
0>
0C
#509750000000
1!
1*
b1 6
19
1>
1C
b1 G
#509760000000
0!
0*
09
0>
0C
#509770000000
1!
1*
b10 6
19
1>
1C
b10 G
#509780000000
0!
0*
09
0>
0C
#509790000000
1!
1*
b11 6
19
1>
1C
b11 G
#509800000000
0!
0*
09
0>
0C
#509810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#509820000000
0!
0*
09
0>
0C
#509830000000
1!
1*
b101 6
19
1>
1C
b101 G
#509840000000
0!
0*
09
0>
0C
#509850000000
1!
1*
b110 6
19
1>
1C
b110 G
#509860000000
0!
0*
09
0>
0C
#509870000000
1!
1*
b111 6
19
1>
1C
b111 G
#509880000000
0!
0*
09
0>
0C
#509890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#509900000000
0!
0*
09
0>
0C
#509910000000
1!
1*
b1 6
19
1>
1C
b1 G
#509920000000
0!
0*
09
0>
0C
#509930000000
1!
1*
b10 6
19
1>
1C
b10 G
#509940000000
0!
0*
09
0>
0C
#509950000000
1!
1*
b11 6
19
1>
1C
b11 G
#509960000000
0!
0*
09
0>
0C
#509970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#509980000000
0!
0*
09
0>
0C
#509990000000
1!
1*
b101 6
19
1>
1C
b101 G
#510000000000
0!
0*
09
0>
0C
#510010000000
1!
1*
b110 6
19
1>
1C
b110 G
#510020000000
0!
0*
09
0>
0C
#510030000000
1!
1*
b111 6
19
1>
1C
b111 G
#510040000000
0!
1"
0*
1+
09
1:
0>
0C
#510050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#510060000000
0!
0*
09
0>
0C
#510070000000
1!
1*
b1 6
19
1>
1C
b1 G
#510080000000
0!
0*
09
0>
0C
#510090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#510100000000
0!
0*
09
0>
0C
#510110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#510120000000
0!
0*
09
0>
0C
#510130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#510140000000
0!
0*
09
0>
0C
#510150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#510160000000
0!
0#
0*
0,
09
0>
0?
0C
#510170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#510180000000
0!
0*
09
0>
0C
#510190000000
1!
1*
19
1>
1C
#510200000000
0!
0*
09
0>
0C
#510210000000
1!
1*
19
1>
1C
#510220000000
0!
0*
09
0>
0C
#510230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#510240000000
0!
0*
09
0>
0C
#510250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#510260000000
0!
0*
09
0>
0C
#510270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#510280000000
0!
0*
09
0>
0C
#510290000000
1!
1*
b10 6
19
1>
1C
b10 G
#510300000000
0!
0*
09
0>
0C
#510310000000
1!
1*
b11 6
19
1>
1C
b11 G
#510320000000
0!
0*
09
0>
0C
#510330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#510340000000
0!
0*
09
0>
0C
#510350000000
1!
1*
b101 6
19
1>
1C
b101 G
#510360000000
0!
0*
09
0>
0C
#510370000000
1!
1*
b110 6
19
1>
1C
b110 G
#510380000000
0!
0*
09
0>
0C
#510390000000
1!
1*
b111 6
19
1>
1C
b111 G
#510400000000
0!
0*
09
0>
0C
#510410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#510420000000
0!
0*
09
0>
0C
#510430000000
1!
1*
b1 6
19
1>
1C
b1 G
#510440000000
0!
0*
09
0>
0C
#510450000000
1!
1*
b10 6
19
1>
1C
b10 G
#510460000000
0!
0*
09
0>
0C
#510470000000
1!
1*
b11 6
19
1>
1C
b11 G
#510480000000
0!
0*
09
0>
0C
#510490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#510500000000
0!
0*
09
0>
0C
#510510000000
1!
1*
b101 6
19
1>
1C
b101 G
#510520000000
0!
0*
09
0>
0C
#510530000000
1!
1*
b110 6
19
1>
1C
b110 G
#510540000000
0!
0*
09
0>
0C
#510550000000
1!
1*
b111 6
19
1>
1C
b111 G
#510560000000
0!
0*
09
0>
0C
#510570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#510580000000
0!
0*
09
0>
0C
#510590000000
1!
1*
b1 6
19
1>
1C
b1 G
#510600000000
0!
0*
09
0>
0C
#510610000000
1!
1*
b10 6
19
1>
1C
b10 G
#510620000000
0!
0*
09
0>
0C
#510630000000
1!
1*
b11 6
19
1>
1C
b11 G
#510640000000
0!
0*
09
0>
0C
#510650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#510660000000
0!
0*
09
0>
0C
#510670000000
1!
1*
b101 6
19
1>
1C
b101 G
#510680000000
0!
0*
09
0>
0C
#510690000000
1!
1*
b110 6
19
1>
1C
b110 G
#510700000000
0!
0*
09
0>
0C
#510710000000
1!
1*
b111 6
19
1>
1C
b111 G
#510720000000
0!
1"
0*
1+
09
1:
0>
0C
#510730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#510740000000
0!
0*
09
0>
0C
#510750000000
1!
1*
b1 6
19
1>
1C
b1 G
#510760000000
0!
0*
09
0>
0C
#510770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#510780000000
0!
0*
09
0>
0C
#510790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#510800000000
0!
0*
09
0>
0C
#510810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#510820000000
0!
0*
09
0>
0C
#510830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#510840000000
0!
0#
0*
0,
09
0>
0?
0C
#510850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#510860000000
0!
0*
09
0>
0C
#510870000000
1!
1*
19
1>
1C
#510880000000
0!
0*
09
0>
0C
#510890000000
1!
1*
19
1>
1C
#510900000000
0!
0*
09
0>
0C
#510910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#510920000000
0!
0*
09
0>
0C
#510930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#510940000000
0!
0*
09
0>
0C
#510950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#510960000000
0!
0*
09
0>
0C
#510970000000
1!
1*
b10 6
19
1>
1C
b10 G
#510980000000
0!
0*
09
0>
0C
#510990000000
1!
1*
b11 6
19
1>
1C
b11 G
#511000000000
0!
0*
09
0>
0C
#511010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#511020000000
0!
0*
09
0>
0C
#511030000000
1!
1*
b101 6
19
1>
1C
b101 G
#511040000000
0!
0*
09
0>
0C
#511050000000
1!
1*
b110 6
19
1>
1C
b110 G
#511060000000
0!
0*
09
0>
0C
#511070000000
1!
1*
b111 6
19
1>
1C
b111 G
#511080000000
0!
0*
09
0>
0C
#511090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#511100000000
0!
0*
09
0>
0C
#511110000000
1!
1*
b1 6
19
1>
1C
b1 G
#511120000000
0!
0*
09
0>
0C
#511130000000
1!
1*
b10 6
19
1>
1C
b10 G
#511140000000
0!
0*
09
0>
0C
#511150000000
1!
1*
b11 6
19
1>
1C
b11 G
#511160000000
0!
0*
09
0>
0C
#511170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#511180000000
0!
0*
09
0>
0C
#511190000000
1!
1*
b101 6
19
1>
1C
b101 G
#511200000000
0!
0*
09
0>
0C
#511210000000
1!
1*
b110 6
19
1>
1C
b110 G
#511220000000
0!
0*
09
0>
0C
#511230000000
1!
1*
b111 6
19
1>
1C
b111 G
#511240000000
0!
0*
09
0>
0C
#511250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#511260000000
0!
0*
09
0>
0C
#511270000000
1!
1*
b1 6
19
1>
1C
b1 G
#511280000000
0!
0*
09
0>
0C
#511290000000
1!
1*
b10 6
19
1>
1C
b10 G
#511300000000
0!
0*
09
0>
0C
#511310000000
1!
1*
b11 6
19
1>
1C
b11 G
#511320000000
0!
0*
09
0>
0C
#511330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#511340000000
0!
0*
09
0>
0C
#511350000000
1!
1*
b101 6
19
1>
1C
b101 G
#511360000000
0!
0*
09
0>
0C
#511370000000
1!
1*
b110 6
19
1>
1C
b110 G
#511380000000
0!
0*
09
0>
0C
#511390000000
1!
1*
b111 6
19
1>
1C
b111 G
#511400000000
0!
1"
0*
1+
09
1:
0>
0C
#511410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#511420000000
0!
0*
09
0>
0C
#511430000000
1!
1*
b1 6
19
1>
1C
b1 G
#511440000000
0!
0*
09
0>
0C
#511450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#511460000000
0!
0*
09
0>
0C
#511470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#511480000000
0!
0*
09
0>
0C
#511490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#511500000000
0!
0*
09
0>
0C
#511510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#511520000000
0!
0#
0*
0,
09
0>
0?
0C
#511530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#511540000000
0!
0*
09
0>
0C
#511550000000
1!
1*
19
1>
1C
#511560000000
0!
0*
09
0>
0C
#511570000000
1!
1*
19
1>
1C
#511580000000
0!
0*
09
0>
0C
#511590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#511600000000
0!
0*
09
0>
0C
#511610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#511620000000
0!
0*
09
0>
0C
#511630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#511640000000
0!
0*
09
0>
0C
#511650000000
1!
1*
b10 6
19
1>
1C
b10 G
#511660000000
0!
0*
09
0>
0C
#511670000000
1!
1*
b11 6
19
1>
1C
b11 G
#511680000000
0!
0*
09
0>
0C
#511690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#511700000000
0!
0*
09
0>
0C
#511710000000
1!
1*
b101 6
19
1>
1C
b101 G
#511720000000
0!
0*
09
0>
0C
#511730000000
1!
1*
b110 6
19
1>
1C
b110 G
#511740000000
0!
0*
09
0>
0C
#511750000000
1!
1*
b111 6
19
1>
1C
b111 G
#511760000000
0!
0*
09
0>
0C
#511770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#511780000000
0!
0*
09
0>
0C
#511790000000
1!
1*
b1 6
19
1>
1C
b1 G
#511800000000
0!
0*
09
0>
0C
#511810000000
1!
1*
b10 6
19
1>
1C
b10 G
#511820000000
0!
0*
09
0>
0C
#511830000000
1!
1*
b11 6
19
1>
1C
b11 G
#511840000000
0!
0*
09
0>
0C
#511850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#511860000000
0!
0*
09
0>
0C
#511870000000
1!
1*
b101 6
19
1>
1C
b101 G
#511880000000
0!
0*
09
0>
0C
#511890000000
1!
1*
b110 6
19
1>
1C
b110 G
#511900000000
0!
0*
09
0>
0C
#511910000000
1!
1*
b111 6
19
1>
1C
b111 G
#511920000000
0!
0*
09
0>
0C
#511930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#511940000000
0!
0*
09
0>
0C
#511950000000
1!
1*
b1 6
19
1>
1C
b1 G
#511960000000
0!
0*
09
0>
0C
#511970000000
1!
1*
b10 6
19
1>
1C
b10 G
#511980000000
0!
0*
09
0>
0C
#511990000000
1!
1*
b11 6
19
1>
1C
b11 G
#512000000000
0!
0*
09
0>
0C
#512010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#512020000000
0!
0*
09
0>
0C
#512030000000
1!
1*
b101 6
19
1>
1C
b101 G
#512040000000
0!
0*
09
0>
0C
#512050000000
1!
1*
b110 6
19
1>
1C
b110 G
#512060000000
0!
0*
09
0>
0C
#512070000000
1!
1*
b111 6
19
1>
1C
b111 G
#512080000000
0!
1"
0*
1+
09
1:
0>
0C
#512090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#512100000000
0!
0*
09
0>
0C
#512110000000
1!
1*
b1 6
19
1>
1C
b1 G
#512120000000
0!
0*
09
0>
0C
#512130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#512140000000
0!
0*
09
0>
0C
#512150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#512160000000
0!
0*
09
0>
0C
#512170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#512180000000
0!
0*
09
0>
0C
#512190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#512200000000
0!
0#
0*
0,
09
0>
0?
0C
#512210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#512220000000
0!
0*
09
0>
0C
#512230000000
1!
1*
19
1>
1C
#512240000000
0!
0*
09
0>
0C
#512250000000
1!
1*
19
1>
1C
#512260000000
0!
0*
09
0>
0C
#512270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#512280000000
0!
0*
09
0>
0C
#512290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#512300000000
0!
0*
09
0>
0C
#512310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#512320000000
0!
0*
09
0>
0C
#512330000000
1!
1*
b10 6
19
1>
1C
b10 G
#512340000000
0!
0*
09
0>
0C
#512350000000
1!
1*
b11 6
19
1>
1C
b11 G
#512360000000
0!
0*
09
0>
0C
#512370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#512380000000
0!
0*
09
0>
0C
#512390000000
1!
1*
b101 6
19
1>
1C
b101 G
#512400000000
0!
0*
09
0>
0C
#512410000000
1!
1*
b110 6
19
1>
1C
b110 G
#512420000000
0!
0*
09
0>
0C
#512430000000
1!
1*
b111 6
19
1>
1C
b111 G
#512440000000
0!
0*
09
0>
0C
#512450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#512460000000
0!
0*
09
0>
0C
#512470000000
1!
1*
b1 6
19
1>
1C
b1 G
#512480000000
0!
0*
09
0>
0C
#512490000000
1!
1*
b10 6
19
1>
1C
b10 G
#512500000000
0!
0*
09
0>
0C
#512510000000
1!
1*
b11 6
19
1>
1C
b11 G
#512520000000
0!
0*
09
0>
0C
#512530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#512540000000
0!
0*
09
0>
0C
#512550000000
1!
1*
b101 6
19
1>
1C
b101 G
#512560000000
0!
0*
09
0>
0C
#512570000000
1!
1*
b110 6
19
1>
1C
b110 G
#512580000000
0!
0*
09
0>
0C
#512590000000
1!
1*
b111 6
19
1>
1C
b111 G
#512600000000
0!
0*
09
0>
0C
#512610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#512620000000
0!
0*
09
0>
0C
#512630000000
1!
1*
b1 6
19
1>
1C
b1 G
#512640000000
0!
0*
09
0>
0C
#512650000000
1!
1*
b10 6
19
1>
1C
b10 G
#512660000000
0!
0*
09
0>
0C
#512670000000
1!
1*
b11 6
19
1>
1C
b11 G
#512680000000
0!
0*
09
0>
0C
#512690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#512700000000
0!
0*
09
0>
0C
#512710000000
1!
1*
b101 6
19
1>
1C
b101 G
#512720000000
0!
0*
09
0>
0C
#512730000000
1!
1*
b110 6
19
1>
1C
b110 G
#512740000000
0!
0*
09
0>
0C
#512750000000
1!
1*
b111 6
19
1>
1C
b111 G
#512760000000
0!
1"
0*
1+
09
1:
0>
0C
#512770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#512780000000
0!
0*
09
0>
0C
#512790000000
1!
1*
b1 6
19
1>
1C
b1 G
#512800000000
0!
0*
09
0>
0C
#512810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#512820000000
0!
0*
09
0>
0C
#512830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#512840000000
0!
0*
09
0>
0C
#512850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#512860000000
0!
0*
09
0>
0C
#512870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#512880000000
0!
0#
0*
0,
09
0>
0?
0C
#512890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#512900000000
0!
0*
09
0>
0C
#512910000000
1!
1*
19
1>
1C
#512920000000
0!
0*
09
0>
0C
#512930000000
1!
1*
19
1>
1C
#512940000000
0!
0*
09
0>
0C
#512950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#512960000000
0!
0*
09
0>
0C
#512970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#512980000000
0!
0*
09
0>
0C
#512990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#513000000000
0!
0*
09
0>
0C
#513010000000
1!
1*
b10 6
19
1>
1C
b10 G
#513020000000
0!
0*
09
0>
0C
#513030000000
1!
1*
b11 6
19
1>
1C
b11 G
#513040000000
0!
0*
09
0>
0C
#513050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#513060000000
0!
0*
09
0>
0C
#513070000000
1!
1*
b101 6
19
1>
1C
b101 G
#513080000000
0!
0*
09
0>
0C
#513090000000
1!
1*
b110 6
19
1>
1C
b110 G
#513100000000
0!
0*
09
0>
0C
#513110000000
1!
1*
b111 6
19
1>
1C
b111 G
#513120000000
0!
0*
09
0>
0C
#513130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#513140000000
0!
0*
09
0>
0C
#513150000000
1!
1*
b1 6
19
1>
1C
b1 G
#513160000000
0!
0*
09
0>
0C
#513170000000
1!
1*
b10 6
19
1>
1C
b10 G
#513180000000
0!
0*
09
0>
0C
#513190000000
1!
1*
b11 6
19
1>
1C
b11 G
#513200000000
0!
0*
09
0>
0C
#513210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#513220000000
0!
0*
09
0>
0C
#513230000000
1!
1*
b101 6
19
1>
1C
b101 G
#513240000000
0!
0*
09
0>
0C
#513250000000
1!
1*
b110 6
19
1>
1C
b110 G
#513260000000
0!
0*
09
0>
0C
#513270000000
1!
1*
b111 6
19
1>
1C
b111 G
#513280000000
0!
0*
09
0>
0C
#513290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#513300000000
0!
0*
09
0>
0C
#513310000000
1!
1*
b1 6
19
1>
1C
b1 G
#513320000000
0!
0*
09
0>
0C
#513330000000
1!
1*
b10 6
19
1>
1C
b10 G
#513340000000
0!
0*
09
0>
0C
#513350000000
1!
1*
b11 6
19
1>
1C
b11 G
#513360000000
0!
0*
09
0>
0C
#513370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#513380000000
0!
0*
09
0>
0C
#513390000000
1!
1*
b101 6
19
1>
1C
b101 G
#513400000000
0!
0*
09
0>
0C
#513410000000
1!
1*
b110 6
19
1>
1C
b110 G
#513420000000
0!
0*
09
0>
0C
#513430000000
1!
1*
b111 6
19
1>
1C
b111 G
#513440000000
0!
1"
0*
1+
09
1:
0>
0C
#513450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#513460000000
0!
0*
09
0>
0C
#513470000000
1!
1*
b1 6
19
1>
1C
b1 G
#513480000000
0!
0*
09
0>
0C
#513490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#513500000000
0!
0*
09
0>
0C
#513510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#513520000000
0!
0*
09
0>
0C
#513530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#513540000000
0!
0*
09
0>
0C
#513550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#513560000000
0!
0#
0*
0,
09
0>
0?
0C
#513570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#513580000000
0!
0*
09
0>
0C
#513590000000
1!
1*
19
1>
1C
#513600000000
0!
0*
09
0>
0C
#513610000000
1!
1*
19
1>
1C
#513620000000
0!
0*
09
0>
0C
#513630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#513640000000
0!
0*
09
0>
0C
#513650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#513660000000
0!
0*
09
0>
0C
#513670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#513680000000
0!
0*
09
0>
0C
#513690000000
1!
1*
b10 6
19
1>
1C
b10 G
#513700000000
0!
0*
09
0>
0C
#513710000000
1!
1*
b11 6
19
1>
1C
b11 G
#513720000000
0!
0*
09
0>
0C
#513730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#513740000000
0!
0*
09
0>
0C
#513750000000
1!
1*
b101 6
19
1>
1C
b101 G
#513760000000
0!
0*
09
0>
0C
#513770000000
1!
1*
b110 6
19
1>
1C
b110 G
#513780000000
0!
0*
09
0>
0C
#513790000000
1!
1*
b111 6
19
1>
1C
b111 G
#513800000000
0!
0*
09
0>
0C
#513810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#513820000000
0!
0*
09
0>
0C
#513830000000
1!
1*
b1 6
19
1>
1C
b1 G
#513840000000
0!
0*
09
0>
0C
#513850000000
1!
1*
b10 6
19
1>
1C
b10 G
#513860000000
0!
0*
09
0>
0C
#513870000000
1!
1*
b11 6
19
1>
1C
b11 G
#513880000000
0!
0*
09
0>
0C
#513890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#513900000000
0!
0*
09
0>
0C
#513910000000
1!
1*
b101 6
19
1>
1C
b101 G
#513920000000
0!
0*
09
0>
0C
#513930000000
1!
1*
b110 6
19
1>
1C
b110 G
#513940000000
0!
0*
09
0>
0C
#513950000000
1!
1*
b111 6
19
1>
1C
b111 G
#513960000000
0!
0*
09
0>
0C
#513970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#513980000000
0!
0*
09
0>
0C
#513990000000
1!
1*
b1 6
19
1>
1C
b1 G
#514000000000
0!
0*
09
0>
0C
#514010000000
1!
1*
b10 6
19
1>
1C
b10 G
#514020000000
0!
0*
09
0>
0C
#514030000000
1!
1*
b11 6
19
1>
1C
b11 G
#514040000000
0!
0*
09
0>
0C
#514050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#514060000000
0!
0*
09
0>
0C
#514070000000
1!
1*
b101 6
19
1>
1C
b101 G
#514080000000
0!
0*
09
0>
0C
#514090000000
1!
1*
b110 6
19
1>
1C
b110 G
#514100000000
0!
0*
09
0>
0C
#514110000000
1!
1*
b111 6
19
1>
1C
b111 G
#514120000000
0!
1"
0*
1+
09
1:
0>
0C
#514130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#514140000000
0!
0*
09
0>
0C
#514150000000
1!
1*
b1 6
19
1>
1C
b1 G
#514160000000
0!
0*
09
0>
0C
#514170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#514180000000
0!
0*
09
0>
0C
#514190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#514200000000
0!
0*
09
0>
0C
#514210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#514220000000
0!
0*
09
0>
0C
#514230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#514240000000
0!
0#
0*
0,
09
0>
0?
0C
#514250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#514260000000
0!
0*
09
0>
0C
#514270000000
1!
1*
19
1>
1C
#514280000000
0!
0*
09
0>
0C
#514290000000
1!
1*
19
1>
1C
#514300000000
0!
0*
09
0>
0C
#514310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#514320000000
0!
0*
09
0>
0C
#514330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#514340000000
0!
0*
09
0>
0C
#514350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#514360000000
0!
0*
09
0>
0C
#514370000000
1!
1*
b10 6
19
1>
1C
b10 G
#514380000000
0!
0*
09
0>
0C
#514390000000
1!
1*
b11 6
19
1>
1C
b11 G
#514400000000
0!
0*
09
0>
0C
#514410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#514420000000
0!
0*
09
0>
0C
#514430000000
1!
1*
b101 6
19
1>
1C
b101 G
#514440000000
0!
0*
09
0>
0C
#514450000000
1!
1*
b110 6
19
1>
1C
b110 G
#514460000000
0!
0*
09
0>
0C
#514470000000
1!
1*
b111 6
19
1>
1C
b111 G
#514480000000
0!
0*
09
0>
0C
#514490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#514500000000
0!
0*
09
0>
0C
#514510000000
1!
1*
b1 6
19
1>
1C
b1 G
#514520000000
0!
0*
09
0>
0C
#514530000000
1!
1*
b10 6
19
1>
1C
b10 G
#514540000000
0!
0*
09
0>
0C
#514550000000
1!
1*
b11 6
19
1>
1C
b11 G
#514560000000
0!
0*
09
0>
0C
#514570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#514580000000
0!
0*
09
0>
0C
#514590000000
1!
1*
b101 6
19
1>
1C
b101 G
#514600000000
0!
0*
09
0>
0C
#514610000000
1!
1*
b110 6
19
1>
1C
b110 G
#514620000000
0!
0*
09
0>
0C
#514630000000
1!
1*
b111 6
19
1>
1C
b111 G
#514640000000
0!
0*
09
0>
0C
#514650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#514660000000
0!
0*
09
0>
0C
#514670000000
1!
1*
b1 6
19
1>
1C
b1 G
#514680000000
0!
0*
09
0>
0C
#514690000000
1!
1*
b10 6
19
1>
1C
b10 G
#514700000000
0!
0*
09
0>
0C
#514710000000
1!
1*
b11 6
19
1>
1C
b11 G
#514720000000
0!
0*
09
0>
0C
#514730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#514740000000
0!
0*
09
0>
0C
#514750000000
1!
1*
b101 6
19
1>
1C
b101 G
#514760000000
0!
0*
09
0>
0C
#514770000000
1!
1*
b110 6
19
1>
1C
b110 G
#514780000000
0!
0*
09
0>
0C
#514790000000
1!
1*
b111 6
19
1>
1C
b111 G
#514800000000
0!
1"
0*
1+
09
1:
0>
0C
#514810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#514820000000
0!
0*
09
0>
0C
#514830000000
1!
1*
b1 6
19
1>
1C
b1 G
#514840000000
0!
0*
09
0>
0C
#514850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#514860000000
0!
0*
09
0>
0C
#514870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#514880000000
0!
0*
09
0>
0C
#514890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#514900000000
0!
0*
09
0>
0C
#514910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#514920000000
0!
0#
0*
0,
09
0>
0?
0C
#514930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#514940000000
0!
0*
09
0>
0C
#514950000000
1!
1*
19
1>
1C
#514960000000
0!
0*
09
0>
0C
#514970000000
1!
1*
19
1>
1C
#514980000000
0!
0*
09
0>
0C
#514990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#515000000000
0!
0*
09
0>
0C
#515010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#515020000000
0!
0*
09
0>
0C
#515030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#515040000000
0!
0*
09
0>
0C
#515050000000
1!
1*
b10 6
19
1>
1C
b10 G
#515060000000
0!
0*
09
0>
0C
#515070000000
1!
1*
b11 6
19
1>
1C
b11 G
#515080000000
0!
0*
09
0>
0C
#515090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#515100000000
0!
0*
09
0>
0C
#515110000000
1!
1*
b101 6
19
1>
1C
b101 G
#515120000000
0!
0*
09
0>
0C
#515130000000
1!
1*
b110 6
19
1>
1C
b110 G
#515140000000
0!
0*
09
0>
0C
#515150000000
1!
1*
b111 6
19
1>
1C
b111 G
#515160000000
0!
0*
09
0>
0C
#515170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#515180000000
0!
0*
09
0>
0C
#515190000000
1!
1*
b1 6
19
1>
1C
b1 G
#515200000000
0!
0*
09
0>
0C
#515210000000
1!
1*
b10 6
19
1>
1C
b10 G
#515220000000
0!
0*
09
0>
0C
#515230000000
1!
1*
b11 6
19
1>
1C
b11 G
#515240000000
0!
0*
09
0>
0C
#515250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#515260000000
0!
0*
09
0>
0C
#515270000000
1!
1*
b101 6
19
1>
1C
b101 G
#515280000000
0!
0*
09
0>
0C
#515290000000
1!
1*
b110 6
19
1>
1C
b110 G
#515300000000
0!
0*
09
0>
0C
#515310000000
1!
1*
b111 6
19
1>
1C
b111 G
#515320000000
0!
0*
09
0>
0C
#515330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#515340000000
0!
0*
09
0>
0C
#515350000000
1!
1*
b1 6
19
1>
1C
b1 G
#515360000000
0!
0*
09
0>
0C
#515370000000
1!
1*
b10 6
19
1>
1C
b10 G
#515380000000
0!
0*
09
0>
0C
#515390000000
1!
1*
b11 6
19
1>
1C
b11 G
#515400000000
0!
0*
09
0>
0C
#515410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#515420000000
0!
0*
09
0>
0C
#515430000000
1!
1*
b101 6
19
1>
1C
b101 G
#515440000000
0!
0*
09
0>
0C
#515450000000
1!
1*
b110 6
19
1>
1C
b110 G
#515460000000
0!
0*
09
0>
0C
#515470000000
1!
1*
b111 6
19
1>
1C
b111 G
#515480000000
0!
1"
0*
1+
09
1:
0>
0C
#515490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#515500000000
0!
0*
09
0>
0C
#515510000000
1!
1*
b1 6
19
1>
1C
b1 G
#515520000000
0!
0*
09
0>
0C
#515530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#515540000000
0!
0*
09
0>
0C
#515550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#515560000000
0!
0*
09
0>
0C
#515570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#515580000000
0!
0*
09
0>
0C
#515590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#515600000000
0!
0#
0*
0,
09
0>
0?
0C
#515610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#515620000000
0!
0*
09
0>
0C
#515630000000
1!
1*
19
1>
1C
#515640000000
0!
0*
09
0>
0C
#515650000000
1!
1*
19
1>
1C
#515660000000
0!
0*
09
0>
0C
#515670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#515680000000
0!
0*
09
0>
0C
#515690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#515700000000
0!
0*
09
0>
0C
#515710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#515720000000
0!
0*
09
0>
0C
#515730000000
1!
1*
b10 6
19
1>
1C
b10 G
#515740000000
0!
0*
09
0>
0C
#515750000000
1!
1*
b11 6
19
1>
1C
b11 G
#515760000000
0!
0*
09
0>
0C
#515770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#515780000000
0!
0*
09
0>
0C
#515790000000
1!
1*
b101 6
19
1>
1C
b101 G
#515800000000
0!
0*
09
0>
0C
#515810000000
1!
1*
b110 6
19
1>
1C
b110 G
#515820000000
0!
0*
09
0>
0C
#515830000000
1!
1*
b111 6
19
1>
1C
b111 G
#515840000000
0!
0*
09
0>
0C
#515850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#515860000000
0!
0*
09
0>
0C
#515870000000
1!
1*
b1 6
19
1>
1C
b1 G
#515880000000
0!
0*
09
0>
0C
#515890000000
1!
1*
b10 6
19
1>
1C
b10 G
#515900000000
0!
0*
09
0>
0C
#515910000000
1!
1*
b11 6
19
1>
1C
b11 G
#515920000000
0!
0*
09
0>
0C
#515930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#515940000000
0!
0*
09
0>
0C
#515950000000
1!
1*
b101 6
19
1>
1C
b101 G
#515960000000
0!
0*
09
0>
0C
#515970000000
1!
1*
b110 6
19
1>
1C
b110 G
#515980000000
0!
0*
09
0>
0C
#515990000000
1!
1*
b111 6
19
1>
1C
b111 G
#516000000000
0!
0*
09
0>
0C
#516010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#516020000000
0!
0*
09
0>
0C
#516030000000
1!
1*
b1 6
19
1>
1C
b1 G
#516040000000
0!
0*
09
0>
0C
#516050000000
1!
1*
b10 6
19
1>
1C
b10 G
#516060000000
0!
0*
09
0>
0C
#516070000000
1!
1*
b11 6
19
1>
1C
b11 G
#516080000000
0!
0*
09
0>
0C
#516090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#516100000000
0!
0*
09
0>
0C
#516110000000
1!
1*
b101 6
19
1>
1C
b101 G
#516120000000
0!
0*
09
0>
0C
#516130000000
1!
1*
b110 6
19
1>
1C
b110 G
#516140000000
0!
0*
09
0>
0C
#516150000000
1!
1*
b111 6
19
1>
1C
b111 G
#516160000000
0!
1"
0*
1+
09
1:
0>
0C
#516170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#516180000000
0!
0*
09
0>
0C
#516190000000
1!
1*
b1 6
19
1>
1C
b1 G
#516200000000
0!
0*
09
0>
0C
#516210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#516220000000
0!
0*
09
0>
0C
#516230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#516240000000
0!
0*
09
0>
0C
#516250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#516260000000
0!
0*
09
0>
0C
#516270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#516280000000
0!
0#
0*
0,
09
0>
0?
0C
#516290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#516300000000
0!
0*
09
0>
0C
#516310000000
1!
1*
19
1>
1C
#516320000000
0!
0*
09
0>
0C
#516330000000
1!
1*
19
1>
1C
#516340000000
0!
0*
09
0>
0C
#516350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#516360000000
0!
0*
09
0>
0C
#516370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#516380000000
0!
0*
09
0>
0C
#516390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#516400000000
0!
0*
09
0>
0C
#516410000000
1!
1*
b10 6
19
1>
1C
b10 G
#516420000000
0!
0*
09
0>
0C
#516430000000
1!
1*
b11 6
19
1>
1C
b11 G
#516440000000
0!
0*
09
0>
0C
#516450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#516460000000
0!
0*
09
0>
0C
#516470000000
1!
1*
b101 6
19
1>
1C
b101 G
#516480000000
0!
0*
09
0>
0C
#516490000000
1!
1*
b110 6
19
1>
1C
b110 G
#516500000000
0!
0*
09
0>
0C
#516510000000
1!
1*
b111 6
19
1>
1C
b111 G
#516520000000
0!
0*
09
0>
0C
#516530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#516540000000
0!
0*
09
0>
0C
#516550000000
1!
1*
b1 6
19
1>
1C
b1 G
#516560000000
0!
0*
09
0>
0C
#516570000000
1!
1*
b10 6
19
1>
1C
b10 G
#516580000000
0!
0*
09
0>
0C
#516590000000
1!
1*
b11 6
19
1>
1C
b11 G
#516600000000
0!
0*
09
0>
0C
#516610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#516620000000
0!
0*
09
0>
0C
#516630000000
1!
1*
b101 6
19
1>
1C
b101 G
#516640000000
0!
0*
09
0>
0C
#516650000000
1!
1*
b110 6
19
1>
1C
b110 G
#516660000000
0!
0*
09
0>
0C
#516670000000
1!
1*
b111 6
19
1>
1C
b111 G
#516680000000
0!
0*
09
0>
0C
#516690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#516700000000
0!
0*
09
0>
0C
#516710000000
1!
1*
b1 6
19
1>
1C
b1 G
#516720000000
0!
0*
09
0>
0C
#516730000000
1!
1*
b10 6
19
1>
1C
b10 G
#516740000000
0!
0*
09
0>
0C
#516750000000
1!
1*
b11 6
19
1>
1C
b11 G
#516760000000
0!
0*
09
0>
0C
#516770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#516780000000
0!
0*
09
0>
0C
#516790000000
1!
1*
b101 6
19
1>
1C
b101 G
#516800000000
0!
0*
09
0>
0C
#516810000000
1!
1*
b110 6
19
1>
1C
b110 G
#516820000000
0!
0*
09
0>
0C
#516830000000
1!
1*
b111 6
19
1>
1C
b111 G
#516840000000
0!
1"
0*
1+
09
1:
0>
0C
#516850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#516860000000
0!
0*
09
0>
0C
#516870000000
1!
1*
b1 6
19
1>
1C
b1 G
#516880000000
0!
0*
09
0>
0C
#516890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#516900000000
0!
0*
09
0>
0C
#516910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#516920000000
0!
0*
09
0>
0C
#516930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#516940000000
0!
0*
09
0>
0C
#516950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#516960000000
0!
0#
0*
0,
09
0>
0?
0C
#516970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#516980000000
0!
0*
09
0>
0C
#516990000000
1!
1*
19
1>
1C
#517000000000
0!
0*
09
0>
0C
#517010000000
1!
1*
19
1>
1C
#517020000000
0!
0*
09
0>
0C
#517030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#517040000000
0!
0*
09
0>
0C
#517050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#517060000000
0!
0*
09
0>
0C
#517070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#517080000000
0!
0*
09
0>
0C
#517090000000
1!
1*
b10 6
19
1>
1C
b10 G
#517100000000
0!
0*
09
0>
0C
#517110000000
1!
1*
b11 6
19
1>
1C
b11 G
#517120000000
0!
0*
09
0>
0C
#517130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#517140000000
0!
0*
09
0>
0C
#517150000000
1!
1*
b101 6
19
1>
1C
b101 G
#517160000000
0!
0*
09
0>
0C
#517170000000
1!
1*
b110 6
19
1>
1C
b110 G
#517180000000
0!
0*
09
0>
0C
#517190000000
1!
1*
b111 6
19
1>
1C
b111 G
#517200000000
0!
0*
09
0>
0C
#517210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#517220000000
0!
0*
09
0>
0C
#517230000000
1!
1*
b1 6
19
1>
1C
b1 G
#517240000000
0!
0*
09
0>
0C
#517250000000
1!
1*
b10 6
19
1>
1C
b10 G
#517260000000
0!
0*
09
0>
0C
#517270000000
1!
1*
b11 6
19
1>
1C
b11 G
#517280000000
0!
0*
09
0>
0C
#517290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#517300000000
0!
0*
09
0>
0C
#517310000000
1!
1*
b101 6
19
1>
1C
b101 G
#517320000000
0!
0*
09
0>
0C
#517330000000
1!
1*
b110 6
19
1>
1C
b110 G
#517340000000
0!
0*
09
0>
0C
#517350000000
1!
1*
b111 6
19
1>
1C
b111 G
#517360000000
0!
0*
09
0>
0C
#517370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#517380000000
0!
0*
09
0>
0C
#517390000000
1!
1*
b1 6
19
1>
1C
b1 G
#517400000000
0!
0*
09
0>
0C
#517410000000
1!
1*
b10 6
19
1>
1C
b10 G
#517420000000
0!
0*
09
0>
0C
#517430000000
1!
1*
b11 6
19
1>
1C
b11 G
#517440000000
0!
0*
09
0>
0C
#517450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#517460000000
0!
0*
09
0>
0C
#517470000000
1!
1*
b101 6
19
1>
1C
b101 G
#517480000000
0!
0*
09
0>
0C
#517490000000
1!
1*
b110 6
19
1>
1C
b110 G
#517500000000
0!
0*
09
0>
0C
#517510000000
1!
1*
b111 6
19
1>
1C
b111 G
#517520000000
0!
1"
0*
1+
09
1:
0>
0C
#517530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#517540000000
0!
0*
09
0>
0C
#517550000000
1!
1*
b1 6
19
1>
1C
b1 G
#517560000000
0!
0*
09
0>
0C
#517570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#517580000000
0!
0*
09
0>
0C
#517590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#517600000000
0!
0*
09
0>
0C
#517610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#517620000000
0!
0*
09
0>
0C
#517630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#517640000000
0!
0#
0*
0,
09
0>
0?
0C
#517650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#517660000000
0!
0*
09
0>
0C
#517670000000
1!
1*
19
1>
1C
#517680000000
0!
0*
09
0>
0C
#517690000000
1!
1*
19
1>
1C
#517700000000
0!
0*
09
0>
0C
#517710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#517720000000
0!
0*
09
0>
0C
#517730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#517740000000
0!
0*
09
0>
0C
#517750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#517760000000
0!
0*
09
0>
0C
#517770000000
1!
1*
b10 6
19
1>
1C
b10 G
#517780000000
0!
0*
09
0>
0C
#517790000000
1!
1*
b11 6
19
1>
1C
b11 G
#517800000000
0!
0*
09
0>
0C
#517810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#517820000000
0!
0*
09
0>
0C
#517830000000
1!
1*
b101 6
19
1>
1C
b101 G
#517840000000
0!
0*
09
0>
0C
#517850000000
1!
1*
b110 6
19
1>
1C
b110 G
#517860000000
0!
0*
09
0>
0C
#517870000000
1!
1*
b111 6
19
1>
1C
b111 G
#517880000000
0!
0*
09
0>
0C
#517890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#517900000000
0!
0*
09
0>
0C
#517910000000
1!
1*
b1 6
19
1>
1C
b1 G
#517920000000
0!
0*
09
0>
0C
#517930000000
1!
1*
b10 6
19
1>
1C
b10 G
#517940000000
0!
0*
09
0>
0C
#517950000000
1!
1*
b11 6
19
1>
1C
b11 G
#517960000000
0!
0*
09
0>
0C
#517970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#517980000000
0!
0*
09
0>
0C
#517990000000
1!
1*
b101 6
19
1>
1C
b101 G
#518000000000
0!
0*
09
0>
0C
#518010000000
1!
1*
b110 6
19
1>
1C
b110 G
#518020000000
0!
0*
09
0>
0C
#518030000000
1!
1*
b111 6
19
1>
1C
b111 G
#518040000000
0!
0*
09
0>
0C
#518050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#518060000000
0!
0*
09
0>
0C
#518070000000
1!
1*
b1 6
19
1>
1C
b1 G
#518080000000
0!
0*
09
0>
0C
#518090000000
1!
1*
b10 6
19
1>
1C
b10 G
#518100000000
0!
0*
09
0>
0C
#518110000000
1!
1*
b11 6
19
1>
1C
b11 G
#518120000000
0!
0*
09
0>
0C
#518130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#518140000000
0!
0*
09
0>
0C
#518150000000
1!
1*
b101 6
19
1>
1C
b101 G
#518160000000
0!
0*
09
0>
0C
#518170000000
1!
1*
b110 6
19
1>
1C
b110 G
#518180000000
0!
0*
09
0>
0C
#518190000000
1!
1*
b111 6
19
1>
1C
b111 G
#518200000000
0!
1"
0*
1+
09
1:
0>
0C
#518210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#518220000000
0!
0*
09
0>
0C
#518230000000
1!
1*
b1 6
19
1>
1C
b1 G
#518240000000
0!
0*
09
0>
0C
#518250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#518260000000
0!
0*
09
0>
0C
#518270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#518280000000
0!
0*
09
0>
0C
#518290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#518300000000
0!
0*
09
0>
0C
#518310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#518320000000
0!
0#
0*
0,
09
0>
0?
0C
#518330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#518340000000
0!
0*
09
0>
0C
#518350000000
1!
1*
19
1>
1C
#518360000000
0!
0*
09
0>
0C
#518370000000
1!
1*
19
1>
1C
#518380000000
0!
0*
09
0>
0C
#518390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#518400000000
0!
0*
09
0>
0C
#518410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#518420000000
0!
0*
09
0>
0C
#518430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#518440000000
0!
0*
09
0>
0C
#518450000000
1!
1*
b10 6
19
1>
1C
b10 G
#518460000000
0!
0*
09
0>
0C
#518470000000
1!
1*
b11 6
19
1>
1C
b11 G
#518480000000
0!
0*
09
0>
0C
#518490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#518500000000
0!
0*
09
0>
0C
#518510000000
1!
1*
b101 6
19
1>
1C
b101 G
#518520000000
0!
0*
09
0>
0C
#518530000000
1!
1*
b110 6
19
1>
1C
b110 G
#518540000000
0!
0*
09
0>
0C
#518550000000
1!
1*
b111 6
19
1>
1C
b111 G
#518560000000
0!
0*
09
0>
0C
#518570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#518580000000
0!
0*
09
0>
0C
#518590000000
1!
1*
b1 6
19
1>
1C
b1 G
#518600000000
0!
0*
09
0>
0C
#518610000000
1!
1*
b10 6
19
1>
1C
b10 G
#518620000000
0!
0*
09
0>
0C
#518630000000
1!
1*
b11 6
19
1>
1C
b11 G
#518640000000
0!
0*
09
0>
0C
#518650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#518660000000
0!
0*
09
0>
0C
#518670000000
1!
1*
b101 6
19
1>
1C
b101 G
#518680000000
0!
0*
09
0>
0C
#518690000000
1!
1*
b110 6
19
1>
1C
b110 G
#518700000000
0!
0*
09
0>
0C
#518710000000
1!
1*
b111 6
19
1>
1C
b111 G
#518720000000
0!
0*
09
0>
0C
#518730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#518740000000
0!
0*
09
0>
0C
#518750000000
1!
1*
b1 6
19
1>
1C
b1 G
#518760000000
0!
0*
09
0>
0C
#518770000000
1!
1*
b10 6
19
1>
1C
b10 G
#518780000000
0!
0*
09
0>
0C
#518790000000
1!
1*
b11 6
19
1>
1C
b11 G
#518800000000
0!
0*
09
0>
0C
#518810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#518820000000
0!
0*
09
0>
0C
#518830000000
1!
1*
b101 6
19
1>
1C
b101 G
#518840000000
0!
0*
09
0>
0C
#518850000000
1!
1*
b110 6
19
1>
1C
b110 G
#518860000000
0!
0*
09
0>
0C
#518870000000
1!
1*
b111 6
19
1>
1C
b111 G
#518880000000
0!
1"
0*
1+
09
1:
0>
0C
#518890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#518900000000
0!
0*
09
0>
0C
#518910000000
1!
1*
b1 6
19
1>
1C
b1 G
#518920000000
0!
0*
09
0>
0C
#518930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#518940000000
0!
0*
09
0>
0C
#518950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#518960000000
0!
0*
09
0>
0C
#518970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#518980000000
0!
0*
09
0>
0C
#518990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#519000000000
0!
0#
0*
0,
09
0>
0?
0C
#519010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#519020000000
0!
0*
09
0>
0C
#519030000000
1!
1*
19
1>
1C
#519040000000
0!
0*
09
0>
0C
#519050000000
1!
1*
19
1>
1C
#519060000000
0!
0*
09
0>
0C
#519070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#519080000000
0!
0*
09
0>
0C
#519090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#519100000000
0!
0*
09
0>
0C
#519110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#519120000000
0!
0*
09
0>
0C
#519130000000
1!
1*
b10 6
19
1>
1C
b10 G
#519140000000
0!
0*
09
0>
0C
#519150000000
1!
1*
b11 6
19
1>
1C
b11 G
#519160000000
0!
0*
09
0>
0C
#519170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#519180000000
0!
0*
09
0>
0C
#519190000000
1!
1*
b101 6
19
1>
1C
b101 G
#519200000000
0!
0*
09
0>
0C
#519210000000
1!
1*
b110 6
19
1>
1C
b110 G
#519220000000
0!
0*
09
0>
0C
#519230000000
1!
1*
b111 6
19
1>
1C
b111 G
#519240000000
0!
0*
09
0>
0C
#519250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#519260000000
0!
0*
09
0>
0C
#519270000000
1!
1*
b1 6
19
1>
1C
b1 G
#519280000000
0!
0*
09
0>
0C
#519290000000
1!
1*
b10 6
19
1>
1C
b10 G
#519300000000
0!
0*
09
0>
0C
#519310000000
1!
1*
b11 6
19
1>
1C
b11 G
#519320000000
0!
0*
09
0>
0C
#519330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#519340000000
0!
0*
09
0>
0C
#519350000000
1!
1*
b101 6
19
1>
1C
b101 G
#519360000000
0!
0*
09
0>
0C
#519370000000
1!
1*
b110 6
19
1>
1C
b110 G
#519380000000
0!
0*
09
0>
0C
#519390000000
1!
1*
b111 6
19
1>
1C
b111 G
#519400000000
0!
0*
09
0>
0C
#519410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#519420000000
0!
0*
09
0>
0C
#519430000000
1!
1*
b1 6
19
1>
1C
b1 G
#519440000000
0!
0*
09
0>
0C
#519450000000
1!
1*
b10 6
19
1>
1C
b10 G
#519460000000
0!
0*
09
0>
0C
#519470000000
1!
1*
b11 6
19
1>
1C
b11 G
#519480000000
0!
0*
09
0>
0C
#519490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#519500000000
0!
0*
09
0>
0C
#519510000000
1!
1*
b101 6
19
1>
1C
b101 G
#519520000000
0!
0*
09
0>
0C
#519530000000
1!
1*
b110 6
19
1>
1C
b110 G
#519540000000
0!
0*
09
0>
0C
#519550000000
1!
1*
b111 6
19
1>
1C
b111 G
#519560000000
0!
1"
0*
1+
09
1:
0>
0C
#519570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#519580000000
0!
0*
09
0>
0C
#519590000000
1!
1*
b1 6
19
1>
1C
b1 G
#519600000000
0!
0*
09
0>
0C
#519610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#519620000000
0!
0*
09
0>
0C
#519630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#519640000000
0!
0*
09
0>
0C
#519650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#519660000000
0!
0*
09
0>
0C
#519670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#519680000000
0!
0#
0*
0,
09
0>
0?
0C
#519690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#519700000000
0!
0*
09
0>
0C
#519710000000
1!
1*
19
1>
1C
#519720000000
0!
0*
09
0>
0C
#519730000000
1!
1*
19
1>
1C
#519740000000
0!
0*
09
0>
0C
#519750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#519760000000
0!
0*
09
0>
0C
#519770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#519780000000
0!
0*
09
0>
0C
#519790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#519800000000
0!
0*
09
0>
0C
#519810000000
1!
1*
b10 6
19
1>
1C
b10 G
#519820000000
0!
0*
09
0>
0C
#519830000000
1!
1*
b11 6
19
1>
1C
b11 G
#519840000000
0!
0*
09
0>
0C
#519850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#519860000000
0!
0*
09
0>
0C
#519870000000
1!
1*
b101 6
19
1>
1C
b101 G
#519880000000
0!
0*
09
0>
0C
#519890000000
1!
1*
b110 6
19
1>
1C
b110 G
#519900000000
0!
0*
09
0>
0C
#519910000000
1!
1*
b111 6
19
1>
1C
b111 G
#519920000000
0!
0*
09
0>
0C
#519930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#519940000000
0!
0*
09
0>
0C
#519950000000
1!
1*
b1 6
19
1>
1C
b1 G
#519960000000
0!
0*
09
0>
0C
#519970000000
1!
1*
b10 6
19
1>
1C
b10 G
#519980000000
0!
0*
09
0>
0C
#519990000000
1!
1*
b11 6
19
1>
1C
b11 G
#520000000000
0!
0*
09
0>
0C
#520010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#520020000000
0!
0*
09
0>
0C
#520030000000
1!
1*
b101 6
19
1>
1C
b101 G
#520040000000
0!
0*
09
0>
0C
#520050000000
1!
1*
b110 6
19
1>
1C
b110 G
#520060000000
0!
0*
09
0>
0C
#520070000000
1!
1*
b111 6
19
1>
1C
b111 G
#520080000000
0!
0*
09
0>
0C
#520090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#520100000000
0!
0*
09
0>
0C
#520110000000
1!
1*
b1 6
19
1>
1C
b1 G
#520120000000
0!
0*
09
0>
0C
#520130000000
1!
1*
b10 6
19
1>
1C
b10 G
#520140000000
0!
0*
09
0>
0C
#520150000000
1!
1*
b11 6
19
1>
1C
b11 G
#520160000000
0!
0*
09
0>
0C
#520170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#520180000000
0!
0*
09
0>
0C
#520190000000
1!
1*
b101 6
19
1>
1C
b101 G
#520200000000
0!
0*
09
0>
0C
#520210000000
1!
1*
b110 6
19
1>
1C
b110 G
#520220000000
0!
0*
09
0>
0C
#520230000000
1!
1*
b111 6
19
1>
1C
b111 G
#520240000000
0!
1"
0*
1+
09
1:
0>
0C
#520250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#520260000000
0!
0*
09
0>
0C
#520270000000
1!
1*
b1 6
19
1>
1C
b1 G
#520280000000
0!
0*
09
0>
0C
#520290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#520300000000
0!
0*
09
0>
0C
#520310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#520320000000
0!
0*
09
0>
0C
#520330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#520340000000
0!
0*
09
0>
0C
#520350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#520360000000
0!
0#
0*
0,
09
0>
0?
0C
#520370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#520380000000
0!
0*
09
0>
0C
#520390000000
1!
1*
19
1>
1C
#520400000000
0!
0*
09
0>
0C
#520410000000
1!
1*
19
1>
1C
#520420000000
0!
0*
09
0>
0C
#520430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#520440000000
0!
0*
09
0>
0C
#520450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#520460000000
0!
0*
09
0>
0C
#520470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#520480000000
0!
0*
09
0>
0C
#520490000000
1!
1*
b10 6
19
1>
1C
b10 G
#520500000000
0!
0*
09
0>
0C
#520510000000
1!
1*
b11 6
19
1>
1C
b11 G
#520520000000
0!
0*
09
0>
0C
#520530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#520540000000
0!
0*
09
0>
0C
#520550000000
1!
1*
b101 6
19
1>
1C
b101 G
#520560000000
0!
0*
09
0>
0C
#520570000000
1!
1*
b110 6
19
1>
1C
b110 G
#520580000000
0!
0*
09
0>
0C
#520590000000
1!
1*
b111 6
19
1>
1C
b111 G
#520600000000
0!
0*
09
0>
0C
#520610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#520620000000
0!
0*
09
0>
0C
#520630000000
1!
1*
b1 6
19
1>
1C
b1 G
#520640000000
0!
0*
09
0>
0C
#520650000000
1!
1*
b10 6
19
1>
1C
b10 G
#520660000000
0!
0*
09
0>
0C
#520670000000
1!
1*
b11 6
19
1>
1C
b11 G
#520680000000
0!
0*
09
0>
0C
#520690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#520700000000
0!
0*
09
0>
0C
#520710000000
1!
1*
b101 6
19
1>
1C
b101 G
#520720000000
0!
0*
09
0>
0C
#520730000000
1!
1*
b110 6
19
1>
1C
b110 G
#520740000000
0!
0*
09
0>
0C
#520750000000
1!
1*
b111 6
19
1>
1C
b111 G
#520760000000
0!
0*
09
0>
0C
#520770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#520780000000
0!
0*
09
0>
0C
#520790000000
1!
1*
b1 6
19
1>
1C
b1 G
#520800000000
0!
0*
09
0>
0C
#520810000000
1!
1*
b10 6
19
1>
1C
b10 G
#520820000000
0!
0*
09
0>
0C
#520830000000
1!
1*
b11 6
19
1>
1C
b11 G
#520840000000
0!
0*
09
0>
0C
#520850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#520860000000
0!
0*
09
0>
0C
#520870000000
1!
1*
b101 6
19
1>
1C
b101 G
#520880000000
0!
0*
09
0>
0C
#520890000000
1!
1*
b110 6
19
1>
1C
b110 G
#520900000000
0!
0*
09
0>
0C
#520910000000
1!
1*
b111 6
19
1>
1C
b111 G
#520920000000
0!
1"
0*
1+
09
1:
0>
0C
#520930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#520940000000
0!
0*
09
0>
0C
#520950000000
1!
1*
b1 6
19
1>
1C
b1 G
#520960000000
0!
0*
09
0>
0C
#520970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#520980000000
0!
0*
09
0>
0C
#520990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#521000000000
0!
0*
09
0>
0C
#521010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#521020000000
0!
0*
09
0>
0C
#521030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#521040000000
0!
0#
0*
0,
09
0>
0?
0C
#521050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#521060000000
0!
0*
09
0>
0C
#521070000000
1!
1*
19
1>
1C
#521080000000
0!
0*
09
0>
0C
#521090000000
1!
1*
19
1>
1C
#521100000000
0!
0*
09
0>
0C
#521110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#521120000000
0!
0*
09
0>
0C
#521130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#521140000000
0!
0*
09
0>
0C
#521150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#521160000000
0!
0*
09
0>
0C
#521170000000
1!
1*
b10 6
19
1>
1C
b10 G
#521180000000
0!
0*
09
0>
0C
#521190000000
1!
1*
b11 6
19
1>
1C
b11 G
#521200000000
0!
0*
09
0>
0C
#521210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#521220000000
0!
0*
09
0>
0C
#521230000000
1!
1*
b101 6
19
1>
1C
b101 G
#521240000000
0!
0*
09
0>
0C
#521250000000
1!
1*
b110 6
19
1>
1C
b110 G
#521260000000
0!
0*
09
0>
0C
#521270000000
1!
1*
b111 6
19
1>
1C
b111 G
#521280000000
0!
0*
09
0>
0C
#521290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#521300000000
0!
0*
09
0>
0C
#521310000000
1!
1*
b1 6
19
1>
1C
b1 G
#521320000000
0!
0*
09
0>
0C
#521330000000
1!
1*
b10 6
19
1>
1C
b10 G
#521340000000
0!
0*
09
0>
0C
#521350000000
1!
1*
b11 6
19
1>
1C
b11 G
#521360000000
0!
0*
09
0>
0C
#521370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#521380000000
0!
0*
09
0>
0C
#521390000000
1!
1*
b101 6
19
1>
1C
b101 G
#521400000000
0!
0*
09
0>
0C
#521410000000
1!
1*
b110 6
19
1>
1C
b110 G
#521420000000
0!
0*
09
0>
0C
#521430000000
1!
1*
b111 6
19
1>
1C
b111 G
#521440000000
0!
0*
09
0>
0C
#521450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#521460000000
0!
0*
09
0>
0C
#521470000000
1!
1*
b1 6
19
1>
1C
b1 G
#521480000000
0!
0*
09
0>
0C
#521490000000
1!
1*
b10 6
19
1>
1C
b10 G
#521500000000
0!
0*
09
0>
0C
#521510000000
1!
1*
b11 6
19
1>
1C
b11 G
#521520000000
0!
0*
09
0>
0C
#521530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#521540000000
0!
0*
09
0>
0C
#521550000000
1!
1*
b101 6
19
1>
1C
b101 G
#521560000000
0!
0*
09
0>
0C
#521570000000
1!
1*
b110 6
19
1>
1C
b110 G
#521580000000
0!
0*
09
0>
0C
#521590000000
1!
1*
b111 6
19
1>
1C
b111 G
#521600000000
0!
1"
0*
1+
09
1:
0>
0C
#521610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#521620000000
0!
0*
09
0>
0C
#521630000000
1!
1*
b1 6
19
1>
1C
b1 G
#521640000000
0!
0*
09
0>
0C
#521650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#521660000000
0!
0*
09
0>
0C
#521670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#521680000000
0!
0*
09
0>
0C
#521690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#521700000000
0!
0*
09
0>
0C
#521710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#521720000000
0!
0#
0*
0,
09
0>
0?
0C
#521730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#521740000000
0!
0*
09
0>
0C
#521750000000
1!
1*
19
1>
1C
#521760000000
0!
0*
09
0>
0C
#521770000000
1!
1*
19
1>
1C
#521780000000
0!
0*
09
0>
0C
#521790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#521800000000
0!
0*
09
0>
0C
#521810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#521820000000
0!
0*
09
0>
0C
#521830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#521840000000
0!
0*
09
0>
0C
#521850000000
1!
1*
b10 6
19
1>
1C
b10 G
#521860000000
0!
0*
09
0>
0C
#521870000000
1!
1*
b11 6
19
1>
1C
b11 G
#521880000000
0!
0*
09
0>
0C
#521890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#521900000000
0!
0*
09
0>
0C
#521910000000
1!
1*
b101 6
19
1>
1C
b101 G
#521920000000
0!
0*
09
0>
0C
#521930000000
1!
1*
b110 6
19
1>
1C
b110 G
#521940000000
0!
0*
09
0>
0C
#521950000000
1!
1*
b111 6
19
1>
1C
b111 G
#521960000000
0!
0*
09
0>
0C
#521970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#521980000000
0!
0*
09
0>
0C
#521990000000
1!
1*
b1 6
19
1>
1C
b1 G
#522000000000
0!
0*
09
0>
0C
#522010000000
1!
1*
b10 6
19
1>
1C
b10 G
#522020000000
0!
0*
09
0>
0C
#522030000000
1!
1*
b11 6
19
1>
1C
b11 G
#522040000000
0!
0*
09
0>
0C
#522050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#522060000000
0!
0*
09
0>
0C
#522070000000
1!
1*
b101 6
19
1>
1C
b101 G
#522080000000
0!
0*
09
0>
0C
#522090000000
1!
1*
b110 6
19
1>
1C
b110 G
#522100000000
0!
0*
09
0>
0C
#522110000000
1!
1*
b111 6
19
1>
1C
b111 G
#522120000000
0!
0*
09
0>
0C
#522130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#522140000000
0!
0*
09
0>
0C
#522150000000
1!
1*
b1 6
19
1>
1C
b1 G
#522160000000
0!
0*
09
0>
0C
#522170000000
1!
1*
b10 6
19
1>
1C
b10 G
#522180000000
0!
0*
09
0>
0C
#522190000000
1!
1*
b11 6
19
1>
1C
b11 G
#522200000000
0!
0*
09
0>
0C
#522210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#522220000000
0!
0*
09
0>
0C
#522230000000
1!
1*
b101 6
19
1>
1C
b101 G
#522240000000
0!
0*
09
0>
0C
#522250000000
1!
1*
b110 6
19
1>
1C
b110 G
#522260000000
0!
0*
09
0>
0C
#522270000000
1!
1*
b111 6
19
1>
1C
b111 G
#522280000000
0!
1"
0*
1+
09
1:
0>
0C
#522290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#522300000000
0!
0*
09
0>
0C
#522310000000
1!
1*
b1 6
19
1>
1C
b1 G
#522320000000
0!
0*
09
0>
0C
#522330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#522340000000
0!
0*
09
0>
0C
#522350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#522360000000
0!
0*
09
0>
0C
#522370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#522380000000
0!
0*
09
0>
0C
#522390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#522400000000
0!
0#
0*
0,
09
0>
0?
0C
#522410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#522420000000
0!
0*
09
0>
0C
#522430000000
1!
1*
19
1>
1C
#522440000000
0!
0*
09
0>
0C
#522450000000
1!
1*
19
1>
1C
#522460000000
0!
0*
09
0>
0C
#522470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#522480000000
0!
0*
09
0>
0C
#522490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#522500000000
0!
0*
09
0>
0C
#522510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#522520000000
0!
0*
09
0>
0C
#522530000000
1!
1*
b10 6
19
1>
1C
b10 G
#522540000000
0!
0*
09
0>
0C
#522550000000
1!
1*
b11 6
19
1>
1C
b11 G
#522560000000
0!
0*
09
0>
0C
#522570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#522580000000
0!
0*
09
0>
0C
#522590000000
1!
1*
b101 6
19
1>
1C
b101 G
#522600000000
0!
0*
09
0>
0C
#522610000000
1!
1*
b110 6
19
1>
1C
b110 G
#522620000000
0!
0*
09
0>
0C
#522630000000
1!
1*
b111 6
19
1>
1C
b111 G
#522640000000
0!
0*
09
0>
0C
#522650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#522660000000
0!
0*
09
0>
0C
#522670000000
1!
1*
b1 6
19
1>
1C
b1 G
#522680000000
0!
0*
09
0>
0C
#522690000000
1!
1*
b10 6
19
1>
1C
b10 G
#522700000000
0!
0*
09
0>
0C
#522710000000
1!
1*
b11 6
19
1>
1C
b11 G
#522720000000
0!
0*
09
0>
0C
#522730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#522740000000
0!
0*
09
0>
0C
#522750000000
1!
1*
b101 6
19
1>
1C
b101 G
#522760000000
0!
0*
09
0>
0C
#522770000000
1!
1*
b110 6
19
1>
1C
b110 G
#522780000000
0!
0*
09
0>
0C
#522790000000
1!
1*
b111 6
19
1>
1C
b111 G
#522800000000
0!
0*
09
0>
0C
#522810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#522820000000
0!
0*
09
0>
0C
#522830000000
1!
1*
b1 6
19
1>
1C
b1 G
#522840000000
0!
0*
09
0>
0C
#522850000000
1!
1*
b10 6
19
1>
1C
b10 G
#522860000000
0!
0*
09
0>
0C
#522870000000
1!
1*
b11 6
19
1>
1C
b11 G
#522880000000
0!
0*
09
0>
0C
#522890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#522900000000
0!
0*
09
0>
0C
#522910000000
1!
1*
b101 6
19
1>
1C
b101 G
#522920000000
0!
0*
09
0>
0C
#522930000000
1!
1*
b110 6
19
1>
1C
b110 G
#522940000000
0!
0*
09
0>
0C
#522950000000
1!
1*
b111 6
19
1>
1C
b111 G
#522960000000
0!
1"
0*
1+
09
1:
0>
0C
#522970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#522980000000
0!
0*
09
0>
0C
#522990000000
1!
1*
b1 6
19
1>
1C
b1 G
#523000000000
0!
0*
09
0>
0C
#523010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#523020000000
0!
0*
09
0>
0C
#523030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#523040000000
0!
0*
09
0>
0C
#523050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#523060000000
0!
0*
09
0>
0C
#523070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#523080000000
0!
0#
0*
0,
09
0>
0?
0C
#523090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#523100000000
0!
0*
09
0>
0C
#523110000000
1!
1*
19
1>
1C
#523120000000
0!
0*
09
0>
0C
#523130000000
1!
1*
19
1>
1C
#523140000000
0!
0*
09
0>
0C
#523150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#523160000000
0!
0*
09
0>
0C
#523170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#523180000000
0!
0*
09
0>
0C
#523190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#523200000000
0!
0*
09
0>
0C
#523210000000
1!
1*
b10 6
19
1>
1C
b10 G
#523220000000
0!
0*
09
0>
0C
#523230000000
1!
1*
b11 6
19
1>
1C
b11 G
#523240000000
0!
0*
09
0>
0C
#523250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#523260000000
0!
0*
09
0>
0C
#523270000000
1!
1*
b101 6
19
1>
1C
b101 G
#523280000000
0!
0*
09
0>
0C
#523290000000
1!
1*
b110 6
19
1>
1C
b110 G
#523300000000
0!
0*
09
0>
0C
#523310000000
1!
1*
b111 6
19
1>
1C
b111 G
#523320000000
0!
0*
09
0>
0C
#523330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#523340000000
0!
0*
09
0>
0C
#523350000000
1!
1*
b1 6
19
1>
1C
b1 G
#523360000000
0!
0*
09
0>
0C
#523370000000
1!
1*
b10 6
19
1>
1C
b10 G
#523380000000
0!
0*
09
0>
0C
#523390000000
1!
1*
b11 6
19
1>
1C
b11 G
#523400000000
0!
0*
09
0>
0C
#523410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#523420000000
0!
0*
09
0>
0C
#523430000000
1!
1*
b101 6
19
1>
1C
b101 G
#523440000000
0!
0*
09
0>
0C
#523450000000
1!
1*
b110 6
19
1>
1C
b110 G
#523460000000
0!
0*
09
0>
0C
#523470000000
1!
1*
b111 6
19
1>
1C
b111 G
#523480000000
0!
0*
09
0>
0C
#523490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#523500000000
0!
0*
09
0>
0C
#523510000000
1!
1*
b1 6
19
1>
1C
b1 G
#523520000000
0!
0*
09
0>
0C
#523530000000
1!
1*
b10 6
19
1>
1C
b10 G
#523540000000
0!
0*
09
0>
0C
#523550000000
1!
1*
b11 6
19
1>
1C
b11 G
#523560000000
0!
0*
09
0>
0C
#523570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#523580000000
0!
0*
09
0>
0C
#523590000000
1!
1*
b101 6
19
1>
1C
b101 G
#523600000000
0!
0*
09
0>
0C
#523610000000
1!
1*
b110 6
19
1>
1C
b110 G
#523620000000
0!
0*
09
0>
0C
#523630000000
1!
1*
b111 6
19
1>
1C
b111 G
#523640000000
0!
1"
0*
1+
09
1:
0>
0C
#523650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#523660000000
0!
0*
09
0>
0C
#523670000000
1!
1*
b1 6
19
1>
1C
b1 G
#523680000000
0!
0*
09
0>
0C
#523690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#523700000000
0!
0*
09
0>
0C
#523710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#523720000000
0!
0*
09
0>
0C
#523730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#523740000000
0!
0*
09
0>
0C
#523750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#523760000000
0!
0#
0*
0,
09
0>
0?
0C
#523770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#523780000000
0!
0*
09
0>
0C
#523790000000
1!
1*
19
1>
1C
#523800000000
0!
0*
09
0>
0C
#523810000000
1!
1*
19
1>
1C
#523820000000
0!
0*
09
0>
0C
#523830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#523840000000
0!
0*
09
0>
0C
#523850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#523860000000
0!
0*
09
0>
0C
#523870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#523880000000
0!
0*
09
0>
0C
#523890000000
1!
1*
b10 6
19
1>
1C
b10 G
#523900000000
0!
0*
09
0>
0C
#523910000000
1!
1*
b11 6
19
1>
1C
b11 G
#523920000000
0!
0*
09
0>
0C
#523930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#523940000000
0!
0*
09
0>
0C
#523950000000
1!
1*
b101 6
19
1>
1C
b101 G
#523960000000
0!
0*
09
0>
0C
#523970000000
1!
1*
b110 6
19
1>
1C
b110 G
#523980000000
0!
0*
09
0>
0C
#523990000000
1!
1*
b111 6
19
1>
1C
b111 G
#524000000000
0!
0*
09
0>
0C
#524010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#524020000000
0!
0*
09
0>
0C
#524030000000
1!
1*
b1 6
19
1>
1C
b1 G
#524040000000
0!
0*
09
0>
0C
#524050000000
1!
1*
b10 6
19
1>
1C
b10 G
#524060000000
0!
0*
09
0>
0C
#524070000000
1!
1*
b11 6
19
1>
1C
b11 G
#524080000000
0!
0*
09
0>
0C
#524090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#524100000000
0!
0*
09
0>
0C
#524110000000
1!
1*
b101 6
19
1>
1C
b101 G
#524120000000
0!
0*
09
0>
0C
#524130000000
1!
1*
b110 6
19
1>
1C
b110 G
#524140000000
0!
0*
09
0>
0C
#524150000000
1!
1*
b111 6
19
1>
1C
b111 G
#524160000000
0!
0*
09
0>
0C
#524170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#524180000000
0!
0*
09
0>
0C
#524190000000
1!
1*
b1 6
19
1>
1C
b1 G
#524200000000
0!
0*
09
0>
0C
#524210000000
1!
1*
b10 6
19
1>
1C
b10 G
#524220000000
0!
0*
09
0>
0C
#524230000000
1!
1*
b11 6
19
1>
1C
b11 G
#524240000000
0!
0*
09
0>
0C
#524250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#524260000000
0!
0*
09
0>
0C
#524270000000
1!
1*
b101 6
19
1>
1C
b101 G
#524280000000
0!
0*
09
0>
0C
#524290000000
1!
1*
b110 6
19
1>
1C
b110 G
#524300000000
0!
0*
09
0>
0C
#524310000000
1!
1*
b111 6
19
1>
1C
b111 G
#524320000000
0!
1"
0*
1+
09
1:
0>
0C
#524330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#524340000000
0!
0*
09
0>
0C
#524350000000
1!
1*
b1 6
19
1>
1C
b1 G
#524360000000
0!
0*
09
0>
0C
#524370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#524380000000
0!
0*
09
0>
0C
#524390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#524400000000
0!
0*
09
0>
0C
#524410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#524420000000
0!
0*
09
0>
0C
#524430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#524440000000
0!
0#
0*
0,
09
0>
0?
0C
#524450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#524460000000
0!
0*
09
0>
0C
#524470000000
1!
1*
19
1>
1C
#524480000000
0!
0*
09
0>
0C
#524490000000
1!
1*
19
1>
1C
#524500000000
0!
0*
09
0>
0C
#524510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#524520000000
0!
0*
09
0>
0C
#524530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#524540000000
0!
0*
09
0>
0C
#524550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#524560000000
0!
0*
09
0>
0C
#524570000000
1!
1*
b10 6
19
1>
1C
b10 G
#524580000000
0!
0*
09
0>
0C
#524590000000
1!
1*
b11 6
19
1>
1C
b11 G
#524600000000
0!
0*
09
0>
0C
#524610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#524620000000
0!
0*
09
0>
0C
#524630000000
1!
1*
b101 6
19
1>
1C
b101 G
#524640000000
0!
0*
09
0>
0C
#524650000000
1!
1*
b110 6
19
1>
1C
b110 G
#524660000000
0!
0*
09
0>
0C
#524670000000
1!
1*
b111 6
19
1>
1C
b111 G
#524680000000
0!
0*
09
0>
0C
#524690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#524700000000
0!
0*
09
0>
0C
#524710000000
1!
1*
b1 6
19
1>
1C
b1 G
#524720000000
0!
0*
09
0>
0C
#524730000000
1!
1*
b10 6
19
1>
1C
b10 G
#524740000000
0!
0*
09
0>
0C
#524750000000
1!
1*
b11 6
19
1>
1C
b11 G
#524760000000
0!
0*
09
0>
0C
#524770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#524780000000
0!
0*
09
0>
0C
#524790000000
1!
1*
b101 6
19
1>
1C
b101 G
#524800000000
0!
0*
09
0>
0C
#524810000000
1!
1*
b110 6
19
1>
1C
b110 G
#524820000000
0!
0*
09
0>
0C
#524830000000
1!
1*
b111 6
19
1>
1C
b111 G
#524840000000
0!
0*
09
0>
0C
#524850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#524860000000
0!
0*
09
0>
0C
#524870000000
1!
1*
b1 6
19
1>
1C
b1 G
#524880000000
0!
0*
09
0>
0C
#524890000000
1!
1*
b10 6
19
1>
1C
b10 G
#524900000000
0!
0*
09
0>
0C
#524910000000
1!
1*
b11 6
19
1>
1C
b11 G
#524920000000
0!
0*
09
0>
0C
#524930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#524940000000
0!
0*
09
0>
0C
#524950000000
1!
1*
b101 6
19
1>
1C
b101 G
#524960000000
0!
0*
09
0>
0C
#524970000000
1!
1*
b110 6
19
1>
1C
b110 G
#524980000000
0!
0*
09
0>
0C
#524990000000
1!
1*
b111 6
19
1>
1C
b111 G
#525000000000
0!
1"
0*
1+
09
1:
0>
0C
#525010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#525020000000
0!
0*
09
0>
0C
#525030000000
1!
1*
b1 6
19
1>
1C
b1 G
#525040000000
0!
0*
09
0>
0C
#525050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#525060000000
0!
0*
09
0>
0C
#525070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#525080000000
0!
0*
09
0>
0C
#525090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#525100000000
0!
0*
09
0>
0C
#525110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#525120000000
0!
0#
0*
0,
09
0>
0?
0C
#525130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#525140000000
0!
0*
09
0>
0C
#525150000000
1!
1*
19
1>
1C
#525160000000
0!
0*
09
0>
0C
#525170000000
1!
1*
19
1>
1C
#525180000000
0!
0*
09
0>
0C
#525190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#525200000000
0!
0*
09
0>
0C
#525210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#525220000000
0!
0*
09
0>
0C
#525230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#525240000000
0!
0*
09
0>
0C
#525250000000
1!
1*
b10 6
19
1>
1C
b10 G
#525260000000
0!
0*
09
0>
0C
#525270000000
1!
1*
b11 6
19
1>
1C
b11 G
#525280000000
0!
0*
09
0>
0C
#525290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#525300000000
0!
0*
09
0>
0C
#525310000000
1!
1*
b101 6
19
1>
1C
b101 G
#525320000000
0!
0*
09
0>
0C
#525330000000
1!
1*
b110 6
19
1>
1C
b110 G
#525340000000
0!
0*
09
0>
0C
#525350000000
1!
1*
b111 6
19
1>
1C
b111 G
#525360000000
0!
0*
09
0>
0C
#525370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#525380000000
0!
0*
09
0>
0C
#525390000000
1!
1*
b1 6
19
1>
1C
b1 G
#525400000000
0!
0*
09
0>
0C
#525410000000
1!
1*
b10 6
19
1>
1C
b10 G
#525420000000
0!
0*
09
0>
0C
#525430000000
1!
1*
b11 6
19
1>
1C
b11 G
#525440000000
0!
0*
09
0>
0C
#525450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#525460000000
0!
0*
09
0>
0C
#525470000000
1!
1*
b101 6
19
1>
1C
b101 G
#525480000000
0!
0*
09
0>
0C
#525490000000
1!
1*
b110 6
19
1>
1C
b110 G
#525500000000
0!
0*
09
0>
0C
#525510000000
1!
1*
b111 6
19
1>
1C
b111 G
#525520000000
0!
0*
09
0>
0C
#525530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#525540000000
0!
0*
09
0>
0C
#525550000000
1!
1*
b1 6
19
1>
1C
b1 G
#525560000000
0!
0*
09
0>
0C
#525570000000
1!
1*
b10 6
19
1>
1C
b10 G
#525580000000
0!
0*
09
0>
0C
#525590000000
1!
1*
b11 6
19
1>
1C
b11 G
#525600000000
0!
0*
09
0>
0C
#525610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#525620000000
0!
0*
09
0>
0C
#525630000000
1!
1*
b101 6
19
1>
1C
b101 G
#525640000000
0!
0*
09
0>
0C
#525650000000
1!
1*
b110 6
19
1>
1C
b110 G
#525660000000
0!
0*
09
0>
0C
#525670000000
1!
1*
b111 6
19
1>
1C
b111 G
#525680000000
0!
1"
0*
1+
09
1:
0>
0C
#525690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#525700000000
0!
0*
09
0>
0C
#525710000000
1!
1*
b1 6
19
1>
1C
b1 G
#525720000000
0!
0*
09
0>
0C
#525730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#525740000000
0!
0*
09
0>
0C
#525750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#525760000000
0!
0*
09
0>
0C
#525770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#525780000000
0!
0*
09
0>
0C
#525790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#525800000000
0!
0#
0*
0,
09
0>
0?
0C
#525810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#525820000000
0!
0*
09
0>
0C
#525830000000
1!
1*
19
1>
1C
#525840000000
0!
0*
09
0>
0C
#525850000000
1!
1*
19
1>
1C
#525860000000
0!
0*
09
0>
0C
#525870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#525880000000
0!
0*
09
0>
0C
#525890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#525900000000
0!
0*
09
0>
0C
#525910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#525920000000
0!
0*
09
0>
0C
#525930000000
1!
1*
b10 6
19
1>
1C
b10 G
#525940000000
0!
0*
09
0>
0C
#525950000000
1!
1*
b11 6
19
1>
1C
b11 G
#525960000000
0!
0*
09
0>
0C
#525970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#525980000000
0!
0*
09
0>
0C
#525990000000
1!
1*
b101 6
19
1>
1C
b101 G
#526000000000
0!
0*
09
0>
0C
#526010000000
1!
1*
b110 6
19
1>
1C
b110 G
#526020000000
0!
0*
09
0>
0C
#526030000000
1!
1*
b111 6
19
1>
1C
b111 G
#526040000000
0!
0*
09
0>
0C
#526050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#526060000000
0!
0*
09
0>
0C
#526070000000
1!
1*
b1 6
19
1>
1C
b1 G
#526080000000
0!
0*
09
0>
0C
#526090000000
1!
1*
b10 6
19
1>
1C
b10 G
#526100000000
0!
0*
09
0>
0C
#526110000000
1!
1*
b11 6
19
1>
1C
b11 G
#526120000000
0!
0*
09
0>
0C
#526130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#526140000000
0!
0*
09
0>
0C
#526150000000
1!
1*
b101 6
19
1>
1C
b101 G
#526160000000
0!
0*
09
0>
0C
#526170000000
1!
1*
b110 6
19
1>
1C
b110 G
#526180000000
0!
0*
09
0>
0C
#526190000000
1!
1*
b111 6
19
1>
1C
b111 G
#526200000000
0!
0*
09
0>
0C
#526210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#526220000000
0!
0*
09
0>
0C
#526230000000
1!
1*
b1 6
19
1>
1C
b1 G
#526240000000
0!
0*
09
0>
0C
#526250000000
1!
1*
b10 6
19
1>
1C
b10 G
#526260000000
0!
0*
09
0>
0C
#526270000000
1!
1*
b11 6
19
1>
1C
b11 G
#526280000000
0!
0*
09
0>
0C
#526290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#526300000000
0!
0*
09
0>
0C
#526310000000
1!
1*
b101 6
19
1>
1C
b101 G
#526320000000
0!
0*
09
0>
0C
#526330000000
1!
1*
b110 6
19
1>
1C
b110 G
#526340000000
0!
0*
09
0>
0C
#526350000000
1!
1*
b111 6
19
1>
1C
b111 G
#526360000000
0!
1"
0*
1+
09
1:
0>
0C
#526370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#526380000000
0!
0*
09
0>
0C
#526390000000
1!
1*
b1 6
19
1>
1C
b1 G
#526400000000
0!
0*
09
0>
0C
#526410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#526420000000
0!
0*
09
0>
0C
#526430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#526440000000
0!
0*
09
0>
0C
#526450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#526460000000
0!
0*
09
0>
0C
#526470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#526480000000
0!
0#
0*
0,
09
0>
0?
0C
#526490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#526500000000
0!
0*
09
0>
0C
#526510000000
1!
1*
19
1>
1C
#526520000000
0!
0*
09
0>
0C
#526530000000
1!
1*
19
1>
1C
#526540000000
0!
0*
09
0>
0C
#526550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#526560000000
0!
0*
09
0>
0C
#526570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#526580000000
0!
0*
09
0>
0C
#526590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#526600000000
0!
0*
09
0>
0C
#526610000000
1!
1*
b10 6
19
1>
1C
b10 G
#526620000000
0!
0*
09
0>
0C
#526630000000
1!
1*
b11 6
19
1>
1C
b11 G
#526640000000
0!
0*
09
0>
0C
#526650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#526660000000
0!
0*
09
0>
0C
#526670000000
1!
1*
b101 6
19
1>
1C
b101 G
#526680000000
0!
0*
09
0>
0C
#526690000000
1!
1*
b110 6
19
1>
1C
b110 G
#526700000000
0!
0*
09
0>
0C
#526710000000
1!
1*
b111 6
19
1>
1C
b111 G
#526720000000
0!
0*
09
0>
0C
#526730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#526740000000
0!
0*
09
0>
0C
#526750000000
1!
1*
b1 6
19
1>
1C
b1 G
#526760000000
0!
0*
09
0>
0C
#526770000000
1!
1*
b10 6
19
1>
1C
b10 G
#526780000000
0!
0*
09
0>
0C
#526790000000
1!
1*
b11 6
19
1>
1C
b11 G
#526800000000
0!
0*
09
0>
0C
#526810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#526820000000
0!
0*
09
0>
0C
#526830000000
1!
1*
b101 6
19
1>
1C
b101 G
#526840000000
0!
0*
09
0>
0C
#526850000000
1!
1*
b110 6
19
1>
1C
b110 G
#526860000000
0!
0*
09
0>
0C
#526870000000
1!
1*
b111 6
19
1>
1C
b111 G
#526880000000
0!
0*
09
0>
0C
#526890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#526900000000
0!
0*
09
0>
0C
#526910000000
1!
1*
b1 6
19
1>
1C
b1 G
#526920000000
0!
0*
09
0>
0C
#526930000000
1!
1*
b10 6
19
1>
1C
b10 G
#526940000000
0!
0*
09
0>
0C
#526950000000
1!
1*
b11 6
19
1>
1C
b11 G
#526960000000
0!
0*
09
0>
0C
#526970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#526980000000
0!
0*
09
0>
0C
#526990000000
1!
1*
b101 6
19
1>
1C
b101 G
#527000000000
0!
0*
09
0>
0C
#527010000000
1!
1*
b110 6
19
1>
1C
b110 G
#527020000000
0!
0*
09
0>
0C
#527030000000
1!
1*
b111 6
19
1>
1C
b111 G
#527040000000
0!
1"
0*
1+
09
1:
0>
0C
#527050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#527060000000
0!
0*
09
0>
0C
#527070000000
1!
1*
b1 6
19
1>
1C
b1 G
#527080000000
0!
0*
09
0>
0C
#527090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#527100000000
0!
0*
09
0>
0C
#527110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#527120000000
0!
0*
09
0>
0C
#527130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#527140000000
0!
0*
09
0>
0C
#527150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#527160000000
0!
0#
0*
0,
09
0>
0?
0C
#527170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#527180000000
0!
0*
09
0>
0C
#527190000000
1!
1*
19
1>
1C
#527200000000
0!
0*
09
0>
0C
#527210000000
1!
1*
19
1>
1C
#527220000000
0!
0*
09
0>
0C
#527230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#527240000000
0!
0*
09
0>
0C
#527250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#527260000000
0!
0*
09
0>
0C
#527270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#527280000000
0!
0*
09
0>
0C
#527290000000
1!
1*
b10 6
19
1>
1C
b10 G
#527300000000
0!
0*
09
0>
0C
#527310000000
1!
1*
b11 6
19
1>
1C
b11 G
#527320000000
0!
0*
09
0>
0C
#527330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#527340000000
0!
0*
09
0>
0C
#527350000000
1!
1*
b101 6
19
1>
1C
b101 G
#527360000000
0!
0*
09
0>
0C
#527370000000
1!
1*
b110 6
19
1>
1C
b110 G
#527380000000
0!
0*
09
0>
0C
#527390000000
1!
1*
b111 6
19
1>
1C
b111 G
#527400000000
0!
0*
09
0>
0C
#527410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#527420000000
0!
0*
09
0>
0C
#527430000000
1!
1*
b1 6
19
1>
1C
b1 G
#527440000000
0!
0*
09
0>
0C
#527450000000
1!
1*
b10 6
19
1>
1C
b10 G
#527460000000
0!
0*
09
0>
0C
#527470000000
1!
1*
b11 6
19
1>
1C
b11 G
#527480000000
0!
0*
09
0>
0C
#527490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#527500000000
0!
0*
09
0>
0C
#527510000000
1!
1*
b101 6
19
1>
1C
b101 G
#527520000000
0!
0*
09
0>
0C
#527530000000
1!
1*
b110 6
19
1>
1C
b110 G
#527540000000
0!
0*
09
0>
0C
#527550000000
1!
1*
b111 6
19
1>
1C
b111 G
#527560000000
0!
0*
09
0>
0C
#527570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#527580000000
0!
0*
09
0>
0C
#527590000000
1!
1*
b1 6
19
1>
1C
b1 G
#527600000000
0!
0*
09
0>
0C
#527610000000
1!
1*
b10 6
19
1>
1C
b10 G
#527620000000
0!
0*
09
0>
0C
#527630000000
1!
1*
b11 6
19
1>
1C
b11 G
#527640000000
0!
0*
09
0>
0C
#527650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#527660000000
0!
0*
09
0>
0C
#527670000000
1!
1*
b101 6
19
1>
1C
b101 G
#527680000000
0!
0*
09
0>
0C
#527690000000
1!
1*
b110 6
19
1>
1C
b110 G
#527700000000
0!
0*
09
0>
0C
#527710000000
1!
1*
b111 6
19
1>
1C
b111 G
#527720000000
0!
1"
0*
1+
09
1:
0>
0C
#527730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#527740000000
0!
0*
09
0>
0C
#527750000000
1!
1*
b1 6
19
1>
1C
b1 G
#527760000000
0!
0*
09
0>
0C
#527770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#527780000000
0!
0*
09
0>
0C
#527790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#527800000000
0!
0*
09
0>
0C
#527810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#527820000000
0!
0*
09
0>
0C
#527830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#527840000000
0!
0#
0*
0,
09
0>
0?
0C
#527850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#527860000000
0!
0*
09
0>
0C
#527870000000
1!
1*
19
1>
1C
#527880000000
0!
0*
09
0>
0C
#527890000000
1!
1*
19
1>
1C
#527900000000
0!
0*
09
0>
0C
#527910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#527920000000
0!
0*
09
0>
0C
#527930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#527940000000
0!
0*
09
0>
0C
#527950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#527960000000
0!
0*
09
0>
0C
#527970000000
1!
1*
b10 6
19
1>
1C
b10 G
#527980000000
0!
0*
09
0>
0C
#527990000000
1!
1*
b11 6
19
1>
1C
b11 G
#528000000000
0!
0*
09
0>
0C
#528010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#528020000000
0!
0*
09
0>
0C
#528030000000
1!
1*
b101 6
19
1>
1C
b101 G
#528040000000
0!
0*
09
0>
0C
#528050000000
1!
1*
b110 6
19
1>
1C
b110 G
#528060000000
0!
0*
09
0>
0C
#528070000000
1!
1*
b111 6
19
1>
1C
b111 G
#528080000000
0!
0*
09
0>
0C
#528090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#528100000000
0!
0*
09
0>
0C
#528110000000
1!
1*
b1 6
19
1>
1C
b1 G
#528120000000
0!
0*
09
0>
0C
#528130000000
1!
1*
b10 6
19
1>
1C
b10 G
#528140000000
0!
0*
09
0>
0C
#528150000000
1!
1*
b11 6
19
1>
1C
b11 G
#528160000000
0!
0*
09
0>
0C
#528170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#528180000000
0!
0*
09
0>
0C
#528190000000
1!
1*
b101 6
19
1>
1C
b101 G
#528200000000
0!
0*
09
0>
0C
#528210000000
1!
1*
b110 6
19
1>
1C
b110 G
#528220000000
0!
0*
09
0>
0C
#528230000000
1!
1*
b111 6
19
1>
1C
b111 G
#528240000000
0!
0*
09
0>
0C
#528250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#528260000000
0!
0*
09
0>
0C
#528270000000
1!
1*
b1 6
19
1>
1C
b1 G
#528280000000
0!
0*
09
0>
0C
#528290000000
1!
1*
b10 6
19
1>
1C
b10 G
#528300000000
0!
0*
09
0>
0C
#528310000000
1!
1*
b11 6
19
1>
1C
b11 G
#528320000000
0!
0*
09
0>
0C
#528330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#528340000000
0!
0*
09
0>
0C
#528350000000
1!
1*
b101 6
19
1>
1C
b101 G
#528360000000
0!
0*
09
0>
0C
#528370000000
1!
1*
b110 6
19
1>
1C
b110 G
#528380000000
0!
0*
09
0>
0C
#528390000000
1!
1*
b111 6
19
1>
1C
b111 G
#528400000000
0!
1"
0*
1+
09
1:
0>
0C
#528410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#528420000000
0!
0*
09
0>
0C
#528430000000
1!
1*
b1 6
19
1>
1C
b1 G
#528440000000
0!
0*
09
0>
0C
#528450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#528460000000
0!
0*
09
0>
0C
#528470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#528480000000
0!
0*
09
0>
0C
#528490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#528500000000
0!
0*
09
0>
0C
#528510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#528520000000
0!
0#
0*
0,
09
0>
0?
0C
#528530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#528540000000
0!
0*
09
0>
0C
#528550000000
1!
1*
19
1>
1C
#528560000000
0!
0*
09
0>
0C
#528570000000
1!
1*
19
1>
1C
#528580000000
0!
0*
09
0>
0C
#528590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#528600000000
0!
0*
09
0>
0C
#528610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#528620000000
0!
0*
09
0>
0C
#528630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#528640000000
0!
0*
09
0>
0C
#528650000000
1!
1*
b10 6
19
1>
1C
b10 G
#528660000000
0!
0*
09
0>
0C
#528670000000
1!
1*
b11 6
19
1>
1C
b11 G
#528680000000
0!
0*
09
0>
0C
#528690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#528700000000
0!
0*
09
0>
0C
#528710000000
1!
1*
b101 6
19
1>
1C
b101 G
#528720000000
0!
0*
09
0>
0C
#528730000000
1!
1*
b110 6
19
1>
1C
b110 G
#528740000000
0!
0*
09
0>
0C
#528750000000
1!
1*
b111 6
19
1>
1C
b111 G
#528760000000
0!
0*
09
0>
0C
#528770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#528780000000
0!
0*
09
0>
0C
#528790000000
1!
1*
b1 6
19
1>
1C
b1 G
#528800000000
0!
0*
09
0>
0C
#528810000000
1!
1*
b10 6
19
1>
1C
b10 G
#528820000000
0!
0*
09
0>
0C
#528830000000
1!
1*
b11 6
19
1>
1C
b11 G
#528840000000
0!
0*
09
0>
0C
#528850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#528860000000
0!
0*
09
0>
0C
#528870000000
1!
1*
b101 6
19
1>
1C
b101 G
#528880000000
0!
0*
09
0>
0C
#528890000000
1!
1*
b110 6
19
1>
1C
b110 G
#528900000000
0!
0*
09
0>
0C
#528910000000
1!
1*
b111 6
19
1>
1C
b111 G
#528920000000
0!
0*
09
0>
0C
#528930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#528940000000
0!
0*
09
0>
0C
#528950000000
1!
1*
b1 6
19
1>
1C
b1 G
#528960000000
0!
0*
09
0>
0C
#528970000000
1!
1*
b10 6
19
1>
1C
b10 G
#528980000000
0!
0*
09
0>
0C
#528990000000
1!
1*
b11 6
19
1>
1C
b11 G
#529000000000
0!
0*
09
0>
0C
#529010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#529020000000
0!
0*
09
0>
0C
#529030000000
1!
1*
b101 6
19
1>
1C
b101 G
#529040000000
0!
0*
09
0>
0C
#529050000000
1!
1*
b110 6
19
1>
1C
b110 G
#529060000000
0!
0*
09
0>
0C
#529070000000
1!
1*
b111 6
19
1>
1C
b111 G
#529080000000
0!
1"
0*
1+
09
1:
0>
0C
#529090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#529100000000
0!
0*
09
0>
0C
#529110000000
1!
1*
b1 6
19
1>
1C
b1 G
#529120000000
0!
0*
09
0>
0C
#529130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#529140000000
0!
0*
09
0>
0C
#529150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#529160000000
0!
0*
09
0>
0C
#529170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#529180000000
0!
0*
09
0>
0C
#529190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#529200000000
0!
0#
0*
0,
09
0>
0?
0C
#529210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#529220000000
0!
0*
09
0>
0C
#529230000000
1!
1*
19
1>
1C
#529240000000
0!
0*
09
0>
0C
#529250000000
1!
1*
19
1>
1C
#529260000000
0!
0*
09
0>
0C
#529270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#529280000000
0!
0*
09
0>
0C
#529290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#529300000000
0!
0*
09
0>
0C
#529310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#529320000000
0!
0*
09
0>
0C
#529330000000
1!
1*
b10 6
19
1>
1C
b10 G
#529340000000
0!
0*
09
0>
0C
#529350000000
1!
1*
b11 6
19
1>
1C
b11 G
#529360000000
0!
0*
09
0>
0C
#529370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#529380000000
0!
0*
09
0>
0C
#529390000000
1!
1*
b101 6
19
1>
1C
b101 G
#529400000000
0!
0*
09
0>
0C
#529410000000
1!
1*
b110 6
19
1>
1C
b110 G
#529420000000
0!
0*
09
0>
0C
#529430000000
1!
1*
b111 6
19
1>
1C
b111 G
#529440000000
0!
0*
09
0>
0C
#529450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#529460000000
0!
0*
09
0>
0C
#529470000000
1!
1*
b1 6
19
1>
1C
b1 G
#529480000000
0!
0*
09
0>
0C
#529490000000
1!
1*
b10 6
19
1>
1C
b10 G
#529500000000
0!
0*
09
0>
0C
#529510000000
1!
1*
b11 6
19
1>
1C
b11 G
#529520000000
0!
0*
09
0>
0C
#529530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#529540000000
0!
0*
09
0>
0C
#529550000000
1!
1*
b101 6
19
1>
1C
b101 G
#529560000000
0!
0*
09
0>
0C
#529570000000
1!
1*
b110 6
19
1>
1C
b110 G
#529580000000
0!
0*
09
0>
0C
#529590000000
1!
1*
b111 6
19
1>
1C
b111 G
#529600000000
0!
0*
09
0>
0C
#529610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#529620000000
0!
0*
09
0>
0C
#529630000000
1!
1*
b1 6
19
1>
1C
b1 G
#529640000000
0!
0*
09
0>
0C
#529650000000
1!
1*
b10 6
19
1>
1C
b10 G
#529660000000
0!
0*
09
0>
0C
#529670000000
1!
1*
b11 6
19
1>
1C
b11 G
#529680000000
0!
0*
09
0>
0C
#529690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#529700000000
0!
0*
09
0>
0C
#529710000000
1!
1*
b101 6
19
1>
1C
b101 G
#529720000000
0!
0*
09
0>
0C
#529730000000
1!
1*
b110 6
19
1>
1C
b110 G
#529740000000
0!
0*
09
0>
0C
#529750000000
1!
1*
b111 6
19
1>
1C
b111 G
#529760000000
0!
1"
0*
1+
09
1:
0>
0C
#529770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#529780000000
0!
0*
09
0>
0C
#529790000000
1!
1*
b1 6
19
1>
1C
b1 G
#529800000000
0!
0*
09
0>
0C
#529810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#529820000000
0!
0*
09
0>
0C
#529830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#529840000000
0!
0*
09
0>
0C
#529850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#529860000000
0!
0*
09
0>
0C
#529870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#529880000000
0!
0#
0*
0,
09
0>
0?
0C
#529890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#529900000000
0!
0*
09
0>
0C
#529910000000
1!
1*
19
1>
1C
#529920000000
0!
0*
09
0>
0C
#529930000000
1!
1*
19
1>
1C
#529940000000
0!
0*
09
0>
0C
#529950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#529960000000
0!
0*
09
0>
0C
#529970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#529980000000
0!
0*
09
0>
0C
#529990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#530000000000
0!
0*
09
0>
0C
#530010000000
1!
1*
b10 6
19
1>
1C
b10 G
#530020000000
0!
0*
09
0>
0C
#530030000000
1!
1*
b11 6
19
1>
1C
b11 G
#530040000000
0!
0*
09
0>
0C
#530050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#530060000000
0!
0*
09
0>
0C
#530070000000
1!
1*
b101 6
19
1>
1C
b101 G
#530080000000
0!
0*
09
0>
0C
#530090000000
1!
1*
b110 6
19
1>
1C
b110 G
#530100000000
0!
0*
09
0>
0C
#530110000000
1!
1*
b111 6
19
1>
1C
b111 G
#530120000000
0!
0*
09
0>
0C
#530130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#530140000000
0!
0*
09
0>
0C
#530150000000
1!
1*
b1 6
19
1>
1C
b1 G
#530160000000
0!
0*
09
0>
0C
#530170000000
1!
1*
b10 6
19
1>
1C
b10 G
#530180000000
0!
0*
09
0>
0C
#530190000000
1!
1*
b11 6
19
1>
1C
b11 G
#530200000000
0!
0*
09
0>
0C
#530210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#530220000000
0!
0*
09
0>
0C
#530230000000
1!
1*
b101 6
19
1>
1C
b101 G
#530240000000
0!
0*
09
0>
0C
#530250000000
1!
1*
b110 6
19
1>
1C
b110 G
#530260000000
0!
0*
09
0>
0C
#530270000000
1!
1*
b111 6
19
1>
1C
b111 G
#530280000000
0!
0*
09
0>
0C
#530290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#530300000000
0!
0*
09
0>
0C
#530310000000
1!
1*
b1 6
19
1>
1C
b1 G
#530320000000
0!
0*
09
0>
0C
#530330000000
1!
1*
b10 6
19
1>
1C
b10 G
#530340000000
0!
0*
09
0>
0C
#530350000000
1!
1*
b11 6
19
1>
1C
b11 G
#530360000000
0!
0*
09
0>
0C
#530370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#530380000000
0!
0*
09
0>
0C
#530390000000
1!
1*
b101 6
19
1>
1C
b101 G
#530400000000
0!
0*
09
0>
0C
#530410000000
1!
1*
b110 6
19
1>
1C
b110 G
#530420000000
0!
0*
09
0>
0C
#530430000000
1!
1*
b111 6
19
1>
1C
b111 G
#530440000000
0!
1"
0*
1+
09
1:
0>
0C
#530450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#530460000000
0!
0*
09
0>
0C
#530470000000
1!
1*
b1 6
19
1>
1C
b1 G
#530480000000
0!
0*
09
0>
0C
#530490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#530500000000
0!
0*
09
0>
0C
#530510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#530520000000
0!
0*
09
0>
0C
#530530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#530540000000
0!
0*
09
0>
0C
#530550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#530560000000
0!
0#
0*
0,
09
0>
0?
0C
#530570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#530580000000
0!
0*
09
0>
0C
#530590000000
1!
1*
19
1>
1C
#530600000000
0!
0*
09
0>
0C
#530610000000
1!
1*
19
1>
1C
#530620000000
0!
0*
09
0>
0C
#530630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#530640000000
0!
0*
09
0>
0C
#530650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#530660000000
0!
0*
09
0>
0C
#530670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#530680000000
0!
0*
09
0>
0C
#530690000000
1!
1*
b10 6
19
1>
1C
b10 G
#530700000000
0!
0*
09
0>
0C
#530710000000
1!
1*
b11 6
19
1>
1C
b11 G
#530720000000
0!
0*
09
0>
0C
#530730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#530740000000
0!
0*
09
0>
0C
#530750000000
1!
1*
b101 6
19
1>
1C
b101 G
#530760000000
0!
0*
09
0>
0C
#530770000000
1!
1*
b110 6
19
1>
1C
b110 G
#530780000000
0!
0*
09
0>
0C
#530790000000
1!
1*
b111 6
19
1>
1C
b111 G
#530800000000
0!
0*
09
0>
0C
#530810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#530820000000
0!
0*
09
0>
0C
#530830000000
1!
1*
b1 6
19
1>
1C
b1 G
#530840000000
0!
0*
09
0>
0C
#530850000000
1!
1*
b10 6
19
1>
1C
b10 G
#530860000000
0!
0*
09
0>
0C
#530870000000
1!
1*
b11 6
19
1>
1C
b11 G
#530880000000
0!
0*
09
0>
0C
#530890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#530900000000
0!
0*
09
0>
0C
#530910000000
1!
1*
b101 6
19
1>
1C
b101 G
#530920000000
0!
0*
09
0>
0C
#530930000000
1!
1*
b110 6
19
1>
1C
b110 G
#530940000000
0!
0*
09
0>
0C
#530950000000
1!
1*
b111 6
19
1>
1C
b111 G
#530960000000
0!
0*
09
0>
0C
#530970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#530980000000
0!
0*
09
0>
0C
#530990000000
1!
1*
b1 6
19
1>
1C
b1 G
#531000000000
0!
0*
09
0>
0C
#531010000000
1!
1*
b10 6
19
1>
1C
b10 G
#531020000000
0!
0*
09
0>
0C
#531030000000
1!
1*
b11 6
19
1>
1C
b11 G
#531040000000
0!
0*
09
0>
0C
#531050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#531060000000
0!
0*
09
0>
0C
#531070000000
1!
1*
b101 6
19
1>
1C
b101 G
#531080000000
0!
0*
09
0>
0C
#531090000000
1!
1*
b110 6
19
1>
1C
b110 G
#531100000000
0!
0*
09
0>
0C
#531110000000
1!
1*
b111 6
19
1>
1C
b111 G
#531120000000
0!
1"
0*
1+
09
1:
0>
0C
#531130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#531140000000
0!
0*
09
0>
0C
#531150000000
1!
1*
b1 6
19
1>
1C
b1 G
#531160000000
0!
0*
09
0>
0C
#531170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#531180000000
0!
0*
09
0>
0C
#531190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#531200000000
0!
0*
09
0>
0C
#531210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#531220000000
0!
0*
09
0>
0C
#531230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#531240000000
0!
0#
0*
0,
09
0>
0?
0C
#531250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#531260000000
0!
0*
09
0>
0C
#531270000000
1!
1*
19
1>
1C
#531280000000
0!
0*
09
0>
0C
#531290000000
1!
1*
19
1>
1C
#531300000000
0!
0*
09
0>
0C
#531310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#531320000000
0!
0*
09
0>
0C
#531330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#531340000000
0!
0*
09
0>
0C
#531350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#531360000000
0!
0*
09
0>
0C
#531370000000
1!
1*
b10 6
19
1>
1C
b10 G
#531380000000
0!
0*
09
0>
0C
#531390000000
1!
1*
b11 6
19
1>
1C
b11 G
#531400000000
0!
0*
09
0>
0C
#531410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#531420000000
0!
0*
09
0>
0C
#531430000000
1!
1*
b101 6
19
1>
1C
b101 G
#531440000000
0!
0*
09
0>
0C
#531450000000
1!
1*
b110 6
19
1>
1C
b110 G
#531460000000
0!
0*
09
0>
0C
#531470000000
1!
1*
b111 6
19
1>
1C
b111 G
#531480000000
0!
0*
09
0>
0C
#531490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#531500000000
0!
0*
09
0>
0C
#531510000000
1!
1*
b1 6
19
1>
1C
b1 G
#531520000000
0!
0*
09
0>
0C
#531530000000
1!
1*
b10 6
19
1>
1C
b10 G
#531540000000
0!
0*
09
0>
0C
#531550000000
1!
1*
b11 6
19
1>
1C
b11 G
#531560000000
0!
0*
09
0>
0C
#531570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#531580000000
0!
0*
09
0>
0C
#531590000000
1!
1*
b101 6
19
1>
1C
b101 G
#531600000000
0!
0*
09
0>
0C
#531610000000
1!
1*
b110 6
19
1>
1C
b110 G
#531620000000
0!
0*
09
0>
0C
#531630000000
1!
1*
b111 6
19
1>
1C
b111 G
#531640000000
0!
0*
09
0>
0C
#531650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#531660000000
0!
0*
09
0>
0C
#531670000000
1!
1*
b1 6
19
1>
1C
b1 G
#531680000000
0!
0*
09
0>
0C
#531690000000
1!
1*
b10 6
19
1>
1C
b10 G
#531700000000
0!
0*
09
0>
0C
#531710000000
1!
1*
b11 6
19
1>
1C
b11 G
#531720000000
0!
0*
09
0>
0C
#531730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#531740000000
0!
0*
09
0>
0C
#531750000000
1!
1*
b101 6
19
1>
1C
b101 G
#531760000000
0!
0*
09
0>
0C
#531770000000
1!
1*
b110 6
19
1>
1C
b110 G
#531780000000
0!
0*
09
0>
0C
#531790000000
1!
1*
b111 6
19
1>
1C
b111 G
#531800000000
0!
1"
0*
1+
09
1:
0>
0C
#531810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#531820000000
0!
0*
09
0>
0C
#531830000000
1!
1*
b1 6
19
1>
1C
b1 G
#531840000000
0!
0*
09
0>
0C
#531850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#531860000000
0!
0*
09
0>
0C
#531870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#531880000000
0!
0*
09
0>
0C
#531890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#531900000000
0!
0*
09
0>
0C
#531910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#531920000000
0!
0#
0*
0,
09
0>
0?
0C
#531930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#531940000000
0!
0*
09
0>
0C
#531950000000
1!
1*
19
1>
1C
#531960000000
0!
0*
09
0>
0C
#531970000000
1!
1*
19
1>
1C
#531980000000
0!
0*
09
0>
0C
#531990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#532000000000
0!
0*
09
0>
0C
#532010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#532020000000
0!
0*
09
0>
0C
#532030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#532040000000
0!
0*
09
0>
0C
#532050000000
1!
1*
b10 6
19
1>
1C
b10 G
#532060000000
0!
0*
09
0>
0C
#532070000000
1!
1*
b11 6
19
1>
1C
b11 G
#532080000000
0!
0*
09
0>
0C
#532090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#532100000000
0!
0*
09
0>
0C
#532110000000
1!
1*
b101 6
19
1>
1C
b101 G
#532120000000
0!
0*
09
0>
0C
#532130000000
1!
1*
b110 6
19
1>
1C
b110 G
#532140000000
0!
0*
09
0>
0C
#532150000000
1!
1*
b111 6
19
1>
1C
b111 G
#532160000000
0!
0*
09
0>
0C
#532170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#532180000000
0!
0*
09
0>
0C
#532190000000
1!
1*
b1 6
19
1>
1C
b1 G
#532200000000
0!
0*
09
0>
0C
#532210000000
1!
1*
b10 6
19
1>
1C
b10 G
#532220000000
0!
0*
09
0>
0C
#532230000000
1!
1*
b11 6
19
1>
1C
b11 G
#532240000000
0!
0*
09
0>
0C
#532250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#532260000000
0!
0*
09
0>
0C
#532270000000
1!
1*
b101 6
19
1>
1C
b101 G
#532280000000
0!
0*
09
0>
0C
#532290000000
1!
1*
b110 6
19
1>
1C
b110 G
#532300000000
0!
0*
09
0>
0C
#532310000000
1!
1*
b111 6
19
1>
1C
b111 G
#532320000000
0!
0*
09
0>
0C
#532330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#532340000000
0!
0*
09
0>
0C
#532350000000
1!
1*
b1 6
19
1>
1C
b1 G
#532360000000
0!
0*
09
0>
0C
#532370000000
1!
1*
b10 6
19
1>
1C
b10 G
#532380000000
0!
0*
09
0>
0C
#532390000000
1!
1*
b11 6
19
1>
1C
b11 G
#532400000000
0!
0*
09
0>
0C
#532410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#532420000000
0!
0*
09
0>
0C
#532430000000
1!
1*
b101 6
19
1>
1C
b101 G
#532440000000
0!
0*
09
0>
0C
#532450000000
1!
1*
b110 6
19
1>
1C
b110 G
#532460000000
0!
0*
09
0>
0C
#532470000000
1!
1*
b111 6
19
1>
1C
b111 G
#532480000000
0!
1"
0*
1+
09
1:
0>
0C
#532490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#532500000000
0!
0*
09
0>
0C
#532510000000
1!
1*
b1 6
19
1>
1C
b1 G
#532520000000
0!
0*
09
0>
0C
#532530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#532540000000
0!
0*
09
0>
0C
#532550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#532560000000
0!
0*
09
0>
0C
#532570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#532580000000
0!
0*
09
0>
0C
#532590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#532600000000
0!
0#
0*
0,
09
0>
0?
0C
#532610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#532620000000
0!
0*
09
0>
0C
#532630000000
1!
1*
19
1>
1C
#532640000000
0!
0*
09
0>
0C
#532650000000
1!
1*
19
1>
1C
#532660000000
0!
0*
09
0>
0C
#532670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#532680000000
0!
0*
09
0>
0C
#532690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#532700000000
0!
0*
09
0>
0C
#532710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#532720000000
0!
0*
09
0>
0C
#532730000000
1!
1*
b10 6
19
1>
1C
b10 G
#532740000000
0!
0*
09
0>
0C
#532750000000
1!
1*
b11 6
19
1>
1C
b11 G
#532760000000
0!
0*
09
0>
0C
#532770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#532780000000
0!
0*
09
0>
0C
#532790000000
1!
1*
b101 6
19
1>
1C
b101 G
#532800000000
0!
0*
09
0>
0C
#532810000000
1!
1*
b110 6
19
1>
1C
b110 G
#532820000000
0!
0*
09
0>
0C
#532830000000
1!
1*
b111 6
19
1>
1C
b111 G
#532840000000
0!
0*
09
0>
0C
#532850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#532860000000
0!
0*
09
0>
0C
#532870000000
1!
1*
b1 6
19
1>
1C
b1 G
#532880000000
0!
0*
09
0>
0C
#532890000000
1!
1*
b10 6
19
1>
1C
b10 G
#532900000000
0!
0*
09
0>
0C
#532910000000
1!
1*
b11 6
19
1>
1C
b11 G
#532920000000
0!
0*
09
0>
0C
#532930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#532940000000
0!
0*
09
0>
0C
#532950000000
1!
1*
b101 6
19
1>
1C
b101 G
#532960000000
0!
0*
09
0>
0C
#532970000000
1!
1*
b110 6
19
1>
1C
b110 G
#532980000000
0!
0*
09
0>
0C
#532990000000
1!
1*
b111 6
19
1>
1C
b111 G
#533000000000
0!
0*
09
0>
0C
#533010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#533020000000
0!
0*
09
0>
0C
#533030000000
1!
1*
b1 6
19
1>
1C
b1 G
#533040000000
0!
0*
09
0>
0C
#533050000000
1!
1*
b10 6
19
1>
1C
b10 G
#533060000000
0!
0*
09
0>
0C
#533070000000
1!
1*
b11 6
19
1>
1C
b11 G
#533080000000
0!
0*
09
0>
0C
#533090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#533100000000
0!
0*
09
0>
0C
#533110000000
1!
1*
b101 6
19
1>
1C
b101 G
#533120000000
0!
0*
09
0>
0C
#533130000000
1!
1*
b110 6
19
1>
1C
b110 G
#533140000000
0!
0*
09
0>
0C
#533150000000
1!
1*
b111 6
19
1>
1C
b111 G
#533160000000
0!
1"
0*
1+
09
1:
0>
0C
#533170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#533180000000
0!
0*
09
0>
0C
#533190000000
1!
1*
b1 6
19
1>
1C
b1 G
#533200000000
0!
0*
09
0>
0C
#533210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#533220000000
0!
0*
09
0>
0C
#533230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#533240000000
0!
0*
09
0>
0C
#533250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#533260000000
0!
0*
09
0>
0C
#533270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#533280000000
0!
0#
0*
0,
09
0>
0?
0C
#533290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#533300000000
0!
0*
09
0>
0C
#533310000000
1!
1*
19
1>
1C
#533320000000
0!
0*
09
0>
0C
#533330000000
1!
1*
19
1>
1C
#533340000000
0!
0*
09
0>
0C
#533350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#533360000000
0!
0*
09
0>
0C
#533370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#533380000000
0!
0*
09
0>
0C
#533390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#533400000000
0!
0*
09
0>
0C
#533410000000
1!
1*
b10 6
19
1>
1C
b10 G
#533420000000
0!
0*
09
0>
0C
#533430000000
1!
1*
b11 6
19
1>
1C
b11 G
#533440000000
0!
0*
09
0>
0C
#533450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#533460000000
0!
0*
09
0>
0C
#533470000000
1!
1*
b101 6
19
1>
1C
b101 G
#533480000000
0!
0*
09
0>
0C
#533490000000
1!
1*
b110 6
19
1>
1C
b110 G
#533500000000
0!
0*
09
0>
0C
#533510000000
1!
1*
b111 6
19
1>
1C
b111 G
#533520000000
0!
0*
09
0>
0C
#533530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#533540000000
0!
0*
09
0>
0C
#533550000000
1!
1*
b1 6
19
1>
1C
b1 G
#533560000000
0!
0*
09
0>
0C
#533570000000
1!
1*
b10 6
19
1>
1C
b10 G
#533580000000
0!
0*
09
0>
0C
#533590000000
1!
1*
b11 6
19
1>
1C
b11 G
#533600000000
0!
0*
09
0>
0C
#533610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#533620000000
0!
0*
09
0>
0C
#533630000000
1!
1*
b101 6
19
1>
1C
b101 G
#533640000000
0!
0*
09
0>
0C
#533650000000
1!
1*
b110 6
19
1>
1C
b110 G
#533660000000
0!
0*
09
0>
0C
#533670000000
1!
1*
b111 6
19
1>
1C
b111 G
#533680000000
0!
0*
09
0>
0C
#533690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#533700000000
0!
0*
09
0>
0C
#533710000000
1!
1*
b1 6
19
1>
1C
b1 G
#533720000000
0!
0*
09
0>
0C
#533730000000
1!
1*
b10 6
19
1>
1C
b10 G
#533740000000
0!
0*
09
0>
0C
#533750000000
1!
1*
b11 6
19
1>
1C
b11 G
#533760000000
0!
0*
09
0>
0C
#533770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#533780000000
0!
0*
09
0>
0C
#533790000000
1!
1*
b101 6
19
1>
1C
b101 G
#533800000000
0!
0*
09
0>
0C
#533810000000
1!
1*
b110 6
19
1>
1C
b110 G
#533820000000
0!
0*
09
0>
0C
#533830000000
1!
1*
b111 6
19
1>
1C
b111 G
#533840000000
0!
1"
0*
1+
09
1:
0>
0C
#533850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#533860000000
0!
0*
09
0>
0C
#533870000000
1!
1*
b1 6
19
1>
1C
b1 G
#533880000000
0!
0*
09
0>
0C
#533890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#533900000000
0!
0*
09
0>
0C
#533910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#533920000000
0!
0*
09
0>
0C
#533930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#533940000000
0!
0*
09
0>
0C
#533950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#533960000000
0!
0#
0*
0,
09
0>
0?
0C
#533970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#533980000000
0!
0*
09
0>
0C
#533990000000
1!
1*
19
1>
1C
#534000000000
0!
0*
09
0>
0C
#534010000000
1!
1*
19
1>
1C
#534020000000
0!
0*
09
0>
0C
#534030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#534040000000
0!
0*
09
0>
0C
#534050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#534060000000
0!
0*
09
0>
0C
#534070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#534080000000
0!
0*
09
0>
0C
#534090000000
1!
1*
b10 6
19
1>
1C
b10 G
#534100000000
0!
0*
09
0>
0C
#534110000000
1!
1*
b11 6
19
1>
1C
b11 G
#534120000000
0!
0*
09
0>
0C
#534130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#534140000000
0!
0*
09
0>
0C
#534150000000
1!
1*
b101 6
19
1>
1C
b101 G
#534160000000
0!
0*
09
0>
0C
#534170000000
1!
1*
b110 6
19
1>
1C
b110 G
#534180000000
0!
0*
09
0>
0C
#534190000000
1!
1*
b111 6
19
1>
1C
b111 G
#534200000000
0!
0*
09
0>
0C
#534210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#534220000000
0!
0*
09
0>
0C
#534230000000
1!
1*
b1 6
19
1>
1C
b1 G
#534240000000
0!
0*
09
0>
0C
#534250000000
1!
1*
b10 6
19
1>
1C
b10 G
#534260000000
0!
0*
09
0>
0C
#534270000000
1!
1*
b11 6
19
1>
1C
b11 G
#534280000000
0!
0*
09
0>
0C
#534290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#534300000000
0!
0*
09
0>
0C
#534310000000
1!
1*
b101 6
19
1>
1C
b101 G
#534320000000
0!
0*
09
0>
0C
#534330000000
1!
1*
b110 6
19
1>
1C
b110 G
#534340000000
0!
0*
09
0>
0C
#534350000000
1!
1*
b111 6
19
1>
1C
b111 G
#534360000000
0!
0*
09
0>
0C
#534370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#534380000000
0!
0*
09
0>
0C
#534390000000
1!
1*
b1 6
19
1>
1C
b1 G
#534400000000
0!
0*
09
0>
0C
#534410000000
1!
1*
b10 6
19
1>
1C
b10 G
#534420000000
0!
0*
09
0>
0C
#534430000000
1!
1*
b11 6
19
1>
1C
b11 G
#534440000000
0!
0*
09
0>
0C
#534450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#534460000000
0!
0*
09
0>
0C
#534470000000
1!
1*
b101 6
19
1>
1C
b101 G
#534480000000
0!
0*
09
0>
0C
#534490000000
1!
1*
b110 6
19
1>
1C
b110 G
#534500000000
0!
0*
09
0>
0C
#534510000000
1!
1*
b111 6
19
1>
1C
b111 G
#534520000000
0!
1"
0*
1+
09
1:
0>
0C
#534530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#534540000000
0!
0*
09
0>
0C
#534550000000
1!
1*
b1 6
19
1>
1C
b1 G
#534560000000
0!
0*
09
0>
0C
#534570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#534580000000
0!
0*
09
0>
0C
#534590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#534600000000
0!
0*
09
0>
0C
#534610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#534620000000
0!
0*
09
0>
0C
#534630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#534640000000
0!
0#
0*
0,
09
0>
0?
0C
#534650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#534660000000
0!
0*
09
0>
0C
#534670000000
1!
1*
19
1>
1C
#534680000000
0!
0*
09
0>
0C
#534690000000
1!
1*
19
1>
1C
#534700000000
0!
0*
09
0>
0C
#534710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#534720000000
0!
0*
09
0>
0C
#534730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#534740000000
0!
0*
09
0>
0C
#534750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#534760000000
0!
0*
09
0>
0C
#534770000000
1!
1*
b10 6
19
1>
1C
b10 G
#534780000000
0!
0*
09
0>
0C
#534790000000
1!
1*
b11 6
19
1>
1C
b11 G
#534800000000
0!
0*
09
0>
0C
#534810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#534820000000
0!
0*
09
0>
0C
#534830000000
1!
1*
b101 6
19
1>
1C
b101 G
#534840000000
0!
0*
09
0>
0C
#534850000000
1!
1*
b110 6
19
1>
1C
b110 G
#534860000000
0!
0*
09
0>
0C
#534870000000
1!
1*
b111 6
19
1>
1C
b111 G
#534880000000
0!
0*
09
0>
0C
#534890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#534900000000
0!
0*
09
0>
0C
#534910000000
1!
1*
b1 6
19
1>
1C
b1 G
#534920000000
0!
0*
09
0>
0C
#534930000000
1!
1*
b10 6
19
1>
1C
b10 G
#534940000000
0!
0*
09
0>
0C
#534950000000
1!
1*
b11 6
19
1>
1C
b11 G
#534960000000
0!
0*
09
0>
0C
#534970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#534980000000
0!
0*
09
0>
0C
#534990000000
1!
1*
b101 6
19
1>
1C
b101 G
#535000000000
0!
0*
09
0>
0C
#535010000000
1!
1*
b110 6
19
1>
1C
b110 G
#535020000000
0!
0*
09
0>
0C
#535030000000
1!
1*
b111 6
19
1>
1C
b111 G
#535040000000
0!
0*
09
0>
0C
#535050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#535060000000
0!
0*
09
0>
0C
#535070000000
1!
1*
b1 6
19
1>
1C
b1 G
#535080000000
0!
0*
09
0>
0C
#535090000000
1!
1*
b10 6
19
1>
1C
b10 G
#535100000000
0!
0*
09
0>
0C
#535110000000
1!
1*
b11 6
19
1>
1C
b11 G
#535120000000
0!
0*
09
0>
0C
#535130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#535140000000
0!
0*
09
0>
0C
#535150000000
1!
1*
b101 6
19
1>
1C
b101 G
#535160000000
0!
0*
09
0>
0C
#535170000000
1!
1*
b110 6
19
1>
1C
b110 G
#535180000000
0!
0*
09
0>
0C
#535190000000
1!
1*
b111 6
19
1>
1C
b111 G
#535200000000
0!
1"
0*
1+
09
1:
0>
0C
#535210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#535220000000
0!
0*
09
0>
0C
#535230000000
1!
1*
b1 6
19
1>
1C
b1 G
#535240000000
0!
0*
09
0>
0C
#535250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#535260000000
0!
0*
09
0>
0C
#535270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#535280000000
0!
0*
09
0>
0C
#535290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#535300000000
0!
0*
09
0>
0C
#535310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#535320000000
0!
0#
0*
0,
09
0>
0?
0C
#535330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#535340000000
0!
0*
09
0>
0C
#535350000000
1!
1*
19
1>
1C
#535360000000
0!
0*
09
0>
0C
#535370000000
1!
1*
19
1>
1C
#535380000000
0!
0*
09
0>
0C
#535390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#535400000000
0!
0*
09
0>
0C
#535410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#535420000000
0!
0*
09
0>
0C
#535430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#535440000000
0!
0*
09
0>
0C
#535450000000
1!
1*
b10 6
19
1>
1C
b10 G
#535460000000
0!
0*
09
0>
0C
#535470000000
1!
1*
b11 6
19
1>
1C
b11 G
#535480000000
0!
0*
09
0>
0C
#535490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#535500000000
0!
0*
09
0>
0C
#535510000000
1!
1*
b101 6
19
1>
1C
b101 G
#535520000000
0!
0*
09
0>
0C
#535530000000
1!
1*
b110 6
19
1>
1C
b110 G
#535540000000
0!
0*
09
0>
0C
#535550000000
1!
1*
b111 6
19
1>
1C
b111 G
#535560000000
0!
0*
09
0>
0C
#535570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#535580000000
0!
0*
09
0>
0C
#535590000000
1!
1*
b1 6
19
1>
1C
b1 G
#535600000000
0!
0*
09
0>
0C
#535610000000
1!
1*
b10 6
19
1>
1C
b10 G
#535620000000
0!
0*
09
0>
0C
#535630000000
1!
1*
b11 6
19
1>
1C
b11 G
#535640000000
0!
0*
09
0>
0C
#535650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#535660000000
0!
0*
09
0>
0C
#535670000000
1!
1*
b101 6
19
1>
1C
b101 G
#535680000000
0!
0*
09
0>
0C
#535690000000
1!
1*
b110 6
19
1>
1C
b110 G
#535700000000
0!
0*
09
0>
0C
#535710000000
1!
1*
b111 6
19
1>
1C
b111 G
#535720000000
0!
0*
09
0>
0C
#535730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#535740000000
0!
0*
09
0>
0C
#535750000000
1!
1*
b1 6
19
1>
1C
b1 G
#535760000000
0!
0*
09
0>
0C
#535770000000
1!
1*
b10 6
19
1>
1C
b10 G
#535780000000
0!
0*
09
0>
0C
#535790000000
1!
1*
b11 6
19
1>
1C
b11 G
#535800000000
0!
0*
09
0>
0C
#535810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#535820000000
0!
0*
09
0>
0C
#535830000000
1!
1*
b101 6
19
1>
1C
b101 G
#535840000000
0!
0*
09
0>
0C
#535850000000
1!
1*
b110 6
19
1>
1C
b110 G
#535860000000
0!
0*
09
0>
0C
#535870000000
1!
1*
b111 6
19
1>
1C
b111 G
#535880000000
0!
1"
0*
1+
09
1:
0>
0C
#535890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#535900000000
0!
0*
09
0>
0C
#535910000000
1!
1*
b1 6
19
1>
1C
b1 G
#535920000000
0!
0*
09
0>
0C
#535930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#535940000000
0!
0*
09
0>
0C
#535950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#535960000000
0!
0*
09
0>
0C
#535970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#535980000000
0!
0*
09
0>
0C
#535990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#536000000000
0!
0#
0*
0,
09
0>
0?
0C
#536010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#536020000000
0!
0*
09
0>
0C
#536030000000
1!
1*
19
1>
1C
#536040000000
0!
0*
09
0>
0C
#536050000000
1!
1*
19
1>
1C
#536060000000
0!
0*
09
0>
0C
#536070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#536080000000
0!
0*
09
0>
0C
#536090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#536100000000
0!
0*
09
0>
0C
#536110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#536120000000
0!
0*
09
0>
0C
#536130000000
1!
1*
b10 6
19
1>
1C
b10 G
#536140000000
0!
0*
09
0>
0C
#536150000000
1!
1*
b11 6
19
1>
1C
b11 G
#536160000000
0!
0*
09
0>
0C
#536170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#536180000000
0!
0*
09
0>
0C
#536190000000
1!
1*
b101 6
19
1>
1C
b101 G
#536200000000
0!
0*
09
0>
0C
#536210000000
1!
1*
b110 6
19
1>
1C
b110 G
#536220000000
0!
0*
09
0>
0C
#536230000000
1!
1*
b111 6
19
1>
1C
b111 G
#536240000000
0!
0*
09
0>
0C
#536250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#536260000000
0!
0*
09
0>
0C
#536270000000
1!
1*
b1 6
19
1>
1C
b1 G
#536280000000
0!
0*
09
0>
0C
#536290000000
1!
1*
b10 6
19
1>
1C
b10 G
#536300000000
0!
0*
09
0>
0C
#536310000000
1!
1*
b11 6
19
1>
1C
b11 G
#536320000000
0!
0*
09
0>
0C
#536330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#536340000000
0!
0*
09
0>
0C
#536350000000
1!
1*
b101 6
19
1>
1C
b101 G
#536360000000
0!
0*
09
0>
0C
#536370000000
1!
1*
b110 6
19
1>
1C
b110 G
#536380000000
0!
0*
09
0>
0C
#536390000000
1!
1*
b111 6
19
1>
1C
b111 G
#536400000000
0!
0*
09
0>
0C
#536410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#536420000000
0!
0*
09
0>
0C
#536430000000
1!
1*
b1 6
19
1>
1C
b1 G
#536440000000
0!
0*
09
0>
0C
#536450000000
1!
1*
b10 6
19
1>
1C
b10 G
#536460000000
0!
0*
09
0>
0C
#536470000000
1!
1*
b11 6
19
1>
1C
b11 G
#536480000000
0!
0*
09
0>
0C
#536490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#536500000000
0!
0*
09
0>
0C
#536510000000
1!
1*
b101 6
19
1>
1C
b101 G
#536520000000
0!
0*
09
0>
0C
#536530000000
1!
1*
b110 6
19
1>
1C
b110 G
#536540000000
0!
0*
09
0>
0C
#536550000000
1!
1*
b111 6
19
1>
1C
b111 G
#536560000000
0!
1"
0*
1+
09
1:
0>
0C
#536570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#536580000000
0!
0*
09
0>
0C
#536590000000
1!
1*
b1 6
19
1>
1C
b1 G
#536600000000
0!
0*
09
0>
0C
#536610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#536620000000
0!
0*
09
0>
0C
#536630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#536640000000
0!
0*
09
0>
0C
#536650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#536660000000
0!
0*
09
0>
0C
#536670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#536680000000
0!
0#
0*
0,
09
0>
0?
0C
#536690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#536700000000
0!
0*
09
0>
0C
#536710000000
1!
1*
19
1>
1C
#536720000000
0!
0*
09
0>
0C
#536730000000
1!
1*
19
1>
1C
#536740000000
0!
0*
09
0>
0C
#536750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#536760000000
0!
0*
09
0>
0C
#536770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#536780000000
0!
0*
09
0>
0C
#536790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#536800000000
0!
0*
09
0>
0C
#536810000000
1!
1*
b10 6
19
1>
1C
b10 G
#536820000000
0!
0*
09
0>
0C
#536830000000
1!
1*
b11 6
19
1>
1C
b11 G
#536840000000
0!
0*
09
0>
0C
#536850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#536860000000
0!
0*
09
0>
0C
#536870000000
1!
1*
b101 6
19
1>
1C
b101 G
#536880000000
0!
0*
09
0>
0C
#536890000000
1!
1*
b110 6
19
1>
1C
b110 G
#536900000000
0!
0*
09
0>
0C
#536910000000
1!
1*
b111 6
19
1>
1C
b111 G
#536920000000
0!
0*
09
0>
0C
#536930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#536940000000
0!
0*
09
0>
0C
#536950000000
1!
1*
b1 6
19
1>
1C
b1 G
#536960000000
0!
0*
09
0>
0C
#536970000000
1!
1*
b10 6
19
1>
1C
b10 G
#536980000000
0!
0*
09
0>
0C
#536990000000
1!
1*
b11 6
19
1>
1C
b11 G
#537000000000
0!
0*
09
0>
0C
#537010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#537020000000
0!
0*
09
0>
0C
#537030000000
1!
1*
b101 6
19
1>
1C
b101 G
#537040000000
0!
0*
09
0>
0C
#537050000000
1!
1*
b110 6
19
1>
1C
b110 G
#537060000000
0!
0*
09
0>
0C
#537070000000
1!
1*
b111 6
19
1>
1C
b111 G
#537080000000
0!
0*
09
0>
0C
#537090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#537100000000
0!
0*
09
0>
0C
#537110000000
1!
1*
b1 6
19
1>
1C
b1 G
#537120000000
0!
0*
09
0>
0C
#537130000000
1!
1*
b10 6
19
1>
1C
b10 G
#537140000000
0!
0*
09
0>
0C
#537150000000
1!
1*
b11 6
19
1>
1C
b11 G
#537160000000
0!
0*
09
0>
0C
#537170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#537180000000
0!
0*
09
0>
0C
#537190000000
1!
1*
b101 6
19
1>
1C
b101 G
#537200000000
0!
0*
09
0>
0C
#537210000000
1!
1*
b110 6
19
1>
1C
b110 G
#537220000000
0!
0*
09
0>
0C
#537230000000
1!
1*
b111 6
19
1>
1C
b111 G
#537240000000
0!
1"
0*
1+
09
1:
0>
0C
#537250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#537260000000
0!
0*
09
0>
0C
#537270000000
1!
1*
b1 6
19
1>
1C
b1 G
#537280000000
0!
0*
09
0>
0C
#537290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#537300000000
0!
0*
09
0>
0C
#537310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#537320000000
0!
0*
09
0>
0C
#537330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#537340000000
0!
0*
09
0>
0C
#537350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#537360000000
0!
0#
0*
0,
09
0>
0?
0C
#537370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#537380000000
0!
0*
09
0>
0C
#537390000000
1!
1*
19
1>
1C
#537400000000
0!
0*
09
0>
0C
#537410000000
1!
1*
19
1>
1C
#537420000000
0!
0*
09
0>
0C
#537430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#537440000000
0!
0*
09
0>
0C
#537450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#537460000000
0!
0*
09
0>
0C
#537470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#537480000000
0!
0*
09
0>
0C
#537490000000
1!
1*
b10 6
19
1>
1C
b10 G
#537500000000
0!
0*
09
0>
0C
#537510000000
1!
1*
b11 6
19
1>
1C
b11 G
#537520000000
0!
0*
09
0>
0C
#537530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#537540000000
0!
0*
09
0>
0C
#537550000000
1!
1*
b101 6
19
1>
1C
b101 G
#537560000000
0!
0*
09
0>
0C
#537570000000
1!
1*
b110 6
19
1>
1C
b110 G
#537580000000
0!
0*
09
0>
0C
#537590000000
1!
1*
b111 6
19
1>
1C
b111 G
#537600000000
0!
0*
09
0>
0C
#537610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#537620000000
0!
0*
09
0>
0C
#537630000000
1!
1*
b1 6
19
1>
1C
b1 G
#537640000000
0!
0*
09
0>
0C
#537650000000
1!
1*
b10 6
19
1>
1C
b10 G
#537660000000
0!
0*
09
0>
0C
#537670000000
1!
1*
b11 6
19
1>
1C
b11 G
#537680000000
0!
0*
09
0>
0C
#537690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#537700000000
0!
0*
09
0>
0C
#537710000000
1!
1*
b101 6
19
1>
1C
b101 G
#537720000000
0!
0*
09
0>
0C
#537730000000
1!
1*
b110 6
19
1>
1C
b110 G
#537740000000
0!
0*
09
0>
0C
#537750000000
1!
1*
b111 6
19
1>
1C
b111 G
#537760000000
0!
0*
09
0>
0C
#537770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#537780000000
0!
0*
09
0>
0C
#537790000000
1!
1*
b1 6
19
1>
1C
b1 G
#537800000000
0!
0*
09
0>
0C
#537810000000
1!
1*
b10 6
19
1>
1C
b10 G
#537820000000
0!
0*
09
0>
0C
#537830000000
1!
1*
b11 6
19
1>
1C
b11 G
#537840000000
0!
0*
09
0>
0C
#537850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#537860000000
0!
0*
09
0>
0C
#537870000000
1!
1*
b101 6
19
1>
1C
b101 G
#537880000000
0!
0*
09
0>
0C
#537890000000
1!
1*
b110 6
19
1>
1C
b110 G
#537900000000
0!
0*
09
0>
0C
#537910000000
1!
1*
b111 6
19
1>
1C
b111 G
#537920000000
0!
1"
0*
1+
09
1:
0>
0C
#537930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#537940000000
0!
0*
09
0>
0C
#537950000000
1!
1*
b1 6
19
1>
1C
b1 G
#537960000000
0!
0*
09
0>
0C
#537970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#537980000000
0!
0*
09
0>
0C
#537990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#538000000000
0!
0*
09
0>
0C
#538010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#538020000000
0!
0*
09
0>
0C
#538030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#538040000000
0!
0#
0*
0,
09
0>
0?
0C
#538050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#538060000000
0!
0*
09
0>
0C
#538070000000
1!
1*
19
1>
1C
#538080000000
0!
0*
09
0>
0C
#538090000000
1!
1*
19
1>
1C
#538100000000
0!
0*
09
0>
0C
#538110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#538120000000
0!
0*
09
0>
0C
#538130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#538140000000
0!
0*
09
0>
0C
#538150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#538160000000
0!
0*
09
0>
0C
#538170000000
1!
1*
b10 6
19
1>
1C
b10 G
#538180000000
0!
0*
09
0>
0C
#538190000000
1!
1*
b11 6
19
1>
1C
b11 G
#538200000000
0!
0*
09
0>
0C
#538210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#538220000000
0!
0*
09
0>
0C
#538230000000
1!
1*
b101 6
19
1>
1C
b101 G
#538240000000
0!
0*
09
0>
0C
#538250000000
1!
1*
b110 6
19
1>
1C
b110 G
#538260000000
0!
0*
09
0>
0C
#538270000000
1!
1*
b111 6
19
1>
1C
b111 G
#538280000000
0!
0*
09
0>
0C
#538290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#538300000000
0!
0*
09
0>
0C
#538310000000
1!
1*
b1 6
19
1>
1C
b1 G
#538320000000
0!
0*
09
0>
0C
#538330000000
1!
1*
b10 6
19
1>
1C
b10 G
#538340000000
0!
0*
09
0>
0C
#538350000000
1!
1*
b11 6
19
1>
1C
b11 G
#538360000000
0!
0*
09
0>
0C
#538370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#538380000000
0!
0*
09
0>
0C
#538390000000
1!
1*
b101 6
19
1>
1C
b101 G
#538400000000
0!
0*
09
0>
0C
#538410000000
1!
1*
b110 6
19
1>
1C
b110 G
#538420000000
0!
0*
09
0>
0C
#538430000000
1!
1*
b111 6
19
1>
1C
b111 G
#538440000000
0!
0*
09
0>
0C
#538450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#538460000000
0!
0*
09
0>
0C
#538470000000
1!
1*
b1 6
19
1>
1C
b1 G
#538480000000
0!
0*
09
0>
0C
#538490000000
1!
1*
b10 6
19
1>
1C
b10 G
#538500000000
0!
0*
09
0>
0C
#538510000000
1!
1*
b11 6
19
1>
1C
b11 G
#538520000000
0!
0*
09
0>
0C
#538530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#538540000000
0!
0*
09
0>
0C
#538550000000
1!
1*
b101 6
19
1>
1C
b101 G
#538560000000
0!
0*
09
0>
0C
#538570000000
1!
1*
b110 6
19
1>
1C
b110 G
#538580000000
0!
0*
09
0>
0C
#538590000000
1!
1*
b111 6
19
1>
1C
b111 G
#538600000000
0!
1"
0*
1+
09
1:
0>
0C
#538610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#538620000000
0!
0*
09
0>
0C
#538630000000
1!
1*
b1 6
19
1>
1C
b1 G
#538640000000
0!
0*
09
0>
0C
#538650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#538660000000
0!
0*
09
0>
0C
#538670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#538680000000
0!
0*
09
0>
0C
#538690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#538700000000
0!
0*
09
0>
0C
#538710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#538720000000
0!
0#
0*
0,
09
0>
0?
0C
#538730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#538740000000
0!
0*
09
0>
0C
#538750000000
1!
1*
19
1>
1C
#538760000000
0!
0*
09
0>
0C
#538770000000
1!
1*
19
1>
1C
#538780000000
0!
0*
09
0>
0C
#538790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#538800000000
0!
0*
09
0>
0C
#538810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#538820000000
0!
0*
09
0>
0C
#538830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#538840000000
0!
0*
09
0>
0C
#538850000000
1!
1*
b10 6
19
1>
1C
b10 G
#538860000000
0!
0*
09
0>
0C
#538870000000
1!
1*
b11 6
19
1>
1C
b11 G
#538880000000
0!
0*
09
0>
0C
#538890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#538900000000
0!
0*
09
0>
0C
#538910000000
1!
1*
b101 6
19
1>
1C
b101 G
#538920000000
0!
0*
09
0>
0C
#538930000000
1!
1*
b110 6
19
1>
1C
b110 G
#538940000000
0!
0*
09
0>
0C
#538950000000
1!
1*
b111 6
19
1>
1C
b111 G
#538960000000
0!
0*
09
0>
0C
#538970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#538980000000
0!
0*
09
0>
0C
#538990000000
1!
1*
b1 6
19
1>
1C
b1 G
#539000000000
0!
0*
09
0>
0C
#539010000000
1!
1*
b10 6
19
1>
1C
b10 G
#539020000000
0!
0*
09
0>
0C
#539030000000
1!
1*
b11 6
19
1>
1C
b11 G
#539040000000
0!
0*
09
0>
0C
#539050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#539060000000
0!
0*
09
0>
0C
#539070000000
1!
1*
b101 6
19
1>
1C
b101 G
#539080000000
0!
0*
09
0>
0C
#539090000000
1!
1*
b110 6
19
1>
1C
b110 G
#539100000000
0!
0*
09
0>
0C
#539110000000
1!
1*
b111 6
19
1>
1C
b111 G
#539120000000
0!
0*
09
0>
0C
#539130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#539140000000
0!
0*
09
0>
0C
#539150000000
1!
1*
b1 6
19
1>
1C
b1 G
#539160000000
0!
0*
09
0>
0C
#539170000000
1!
1*
b10 6
19
1>
1C
b10 G
#539180000000
0!
0*
09
0>
0C
#539190000000
1!
1*
b11 6
19
1>
1C
b11 G
#539200000000
0!
0*
09
0>
0C
#539210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#539220000000
0!
0*
09
0>
0C
#539230000000
1!
1*
b101 6
19
1>
1C
b101 G
#539240000000
0!
0*
09
0>
0C
#539250000000
1!
1*
b110 6
19
1>
1C
b110 G
#539260000000
0!
0*
09
0>
0C
#539270000000
1!
1*
b111 6
19
1>
1C
b111 G
#539280000000
0!
1"
0*
1+
09
1:
0>
0C
#539290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#539300000000
0!
0*
09
0>
0C
#539310000000
1!
1*
b1 6
19
1>
1C
b1 G
#539320000000
0!
0*
09
0>
0C
#539330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#539340000000
0!
0*
09
0>
0C
#539350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#539360000000
0!
0*
09
0>
0C
#539370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#539380000000
0!
0*
09
0>
0C
#539390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#539400000000
0!
0#
0*
0,
09
0>
0?
0C
#539410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#539420000000
0!
0*
09
0>
0C
#539430000000
1!
1*
19
1>
1C
#539440000000
0!
0*
09
0>
0C
#539450000000
1!
1*
19
1>
1C
#539460000000
0!
0*
09
0>
0C
#539470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#539480000000
0!
0*
09
0>
0C
#539490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#539500000000
0!
0*
09
0>
0C
#539510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#539520000000
0!
0*
09
0>
0C
#539530000000
1!
1*
b10 6
19
1>
1C
b10 G
#539540000000
0!
0*
09
0>
0C
#539550000000
1!
1*
b11 6
19
1>
1C
b11 G
#539560000000
0!
0*
09
0>
0C
#539570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#539580000000
0!
0*
09
0>
0C
#539590000000
1!
1*
b101 6
19
1>
1C
b101 G
#539600000000
0!
0*
09
0>
0C
#539610000000
1!
1*
b110 6
19
1>
1C
b110 G
#539620000000
0!
0*
09
0>
0C
#539630000000
1!
1*
b111 6
19
1>
1C
b111 G
#539640000000
0!
0*
09
0>
0C
#539650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#539660000000
0!
0*
09
0>
0C
#539670000000
1!
1*
b1 6
19
1>
1C
b1 G
#539680000000
0!
0*
09
0>
0C
#539690000000
1!
1*
b10 6
19
1>
1C
b10 G
#539700000000
0!
0*
09
0>
0C
#539710000000
1!
1*
b11 6
19
1>
1C
b11 G
#539720000000
0!
0*
09
0>
0C
#539730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#539740000000
0!
0*
09
0>
0C
#539750000000
1!
1*
b101 6
19
1>
1C
b101 G
#539760000000
0!
0*
09
0>
0C
#539770000000
1!
1*
b110 6
19
1>
1C
b110 G
#539780000000
0!
0*
09
0>
0C
#539790000000
1!
1*
b111 6
19
1>
1C
b111 G
#539800000000
0!
0*
09
0>
0C
#539810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#539820000000
0!
0*
09
0>
0C
#539830000000
1!
1*
b1 6
19
1>
1C
b1 G
#539840000000
0!
0*
09
0>
0C
#539850000000
1!
1*
b10 6
19
1>
1C
b10 G
#539860000000
0!
0*
09
0>
0C
#539870000000
1!
1*
b11 6
19
1>
1C
b11 G
#539880000000
0!
0*
09
0>
0C
#539890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#539900000000
0!
0*
09
0>
0C
#539910000000
1!
1*
b101 6
19
1>
1C
b101 G
#539920000000
0!
0*
09
0>
0C
#539930000000
1!
1*
b110 6
19
1>
1C
b110 G
#539940000000
0!
0*
09
0>
0C
#539950000000
1!
1*
b111 6
19
1>
1C
b111 G
#539960000000
0!
1"
0*
1+
09
1:
0>
0C
#539970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#539980000000
0!
0*
09
0>
0C
#539990000000
1!
1*
b1 6
19
1>
1C
b1 G
#540000000000
0!
0*
09
0>
0C
#540010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#540020000000
0!
0*
09
0>
0C
#540030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#540040000000
0!
0*
09
0>
0C
#540050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#540060000000
0!
0*
09
0>
0C
#540070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#540080000000
0!
0#
0*
0,
09
0>
0?
0C
#540090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#540100000000
0!
0*
09
0>
0C
#540110000000
1!
1*
19
1>
1C
#540120000000
0!
0*
09
0>
0C
#540130000000
1!
1*
19
1>
1C
#540140000000
0!
0*
09
0>
0C
#540150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#540160000000
0!
0*
09
0>
0C
#540170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#540180000000
0!
0*
09
0>
0C
#540190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#540200000000
0!
0*
09
0>
0C
#540210000000
1!
1*
b10 6
19
1>
1C
b10 G
#540220000000
0!
0*
09
0>
0C
#540230000000
1!
1*
b11 6
19
1>
1C
b11 G
#540240000000
0!
0*
09
0>
0C
#540250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#540260000000
0!
0*
09
0>
0C
#540270000000
1!
1*
b101 6
19
1>
1C
b101 G
#540280000000
0!
0*
09
0>
0C
#540290000000
1!
1*
b110 6
19
1>
1C
b110 G
#540300000000
0!
0*
09
0>
0C
#540310000000
1!
1*
b111 6
19
1>
1C
b111 G
#540320000000
0!
0*
09
0>
0C
#540330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#540340000000
0!
0*
09
0>
0C
#540350000000
1!
1*
b1 6
19
1>
1C
b1 G
#540360000000
0!
0*
09
0>
0C
#540370000000
1!
1*
b10 6
19
1>
1C
b10 G
#540380000000
0!
0*
09
0>
0C
#540390000000
1!
1*
b11 6
19
1>
1C
b11 G
#540400000000
0!
0*
09
0>
0C
#540410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#540420000000
0!
0*
09
0>
0C
#540430000000
1!
1*
b101 6
19
1>
1C
b101 G
#540440000000
0!
0*
09
0>
0C
#540450000000
1!
1*
b110 6
19
1>
1C
b110 G
#540460000000
0!
0*
09
0>
0C
#540470000000
1!
1*
b111 6
19
1>
1C
b111 G
#540480000000
0!
0*
09
0>
0C
#540490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#540500000000
0!
0*
09
0>
0C
#540510000000
1!
1*
b1 6
19
1>
1C
b1 G
#540520000000
0!
0*
09
0>
0C
#540530000000
1!
1*
b10 6
19
1>
1C
b10 G
#540540000000
0!
0*
09
0>
0C
#540550000000
1!
1*
b11 6
19
1>
1C
b11 G
#540560000000
0!
0*
09
0>
0C
#540570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#540580000000
0!
0*
09
0>
0C
#540590000000
1!
1*
b101 6
19
1>
1C
b101 G
#540600000000
0!
0*
09
0>
0C
#540610000000
1!
1*
b110 6
19
1>
1C
b110 G
#540620000000
0!
0*
09
0>
0C
#540630000000
1!
1*
b111 6
19
1>
1C
b111 G
#540640000000
0!
1"
0*
1+
09
1:
0>
0C
#540650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#540660000000
0!
0*
09
0>
0C
#540670000000
1!
1*
b1 6
19
1>
1C
b1 G
#540680000000
0!
0*
09
0>
0C
#540690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#540700000000
0!
0*
09
0>
0C
#540710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#540720000000
0!
0*
09
0>
0C
#540730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#540740000000
0!
0*
09
0>
0C
#540750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#540760000000
0!
0#
0*
0,
09
0>
0?
0C
#540770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#540780000000
0!
0*
09
0>
0C
#540790000000
1!
1*
19
1>
1C
#540800000000
0!
0*
09
0>
0C
#540810000000
1!
1*
19
1>
1C
#540820000000
0!
0*
09
0>
0C
#540830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#540840000000
0!
0*
09
0>
0C
#540850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#540860000000
0!
0*
09
0>
0C
#540870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#540880000000
0!
0*
09
0>
0C
#540890000000
1!
1*
b10 6
19
1>
1C
b10 G
#540900000000
0!
0*
09
0>
0C
#540910000000
1!
1*
b11 6
19
1>
1C
b11 G
#540920000000
0!
0*
09
0>
0C
#540930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#540940000000
0!
0*
09
0>
0C
#540950000000
1!
1*
b101 6
19
1>
1C
b101 G
#540960000000
0!
0*
09
0>
0C
#540970000000
1!
1*
b110 6
19
1>
1C
b110 G
#540980000000
0!
0*
09
0>
0C
#540990000000
1!
1*
b111 6
19
1>
1C
b111 G
#541000000000
0!
0*
09
0>
0C
#541010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#541020000000
0!
0*
09
0>
0C
#541030000000
1!
1*
b1 6
19
1>
1C
b1 G
#541040000000
0!
0*
09
0>
0C
#541050000000
1!
1*
b10 6
19
1>
1C
b10 G
#541060000000
0!
0*
09
0>
0C
#541070000000
1!
1*
b11 6
19
1>
1C
b11 G
#541080000000
0!
0*
09
0>
0C
#541090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#541100000000
0!
0*
09
0>
0C
#541110000000
1!
1*
b101 6
19
1>
1C
b101 G
#541120000000
0!
0*
09
0>
0C
#541130000000
1!
1*
b110 6
19
1>
1C
b110 G
#541140000000
0!
0*
09
0>
0C
#541150000000
1!
1*
b111 6
19
1>
1C
b111 G
#541160000000
0!
0*
09
0>
0C
#541170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#541180000000
0!
0*
09
0>
0C
#541190000000
1!
1*
b1 6
19
1>
1C
b1 G
#541200000000
0!
0*
09
0>
0C
#541210000000
1!
1*
b10 6
19
1>
1C
b10 G
#541220000000
0!
0*
09
0>
0C
#541230000000
1!
1*
b11 6
19
1>
1C
b11 G
#541240000000
0!
0*
09
0>
0C
#541250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#541260000000
0!
0*
09
0>
0C
#541270000000
1!
1*
b101 6
19
1>
1C
b101 G
#541280000000
0!
0*
09
0>
0C
#541290000000
1!
1*
b110 6
19
1>
1C
b110 G
#541300000000
0!
0*
09
0>
0C
#541310000000
1!
1*
b111 6
19
1>
1C
b111 G
#541320000000
0!
1"
0*
1+
09
1:
0>
0C
#541330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#541340000000
0!
0*
09
0>
0C
#541350000000
1!
1*
b1 6
19
1>
1C
b1 G
#541360000000
0!
0*
09
0>
0C
#541370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#541380000000
0!
0*
09
0>
0C
#541390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#541400000000
0!
0*
09
0>
0C
#541410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#541420000000
0!
0*
09
0>
0C
#541430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#541440000000
0!
0#
0*
0,
09
0>
0?
0C
#541450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#541460000000
0!
0*
09
0>
0C
#541470000000
1!
1*
19
1>
1C
#541480000000
0!
0*
09
0>
0C
#541490000000
1!
1*
19
1>
1C
#541500000000
0!
0*
09
0>
0C
#541510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#541520000000
0!
0*
09
0>
0C
#541530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#541540000000
0!
0*
09
0>
0C
#541550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#541560000000
0!
0*
09
0>
0C
#541570000000
1!
1*
b10 6
19
1>
1C
b10 G
#541580000000
0!
0*
09
0>
0C
#541590000000
1!
1*
b11 6
19
1>
1C
b11 G
#541600000000
0!
0*
09
0>
0C
#541610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#541620000000
0!
0*
09
0>
0C
#541630000000
1!
1*
b101 6
19
1>
1C
b101 G
#541640000000
0!
0*
09
0>
0C
#541650000000
1!
1*
b110 6
19
1>
1C
b110 G
#541660000000
0!
0*
09
0>
0C
#541670000000
1!
1*
b111 6
19
1>
1C
b111 G
#541680000000
0!
0*
09
0>
0C
#541690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#541700000000
0!
0*
09
0>
0C
#541710000000
1!
1*
b1 6
19
1>
1C
b1 G
#541720000000
0!
0*
09
0>
0C
#541730000000
1!
1*
b10 6
19
1>
1C
b10 G
#541740000000
0!
0*
09
0>
0C
#541750000000
1!
1*
b11 6
19
1>
1C
b11 G
#541760000000
0!
0*
09
0>
0C
#541770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#541780000000
0!
0*
09
0>
0C
#541790000000
1!
1*
b101 6
19
1>
1C
b101 G
#541800000000
0!
0*
09
0>
0C
#541810000000
1!
1*
b110 6
19
1>
1C
b110 G
#541820000000
0!
0*
09
0>
0C
#541830000000
1!
1*
b111 6
19
1>
1C
b111 G
#541840000000
0!
0*
09
0>
0C
#541850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#541860000000
0!
0*
09
0>
0C
#541870000000
1!
1*
b1 6
19
1>
1C
b1 G
#541880000000
0!
0*
09
0>
0C
#541890000000
1!
1*
b10 6
19
1>
1C
b10 G
#541900000000
0!
0*
09
0>
0C
#541910000000
1!
1*
b11 6
19
1>
1C
b11 G
#541920000000
0!
0*
09
0>
0C
#541930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#541940000000
0!
0*
09
0>
0C
#541950000000
1!
1*
b101 6
19
1>
1C
b101 G
#541960000000
0!
0*
09
0>
0C
#541970000000
1!
1*
b110 6
19
1>
1C
b110 G
#541980000000
0!
0*
09
0>
0C
#541990000000
1!
1*
b111 6
19
1>
1C
b111 G
#542000000000
0!
1"
0*
1+
09
1:
0>
0C
#542010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#542020000000
0!
0*
09
0>
0C
#542030000000
1!
1*
b1 6
19
1>
1C
b1 G
#542040000000
0!
0*
09
0>
0C
#542050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#542060000000
0!
0*
09
0>
0C
#542070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#542080000000
0!
0*
09
0>
0C
#542090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#542100000000
0!
0*
09
0>
0C
#542110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#542120000000
0!
0#
0*
0,
09
0>
0?
0C
#542130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#542140000000
0!
0*
09
0>
0C
#542150000000
1!
1*
19
1>
1C
#542160000000
0!
0*
09
0>
0C
#542170000000
1!
1*
19
1>
1C
#542180000000
0!
0*
09
0>
0C
#542190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#542200000000
0!
0*
09
0>
0C
#542210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#542220000000
0!
0*
09
0>
0C
#542230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#542240000000
0!
0*
09
0>
0C
#542250000000
1!
1*
b10 6
19
1>
1C
b10 G
#542260000000
0!
0*
09
0>
0C
#542270000000
1!
1*
b11 6
19
1>
1C
b11 G
#542280000000
0!
0*
09
0>
0C
#542290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#542300000000
0!
0*
09
0>
0C
#542310000000
1!
1*
b101 6
19
1>
1C
b101 G
#542320000000
0!
0*
09
0>
0C
#542330000000
1!
1*
b110 6
19
1>
1C
b110 G
#542340000000
0!
0*
09
0>
0C
#542350000000
1!
1*
b111 6
19
1>
1C
b111 G
#542360000000
0!
0*
09
0>
0C
#542370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#542380000000
0!
0*
09
0>
0C
#542390000000
1!
1*
b1 6
19
1>
1C
b1 G
#542400000000
0!
0*
09
0>
0C
#542410000000
1!
1*
b10 6
19
1>
1C
b10 G
#542420000000
0!
0*
09
0>
0C
#542430000000
1!
1*
b11 6
19
1>
1C
b11 G
#542440000000
0!
0*
09
0>
0C
#542450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#542460000000
0!
0*
09
0>
0C
#542470000000
1!
1*
b101 6
19
1>
1C
b101 G
#542480000000
0!
0*
09
0>
0C
#542490000000
1!
1*
b110 6
19
1>
1C
b110 G
#542500000000
0!
0*
09
0>
0C
#542510000000
1!
1*
b111 6
19
1>
1C
b111 G
#542520000000
0!
0*
09
0>
0C
#542530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#542540000000
0!
0*
09
0>
0C
#542550000000
1!
1*
b1 6
19
1>
1C
b1 G
#542560000000
0!
0*
09
0>
0C
#542570000000
1!
1*
b10 6
19
1>
1C
b10 G
#542580000000
0!
0*
09
0>
0C
#542590000000
1!
1*
b11 6
19
1>
1C
b11 G
#542600000000
0!
0*
09
0>
0C
#542610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#542620000000
0!
0*
09
0>
0C
#542630000000
1!
1*
b101 6
19
1>
1C
b101 G
#542640000000
0!
0*
09
0>
0C
#542650000000
1!
1*
b110 6
19
1>
1C
b110 G
#542660000000
0!
0*
09
0>
0C
#542670000000
1!
1*
b111 6
19
1>
1C
b111 G
#542680000000
0!
1"
0*
1+
09
1:
0>
0C
#542690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#542700000000
0!
0*
09
0>
0C
#542710000000
1!
1*
b1 6
19
1>
1C
b1 G
#542720000000
0!
0*
09
0>
0C
#542730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#542740000000
0!
0*
09
0>
0C
#542750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#542760000000
0!
0*
09
0>
0C
#542770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#542780000000
0!
0*
09
0>
0C
#542790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#542800000000
0!
0#
0*
0,
09
0>
0?
0C
#542810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#542820000000
0!
0*
09
0>
0C
#542830000000
1!
1*
19
1>
1C
#542840000000
0!
0*
09
0>
0C
#542850000000
1!
1*
19
1>
1C
#542860000000
0!
0*
09
0>
0C
#542870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#542880000000
0!
0*
09
0>
0C
#542890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#542900000000
0!
0*
09
0>
0C
#542910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#542920000000
0!
0*
09
0>
0C
#542930000000
1!
1*
b10 6
19
1>
1C
b10 G
#542940000000
0!
0*
09
0>
0C
#542950000000
1!
1*
b11 6
19
1>
1C
b11 G
#542960000000
0!
0*
09
0>
0C
#542970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#542980000000
0!
0*
09
0>
0C
#542990000000
1!
1*
b101 6
19
1>
1C
b101 G
#543000000000
0!
0*
09
0>
0C
#543010000000
1!
1*
b110 6
19
1>
1C
b110 G
#543020000000
0!
0*
09
0>
0C
#543030000000
1!
1*
b111 6
19
1>
1C
b111 G
#543040000000
0!
0*
09
0>
0C
#543050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#543060000000
0!
0*
09
0>
0C
#543070000000
1!
1*
b1 6
19
1>
1C
b1 G
#543080000000
0!
0*
09
0>
0C
#543090000000
1!
1*
b10 6
19
1>
1C
b10 G
#543100000000
0!
0*
09
0>
0C
#543110000000
1!
1*
b11 6
19
1>
1C
b11 G
#543120000000
0!
0*
09
0>
0C
#543130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#543140000000
0!
0*
09
0>
0C
#543150000000
1!
1*
b101 6
19
1>
1C
b101 G
#543160000000
0!
0*
09
0>
0C
#543170000000
1!
1*
b110 6
19
1>
1C
b110 G
#543180000000
0!
0*
09
0>
0C
#543190000000
1!
1*
b111 6
19
1>
1C
b111 G
#543200000000
0!
0*
09
0>
0C
#543210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#543220000000
0!
0*
09
0>
0C
#543230000000
1!
1*
b1 6
19
1>
1C
b1 G
#543240000000
0!
0*
09
0>
0C
#543250000000
1!
1*
b10 6
19
1>
1C
b10 G
#543260000000
0!
0*
09
0>
0C
#543270000000
1!
1*
b11 6
19
1>
1C
b11 G
#543280000000
0!
0*
09
0>
0C
#543290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#543300000000
0!
0*
09
0>
0C
#543310000000
1!
1*
b101 6
19
1>
1C
b101 G
#543320000000
0!
0*
09
0>
0C
#543330000000
1!
1*
b110 6
19
1>
1C
b110 G
#543340000000
0!
0*
09
0>
0C
#543350000000
1!
1*
b111 6
19
1>
1C
b111 G
#543360000000
0!
1"
0*
1+
09
1:
0>
0C
#543370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#543380000000
0!
0*
09
0>
0C
#543390000000
1!
1*
b1 6
19
1>
1C
b1 G
#543400000000
0!
0*
09
0>
0C
#543410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#543420000000
0!
0*
09
0>
0C
#543430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#543440000000
0!
0*
09
0>
0C
#543450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#543460000000
0!
0*
09
0>
0C
#543470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#543480000000
0!
0#
0*
0,
09
0>
0?
0C
#543490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#543500000000
0!
0*
09
0>
0C
#543510000000
1!
1*
19
1>
1C
#543520000000
0!
0*
09
0>
0C
#543530000000
1!
1*
19
1>
1C
#543540000000
0!
0*
09
0>
0C
#543550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#543560000000
0!
0*
09
0>
0C
#543570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#543580000000
0!
0*
09
0>
0C
#543590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#543600000000
0!
0*
09
0>
0C
#543610000000
1!
1*
b10 6
19
1>
1C
b10 G
#543620000000
0!
0*
09
0>
0C
#543630000000
1!
1*
b11 6
19
1>
1C
b11 G
#543640000000
0!
0*
09
0>
0C
#543650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#543660000000
0!
0*
09
0>
0C
#543670000000
1!
1*
b101 6
19
1>
1C
b101 G
#543680000000
0!
0*
09
0>
0C
#543690000000
1!
1*
b110 6
19
1>
1C
b110 G
#543700000000
0!
0*
09
0>
0C
#543710000000
1!
1*
b111 6
19
1>
1C
b111 G
#543720000000
0!
0*
09
0>
0C
#543730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#543740000000
0!
0*
09
0>
0C
#543750000000
1!
1*
b1 6
19
1>
1C
b1 G
#543760000000
0!
0*
09
0>
0C
#543770000000
1!
1*
b10 6
19
1>
1C
b10 G
#543780000000
0!
0*
09
0>
0C
#543790000000
1!
1*
b11 6
19
1>
1C
b11 G
#543800000000
0!
0*
09
0>
0C
#543810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#543820000000
0!
0*
09
0>
0C
#543830000000
1!
1*
b101 6
19
1>
1C
b101 G
#543840000000
0!
0*
09
0>
0C
#543850000000
1!
1*
b110 6
19
1>
1C
b110 G
#543860000000
0!
0*
09
0>
0C
#543870000000
1!
1*
b111 6
19
1>
1C
b111 G
#543880000000
0!
0*
09
0>
0C
#543890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#543900000000
0!
0*
09
0>
0C
#543910000000
1!
1*
b1 6
19
1>
1C
b1 G
#543920000000
0!
0*
09
0>
0C
#543930000000
1!
1*
b10 6
19
1>
1C
b10 G
#543940000000
0!
0*
09
0>
0C
#543950000000
1!
1*
b11 6
19
1>
1C
b11 G
#543960000000
0!
0*
09
0>
0C
#543970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#543980000000
0!
0*
09
0>
0C
#543990000000
1!
1*
b101 6
19
1>
1C
b101 G
#544000000000
0!
0*
09
0>
0C
#544010000000
1!
1*
b110 6
19
1>
1C
b110 G
#544020000000
0!
0*
09
0>
0C
#544030000000
1!
1*
b111 6
19
1>
1C
b111 G
#544040000000
0!
1"
0*
1+
09
1:
0>
0C
#544050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#544060000000
0!
0*
09
0>
0C
#544070000000
1!
1*
b1 6
19
1>
1C
b1 G
#544080000000
0!
0*
09
0>
0C
#544090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#544100000000
0!
0*
09
0>
0C
#544110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#544120000000
0!
0*
09
0>
0C
#544130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#544140000000
0!
0*
09
0>
0C
#544150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#544160000000
0!
0#
0*
0,
09
0>
0?
0C
#544170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#544180000000
0!
0*
09
0>
0C
#544190000000
1!
1*
19
1>
1C
#544200000000
0!
0*
09
0>
0C
#544210000000
1!
1*
19
1>
1C
#544220000000
0!
0*
09
0>
0C
#544230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#544240000000
0!
0*
09
0>
0C
#544250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#544260000000
0!
0*
09
0>
0C
#544270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#544280000000
0!
0*
09
0>
0C
#544290000000
1!
1*
b10 6
19
1>
1C
b10 G
#544300000000
0!
0*
09
0>
0C
#544310000000
1!
1*
b11 6
19
1>
1C
b11 G
#544320000000
0!
0*
09
0>
0C
#544330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#544340000000
0!
0*
09
0>
0C
#544350000000
1!
1*
b101 6
19
1>
1C
b101 G
#544360000000
0!
0*
09
0>
0C
#544370000000
1!
1*
b110 6
19
1>
1C
b110 G
#544380000000
0!
0*
09
0>
0C
#544390000000
1!
1*
b111 6
19
1>
1C
b111 G
#544400000000
0!
0*
09
0>
0C
#544410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#544420000000
0!
0*
09
0>
0C
#544430000000
1!
1*
b1 6
19
1>
1C
b1 G
#544440000000
0!
0*
09
0>
0C
#544450000000
1!
1*
b10 6
19
1>
1C
b10 G
#544460000000
0!
0*
09
0>
0C
#544470000000
1!
1*
b11 6
19
1>
1C
b11 G
#544480000000
0!
0*
09
0>
0C
#544490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#544500000000
0!
0*
09
0>
0C
#544510000000
1!
1*
b101 6
19
1>
1C
b101 G
#544520000000
0!
0*
09
0>
0C
#544530000000
1!
1*
b110 6
19
1>
1C
b110 G
#544540000000
0!
0*
09
0>
0C
#544550000000
1!
1*
b111 6
19
1>
1C
b111 G
#544560000000
0!
0*
09
0>
0C
#544570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#544580000000
0!
0*
09
0>
0C
#544590000000
1!
1*
b1 6
19
1>
1C
b1 G
#544600000000
0!
0*
09
0>
0C
#544610000000
1!
1*
b10 6
19
1>
1C
b10 G
#544620000000
0!
0*
09
0>
0C
#544630000000
1!
1*
b11 6
19
1>
1C
b11 G
#544640000000
0!
0*
09
0>
0C
#544650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#544660000000
0!
0*
09
0>
0C
#544670000000
1!
1*
b101 6
19
1>
1C
b101 G
#544680000000
0!
0*
09
0>
0C
#544690000000
1!
1*
b110 6
19
1>
1C
b110 G
#544700000000
0!
0*
09
0>
0C
#544710000000
1!
1*
b111 6
19
1>
1C
b111 G
#544720000000
0!
1"
0*
1+
09
1:
0>
0C
#544730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#544740000000
0!
0*
09
0>
0C
#544750000000
1!
1*
b1 6
19
1>
1C
b1 G
#544760000000
0!
0*
09
0>
0C
#544770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#544780000000
0!
0*
09
0>
0C
#544790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#544800000000
0!
0*
09
0>
0C
#544810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#544820000000
0!
0*
09
0>
0C
#544830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#544840000000
0!
0#
0*
0,
09
0>
0?
0C
#544850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#544860000000
0!
0*
09
0>
0C
#544870000000
1!
1*
19
1>
1C
#544880000000
0!
0*
09
0>
0C
#544890000000
1!
1*
19
1>
1C
#544900000000
0!
0*
09
0>
0C
#544910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#544920000000
0!
0*
09
0>
0C
#544930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#544940000000
0!
0*
09
0>
0C
#544950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#544960000000
0!
0*
09
0>
0C
#544970000000
1!
1*
b10 6
19
1>
1C
b10 G
#544980000000
0!
0*
09
0>
0C
#544990000000
1!
1*
b11 6
19
1>
1C
b11 G
#545000000000
0!
0*
09
0>
0C
#545010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#545020000000
0!
0*
09
0>
0C
#545030000000
1!
1*
b101 6
19
1>
1C
b101 G
#545040000000
0!
0*
09
0>
0C
#545050000000
1!
1*
b110 6
19
1>
1C
b110 G
#545060000000
0!
0*
09
0>
0C
#545070000000
1!
1*
b111 6
19
1>
1C
b111 G
#545080000000
0!
0*
09
0>
0C
#545090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#545100000000
0!
0*
09
0>
0C
#545110000000
1!
1*
b1 6
19
1>
1C
b1 G
#545120000000
0!
0*
09
0>
0C
#545130000000
1!
1*
b10 6
19
1>
1C
b10 G
#545140000000
0!
0*
09
0>
0C
#545150000000
1!
1*
b11 6
19
1>
1C
b11 G
#545160000000
0!
0*
09
0>
0C
#545170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#545180000000
0!
0*
09
0>
0C
#545190000000
1!
1*
b101 6
19
1>
1C
b101 G
#545200000000
0!
0*
09
0>
0C
#545210000000
1!
1*
b110 6
19
1>
1C
b110 G
#545220000000
0!
0*
09
0>
0C
#545230000000
1!
1*
b111 6
19
1>
1C
b111 G
#545240000000
0!
0*
09
0>
0C
#545250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#545260000000
0!
0*
09
0>
0C
#545270000000
1!
1*
b1 6
19
1>
1C
b1 G
#545280000000
0!
0*
09
0>
0C
#545290000000
1!
1*
b10 6
19
1>
1C
b10 G
#545300000000
0!
0*
09
0>
0C
#545310000000
1!
1*
b11 6
19
1>
1C
b11 G
#545320000000
0!
0*
09
0>
0C
#545330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#545340000000
0!
0*
09
0>
0C
#545350000000
1!
1*
b101 6
19
1>
1C
b101 G
#545360000000
0!
0*
09
0>
0C
#545370000000
1!
1*
b110 6
19
1>
1C
b110 G
#545380000000
0!
0*
09
0>
0C
#545390000000
1!
1*
b111 6
19
1>
1C
b111 G
#545400000000
0!
1"
0*
1+
09
1:
0>
0C
#545410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#545420000000
0!
0*
09
0>
0C
#545430000000
1!
1*
b1 6
19
1>
1C
b1 G
#545440000000
0!
0*
09
0>
0C
#545450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#545460000000
0!
0*
09
0>
0C
#545470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#545480000000
0!
0*
09
0>
0C
#545490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#545500000000
0!
0*
09
0>
0C
#545510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#545520000000
0!
0#
0*
0,
09
0>
0?
0C
#545530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#545540000000
0!
0*
09
0>
0C
#545550000000
1!
1*
19
1>
1C
#545560000000
0!
0*
09
0>
0C
#545570000000
1!
1*
19
1>
1C
#545580000000
0!
0*
09
0>
0C
#545590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#545600000000
0!
0*
09
0>
0C
#545610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#545620000000
0!
0*
09
0>
0C
#545630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#545640000000
0!
0*
09
0>
0C
#545650000000
1!
1*
b10 6
19
1>
1C
b10 G
#545660000000
0!
0*
09
0>
0C
#545670000000
1!
1*
b11 6
19
1>
1C
b11 G
#545680000000
0!
0*
09
0>
0C
#545690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#545700000000
0!
0*
09
0>
0C
#545710000000
1!
1*
b101 6
19
1>
1C
b101 G
#545720000000
0!
0*
09
0>
0C
#545730000000
1!
1*
b110 6
19
1>
1C
b110 G
#545740000000
0!
0*
09
0>
0C
#545750000000
1!
1*
b111 6
19
1>
1C
b111 G
#545760000000
0!
0*
09
0>
0C
#545770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#545780000000
0!
0*
09
0>
0C
#545790000000
1!
1*
b1 6
19
1>
1C
b1 G
#545800000000
0!
0*
09
0>
0C
#545810000000
1!
1*
b10 6
19
1>
1C
b10 G
#545820000000
0!
0*
09
0>
0C
#545830000000
1!
1*
b11 6
19
1>
1C
b11 G
#545840000000
0!
0*
09
0>
0C
#545850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#545860000000
0!
0*
09
0>
0C
#545870000000
1!
1*
b101 6
19
1>
1C
b101 G
#545880000000
0!
0*
09
0>
0C
#545890000000
1!
1*
b110 6
19
1>
1C
b110 G
#545900000000
0!
0*
09
0>
0C
#545910000000
1!
1*
b111 6
19
1>
1C
b111 G
#545920000000
0!
0*
09
0>
0C
#545930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#545940000000
0!
0*
09
0>
0C
#545950000000
1!
1*
b1 6
19
1>
1C
b1 G
#545960000000
0!
0*
09
0>
0C
#545970000000
1!
1*
b10 6
19
1>
1C
b10 G
#545980000000
0!
0*
09
0>
0C
#545990000000
1!
1*
b11 6
19
1>
1C
b11 G
#546000000000
0!
0*
09
0>
0C
#546010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#546020000000
0!
0*
09
0>
0C
#546030000000
1!
1*
b101 6
19
1>
1C
b101 G
#546040000000
0!
0*
09
0>
0C
#546050000000
1!
1*
b110 6
19
1>
1C
b110 G
#546060000000
0!
0*
09
0>
0C
#546070000000
1!
1*
b111 6
19
1>
1C
b111 G
#546080000000
0!
1"
0*
1+
09
1:
0>
0C
#546090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#546100000000
0!
0*
09
0>
0C
#546110000000
1!
1*
b1 6
19
1>
1C
b1 G
#546120000000
0!
0*
09
0>
0C
#546130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#546140000000
0!
0*
09
0>
0C
#546150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#546160000000
0!
0*
09
0>
0C
#546170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#546180000000
0!
0*
09
0>
0C
#546190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#546200000000
0!
0#
0*
0,
09
0>
0?
0C
#546210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#546220000000
0!
0*
09
0>
0C
#546230000000
1!
1*
19
1>
1C
#546240000000
0!
0*
09
0>
0C
#546250000000
1!
1*
19
1>
1C
#546260000000
0!
0*
09
0>
0C
#546270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#546280000000
0!
0*
09
0>
0C
#546290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#546300000000
0!
0*
09
0>
0C
#546310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#546320000000
0!
0*
09
0>
0C
#546330000000
1!
1*
b10 6
19
1>
1C
b10 G
#546340000000
0!
0*
09
0>
0C
#546350000000
1!
1*
b11 6
19
1>
1C
b11 G
#546360000000
0!
0*
09
0>
0C
#546370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#546380000000
0!
0*
09
0>
0C
#546390000000
1!
1*
b101 6
19
1>
1C
b101 G
#546400000000
0!
0*
09
0>
0C
#546410000000
1!
1*
b110 6
19
1>
1C
b110 G
#546420000000
0!
0*
09
0>
0C
#546430000000
1!
1*
b111 6
19
1>
1C
b111 G
#546440000000
0!
0*
09
0>
0C
#546450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#546460000000
0!
0*
09
0>
0C
#546470000000
1!
1*
b1 6
19
1>
1C
b1 G
#546480000000
0!
0*
09
0>
0C
#546490000000
1!
1*
b10 6
19
1>
1C
b10 G
#546500000000
0!
0*
09
0>
0C
#546510000000
1!
1*
b11 6
19
1>
1C
b11 G
#546520000000
0!
0*
09
0>
0C
#546530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#546540000000
0!
0*
09
0>
0C
#546550000000
1!
1*
b101 6
19
1>
1C
b101 G
#546560000000
0!
0*
09
0>
0C
#546570000000
1!
1*
b110 6
19
1>
1C
b110 G
#546580000000
0!
0*
09
0>
0C
#546590000000
1!
1*
b111 6
19
1>
1C
b111 G
#546600000000
0!
0*
09
0>
0C
#546610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#546620000000
0!
0*
09
0>
0C
#546630000000
1!
1*
b1 6
19
1>
1C
b1 G
#546640000000
0!
0*
09
0>
0C
#546650000000
1!
1*
b10 6
19
1>
1C
b10 G
#546660000000
0!
0*
09
0>
0C
#546670000000
1!
1*
b11 6
19
1>
1C
b11 G
#546680000000
0!
0*
09
0>
0C
#546690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#546700000000
0!
0*
09
0>
0C
#546710000000
1!
1*
b101 6
19
1>
1C
b101 G
#546720000000
0!
0*
09
0>
0C
#546730000000
1!
1*
b110 6
19
1>
1C
b110 G
#546740000000
0!
0*
09
0>
0C
#546750000000
1!
1*
b111 6
19
1>
1C
b111 G
#546760000000
0!
1"
0*
1+
09
1:
0>
0C
#546770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#546780000000
0!
0*
09
0>
0C
#546790000000
1!
1*
b1 6
19
1>
1C
b1 G
#546800000000
0!
0*
09
0>
0C
#546810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#546820000000
0!
0*
09
0>
0C
#546830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#546840000000
0!
0*
09
0>
0C
#546850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#546860000000
0!
0*
09
0>
0C
#546870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#546880000000
0!
0#
0*
0,
09
0>
0?
0C
#546890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#546900000000
0!
0*
09
0>
0C
#546910000000
1!
1*
19
1>
1C
#546920000000
0!
0*
09
0>
0C
#546930000000
1!
1*
19
1>
1C
#546940000000
0!
0*
09
0>
0C
#546950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#546960000000
0!
0*
09
0>
0C
#546970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#546980000000
0!
0*
09
0>
0C
#546990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#547000000000
0!
0*
09
0>
0C
#547010000000
1!
1*
b10 6
19
1>
1C
b10 G
#547020000000
0!
0*
09
0>
0C
#547030000000
1!
1*
b11 6
19
1>
1C
b11 G
#547040000000
0!
0*
09
0>
0C
#547050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#547060000000
0!
0*
09
0>
0C
#547070000000
1!
1*
b101 6
19
1>
1C
b101 G
#547080000000
0!
0*
09
0>
0C
#547090000000
1!
1*
b110 6
19
1>
1C
b110 G
#547100000000
0!
0*
09
0>
0C
#547110000000
1!
1*
b111 6
19
1>
1C
b111 G
#547120000000
0!
0*
09
0>
0C
#547130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#547140000000
0!
0*
09
0>
0C
#547150000000
1!
1*
b1 6
19
1>
1C
b1 G
#547160000000
0!
0*
09
0>
0C
#547170000000
1!
1*
b10 6
19
1>
1C
b10 G
#547180000000
0!
0*
09
0>
0C
#547190000000
1!
1*
b11 6
19
1>
1C
b11 G
#547200000000
0!
0*
09
0>
0C
#547210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#547220000000
0!
0*
09
0>
0C
#547230000000
1!
1*
b101 6
19
1>
1C
b101 G
#547240000000
0!
0*
09
0>
0C
#547250000000
1!
1*
b110 6
19
1>
1C
b110 G
#547260000000
0!
0*
09
0>
0C
#547270000000
1!
1*
b111 6
19
1>
1C
b111 G
#547280000000
0!
0*
09
0>
0C
#547290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#547300000000
0!
0*
09
0>
0C
#547310000000
1!
1*
b1 6
19
1>
1C
b1 G
#547320000000
0!
0*
09
0>
0C
#547330000000
1!
1*
b10 6
19
1>
1C
b10 G
#547340000000
0!
0*
09
0>
0C
#547350000000
1!
1*
b11 6
19
1>
1C
b11 G
#547360000000
0!
0*
09
0>
0C
#547370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#547380000000
0!
0*
09
0>
0C
#547390000000
1!
1*
b101 6
19
1>
1C
b101 G
#547400000000
0!
0*
09
0>
0C
#547410000000
1!
1*
b110 6
19
1>
1C
b110 G
#547420000000
0!
0*
09
0>
0C
#547430000000
1!
1*
b111 6
19
1>
1C
b111 G
#547440000000
0!
1"
0*
1+
09
1:
0>
0C
#547450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#547460000000
0!
0*
09
0>
0C
#547470000000
1!
1*
b1 6
19
1>
1C
b1 G
#547480000000
0!
0*
09
0>
0C
#547490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#547500000000
0!
0*
09
0>
0C
#547510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#547520000000
0!
0*
09
0>
0C
#547530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#547540000000
0!
0*
09
0>
0C
#547550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#547560000000
0!
0#
0*
0,
09
0>
0?
0C
#547570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#547580000000
0!
0*
09
0>
0C
#547590000000
1!
1*
19
1>
1C
#547600000000
0!
0*
09
0>
0C
#547610000000
1!
1*
19
1>
1C
#547620000000
0!
0*
09
0>
0C
#547630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#547640000000
0!
0*
09
0>
0C
#547650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#547660000000
0!
0*
09
0>
0C
#547670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#547680000000
0!
0*
09
0>
0C
#547690000000
1!
1*
b10 6
19
1>
1C
b10 G
#547700000000
0!
0*
09
0>
0C
#547710000000
1!
1*
b11 6
19
1>
1C
b11 G
#547720000000
0!
0*
09
0>
0C
#547730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#547740000000
0!
0*
09
0>
0C
#547750000000
1!
1*
b101 6
19
1>
1C
b101 G
#547760000000
0!
0*
09
0>
0C
#547770000000
1!
1*
b110 6
19
1>
1C
b110 G
#547780000000
0!
0*
09
0>
0C
#547790000000
1!
1*
b111 6
19
1>
1C
b111 G
#547800000000
0!
0*
09
0>
0C
#547810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#547820000000
0!
0*
09
0>
0C
#547830000000
1!
1*
b1 6
19
1>
1C
b1 G
#547840000000
0!
0*
09
0>
0C
#547850000000
1!
1*
b10 6
19
1>
1C
b10 G
#547860000000
0!
0*
09
0>
0C
#547870000000
1!
1*
b11 6
19
1>
1C
b11 G
#547880000000
0!
0*
09
0>
0C
#547890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#547900000000
0!
0*
09
0>
0C
#547910000000
1!
1*
b101 6
19
1>
1C
b101 G
#547920000000
0!
0*
09
0>
0C
#547930000000
1!
1*
b110 6
19
1>
1C
b110 G
#547940000000
0!
0*
09
0>
0C
#547950000000
1!
1*
b111 6
19
1>
1C
b111 G
#547960000000
0!
0*
09
0>
0C
#547970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#547980000000
0!
0*
09
0>
0C
#547990000000
1!
1*
b1 6
19
1>
1C
b1 G
#548000000000
0!
0*
09
0>
0C
#548010000000
1!
1*
b10 6
19
1>
1C
b10 G
#548020000000
0!
0*
09
0>
0C
#548030000000
1!
1*
b11 6
19
1>
1C
b11 G
#548040000000
0!
0*
09
0>
0C
#548050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#548060000000
0!
0*
09
0>
0C
#548070000000
1!
1*
b101 6
19
1>
1C
b101 G
#548080000000
0!
0*
09
0>
0C
#548090000000
1!
1*
b110 6
19
1>
1C
b110 G
#548100000000
0!
0*
09
0>
0C
#548110000000
1!
1*
b111 6
19
1>
1C
b111 G
#548120000000
0!
1"
0*
1+
09
1:
0>
0C
#548130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#548140000000
0!
0*
09
0>
0C
#548150000000
1!
1*
b1 6
19
1>
1C
b1 G
#548160000000
0!
0*
09
0>
0C
#548170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#548180000000
0!
0*
09
0>
0C
#548190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#548200000000
0!
0*
09
0>
0C
#548210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#548220000000
0!
0*
09
0>
0C
#548230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#548240000000
0!
0#
0*
0,
09
0>
0?
0C
#548250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#548260000000
0!
0*
09
0>
0C
#548270000000
1!
1*
19
1>
1C
#548280000000
0!
0*
09
0>
0C
#548290000000
1!
1*
19
1>
1C
#548300000000
0!
0*
09
0>
0C
#548310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#548320000000
0!
0*
09
0>
0C
#548330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#548340000000
0!
0*
09
0>
0C
#548350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#548360000000
0!
0*
09
0>
0C
#548370000000
1!
1*
b10 6
19
1>
1C
b10 G
#548380000000
0!
0*
09
0>
0C
#548390000000
1!
1*
b11 6
19
1>
1C
b11 G
#548400000000
0!
0*
09
0>
0C
#548410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#548420000000
0!
0*
09
0>
0C
#548430000000
1!
1*
b101 6
19
1>
1C
b101 G
#548440000000
0!
0*
09
0>
0C
#548450000000
1!
1*
b110 6
19
1>
1C
b110 G
#548460000000
0!
0*
09
0>
0C
#548470000000
1!
1*
b111 6
19
1>
1C
b111 G
#548480000000
0!
0*
09
0>
0C
#548490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#548500000000
0!
0*
09
0>
0C
#548510000000
1!
1*
b1 6
19
1>
1C
b1 G
#548520000000
0!
0*
09
0>
0C
#548530000000
1!
1*
b10 6
19
1>
1C
b10 G
#548540000000
0!
0*
09
0>
0C
#548550000000
1!
1*
b11 6
19
1>
1C
b11 G
#548560000000
0!
0*
09
0>
0C
#548570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#548580000000
0!
0*
09
0>
0C
#548590000000
1!
1*
b101 6
19
1>
1C
b101 G
#548600000000
0!
0*
09
0>
0C
#548610000000
1!
1*
b110 6
19
1>
1C
b110 G
#548620000000
0!
0*
09
0>
0C
#548630000000
1!
1*
b111 6
19
1>
1C
b111 G
#548640000000
0!
0*
09
0>
0C
#548650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#548660000000
0!
0*
09
0>
0C
#548670000000
1!
1*
b1 6
19
1>
1C
b1 G
#548680000000
0!
0*
09
0>
0C
#548690000000
1!
1*
b10 6
19
1>
1C
b10 G
#548700000000
0!
0*
09
0>
0C
#548710000000
1!
1*
b11 6
19
1>
1C
b11 G
#548720000000
0!
0*
09
0>
0C
#548730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#548740000000
0!
0*
09
0>
0C
#548750000000
1!
1*
b101 6
19
1>
1C
b101 G
#548760000000
0!
0*
09
0>
0C
#548770000000
1!
1*
b110 6
19
1>
1C
b110 G
#548780000000
0!
0*
09
0>
0C
#548790000000
1!
1*
b111 6
19
1>
1C
b111 G
#548800000000
0!
1"
0*
1+
09
1:
0>
0C
#548810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#548820000000
0!
0*
09
0>
0C
#548830000000
1!
1*
b1 6
19
1>
1C
b1 G
#548840000000
0!
0*
09
0>
0C
#548850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#548860000000
0!
0*
09
0>
0C
#548870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#548880000000
0!
0*
09
0>
0C
#548890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#548900000000
0!
0*
09
0>
0C
#548910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#548920000000
0!
0#
0*
0,
09
0>
0?
0C
#548930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#548940000000
0!
0*
09
0>
0C
#548950000000
1!
1*
19
1>
1C
#548960000000
0!
0*
09
0>
0C
#548970000000
1!
1*
19
1>
1C
#548980000000
0!
0*
09
0>
0C
#548990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#549000000000
0!
0*
09
0>
0C
#549010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#549020000000
0!
0*
09
0>
0C
#549030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#549040000000
0!
0*
09
0>
0C
#549050000000
1!
1*
b10 6
19
1>
1C
b10 G
#549060000000
0!
0*
09
0>
0C
#549070000000
1!
1*
b11 6
19
1>
1C
b11 G
#549080000000
0!
0*
09
0>
0C
#549090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#549100000000
0!
0*
09
0>
0C
#549110000000
1!
1*
b101 6
19
1>
1C
b101 G
#549120000000
0!
0*
09
0>
0C
#549130000000
1!
1*
b110 6
19
1>
1C
b110 G
#549140000000
0!
0*
09
0>
0C
#549150000000
1!
1*
b111 6
19
1>
1C
b111 G
#549160000000
0!
0*
09
0>
0C
#549170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#549180000000
0!
0*
09
0>
0C
#549190000000
1!
1*
b1 6
19
1>
1C
b1 G
#549200000000
0!
0*
09
0>
0C
#549210000000
1!
1*
b10 6
19
1>
1C
b10 G
#549220000000
0!
0*
09
0>
0C
#549230000000
1!
1*
b11 6
19
1>
1C
b11 G
#549240000000
0!
0*
09
0>
0C
#549250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#549260000000
0!
0*
09
0>
0C
#549270000000
1!
1*
b101 6
19
1>
1C
b101 G
#549280000000
0!
0*
09
0>
0C
#549290000000
1!
1*
b110 6
19
1>
1C
b110 G
#549300000000
0!
0*
09
0>
0C
#549310000000
1!
1*
b111 6
19
1>
1C
b111 G
#549320000000
0!
0*
09
0>
0C
#549330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#549340000000
0!
0*
09
0>
0C
#549350000000
1!
1*
b1 6
19
1>
1C
b1 G
#549360000000
0!
0*
09
0>
0C
#549370000000
1!
1*
b10 6
19
1>
1C
b10 G
#549380000000
0!
0*
09
0>
0C
#549390000000
1!
1*
b11 6
19
1>
1C
b11 G
#549400000000
0!
0*
09
0>
0C
#549410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#549420000000
0!
0*
09
0>
0C
#549430000000
1!
1*
b101 6
19
1>
1C
b101 G
#549440000000
0!
0*
09
0>
0C
#549450000000
1!
1*
b110 6
19
1>
1C
b110 G
#549460000000
0!
0*
09
0>
0C
#549470000000
1!
1*
b111 6
19
1>
1C
b111 G
#549480000000
0!
1"
0*
1+
09
1:
0>
0C
#549490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#549500000000
0!
0*
09
0>
0C
#549510000000
1!
1*
b1 6
19
1>
1C
b1 G
#549520000000
0!
0*
09
0>
0C
#549530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#549540000000
0!
0*
09
0>
0C
#549550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#549560000000
0!
0*
09
0>
0C
#549570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#549580000000
0!
0*
09
0>
0C
#549590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#549600000000
0!
0#
0*
0,
09
0>
0?
0C
#549610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#549620000000
0!
0*
09
0>
0C
#549630000000
1!
1*
19
1>
1C
#549640000000
0!
0*
09
0>
0C
#549650000000
1!
1*
19
1>
1C
#549660000000
0!
0*
09
0>
0C
#549670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#549680000000
0!
0*
09
0>
0C
#549690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#549700000000
0!
0*
09
0>
0C
#549710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#549720000000
0!
0*
09
0>
0C
#549730000000
1!
1*
b10 6
19
1>
1C
b10 G
#549740000000
0!
0*
09
0>
0C
#549750000000
1!
1*
b11 6
19
1>
1C
b11 G
#549760000000
0!
0*
09
0>
0C
#549770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#549780000000
0!
0*
09
0>
0C
#549790000000
1!
1*
b101 6
19
1>
1C
b101 G
#549800000000
0!
0*
09
0>
0C
#549810000000
1!
1*
b110 6
19
1>
1C
b110 G
#549820000000
0!
0*
09
0>
0C
#549830000000
1!
1*
b111 6
19
1>
1C
b111 G
#549840000000
0!
0*
09
0>
0C
#549850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#549860000000
0!
0*
09
0>
0C
#549870000000
1!
1*
b1 6
19
1>
1C
b1 G
#549880000000
0!
0*
09
0>
0C
#549890000000
1!
1*
b10 6
19
1>
1C
b10 G
#549900000000
0!
0*
09
0>
0C
#549910000000
1!
1*
b11 6
19
1>
1C
b11 G
#549920000000
0!
0*
09
0>
0C
#549930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#549940000000
0!
0*
09
0>
0C
#549950000000
1!
1*
b101 6
19
1>
1C
b101 G
#549960000000
0!
0*
09
0>
0C
#549970000000
1!
1*
b110 6
19
1>
1C
b110 G
#549980000000
0!
0*
09
0>
0C
#549990000000
1!
1*
b111 6
19
1>
1C
b111 G
#550000000000
0!
0*
09
0>
0C
#550010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#550020000000
0!
0*
09
0>
0C
#550030000000
1!
1*
b1 6
19
1>
1C
b1 G
#550040000000
0!
0*
09
0>
0C
#550050000000
1!
1*
b10 6
19
1>
1C
b10 G
#550060000000
0!
0*
09
0>
0C
#550070000000
1!
1*
b11 6
19
1>
1C
b11 G
#550080000000
0!
0*
09
0>
0C
#550090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#550100000000
0!
0*
09
0>
0C
#550110000000
1!
1*
b101 6
19
1>
1C
b101 G
#550120000000
0!
0*
09
0>
0C
#550130000000
1!
1*
b110 6
19
1>
1C
b110 G
#550140000000
0!
0*
09
0>
0C
#550150000000
1!
1*
b111 6
19
1>
1C
b111 G
#550160000000
0!
1"
0*
1+
09
1:
0>
0C
#550170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#550180000000
0!
0*
09
0>
0C
#550190000000
1!
1*
b1 6
19
1>
1C
b1 G
#550200000000
0!
0*
09
0>
0C
#550210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#550220000000
0!
0*
09
0>
0C
#550230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#550240000000
0!
0*
09
0>
0C
#550250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#550260000000
0!
0*
09
0>
0C
#550270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#550280000000
0!
0#
0*
0,
09
0>
0?
0C
#550290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#550300000000
0!
0*
09
0>
0C
#550310000000
1!
1*
19
1>
1C
#550320000000
0!
0*
09
0>
0C
#550330000000
1!
1*
19
1>
1C
#550340000000
0!
0*
09
0>
0C
#550350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#550360000000
0!
0*
09
0>
0C
#550370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#550380000000
0!
0*
09
0>
0C
#550390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#550400000000
0!
0*
09
0>
0C
#550410000000
1!
1*
b10 6
19
1>
1C
b10 G
#550420000000
0!
0*
09
0>
0C
#550430000000
1!
1*
b11 6
19
1>
1C
b11 G
#550440000000
0!
0*
09
0>
0C
#550450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#550460000000
0!
0*
09
0>
0C
#550470000000
1!
1*
b101 6
19
1>
1C
b101 G
#550480000000
0!
0*
09
0>
0C
#550490000000
1!
1*
b110 6
19
1>
1C
b110 G
#550500000000
0!
0*
09
0>
0C
#550510000000
1!
1*
b111 6
19
1>
1C
b111 G
#550520000000
0!
0*
09
0>
0C
#550530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#550540000000
0!
0*
09
0>
0C
#550550000000
1!
1*
b1 6
19
1>
1C
b1 G
#550560000000
0!
0*
09
0>
0C
#550570000000
1!
1*
b10 6
19
1>
1C
b10 G
#550580000000
0!
0*
09
0>
0C
#550590000000
1!
1*
b11 6
19
1>
1C
b11 G
#550600000000
0!
0*
09
0>
0C
#550610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#550620000000
0!
0*
09
0>
0C
#550630000000
1!
1*
b101 6
19
1>
1C
b101 G
#550640000000
0!
0*
09
0>
0C
#550650000000
1!
1*
b110 6
19
1>
1C
b110 G
#550660000000
0!
0*
09
0>
0C
#550670000000
1!
1*
b111 6
19
1>
1C
b111 G
#550680000000
0!
0*
09
0>
0C
#550690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#550700000000
0!
0*
09
0>
0C
#550710000000
1!
1*
b1 6
19
1>
1C
b1 G
#550720000000
0!
0*
09
0>
0C
#550730000000
1!
1*
b10 6
19
1>
1C
b10 G
#550740000000
0!
0*
09
0>
0C
#550750000000
1!
1*
b11 6
19
1>
1C
b11 G
#550760000000
0!
0*
09
0>
0C
#550770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#550780000000
0!
0*
09
0>
0C
#550790000000
1!
1*
b101 6
19
1>
1C
b101 G
#550800000000
0!
0*
09
0>
0C
#550810000000
1!
1*
b110 6
19
1>
1C
b110 G
#550820000000
0!
0*
09
0>
0C
#550830000000
1!
1*
b111 6
19
1>
1C
b111 G
#550840000000
0!
1"
0*
1+
09
1:
0>
0C
#550850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#550860000000
0!
0*
09
0>
0C
#550870000000
1!
1*
b1 6
19
1>
1C
b1 G
#550880000000
0!
0*
09
0>
0C
#550890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#550900000000
0!
0*
09
0>
0C
#550910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#550920000000
0!
0*
09
0>
0C
#550930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#550940000000
0!
0*
09
0>
0C
#550950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#550960000000
0!
0#
0*
0,
09
0>
0?
0C
#550970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#550980000000
0!
0*
09
0>
0C
#550990000000
1!
1*
19
1>
1C
#551000000000
0!
0*
09
0>
0C
#551010000000
1!
1*
19
1>
1C
#551020000000
0!
0*
09
0>
0C
#551030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#551040000000
0!
0*
09
0>
0C
#551050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#551060000000
0!
0*
09
0>
0C
#551070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#551080000000
0!
0*
09
0>
0C
#551090000000
1!
1*
b10 6
19
1>
1C
b10 G
#551100000000
0!
0*
09
0>
0C
#551110000000
1!
1*
b11 6
19
1>
1C
b11 G
#551120000000
0!
0*
09
0>
0C
#551130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#551140000000
0!
0*
09
0>
0C
#551150000000
1!
1*
b101 6
19
1>
1C
b101 G
#551160000000
0!
0*
09
0>
0C
#551170000000
1!
1*
b110 6
19
1>
1C
b110 G
#551180000000
0!
0*
09
0>
0C
#551190000000
1!
1*
b111 6
19
1>
1C
b111 G
#551200000000
0!
0*
09
0>
0C
#551210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#551220000000
0!
0*
09
0>
0C
#551230000000
1!
1*
b1 6
19
1>
1C
b1 G
#551240000000
0!
0*
09
0>
0C
#551250000000
1!
1*
b10 6
19
1>
1C
b10 G
#551260000000
0!
0*
09
0>
0C
#551270000000
1!
1*
b11 6
19
1>
1C
b11 G
#551280000000
0!
0*
09
0>
0C
#551290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#551300000000
0!
0*
09
0>
0C
#551310000000
1!
1*
b101 6
19
1>
1C
b101 G
#551320000000
0!
0*
09
0>
0C
#551330000000
1!
1*
b110 6
19
1>
1C
b110 G
#551340000000
0!
0*
09
0>
0C
#551350000000
1!
1*
b111 6
19
1>
1C
b111 G
#551360000000
0!
0*
09
0>
0C
#551370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#551380000000
0!
0*
09
0>
0C
#551390000000
1!
1*
b1 6
19
1>
1C
b1 G
#551400000000
0!
0*
09
0>
0C
#551410000000
1!
1*
b10 6
19
1>
1C
b10 G
#551420000000
0!
0*
09
0>
0C
#551430000000
1!
1*
b11 6
19
1>
1C
b11 G
#551440000000
0!
0*
09
0>
0C
#551450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#551460000000
0!
0*
09
0>
0C
#551470000000
1!
1*
b101 6
19
1>
1C
b101 G
#551480000000
0!
0*
09
0>
0C
#551490000000
1!
1*
b110 6
19
1>
1C
b110 G
#551500000000
0!
0*
09
0>
0C
#551510000000
1!
1*
b111 6
19
1>
1C
b111 G
#551520000000
0!
1"
0*
1+
09
1:
0>
0C
#551530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#551540000000
0!
0*
09
0>
0C
#551550000000
1!
1*
b1 6
19
1>
1C
b1 G
#551560000000
0!
0*
09
0>
0C
#551570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#551580000000
0!
0*
09
0>
0C
#551590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#551600000000
0!
0*
09
0>
0C
#551610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#551620000000
0!
0*
09
0>
0C
#551630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#551640000000
0!
0#
0*
0,
09
0>
0?
0C
#551650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#551660000000
0!
0*
09
0>
0C
#551670000000
1!
1*
19
1>
1C
#551680000000
0!
0*
09
0>
0C
#551690000000
1!
1*
19
1>
1C
#551700000000
0!
0*
09
0>
0C
#551710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#551720000000
0!
0*
09
0>
0C
#551730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#551740000000
0!
0*
09
0>
0C
#551750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#551760000000
0!
0*
09
0>
0C
#551770000000
1!
1*
b10 6
19
1>
1C
b10 G
#551780000000
0!
0*
09
0>
0C
#551790000000
1!
1*
b11 6
19
1>
1C
b11 G
#551800000000
0!
0*
09
0>
0C
#551810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#551820000000
0!
0*
09
0>
0C
#551830000000
1!
1*
b101 6
19
1>
1C
b101 G
#551840000000
0!
0*
09
0>
0C
#551850000000
1!
1*
b110 6
19
1>
1C
b110 G
#551860000000
0!
0*
09
0>
0C
#551870000000
1!
1*
b111 6
19
1>
1C
b111 G
#551880000000
0!
0*
09
0>
0C
#551890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#551900000000
0!
0*
09
0>
0C
#551910000000
1!
1*
b1 6
19
1>
1C
b1 G
#551920000000
0!
0*
09
0>
0C
#551930000000
1!
1*
b10 6
19
1>
1C
b10 G
#551940000000
0!
0*
09
0>
0C
#551950000000
1!
1*
b11 6
19
1>
1C
b11 G
#551960000000
0!
0*
09
0>
0C
#551970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#551980000000
0!
0*
09
0>
0C
#551990000000
1!
1*
b101 6
19
1>
1C
b101 G
#552000000000
0!
0*
09
0>
0C
#552010000000
1!
1*
b110 6
19
1>
1C
b110 G
#552020000000
0!
0*
09
0>
0C
#552030000000
1!
1*
b111 6
19
1>
1C
b111 G
#552040000000
0!
0*
09
0>
0C
#552050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#552060000000
0!
0*
09
0>
0C
#552070000000
1!
1*
b1 6
19
1>
1C
b1 G
#552080000000
0!
0*
09
0>
0C
#552090000000
1!
1*
b10 6
19
1>
1C
b10 G
#552100000000
0!
0*
09
0>
0C
#552110000000
1!
1*
b11 6
19
1>
1C
b11 G
#552120000000
0!
0*
09
0>
0C
#552130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#552140000000
0!
0*
09
0>
0C
#552150000000
1!
1*
b101 6
19
1>
1C
b101 G
#552160000000
0!
0*
09
0>
0C
#552170000000
1!
1*
b110 6
19
1>
1C
b110 G
#552180000000
0!
0*
09
0>
0C
#552190000000
1!
1*
b111 6
19
1>
1C
b111 G
#552200000000
0!
1"
0*
1+
09
1:
0>
0C
#552210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#552220000000
0!
0*
09
0>
0C
#552230000000
1!
1*
b1 6
19
1>
1C
b1 G
#552240000000
0!
0*
09
0>
0C
#552250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#552260000000
0!
0*
09
0>
0C
#552270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#552280000000
0!
0*
09
0>
0C
#552290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#552300000000
0!
0*
09
0>
0C
#552310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#552320000000
0!
0#
0*
0,
09
0>
0?
0C
#552330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#552340000000
0!
0*
09
0>
0C
#552350000000
1!
1*
19
1>
1C
#552360000000
0!
0*
09
0>
0C
#552370000000
1!
1*
19
1>
1C
#552380000000
0!
0*
09
0>
0C
#552390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#552400000000
0!
0*
09
0>
0C
#552410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#552420000000
0!
0*
09
0>
0C
#552430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#552440000000
0!
0*
09
0>
0C
#552450000000
1!
1*
b10 6
19
1>
1C
b10 G
#552460000000
0!
0*
09
0>
0C
#552470000000
1!
1*
b11 6
19
1>
1C
b11 G
#552480000000
0!
0*
09
0>
0C
#552490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#552500000000
0!
0*
09
0>
0C
#552510000000
1!
1*
b101 6
19
1>
1C
b101 G
#552520000000
0!
0*
09
0>
0C
#552530000000
1!
1*
b110 6
19
1>
1C
b110 G
#552540000000
0!
0*
09
0>
0C
#552550000000
1!
1*
b111 6
19
1>
1C
b111 G
#552560000000
0!
0*
09
0>
0C
#552570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#552580000000
0!
0*
09
0>
0C
#552590000000
1!
1*
b1 6
19
1>
1C
b1 G
#552600000000
0!
0*
09
0>
0C
#552610000000
1!
1*
b10 6
19
1>
1C
b10 G
#552620000000
0!
0*
09
0>
0C
#552630000000
1!
1*
b11 6
19
1>
1C
b11 G
#552640000000
0!
0*
09
0>
0C
#552650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#552660000000
0!
0*
09
0>
0C
#552670000000
1!
1*
b101 6
19
1>
1C
b101 G
#552680000000
0!
0*
09
0>
0C
#552690000000
1!
1*
b110 6
19
1>
1C
b110 G
#552700000000
0!
0*
09
0>
0C
#552710000000
1!
1*
b111 6
19
1>
1C
b111 G
#552720000000
0!
0*
09
0>
0C
#552730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#552740000000
0!
0*
09
0>
0C
#552750000000
1!
1*
b1 6
19
1>
1C
b1 G
#552760000000
0!
0*
09
0>
0C
#552770000000
1!
1*
b10 6
19
1>
1C
b10 G
#552780000000
0!
0*
09
0>
0C
#552790000000
1!
1*
b11 6
19
1>
1C
b11 G
#552800000000
0!
0*
09
0>
0C
#552810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#552820000000
0!
0*
09
0>
0C
#552830000000
1!
1*
b101 6
19
1>
1C
b101 G
#552840000000
0!
0*
09
0>
0C
#552850000000
1!
1*
b110 6
19
1>
1C
b110 G
#552860000000
0!
0*
09
0>
0C
#552870000000
1!
1*
b111 6
19
1>
1C
b111 G
#552880000000
0!
1"
0*
1+
09
1:
0>
0C
#552890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#552900000000
0!
0*
09
0>
0C
#552910000000
1!
1*
b1 6
19
1>
1C
b1 G
#552920000000
0!
0*
09
0>
0C
#552930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#552940000000
0!
0*
09
0>
0C
#552950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#552960000000
0!
0*
09
0>
0C
#552970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#552980000000
0!
0*
09
0>
0C
#552990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#553000000000
0!
0#
0*
0,
09
0>
0?
0C
#553010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#553020000000
0!
0*
09
0>
0C
#553030000000
1!
1*
19
1>
1C
#553040000000
0!
0*
09
0>
0C
#553050000000
1!
1*
19
1>
1C
#553060000000
0!
0*
09
0>
0C
#553070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#553080000000
0!
0*
09
0>
0C
#553090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#553100000000
0!
0*
09
0>
0C
#553110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#553120000000
0!
0*
09
0>
0C
#553130000000
1!
1*
b10 6
19
1>
1C
b10 G
#553140000000
0!
0*
09
0>
0C
#553150000000
1!
1*
b11 6
19
1>
1C
b11 G
#553160000000
0!
0*
09
0>
0C
#553170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#553180000000
0!
0*
09
0>
0C
#553190000000
1!
1*
b101 6
19
1>
1C
b101 G
#553200000000
0!
0*
09
0>
0C
#553210000000
1!
1*
b110 6
19
1>
1C
b110 G
#553220000000
0!
0*
09
0>
0C
#553230000000
1!
1*
b111 6
19
1>
1C
b111 G
#553240000000
0!
0*
09
0>
0C
#553250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#553260000000
0!
0*
09
0>
0C
#553270000000
1!
1*
b1 6
19
1>
1C
b1 G
#553280000000
0!
0*
09
0>
0C
#553290000000
1!
1*
b10 6
19
1>
1C
b10 G
#553300000000
0!
0*
09
0>
0C
#553310000000
1!
1*
b11 6
19
1>
1C
b11 G
#553320000000
0!
0*
09
0>
0C
#553330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#553340000000
0!
0*
09
0>
0C
#553350000000
1!
1*
b101 6
19
1>
1C
b101 G
#553360000000
0!
0*
09
0>
0C
#553370000000
1!
1*
b110 6
19
1>
1C
b110 G
#553380000000
0!
0*
09
0>
0C
#553390000000
1!
1*
b111 6
19
1>
1C
b111 G
#553400000000
0!
0*
09
0>
0C
#553410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#553420000000
0!
0*
09
0>
0C
#553430000000
1!
1*
b1 6
19
1>
1C
b1 G
#553440000000
0!
0*
09
0>
0C
#553450000000
1!
1*
b10 6
19
1>
1C
b10 G
#553460000000
0!
0*
09
0>
0C
#553470000000
1!
1*
b11 6
19
1>
1C
b11 G
#553480000000
0!
0*
09
0>
0C
#553490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#553500000000
0!
0*
09
0>
0C
#553510000000
1!
1*
b101 6
19
1>
1C
b101 G
#553520000000
0!
0*
09
0>
0C
#553530000000
1!
1*
b110 6
19
1>
1C
b110 G
#553540000000
0!
0*
09
0>
0C
#553550000000
1!
1*
b111 6
19
1>
1C
b111 G
#553560000000
0!
1"
0*
1+
09
1:
0>
0C
#553570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#553580000000
0!
0*
09
0>
0C
#553590000000
1!
1*
b1 6
19
1>
1C
b1 G
#553600000000
0!
0*
09
0>
0C
#553610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#553620000000
0!
0*
09
0>
0C
#553630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#553640000000
0!
0*
09
0>
0C
#553650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#553660000000
0!
0*
09
0>
0C
#553670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#553680000000
0!
0#
0*
0,
09
0>
0?
0C
#553690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#553700000000
0!
0*
09
0>
0C
#553710000000
1!
1*
19
1>
1C
#553720000000
0!
0*
09
0>
0C
#553730000000
1!
1*
19
1>
1C
#553740000000
0!
0*
09
0>
0C
#553750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#553760000000
0!
0*
09
0>
0C
#553770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#553780000000
0!
0*
09
0>
0C
#553790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#553800000000
0!
0*
09
0>
0C
#553810000000
1!
1*
b10 6
19
1>
1C
b10 G
#553820000000
0!
0*
09
0>
0C
#553830000000
1!
1*
b11 6
19
1>
1C
b11 G
#553840000000
0!
0*
09
0>
0C
#553850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#553860000000
0!
0*
09
0>
0C
#553870000000
1!
1*
b101 6
19
1>
1C
b101 G
#553880000000
0!
0*
09
0>
0C
#553890000000
1!
1*
b110 6
19
1>
1C
b110 G
#553900000000
0!
0*
09
0>
0C
#553910000000
1!
1*
b111 6
19
1>
1C
b111 G
#553920000000
0!
0*
09
0>
0C
#553930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#553940000000
0!
0*
09
0>
0C
#553950000000
1!
1*
b1 6
19
1>
1C
b1 G
#553960000000
0!
0*
09
0>
0C
#553970000000
1!
1*
b10 6
19
1>
1C
b10 G
#553980000000
0!
0*
09
0>
0C
#553990000000
1!
1*
b11 6
19
1>
1C
b11 G
#554000000000
0!
0*
09
0>
0C
#554010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#554020000000
0!
0*
09
0>
0C
#554030000000
1!
1*
b101 6
19
1>
1C
b101 G
#554040000000
0!
0*
09
0>
0C
#554050000000
1!
1*
b110 6
19
1>
1C
b110 G
#554060000000
0!
0*
09
0>
0C
#554070000000
1!
1*
b111 6
19
1>
1C
b111 G
#554080000000
0!
0*
09
0>
0C
#554090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#554100000000
0!
0*
09
0>
0C
#554110000000
1!
1*
b1 6
19
1>
1C
b1 G
#554120000000
0!
0*
09
0>
0C
#554130000000
1!
1*
b10 6
19
1>
1C
b10 G
#554140000000
0!
0*
09
0>
0C
#554150000000
1!
1*
b11 6
19
1>
1C
b11 G
#554160000000
0!
0*
09
0>
0C
#554170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#554180000000
0!
0*
09
0>
0C
#554190000000
1!
1*
b101 6
19
1>
1C
b101 G
#554200000000
0!
0*
09
0>
0C
#554210000000
1!
1*
b110 6
19
1>
1C
b110 G
#554220000000
0!
0*
09
0>
0C
#554230000000
1!
1*
b111 6
19
1>
1C
b111 G
#554240000000
0!
1"
0*
1+
09
1:
0>
0C
#554250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#554260000000
0!
0*
09
0>
0C
#554270000000
1!
1*
b1 6
19
1>
1C
b1 G
#554280000000
0!
0*
09
0>
0C
#554290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#554300000000
0!
0*
09
0>
0C
#554310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#554320000000
0!
0*
09
0>
0C
#554330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#554340000000
0!
0*
09
0>
0C
#554350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#554360000000
0!
0#
0*
0,
09
0>
0?
0C
#554370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#554380000000
0!
0*
09
0>
0C
#554390000000
1!
1*
19
1>
1C
#554400000000
0!
0*
09
0>
0C
#554410000000
1!
1*
19
1>
1C
#554420000000
0!
0*
09
0>
0C
#554430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#554440000000
0!
0*
09
0>
0C
#554450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#554460000000
0!
0*
09
0>
0C
#554470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#554480000000
0!
0*
09
0>
0C
#554490000000
1!
1*
b10 6
19
1>
1C
b10 G
#554500000000
0!
0*
09
0>
0C
#554510000000
1!
1*
b11 6
19
1>
1C
b11 G
#554520000000
0!
0*
09
0>
0C
#554530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#554540000000
0!
0*
09
0>
0C
#554550000000
1!
1*
b101 6
19
1>
1C
b101 G
#554560000000
0!
0*
09
0>
0C
#554570000000
1!
1*
b110 6
19
1>
1C
b110 G
#554580000000
0!
0*
09
0>
0C
#554590000000
1!
1*
b111 6
19
1>
1C
b111 G
#554600000000
0!
0*
09
0>
0C
#554610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#554620000000
0!
0*
09
0>
0C
#554630000000
1!
1*
b1 6
19
1>
1C
b1 G
#554640000000
0!
0*
09
0>
0C
#554650000000
1!
1*
b10 6
19
1>
1C
b10 G
#554660000000
0!
0*
09
0>
0C
#554670000000
1!
1*
b11 6
19
1>
1C
b11 G
#554680000000
0!
0*
09
0>
0C
#554690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#554700000000
0!
0*
09
0>
0C
#554710000000
1!
1*
b101 6
19
1>
1C
b101 G
#554720000000
0!
0*
09
0>
0C
#554730000000
1!
1*
b110 6
19
1>
1C
b110 G
#554740000000
0!
0*
09
0>
0C
#554750000000
1!
1*
b111 6
19
1>
1C
b111 G
#554760000000
0!
0*
09
0>
0C
#554770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#554780000000
0!
0*
09
0>
0C
#554790000000
1!
1*
b1 6
19
1>
1C
b1 G
#554800000000
0!
0*
09
0>
0C
#554810000000
1!
1*
b10 6
19
1>
1C
b10 G
#554820000000
0!
0*
09
0>
0C
#554830000000
1!
1*
b11 6
19
1>
1C
b11 G
#554840000000
0!
0*
09
0>
0C
#554850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#554860000000
0!
0*
09
0>
0C
#554870000000
1!
1*
b101 6
19
1>
1C
b101 G
#554880000000
0!
0*
09
0>
0C
#554890000000
1!
1*
b110 6
19
1>
1C
b110 G
#554900000000
0!
0*
09
0>
0C
#554910000000
1!
1*
b111 6
19
1>
1C
b111 G
#554920000000
0!
1"
0*
1+
09
1:
0>
0C
#554930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#554940000000
0!
0*
09
0>
0C
#554950000000
1!
1*
b1 6
19
1>
1C
b1 G
#554960000000
0!
0*
09
0>
0C
#554970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#554980000000
0!
0*
09
0>
0C
#554990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#555000000000
0!
0*
09
0>
0C
#555010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#555020000000
0!
0*
09
0>
0C
#555030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#555040000000
0!
0#
0*
0,
09
0>
0?
0C
#555050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#555060000000
0!
0*
09
0>
0C
#555070000000
1!
1*
19
1>
1C
#555080000000
0!
0*
09
0>
0C
#555090000000
1!
1*
19
1>
1C
#555100000000
0!
0*
09
0>
0C
#555110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#555120000000
0!
0*
09
0>
0C
#555130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#555140000000
0!
0*
09
0>
0C
#555150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#555160000000
0!
0*
09
0>
0C
#555170000000
1!
1*
b10 6
19
1>
1C
b10 G
#555180000000
0!
0*
09
0>
0C
#555190000000
1!
1*
b11 6
19
1>
1C
b11 G
#555200000000
0!
0*
09
0>
0C
#555210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#555220000000
0!
0*
09
0>
0C
#555230000000
1!
1*
b101 6
19
1>
1C
b101 G
#555240000000
0!
0*
09
0>
0C
#555250000000
1!
1*
b110 6
19
1>
1C
b110 G
#555260000000
0!
0*
09
0>
0C
#555270000000
1!
1*
b111 6
19
1>
1C
b111 G
#555280000000
0!
0*
09
0>
0C
#555290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#555300000000
0!
0*
09
0>
0C
#555310000000
1!
1*
b1 6
19
1>
1C
b1 G
#555320000000
0!
0*
09
0>
0C
#555330000000
1!
1*
b10 6
19
1>
1C
b10 G
#555340000000
0!
0*
09
0>
0C
#555350000000
1!
1*
b11 6
19
1>
1C
b11 G
#555360000000
0!
0*
09
0>
0C
#555370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#555380000000
0!
0*
09
0>
0C
#555390000000
1!
1*
b101 6
19
1>
1C
b101 G
#555400000000
0!
0*
09
0>
0C
#555410000000
1!
1*
b110 6
19
1>
1C
b110 G
#555420000000
0!
0*
09
0>
0C
#555430000000
1!
1*
b111 6
19
1>
1C
b111 G
#555440000000
0!
0*
09
0>
0C
#555450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#555460000000
0!
0*
09
0>
0C
#555470000000
1!
1*
b1 6
19
1>
1C
b1 G
#555480000000
0!
0*
09
0>
0C
#555490000000
1!
1*
b10 6
19
1>
1C
b10 G
#555500000000
0!
0*
09
0>
0C
#555510000000
1!
1*
b11 6
19
1>
1C
b11 G
#555520000000
0!
0*
09
0>
0C
#555530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#555540000000
0!
0*
09
0>
0C
#555550000000
1!
1*
b101 6
19
1>
1C
b101 G
#555560000000
0!
0*
09
0>
0C
#555570000000
1!
1*
b110 6
19
1>
1C
b110 G
#555580000000
0!
0*
09
0>
0C
#555590000000
1!
1*
b111 6
19
1>
1C
b111 G
#555600000000
0!
1"
0*
1+
09
1:
0>
0C
#555610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#555620000000
0!
0*
09
0>
0C
#555630000000
1!
1*
b1 6
19
1>
1C
b1 G
#555640000000
0!
0*
09
0>
0C
#555650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#555660000000
0!
0*
09
0>
0C
#555670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#555680000000
0!
0*
09
0>
0C
#555690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#555700000000
0!
0*
09
0>
0C
#555710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#555720000000
0!
0#
0*
0,
09
0>
0?
0C
#555730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#555740000000
0!
0*
09
0>
0C
#555750000000
1!
1*
19
1>
1C
#555760000000
0!
0*
09
0>
0C
#555770000000
1!
1*
19
1>
1C
#555780000000
0!
0*
09
0>
0C
#555790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#555800000000
0!
0*
09
0>
0C
#555810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#555820000000
0!
0*
09
0>
0C
#555830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#555840000000
0!
0*
09
0>
0C
#555850000000
1!
1*
b10 6
19
1>
1C
b10 G
#555860000000
0!
0*
09
0>
0C
#555870000000
1!
1*
b11 6
19
1>
1C
b11 G
#555880000000
0!
0*
09
0>
0C
#555890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#555900000000
0!
0*
09
0>
0C
#555910000000
1!
1*
b101 6
19
1>
1C
b101 G
#555920000000
0!
0*
09
0>
0C
#555930000000
1!
1*
b110 6
19
1>
1C
b110 G
#555940000000
0!
0*
09
0>
0C
#555950000000
1!
1*
b111 6
19
1>
1C
b111 G
#555960000000
0!
0*
09
0>
0C
#555970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#555980000000
0!
0*
09
0>
0C
#555990000000
1!
1*
b1 6
19
1>
1C
b1 G
#556000000000
0!
0*
09
0>
0C
#556010000000
1!
1*
b10 6
19
1>
1C
b10 G
#556020000000
0!
0*
09
0>
0C
#556030000000
1!
1*
b11 6
19
1>
1C
b11 G
#556040000000
0!
0*
09
0>
0C
#556050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#556060000000
0!
0*
09
0>
0C
#556070000000
1!
1*
b101 6
19
1>
1C
b101 G
#556080000000
0!
0*
09
0>
0C
#556090000000
1!
1*
b110 6
19
1>
1C
b110 G
#556100000000
0!
0*
09
0>
0C
#556110000000
1!
1*
b111 6
19
1>
1C
b111 G
#556120000000
0!
0*
09
0>
0C
#556130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#556140000000
0!
0*
09
0>
0C
#556150000000
1!
1*
b1 6
19
1>
1C
b1 G
#556160000000
0!
0*
09
0>
0C
#556170000000
1!
1*
b10 6
19
1>
1C
b10 G
#556180000000
0!
0*
09
0>
0C
#556190000000
1!
1*
b11 6
19
1>
1C
b11 G
#556200000000
0!
0*
09
0>
0C
#556210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#556220000000
0!
0*
09
0>
0C
#556230000000
1!
1*
b101 6
19
1>
1C
b101 G
#556240000000
0!
0*
09
0>
0C
#556250000000
1!
1*
b110 6
19
1>
1C
b110 G
#556260000000
0!
0*
09
0>
0C
#556270000000
1!
1*
b111 6
19
1>
1C
b111 G
#556280000000
0!
1"
0*
1+
09
1:
0>
0C
#556290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#556300000000
0!
0*
09
0>
0C
#556310000000
1!
1*
b1 6
19
1>
1C
b1 G
#556320000000
0!
0*
09
0>
0C
#556330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#556340000000
0!
0*
09
0>
0C
#556350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#556360000000
0!
0*
09
0>
0C
#556370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#556380000000
0!
0*
09
0>
0C
#556390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#556400000000
0!
0#
0*
0,
09
0>
0?
0C
#556410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#556420000000
0!
0*
09
0>
0C
#556430000000
1!
1*
19
1>
1C
#556440000000
0!
0*
09
0>
0C
#556450000000
1!
1*
19
1>
1C
#556460000000
0!
0*
09
0>
0C
#556470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#556480000000
0!
0*
09
0>
0C
#556490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#556500000000
0!
0*
09
0>
0C
#556510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#556520000000
0!
0*
09
0>
0C
#556530000000
1!
1*
b10 6
19
1>
1C
b10 G
#556540000000
0!
0*
09
0>
0C
#556550000000
1!
1*
b11 6
19
1>
1C
b11 G
#556560000000
0!
0*
09
0>
0C
#556570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#556580000000
0!
0*
09
0>
0C
#556590000000
1!
1*
b101 6
19
1>
1C
b101 G
#556600000000
0!
0*
09
0>
0C
#556610000000
1!
1*
b110 6
19
1>
1C
b110 G
#556620000000
0!
0*
09
0>
0C
#556630000000
1!
1*
b111 6
19
1>
1C
b111 G
#556640000000
0!
0*
09
0>
0C
#556650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#556660000000
0!
0*
09
0>
0C
#556670000000
1!
1*
b1 6
19
1>
1C
b1 G
#556680000000
0!
0*
09
0>
0C
#556690000000
1!
1*
b10 6
19
1>
1C
b10 G
#556700000000
0!
0*
09
0>
0C
#556710000000
1!
1*
b11 6
19
1>
1C
b11 G
#556720000000
0!
0*
09
0>
0C
#556730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#556740000000
0!
0*
09
0>
0C
#556750000000
1!
1*
b101 6
19
1>
1C
b101 G
#556760000000
0!
0*
09
0>
0C
#556770000000
1!
1*
b110 6
19
1>
1C
b110 G
#556780000000
0!
0*
09
0>
0C
#556790000000
1!
1*
b111 6
19
1>
1C
b111 G
#556800000000
0!
0*
09
0>
0C
#556810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#556820000000
0!
0*
09
0>
0C
#556830000000
1!
1*
b1 6
19
1>
1C
b1 G
#556840000000
0!
0*
09
0>
0C
#556850000000
1!
1*
b10 6
19
1>
1C
b10 G
#556860000000
0!
0*
09
0>
0C
#556870000000
1!
1*
b11 6
19
1>
1C
b11 G
#556880000000
0!
0*
09
0>
0C
#556890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#556900000000
0!
0*
09
0>
0C
#556910000000
1!
1*
b101 6
19
1>
1C
b101 G
#556920000000
0!
0*
09
0>
0C
#556930000000
1!
1*
b110 6
19
1>
1C
b110 G
#556940000000
0!
0*
09
0>
0C
#556950000000
1!
1*
b111 6
19
1>
1C
b111 G
#556960000000
0!
1"
0*
1+
09
1:
0>
0C
#556970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#556980000000
0!
0*
09
0>
0C
#556990000000
1!
1*
b1 6
19
1>
1C
b1 G
#557000000000
0!
0*
09
0>
0C
#557010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#557020000000
0!
0*
09
0>
0C
#557030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#557040000000
0!
0*
09
0>
0C
#557050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#557060000000
0!
0*
09
0>
0C
#557070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#557080000000
0!
0#
0*
0,
09
0>
0?
0C
#557090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#557100000000
0!
0*
09
0>
0C
#557110000000
1!
1*
19
1>
1C
#557120000000
0!
0*
09
0>
0C
#557130000000
1!
1*
19
1>
1C
#557140000000
0!
0*
09
0>
0C
#557150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#557160000000
0!
0*
09
0>
0C
#557170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#557180000000
0!
0*
09
0>
0C
#557190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#557200000000
0!
0*
09
0>
0C
#557210000000
1!
1*
b10 6
19
1>
1C
b10 G
#557220000000
0!
0*
09
0>
0C
#557230000000
1!
1*
b11 6
19
1>
1C
b11 G
#557240000000
0!
0*
09
0>
0C
#557250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#557260000000
0!
0*
09
0>
0C
#557270000000
1!
1*
b101 6
19
1>
1C
b101 G
#557280000000
0!
0*
09
0>
0C
#557290000000
1!
1*
b110 6
19
1>
1C
b110 G
#557300000000
0!
0*
09
0>
0C
#557310000000
1!
1*
b111 6
19
1>
1C
b111 G
#557320000000
0!
0*
09
0>
0C
#557330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#557340000000
0!
0*
09
0>
0C
#557350000000
1!
1*
b1 6
19
1>
1C
b1 G
#557360000000
0!
0*
09
0>
0C
#557370000000
1!
1*
b10 6
19
1>
1C
b10 G
#557380000000
0!
0*
09
0>
0C
#557390000000
1!
1*
b11 6
19
1>
1C
b11 G
#557400000000
0!
0*
09
0>
0C
#557410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#557420000000
0!
0*
09
0>
0C
#557430000000
1!
1*
b101 6
19
1>
1C
b101 G
#557440000000
0!
0*
09
0>
0C
#557450000000
1!
1*
b110 6
19
1>
1C
b110 G
#557460000000
0!
0*
09
0>
0C
#557470000000
1!
1*
b111 6
19
1>
1C
b111 G
#557480000000
0!
0*
09
0>
0C
#557490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#557500000000
0!
0*
09
0>
0C
#557510000000
1!
1*
b1 6
19
1>
1C
b1 G
#557520000000
0!
0*
09
0>
0C
#557530000000
1!
1*
b10 6
19
1>
1C
b10 G
#557540000000
0!
0*
09
0>
0C
#557550000000
1!
1*
b11 6
19
1>
1C
b11 G
#557560000000
0!
0*
09
0>
0C
#557570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#557580000000
0!
0*
09
0>
0C
#557590000000
1!
1*
b101 6
19
1>
1C
b101 G
#557600000000
0!
0*
09
0>
0C
#557610000000
1!
1*
b110 6
19
1>
1C
b110 G
#557620000000
0!
0*
09
0>
0C
#557630000000
1!
1*
b111 6
19
1>
1C
b111 G
#557640000000
0!
1"
0*
1+
09
1:
0>
0C
#557650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#557660000000
0!
0*
09
0>
0C
#557670000000
1!
1*
b1 6
19
1>
1C
b1 G
#557680000000
0!
0*
09
0>
0C
#557690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#557700000000
0!
0*
09
0>
0C
#557710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#557720000000
0!
0*
09
0>
0C
#557730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#557740000000
0!
0*
09
0>
0C
#557750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#557760000000
0!
0#
0*
0,
09
0>
0?
0C
#557770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#557780000000
0!
0*
09
0>
0C
#557790000000
1!
1*
19
1>
1C
#557800000000
0!
0*
09
0>
0C
#557810000000
1!
1*
19
1>
1C
#557820000000
0!
0*
09
0>
0C
#557830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#557840000000
0!
0*
09
0>
0C
#557850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#557860000000
0!
0*
09
0>
0C
#557870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#557880000000
0!
0*
09
0>
0C
#557890000000
1!
1*
b10 6
19
1>
1C
b10 G
#557900000000
0!
0*
09
0>
0C
#557910000000
1!
1*
b11 6
19
1>
1C
b11 G
#557920000000
0!
0*
09
0>
0C
#557930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#557940000000
0!
0*
09
0>
0C
#557950000000
1!
1*
b101 6
19
1>
1C
b101 G
#557960000000
0!
0*
09
0>
0C
#557970000000
1!
1*
b110 6
19
1>
1C
b110 G
#557980000000
0!
0*
09
0>
0C
#557990000000
1!
1*
b111 6
19
1>
1C
b111 G
#558000000000
0!
0*
09
0>
0C
#558010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#558020000000
0!
0*
09
0>
0C
#558030000000
1!
1*
b1 6
19
1>
1C
b1 G
#558040000000
0!
0*
09
0>
0C
#558050000000
1!
1*
b10 6
19
1>
1C
b10 G
#558060000000
0!
0*
09
0>
0C
#558070000000
1!
1*
b11 6
19
1>
1C
b11 G
#558080000000
0!
0*
09
0>
0C
#558090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#558100000000
0!
0*
09
0>
0C
#558110000000
1!
1*
b101 6
19
1>
1C
b101 G
#558120000000
0!
0*
09
0>
0C
#558130000000
1!
1*
b110 6
19
1>
1C
b110 G
#558140000000
0!
0*
09
0>
0C
#558150000000
1!
1*
b111 6
19
1>
1C
b111 G
#558160000000
0!
0*
09
0>
0C
#558170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#558180000000
0!
0*
09
0>
0C
#558190000000
1!
1*
b1 6
19
1>
1C
b1 G
#558200000000
0!
0*
09
0>
0C
#558210000000
1!
1*
b10 6
19
1>
1C
b10 G
#558220000000
0!
0*
09
0>
0C
#558230000000
1!
1*
b11 6
19
1>
1C
b11 G
#558240000000
0!
0*
09
0>
0C
#558250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#558260000000
0!
0*
09
0>
0C
#558270000000
1!
1*
b101 6
19
1>
1C
b101 G
#558280000000
0!
0*
09
0>
0C
#558290000000
1!
1*
b110 6
19
1>
1C
b110 G
#558300000000
0!
0*
09
0>
0C
#558310000000
1!
1*
b111 6
19
1>
1C
b111 G
#558320000000
0!
1"
0*
1+
09
1:
0>
0C
#558330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#558340000000
0!
0*
09
0>
0C
#558350000000
1!
1*
b1 6
19
1>
1C
b1 G
#558360000000
0!
0*
09
0>
0C
#558370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#558380000000
0!
0*
09
0>
0C
#558390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#558400000000
0!
0*
09
0>
0C
#558410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#558420000000
0!
0*
09
0>
0C
#558430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#558440000000
0!
0#
0*
0,
09
0>
0?
0C
#558450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#558460000000
0!
0*
09
0>
0C
#558470000000
1!
1*
19
1>
1C
#558480000000
0!
0*
09
0>
0C
#558490000000
1!
1*
19
1>
1C
#558500000000
0!
0*
09
0>
0C
#558510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#558520000000
0!
0*
09
0>
0C
#558530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#558540000000
0!
0*
09
0>
0C
#558550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#558560000000
0!
0*
09
0>
0C
#558570000000
1!
1*
b10 6
19
1>
1C
b10 G
#558580000000
0!
0*
09
0>
0C
#558590000000
1!
1*
b11 6
19
1>
1C
b11 G
#558600000000
0!
0*
09
0>
0C
#558610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#558620000000
0!
0*
09
0>
0C
#558630000000
1!
1*
b101 6
19
1>
1C
b101 G
#558640000000
0!
0*
09
0>
0C
#558650000000
1!
1*
b110 6
19
1>
1C
b110 G
#558660000000
0!
0*
09
0>
0C
#558670000000
1!
1*
b111 6
19
1>
1C
b111 G
#558680000000
0!
0*
09
0>
0C
#558690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#558700000000
0!
0*
09
0>
0C
#558710000000
1!
1*
b1 6
19
1>
1C
b1 G
#558720000000
0!
0*
09
0>
0C
#558730000000
1!
1*
b10 6
19
1>
1C
b10 G
#558740000000
0!
0*
09
0>
0C
#558750000000
1!
1*
b11 6
19
1>
1C
b11 G
#558760000000
0!
0*
09
0>
0C
#558770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#558780000000
0!
0*
09
0>
0C
#558790000000
1!
1*
b101 6
19
1>
1C
b101 G
#558800000000
0!
0*
09
0>
0C
#558810000000
1!
1*
b110 6
19
1>
1C
b110 G
#558820000000
0!
0*
09
0>
0C
#558830000000
1!
1*
b111 6
19
1>
1C
b111 G
#558840000000
0!
0*
09
0>
0C
#558850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#558860000000
0!
0*
09
0>
0C
#558870000000
1!
1*
b1 6
19
1>
1C
b1 G
#558880000000
0!
0*
09
0>
0C
#558890000000
1!
1*
b10 6
19
1>
1C
b10 G
#558900000000
0!
0*
09
0>
0C
#558910000000
1!
1*
b11 6
19
1>
1C
b11 G
#558920000000
0!
0*
09
0>
0C
#558930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#558940000000
0!
0*
09
0>
0C
#558950000000
1!
1*
b101 6
19
1>
1C
b101 G
#558960000000
0!
0*
09
0>
0C
#558970000000
1!
1*
b110 6
19
1>
1C
b110 G
#558980000000
0!
0*
09
0>
0C
#558990000000
1!
1*
b111 6
19
1>
1C
b111 G
#559000000000
0!
1"
0*
1+
09
1:
0>
0C
#559010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#559020000000
0!
0*
09
0>
0C
#559030000000
1!
1*
b1 6
19
1>
1C
b1 G
#559040000000
0!
0*
09
0>
0C
#559050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#559060000000
0!
0*
09
0>
0C
#559070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#559080000000
0!
0*
09
0>
0C
#559090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#559100000000
0!
0*
09
0>
0C
#559110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#559120000000
0!
0#
0*
0,
09
0>
0?
0C
#559130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#559140000000
0!
0*
09
0>
0C
#559150000000
1!
1*
19
1>
1C
#559160000000
0!
0*
09
0>
0C
#559170000000
1!
1*
19
1>
1C
#559180000000
0!
0*
09
0>
0C
#559190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#559200000000
0!
0*
09
0>
0C
#559210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#559220000000
0!
0*
09
0>
0C
#559230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#559240000000
0!
0*
09
0>
0C
#559250000000
1!
1*
b10 6
19
1>
1C
b10 G
#559260000000
0!
0*
09
0>
0C
#559270000000
1!
1*
b11 6
19
1>
1C
b11 G
#559280000000
0!
0*
09
0>
0C
#559290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#559300000000
0!
0*
09
0>
0C
#559310000000
1!
1*
b101 6
19
1>
1C
b101 G
#559320000000
0!
0*
09
0>
0C
#559330000000
1!
1*
b110 6
19
1>
1C
b110 G
#559340000000
0!
0*
09
0>
0C
#559350000000
1!
1*
b111 6
19
1>
1C
b111 G
#559360000000
0!
0*
09
0>
0C
#559370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#559380000000
0!
0*
09
0>
0C
#559390000000
1!
1*
b1 6
19
1>
1C
b1 G
#559400000000
0!
0*
09
0>
0C
#559410000000
1!
1*
b10 6
19
1>
1C
b10 G
#559420000000
0!
0*
09
0>
0C
#559430000000
1!
1*
b11 6
19
1>
1C
b11 G
#559440000000
0!
0*
09
0>
0C
#559450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#559460000000
0!
0*
09
0>
0C
#559470000000
1!
1*
b101 6
19
1>
1C
b101 G
#559480000000
0!
0*
09
0>
0C
#559490000000
1!
1*
b110 6
19
1>
1C
b110 G
#559500000000
0!
0*
09
0>
0C
#559510000000
1!
1*
b111 6
19
1>
1C
b111 G
#559520000000
0!
0*
09
0>
0C
#559530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#559540000000
0!
0*
09
0>
0C
#559550000000
1!
1*
b1 6
19
1>
1C
b1 G
#559560000000
0!
0*
09
0>
0C
#559570000000
1!
1*
b10 6
19
1>
1C
b10 G
#559580000000
0!
0*
09
0>
0C
#559590000000
1!
1*
b11 6
19
1>
1C
b11 G
#559600000000
0!
0*
09
0>
0C
#559610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#559620000000
0!
0*
09
0>
0C
#559630000000
1!
1*
b101 6
19
1>
1C
b101 G
#559640000000
0!
0*
09
0>
0C
#559650000000
1!
1*
b110 6
19
1>
1C
b110 G
#559660000000
0!
0*
09
0>
0C
#559670000000
1!
1*
b111 6
19
1>
1C
b111 G
#559680000000
0!
1"
0*
1+
09
1:
0>
0C
#559690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#559700000000
0!
0*
09
0>
0C
#559710000000
1!
1*
b1 6
19
1>
1C
b1 G
#559720000000
0!
0*
09
0>
0C
#559730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#559740000000
0!
0*
09
0>
0C
#559750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#559760000000
0!
0*
09
0>
0C
#559770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#559780000000
0!
0*
09
0>
0C
#559790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#559800000000
0!
0#
0*
0,
09
0>
0?
0C
#559810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#559820000000
0!
0*
09
0>
0C
#559830000000
1!
1*
19
1>
1C
#559840000000
0!
0*
09
0>
0C
#559850000000
1!
1*
19
1>
1C
#559860000000
0!
0*
09
0>
0C
#559870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#559880000000
0!
0*
09
0>
0C
#559890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#559900000000
0!
0*
09
0>
0C
#559910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#559920000000
0!
0*
09
0>
0C
#559930000000
1!
1*
b10 6
19
1>
1C
b10 G
#559940000000
0!
0*
09
0>
0C
#559950000000
1!
1*
b11 6
19
1>
1C
b11 G
#559960000000
0!
0*
09
0>
0C
#559970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#559980000000
0!
0*
09
0>
0C
#559990000000
1!
1*
b101 6
19
1>
1C
b101 G
#560000000000
0!
0*
09
0>
0C
#560010000000
1!
1*
b110 6
19
1>
1C
b110 G
#560020000000
0!
0*
09
0>
0C
#560030000000
1!
1*
b111 6
19
1>
1C
b111 G
#560040000000
0!
0*
09
0>
0C
#560050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#560060000000
0!
0*
09
0>
0C
#560070000000
1!
1*
b1 6
19
1>
1C
b1 G
#560080000000
0!
0*
09
0>
0C
#560090000000
1!
1*
b10 6
19
1>
1C
b10 G
#560100000000
0!
0*
09
0>
0C
#560110000000
1!
1*
b11 6
19
1>
1C
b11 G
#560120000000
0!
0*
09
0>
0C
#560130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#560140000000
0!
0*
09
0>
0C
#560150000000
1!
1*
b101 6
19
1>
1C
b101 G
#560160000000
0!
0*
09
0>
0C
#560170000000
1!
1*
b110 6
19
1>
1C
b110 G
#560180000000
0!
0*
09
0>
0C
#560190000000
1!
1*
b111 6
19
1>
1C
b111 G
#560200000000
0!
0*
09
0>
0C
#560210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#560220000000
0!
0*
09
0>
0C
#560230000000
1!
1*
b1 6
19
1>
1C
b1 G
#560240000000
0!
0*
09
0>
0C
#560250000000
1!
1*
b10 6
19
1>
1C
b10 G
#560260000000
0!
0*
09
0>
0C
#560270000000
1!
1*
b11 6
19
1>
1C
b11 G
#560280000000
0!
0*
09
0>
0C
#560290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#560300000000
0!
0*
09
0>
0C
#560310000000
1!
1*
b101 6
19
1>
1C
b101 G
#560320000000
0!
0*
09
0>
0C
#560330000000
1!
1*
b110 6
19
1>
1C
b110 G
#560340000000
0!
0*
09
0>
0C
#560350000000
1!
1*
b111 6
19
1>
1C
b111 G
#560360000000
0!
1"
0*
1+
09
1:
0>
0C
#560370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#560380000000
0!
0*
09
0>
0C
#560390000000
1!
1*
b1 6
19
1>
1C
b1 G
#560400000000
0!
0*
09
0>
0C
#560410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#560420000000
0!
0*
09
0>
0C
#560430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#560440000000
0!
0*
09
0>
0C
#560450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#560460000000
0!
0*
09
0>
0C
#560470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#560480000000
0!
0#
0*
0,
09
0>
0?
0C
#560490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#560500000000
0!
0*
09
0>
0C
#560510000000
1!
1*
19
1>
1C
#560520000000
0!
0*
09
0>
0C
#560530000000
1!
1*
19
1>
1C
#560540000000
0!
0*
09
0>
0C
#560550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#560560000000
0!
0*
09
0>
0C
#560570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#560580000000
0!
0*
09
0>
0C
#560590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#560600000000
0!
0*
09
0>
0C
#560610000000
1!
1*
b10 6
19
1>
1C
b10 G
#560620000000
0!
0*
09
0>
0C
#560630000000
1!
1*
b11 6
19
1>
1C
b11 G
#560640000000
0!
0*
09
0>
0C
#560650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#560660000000
0!
0*
09
0>
0C
#560670000000
1!
1*
b101 6
19
1>
1C
b101 G
#560680000000
0!
0*
09
0>
0C
#560690000000
1!
1*
b110 6
19
1>
1C
b110 G
#560700000000
0!
0*
09
0>
0C
#560710000000
1!
1*
b111 6
19
1>
1C
b111 G
#560720000000
0!
0*
09
0>
0C
#560730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#560740000000
0!
0*
09
0>
0C
#560750000000
1!
1*
b1 6
19
1>
1C
b1 G
#560760000000
0!
0*
09
0>
0C
#560770000000
1!
1*
b10 6
19
1>
1C
b10 G
#560780000000
0!
0*
09
0>
0C
#560790000000
1!
1*
b11 6
19
1>
1C
b11 G
#560800000000
0!
0*
09
0>
0C
#560810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#560820000000
0!
0*
09
0>
0C
#560830000000
1!
1*
b101 6
19
1>
1C
b101 G
#560840000000
0!
0*
09
0>
0C
#560850000000
1!
1*
b110 6
19
1>
1C
b110 G
#560860000000
0!
0*
09
0>
0C
#560870000000
1!
1*
b111 6
19
1>
1C
b111 G
#560880000000
0!
0*
09
0>
0C
#560890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#560900000000
0!
0*
09
0>
0C
#560910000000
1!
1*
b1 6
19
1>
1C
b1 G
#560920000000
0!
0*
09
0>
0C
#560930000000
1!
1*
b10 6
19
1>
1C
b10 G
#560940000000
0!
0*
09
0>
0C
#560950000000
1!
1*
b11 6
19
1>
1C
b11 G
#560960000000
0!
0*
09
0>
0C
#560970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#560980000000
0!
0*
09
0>
0C
#560990000000
1!
1*
b101 6
19
1>
1C
b101 G
#561000000000
0!
0*
09
0>
0C
#561010000000
1!
1*
b110 6
19
1>
1C
b110 G
#561020000000
0!
0*
09
0>
0C
#561030000000
1!
1*
b111 6
19
1>
1C
b111 G
#561040000000
0!
1"
0*
1+
09
1:
0>
0C
#561050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#561060000000
0!
0*
09
0>
0C
#561070000000
1!
1*
b1 6
19
1>
1C
b1 G
#561080000000
0!
0*
09
0>
0C
#561090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#561100000000
0!
0*
09
0>
0C
#561110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#561120000000
0!
0*
09
0>
0C
#561130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#561140000000
0!
0*
09
0>
0C
#561150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#561160000000
0!
0#
0*
0,
09
0>
0?
0C
#561170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#561180000000
0!
0*
09
0>
0C
#561190000000
1!
1*
19
1>
1C
#561200000000
0!
0*
09
0>
0C
#561210000000
1!
1*
19
1>
1C
#561220000000
0!
0*
09
0>
0C
#561230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#561240000000
0!
0*
09
0>
0C
#561250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#561260000000
0!
0*
09
0>
0C
#561270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#561280000000
0!
0*
09
0>
0C
#561290000000
1!
1*
b10 6
19
1>
1C
b10 G
#561300000000
0!
0*
09
0>
0C
#561310000000
1!
1*
b11 6
19
1>
1C
b11 G
#561320000000
0!
0*
09
0>
0C
#561330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#561340000000
0!
0*
09
0>
0C
#561350000000
1!
1*
b101 6
19
1>
1C
b101 G
#561360000000
0!
0*
09
0>
0C
#561370000000
1!
1*
b110 6
19
1>
1C
b110 G
#561380000000
0!
0*
09
0>
0C
#561390000000
1!
1*
b111 6
19
1>
1C
b111 G
#561400000000
0!
0*
09
0>
0C
#561410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#561420000000
0!
0*
09
0>
0C
#561430000000
1!
1*
b1 6
19
1>
1C
b1 G
#561440000000
0!
0*
09
0>
0C
#561450000000
1!
1*
b10 6
19
1>
1C
b10 G
#561460000000
0!
0*
09
0>
0C
#561470000000
1!
1*
b11 6
19
1>
1C
b11 G
#561480000000
0!
0*
09
0>
0C
#561490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#561500000000
0!
0*
09
0>
0C
#561510000000
1!
1*
b101 6
19
1>
1C
b101 G
#561520000000
0!
0*
09
0>
0C
#561530000000
1!
1*
b110 6
19
1>
1C
b110 G
#561540000000
0!
0*
09
0>
0C
#561550000000
1!
1*
b111 6
19
1>
1C
b111 G
#561560000000
0!
0*
09
0>
0C
#561570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#561580000000
0!
0*
09
0>
0C
#561590000000
1!
1*
b1 6
19
1>
1C
b1 G
#561600000000
0!
0*
09
0>
0C
#561610000000
1!
1*
b10 6
19
1>
1C
b10 G
#561620000000
0!
0*
09
0>
0C
#561630000000
1!
1*
b11 6
19
1>
1C
b11 G
#561640000000
0!
0*
09
0>
0C
#561650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#561660000000
0!
0*
09
0>
0C
#561670000000
1!
1*
b101 6
19
1>
1C
b101 G
#561680000000
0!
0*
09
0>
0C
#561690000000
1!
1*
b110 6
19
1>
1C
b110 G
#561700000000
0!
0*
09
0>
0C
#561710000000
1!
1*
b111 6
19
1>
1C
b111 G
#561720000000
0!
1"
0*
1+
09
1:
0>
0C
#561730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#561740000000
0!
0*
09
0>
0C
#561750000000
1!
1*
b1 6
19
1>
1C
b1 G
#561760000000
0!
0*
09
0>
0C
#561770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#561780000000
0!
0*
09
0>
0C
#561790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#561800000000
0!
0*
09
0>
0C
#561810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#561820000000
0!
0*
09
0>
0C
#561830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#561840000000
0!
0#
0*
0,
09
0>
0?
0C
#561850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#561860000000
0!
0*
09
0>
0C
#561870000000
1!
1*
19
1>
1C
#561880000000
0!
0*
09
0>
0C
#561890000000
1!
1*
19
1>
1C
#561900000000
0!
0*
09
0>
0C
#561910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#561920000000
0!
0*
09
0>
0C
#561930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#561940000000
0!
0*
09
0>
0C
#561950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#561960000000
0!
0*
09
0>
0C
#561970000000
1!
1*
b10 6
19
1>
1C
b10 G
#561980000000
0!
0*
09
0>
0C
#561990000000
1!
1*
b11 6
19
1>
1C
b11 G
#562000000000
0!
0*
09
0>
0C
#562010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#562020000000
0!
0*
09
0>
0C
#562030000000
1!
1*
b101 6
19
1>
1C
b101 G
#562040000000
0!
0*
09
0>
0C
#562050000000
1!
1*
b110 6
19
1>
1C
b110 G
#562060000000
0!
0*
09
0>
0C
#562070000000
1!
1*
b111 6
19
1>
1C
b111 G
#562080000000
0!
0*
09
0>
0C
#562090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#562100000000
0!
0*
09
0>
0C
#562110000000
1!
1*
b1 6
19
1>
1C
b1 G
#562120000000
0!
0*
09
0>
0C
#562130000000
1!
1*
b10 6
19
1>
1C
b10 G
#562140000000
0!
0*
09
0>
0C
#562150000000
1!
1*
b11 6
19
1>
1C
b11 G
#562160000000
0!
0*
09
0>
0C
#562170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#562180000000
0!
0*
09
0>
0C
#562190000000
1!
1*
b101 6
19
1>
1C
b101 G
#562200000000
0!
0*
09
0>
0C
#562210000000
1!
1*
b110 6
19
1>
1C
b110 G
#562220000000
0!
0*
09
0>
0C
#562230000000
1!
1*
b111 6
19
1>
1C
b111 G
#562240000000
0!
0*
09
0>
0C
#562250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#562260000000
0!
0*
09
0>
0C
#562270000000
1!
1*
b1 6
19
1>
1C
b1 G
#562280000000
0!
0*
09
0>
0C
#562290000000
1!
1*
b10 6
19
1>
1C
b10 G
#562300000000
0!
0*
09
0>
0C
#562310000000
1!
1*
b11 6
19
1>
1C
b11 G
#562320000000
0!
0*
09
0>
0C
#562330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#562340000000
0!
0*
09
0>
0C
#562350000000
1!
1*
b101 6
19
1>
1C
b101 G
#562360000000
0!
0*
09
0>
0C
#562370000000
1!
1*
b110 6
19
1>
1C
b110 G
#562380000000
0!
0*
09
0>
0C
#562390000000
1!
1*
b111 6
19
1>
1C
b111 G
#562400000000
0!
1"
0*
1+
09
1:
0>
0C
#562410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#562420000000
0!
0*
09
0>
0C
#562430000000
1!
1*
b1 6
19
1>
1C
b1 G
#562440000000
0!
0*
09
0>
0C
#562450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#562460000000
0!
0*
09
0>
0C
#562470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#562480000000
0!
0*
09
0>
0C
#562490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#562500000000
0!
0*
09
0>
0C
#562510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#562520000000
0!
0#
0*
0,
09
0>
0?
0C
#562530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#562540000000
0!
0*
09
0>
0C
#562550000000
1!
1*
19
1>
1C
#562560000000
0!
0*
09
0>
0C
#562570000000
1!
1*
19
1>
1C
#562580000000
0!
0*
09
0>
0C
#562590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#562600000000
0!
0*
09
0>
0C
#562610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#562620000000
0!
0*
09
0>
0C
#562630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#562640000000
0!
0*
09
0>
0C
#562650000000
1!
1*
b10 6
19
1>
1C
b10 G
#562660000000
0!
0*
09
0>
0C
#562670000000
1!
1*
b11 6
19
1>
1C
b11 G
#562680000000
0!
0*
09
0>
0C
#562690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#562700000000
0!
0*
09
0>
0C
#562710000000
1!
1*
b101 6
19
1>
1C
b101 G
#562720000000
0!
0*
09
0>
0C
#562730000000
1!
1*
b110 6
19
1>
1C
b110 G
#562740000000
0!
0*
09
0>
0C
#562750000000
1!
1*
b111 6
19
1>
1C
b111 G
#562760000000
0!
0*
09
0>
0C
#562770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#562780000000
0!
0*
09
0>
0C
#562790000000
1!
1*
b1 6
19
1>
1C
b1 G
#562800000000
0!
0*
09
0>
0C
#562810000000
1!
1*
b10 6
19
1>
1C
b10 G
#562820000000
0!
0*
09
0>
0C
#562830000000
1!
1*
b11 6
19
1>
1C
b11 G
#562840000000
0!
0*
09
0>
0C
#562850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#562860000000
0!
0*
09
0>
0C
#562870000000
1!
1*
b101 6
19
1>
1C
b101 G
#562880000000
0!
0*
09
0>
0C
#562890000000
1!
1*
b110 6
19
1>
1C
b110 G
#562900000000
0!
0*
09
0>
0C
#562910000000
1!
1*
b111 6
19
1>
1C
b111 G
#562920000000
0!
0*
09
0>
0C
#562930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#562940000000
0!
0*
09
0>
0C
#562950000000
1!
1*
b1 6
19
1>
1C
b1 G
#562960000000
0!
0*
09
0>
0C
#562970000000
1!
1*
b10 6
19
1>
1C
b10 G
#562980000000
0!
0*
09
0>
0C
#562990000000
1!
1*
b11 6
19
1>
1C
b11 G
#563000000000
0!
0*
09
0>
0C
#563010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#563020000000
0!
0*
09
0>
0C
#563030000000
1!
1*
b101 6
19
1>
1C
b101 G
#563040000000
0!
0*
09
0>
0C
#563050000000
1!
1*
b110 6
19
1>
1C
b110 G
#563060000000
0!
0*
09
0>
0C
#563070000000
1!
1*
b111 6
19
1>
1C
b111 G
#563080000000
0!
1"
0*
1+
09
1:
0>
0C
#563090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#563100000000
0!
0*
09
0>
0C
#563110000000
1!
1*
b1 6
19
1>
1C
b1 G
#563120000000
0!
0*
09
0>
0C
#563130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#563140000000
0!
0*
09
0>
0C
#563150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#563160000000
0!
0*
09
0>
0C
#563170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#563180000000
0!
0*
09
0>
0C
#563190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#563200000000
0!
0#
0*
0,
09
0>
0?
0C
#563210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#563220000000
0!
0*
09
0>
0C
#563230000000
1!
1*
19
1>
1C
#563240000000
0!
0*
09
0>
0C
#563250000000
1!
1*
19
1>
1C
#563260000000
0!
0*
09
0>
0C
#563270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#563280000000
0!
0*
09
0>
0C
#563290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#563300000000
0!
0*
09
0>
0C
#563310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#563320000000
0!
0*
09
0>
0C
#563330000000
1!
1*
b10 6
19
1>
1C
b10 G
#563340000000
0!
0*
09
0>
0C
#563350000000
1!
1*
b11 6
19
1>
1C
b11 G
#563360000000
0!
0*
09
0>
0C
#563370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#563380000000
0!
0*
09
0>
0C
#563390000000
1!
1*
b101 6
19
1>
1C
b101 G
#563400000000
0!
0*
09
0>
0C
#563410000000
1!
1*
b110 6
19
1>
1C
b110 G
#563420000000
0!
0*
09
0>
0C
#563430000000
1!
1*
b111 6
19
1>
1C
b111 G
#563440000000
0!
0*
09
0>
0C
#563450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#563460000000
0!
0*
09
0>
0C
#563470000000
1!
1*
b1 6
19
1>
1C
b1 G
#563480000000
0!
0*
09
0>
0C
#563490000000
1!
1*
b10 6
19
1>
1C
b10 G
#563500000000
0!
0*
09
0>
0C
#563510000000
1!
1*
b11 6
19
1>
1C
b11 G
#563520000000
0!
0*
09
0>
0C
#563530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#563540000000
0!
0*
09
0>
0C
#563550000000
1!
1*
b101 6
19
1>
1C
b101 G
#563560000000
0!
0*
09
0>
0C
#563570000000
1!
1*
b110 6
19
1>
1C
b110 G
#563580000000
0!
0*
09
0>
0C
#563590000000
1!
1*
b111 6
19
1>
1C
b111 G
#563600000000
0!
0*
09
0>
0C
#563610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#563620000000
0!
0*
09
0>
0C
#563630000000
1!
1*
b1 6
19
1>
1C
b1 G
#563640000000
0!
0*
09
0>
0C
#563650000000
1!
1*
b10 6
19
1>
1C
b10 G
#563660000000
0!
0*
09
0>
0C
#563670000000
1!
1*
b11 6
19
1>
1C
b11 G
#563680000000
0!
0*
09
0>
0C
#563690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#563700000000
0!
0*
09
0>
0C
#563710000000
1!
1*
b101 6
19
1>
1C
b101 G
#563720000000
0!
0*
09
0>
0C
#563730000000
1!
1*
b110 6
19
1>
1C
b110 G
#563740000000
0!
0*
09
0>
0C
#563750000000
1!
1*
b111 6
19
1>
1C
b111 G
#563760000000
0!
1"
0*
1+
09
1:
0>
0C
#563770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#563780000000
0!
0*
09
0>
0C
#563790000000
1!
1*
b1 6
19
1>
1C
b1 G
#563800000000
0!
0*
09
0>
0C
#563810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#563820000000
0!
0*
09
0>
0C
#563830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#563840000000
0!
0*
09
0>
0C
#563850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#563860000000
0!
0*
09
0>
0C
#563870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#563880000000
0!
0#
0*
0,
09
0>
0?
0C
#563890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#563900000000
0!
0*
09
0>
0C
#563910000000
1!
1*
19
1>
1C
#563920000000
0!
0*
09
0>
0C
#563930000000
1!
1*
19
1>
1C
#563940000000
0!
0*
09
0>
0C
#563950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#563960000000
0!
0*
09
0>
0C
#563970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#563980000000
0!
0*
09
0>
0C
#563990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#564000000000
0!
0*
09
0>
0C
#564010000000
1!
1*
b10 6
19
1>
1C
b10 G
#564020000000
0!
0*
09
0>
0C
#564030000000
1!
1*
b11 6
19
1>
1C
b11 G
#564040000000
0!
0*
09
0>
0C
#564050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#564060000000
0!
0*
09
0>
0C
#564070000000
1!
1*
b101 6
19
1>
1C
b101 G
#564080000000
0!
0*
09
0>
0C
#564090000000
1!
1*
b110 6
19
1>
1C
b110 G
#564100000000
0!
0*
09
0>
0C
#564110000000
1!
1*
b111 6
19
1>
1C
b111 G
#564120000000
0!
0*
09
0>
0C
#564130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#564140000000
0!
0*
09
0>
0C
#564150000000
1!
1*
b1 6
19
1>
1C
b1 G
#564160000000
0!
0*
09
0>
0C
#564170000000
1!
1*
b10 6
19
1>
1C
b10 G
#564180000000
0!
0*
09
0>
0C
#564190000000
1!
1*
b11 6
19
1>
1C
b11 G
#564200000000
0!
0*
09
0>
0C
#564210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#564220000000
0!
0*
09
0>
0C
#564230000000
1!
1*
b101 6
19
1>
1C
b101 G
#564240000000
0!
0*
09
0>
0C
#564250000000
1!
1*
b110 6
19
1>
1C
b110 G
#564260000000
0!
0*
09
0>
0C
#564270000000
1!
1*
b111 6
19
1>
1C
b111 G
#564280000000
0!
0*
09
0>
0C
#564290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#564300000000
0!
0*
09
0>
0C
#564310000000
1!
1*
b1 6
19
1>
1C
b1 G
#564320000000
0!
0*
09
0>
0C
#564330000000
1!
1*
b10 6
19
1>
1C
b10 G
#564340000000
0!
0*
09
0>
0C
#564350000000
1!
1*
b11 6
19
1>
1C
b11 G
#564360000000
0!
0*
09
0>
0C
#564370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#564380000000
0!
0*
09
0>
0C
#564390000000
1!
1*
b101 6
19
1>
1C
b101 G
#564400000000
0!
0*
09
0>
0C
#564410000000
1!
1*
b110 6
19
1>
1C
b110 G
#564420000000
0!
0*
09
0>
0C
#564430000000
1!
1*
b111 6
19
1>
1C
b111 G
#564440000000
0!
1"
0*
1+
09
1:
0>
0C
#564450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#564460000000
0!
0*
09
0>
0C
#564470000000
1!
1*
b1 6
19
1>
1C
b1 G
#564480000000
0!
0*
09
0>
0C
#564490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#564500000000
0!
0*
09
0>
0C
#564510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#564520000000
0!
0*
09
0>
0C
#564530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#564540000000
0!
0*
09
0>
0C
#564550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#564560000000
0!
0#
0*
0,
09
0>
0?
0C
#564570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#564580000000
0!
0*
09
0>
0C
#564590000000
1!
1*
19
1>
1C
#564600000000
0!
0*
09
0>
0C
#564610000000
1!
1*
19
1>
1C
#564620000000
0!
0*
09
0>
0C
#564630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#564640000000
0!
0*
09
0>
0C
#564650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#564660000000
0!
0*
09
0>
0C
#564670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#564680000000
0!
0*
09
0>
0C
#564690000000
1!
1*
b10 6
19
1>
1C
b10 G
#564700000000
0!
0*
09
0>
0C
#564710000000
1!
1*
b11 6
19
1>
1C
b11 G
#564720000000
0!
0*
09
0>
0C
#564730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#564740000000
0!
0*
09
0>
0C
#564750000000
1!
1*
b101 6
19
1>
1C
b101 G
#564760000000
0!
0*
09
0>
0C
#564770000000
1!
1*
b110 6
19
1>
1C
b110 G
#564780000000
0!
0*
09
0>
0C
#564790000000
1!
1*
b111 6
19
1>
1C
b111 G
#564800000000
0!
0*
09
0>
0C
#564810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#564820000000
0!
0*
09
0>
0C
#564830000000
1!
1*
b1 6
19
1>
1C
b1 G
#564840000000
0!
0*
09
0>
0C
#564850000000
1!
1*
b10 6
19
1>
1C
b10 G
#564860000000
0!
0*
09
0>
0C
#564870000000
1!
1*
b11 6
19
1>
1C
b11 G
#564880000000
0!
0*
09
0>
0C
#564890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#564900000000
0!
0*
09
0>
0C
#564910000000
1!
1*
b101 6
19
1>
1C
b101 G
#564920000000
0!
0*
09
0>
0C
#564930000000
1!
1*
b110 6
19
1>
1C
b110 G
#564940000000
0!
0*
09
0>
0C
#564950000000
1!
1*
b111 6
19
1>
1C
b111 G
#564960000000
0!
0*
09
0>
0C
#564970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#564980000000
0!
0*
09
0>
0C
#564990000000
1!
1*
b1 6
19
1>
1C
b1 G
#565000000000
0!
0*
09
0>
0C
#565010000000
1!
1*
b10 6
19
1>
1C
b10 G
#565020000000
0!
0*
09
0>
0C
#565030000000
1!
1*
b11 6
19
1>
1C
b11 G
#565040000000
0!
0*
09
0>
0C
#565050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#565060000000
0!
0*
09
0>
0C
#565070000000
1!
1*
b101 6
19
1>
1C
b101 G
#565080000000
0!
0*
09
0>
0C
#565090000000
1!
1*
b110 6
19
1>
1C
b110 G
#565100000000
0!
0*
09
0>
0C
#565110000000
1!
1*
b111 6
19
1>
1C
b111 G
#565120000000
0!
1"
0*
1+
09
1:
0>
0C
#565130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#565140000000
0!
0*
09
0>
0C
#565150000000
1!
1*
b1 6
19
1>
1C
b1 G
#565160000000
0!
0*
09
0>
0C
#565170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#565180000000
0!
0*
09
0>
0C
#565190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#565200000000
0!
0*
09
0>
0C
#565210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#565220000000
0!
0*
09
0>
0C
#565230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#565240000000
0!
0#
0*
0,
09
0>
0?
0C
#565250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#565260000000
0!
0*
09
0>
0C
#565270000000
1!
1*
19
1>
1C
#565280000000
0!
0*
09
0>
0C
#565290000000
1!
1*
19
1>
1C
#565300000000
0!
0*
09
0>
0C
#565310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#565320000000
0!
0*
09
0>
0C
#565330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#565340000000
0!
0*
09
0>
0C
#565350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#565360000000
0!
0*
09
0>
0C
#565370000000
1!
1*
b10 6
19
1>
1C
b10 G
#565380000000
0!
0*
09
0>
0C
#565390000000
1!
1*
b11 6
19
1>
1C
b11 G
#565400000000
0!
0*
09
0>
0C
#565410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#565420000000
0!
0*
09
0>
0C
#565430000000
1!
1*
b101 6
19
1>
1C
b101 G
#565440000000
0!
0*
09
0>
0C
#565450000000
1!
1*
b110 6
19
1>
1C
b110 G
#565460000000
0!
0*
09
0>
0C
#565470000000
1!
1*
b111 6
19
1>
1C
b111 G
#565480000000
0!
0*
09
0>
0C
#565490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#565500000000
0!
0*
09
0>
0C
#565510000000
1!
1*
b1 6
19
1>
1C
b1 G
#565520000000
0!
0*
09
0>
0C
#565530000000
1!
1*
b10 6
19
1>
1C
b10 G
#565540000000
0!
0*
09
0>
0C
#565550000000
1!
1*
b11 6
19
1>
1C
b11 G
#565560000000
0!
0*
09
0>
0C
#565570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#565580000000
0!
0*
09
0>
0C
#565590000000
1!
1*
b101 6
19
1>
1C
b101 G
#565600000000
0!
0*
09
0>
0C
#565610000000
1!
1*
b110 6
19
1>
1C
b110 G
#565620000000
0!
0*
09
0>
0C
#565630000000
1!
1*
b111 6
19
1>
1C
b111 G
#565640000000
0!
0*
09
0>
0C
#565650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#565660000000
0!
0*
09
0>
0C
#565670000000
1!
1*
b1 6
19
1>
1C
b1 G
#565680000000
0!
0*
09
0>
0C
#565690000000
1!
1*
b10 6
19
1>
1C
b10 G
#565700000000
0!
0*
09
0>
0C
#565710000000
1!
1*
b11 6
19
1>
1C
b11 G
#565720000000
0!
0*
09
0>
0C
#565730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#565740000000
0!
0*
09
0>
0C
#565750000000
1!
1*
b101 6
19
1>
1C
b101 G
#565760000000
0!
0*
09
0>
0C
#565770000000
1!
1*
b110 6
19
1>
1C
b110 G
#565780000000
0!
0*
09
0>
0C
#565790000000
1!
1*
b111 6
19
1>
1C
b111 G
#565800000000
0!
1"
0*
1+
09
1:
0>
0C
#565810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#565820000000
0!
0*
09
0>
0C
#565830000000
1!
1*
b1 6
19
1>
1C
b1 G
#565840000000
0!
0*
09
0>
0C
#565850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#565860000000
0!
0*
09
0>
0C
#565870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#565880000000
0!
0*
09
0>
0C
#565890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#565900000000
0!
0*
09
0>
0C
#565910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#565920000000
0!
0#
0*
0,
09
0>
0?
0C
#565930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#565940000000
0!
0*
09
0>
0C
#565950000000
1!
1*
19
1>
1C
#565960000000
0!
0*
09
0>
0C
#565970000000
1!
1*
19
1>
1C
#565980000000
0!
0*
09
0>
0C
#565990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#566000000000
0!
0*
09
0>
0C
#566010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#566020000000
0!
0*
09
0>
0C
#566030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#566040000000
0!
0*
09
0>
0C
#566050000000
1!
1*
b10 6
19
1>
1C
b10 G
#566060000000
0!
0*
09
0>
0C
#566070000000
1!
1*
b11 6
19
1>
1C
b11 G
#566080000000
0!
0*
09
0>
0C
#566090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#566100000000
0!
0*
09
0>
0C
#566110000000
1!
1*
b101 6
19
1>
1C
b101 G
#566120000000
0!
0*
09
0>
0C
#566130000000
1!
1*
b110 6
19
1>
1C
b110 G
#566140000000
0!
0*
09
0>
0C
#566150000000
1!
1*
b111 6
19
1>
1C
b111 G
#566160000000
0!
0*
09
0>
0C
#566170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#566180000000
0!
0*
09
0>
0C
#566190000000
1!
1*
b1 6
19
1>
1C
b1 G
#566200000000
0!
0*
09
0>
0C
#566210000000
1!
1*
b10 6
19
1>
1C
b10 G
#566220000000
0!
0*
09
0>
0C
#566230000000
1!
1*
b11 6
19
1>
1C
b11 G
#566240000000
0!
0*
09
0>
0C
#566250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#566260000000
0!
0*
09
0>
0C
#566270000000
1!
1*
b101 6
19
1>
1C
b101 G
#566280000000
0!
0*
09
0>
0C
#566290000000
1!
1*
b110 6
19
1>
1C
b110 G
#566300000000
0!
0*
09
0>
0C
#566310000000
1!
1*
b111 6
19
1>
1C
b111 G
#566320000000
0!
0*
09
0>
0C
#566330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#566340000000
0!
0*
09
0>
0C
#566350000000
1!
1*
b1 6
19
1>
1C
b1 G
#566360000000
0!
0*
09
0>
0C
#566370000000
1!
1*
b10 6
19
1>
1C
b10 G
#566380000000
0!
0*
09
0>
0C
#566390000000
1!
1*
b11 6
19
1>
1C
b11 G
#566400000000
0!
0*
09
0>
0C
#566410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#566420000000
0!
0*
09
0>
0C
#566430000000
1!
1*
b101 6
19
1>
1C
b101 G
#566440000000
0!
0*
09
0>
0C
#566450000000
1!
1*
b110 6
19
1>
1C
b110 G
#566460000000
0!
0*
09
0>
0C
#566470000000
1!
1*
b111 6
19
1>
1C
b111 G
#566480000000
0!
1"
0*
1+
09
1:
0>
0C
#566490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#566500000000
0!
0*
09
0>
0C
#566510000000
1!
1*
b1 6
19
1>
1C
b1 G
#566520000000
0!
0*
09
0>
0C
#566530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#566540000000
0!
0*
09
0>
0C
#566550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#566560000000
0!
0*
09
0>
0C
#566570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#566580000000
0!
0*
09
0>
0C
#566590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#566600000000
0!
0#
0*
0,
09
0>
0?
0C
#566610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#566620000000
0!
0*
09
0>
0C
#566630000000
1!
1*
19
1>
1C
#566640000000
0!
0*
09
0>
0C
#566650000000
1!
1*
19
1>
1C
#566660000000
0!
0*
09
0>
0C
#566670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#566680000000
0!
0*
09
0>
0C
#566690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#566700000000
0!
0*
09
0>
0C
#566710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#566720000000
0!
0*
09
0>
0C
#566730000000
1!
1*
b10 6
19
1>
1C
b10 G
#566740000000
0!
0*
09
0>
0C
#566750000000
1!
1*
b11 6
19
1>
1C
b11 G
#566760000000
0!
0*
09
0>
0C
#566770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#566780000000
0!
0*
09
0>
0C
#566790000000
1!
1*
b101 6
19
1>
1C
b101 G
#566800000000
0!
0*
09
0>
0C
#566810000000
1!
1*
b110 6
19
1>
1C
b110 G
#566820000000
0!
0*
09
0>
0C
#566830000000
1!
1*
b111 6
19
1>
1C
b111 G
#566840000000
0!
0*
09
0>
0C
#566850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#566860000000
0!
0*
09
0>
0C
#566870000000
1!
1*
b1 6
19
1>
1C
b1 G
#566880000000
0!
0*
09
0>
0C
#566890000000
1!
1*
b10 6
19
1>
1C
b10 G
#566900000000
0!
0*
09
0>
0C
#566910000000
1!
1*
b11 6
19
1>
1C
b11 G
#566920000000
0!
0*
09
0>
0C
#566930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#566940000000
0!
0*
09
0>
0C
#566950000000
1!
1*
b101 6
19
1>
1C
b101 G
#566960000000
0!
0*
09
0>
0C
#566970000000
1!
1*
b110 6
19
1>
1C
b110 G
#566980000000
0!
0*
09
0>
0C
#566990000000
1!
1*
b111 6
19
1>
1C
b111 G
#567000000000
0!
0*
09
0>
0C
#567010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#567020000000
0!
0*
09
0>
0C
#567030000000
1!
1*
b1 6
19
1>
1C
b1 G
#567040000000
0!
0*
09
0>
0C
#567050000000
1!
1*
b10 6
19
1>
1C
b10 G
#567060000000
0!
0*
09
0>
0C
#567070000000
1!
1*
b11 6
19
1>
1C
b11 G
#567080000000
0!
0*
09
0>
0C
#567090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#567100000000
0!
0*
09
0>
0C
#567110000000
1!
1*
b101 6
19
1>
1C
b101 G
#567120000000
0!
0*
09
0>
0C
#567130000000
1!
1*
b110 6
19
1>
1C
b110 G
#567140000000
0!
0*
09
0>
0C
#567150000000
1!
1*
b111 6
19
1>
1C
b111 G
#567160000000
0!
1"
0*
1+
09
1:
0>
0C
#567170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#567180000000
0!
0*
09
0>
0C
#567190000000
1!
1*
b1 6
19
1>
1C
b1 G
#567200000000
0!
0*
09
0>
0C
#567210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#567220000000
0!
0*
09
0>
0C
#567230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#567240000000
0!
0*
09
0>
0C
#567250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#567260000000
0!
0*
09
0>
0C
#567270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#567280000000
0!
0#
0*
0,
09
0>
0?
0C
#567290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#567300000000
0!
0*
09
0>
0C
#567310000000
1!
1*
19
1>
1C
#567320000000
0!
0*
09
0>
0C
#567330000000
1!
1*
19
1>
1C
#567340000000
0!
0*
09
0>
0C
#567350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#567360000000
0!
0*
09
0>
0C
#567370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#567380000000
0!
0*
09
0>
0C
#567390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#567400000000
0!
0*
09
0>
0C
#567410000000
1!
1*
b10 6
19
1>
1C
b10 G
#567420000000
0!
0*
09
0>
0C
#567430000000
1!
1*
b11 6
19
1>
1C
b11 G
#567440000000
0!
0*
09
0>
0C
#567450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#567460000000
0!
0*
09
0>
0C
#567470000000
1!
1*
b101 6
19
1>
1C
b101 G
#567480000000
0!
0*
09
0>
0C
#567490000000
1!
1*
b110 6
19
1>
1C
b110 G
#567500000000
0!
0*
09
0>
0C
#567510000000
1!
1*
b111 6
19
1>
1C
b111 G
#567520000000
0!
0*
09
0>
0C
#567530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#567540000000
0!
0*
09
0>
0C
#567550000000
1!
1*
b1 6
19
1>
1C
b1 G
#567560000000
0!
0*
09
0>
0C
#567570000000
1!
1*
b10 6
19
1>
1C
b10 G
#567580000000
0!
0*
09
0>
0C
#567590000000
1!
1*
b11 6
19
1>
1C
b11 G
#567600000000
0!
0*
09
0>
0C
#567610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#567620000000
0!
0*
09
0>
0C
#567630000000
1!
1*
b101 6
19
1>
1C
b101 G
#567640000000
0!
0*
09
0>
0C
#567650000000
1!
1*
b110 6
19
1>
1C
b110 G
#567660000000
0!
0*
09
0>
0C
#567670000000
1!
1*
b111 6
19
1>
1C
b111 G
#567680000000
0!
0*
09
0>
0C
#567690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#567700000000
0!
0*
09
0>
0C
#567710000000
1!
1*
b1 6
19
1>
1C
b1 G
#567720000000
0!
0*
09
0>
0C
#567730000000
1!
1*
b10 6
19
1>
1C
b10 G
#567740000000
0!
0*
09
0>
0C
#567750000000
1!
1*
b11 6
19
1>
1C
b11 G
#567760000000
0!
0*
09
0>
0C
#567770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#567780000000
0!
0*
09
0>
0C
#567790000000
1!
1*
b101 6
19
1>
1C
b101 G
#567800000000
0!
0*
09
0>
0C
#567810000000
1!
1*
b110 6
19
1>
1C
b110 G
#567820000000
0!
0*
09
0>
0C
#567830000000
1!
1*
b111 6
19
1>
1C
b111 G
#567840000000
0!
1"
0*
1+
09
1:
0>
0C
#567850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#567860000000
0!
0*
09
0>
0C
#567870000000
1!
1*
b1 6
19
1>
1C
b1 G
#567880000000
0!
0*
09
0>
0C
#567890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#567900000000
0!
0*
09
0>
0C
#567910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#567920000000
0!
0*
09
0>
0C
#567930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#567940000000
0!
0*
09
0>
0C
#567950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#567960000000
0!
0#
0*
0,
09
0>
0?
0C
#567970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#567980000000
0!
0*
09
0>
0C
#567990000000
1!
1*
19
1>
1C
#568000000000
0!
0*
09
0>
0C
#568010000000
1!
1*
19
1>
1C
#568020000000
0!
0*
09
0>
0C
#568030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#568040000000
0!
0*
09
0>
0C
#568050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#568060000000
0!
0*
09
0>
0C
#568070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#568080000000
0!
0*
09
0>
0C
#568090000000
1!
1*
b10 6
19
1>
1C
b10 G
#568100000000
0!
0*
09
0>
0C
#568110000000
1!
1*
b11 6
19
1>
1C
b11 G
#568120000000
0!
0*
09
0>
0C
#568130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#568140000000
0!
0*
09
0>
0C
#568150000000
1!
1*
b101 6
19
1>
1C
b101 G
#568160000000
0!
0*
09
0>
0C
#568170000000
1!
1*
b110 6
19
1>
1C
b110 G
#568180000000
0!
0*
09
0>
0C
#568190000000
1!
1*
b111 6
19
1>
1C
b111 G
#568200000000
0!
0*
09
0>
0C
#568210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#568220000000
0!
0*
09
0>
0C
#568230000000
1!
1*
b1 6
19
1>
1C
b1 G
#568240000000
0!
0*
09
0>
0C
#568250000000
1!
1*
b10 6
19
1>
1C
b10 G
#568260000000
0!
0*
09
0>
0C
#568270000000
1!
1*
b11 6
19
1>
1C
b11 G
#568280000000
0!
0*
09
0>
0C
#568290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#568300000000
0!
0*
09
0>
0C
#568310000000
1!
1*
b101 6
19
1>
1C
b101 G
#568320000000
0!
0*
09
0>
0C
#568330000000
1!
1*
b110 6
19
1>
1C
b110 G
#568340000000
0!
0*
09
0>
0C
#568350000000
1!
1*
b111 6
19
1>
1C
b111 G
#568360000000
0!
0*
09
0>
0C
#568370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#568380000000
0!
0*
09
0>
0C
#568390000000
1!
1*
b1 6
19
1>
1C
b1 G
#568400000000
0!
0*
09
0>
0C
#568410000000
1!
1*
b10 6
19
1>
1C
b10 G
#568420000000
0!
0*
09
0>
0C
#568430000000
1!
1*
b11 6
19
1>
1C
b11 G
#568440000000
0!
0*
09
0>
0C
#568450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#568460000000
0!
0*
09
0>
0C
#568470000000
1!
1*
b101 6
19
1>
1C
b101 G
#568480000000
0!
0*
09
0>
0C
#568490000000
1!
1*
b110 6
19
1>
1C
b110 G
#568500000000
0!
0*
09
0>
0C
#568510000000
1!
1*
b111 6
19
1>
1C
b111 G
#568520000000
0!
1"
0*
1+
09
1:
0>
0C
#568530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#568540000000
0!
0*
09
0>
0C
#568550000000
1!
1*
b1 6
19
1>
1C
b1 G
#568560000000
0!
0*
09
0>
0C
#568570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#568580000000
0!
0*
09
0>
0C
#568590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#568600000000
0!
0*
09
0>
0C
#568610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#568620000000
0!
0*
09
0>
0C
#568630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#568640000000
0!
0#
0*
0,
09
0>
0?
0C
#568650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#568660000000
0!
0*
09
0>
0C
#568670000000
1!
1*
19
1>
1C
#568680000000
0!
0*
09
0>
0C
#568690000000
1!
1*
19
1>
1C
#568700000000
0!
0*
09
0>
0C
#568710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#568720000000
0!
0*
09
0>
0C
#568730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#568740000000
0!
0*
09
0>
0C
#568750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#568760000000
0!
0*
09
0>
0C
#568770000000
1!
1*
b10 6
19
1>
1C
b10 G
#568780000000
0!
0*
09
0>
0C
#568790000000
1!
1*
b11 6
19
1>
1C
b11 G
#568800000000
0!
0*
09
0>
0C
#568810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#568820000000
0!
0*
09
0>
0C
#568830000000
1!
1*
b101 6
19
1>
1C
b101 G
#568840000000
0!
0*
09
0>
0C
#568850000000
1!
1*
b110 6
19
1>
1C
b110 G
#568860000000
0!
0*
09
0>
0C
#568870000000
1!
1*
b111 6
19
1>
1C
b111 G
#568880000000
0!
0*
09
0>
0C
#568890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#568900000000
0!
0*
09
0>
0C
#568910000000
1!
1*
b1 6
19
1>
1C
b1 G
#568920000000
0!
0*
09
0>
0C
#568930000000
1!
1*
b10 6
19
1>
1C
b10 G
#568940000000
0!
0*
09
0>
0C
#568950000000
1!
1*
b11 6
19
1>
1C
b11 G
#568960000000
0!
0*
09
0>
0C
#568970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#568980000000
0!
0*
09
0>
0C
#568990000000
1!
1*
b101 6
19
1>
1C
b101 G
#569000000000
0!
0*
09
0>
0C
#569010000000
1!
1*
b110 6
19
1>
1C
b110 G
#569020000000
0!
0*
09
0>
0C
#569030000000
1!
1*
b111 6
19
1>
1C
b111 G
#569040000000
0!
0*
09
0>
0C
#569050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#569060000000
0!
0*
09
0>
0C
#569070000000
1!
1*
b1 6
19
1>
1C
b1 G
#569080000000
0!
0*
09
0>
0C
#569090000000
1!
1*
b10 6
19
1>
1C
b10 G
#569100000000
0!
0*
09
0>
0C
#569110000000
1!
1*
b11 6
19
1>
1C
b11 G
#569120000000
0!
0*
09
0>
0C
#569130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#569140000000
0!
0*
09
0>
0C
#569150000000
1!
1*
b101 6
19
1>
1C
b101 G
#569160000000
0!
0*
09
0>
0C
#569170000000
1!
1*
b110 6
19
1>
1C
b110 G
#569180000000
0!
0*
09
0>
0C
#569190000000
1!
1*
b111 6
19
1>
1C
b111 G
#569200000000
0!
1"
0*
1+
09
1:
0>
0C
#569210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#569220000000
0!
0*
09
0>
0C
#569230000000
1!
1*
b1 6
19
1>
1C
b1 G
#569240000000
0!
0*
09
0>
0C
#569250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#569260000000
0!
0*
09
0>
0C
#569270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#569280000000
0!
0*
09
0>
0C
#569290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#569300000000
0!
0*
09
0>
0C
#569310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#569320000000
0!
0#
0*
0,
09
0>
0?
0C
#569330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#569340000000
0!
0*
09
0>
0C
#569350000000
1!
1*
19
1>
1C
#569360000000
0!
0*
09
0>
0C
#569370000000
1!
1*
19
1>
1C
#569380000000
0!
0*
09
0>
0C
#569390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#569400000000
0!
0*
09
0>
0C
#569410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#569420000000
0!
0*
09
0>
0C
#569430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#569440000000
0!
0*
09
0>
0C
#569450000000
1!
1*
b10 6
19
1>
1C
b10 G
#569460000000
0!
0*
09
0>
0C
#569470000000
1!
1*
b11 6
19
1>
1C
b11 G
#569480000000
0!
0*
09
0>
0C
#569490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#569500000000
0!
0*
09
0>
0C
#569510000000
1!
1*
b101 6
19
1>
1C
b101 G
#569520000000
0!
0*
09
0>
0C
#569530000000
1!
1*
b110 6
19
1>
1C
b110 G
#569540000000
0!
0*
09
0>
0C
#569550000000
1!
1*
b111 6
19
1>
1C
b111 G
#569560000000
0!
0*
09
0>
0C
#569570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#569580000000
0!
0*
09
0>
0C
#569590000000
1!
1*
b1 6
19
1>
1C
b1 G
#569600000000
0!
0*
09
0>
0C
#569610000000
1!
1*
b10 6
19
1>
1C
b10 G
#569620000000
0!
0*
09
0>
0C
#569630000000
1!
1*
b11 6
19
1>
1C
b11 G
#569640000000
0!
0*
09
0>
0C
#569650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#569660000000
0!
0*
09
0>
0C
#569670000000
1!
1*
b101 6
19
1>
1C
b101 G
#569680000000
0!
0*
09
0>
0C
#569690000000
1!
1*
b110 6
19
1>
1C
b110 G
#569700000000
0!
0*
09
0>
0C
#569710000000
1!
1*
b111 6
19
1>
1C
b111 G
#569720000000
0!
0*
09
0>
0C
#569730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#569740000000
0!
0*
09
0>
0C
#569750000000
1!
1*
b1 6
19
1>
1C
b1 G
#569760000000
0!
0*
09
0>
0C
#569770000000
1!
1*
b10 6
19
1>
1C
b10 G
#569780000000
0!
0*
09
0>
0C
#569790000000
1!
1*
b11 6
19
1>
1C
b11 G
#569800000000
0!
0*
09
0>
0C
#569810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#569820000000
0!
0*
09
0>
0C
#569830000000
1!
1*
b101 6
19
1>
1C
b101 G
#569840000000
0!
0*
09
0>
0C
#569850000000
1!
1*
b110 6
19
1>
1C
b110 G
#569860000000
0!
0*
09
0>
0C
#569870000000
1!
1*
b111 6
19
1>
1C
b111 G
#569880000000
0!
1"
0*
1+
09
1:
0>
0C
#569890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#569900000000
0!
0*
09
0>
0C
#569910000000
1!
1*
b1 6
19
1>
1C
b1 G
#569920000000
0!
0*
09
0>
0C
#569930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#569940000000
0!
0*
09
0>
0C
#569950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#569960000000
0!
0*
09
0>
0C
#569970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#569980000000
0!
0*
09
0>
0C
#569990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#570000000000
0!
0#
0*
0,
09
0>
0?
0C
#570010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#570020000000
0!
0*
09
0>
0C
#570030000000
1!
1*
19
1>
1C
#570040000000
0!
0*
09
0>
0C
#570050000000
1!
1*
19
1>
1C
#570060000000
0!
0*
09
0>
0C
#570070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#570080000000
0!
0*
09
0>
0C
#570090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#570100000000
0!
0*
09
0>
0C
#570110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#570120000000
0!
0*
09
0>
0C
#570130000000
1!
1*
b10 6
19
1>
1C
b10 G
#570140000000
0!
0*
09
0>
0C
#570150000000
1!
1*
b11 6
19
1>
1C
b11 G
#570160000000
0!
0*
09
0>
0C
#570170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#570180000000
0!
0*
09
0>
0C
#570190000000
1!
1*
b101 6
19
1>
1C
b101 G
#570200000000
0!
0*
09
0>
0C
#570210000000
1!
1*
b110 6
19
1>
1C
b110 G
#570220000000
0!
0*
09
0>
0C
#570230000000
1!
1*
b111 6
19
1>
1C
b111 G
#570240000000
0!
0*
09
0>
0C
#570250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#570260000000
0!
0*
09
0>
0C
#570270000000
1!
1*
b1 6
19
1>
1C
b1 G
#570280000000
0!
0*
09
0>
0C
#570290000000
1!
1*
b10 6
19
1>
1C
b10 G
#570300000000
0!
0*
09
0>
0C
#570310000000
1!
1*
b11 6
19
1>
1C
b11 G
#570320000000
0!
0*
09
0>
0C
#570330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#570340000000
0!
0*
09
0>
0C
#570350000000
1!
1*
b101 6
19
1>
1C
b101 G
#570360000000
0!
0*
09
0>
0C
#570370000000
1!
1*
b110 6
19
1>
1C
b110 G
#570380000000
0!
0*
09
0>
0C
#570390000000
1!
1*
b111 6
19
1>
1C
b111 G
#570400000000
0!
0*
09
0>
0C
#570410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#570420000000
0!
0*
09
0>
0C
#570430000000
1!
1*
b1 6
19
1>
1C
b1 G
#570440000000
0!
0*
09
0>
0C
#570450000000
1!
1*
b10 6
19
1>
1C
b10 G
#570460000000
0!
0*
09
0>
0C
#570470000000
1!
1*
b11 6
19
1>
1C
b11 G
#570480000000
0!
0*
09
0>
0C
#570490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#570500000000
0!
0*
09
0>
0C
#570510000000
1!
1*
b101 6
19
1>
1C
b101 G
#570520000000
0!
0*
09
0>
0C
#570530000000
1!
1*
b110 6
19
1>
1C
b110 G
#570540000000
0!
0*
09
0>
0C
#570550000000
1!
1*
b111 6
19
1>
1C
b111 G
#570560000000
0!
1"
0*
1+
09
1:
0>
0C
#570570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#570580000000
0!
0*
09
0>
0C
#570590000000
1!
1*
b1 6
19
1>
1C
b1 G
#570600000000
0!
0*
09
0>
0C
#570610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#570620000000
0!
0*
09
0>
0C
#570630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#570640000000
0!
0*
09
0>
0C
#570650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#570660000000
0!
0*
09
0>
0C
#570670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#570680000000
0!
0#
0*
0,
09
0>
0?
0C
#570690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#570700000000
0!
0*
09
0>
0C
#570710000000
1!
1*
19
1>
1C
#570720000000
0!
0*
09
0>
0C
#570730000000
1!
1*
19
1>
1C
#570740000000
0!
0*
09
0>
0C
#570750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#570760000000
0!
0*
09
0>
0C
#570770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#570780000000
0!
0*
09
0>
0C
#570790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#570800000000
0!
0*
09
0>
0C
#570810000000
1!
1*
b10 6
19
1>
1C
b10 G
#570820000000
0!
0*
09
0>
0C
#570830000000
1!
1*
b11 6
19
1>
1C
b11 G
#570840000000
0!
0*
09
0>
0C
#570850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#570860000000
0!
0*
09
0>
0C
#570870000000
1!
1*
b101 6
19
1>
1C
b101 G
#570880000000
0!
0*
09
0>
0C
#570890000000
1!
1*
b110 6
19
1>
1C
b110 G
#570900000000
0!
0*
09
0>
0C
#570910000000
1!
1*
b111 6
19
1>
1C
b111 G
#570920000000
0!
0*
09
0>
0C
#570930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#570940000000
0!
0*
09
0>
0C
#570950000000
1!
1*
b1 6
19
1>
1C
b1 G
#570960000000
0!
0*
09
0>
0C
#570970000000
1!
1*
b10 6
19
1>
1C
b10 G
#570980000000
0!
0*
09
0>
0C
#570990000000
1!
1*
b11 6
19
1>
1C
b11 G
#571000000000
0!
0*
09
0>
0C
#571010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#571020000000
0!
0*
09
0>
0C
#571030000000
1!
1*
b101 6
19
1>
1C
b101 G
#571040000000
0!
0*
09
0>
0C
#571050000000
1!
1*
b110 6
19
1>
1C
b110 G
#571060000000
0!
0*
09
0>
0C
#571070000000
1!
1*
b111 6
19
1>
1C
b111 G
#571080000000
0!
0*
09
0>
0C
#571090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#571100000000
0!
0*
09
0>
0C
#571110000000
1!
1*
b1 6
19
1>
1C
b1 G
#571120000000
0!
0*
09
0>
0C
#571130000000
1!
1*
b10 6
19
1>
1C
b10 G
#571140000000
0!
0*
09
0>
0C
#571150000000
1!
1*
b11 6
19
1>
1C
b11 G
#571160000000
0!
0*
09
0>
0C
#571170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#571180000000
0!
0*
09
0>
0C
#571190000000
1!
1*
b101 6
19
1>
1C
b101 G
#571200000000
0!
0*
09
0>
0C
#571210000000
1!
1*
b110 6
19
1>
1C
b110 G
#571220000000
0!
0*
09
0>
0C
#571230000000
1!
1*
b111 6
19
1>
1C
b111 G
#571240000000
0!
1"
0*
1+
09
1:
0>
0C
#571250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#571260000000
0!
0*
09
0>
0C
#571270000000
1!
1*
b1 6
19
1>
1C
b1 G
#571280000000
0!
0*
09
0>
0C
#571290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#571300000000
0!
0*
09
0>
0C
#571310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#571320000000
0!
0*
09
0>
0C
#571330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#571340000000
0!
0*
09
0>
0C
#571350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#571360000000
0!
0#
0*
0,
09
0>
0?
0C
#571370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#571380000000
0!
0*
09
0>
0C
#571390000000
1!
1*
19
1>
1C
#571400000000
0!
0*
09
0>
0C
#571410000000
1!
1*
19
1>
1C
#571420000000
0!
0*
09
0>
0C
#571430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#571440000000
0!
0*
09
0>
0C
#571450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#571460000000
0!
0*
09
0>
0C
#571470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#571480000000
0!
0*
09
0>
0C
#571490000000
1!
1*
b10 6
19
1>
1C
b10 G
#571500000000
0!
0*
09
0>
0C
#571510000000
1!
1*
b11 6
19
1>
1C
b11 G
#571520000000
0!
0*
09
0>
0C
#571530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#571540000000
0!
0*
09
0>
0C
#571550000000
1!
1*
b101 6
19
1>
1C
b101 G
#571560000000
0!
0*
09
0>
0C
#571570000000
1!
1*
b110 6
19
1>
1C
b110 G
#571580000000
0!
0*
09
0>
0C
#571590000000
1!
1*
b111 6
19
1>
1C
b111 G
#571600000000
0!
0*
09
0>
0C
#571610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#571620000000
0!
0*
09
0>
0C
#571630000000
1!
1*
b1 6
19
1>
1C
b1 G
#571640000000
0!
0*
09
0>
0C
#571650000000
1!
1*
b10 6
19
1>
1C
b10 G
#571660000000
0!
0*
09
0>
0C
#571670000000
1!
1*
b11 6
19
1>
1C
b11 G
#571680000000
0!
0*
09
0>
0C
#571690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#571700000000
0!
0*
09
0>
0C
#571710000000
1!
1*
b101 6
19
1>
1C
b101 G
#571720000000
0!
0*
09
0>
0C
#571730000000
1!
1*
b110 6
19
1>
1C
b110 G
#571740000000
0!
0*
09
0>
0C
#571750000000
1!
1*
b111 6
19
1>
1C
b111 G
#571760000000
0!
0*
09
0>
0C
#571770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#571780000000
0!
0*
09
0>
0C
#571790000000
1!
1*
b1 6
19
1>
1C
b1 G
#571800000000
0!
0*
09
0>
0C
#571810000000
1!
1*
b10 6
19
1>
1C
b10 G
#571820000000
0!
0*
09
0>
0C
#571830000000
1!
1*
b11 6
19
1>
1C
b11 G
#571840000000
0!
0*
09
0>
0C
#571850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#571860000000
0!
0*
09
0>
0C
#571870000000
1!
1*
b101 6
19
1>
1C
b101 G
#571880000000
0!
0*
09
0>
0C
#571890000000
1!
1*
b110 6
19
1>
1C
b110 G
#571900000000
0!
0*
09
0>
0C
#571910000000
1!
1*
b111 6
19
1>
1C
b111 G
#571920000000
0!
1"
0*
1+
09
1:
0>
0C
#571930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#571940000000
0!
0*
09
0>
0C
#571950000000
1!
1*
b1 6
19
1>
1C
b1 G
#571960000000
0!
0*
09
0>
0C
#571970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#571980000000
0!
0*
09
0>
0C
#571990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#572000000000
0!
0*
09
0>
0C
#572010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#572020000000
0!
0*
09
0>
0C
#572030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#572040000000
0!
0#
0*
0,
09
0>
0?
0C
#572050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#572060000000
0!
0*
09
0>
0C
#572070000000
1!
1*
19
1>
1C
#572080000000
0!
0*
09
0>
0C
#572090000000
1!
1*
19
1>
1C
#572100000000
0!
0*
09
0>
0C
#572110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#572120000000
0!
0*
09
0>
0C
#572130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#572140000000
0!
0*
09
0>
0C
#572150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#572160000000
0!
0*
09
0>
0C
#572170000000
1!
1*
b10 6
19
1>
1C
b10 G
#572180000000
0!
0*
09
0>
0C
#572190000000
1!
1*
b11 6
19
1>
1C
b11 G
#572200000000
0!
0*
09
0>
0C
#572210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#572220000000
0!
0*
09
0>
0C
#572230000000
1!
1*
b101 6
19
1>
1C
b101 G
#572240000000
0!
0*
09
0>
0C
#572250000000
1!
1*
b110 6
19
1>
1C
b110 G
#572260000000
0!
0*
09
0>
0C
#572270000000
1!
1*
b111 6
19
1>
1C
b111 G
#572280000000
0!
0*
09
0>
0C
#572290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#572300000000
0!
0*
09
0>
0C
#572310000000
1!
1*
b1 6
19
1>
1C
b1 G
#572320000000
0!
0*
09
0>
0C
#572330000000
1!
1*
b10 6
19
1>
1C
b10 G
#572340000000
0!
0*
09
0>
0C
#572350000000
1!
1*
b11 6
19
1>
1C
b11 G
#572360000000
0!
0*
09
0>
0C
#572370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#572380000000
0!
0*
09
0>
0C
#572390000000
1!
1*
b101 6
19
1>
1C
b101 G
#572400000000
0!
0*
09
0>
0C
#572410000000
1!
1*
b110 6
19
1>
1C
b110 G
#572420000000
0!
0*
09
0>
0C
#572430000000
1!
1*
b111 6
19
1>
1C
b111 G
#572440000000
0!
0*
09
0>
0C
#572450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#572460000000
0!
0*
09
0>
0C
#572470000000
1!
1*
b1 6
19
1>
1C
b1 G
#572480000000
0!
0*
09
0>
0C
#572490000000
1!
1*
b10 6
19
1>
1C
b10 G
#572500000000
0!
0*
09
0>
0C
#572510000000
1!
1*
b11 6
19
1>
1C
b11 G
#572520000000
0!
0*
09
0>
0C
#572530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#572540000000
0!
0*
09
0>
0C
#572550000000
1!
1*
b101 6
19
1>
1C
b101 G
#572560000000
0!
0*
09
0>
0C
#572570000000
1!
1*
b110 6
19
1>
1C
b110 G
#572580000000
0!
0*
09
0>
0C
#572590000000
1!
1*
b111 6
19
1>
1C
b111 G
#572600000000
0!
1"
0*
1+
09
1:
0>
0C
#572610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#572620000000
0!
0*
09
0>
0C
#572630000000
1!
1*
b1 6
19
1>
1C
b1 G
#572640000000
0!
0*
09
0>
0C
#572650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#572660000000
0!
0*
09
0>
0C
#572670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#572680000000
0!
0*
09
0>
0C
#572690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#572700000000
0!
0*
09
0>
0C
#572710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#572720000000
0!
0#
0*
0,
09
0>
0?
0C
#572730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#572740000000
0!
0*
09
0>
0C
#572750000000
1!
1*
19
1>
1C
#572760000000
0!
0*
09
0>
0C
#572770000000
1!
1*
19
1>
1C
#572780000000
0!
0*
09
0>
0C
#572790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#572800000000
0!
0*
09
0>
0C
#572810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#572820000000
0!
0*
09
0>
0C
#572830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#572840000000
0!
0*
09
0>
0C
#572850000000
1!
1*
b10 6
19
1>
1C
b10 G
#572860000000
0!
0*
09
0>
0C
#572870000000
1!
1*
b11 6
19
1>
1C
b11 G
#572880000000
0!
0*
09
0>
0C
#572890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#572900000000
0!
0*
09
0>
0C
#572910000000
1!
1*
b101 6
19
1>
1C
b101 G
#572920000000
0!
0*
09
0>
0C
#572930000000
1!
1*
b110 6
19
1>
1C
b110 G
#572940000000
0!
0*
09
0>
0C
#572950000000
1!
1*
b111 6
19
1>
1C
b111 G
#572960000000
0!
0*
09
0>
0C
#572970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#572980000000
0!
0*
09
0>
0C
#572990000000
1!
1*
b1 6
19
1>
1C
b1 G
#573000000000
0!
0*
09
0>
0C
#573010000000
1!
1*
b10 6
19
1>
1C
b10 G
#573020000000
0!
0*
09
0>
0C
#573030000000
1!
1*
b11 6
19
1>
1C
b11 G
#573040000000
0!
0*
09
0>
0C
#573050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#573060000000
0!
0*
09
0>
0C
#573070000000
1!
1*
b101 6
19
1>
1C
b101 G
#573080000000
0!
0*
09
0>
0C
#573090000000
1!
1*
b110 6
19
1>
1C
b110 G
#573100000000
0!
0*
09
0>
0C
#573110000000
1!
1*
b111 6
19
1>
1C
b111 G
#573120000000
0!
0*
09
0>
0C
#573130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#573140000000
0!
0*
09
0>
0C
#573150000000
1!
1*
b1 6
19
1>
1C
b1 G
#573160000000
0!
0*
09
0>
0C
#573170000000
1!
1*
b10 6
19
1>
1C
b10 G
#573180000000
0!
0*
09
0>
0C
#573190000000
1!
1*
b11 6
19
1>
1C
b11 G
#573200000000
0!
0*
09
0>
0C
#573210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#573220000000
0!
0*
09
0>
0C
#573230000000
1!
1*
b101 6
19
1>
1C
b101 G
#573240000000
0!
0*
09
0>
0C
#573250000000
1!
1*
b110 6
19
1>
1C
b110 G
#573260000000
0!
0*
09
0>
0C
#573270000000
1!
1*
b111 6
19
1>
1C
b111 G
#573280000000
0!
1"
0*
1+
09
1:
0>
0C
#573290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#573300000000
0!
0*
09
0>
0C
#573310000000
1!
1*
b1 6
19
1>
1C
b1 G
#573320000000
0!
0*
09
0>
0C
#573330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#573340000000
0!
0*
09
0>
0C
#573350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#573360000000
0!
0*
09
0>
0C
#573370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#573380000000
0!
0*
09
0>
0C
#573390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#573400000000
0!
0#
0*
0,
09
0>
0?
0C
#573410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#573420000000
0!
0*
09
0>
0C
#573430000000
1!
1*
19
1>
1C
#573440000000
0!
0*
09
0>
0C
#573450000000
1!
1*
19
1>
1C
#573460000000
0!
0*
09
0>
0C
#573470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#573480000000
0!
0*
09
0>
0C
#573490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#573500000000
0!
0*
09
0>
0C
#573510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#573520000000
0!
0*
09
0>
0C
#573530000000
1!
1*
b10 6
19
1>
1C
b10 G
#573540000000
0!
0*
09
0>
0C
#573550000000
1!
1*
b11 6
19
1>
1C
b11 G
#573560000000
0!
0*
09
0>
0C
#573570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#573580000000
0!
0*
09
0>
0C
#573590000000
1!
1*
b101 6
19
1>
1C
b101 G
#573600000000
0!
0*
09
0>
0C
#573610000000
1!
1*
b110 6
19
1>
1C
b110 G
#573620000000
0!
0*
09
0>
0C
#573630000000
1!
1*
b111 6
19
1>
1C
b111 G
#573640000000
0!
0*
09
0>
0C
#573650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#573660000000
0!
0*
09
0>
0C
#573670000000
1!
1*
b1 6
19
1>
1C
b1 G
#573680000000
0!
0*
09
0>
0C
#573690000000
1!
1*
b10 6
19
1>
1C
b10 G
#573700000000
0!
0*
09
0>
0C
#573710000000
1!
1*
b11 6
19
1>
1C
b11 G
#573720000000
0!
0*
09
0>
0C
#573730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#573740000000
0!
0*
09
0>
0C
#573750000000
1!
1*
b101 6
19
1>
1C
b101 G
#573760000000
0!
0*
09
0>
0C
#573770000000
1!
1*
b110 6
19
1>
1C
b110 G
#573780000000
0!
0*
09
0>
0C
#573790000000
1!
1*
b111 6
19
1>
1C
b111 G
#573800000000
0!
0*
09
0>
0C
#573810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#573820000000
0!
0*
09
0>
0C
#573830000000
1!
1*
b1 6
19
1>
1C
b1 G
#573840000000
0!
0*
09
0>
0C
#573850000000
1!
1*
b10 6
19
1>
1C
b10 G
#573860000000
0!
0*
09
0>
0C
#573870000000
1!
1*
b11 6
19
1>
1C
b11 G
#573880000000
0!
0*
09
0>
0C
#573890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#573900000000
0!
0*
09
0>
0C
#573910000000
1!
1*
b101 6
19
1>
1C
b101 G
#573920000000
0!
0*
09
0>
0C
#573930000000
1!
1*
b110 6
19
1>
1C
b110 G
#573940000000
0!
0*
09
0>
0C
#573950000000
1!
1*
b111 6
19
1>
1C
b111 G
#573960000000
0!
1"
0*
1+
09
1:
0>
0C
#573970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#573980000000
0!
0*
09
0>
0C
#573990000000
1!
1*
b1 6
19
1>
1C
b1 G
#574000000000
0!
0*
09
0>
0C
#574010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#574020000000
0!
0*
09
0>
0C
#574030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#574040000000
0!
0*
09
0>
0C
#574050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#574060000000
0!
0*
09
0>
0C
#574070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#574080000000
0!
0#
0*
0,
09
0>
0?
0C
#574090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#574100000000
0!
0*
09
0>
0C
#574110000000
1!
1*
19
1>
1C
#574120000000
0!
0*
09
0>
0C
#574130000000
1!
1*
19
1>
1C
#574140000000
0!
0*
09
0>
0C
#574150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#574160000000
0!
0*
09
0>
0C
#574170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#574180000000
0!
0*
09
0>
0C
#574190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#574200000000
0!
0*
09
0>
0C
#574210000000
1!
1*
b10 6
19
1>
1C
b10 G
#574220000000
0!
0*
09
0>
0C
#574230000000
1!
1*
b11 6
19
1>
1C
b11 G
#574240000000
0!
0*
09
0>
0C
#574250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#574260000000
0!
0*
09
0>
0C
#574270000000
1!
1*
b101 6
19
1>
1C
b101 G
#574280000000
0!
0*
09
0>
0C
#574290000000
1!
1*
b110 6
19
1>
1C
b110 G
#574300000000
0!
0*
09
0>
0C
#574310000000
1!
1*
b111 6
19
1>
1C
b111 G
#574320000000
0!
0*
09
0>
0C
#574330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#574340000000
0!
0*
09
0>
0C
#574350000000
1!
1*
b1 6
19
1>
1C
b1 G
#574360000000
0!
0*
09
0>
0C
#574370000000
1!
1*
b10 6
19
1>
1C
b10 G
#574380000000
0!
0*
09
0>
0C
#574390000000
1!
1*
b11 6
19
1>
1C
b11 G
#574400000000
0!
0*
09
0>
0C
#574410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#574420000000
0!
0*
09
0>
0C
#574430000000
1!
1*
b101 6
19
1>
1C
b101 G
#574440000000
0!
0*
09
0>
0C
#574450000000
1!
1*
b110 6
19
1>
1C
b110 G
#574460000000
0!
0*
09
0>
0C
#574470000000
1!
1*
b111 6
19
1>
1C
b111 G
#574480000000
0!
0*
09
0>
0C
#574490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#574500000000
0!
0*
09
0>
0C
#574510000000
1!
1*
b1 6
19
1>
1C
b1 G
#574520000000
0!
0*
09
0>
0C
#574530000000
1!
1*
b10 6
19
1>
1C
b10 G
#574540000000
0!
0*
09
0>
0C
#574550000000
1!
1*
b11 6
19
1>
1C
b11 G
#574560000000
0!
0*
09
0>
0C
#574570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#574580000000
0!
0*
09
0>
0C
#574590000000
1!
1*
b101 6
19
1>
1C
b101 G
#574600000000
0!
0*
09
0>
0C
#574610000000
1!
1*
b110 6
19
1>
1C
b110 G
#574620000000
0!
0*
09
0>
0C
#574630000000
1!
1*
b111 6
19
1>
1C
b111 G
#574640000000
0!
1"
0*
1+
09
1:
0>
0C
#574650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#574660000000
0!
0*
09
0>
0C
#574670000000
1!
1*
b1 6
19
1>
1C
b1 G
#574680000000
0!
0*
09
0>
0C
#574690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#574700000000
0!
0*
09
0>
0C
#574710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#574720000000
0!
0*
09
0>
0C
#574730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#574740000000
0!
0*
09
0>
0C
#574750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#574760000000
0!
0#
0*
0,
09
0>
0?
0C
#574770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#574780000000
0!
0*
09
0>
0C
#574790000000
1!
1*
19
1>
1C
#574800000000
0!
0*
09
0>
0C
#574810000000
1!
1*
19
1>
1C
#574820000000
0!
0*
09
0>
0C
#574830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#574840000000
0!
0*
09
0>
0C
#574850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#574860000000
0!
0*
09
0>
0C
#574870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#574880000000
0!
0*
09
0>
0C
#574890000000
1!
1*
b10 6
19
1>
1C
b10 G
#574900000000
0!
0*
09
0>
0C
#574910000000
1!
1*
b11 6
19
1>
1C
b11 G
#574920000000
0!
0*
09
0>
0C
#574930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#574940000000
0!
0*
09
0>
0C
#574950000000
1!
1*
b101 6
19
1>
1C
b101 G
#574960000000
0!
0*
09
0>
0C
#574970000000
1!
1*
b110 6
19
1>
1C
b110 G
#574980000000
0!
0*
09
0>
0C
#574990000000
1!
1*
b111 6
19
1>
1C
b111 G
#575000000000
0!
0*
09
0>
0C
#575010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#575020000000
0!
0*
09
0>
0C
#575030000000
1!
1*
b1 6
19
1>
1C
b1 G
#575040000000
0!
0*
09
0>
0C
#575050000000
1!
1*
b10 6
19
1>
1C
b10 G
#575060000000
0!
0*
09
0>
0C
#575070000000
1!
1*
b11 6
19
1>
1C
b11 G
#575080000000
0!
0*
09
0>
0C
#575090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#575100000000
0!
0*
09
0>
0C
#575110000000
1!
1*
b101 6
19
1>
1C
b101 G
#575120000000
0!
0*
09
0>
0C
#575130000000
1!
1*
b110 6
19
1>
1C
b110 G
#575140000000
0!
0*
09
0>
0C
#575150000000
1!
1*
b111 6
19
1>
1C
b111 G
#575160000000
0!
0*
09
0>
0C
#575170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#575180000000
0!
0*
09
0>
0C
#575190000000
1!
1*
b1 6
19
1>
1C
b1 G
#575200000000
0!
0*
09
0>
0C
#575210000000
1!
1*
b10 6
19
1>
1C
b10 G
#575220000000
0!
0*
09
0>
0C
#575230000000
1!
1*
b11 6
19
1>
1C
b11 G
#575240000000
0!
0*
09
0>
0C
#575250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#575260000000
0!
0*
09
0>
0C
#575270000000
1!
1*
b101 6
19
1>
1C
b101 G
#575280000000
0!
0*
09
0>
0C
#575290000000
1!
1*
b110 6
19
1>
1C
b110 G
#575300000000
0!
0*
09
0>
0C
#575310000000
1!
1*
b111 6
19
1>
1C
b111 G
#575320000000
0!
1"
0*
1+
09
1:
0>
0C
#575330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#575340000000
0!
0*
09
0>
0C
#575350000000
1!
1*
b1 6
19
1>
1C
b1 G
#575360000000
0!
0*
09
0>
0C
#575370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#575380000000
0!
0*
09
0>
0C
#575390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#575400000000
0!
0*
09
0>
0C
#575410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#575420000000
0!
0*
09
0>
0C
#575430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#575440000000
0!
0#
0*
0,
09
0>
0?
0C
#575450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#575460000000
0!
0*
09
0>
0C
#575470000000
1!
1*
19
1>
1C
#575480000000
0!
0*
09
0>
0C
#575490000000
1!
1*
19
1>
1C
#575500000000
0!
0*
09
0>
0C
#575510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#575520000000
0!
0*
09
0>
0C
#575530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#575540000000
0!
0*
09
0>
0C
#575550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#575560000000
0!
0*
09
0>
0C
#575570000000
1!
1*
b10 6
19
1>
1C
b10 G
#575580000000
0!
0*
09
0>
0C
#575590000000
1!
1*
b11 6
19
1>
1C
b11 G
#575600000000
0!
0*
09
0>
0C
#575610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#575620000000
0!
0*
09
0>
0C
#575630000000
1!
1*
b101 6
19
1>
1C
b101 G
#575640000000
0!
0*
09
0>
0C
#575650000000
1!
1*
b110 6
19
1>
1C
b110 G
#575660000000
0!
0*
09
0>
0C
#575670000000
1!
1*
b111 6
19
1>
1C
b111 G
#575680000000
0!
0*
09
0>
0C
#575690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#575700000000
0!
0*
09
0>
0C
#575710000000
1!
1*
b1 6
19
1>
1C
b1 G
#575720000000
0!
0*
09
0>
0C
#575730000000
1!
1*
b10 6
19
1>
1C
b10 G
#575740000000
0!
0*
09
0>
0C
#575750000000
1!
1*
b11 6
19
1>
1C
b11 G
#575760000000
0!
0*
09
0>
0C
#575770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#575780000000
0!
0*
09
0>
0C
#575790000000
1!
1*
b101 6
19
1>
1C
b101 G
#575800000000
0!
0*
09
0>
0C
#575810000000
1!
1*
b110 6
19
1>
1C
b110 G
#575820000000
0!
0*
09
0>
0C
#575830000000
1!
1*
b111 6
19
1>
1C
b111 G
#575840000000
0!
0*
09
0>
0C
#575850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#575860000000
0!
0*
09
0>
0C
#575870000000
1!
1*
b1 6
19
1>
1C
b1 G
#575880000000
0!
0*
09
0>
0C
#575890000000
1!
1*
b10 6
19
1>
1C
b10 G
#575900000000
0!
0*
09
0>
0C
#575910000000
1!
1*
b11 6
19
1>
1C
b11 G
#575920000000
0!
0*
09
0>
0C
#575930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#575940000000
0!
0*
09
0>
0C
#575950000000
1!
1*
b101 6
19
1>
1C
b101 G
#575960000000
0!
0*
09
0>
0C
#575970000000
1!
1*
b110 6
19
1>
1C
b110 G
#575980000000
0!
0*
09
0>
0C
#575990000000
1!
1*
b111 6
19
1>
1C
b111 G
#576000000000
0!
1"
0*
1+
09
1:
0>
0C
#576010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#576020000000
0!
0*
09
0>
0C
#576030000000
1!
1*
b1 6
19
1>
1C
b1 G
#576040000000
0!
0*
09
0>
0C
#576050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#576060000000
0!
0*
09
0>
0C
#576070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#576080000000
0!
0*
09
0>
0C
#576090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#576100000000
0!
0*
09
0>
0C
#576110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#576120000000
0!
0#
0*
0,
09
0>
0?
0C
#576130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#576140000000
0!
0*
09
0>
0C
#576150000000
1!
1*
19
1>
1C
#576160000000
0!
0*
09
0>
0C
#576170000000
1!
1*
19
1>
1C
#576180000000
0!
0*
09
0>
0C
#576190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#576200000000
0!
0*
09
0>
0C
#576210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#576220000000
0!
0*
09
0>
0C
#576230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#576240000000
0!
0*
09
0>
0C
#576250000000
1!
1*
b10 6
19
1>
1C
b10 G
#576260000000
0!
0*
09
0>
0C
#576270000000
1!
1*
b11 6
19
1>
1C
b11 G
#576280000000
0!
0*
09
0>
0C
#576290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#576300000000
0!
0*
09
0>
0C
#576310000000
1!
1*
b101 6
19
1>
1C
b101 G
#576320000000
0!
0*
09
0>
0C
#576330000000
1!
1*
b110 6
19
1>
1C
b110 G
#576340000000
0!
0*
09
0>
0C
#576350000000
1!
1*
b111 6
19
1>
1C
b111 G
#576360000000
0!
0*
09
0>
0C
#576370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#576380000000
0!
0*
09
0>
0C
#576390000000
1!
1*
b1 6
19
1>
1C
b1 G
#576400000000
0!
0*
09
0>
0C
#576410000000
1!
1*
b10 6
19
1>
1C
b10 G
#576420000000
0!
0*
09
0>
0C
#576430000000
1!
1*
b11 6
19
1>
1C
b11 G
#576440000000
0!
0*
09
0>
0C
#576450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#576460000000
0!
0*
09
0>
0C
#576470000000
1!
1*
b101 6
19
1>
1C
b101 G
#576480000000
0!
0*
09
0>
0C
#576490000000
1!
1*
b110 6
19
1>
1C
b110 G
#576500000000
0!
0*
09
0>
0C
#576510000000
1!
1*
b111 6
19
1>
1C
b111 G
#576520000000
0!
0*
09
0>
0C
#576530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#576540000000
0!
0*
09
0>
0C
#576550000000
1!
1*
b1 6
19
1>
1C
b1 G
#576560000000
0!
0*
09
0>
0C
#576570000000
1!
1*
b10 6
19
1>
1C
b10 G
#576580000000
0!
0*
09
0>
0C
#576590000000
1!
1*
b11 6
19
1>
1C
b11 G
#576600000000
0!
0*
09
0>
0C
#576610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#576620000000
0!
0*
09
0>
0C
#576630000000
1!
1*
b101 6
19
1>
1C
b101 G
#576640000000
0!
0*
09
0>
0C
#576650000000
1!
1*
b110 6
19
1>
1C
b110 G
#576660000000
0!
0*
09
0>
0C
#576670000000
1!
1*
b111 6
19
1>
1C
b111 G
#576680000000
0!
1"
0*
1+
09
1:
0>
0C
#576690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#576700000000
0!
0*
09
0>
0C
#576710000000
1!
1*
b1 6
19
1>
1C
b1 G
#576720000000
0!
0*
09
0>
0C
#576730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#576740000000
0!
0*
09
0>
0C
#576750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#576760000000
0!
0*
09
0>
0C
#576770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#576780000000
0!
0*
09
0>
0C
#576790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#576800000000
0!
0#
0*
0,
09
0>
0?
0C
#576810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#576820000000
0!
0*
09
0>
0C
#576830000000
1!
1*
19
1>
1C
#576840000000
0!
0*
09
0>
0C
#576850000000
1!
1*
19
1>
1C
#576860000000
0!
0*
09
0>
0C
#576870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#576880000000
0!
0*
09
0>
0C
#576890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#576900000000
0!
0*
09
0>
0C
#576910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#576920000000
0!
0*
09
0>
0C
#576930000000
1!
1*
b10 6
19
1>
1C
b10 G
#576940000000
0!
0*
09
0>
0C
#576950000000
1!
1*
b11 6
19
1>
1C
b11 G
#576960000000
0!
0*
09
0>
0C
#576970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#576980000000
0!
0*
09
0>
0C
#576990000000
1!
1*
b101 6
19
1>
1C
b101 G
#577000000000
0!
0*
09
0>
0C
#577010000000
1!
1*
b110 6
19
1>
1C
b110 G
#577020000000
0!
0*
09
0>
0C
#577030000000
1!
1*
b111 6
19
1>
1C
b111 G
#577040000000
0!
0*
09
0>
0C
#577050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#577060000000
0!
0*
09
0>
0C
#577070000000
1!
1*
b1 6
19
1>
1C
b1 G
#577080000000
0!
0*
09
0>
0C
#577090000000
1!
1*
b10 6
19
1>
1C
b10 G
#577100000000
0!
0*
09
0>
0C
#577110000000
1!
1*
b11 6
19
1>
1C
b11 G
#577120000000
0!
0*
09
0>
0C
#577130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#577140000000
0!
0*
09
0>
0C
#577150000000
1!
1*
b101 6
19
1>
1C
b101 G
#577160000000
0!
0*
09
0>
0C
#577170000000
1!
1*
b110 6
19
1>
1C
b110 G
#577180000000
0!
0*
09
0>
0C
#577190000000
1!
1*
b111 6
19
1>
1C
b111 G
#577200000000
0!
0*
09
0>
0C
#577210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#577220000000
0!
0*
09
0>
0C
#577230000000
1!
1*
b1 6
19
1>
1C
b1 G
#577240000000
0!
0*
09
0>
0C
#577250000000
1!
1*
b10 6
19
1>
1C
b10 G
#577260000000
0!
0*
09
0>
0C
#577270000000
1!
1*
b11 6
19
1>
1C
b11 G
#577280000000
0!
0*
09
0>
0C
#577290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#577300000000
0!
0*
09
0>
0C
#577310000000
1!
1*
b101 6
19
1>
1C
b101 G
#577320000000
0!
0*
09
0>
0C
#577330000000
1!
1*
b110 6
19
1>
1C
b110 G
#577340000000
0!
0*
09
0>
0C
#577350000000
1!
1*
b111 6
19
1>
1C
b111 G
#577360000000
0!
1"
0*
1+
09
1:
0>
0C
#577370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#577380000000
0!
0*
09
0>
0C
#577390000000
1!
1*
b1 6
19
1>
1C
b1 G
#577400000000
0!
0*
09
0>
0C
#577410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#577420000000
0!
0*
09
0>
0C
#577430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#577440000000
0!
0*
09
0>
0C
#577450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#577460000000
0!
0*
09
0>
0C
#577470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#577480000000
0!
0#
0*
0,
09
0>
0?
0C
#577490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#577500000000
0!
0*
09
0>
0C
#577510000000
1!
1*
19
1>
1C
#577520000000
0!
0*
09
0>
0C
#577530000000
1!
1*
19
1>
1C
#577540000000
0!
0*
09
0>
0C
#577550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#577560000000
0!
0*
09
0>
0C
#577570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#577580000000
0!
0*
09
0>
0C
#577590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#577600000000
0!
0*
09
0>
0C
#577610000000
1!
1*
b10 6
19
1>
1C
b10 G
#577620000000
0!
0*
09
0>
0C
#577630000000
1!
1*
b11 6
19
1>
1C
b11 G
#577640000000
0!
0*
09
0>
0C
#577650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#577660000000
0!
0*
09
0>
0C
#577670000000
1!
1*
b101 6
19
1>
1C
b101 G
#577680000000
0!
0*
09
0>
0C
#577690000000
1!
1*
b110 6
19
1>
1C
b110 G
#577700000000
0!
0*
09
0>
0C
#577710000000
1!
1*
b111 6
19
1>
1C
b111 G
#577720000000
0!
0*
09
0>
0C
#577730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#577740000000
0!
0*
09
0>
0C
#577750000000
1!
1*
b1 6
19
1>
1C
b1 G
#577760000000
0!
0*
09
0>
0C
#577770000000
1!
1*
b10 6
19
1>
1C
b10 G
#577780000000
0!
0*
09
0>
0C
#577790000000
1!
1*
b11 6
19
1>
1C
b11 G
#577800000000
0!
0*
09
0>
0C
#577810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#577820000000
0!
0*
09
0>
0C
#577830000000
1!
1*
b101 6
19
1>
1C
b101 G
#577840000000
0!
0*
09
0>
0C
#577850000000
1!
1*
b110 6
19
1>
1C
b110 G
#577860000000
0!
0*
09
0>
0C
#577870000000
1!
1*
b111 6
19
1>
1C
b111 G
#577880000000
0!
0*
09
0>
0C
#577890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#577900000000
0!
0*
09
0>
0C
#577910000000
1!
1*
b1 6
19
1>
1C
b1 G
#577920000000
0!
0*
09
0>
0C
#577930000000
1!
1*
b10 6
19
1>
1C
b10 G
#577940000000
0!
0*
09
0>
0C
#577950000000
1!
1*
b11 6
19
1>
1C
b11 G
#577960000000
0!
0*
09
0>
0C
#577970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#577980000000
0!
0*
09
0>
0C
#577990000000
1!
1*
b101 6
19
1>
1C
b101 G
#578000000000
0!
0*
09
0>
0C
#578010000000
1!
1*
b110 6
19
1>
1C
b110 G
#578020000000
0!
0*
09
0>
0C
#578030000000
1!
1*
b111 6
19
1>
1C
b111 G
#578040000000
0!
1"
0*
1+
09
1:
0>
0C
#578050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#578060000000
0!
0*
09
0>
0C
#578070000000
1!
1*
b1 6
19
1>
1C
b1 G
#578080000000
0!
0*
09
0>
0C
#578090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#578100000000
0!
0*
09
0>
0C
#578110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#578120000000
0!
0*
09
0>
0C
#578130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#578140000000
0!
0*
09
0>
0C
#578150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#578160000000
0!
0#
0*
0,
09
0>
0?
0C
#578170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#578180000000
0!
0*
09
0>
0C
#578190000000
1!
1*
19
1>
1C
#578200000000
0!
0*
09
0>
0C
#578210000000
1!
1*
19
1>
1C
#578220000000
0!
0*
09
0>
0C
#578230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#578240000000
0!
0*
09
0>
0C
#578250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#578260000000
0!
0*
09
0>
0C
#578270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#578280000000
0!
0*
09
0>
0C
#578290000000
1!
1*
b10 6
19
1>
1C
b10 G
#578300000000
0!
0*
09
0>
0C
#578310000000
1!
1*
b11 6
19
1>
1C
b11 G
#578320000000
0!
0*
09
0>
0C
#578330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#578340000000
0!
0*
09
0>
0C
#578350000000
1!
1*
b101 6
19
1>
1C
b101 G
#578360000000
0!
0*
09
0>
0C
#578370000000
1!
1*
b110 6
19
1>
1C
b110 G
#578380000000
0!
0*
09
0>
0C
#578390000000
1!
1*
b111 6
19
1>
1C
b111 G
#578400000000
0!
0*
09
0>
0C
#578410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#578420000000
0!
0*
09
0>
0C
#578430000000
1!
1*
b1 6
19
1>
1C
b1 G
#578440000000
0!
0*
09
0>
0C
#578450000000
1!
1*
b10 6
19
1>
1C
b10 G
#578460000000
0!
0*
09
0>
0C
#578470000000
1!
1*
b11 6
19
1>
1C
b11 G
#578480000000
0!
0*
09
0>
0C
#578490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#578500000000
0!
0*
09
0>
0C
#578510000000
1!
1*
b101 6
19
1>
1C
b101 G
#578520000000
0!
0*
09
0>
0C
#578530000000
1!
1*
b110 6
19
1>
1C
b110 G
#578540000000
0!
0*
09
0>
0C
#578550000000
1!
1*
b111 6
19
1>
1C
b111 G
#578560000000
0!
0*
09
0>
0C
#578570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#578580000000
0!
0*
09
0>
0C
#578590000000
1!
1*
b1 6
19
1>
1C
b1 G
#578600000000
0!
0*
09
0>
0C
#578610000000
1!
1*
b10 6
19
1>
1C
b10 G
#578620000000
0!
0*
09
0>
0C
#578630000000
1!
1*
b11 6
19
1>
1C
b11 G
#578640000000
0!
0*
09
0>
0C
#578650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#578660000000
0!
0*
09
0>
0C
#578670000000
1!
1*
b101 6
19
1>
1C
b101 G
#578680000000
0!
0*
09
0>
0C
#578690000000
1!
1*
b110 6
19
1>
1C
b110 G
#578700000000
0!
0*
09
0>
0C
#578710000000
1!
1*
b111 6
19
1>
1C
b111 G
#578720000000
0!
1"
0*
1+
09
1:
0>
0C
#578730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#578740000000
0!
0*
09
0>
0C
#578750000000
1!
1*
b1 6
19
1>
1C
b1 G
#578760000000
0!
0*
09
0>
0C
#578770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#578780000000
0!
0*
09
0>
0C
#578790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#578800000000
0!
0*
09
0>
0C
#578810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#578820000000
0!
0*
09
0>
0C
#578830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#578840000000
0!
0#
0*
0,
09
0>
0?
0C
#578850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#578860000000
0!
0*
09
0>
0C
#578870000000
1!
1*
19
1>
1C
#578880000000
0!
0*
09
0>
0C
#578890000000
1!
1*
19
1>
1C
#578900000000
0!
0*
09
0>
0C
#578910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#578920000000
0!
0*
09
0>
0C
#578930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#578940000000
0!
0*
09
0>
0C
#578950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#578960000000
0!
0*
09
0>
0C
#578970000000
1!
1*
b10 6
19
1>
1C
b10 G
#578980000000
0!
0*
09
0>
0C
#578990000000
1!
1*
b11 6
19
1>
1C
b11 G
#579000000000
0!
0*
09
0>
0C
#579010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#579020000000
0!
0*
09
0>
0C
#579030000000
1!
1*
b101 6
19
1>
1C
b101 G
#579040000000
0!
0*
09
0>
0C
#579050000000
1!
1*
b110 6
19
1>
1C
b110 G
#579060000000
0!
0*
09
0>
0C
#579070000000
1!
1*
b111 6
19
1>
1C
b111 G
#579080000000
0!
0*
09
0>
0C
#579090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#579100000000
0!
0*
09
0>
0C
#579110000000
1!
1*
b1 6
19
1>
1C
b1 G
#579120000000
0!
0*
09
0>
0C
#579130000000
1!
1*
b10 6
19
1>
1C
b10 G
#579140000000
0!
0*
09
0>
0C
#579150000000
1!
1*
b11 6
19
1>
1C
b11 G
#579160000000
0!
0*
09
0>
0C
#579170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#579180000000
0!
0*
09
0>
0C
#579190000000
1!
1*
b101 6
19
1>
1C
b101 G
#579200000000
0!
0*
09
0>
0C
#579210000000
1!
1*
b110 6
19
1>
1C
b110 G
#579220000000
0!
0*
09
0>
0C
#579230000000
1!
1*
b111 6
19
1>
1C
b111 G
#579240000000
0!
0*
09
0>
0C
#579250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#579260000000
0!
0*
09
0>
0C
#579270000000
1!
1*
b1 6
19
1>
1C
b1 G
#579280000000
0!
0*
09
0>
0C
#579290000000
1!
1*
b10 6
19
1>
1C
b10 G
#579300000000
0!
0*
09
0>
0C
#579310000000
1!
1*
b11 6
19
1>
1C
b11 G
#579320000000
0!
0*
09
0>
0C
#579330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#579340000000
0!
0*
09
0>
0C
#579350000000
1!
1*
b101 6
19
1>
1C
b101 G
#579360000000
0!
0*
09
0>
0C
#579370000000
1!
1*
b110 6
19
1>
1C
b110 G
#579380000000
0!
0*
09
0>
0C
#579390000000
1!
1*
b111 6
19
1>
1C
b111 G
#579400000000
0!
1"
0*
1+
09
1:
0>
0C
#579410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#579420000000
0!
0*
09
0>
0C
#579430000000
1!
1*
b1 6
19
1>
1C
b1 G
#579440000000
0!
0*
09
0>
0C
#579450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#579460000000
0!
0*
09
0>
0C
#579470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#579480000000
0!
0*
09
0>
0C
#579490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#579500000000
0!
0*
09
0>
0C
#579510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#579520000000
0!
0#
0*
0,
09
0>
0?
0C
#579530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#579540000000
0!
0*
09
0>
0C
#579550000000
1!
1*
19
1>
1C
#579560000000
0!
0*
09
0>
0C
#579570000000
1!
1*
19
1>
1C
#579580000000
0!
0*
09
0>
0C
#579590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#579600000000
0!
0*
09
0>
0C
#579610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#579620000000
0!
0*
09
0>
0C
#579630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#579640000000
0!
0*
09
0>
0C
#579650000000
1!
1*
b10 6
19
1>
1C
b10 G
#579660000000
0!
0*
09
0>
0C
#579670000000
1!
1*
b11 6
19
1>
1C
b11 G
#579680000000
0!
0*
09
0>
0C
#579690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#579700000000
0!
0*
09
0>
0C
#579710000000
1!
1*
b101 6
19
1>
1C
b101 G
#579720000000
0!
0*
09
0>
0C
#579730000000
1!
1*
b110 6
19
1>
1C
b110 G
#579740000000
0!
0*
09
0>
0C
#579750000000
1!
1*
b111 6
19
1>
1C
b111 G
#579760000000
0!
0*
09
0>
0C
#579770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#579780000000
0!
0*
09
0>
0C
#579790000000
1!
1*
b1 6
19
1>
1C
b1 G
#579800000000
0!
0*
09
0>
0C
#579810000000
1!
1*
b10 6
19
1>
1C
b10 G
#579820000000
0!
0*
09
0>
0C
#579830000000
1!
1*
b11 6
19
1>
1C
b11 G
#579840000000
0!
0*
09
0>
0C
#579850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#579860000000
0!
0*
09
0>
0C
#579870000000
1!
1*
b101 6
19
1>
1C
b101 G
#579880000000
0!
0*
09
0>
0C
#579890000000
1!
1*
b110 6
19
1>
1C
b110 G
#579900000000
0!
0*
09
0>
0C
#579910000000
1!
1*
b111 6
19
1>
1C
b111 G
#579920000000
0!
0*
09
0>
0C
#579930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#579940000000
0!
0*
09
0>
0C
#579950000000
1!
1*
b1 6
19
1>
1C
b1 G
#579960000000
0!
0*
09
0>
0C
#579970000000
1!
1*
b10 6
19
1>
1C
b10 G
#579980000000
0!
0*
09
0>
0C
#579990000000
1!
1*
b11 6
19
1>
1C
b11 G
#580000000000
0!
0*
09
0>
0C
#580010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#580020000000
0!
0*
09
0>
0C
#580030000000
1!
1*
b101 6
19
1>
1C
b101 G
#580040000000
0!
0*
09
0>
0C
#580050000000
1!
1*
b110 6
19
1>
1C
b110 G
#580060000000
0!
0*
09
0>
0C
#580070000000
1!
1*
b111 6
19
1>
1C
b111 G
#580080000000
0!
1"
0*
1+
09
1:
0>
0C
#580090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#580100000000
0!
0*
09
0>
0C
#580110000000
1!
1*
b1 6
19
1>
1C
b1 G
#580120000000
0!
0*
09
0>
0C
#580130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#580140000000
0!
0*
09
0>
0C
#580150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#580160000000
0!
0*
09
0>
0C
#580170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#580180000000
0!
0*
09
0>
0C
#580190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#580200000000
0!
0#
0*
0,
09
0>
0?
0C
#580210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#580220000000
0!
0*
09
0>
0C
#580230000000
1!
1*
19
1>
1C
#580240000000
0!
0*
09
0>
0C
#580250000000
1!
1*
19
1>
1C
#580260000000
0!
0*
09
0>
0C
#580270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#580280000000
0!
0*
09
0>
0C
#580290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#580300000000
0!
0*
09
0>
0C
#580310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#580320000000
0!
0*
09
0>
0C
#580330000000
1!
1*
b10 6
19
1>
1C
b10 G
#580340000000
0!
0*
09
0>
0C
#580350000000
1!
1*
b11 6
19
1>
1C
b11 G
#580360000000
0!
0*
09
0>
0C
#580370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#580380000000
0!
0*
09
0>
0C
#580390000000
1!
1*
b101 6
19
1>
1C
b101 G
#580400000000
0!
0*
09
0>
0C
#580410000000
1!
1*
b110 6
19
1>
1C
b110 G
#580420000000
0!
0*
09
0>
0C
#580430000000
1!
1*
b111 6
19
1>
1C
b111 G
#580440000000
0!
0*
09
0>
0C
#580450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#580460000000
0!
0*
09
0>
0C
#580470000000
1!
1*
b1 6
19
1>
1C
b1 G
#580480000000
0!
0*
09
0>
0C
#580490000000
1!
1*
b10 6
19
1>
1C
b10 G
#580500000000
0!
0*
09
0>
0C
#580510000000
1!
1*
b11 6
19
1>
1C
b11 G
#580520000000
0!
0*
09
0>
0C
#580530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#580540000000
0!
0*
09
0>
0C
#580550000000
1!
1*
b101 6
19
1>
1C
b101 G
#580560000000
0!
0*
09
0>
0C
#580570000000
1!
1*
b110 6
19
1>
1C
b110 G
#580580000000
0!
0*
09
0>
0C
#580590000000
1!
1*
b111 6
19
1>
1C
b111 G
#580600000000
0!
0*
09
0>
0C
#580610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#580620000000
0!
0*
09
0>
0C
#580630000000
1!
1*
b1 6
19
1>
1C
b1 G
#580640000000
0!
0*
09
0>
0C
#580650000000
1!
1*
b10 6
19
1>
1C
b10 G
#580660000000
0!
0*
09
0>
0C
#580670000000
1!
1*
b11 6
19
1>
1C
b11 G
#580680000000
0!
0*
09
0>
0C
#580690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#580700000000
0!
0*
09
0>
0C
#580710000000
1!
1*
b101 6
19
1>
1C
b101 G
#580720000000
0!
0*
09
0>
0C
#580730000000
1!
1*
b110 6
19
1>
1C
b110 G
#580740000000
0!
0*
09
0>
0C
#580750000000
1!
1*
b111 6
19
1>
1C
b111 G
#580760000000
0!
1"
0*
1+
09
1:
0>
0C
#580770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#580780000000
0!
0*
09
0>
0C
#580790000000
1!
1*
b1 6
19
1>
1C
b1 G
#580800000000
0!
0*
09
0>
0C
#580810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#580820000000
0!
0*
09
0>
0C
#580830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#580840000000
0!
0*
09
0>
0C
#580850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#580860000000
0!
0*
09
0>
0C
#580870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#580880000000
0!
0#
0*
0,
09
0>
0?
0C
#580890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#580900000000
0!
0*
09
0>
0C
#580910000000
1!
1*
19
1>
1C
#580920000000
0!
0*
09
0>
0C
#580930000000
1!
1*
19
1>
1C
#580940000000
0!
0*
09
0>
0C
#580950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#580960000000
0!
0*
09
0>
0C
#580970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#580980000000
0!
0*
09
0>
0C
#580990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#581000000000
0!
0*
09
0>
0C
#581010000000
1!
1*
b10 6
19
1>
1C
b10 G
#581020000000
0!
0*
09
0>
0C
#581030000000
1!
1*
b11 6
19
1>
1C
b11 G
#581040000000
0!
0*
09
0>
0C
#581050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#581060000000
0!
0*
09
0>
0C
#581070000000
1!
1*
b101 6
19
1>
1C
b101 G
#581080000000
0!
0*
09
0>
0C
#581090000000
1!
1*
b110 6
19
1>
1C
b110 G
#581100000000
0!
0*
09
0>
0C
#581110000000
1!
1*
b111 6
19
1>
1C
b111 G
#581120000000
0!
0*
09
0>
0C
#581130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#581140000000
0!
0*
09
0>
0C
#581150000000
1!
1*
b1 6
19
1>
1C
b1 G
#581160000000
0!
0*
09
0>
0C
#581170000000
1!
1*
b10 6
19
1>
1C
b10 G
#581180000000
0!
0*
09
0>
0C
#581190000000
1!
1*
b11 6
19
1>
1C
b11 G
#581200000000
0!
0*
09
0>
0C
#581210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#581220000000
0!
0*
09
0>
0C
#581230000000
1!
1*
b101 6
19
1>
1C
b101 G
#581240000000
0!
0*
09
0>
0C
#581250000000
1!
1*
b110 6
19
1>
1C
b110 G
#581260000000
0!
0*
09
0>
0C
#581270000000
1!
1*
b111 6
19
1>
1C
b111 G
#581280000000
0!
0*
09
0>
0C
#581290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#581300000000
0!
0*
09
0>
0C
#581310000000
1!
1*
b1 6
19
1>
1C
b1 G
#581320000000
0!
0*
09
0>
0C
#581330000000
1!
1*
b10 6
19
1>
1C
b10 G
#581340000000
0!
0*
09
0>
0C
#581350000000
1!
1*
b11 6
19
1>
1C
b11 G
#581360000000
0!
0*
09
0>
0C
#581370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#581380000000
0!
0*
09
0>
0C
#581390000000
1!
1*
b101 6
19
1>
1C
b101 G
#581400000000
0!
0*
09
0>
0C
#581410000000
1!
1*
b110 6
19
1>
1C
b110 G
#581420000000
0!
0*
09
0>
0C
#581430000000
1!
1*
b111 6
19
1>
1C
b111 G
#581440000000
0!
1"
0*
1+
09
1:
0>
0C
#581450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#581460000000
0!
0*
09
0>
0C
#581470000000
1!
1*
b1 6
19
1>
1C
b1 G
#581480000000
0!
0*
09
0>
0C
#581490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#581500000000
0!
0*
09
0>
0C
#581510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#581520000000
0!
0*
09
0>
0C
#581530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#581540000000
0!
0*
09
0>
0C
#581550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#581560000000
0!
0#
0*
0,
09
0>
0?
0C
#581570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#581580000000
0!
0*
09
0>
0C
#581590000000
1!
1*
19
1>
1C
#581600000000
0!
0*
09
0>
0C
#581610000000
1!
1*
19
1>
1C
#581620000000
0!
0*
09
0>
0C
#581630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#581640000000
0!
0*
09
0>
0C
#581650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#581660000000
0!
0*
09
0>
0C
#581670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#581680000000
0!
0*
09
0>
0C
#581690000000
1!
1*
b10 6
19
1>
1C
b10 G
#581700000000
0!
0*
09
0>
0C
#581710000000
1!
1*
b11 6
19
1>
1C
b11 G
#581720000000
0!
0*
09
0>
0C
#581730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#581740000000
0!
0*
09
0>
0C
#581750000000
1!
1*
b101 6
19
1>
1C
b101 G
#581760000000
0!
0*
09
0>
0C
#581770000000
1!
1*
b110 6
19
1>
1C
b110 G
#581780000000
0!
0*
09
0>
0C
#581790000000
1!
1*
b111 6
19
1>
1C
b111 G
#581800000000
0!
0*
09
0>
0C
#581810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#581820000000
0!
0*
09
0>
0C
#581830000000
1!
1*
b1 6
19
1>
1C
b1 G
#581840000000
0!
0*
09
0>
0C
#581850000000
1!
1*
b10 6
19
1>
1C
b10 G
#581860000000
0!
0*
09
0>
0C
#581870000000
1!
1*
b11 6
19
1>
1C
b11 G
#581880000000
0!
0*
09
0>
0C
#581890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#581900000000
0!
0*
09
0>
0C
#581910000000
1!
1*
b101 6
19
1>
1C
b101 G
#581920000000
0!
0*
09
0>
0C
#581930000000
1!
1*
b110 6
19
1>
1C
b110 G
#581940000000
0!
0*
09
0>
0C
#581950000000
1!
1*
b111 6
19
1>
1C
b111 G
#581960000000
0!
0*
09
0>
0C
#581970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#581980000000
0!
0*
09
0>
0C
#581990000000
1!
1*
b1 6
19
1>
1C
b1 G
#582000000000
0!
0*
09
0>
0C
#582010000000
1!
1*
b10 6
19
1>
1C
b10 G
#582020000000
0!
0*
09
0>
0C
#582030000000
1!
1*
b11 6
19
1>
1C
b11 G
#582040000000
0!
0*
09
0>
0C
#582050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#582060000000
0!
0*
09
0>
0C
#582070000000
1!
1*
b101 6
19
1>
1C
b101 G
#582080000000
0!
0*
09
0>
0C
#582090000000
1!
1*
b110 6
19
1>
1C
b110 G
#582100000000
0!
0*
09
0>
0C
#582110000000
1!
1*
b111 6
19
1>
1C
b111 G
#582120000000
0!
1"
0*
1+
09
1:
0>
0C
#582130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#582140000000
0!
0*
09
0>
0C
#582150000000
1!
1*
b1 6
19
1>
1C
b1 G
#582160000000
0!
0*
09
0>
0C
#582170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#582180000000
0!
0*
09
0>
0C
#582190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#582200000000
0!
0*
09
0>
0C
#582210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#582220000000
0!
0*
09
0>
0C
#582230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#582240000000
0!
0#
0*
0,
09
0>
0?
0C
#582250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#582260000000
0!
0*
09
0>
0C
#582270000000
1!
1*
19
1>
1C
#582280000000
0!
0*
09
0>
0C
#582290000000
1!
1*
19
1>
1C
#582300000000
0!
0*
09
0>
0C
#582310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#582320000000
0!
0*
09
0>
0C
#582330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#582340000000
0!
0*
09
0>
0C
#582350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#582360000000
0!
0*
09
0>
0C
#582370000000
1!
1*
b10 6
19
1>
1C
b10 G
#582380000000
0!
0*
09
0>
0C
#582390000000
1!
1*
b11 6
19
1>
1C
b11 G
#582400000000
0!
0*
09
0>
0C
#582410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#582420000000
0!
0*
09
0>
0C
#582430000000
1!
1*
b101 6
19
1>
1C
b101 G
#582440000000
0!
0*
09
0>
0C
#582450000000
1!
1*
b110 6
19
1>
1C
b110 G
#582460000000
0!
0*
09
0>
0C
#582470000000
1!
1*
b111 6
19
1>
1C
b111 G
#582480000000
0!
0*
09
0>
0C
#582490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#582500000000
0!
0*
09
0>
0C
#582510000000
1!
1*
b1 6
19
1>
1C
b1 G
#582520000000
0!
0*
09
0>
0C
#582530000000
1!
1*
b10 6
19
1>
1C
b10 G
#582540000000
0!
0*
09
0>
0C
#582550000000
1!
1*
b11 6
19
1>
1C
b11 G
#582560000000
0!
0*
09
0>
0C
#582570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#582580000000
0!
0*
09
0>
0C
#582590000000
1!
1*
b101 6
19
1>
1C
b101 G
#582600000000
0!
0*
09
0>
0C
#582610000000
1!
1*
b110 6
19
1>
1C
b110 G
#582620000000
0!
0*
09
0>
0C
#582630000000
1!
1*
b111 6
19
1>
1C
b111 G
#582640000000
0!
0*
09
0>
0C
#582650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#582660000000
0!
0*
09
0>
0C
#582670000000
1!
1*
b1 6
19
1>
1C
b1 G
#582680000000
0!
0*
09
0>
0C
#582690000000
1!
1*
b10 6
19
1>
1C
b10 G
#582700000000
0!
0*
09
0>
0C
#582710000000
1!
1*
b11 6
19
1>
1C
b11 G
#582720000000
0!
0*
09
0>
0C
#582730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#582740000000
0!
0*
09
0>
0C
#582750000000
1!
1*
b101 6
19
1>
1C
b101 G
#582760000000
0!
0*
09
0>
0C
#582770000000
1!
1*
b110 6
19
1>
1C
b110 G
#582780000000
0!
0*
09
0>
0C
#582790000000
1!
1*
b111 6
19
1>
1C
b111 G
#582800000000
0!
1"
0*
1+
09
1:
0>
0C
#582810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#582820000000
0!
0*
09
0>
0C
#582830000000
1!
1*
b1 6
19
1>
1C
b1 G
#582840000000
0!
0*
09
0>
0C
#582850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#582860000000
0!
0*
09
0>
0C
#582870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#582880000000
0!
0*
09
0>
0C
#582890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#582900000000
0!
0*
09
0>
0C
#582910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#582920000000
0!
0#
0*
0,
09
0>
0?
0C
#582930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#582940000000
0!
0*
09
0>
0C
#582950000000
1!
1*
19
1>
1C
#582960000000
0!
0*
09
0>
0C
#582970000000
1!
1*
19
1>
1C
#582980000000
0!
0*
09
0>
0C
#582990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#583000000000
0!
0*
09
0>
0C
#583010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#583020000000
0!
0*
09
0>
0C
#583030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#583040000000
0!
0*
09
0>
0C
#583050000000
1!
1*
b10 6
19
1>
1C
b10 G
#583060000000
0!
0*
09
0>
0C
#583070000000
1!
1*
b11 6
19
1>
1C
b11 G
#583080000000
0!
0*
09
0>
0C
#583090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#583100000000
0!
0*
09
0>
0C
#583110000000
1!
1*
b101 6
19
1>
1C
b101 G
#583120000000
0!
0*
09
0>
0C
#583130000000
1!
1*
b110 6
19
1>
1C
b110 G
#583140000000
0!
0*
09
0>
0C
#583150000000
1!
1*
b111 6
19
1>
1C
b111 G
#583160000000
0!
0*
09
0>
0C
#583170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#583180000000
0!
0*
09
0>
0C
#583190000000
1!
1*
b1 6
19
1>
1C
b1 G
#583200000000
0!
0*
09
0>
0C
#583210000000
1!
1*
b10 6
19
1>
1C
b10 G
#583220000000
0!
0*
09
0>
0C
#583230000000
1!
1*
b11 6
19
1>
1C
b11 G
#583240000000
0!
0*
09
0>
0C
#583250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#583260000000
0!
0*
09
0>
0C
#583270000000
1!
1*
b101 6
19
1>
1C
b101 G
#583280000000
0!
0*
09
0>
0C
#583290000000
1!
1*
b110 6
19
1>
1C
b110 G
#583300000000
0!
0*
09
0>
0C
#583310000000
1!
1*
b111 6
19
1>
1C
b111 G
#583320000000
0!
0*
09
0>
0C
#583330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#583340000000
0!
0*
09
0>
0C
#583350000000
1!
1*
b1 6
19
1>
1C
b1 G
#583360000000
0!
0*
09
0>
0C
#583370000000
1!
1*
b10 6
19
1>
1C
b10 G
#583380000000
0!
0*
09
0>
0C
#583390000000
1!
1*
b11 6
19
1>
1C
b11 G
#583400000000
0!
0*
09
0>
0C
#583410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#583420000000
0!
0*
09
0>
0C
#583430000000
1!
1*
b101 6
19
1>
1C
b101 G
#583440000000
0!
0*
09
0>
0C
#583450000000
1!
1*
b110 6
19
1>
1C
b110 G
#583460000000
0!
0*
09
0>
0C
#583470000000
1!
1*
b111 6
19
1>
1C
b111 G
#583480000000
0!
1"
0*
1+
09
1:
0>
0C
#583490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#583500000000
0!
0*
09
0>
0C
#583510000000
1!
1*
b1 6
19
1>
1C
b1 G
#583520000000
0!
0*
09
0>
0C
#583530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#583540000000
0!
0*
09
0>
0C
#583550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#583560000000
0!
0*
09
0>
0C
#583570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#583580000000
0!
0*
09
0>
0C
#583590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#583600000000
0!
0#
0*
0,
09
0>
0?
0C
#583610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#583620000000
0!
0*
09
0>
0C
#583630000000
1!
1*
19
1>
1C
#583640000000
0!
0*
09
0>
0C
#583650000000
1!
1*
19
1>
1C
#583660000000
0!
0*
09
0>
0C
#583670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#583680000000
0!
0*
09
0>
0C
#583690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#583700000000
0!
0*
09
0>
0C
#583710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#583720000000
0!
0*
09
0>
0C
#583730000000
1!
1*
b10 6
19
1>
1C
b10 G
#583740000000
0!
0*
09
0>
0C
#583750000000
1!
1*
b11 6
19
1>
1C
b11 G
#583760000000
0!
0*
09
0>
0C
#583770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#583780000000
0!
0*
09
0>
0C
#583790000000
1!
1*
b101 6
19
1>
1C
b101 G
#583800000000
0!
0*
09
0>
0C
#583810000000
1!
1*
b110 6
19
1>
1C
b110 G
#583820000000
0!
0*
09
0>
0C
#583830000000
1!
1*
b111 6
19
1>
1C
b111 G
#583840000000
0!
0*
09
0>
0C
#583850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#583860000000
0!
0*
09
0>
0C
#583870000000
1!
1*
b1 6
19
1>
1C
b1 G
#583880000000
0!
0*
09
0>
0C
#583890000000
1!
1*
b10 6
19
1>
1C
b10 G
#583900000000
0!
0*
09
0>
0C
#583910000000
1!
1*
b11 6
19
1>
1C
b11 G
#583920000000
0!
0*
09
0>
0C
#583930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#583940000000
0!
0*
09
0>
0C
#583950000000
1!
1*
b101 6
19
1>
1C
b101 G
#583960000000
0!
0*
09
0>
0C
#583970000000
1!
1*
b110 6
19
1>
1C
b110 G
#583980000000
0!
0*
09
0>
0C
#583990000000
1!
1*
b111 6
19
1>
1C
b111 G
#584000000000
0!
0*
09
0>
0C
#584010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#584020000000
0!
0*
09
0>
0C
#584030000000
1!
1*
b1 6
19
1>
1C
b1 G
#584040000000
0!
0*
09
0>
0C
#584050000000
1!
1*
b10 6
19
1>
1C
b10 G
#584060000000
0!
0*
09
0>
0C
#584070000000
1!
1*
b11 6
19
1>
1C
b11 G
#584080000000
0!
0*
09
0>
0C
#584090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#584100000000
0!
0*
09
0>
0C
#584110000000
1!
1*
b101 6
19
1>
1C
b101 G
#584120000000
0!
0*
09
0>
0C
#584130000000
1!
1*
b110 6
19
1>
1C
b110 G
#584140000000
0!
0*
09
0>
0C
#584150000000
1!
1*
b111 6
19
1>
1C
b111 G
#584160000000
0!
1"
0*
1+
09
1:
0>
0C
#584170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#584180000000
0!
0*
09
0>
0C
#584190000000
1!
1*
b1 6
19
1>
1C
b1 G
#584200000000
0!
0*
09
0>
0C
#584210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#584220000000
0!
0*
09
0>
0C
#584230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#584240000000
0!
0*
09
0>
0C
#584250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#584260000000
0!
0*
09
0>
0C
#584270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#584280000000
0!
0#
0*
0,
09
0>
0?
0C
#584290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#584300000000
0!
0*
09
0>
0C
#584310000000
1!
1*
19
1>
1C
#584320000000
0!
0*
09
0>
0C
#584330000000
1!
1*
19
1>
1C
#584340000000
0!
0*
09
0>
0C
#584350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#584360000000
0!
0*
09
0>
0C
#584370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#584380000000
0!
0*
09
0>
0C
#584390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#584400000000
0!
0*
09
0>
0C
#584410000000
1!
1*
b10 6
19
1>
1C
b10 G
#584420000000
0!
0*
09
0>
0C
#584430000000
1!
1*
b11 6
19
1>
1C
b11 G
#584440000000
0!
0*
09
0>
0C
#584450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#584460000000
0!
0*
09
0>
0C
#584470000000
1!
1*
b101 6
19
1>
1C
b101 G
#584480000000
0!
0*
09
0>
0C
#584490000000
1!
1*
b110 6
19
1>
1C
b110 G
#584500000000
0!
0*
09
0>
0C
#584510000000
1!
1*
b111 6
19
1>
1C
b111 G
#584520000000
0!
0*
09
0>
0C
#584530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#584540000000
0!
0*
09
0>
0C
#584550000000
1!
1*
b1 6
19
1>
1C
b1 G
#584560000000
0!
0*
09
0>
0C
#584570000000
1!
1*
b10 6
19
1>
1C
b10 G
#584580000000
0!
0*
09
0>
0C
#584590000000
1!
1*
b11 6
19
1>
1C
b11 G
#584600000000
0!
0*
09
0>
0C
#584610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#584620000000
0!
0*
09
0>
0C
#584630000000
1!
1*
b101 6
19
1>
1C
b101 G
#584640000000
0!
0*
09
0>
0C
#584650000000
1!
1*
b110 6
19
1>
1C
b110 G
#584660000000
0!
0*
09
0>
0C
#584670000000
1!
1*
b111 6
19
1>
1C
b111 G
#584680000000
0!
0*
09
0>
0C
#584690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#584700000000
0!
0*
09
0>
0C
#584710000000
1!
1*
b1 6
19
1>
1C
b1 G
#584720000000
0!
0*
09
0>
0C
#584730000000
1!
1*
b10 6
19
1>
1C
b10 G
#584740000000
0!
0*
09
0>
0C
#584750000000
1!
1*
b11 6
19
1>
1C
b11 G
#584760000000
0!
0*
09
0>
0C
#584770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#584780000000
0!
0*
09
0>
0C
#584790000000
1!
1*
b101 6
19
1>
1C
b101 G
#584800000000
0!
0*
09
0>
0C
#584810000000
1!
1*
b110 6
19
1>
1C
b110 G
#584820000000
0!
0*
09
0>
0C
#584830000000
1!
1*
b111 6
19
1>
1C
b111 G
#584840000000
0!
1"
0*
1+
09
1:
0>
0C
#584850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#584860000000
0!
0*
09
0>
0C
#584870000000
1!
1*
b1 6
19
1>
1C
b1 G
#584880000000
0!
0*
09
0>
0C
#584890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#584900000000
0!
0*
09
0>
0C
#584910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#584920000000
0!
0*
09
0>
0C
#584930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#584940000000
0!
0*
09
0>
0C
#584950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#584960000000
0!
0#
0*
0,
09
0>
0?
0C
#584970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#584980000000
0!
0*
09
0>
0C
#584990000000
1!
1*
19
1>
1C
#585000000000
0!
0*
09
0>
0C
#585010000000
1!
1*
19
1>
1C
#585020000000
0!
0*
09
0>
0C
#585030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#585040000000
0!
0*
09
0>
0C
#585050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#585060000000
0!
0*
09
0>
0C
#585070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#585080000000
0!
0*
09
0>
0C
#585090000000
1!
1*
b10 6
19
1>
1C
b10 G
#585100000000
0!
0*
09
0>
0C
#585110000000
1!
1*
b11 6
19
1>
1C
b11 G
#585120000000
0!
0*
09
0>
0C
#585130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#585140000000
0!
0*
09
0>
0C
#585150000000
1!
1*
b101 6
19
1>
1C
b101 G
#585160000000
0!
0*
09
0>
0C
#585170000000
1!
1*
b110 6
19
1>
1C
b110 G
#585180000000
0!
0*
09
0>
0C
#585190000000
1!
1*
b111 6
19
1>
1C
b111 G
#585200000000
0!
0*
09
0>
0C
#585210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#585220000000
0!
0*
09
0>
0C
#585230000000
1!
1*
b1 6
19
1>
1C
b1 G
#585240000000
0!
0*
09
0>
0C
#585250000000
1!
1*
b10 6
19
1>
1C
b10 G
#585260000000
0!
0*
09
0>
0C
#585270000000
1!
1*
b11 6
19
1>
1C
b11 G
#585280000000
0!
0*
09
0>
0C
#585290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#585300000000
0!
0*
09
0>
0C
#585310000000
1!
1*
b101 6
19
1>
1C
b101 G
#585320000000
0!
0*
09
0>
0C
#585330000000
1!
1*
b110 6
19
1>
1C
b110 G
#585340000000
0!
0*
09
0>
0C
#585350000000
1!
1*
b111 6
19
1>
1C
b111 G
#585360000000
0!
0*
09
0>
0C
#585370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#585380000000
0!
0*
09
0>
0C
#585390000000
1!
1*
b1 6
19
1>
1C
b1 G
#585400000000
0!
0*
09
0>
0C
#585410000000
1!
1*
b10 6
19
1>
1C
b10 G
#585420000000
0!
0*
09
0>
0C
#585430000000
1!
1*
b11 6
19
1>
1C
b11 G
#585440000000
0!
0*
09
0>
0C
#585450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#585460000000
0!
0*
09
0>
0C
#585470000000
1!
1*
b101 6
19
1>
1C
b101 G
#585480000000
0!
0*
09
0>
0C
#585490000000
1!
1*
b110 6
19
1>
1C
b110 G
#585500000000
0!
0*
09
0>
0C
#585510000000
1!
1*
b111 6
19
1>
1C
b111 G
#585520000000
0!
1"
0*
1+
09
1:
0>
0C
#585530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#585540000000
0!
0*
09
0>
0C
#585550000000
1!
1*
b1 6
19
1>
1C
b1 G
#585560000000
0!
0*
09
0>
0C
#585570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#585580000000
0!
0*
09
0>
0C
#585590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#585600000000
0!
0*
09
0>
0C
#585610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#585620000000
0!
0*
09
0>
0C
#585630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#585640000000
0!
0#
0*
0,
09
0>
0?
0C
#585650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#585660000000
0!
0*
09
0>
0C
#585670000000
1!
1*
19
1>
1C
#585680000000
0!
0*
09
0>
0C
#585690000000
1!
1*
19
1>
1C
#585700000000
0!
0*
09
0>
0C
#585710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#585720000000
0!
0*
09
0>
0C
#585730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#585740000000
0!
0*
09
0>
0C
#585750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#585760000000
0!
0*
09
0>
0C
#585770000000
1!
1*
b10 6
19
1>
1C
b10 G
#585780000000
0!
0*
09
0>
0C
#585790000000
1!
1*
b11 6
19
1>
1C
b11 G
#585800000000
0!
0*
09
0>
0C
#585810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#585820000000
0!
0*
09
0>
0C
#585830000000
1!
1*
b101 6
19
1>
1C
b101 G
#585840000000
0!
0*
09
0>
0C
#585850000000
1!
1*
b110 6
19
1>
1C
b110 G
#585860000000
0!
0*
09
0>
0C
#585870000000
1!
1*
b111 6
19
1>
1C
b111 G
#585880000000
0!
0*
09
0>
0C
#585890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#585900000000
0!
0*
09
0>
0C
#585910000000
1!
1*
b1 6
19
1>
1C
b1 G
#585920000000
0!
0*
09
0>
0C
#585930000000
1!
1*
b10 6
19
1>
1C
b10 G
#585940000000
0!
0*
09
0>
0C
#585950000000
1!
1*
b11 6
19
1>
1C
b11 G
#585960000000
0!
0*
09
0>
0C
#585970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#585980000000
0!
0*
09
0>
0C
#585990000000
1!
1*
b101 6
19
1>
1C
b101 G
#586000000000
0!
0*
09
0>
0C
#586010000000
1!
1*
b110 6
19
1>
1C
b110 G
#586020000000
0!
0*
09
0>
0C
#586030000000
1!
1*
b111 6
19
1>
1C
b111 G
#586040000000
0!
0*
09
0>
0C
#586050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#586060000000
0!
0*
09
0>
0C
#586070000000
1!
1*
b1 6
19
1>
1C
b1 G
#586080000000
0!
0*
09
0>
0C
#586090000000
1!
1*
b10 6
19
1>
1C
b10 G
#586100000000
0!
0*
09
0>
0C
#586110000000
1!
1*
b11 6
19
1>
1C
b11 G
#586120000000
0!
0*
09
0>
0C
#586130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#586140000000
0!
0*
09
0>
0C
#586150000000
1!
1*
b101 6
19
1>
1C
b101 G
#586160000000
0!
0*
09
0>
0C
#586170000000
1!
1*
b110 6
19
1>
1C
b110 G
#586180000000
0!
0*
09
0>
0C
#586190000000
1!
1*
b111 6
19
1>
1C
b111 G
#586200000000
0!
1"
0*
1+
09
1:
0>
0C
#586210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#586220000000
0!
0*
09
0>
0C
#586230000000
1!
1*
b1 6
19
1>
1C
b1 G
#586240000000
0!
0*
09
0>
0C
#586250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#586260000000
0!
0*
09
0>
0C
#586270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#586280000000
0!
0*
09
0>
0C
#586290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#586300000000
0!
0*
09
0>
0C
#586310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#586320000000
0!
0#
0*
0,
09
0>
0?
0C
#586330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#586340000000
0!
0*
09
0>
0C
#586350000000
1!
1*
19
1>
1C
#586360000000
0!
0*
09
0>
0C
#586370000000
1!
1*
19
1>
1C
#586380000000
0!
0*
09
0>
0C
#586390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#586400000000
0!
0*
09
0>
0C
#586410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#586420000000
0!
0*
09
0>
0C
#586430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#586440000000
0!
0*
09
0>
0C
#586450000000
1!
1*
b10 6
19
1>
1C
b10 G
#586460000000
0!
0*
09
0>
0C
#586470000000
1!
1*
b11 6
19
1>
1C
b11 G
#586480000000
0!
0*
09
0>
0C
#586490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#586500000000
0!
0*
09
0>
0C
#586510000000
1!
1*
b101 6
19
1>
1C
b101 G
#586520000000
0!
0*
09
0>
0C
#586530000000
1!
1*
b110 6
19
1>
1C
b110 G
#586540000000
0!
0*
09
0>
0C
#586550000000
1!
1*
b111 6
19
1>
1C
b111 G
#586560000000
0!
0*
09
0>
0C
#586570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#586580000000
0!
0*
09
0>
0C
#586590000000
1!
1*
b1 6
19
1>
1C
b1 G
#586600000000
0!
0*
09
0>
0C
#586610000000
1!
1*
b10 6
19
1>
1C
b10 G
#586620000000
0!
0*
09
0>
0C
#586630000000
1!
1*
b11 6
19
1>
1C
b11 G
#586640000000
0!
0*
09
0>
0C
#586650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#586660000000
0!
0*
09
0>
0C
#586670000000
1!
1*
b101 6
19
1>
1C
b101 G
#586680000000
0!
0*
09
0>
0C
#586690000000
1!
1*
b110 6
19
1>
1C
b110 G
#586700000000
0!
0*
09
0>
0C
#586710000000
1!
1*
b111 6
19
1>
1C
b111 G
#586720000000
0!
0*
09
0>
0C
#586730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#586740000000
0!
0*
09
0>
0C
#586750000000
1!
1*
b1 6
19
1>
1C
b1 G
#586760000000
0!
0*
09
0>
0C
#586770000000
1!
1*
b10 6
19
1>
1C
b10 G
#586780000000
0!
0*
09
0>
0C
#586790000000
1!
1*
b11 6
19
1>
1C
b11 G
#586800000000
0!
0*
09
0>
0C
#586810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#586820000000
0!
0*
09
0>
0C
#586830000000
1!
1*
b101 6
19
1>
1C
b101 G
#586840000000
0!
0*
09
0>
0C
#586850000000
1!
1*
b110 6
19
1>
1C
b110 G
#586860000000
0!
0*
09
0>
0C
#586870000000
1!
1*
b111 6
19
1>
1C
b111 G
#586880000000
0!
1"
0*
1+
09
1:
0>
0C
#586890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#586900000000
0!
0*
09
0>
0C
#586910000000
1!
1*
b1 6
19
1>
1C
b1 G
#586920000000
0!
0*
09
0>
0C
#586930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#586940000000
0!
0*
09
0>
0C
#586950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#586960000000
0!
0*
09
0>
0C
#586970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#586980000000
0!
0*
09
0>
0C
#586990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#587000000000
0!
0#
0*
0,
09
0>
0?
0C
#587010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#587020000000
0!
0*
09
0>
0C
#587030000000
1!
1*
19
1>
1C
#587040000000
0!
0*
09
0>
0C
#587050000000
1!
1*
19
1>
1C
#587060000000
0!
0*
09
0>
0C
#587070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#587080000000
0!
0*
09
0>
0C
#587090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#587100000000
0!
0*
09
0>
0C
#587110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#587120000000
0!
0*
09
0>
0C
#587130000000
1!
1*
b10 6
19
1>
1C
b10 G
#587140000000
0!
0*
09
0>
0C
#587150000000
1!
1*
b11 6
19
1>
1C
b11 G
#587160000000
0!
0*
09
0>
0C
#587170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#587180000000
0!
0*
09
0>
0C
#587190000000
1!
1*
b101 6
19
1>
1C
b101 G
#587200000000
0!
0*
09
0>
0C
#587210000000
1!
1*
b110 6
19
1>
1C
b110 G
#587220000000
0!
0*
09
0>
0C
#587230000000
1!
1*
b111 6
19
1>
1C
b111 G
#587240000000
0!
0*
09
0>
0C
#587250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#587260000000
0!
0*
09
0>
0C
#587270000000
1!
1*
b1 6
19
1>
1C
b1 G
#587280000000
0!
0*
09
0>
0C
#587290000000
1!
1*
b10 6
19
1>
1C
b10 G
#587300000000
0!
0*
09
0>
0C
#587310000000
1!
1*
b11 6
19
1>
1C
b11 G
#587320000000
0!
0*
09
0>
0C
#587330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#587340000000
0!
0*
09
0>
0C
#587350000000
1!
1*
b101 6
19
1>
1C
b101 G
#587360000000
0!
0*
09
0>
0C
#587370000000
1!
1*
b110 6
19
1>
1C
b110 G
#587380000000
0!
0*
09
0>
0C
#587390000000
1!
1*
b111 6
19
1>
1C
b111 G
#587400000000
0!
0*
09
0>
0C
#587410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#587420000000
0!
0*
09
0>
0C
#587430000000
1!
1*
b1 6
19
1>
1C
b1 G
#587440000000
0!
0*
09
0>
0C
#587450000000
1!
1*
b10 6
19
1>
1C
b10 G
#587460000000
0!
0*
09
0>
0C
#587470000000
1!
1*
b11 6
19
1>
1C
b11 G
#587480000000
0!
0*
09
0>
0C
#587490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#587500000000
0!
0*
09
0>
0C
#587510000000
1!
1*
b101 6
19
1>
1C
b101 G
#587520000000
0!
0*
09
0>
0C
#587530000000
1!
1*
b110 6
19
1>
1C
b110 G
#587540000000
0!
0*
09
0>
0C
#587550000000
1!
1*
b111 6
19
1>
1C
b111 G
#587560000000
0!
1"
0*
1+
09
1:
0>
0C
#587570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#587580000000
0!
0*
09
0>
0C
#587590000000
1!
1*
b1 6
19
1>
1C
b1 G
#587600000000
0!
0*
09
0>
0C
#587610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#587620000000
0!
0*
09
0>
0C
#587630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#587640000000
0!
0*
09
0>
0C
#587650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#587660000000
0!
0*
09
0>
0C
#587670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#587680000000
0!
0#
0*
0,
09
0>
0?
0C
#587690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#587700000000
0!
0*
09
0>
0C
#587710000000
1!
1*
19
1>
1C
#587720000000
0!
0*
09
0>
0C
#587730000000
1!
1*
19
1>
1C
#587740000000
0!
0*
09
0>
0C
#587750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#587760000000
0!
0*
09
0>
0C
#587770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#587780000000
0!
0*
09
0>
0C
#587790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#587800000000
0!
0*
09
0>
0C
#587810000000
1!
1*
b10 6
19
1>
1C
b10 G
#587820000000
0!
0*
09
0>
0C
#587830000000
1!
1*
b11 6
19
1>
1C
b11 G
#587840000000
0!
0*
09
0>
0C
#587850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#587860000000
0!
0*
09
0>
0C
#587870000000
1!
1*
b101 6
19
1>
1C
b101 G
#587880000000
0!
0*
09
0>
0C
#587890000000
1!
1*
b110 6
19
1>
1C
b110 G
#587900000000
0!
0*
09
0>
0C
#587910000000
1!
1*
b111 6
19
1>
1C
b111 G
#587920000000
0!
0*
09
0>
0C
#587930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#587940000000
0!
0*
09
0>
0C
#587950000000
1!
1*
b1 6
19
1>
1C
b1 G
#587960000000
0!
0*
09
0>
0C
#587970000000
1!
1*
b10 6
19
1>
1C
b10 G
#587980000000
0!
0*
09
0>
0C
#587990000000
1!
1*
b11 6
19
1>
1C
b11 G
#588000000000
0!
0*
09
0>
0C
#588010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#588020000000
0!
0*
09
0>
0C
#588030000000
1!
1*
b101 6
19
1>
1C
b101 G
#588040000000
0!
0*
09
0>
0C
#588050000000
1!
1*
b110 6
19
1>
1C
b110 G
#588060000000
0!
0*
09
0>
0C
#588070000000
1!
1*
b111 6
19
1>
1C
b111 G
#588080000000
0!
0*
09
0>
0C
#588090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#588100000000
0!
0*
09
0>
0C
#588110000000
1!
1*
b1 6
19
1>
1C
b1 G
#588120000000
0!
0*
09
0>
0C
#588130000000
1!
1*
b10 6
19
1>
1C
b10 G
#588140000000
0!
0*
09
0>
0C
#588150000000
1!
1*
b11 6
19
1>
1C
b11 G
#588160000000
0!
0*
09
0>
0C
#588170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#588180000000
0!
0*
09
0>
0C
#588190000000
1!
1*
b101 6
19
1>
1C
b101 G
#588200000000
0!
0*
09
0>
0C
#588210000000
1!
1*
b110 6
19
1>
1C
b110 G
#588220000000
0!
0*
09
0>
0C
#588230000000
1!
1*
b111 6
19
1>
1C
b111 G
#588240000000
0!
1"
0*
1+
09
1:
0>
0C
#588250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#588260000000
0!
0*
09
0>
0C
#588270000000
1!
1*
b1 6
19
1>
1C
b1 G
#588280000000
0!
0*
09
0>
0C
#588290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#588300000000
0!
0*
09
0>
0C
#588310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#588320000000
0!
0*
09
0>
0C
#588330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#588340000000
0!
0*
09
0>
0C
#588350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#588360000000
0!
0#
0*
0,
09
0>
0?
0C
#588370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#588380000000
0!
0*
09
0>
0C
#588390000000
1!
1*
19
1>
1C
#588400000000
0!
0*
09
0>
0C
#588410000000
1!
1*
19
1>
1C
#588420000000
0!
0*
09
0>
0C
#588430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#588440000000
0!
0*
09
0>
0C
#588450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#588460000000
0!
0*
09
0>
0C
#588470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#588480000000
0!
0*
09
0>
0C
#588490000000
1!
1*
b10 6
19
1>
1C
b10 G
#588500000000
0!
0*
09
0>
0C
#588510000000
1!
1*
b11 6
19
1>
1C
b11 G
#588520000000
0!
0*
09
0>
0C
#588530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#588540000000
0!
0*
09
0>
0C
#588550000000
1!
1*
b101 6
19
1>
1C
b101 G
#588560000000
0!
0*
09
0>
0C
#588570000000
1!
1*
b110 6
19
1>
1C
b110 G
#588580000000
0!
0*
09
0>
0C
#588590000000
1!
1*
b111 6
19
1>
1C
b111 G
#588600000000
0!
0*
09
0>
0C
#588610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#588620000000
0!
0*
09
0>
0C
#588630000000
1!
1*
b1 6
19
1>
1C
b1 G
#588640000000
0!
0*
09
0>
0C
#588650000000
1!
1*
b10 6
19
1>
1C
b10 G
#588660000000
0!
0*
09
0>
0C
#588670000000
1!
1*
b11 6
19
1>
1C
b11 G
#588680000000
0!
0*
09
0>
0C
#588690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#588700000000
0!
0*
09
0>
0C
#588710000000
1!
1*
b101 6
19
1>
1C
b101 G
#588720000000
0!
0*
09
0>
0C
#588730000000
1!
1*
b110 6
19
1>
1C
b110 G
#588740000000
0!
0*
09
0>
0C
#588750000000
1!
1*
b111 6
19
1>
1C
b111 G
#588760000000
0!
0*
09
0>
0C
#588770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#588780000000
0!
0*
09
0>
0C
#588790000000
1!
1*
b1 6
19
1>
1C
b1 G
#588800000000
0!
0*
09
0>
0C
#588810000000
1!
1*
b10 6
19
1>
1C
b10 G
#588820000000
0!
0*
09
0>
0C
#588830000000
1!
1*
b11 6
19
1>
1C
b11 G
#588840000000
0!
0*
09
0>
0C
#588850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#588860000000
0!
0*
09
0>
0C
#588870000000
1!
1*
b101 6
19
1>
1C
b101 G
#588880000000
0!
0*
09
0>
0C
#588890000000
1!
1*
b110 6
19
1>
1C
b110 G
#588900000000
0!
0*
09
0>
0C
#588910000000
1!
1*
b111 6
19
1>
1C
b111 G
#588920000000
0!
1"
0*
1+
09
1:
0>
0C
#588930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#588940000000
0!
0*
09
0>
0C
#588950000000
1!
1*
b1 6
19
1>
1C
b1 G
#588960000000
0!
0*
09
0>
0C
#588970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#588980000000
0!
0*
09
0>
0C
#588990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#589000000000
0!
0*
09
0>
0C
#589010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#589020000000
0!
0*
09
0>
0C
#589030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#589040000000
0!
0#
0*
0,
09
0>
0?
0C
#589050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#589060000000
0!
0*
09
0>
0C
#589070000000
1!
1*
19
1>
1C
#589080000000
0!
0*
09
0>
0C
#589090000000
1!
1*
19
1>
1C
#589100000000
0!
0*
09
0>
0C
#589110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#589120000000
0!
0*
09
0>
0C
#589130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#589140000000
0!
0*
09
0>
0C
#589150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#589160000000
0!
0*
09
0>
0C
#589170000000
1!
1*
b10 6
19
1>
1C
b10 G
#589180000000
0!
0*
09
0>
0C
#589190000000
1!
1*
b11 6
19
1>
1C
b11 G
#589200000000
0!
0*
09
0>
0C
#589210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#589220000000
0!
0*
09
0>
0C
#589230000000
1!
1*
b101 6
19
1>
1C
b101 G
#589240000000
0!
0*
09
0>
0C
#589250000000
1!
1*
b110 6
19
1>
1C
b110 G
#589260000000
0!
0*
09
0>
0C
#589270000000
1!
1*
b111 6
19
1>
1C
b111 G
#589280000000
0!
0*
09
0>
0C
#589290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#589300000000
0!
0*
09
0>
0C
#589310000000
1!
1*
b1 6
19
1>
1C
b1 G
#589320000000
0!
0*
09
0>
0C
#589330000000
1!
1*
b10 6
19
1>
1C
b10 G
#589340000000
0!
0*
09
0>
0C
#589350000000
1!
1*
b11 6
19
1>
1C
b11 G
#589360000000
0!
0*
09
0>
0C
#589370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#589380000000
0!
0*
09
0>
0C
#589390000000
1!
1*
b101 6
19
1>
1C
b101 G
#589400000000
0!
0*
09
0>
0C
#589410000000
1!
1*
b110 6
19
1>
1C
b110 G
#589420000000
0!
0*
09
0>
0C
#589430000000
1!
1*
b111 6
19
1>
1C
b111 G
#589440000000
0!
0*
09
0>
0C
#589450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#589460000000
0!
0*
09
0>
0C
#589470000000
1!
1*
b1 6
19
1>
1C
b1 G
#589480000000
0!
0*
09
0>
0C
#589490000000
1!
1*
b10 6
19
1>
1C
b10 G
#589500000000
0!
0*
09
0>
0C
#589510000000
1!
1*
b11 6
19
1>
1C
b11 G
#589520000000
0!
0*
09
0>
0C
#589530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#589540000000
0!
0*
09
0>
0C
#589550000000
1!
1*
b101 6
19
1>
1C
b101 G
#589560000000
0!
0*
09
0>
0C
#589570000000
1!
1*
b110 6
19
1>
1C
b110 G
#589580000000
0!
0*
09
0>
0C
#589590000000
1!
1*
b111 6
19
1>
1C
b111 G
#589600000000
0!
1"
0*
1+
09
1:
0>
0C
#589610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#589620000000
0!
0*
09
0>
0C
#589630000000
1!
1*
b1 6
19
1>
1C
b1 G
#589640000000
0!
0*
09
0>
0C
#589650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#589660000000
0!
0*
09
0>
0C
#589670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#589680000000
0!
0*
09
0>
0C
#589690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#589700000000
0!
0*
09
0>
0C
#589710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#589720000000
0!
0#
0*
0,
09
0>
0?
0C
#589730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#589740000000
0!
0*
09
0>
0C
#589750000000
1!
1*
19
1>
1C
#589760000000
0!
0*
09
0>
0C
#589770000000
1!
1*
19
1>
1C
#589780000000
0!
0*
09
0>
0C
#589790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#589800000000
0!
0*
09
0>
0C
#589810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#589820000000
0!
0*
09
0>
0C
#589830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#589840000000
0!
0*
09
0>
0C
#589850000000
1!
1*
b10 6
19
1>
1C
b10 G
#589860000000
0!
0*
09
0>
0C
#589870000000
1!
1*
b11 6
19
1>
1C
b11 G
#589880000000
0!
0*
09
0>
0C
#589890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#589900000000
0!
0*
09
0>
0C
#589910000000
1!
1*
b101 6
19
1>
1C
b101 G
#589920000000
0!
0*
09
0>
0C
#589930000000
1!
1*
b110 6
19
1>
1C
b110 G
#589940000000
0!
0*
09
0>
0C
#589950000000
1!
1*
b111 6
19
1>
1C
b111 G
#589960000000
0!
0*
09
0>
0C
#589970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#589980000000
0!
0*
09
0>
0C
#589990000000
1!
1*
b1 6
19
1>
1C
b1 G
#590000000000
0!
0*
09
0>
0C
#590010000000
1!
1*
b10 6
19
1>
1C
b10 G
#590020000000
0!
0*
09
0>
0C
#590030000000
1!
1*
b11 6
19
1>
1C
b11 G
#590040000000
0!
0*
09
0>
0C
#590050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#590060000000
0!
0*
09
0>
0C
#590070000000
1!
1*
b101 6
19
1>
1C
b101 G
#590080000000
0!
0*
09
0>
0C
#590090000000
1!
1*
b110 6
19
1>
1C
b110 G
#590100000000
0!
0*
09
0>
0C
#590110000000
1!
1*
b111 6
19
1>
1C
b111 G
#590120000000
0!
0*
09
0>
0C
#590130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#590140000000
0!
0*
09
0>
0C
#590150000000
1!
1*
b1 6
19
1>
1C
b1 G
#590160000000
0!
0*
09
0>
0C
#590170000000
1!
1*
b10 6
19
1>
1C
b10 G
#590180000000
0!
0*
09
0>
0C
#590190000000
1!
1*
b11 6
19
1>
1C
b11 G
#590200000000
0!
0*
09
0>
0C
#590210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#590220000000
0!
0*
09
0>
0C
#590230000000
1!
1*
b101 6
19
1>
1C
b101 G
#590240000000
0!
0*
09
0>
0C
#590250000000
1!
1*
b110 6
19
1>
1C
b110 G
#590260000000
0!
0*
09
0>
0C
#590270000000
1!
1*
b111 6
19
1>
1C
b111 G
#590280000000
0!
1"
0*
1+
09
1:
0>
0C
#590290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#590300000000
0!
0*
09
0>
0C
#590310000000
1!
1*
b1 6
19
1>
1C
b1 G
#590320000000
0!
0*
09
0>
0C
#590330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#590340000000
0!
0*
09
0>
0C
#590350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#590360000000
0!
0*
09
0>
0C
#590370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#590380000000
0!
0*
09
0>
0C
#590390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#590400000000
0!
0#
0*
0,
09
0>
0?
0C
#590410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#590420000000
0!
0*
09
0>
0C
#590430000000
1!
1*
19
1>
1C
#590440000000
0!
0*
09
0>
0C
#590450000000
1!
1*
19
1>
1C
#590460000000
0!
0*
09
0>
0C
#590470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#590480000000
0!
0*
09
0>
0C
#590490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#590500000000
0!
0*
09
0>
0C
#590510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#590520000000
0!
0*
09
0>
0C
#590530000000
1!
1*
b10 6
19
1>
1C
b10 G
#590540000000
0!
0*
09
0>
0C
#590550000000
1!
1*
b11 6
19
1>
1C
b11 G
#590560000000
0!
0*
09
0>
0C
#590570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#590580000000
0!
0*
09
0>
0C
#590590000000
1!
1*
b101 6
19
1>
1C
b101 G
#590600000000
0!
0*
09
0>
0C
#590610000000
1!
1*
b110 6
19
1>
1C
b110 G
#590620000000
0!
0*
09
0>
0C
#590630000000
1!
1*
b111 6
19
1>
1C
b111 G
#590640000000
0!
0*
09
0>
0C
#590650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#590660000000
0!
0*
09
0>
0C
#590670000000
1!
1*
b1 6
19
1>
1C
b1 G
#590680000000
0!
0*
09
0>
0C
#590690000000
1!
1*
b10 6
19
1>
1C
b10 G
#590700000000
0!
0*
09
0>
0C
#590710000000
1!
1*
b11 6
19
1>
1C
b11 G
#590720000000
0!
0*
09
0>
0C
#590730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#590740000000
0!
0*
09
0>
0C
#590750000000
1!
1*
b101 6
19
1>
1C
b101 G
#590760000000
0!
0*
09
0>
0C
#590770000000
1!
1*
b110 6
19
1>
1C
b110 G
#590780000000
0!
0*
09
0>
0C
#590790000000
1!
1*
b111 6
19
1>
1C
b111 G
#590800000000
0!
0*
09
0>
0C
#590810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#590820000000
0!
0*
09
0>
0C
#590830000000
1!
1*
b1 6
19
1>
1C
b1 G
#590840000000
0!
0*
09
0>
0C
#590850000000
1!
1*
b10 6
19
1>
1C
b10 G
#590860000000
0!
0*
09
0>
0C
#590870000000
1!
1*
b11 6
19
1>
1C
b11 G
#590880000000
0!
0*
09
0>
0C
#590890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#590900000000
0!
0*
09
0>
0C
#590910000000
1!
1*
b101 6
19
1>
1C
b101 G
#590920000000
0!
0*
09
0>
0C
#590930000000
1!
1*
b110 6
19
1>
1C
b110 G
#590940000000
0!
0*
09
0>
0C
#590950000000
1!
1*
b111 6
19
1>
1C
b111 G
#590960000000
0!
1"
0*
1+
09
1:
0>
0C
#590970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#590980000000
0!
0*
09
0>
0C
#590990000000
1!
1*
b1 6
19
1>
1C
b1 G
#591000000000
0!
0*
09
0>
0C
#591010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#591020000000
0!
0*
09
0>
0C
#591030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#591040000000
0!
0*
09
0>
0C
#591050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#591060000000
0!
0*
09
0>
0C
#591070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#591080000000
0!
0#
0*
0,
09
0>
0?
0C
#591090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#591100000000
0!
0*
09
0>
0C
#591110000000
1!
1*
19
1>
1C
#591120000000
0!
0*
09
0>
0C
#591130000000
1!
1*
19
1>
1C
#591140000000
0!
0*
09
0>
0C
#591150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#591160000000
0!
0*
09
0>
0C
#591170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#591180000000
0!
0*
09
0>
0C
#591190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#591200000000
0!
0*
09
0>
0C
#591210000000
1!
1*
b10 6
19
1>
1C
b10 G
#591220000000
0!
0*
09
0>
0C
#591230000000
1!
1*
b11 6
19
1>
1C
b11 G
#591240000000
0!
0*
09
0>
0C
#591250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#591260000000
0!
0*
09
0>
0C
#591270000000
1!
1*
b101 6
19
1>
1C
b101 G
#591280000000
0!
0*
09
0>
0C
#591290000000
1!
1*
b110 6
19
1>
1C
b110 G
#591300000000
0!
0*
09
0>
0C
#591310000000
1!
1*
b111 6
19
1>
1C
b111 G
#591320000000
0!
0*
09
0>
0C
#591330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#591340000000
0!
0*
09
0>
0C
#591350000000
1!
1*
b1 6
19
1>
1C
b1 G
#591360000000
0!
0*
09
0>
0C
#591370000000
1!
1*
b10 6
19
1>
1C
b10 G
#591380000000
0!
0*
09
0>
0C
#591390000000
1!
1*
b11 6
19
1>
1C
b11 G
#591400000000
0!
0*
09
0>
0C
#591410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#591420000000
0!
0*
09
0>
0C
#591430000000
1!
1*
b101 6
19
1>
1C
b101 G
#591440000000
0!
0*
09
0>
0C
#591450000000
1!
1*
b110 6
19
1>
1C
b110 G
#591460000000
0!
0*
09
0>
0C
#591470000000
1!
1*
b111 6
19
1>
1C
b111 G
#591480000000
0!
0*
09
0>
0C
#591490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#591500000000
0!
0*
09
0>
0C
#591510000000
1!
1*
b1 6
19
1>
1C
b1 G
#591520000000
0!
0*
09
0>
0C
#591530000000
1!
1*
b10 6
19
1>
1C
b10 G
#591540000000
0!
0*
09
0>
0C
#591550000000
1!
1*
b11 6
19
1>
1C
b11 G
#591560000000
0!
0*
09
0>
0C
#591570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#591580000000
0!
0*
09
0>
0C
#591590000000
1!
1*
b101 6
19
1>
1C
b101 G
#591600000000
0!
0*
09
0>
0C
#591610000000
1!
1*
b110 6
19
1>
1C
b110 G
#591620000000
0!
0*
09
0>
0C
#591630000000
1!
1*
b111 6
19
1>
1C
b111 G
#591640000000
0!
1"
0*
1+
09
1:
0>
0C
#591650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#591660000000
0!
0*
09
0>
0C
#591670000000
1!
1*
b1 6
19
1>
1C
b1 G
#591680000000
0!
0*
09
0>
0C
#591690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#591700000000
0!
0*
09
0>
0C
#591710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#591720000000
0!
0*
09
0>
0C
#591730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#591740000000
0!
0*
09
0>
0C
#591750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#591760000000
0!
0#
0*
0,
09
0>
0?
0C
#591770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#591780000000
0!
0*
09
0>
0C
#591790000000
1!
1*
19
1>
1C
#591800000000
0!
0*
09
0>
0C
#591810000000
1!
1*
19
1>
1C
#591820000000
0!
0*
09
0>
0C
#591830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#591840000000
0!
0*
09
0>
0C
#591850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#591860000000
0!
0*
09
0>
0C
#591870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#591880000000
0!
0*
09
0>
0C
#591890000000
1!
1*
b10 6
19
1>
1C
b10 G
#591900000000
0!
0*
09
0>
0C
#591910000000
1!
1*
b11 6
19
1>
1C
b11 G
#591920000000
0!
0*
09
0>
0C
#591930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#591940000000
0!
0*
09
0>
0C
#591950000000
1!
1*
b101 6
19
1>
1C
b101 G
#591960000000
0!
0*
09
0>
0C
#591970000000
1!
1*
b110 6
19
1>
1C
b110 G
#591980000000
0!
0*
09
0>
0C
#591990000000
1!
1*
b111 6
19
1>
1C
b111 G
#592000000000
0!
0*
09
0>
0C
#592010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#592020000000
0!
0*
09
0>
0C
#592030000000
1!
1*
b1 6
19
1>
1C
b1 G
#592040000000
0!
0*
09
0>
0C
#592050000000
1!
1*
b10 6
19
1>
1C
b10 G
#592060000000
0!
0*
09
0>
0C
#592070000000
1!
1*
b11 6
19
1>
1C
b11 G
#592080000000
0!
0*
09
0>
0C
#592090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#592100000000
0!
0*
09
0>
0C
#592110000000
1!
1*
b101 6
19
1>
1C
b101 G
#592120000000
0!
0*
09
0>
0C
#592130000000
1!
1*
b110 6
19
1>
1C
b110 G
#592140000000
0!
0*
09
0>
0C
#592150000000
1!
1*
b111 6
19
1>
1C
b111 G
#592160000000
0!
0*
09
0>
0C
#592170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#592180000000
0!
0*
09
0>
0C
#592190000000
1!
1*
b1 6
19
1>
1C
b1 G
#592200000000
0!
0*
09
0>
0C
#592210000000
1!
1*
b10 6
19
1>
1C
b10 G
#592220000000
0!
0*
09
0>
0C
#592230000000
1!
1*
b11 6
19
1>
1C
b11 G
#592240000000
0!
0*
09
0>
0C
#592250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#592260000000
0!
0*
09
0>
0C
#592270000000
1!
1*
b101 6
19
1>
1C
b101 G
#592280000000
0!
0*
09
0>
0C
#592290000000
1!
1*
b110 6
19
1>
1C
b110 G
#592300000000
0!
0*
09
0>
0C
#592310000000
1!
1*
b111 6
19
1>
1C
b111 G
#592320000000
0!
1"
0*
1+
09
1:
0>
0C
#592330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#592340000000
0!
0*
09
0>
0C
#592350000000
1!
1*
b1 6
19
1>
1C
b1 G
#592360000000
0!
0*
09
0>
0C
#592370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#592380000000
0!
0*
09
0>
0C
#592390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#592400000000
0!
0*
09
0>
0C
#592410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#592420000000
0!
0*
09
0>
0C
#592430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#592440000000
0!
0#
0*
0,
09
0>
0?
0C
#592450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#592460000000
0!
0*
09
0>
0C
#592470000000
1!
1*
19
1>
1C
#592480000000
0!
0*
09
0>
0C
#592490000000
1!
1*
19
1>
1C
#592500000000
0!
0*
09
0>
0C
#592510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#592520000000
0!
0*
09
0>
0C
#592530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#592540000000
0!
0*
09
0>
0C
#592550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#592560000000
0!
0*
09
0>
0C
#592570000000
1!
1*
b10 6
19
1>
1C
b10 G
#592580000000
0!
0*
09
0>
0C
#592590000000
1!
1*
b11 6
19
1>
1C
b11 G
#592600000000
0!
0*
09
0>
0C
#592610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#592620000000
0!
0*
09
0>
0C
#592630000000
1!
1*
b101 6
19
1>
1C
b101 G
#592640000000
0!
0*
09
0>
0C
#592650000000
1!
1*
b110 6
19
1>
1C
b110 G
#592660000000
0!
0*
09
0>
0C
#592670000000
1!
1*
b111 6
19
1>
1C
b111 G
#592680000000
0!
0*
09
0>
0C
#592690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#592700000000
0!
0*
09
0>
0C
#592710000000
1!
1*
b1 6
19
1>
1C
b1 G
#592720000000
0!
0*
09
0>
0C
#592730000000
1!
1*
b10 6
19
1>
1C
b10 G
#592740000000
0!
0*
09
0>
0C
#592750000000
1!
1*
b11 6
19
1>
1C
b11 G
#592760000000
0!
0*
09
0>
0C
#592770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#592780000000
0!
0*
09
0>
0C
#592790000000
1!
1*
b101 6
19
1>
1C
b101 G
#592800000000
0!
0*
09
0>
0C
#592810000000
1!
1*
b110 6
19
1>
1C
b110 G
#592820000000
0!
0*
09
0>
0C
#592830000000
1!
1*
b111 6
19
1>
1C
b111 G
#592840000000
0!
0*
09
0>
0C
#592850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#592860000000
0!
0*
09
0>
0C
#592870000000
1!
1*
b1 6
19
1>
1C
b1 G
#592880000000
0!
0*
09
0>
0C
#592890000000
1!
1*
b10 6
19
1>
1C
b10 G
#592900000000
0!
0*
09
0>
0C
#592910000000
1!
1*
b11 6
19
1>
1C
b11 G
#592920000000
0!
0*
09
0>
0C
#592930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#592940000000
0!
0*
09
0>
0C
#592950000000
1!
1*
b101 6
19
1>
1C
b101 G
#592960000000
0!
0*
09
0>
0C
#592970000000
1!
1*
b110 6
19
1>
1C
b110 G
#592980000000
0!
0*
09
0>
0C
#592990000000
1!
1*
b111 6
19
1>
1C
b111 G
#593000000000
0!
1"
0*
1+
09
1:
0>
0C
#593010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#593020000000
0!
0*
09
0>
0C
#593030000000
1!
1*
b1 6
19
1>
1C
b1 G
#593040000000
0!
0*
09
0>
0C
#593050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#593060000000
0!
0*
09
0>
0C
#593070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#593080000000
0!
0*
09
0>
0C
#593090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#593100000000
0!
0*
09
0>
0C
#593110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#593120000000
0!
0#
0*
0,
09
0>
0?
0C
#593130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#593140000000
0!
0*
09
0>
0C
#593150000000
1!
1*
19
1>
1C
#593160000000
0!
0*
09
0>
0C
#593170000000
1!
1*
19
1>
1C
#593180000000
0!
0*
09
0>
0C
#593190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#593200000000
0!
0*
09
0>
0C
#593210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#593220000000
0!
0*
09
0>
0C
#593230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#593240000000
0!
0*
09
0>
0C
#593250000000
1!
1*
b10 6
19
1>
1C
b10 G
#593260000000
0!
0*
09
0>
0C
#593270000000
1!
1*
b11 6
19
1>
1C
b11 G
#593280000000
0!
0*
09
0>
0C
#593290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#593300000000
0!
0*
09
0>
0C
#593310000000
1!
1*
b101 6
19
1>
1C
b101 G
#593320000000
0!
0*
09
0>
0C
#593330000000
1!
1*
b110 6
19
1>
1C
b110 G
#593340000000
0!
0*
09
0>
0C
#593350000000
1!
1*
b111 6
19
1>
1C
b111 G
#593360000000
0!
0*
09
0>
0C
#593370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#593380000000
0!
0*
09
0>
0C
#593390000000
1!
1*
b1 6
19
1>
1C
b1 G
#593400000000
0!
0*
09
0>
0C
#593410000000
1!
1*
b10 6
19
1>
1C
b10 G
#593420000000
0!
0*
09
0>
0C
#593430000000
1!
1*
b11 6
19
1>
1C
b11 G
#593440000000
0!
0*
09
0>
0C
#593450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#593460000000
0!
0*
09
0>
0C
#593470000000
1!
1*
b101 6
19
1>
1C
b101 G
#593480000000
0!
0*
09
0>
0C
#593490000000
1!
1*
b110 6
19
1>
1C
b110 G
#593500000000
0!
0*
09
0>
0C
#593510000000
1!
1*
b111 6
19
1>
1C
b111 G
#593520000000
0!
0*
09
0>
0C
#593530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#593540000000
0!
0*
09
0>
0C
#593550000000
1!
1*
b1 6
19
1>
1C
b1 G
#593560000000
0!
0*
09
0>
0C
#593570000000
1!
1*
b10 6
19
1>
1C
b10 G
#593580000000
0!
0*
09
0>
0C
#593590000000
1!
1*
b11 6
19
1>
1C
b11 G
#593600000000
0!
0*
09
0>
0C
#593610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#593620000000
0!
0*
09
0>
0C
#593630000000
1!
1*
b101 6
19
1>
1C
b101 G
#593640000000
0!
0*
09
0>
0C
#593650000000
1!
1*
b110 6
19
1>
1C
b110 G
#593660000000
0!
0*
09
0>
0C
#593670000000
1!
1*
b111 6
19
1>
1C
b111 G
#593680000000
0!
1"
0*
1+
09
1:
0>
0C
#593690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#593700000000
0!
0*
09
0>
0C
#593710000000
1!
1*
b1 6
19
1>
1C
b1 G
#593720000000
0!
0*
09
0>
0C
#593730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#593740000000
0!
0*
09
0>
0C
#593750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#593760000000
0!
0*
09
0>
0C
#593770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#593780000000
0!
0*
09
0>
0C
#593790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#593800000000
0!
0#
0*
0,
09
0>
0?
0C
#593810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#593820000000
0!
0*
09
0>
0C
#593830000000
1!
1*
19
1>
1C
#593840000000
0!
0*
09
0>
0C
#593850000000
1!
1*
19
1>
1C
#593860000000
0!
0*
09
0>
0C
#593870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#593880000000
0!
0*
09
0>
0C
#593890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#593900000000
0!
0*
09
0>
0C
#593910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#593920000000
0!
0*
09
0>
0C
#593930000000
1!
1*
b10 6
19
1>
1C
b10 G
#593940000000
0!
0*
09
0>
0C
#593950000000
1!
1*
b11 6
19
1>
1C
b11 G
#593960000000
0!
0*
09
0>
0C
#593970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#593980000000
0!
0*
09
0>
0C
#593990000000
1!
1*
b101 6
19
1>
1C
b101 G
#594000000000
0!
0*
09
0>
0C
#594010000000
1!
1*
b110 6
19
1>
1C
b110 G
#594020000000
0!
0*
09
0>
0C
#594030000000
1!
1*
b111 6
19
1>
1C
b111 G
#594040000000
0!
0*
09
0>
0C
#594050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#594060000000
0!
0*
09
0>
0C
#594070000000
1!
1*
b1 6
19
1>
1C
b1 G
#594080000000
0!
0*
09
0>
0C
#594090000000
1!
1*
b10 6
19
1>
1C
b10 G
#594100000000
0!
0*
09
0>
0C
#594110000000
1!
1*
b11 6
19
1>
1C
b11 G
#594120000000
0!
0*
09
0>
0C
#594130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#594140000000
0!
0*
09
0>
0C
#594150000000
1!
1*
b101 6
19
1>
1C
b101 G
#594160000000
0!
0*
09
0>
0C
#594170000000
1!
1*
b110 6
19
1>
1C
b110 G
#594180000000
0!
0*
09
0>
0C
#594190000000
1!
1*
b111 6
19
1>
1C
b111 G
#594200000000
0!
0*
09
0>
0C
#594210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#594220000000
0!
0*
09
0>
0C
#594230000000
1!
1*
b1 6
19
1>
1C
b1 G
#594240000000
0!
0*
09
0>
0C
#594250000000
1!
1*
b10 6
19
1>
1C
b10 G
#594260000000
0!
0*
09
0>
0C
#594270000000
1!
1*
b11 6
19
1>
1C
b11 G
#594280000000
0!
0*
09
0>
0C
#594290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#594300000000
0!
0*
09
0>
0C
#594310000000
1!
1*
b101 6
19
1>
1C
b101 G
#594320000000
0!
0*
09
0>
0C
#594330000000
1!
1*
b110 6
19
1>
1C
b110 G
#594340000000
0!
0*
09
0>
0C
#594350000000
1!
1*
b111 6
19
1>
1C
b111 G
#594360000000
0!
1"
0*
1+
09
1:
0>
0C
#594370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#594380000000
0!
0*
09
0>
0C
#594390000000
1!
1*
b1 6
19
1>
1C
b1 G
#594400000000
0!
0*
09
0>
0C
#594410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#594420000000
0!
0*
09
0>
0C
#594430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#594440000000
0!
0*
09
0>
0C
#594450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#594460000000
0!
0*
09
0>
0C
#594470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#594480000000
0!
0#
0*
0,
09
0>
0?
0C
#594490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#594500000000
0!
0*
09
0>
0C
#594510000000
1!
1*
19
1>
1C
#594520000000
0!
0*
09
0>
0C
#594530000000
1!
1*
19
1>
1C
#594540000000
0!
0*
09
0>
0C
#594550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#594560000000
0!
0*
09
0>
0C
#594570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#594580000000
0!
0*
09
0>
0C
#594590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#594600000000
0!
0*
09
0>
0C
#594610000000
1!
1*
b10 6
19
1>
1C
b10 G
#594620000000
0!
0*
09
0>
0C
#594630000000
1!
1*
b11 6
19
1>
1C
b11 G
#594640000000
0!
0*
09
0>
0C
#594650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#594660000000
0!
0*
09
0>
0C
#594670000000
1!
1*
b101 6
19
1>
1C
b101 G
#594680000000
0!
0*
09
0>
0C
#594690000000
1!
1*
b110 6
19
1>
1C
b110 G
#594700000000
0!
0*
09
0>
0C
#594710000000
1!
1*
b111 6
19
1>
1C
b111 G
#594720000000
0!
0*
09
0>
0C
#594730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#594740000000
0!
0*
09
0>
0C
#594750000000
1!
1*
b1 6
19
1>
1C
b1 G
#594760000000
0!
0*
09
0>
0C
#594770000000
1!
1*
b10 6
19
1>
1C
b10 G
#594780000000
0!
0*
09
0>
0C
#594790000000
1!
1*
b11 6
19
1>
1C
b11 G
#594800000000
0!
0*
09
0>
0C
#594810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#594820000000
0!
0*
09
0>
0C
#594830000000
1!
1*
b101 6
19
1>
1C
b101 G
#594840000000
0!
0*
09
0>
0C
#594850000000
1!
1*
b110 6
19
1>
1C
b110 G
#594860000000
0!
0*
09
0>
0C
#594870000000
1!
1*
b111 6
19
1>
1C
b111 G
#594880000000
0!
0*
09
0>
0C
#594890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#594900000000
0!
0*
09
0>
0C
#594910000000
1!
1*
b1 6
19
1>
1C
b1 G
#594920000000
0!
0*
09
0>
0C
#594930000000
1!
1*
b10 6
19
1>
1C
b10 G
#594940000000
0!
0*
09
0>
0C
#594950000000
1!
1*
b11 6
19
1>
1C
b11 G
#594960000000
0!
0*
09
0>
0C
#594970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#594980000000
0!
0*
09
0>
0C
#594990000000
1!
1*
b101 6
19
1>
1C
b101 G
#595000000000
0!
0*
09
0>
0C
#595010000000
1!
1*
b110 6
19
1>
1C
b110 G
#595020000000
0!
0*
09
0>
0C
#595030000000
1!
1*
b111 6
19
1>
1C
b111 G
#595040000000
0!
1"
0*
1+
09
1:
0>
0C
#595050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#595060000000
0!
0*
09
0>
0C
#595070000000
1!
1*
b1 6
19
1>
1C
b1 G
#595080000000
0!
0*
09
0>
0C
#595090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#595100000000
0!
0*
09
0>
0C
#595110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#595120000000
0!
0*
09
0>
0C
#595130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#595140000000
0!
0*
09
0>
0C
#595150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#595160000000
0!
0#
0*
0,
09
0>
0?
0C
#595170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#595180000000
0!
0*
09
0>
0C
#595190000000
1!
1*
19
1>
1C
#595200000000
0!
0*
09
0>
0C
#595210000000
1!
1*
19
1>
1C
#595220000000
0!
0*
09
0>
0C
#595230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#595240000000
0!
0*
09
0>
0C
#595250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#595260000000
0!
0*
09
0>
0C
#595270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#595280000000
0!
0*
09
0>
0C
#595290000000
1!
1*
b10 6
19
1>
1C
b10 G
#595300000000
0!
0*
09
0>
0C
#595310000000
1!
1*
b11 6
19
1>
1C
b11 G
#595320000000
0!
0*
09
0>
0C
#595330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#595340000000
0!
0*
09
0>
0C
#595350000000
1!
1*
b101 6
19
1>
1C
b101 G
#595360000000
0!
0*
09
0>
0C
#595370000000
1!
1*
b110 6
19
1>
1C
b110 G
#595380000000
0!
0*
09
0>
0C
#595390000000
1!
1*
b111 6
19
1>
1C
b111 G
#595400000000
0!
0*
09
0>
0C
#595410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#595420000000
0!
0*
09
0>
0C
#595430000000
1!
1*
b1 6
19
1>
1C
b1 G
#595440000000
0!
0*
09
0>
0C
#595450000000
1!
1*
b10 6
19
1>
1C
b10 G
#595460000000
0!
0*
09
0>
0C
#595470000000
1!
1*
b11 6
19
1>
1C
b11 G
#595480000000
0!
0*
09
0>
0C
#595490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#595500000000
0!
0*
09
0>
0C
#595510000000
1!
1*
b101 6
19
1>
1C
b101 G
#595520000000
0!
0*
09
0>
0C
#595530000000
1!
1*
b110 6
19
1>
1C
b110 G
#595540000000
0!
0*
09
0>
0C
#595550000000
1!
1*
b111 6
19
1>
1C
b111 G
#595560000000
0!
0*
09
0>
0C
#595570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#595580000000
0!
0*
09
0>
0C
#595590000000
1!
1*
b1 6
19
1>
1C
b1 G
#595600000000
0!
0*
09
0>
0C
#595610000000
1!
1*
b10 6
19
1>
1C
b10 G
#595620000000
0!
0*
09
0>
0C
#595630000000
1!
1*
b11 6
19
1>
1C
b11 G
#595640000000
0!
0*
09
0>
0C
#595650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#595660000000
0!
0*
09
0>
0C
#595670000000
1!
1*
b101 6
19
1>
1C
b101 G
#595680000000
0!
0*
09
0>
0C
#595690000000
1!
1*
b110 6
19
1>
1C
b110 G
#595700000000
0!
0*
09
0>
0C
#595710000000
1!
1*
b111 6
19
1>
1C
b111 G
#595720000000
0!
1"
0*
1+
09
1:
0>
0C
#595730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#595740000000
0!
0*
09
0>
0C
#595750000000
1!
1*
b1 6
19
1>
1C
b1 G
#595760000000
0!
0*
09
0>
0C
#595770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#595780000000
0!
0*
09
0>
0C
#595790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#595800000000
0!
0*
09
0>
0C
#595810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#595820000000
0!
0*
09
0>
0C
#595830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#595840000000
0!
0#
0*
0,
09
0>
0?
0C
#595850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#595860000000
0!
0*
09
0>
0C
#595870000000
1!
1*
19
1>
1C
#595880000000
0!
0*
09
0>
0C
#595890000000
1!
1*
19
1>
1C
#595900000000
0!
0*
09
0>
0C
#595910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#595920000000
0!
0*
09
0>
0C
#595930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#595940000000
0!
0*
09
0>
0C
#595950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#595960000000
0!
0*
09
0>
0C
#595970000000
1!
1*
b10 6
19
1>
1C
b10 G
#595980000000
0!
0*
09
0>
0C
#595990000000
1!
1*
b11 6
19
1>
1C
b11 G
#596000000000
0!
0*
09
0>
0C
#596010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#596020000000
0!
0*
09
0>
0C
#596030000000
1!
1*
b101 6
19
1>
1C
b101 G
#596040000000
0!
0*
09
0>
0C
#596050000000
1!
1*
b110 6
19
1>
1C
b110 G
#596060000000
0!
0*
09
0>
0C
#596070000000
1!
1*
b111 6
19
1>
1C
b111 G
#596080000000
0!
0*
09
0>
0C
#596090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#596100000000
0!
0*
09
0>
0C
#596110000000
1!
1*
b1 6
19
1>
1C
b1 G
#596120000000
0!
0*
09
0>
0C
#596130000000
1!
1*
b10 6
19
1>
1C
b10 G
#596140000000
0!
0*
09
0>
0C
#596150000000
1!
1*
b11 6
19
1>
1C
b11 G
#596160000000
0!
0*
09
0>
0C
#596170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#596180000000
0!
0*
09
0>
0C
#596190000000
1!
1*
b101 6
19
1>
1C
b101 G
#596200000000
0!
0*
09
0>
0C
#596210000000
1!
1*
b110 6
19
1>
1C
b110 G
#596220000000
0!
0*
09
0>
0C
#596230000000
1!
1*
b111 6
19
1>
1C
b111 G
#596240000000
0!
0*
09
0>
0C
#596250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#596260000000
0!
0*
09
0>
0C
#596270000000
1!
1*
b1 6
19
1>
1C
b1 G
#596280000000
0!
0*
09
0>
0C
#596290000000
1!
1*
b10 6
19
1>
1C
b10 G
#596300000000
0!
0*
09
0>
0C
#596310000000
1!
1*
b11 6
19
1>
1C
b11 G
#596320000000
0!
0*
09
0>
0C
#596330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#596340000000
0!
0*
09
0>
0C
#596350000000
1!
1*
b101 6
19
1>
1C
b101 G
#596360000000
0!
0*
09
0>
0C
#596370000000
1!
1*
b110 6
19
1>
1C
b110 G
#596380000000
0!
0*
09
0>
0C
#596390000000
1!
1*
b111 6
19
1>
1C
b111 G
#596400000000
0!
1"
0*
1+
09
1:
0>
0C
#596410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#596420000000
0!
0*
09
0>
0C
#596430000000
1!
1*
b1 6
19
1>
1C
b1 G
#596440000000
0!
0*
09
0>
0C
#596450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#596460000000
0!
0*
09
0>
0C
#596470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#596480000000
0!
0*
09
0>
0C
#596490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#596500000000
0!
0*
09
0>
0C
#596510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#596520000000
0!
0#
0*
0,
09
0>
0?
0C
#596530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#596540000000
0!
0*
09
0>
0C
#596550000000
1!
1*
19
1>
1C
#596560000000
0!
0*
09
0>
0C
#596570000000
1!
1*
19
1>
1C
#596580000000
0!
0*
09
0>
0C
#596590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#596600000000
0!
0*
09
0>
0C
#596610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#596620000000
0!
0*
09
0>
0C
#596630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#596640000000
0!
0*
09
0>
0C
#596650000000
1!
1*
b10 6
19
1>
1C
b10 G
#596660000000
0!
0*
09
0>
0C
#596670000000
1!
1*
b11 6
19
1>
1C
b11 G
#596680000000
0!
0*
09
0>
0C
#596690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#596700000000
0!
0*
09
0>
0C
#596710000000
1!
1*
b101 6
19
1>
1C
b101 G
#596720000000
0!
0*
09
0>
0C
#596730000000
1!
1*
b110 6
19
1>
1C
b110 G
#596740000000
0!
0*
09
0>
0C
#596750000000
1!
1*
b111 6
19
1>
1C
b111 G
#596760000000
0!
0*
09
0>
0C
#596770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#596780000000
0!
0*
09
0>
0C
#596790000000
1!
1*
b1 6
19
1>
1C
b1 G
#596800000000
0!
0*
09
0>
0C
#596810000000
1!
1*
b10 6
19
1>
1C
b10 G
#596820000000
0!
0*
09
0>
0C
#596830000000
1!
1*
b11 6
19
1>
1C
b11 G
#596840000000
0!
0*
09
0>
0C
#596850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#596860000000
0!
0*
09
0>
0C
#596870000000
1!
1*
b101 6
19
1>
1C
b101 G
#596880000000
0!
0*
09
0>
0C
#596890000000
1!
1*
b110 6
19
1>
1C
b110 G
#596900000000
0!
0*
09
0>
0C
#596910000000
1!
1*
b111 6
19
1>
1C
b111 G
#596920000000
0!
0*
09
0>
0C
#596930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#596940000000
0!
0*
09
0>
0C
#596950000000
1!
1*
b1 6
19
1>
1C
b1 G
#596960000000
0!
0*
09
0>
0C
#596970000000
1!
1*
b10 6
19
1>
1C
b10 G
#596980000000
0!
0*
09
0>
0C
#596990000000
1!
1*
b11 6
19
1>
1C
b11 G
#597000000000
0!
0*
09
0>
0C
#597010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#597020000000
0!
0*
09
0>
0C
#597030000000
1!
1*
b101 6
19
1>
1C
b101 G
#597040000000
0!
0*
09
0>
0C
#597050000000
1!
1*
b110 6
19
1>
1C
b110 G
#597060000000
0!
0*
09
0>
0C
#597070000000
1!
1*
b111 6
19
1>
1C
b111 G
#597080000000
0!
1"
0*
1+
09
1:
0>
0C
#597090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#597100000000
0!
0*
09
0>
0C
#597110000000
1!
1*
b1 6
19
1>
1C
b1 G
#597120000000
0!
0*
09
0>
0C
#597130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#597140000000
0!
0*
09
0>
0C
#597150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#597160000000
0!
0*
09
0>
0C
#597170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#597180000000
0!
0*
09
0>
0C
#597190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#597200000000
0!
0#
0*
0,
09
0>
0?
0C
#597210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#597220000000
0!
0*
09
0>
0C
#597230000000
1!
1*
19
1>
1C
#597240000000
0!
0*
09
0>
0C
#597250000000
1!
1*
19
1>
1C
#597260000000
0!
0*
09
0>
0C
#597270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#597280000000
0!
0*
09
0>
0C
#597290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#597300000000
0!
0*
09
0>
0C
#597310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#597320000000
0!
0*
09
0>
0C
#597330000000
1!
1*
b10 6
19
1>
1C
b10 G
#597340000000
0!
0*
09
0>
0C
#597350000000
1!
1*
b11 6
19
1>
1C
b11 G
#597360000000
0!
0*
09
0>
0C
#597370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#597380000000
0!
0*
09
0>
0C
#597390000000
1!
1*
b101 6
19
1>
1C
b101 G
#597400000000
0!
0*
09
0>
0C
#597410000000
1!
1*
b110 6
19
1>
1C
b110 G
#597420000000
0!
0*
09
0>
0C
#597430000000
1!
1*
b111 6
19
1>
1C
b111 G
#597440000000
0!
0*
09
0>
0C
#597450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#597460000000
0!
0*
09
0>
0C
#597470000000
1!
1*
b1 6
19
1>
1C
b1 G
#597480000000
0!
0*
09
0>
0C
#597490000000
1!
1*
b10 6
19
1>
1C
b10 G
#597500000000
0!
0*
09
0>
0C
#597510000000
1!
1*
b11 6
19
1>
1C
b11 G
#597520000000
0!
0*
09
0>
0C
#597530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#597540000000
0!
0*
09
0>
0C
#597550000000
1!
1*
b101 6
19
1>
1C
b101 G
#597560000000
0!
0*
09
0>
0C
#597570000000
1!
1*
b110 6
19
1>
1C
b110 G
#597580000000
0!
0*
09
0>
0C
#597590000000
1!
1*
b111 6
19
1>
1C
b111 G
#597600000000
0!
0*
09
0>
0C
#597610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#597620000000
0!
0*
09
0>
0C
#597630000000
1!
1*
b1 6
19
1>
1C
b1 G
#597640000000
0!
0*
09
0>
0C
#597650000000
1!
1*
b10 6
19
1>
1C
b10 G
#597660000000
0!
0*
09
0>
0C
#597670000000
1!
1*
b11 6
19
1>
1C
b11 G
#597680000000
0!
0*
09
0>
0C
#597690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#597700000000
0!
0*
09
0>
0C
#597710000000
1!
1*
b101 6
19
1>
1C
b101 G
#597720000000
0!
0*
09
0>
0C
#597730000000
1!
1*
b110 6
19
1>
1C
b110 G
#597740000000
0!
0*
09
0>
0C
#597750000000
1!
1*
b111 6
19
1>
1C
b111 G
#597760000000
0!
1"
0*
1+
09
1:
0>
0C
#597770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#597780000000
0!
0*
09
0>
0C
#597790000000
1!
1*
b1 6
19
1>
1C
b1 G
#597800000000
0!
0*
09
0>
0C
#597810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#597820000000
0!
0*
09
0>
0C
#597830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#597840000000
0!
0*
09
0>
0C
#597850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#597860000000
0!
0*
09
0>
0C
#597870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#597880000000
0!
0#
0*
0,
09
0>
0?
0C
#597890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#597900000000
0!
0*
09
0>
0C
#597910000000
1!
1*
19
1>
1C
#597920000000
0!
0*
09
0>
0C
#597930000000
1!
1*
19
1>
1C
#597940000000
0!
0*
09
0>
0C
#597950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#597960000000
0!
0*
09
0>
0C
#597970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#597980000000
0!
0*
09
0>
0C
#597990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#598000000000
0!
0*
09
0>
0C
#598010000000
1!
1*
b10 6
19
1>
1C
b10 G
#598020000000
0!
0*
09
0>
0C
#598030000000
1!
1*
b11 6
19
1>
1C
b11 G
#598040000000
0!
0*
09
0>
0C
#598050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#598060000000
0!
0*
09
0>
0C
#598070000000
1!
1*
b101 6
19
1>
1C
b101 G
#598080000000
0!
0*
09
0>
0C
#598090000000
1!
1*
b110 6
19
1>
1C
b110 G
#598100000000
0!
0*
09
0>
0C
#598110000000
1!
1*
b111 6
19
1>
1C
b111 G
#598120000000
0!
0*
09
0>
0C
#598130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#598140000000
0!
0*
09
0>
0C
#598150000000
1!
1*
b1 6
19
1>
1C
b1 G
#598160000000
0!
0*
09
0>
0C
#598170000000
1!
1*
b10 6
19
1>
1C
b10 G
#598180000000
0!
0*
09
0>
0C
#598190000000
1!
1*
b11 6
19
1>
1C
b11 G
#598200000000
0!
0*
09
0>
0C
#598210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#598220000000
0!
0*
09
0>
0C
#598230000000
1!
1*
b101 6
19
1>
1C
b101 G
#598240000000
0!
0*
09
0>
0C
#598250000000
1!
1*
b110 6
19
1>
1C
b110 G
#598260000000
0!
0*
09
0>
0C
#598270000000
1!
1*
b111 6
19
1>
1C
b111 G
#598280000000
0!
0*
09
0>
0C
#598290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#598300000000
0!
0*
09
0>
0C
#598310000000
1!
1*
b1 6
19
1>
1C
b1 G
#598320000000
0!
0*
09
0>
0C
#598330000000
1!
1*
b10 6
19
1>
1C
b10 G
#598340000000
0!
0*
09
0>
0C
#598350000000
1!
1*
b11 6
19
1>
1C
b11 G
#598360000000
0!
0*
09
0>
0C
#598370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#598380000000
0!
0*
09
0>
0C
#598390000000
1!
1*
b101 6
19
1>
1C
b101 G
#598400000000
0!
0*
09
0>
0C
#598410000000
1!
1*
b110 6
19
1>
1C
b110 G
#598420000000
0!
0*
09
0>
0C
#598430000000
1!
1*
b111 6
19
1>
1C
b111 G
#598440000000
0!
1"
0*
1+
09
1:
0>
0C
#598450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#598460000000
0!
0*
09
0>
0C
#598470000000
1!
1*
b1 6
19
1>
1C
b1 G
#598480000000
0!
0*
09
0>
0C
#598490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#598500000000
0!
0*
09
0>
0C
#598510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#598520000000
0!
0*
09
0>
0C
#598530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#598540000000
0!
0*
09
0>
0C
#598550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#598560000000
0!
0#
0*
0,
09
0>
0?
0C
#598570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#598580000000
0!
0*
09
0>
0C
#598590000000
1!
1*
19
1>
1C
#598600000000
0!
0*
09
0>
0C
#598610000000
1!
1*
19
1>
1C
#598620000000
0!
0*
09
0>
0C
#598630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#598640000000
0!
0*
09
0>
0C
#598650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#598660000000
0!
0*
09
0>
0C
#598670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#598680000000
0!
0*
09
0>
0C
#598690000000
1!
1*
b10 6
19
1>
1C
b10 G
#598700000000
0!
0*
09
0>
0C
#598710000000
1!
1*
b11 6
19
1>
1C
b11 G
#598720000000
0!
0*
09
0>
0C
#598730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#598740000000
0!
0*
09
0>
0C
#598750000000
1!
1*
b101 6
19
1>
1C
b101 G
#598760000000
0!
0*
09
0>
0C
#598770000000
1!
1*
b110 6
19
1>
1C
b110 G
#598780000000
0!
0*
09
0>
0C
#598790000000
1!
1*
b111 6
19
1>
1C
b111 G
#598800000000
0!
0*
09
0>
0C
#598810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#598820000000
0!
0*
09
0>
0C
#598830000000
1!
1*
b1 6
19
1>
1C
b1 G
#598840000000
0!
0*
09
0>
0C
#598850000000
1!
1*
b10 6
19
1>
1C
b10 G
#598860000000
0!
0*
09
0>
0C
#598870000000
1!
1*
b11 6
19
1>
1C
b11 G
#598880000000
0!
0*
09
0>
0C
#598890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#598900000000
0!
0*
09
0>
0C
#598910000000
1!
1*
b101 6
19
1>
1C
b101 G
#598920000000
0!
0*
09
0>
0C
#598930000000
1!
1*
b110 6
19
1>
1C
b110 G
#598940000000
0!
0*
09
0>
0C
#598950000000
1!
1*
b111 6
19
1>
1C
b111 G
#598960000000
0!
0*
09
0>
0C
#598970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#598980000000
0!
0*
09
0>
0C
#598990000000
1!
1*
b1 6
19
1>
1C
b1 G
#599000000000
0!
0*
09
0>
0C
#599010000000
1!
1*
b10 6
19
1>
1C
b10 G
#599020000000
0!
0*
09
0>
0C
#599030000000
1!
1*
b11 6
19
1>
1C
b11 G
#599040000000
0!
0*
09
0>
0C
#599050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#599060000000
0!
0*
09
0>
0C
#599070000000
1!
1*
b101 6
19
1>
1C
b101 G
#599080000000
0!
0*
09
0>
0C
#599090000000
1!
1*
b110 6
19
1>
1C
b110 G
#599100000000
0!
0*
09
0>
0C
#599110000000
1!
1*
b111 6
19
1>
1C
b111 G
#599120000000
0!
1"
0*
1+
09
1:
0>
0C
#599130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#599140000000
0!
0*
09
0>
0C
#599150000000
1!
1*
b1 6
19
1>
1C
b1 G
#599160000000
0!
0*
09
0>
0C
#599170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#599180000000
0!
0*
09
0>
0C
#599190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#599200000000
0!
0*
09
0>
0C
#599210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#599220000000
0!
0*
09
0>
0C
#599230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#599240000000
0!
0#
0*
0,
09
0>
0?
0C
#599250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#599260000000
0!
0*
09
0>
0C
#599270000000
1!
1*
19
1>
1C
#599280000000
0!
0*
09
0>
0C
#599290000000
1!
1*
19
1>
1C
#599300000000
0!
0*
09
0>
0C
#599310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#599320000000
0!
0*
09
0>
0C
#599330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#599340000000
0!
0*
09
0>
0C
#599350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#599360000000
0!
0*
09
0>
0C
#599370000000
1!
1*
b10 6
19
1>
1C
b10 G
#599380000000
0!
0*
09
0>
0C
#599390000000
1!
1*
b11 6
19
1>
1C
b11 G
#599400000000
0!
0*
09
0>
0C
#599410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#599420000000
0!
0*
09
0>
0C
#599430000000
1!
1*
b101 6
19
1>
1C
b101 G
#599440000000
0!
0*
09
0>
0C
#599450000000
1!
1*
b110 6
19
1>
1C
b110 G
#599460000000
0!
0*
09
0>
0C
#599470000000
1!
1*
b111 6
19
1>
1C
b111 G
#599480000000
0!
0*
09
0>
0C
#599490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#599500000000
0!
0*
09
0>
0C
#599510000000
1!
1*
b1 6
19
1>
1C
b1 G
#599520000000
0!
0*
09
0>
0C
#599530000000
1!
1*
b10 6
19
1>
1C
b10 G
#599540000000
0!
0*
09
0>
0C
#599550000000
1!
1*
b11 6
19
1>
1C
b11 G
#599560000000
0!
0*
09
0>
0C
#599570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#599580000000
0!
0*
09
0>
0C
#599590000000
1!
1*
b101 6
19
1>
1C
b101 G
#599600000000
0!
0*
09
0>
0C
#599610000000
1!
1*
b110 6
19
1>
1C
b110 G
#599620000000
0!
0*
09
0>
0C
#599630000000
1!
1*
b111 6
19
1>
1C
b111 G
#599640000000
0!
0*
09
0>
0C
#599650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#599660000000
0!
0*
09
0>
0C
#599670000000
1!
1*
b1 6
19
1>
1C
b1 G
#599680000000
0!
0*
09
0>
0C
#599690000000
1!
1*
b10 6
19
1>
1C
b10 G
#599700000000
0!
0*
09
0>
0C
#599710000000
1!
1*
b11 6
19
1>
1C
b11 G
#599720000000
0!
0*
09
0>
0C
#599730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#599740000000
0!
0*
09
0>
0C
#599750000000
1!
1*
b101 6
19
1>
1C
b101 G
#599760000000
0!
0*
09
0>
0C
#599770000000
1!
1*
b110 6
19
1>
1C
b110 G
#599780000000
0!
0*
09
0>
0C
#599790000000
1!
1*
b111 6
19
1>
1C
b111 G
#599800000000
0!
1"
0*
1+
09
1:
0>
0C
#599810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#599820000000
0!
0*
09
0>
0C
#599830000000
1!
1*
b1 6
19
1>
1C
b1 G
#599840000000
0!
0*
09
0>
0C
#599850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#599860000000
0!
0*
09
0>
0C
#599870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#599880000000
0!
0*
09
0>
0C
#599890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#599900000000
0!
0*
09
0>
0C
#599910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#599920000000
0!
0#
0*
0,
09
0>
0?
0C
#599930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#599940000000
0!
0*
09
0>
0C
#599950000000
1!
1*
19
1>
1C
#599960000000
0!
0*
09
0>
0C
#599970000000
1!
1*
19
1>
1C
#599980000000
0!
0*
09
0>
0C
#599990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#600000000000
0!
0*
09
0>
0C
#600010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#600020000000
0!
0*
09
0>
0C
#600030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#600040000000
0!
0*
09
0>
0C
#600050000000
1!
1*
b10 6
19
1>
1C
b10 G
#600060000000
0!
0*
09
0>
0C
#600070000000
1!
1*
b11 6
19
1>
1C
b11 G
#600080000000
0!
0*
09
0>
0C
#600090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#600100000000
0!
0*
09
0>
0C
#600110000000
1!
1*
b101 6
19
1>
1C
b101 G
#600120000000
0!
0*
09
0>
0C
#600130000000
1!
1*
b110 6
19
1>
1C
b110 G
#600140000000
0!
0*
09
0>
0C
#600150000000
1!
1*
b111 6
19
1>
1C
b111 G
#600160000000
0!
0*
09
0>
0C
#600170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#600180000000
0!
0*
09
0>
0C
#600190000000
1!
1*
b1 6
19
1>
1C
b1 G
#600200000000
0!
0*
09
0>
0C
#600210000000
1!
1*
b10 6
19
1>
1C
b10 G
#600220000000
0!
0*
09
0>
0C
#600230000000
1!
1*
b11 6
19
1>
1C
b11 G
#600240000000
0!
0*
09
0>
0C
#600250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#600260000000
0!
0*
09
0>
0C
#600270000000
1!
1*
b101 6
19
1>
1C
b101 G
#600280000000
0!
0*
09
0>
0C
#600290000000
1!
1*
b110 6
19
1>
1C
b110 G
#600300000000
0!
0*
09
0>
0C
#600310000000
1!
1*
b111 6
19
1>
1C
b111 G
#600320000000
0!
0*
09
0>
0C
#600330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#600340000000
0!
0*
09
0>
0C
#600350000000
1!
1*
b1 6
19
1>
1C
b1 G
#600360000000
0!
0*
09
0>
0C
#600370000000
1!
1*
b10 6
19
1>
1C
b10 G
#600380000000
0!
0*
09
0>
0C
#600390000000
1!
1*
b11 6
19
1>
1C
b11 G
#600400000000
0!
0*
09
0>
0C
#600410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#600420000000
0!
0*
09
0>
0C
#600430000000
1!
1*
b101 6
19
1>
1C
b101 G
#600440000000
0!
0*
09
0>
0C
#600450000000
1!
1*
b110 6
19
1>
1C
b110 G
#600460000000
0!
0*
09
0>
0C
#600470000000
1!
1*
b111 6
19
1>
1C
b111 G
#600480000000
0!
1"
0*
1+
09
1:
0>
0C
#600490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#600500000000
0!
0*
09
0>
0C
#600510000000
1!
1*
b1 6
19
1>
1C
b1 G
#600520000000
0!
0*
09
0>
0C
#600530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#600540000000
0!
0*
09
0>
0C
#600550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#600560000000
0!
0*
09
0>
0C
#600570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#600580000000
0!
0*
09
0>
0C
#600590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#600600000000
0!
0#
0*
0,
09
0>
0?
0C
#600610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#600620000000
0!
0*
09
0>
0C
#600630000000
1!
1*
19
1>
1C
#600640000000
0!
0*
09
0>
0C
#600650000000
1!
1*
19
1>
1C
#600660000000
0!
0*
09
0>
0C
#600670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#600680000000
0!
0*
09
0>
0C
#600690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#600700000000
0!
0*
09
0>
0C
#600710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#600720000000
0!
0*
09
0>
0C
#600730000000
1!
1*
b10 6
19
1>
1C
b10 G
#600740000000
0!
0*
09
0>
0C
#600750000000
1!
1*
b11 6
19
1>
1C
b11 G
#600760000000
0!
0*
09
0>
0C
#600770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#600780000000
0!
0*
09
0>
0C
#600790000000
1!
1*
b101 6
19
1>
1C
b101 G
#600800000000
0!
0*
09
0>
0C
#600810000000
1!
1*
b110 6
19
1>
1C
b110 G
#600820000000
0!
0*
09
0>
0C
#600830000000
1!
1*
b111 6
19
1>
1C
b111 G
#600840000000
0!
0*
09
0>
0C
#600850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#600860000000
0!
0*
09
0>
0C
#600870000000
1!
1*
b1 6
19
1>
1C
b1 G
#600880000000
0!
0*
09
0>
0C
#600890000000
1!
1*
b10 6
19
1>
1C
b10 G
#600900000000
0!
0*
09
0>
0C
#600910000000
1!
1*
b11 6
19
1>
1C
b11 G
#600920000000
0!
0*
09
0>
0C
#600930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#600940000000
0!
0*
09
0>
0C
#600950000000
1!
1*
b101 6
19
1>
1C
b101 G
#600960000000
0!
0*
09
0>
0C
#600970000000
1!
1*
b110 6
19
1>
1C
b110 G
#600980000000
0!
0*
09
0>
0C
#600990000000
1!
1*
b111 6
19
1>
1C
b111 G
#601000000000
0!
0*
09
0>
0C
#601010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#601020000000
0!
0*
09
0>
0C
#601030000000
1!
1*
b1 6
19
1>
1C
b1 G
#601040000000
0!
0*
09
0>
0C
#601050000000
1!
1*
b10 6
19
1>
1C
b10 G
#601060000000
0!
0*
09
0>
0C
#601070000000
1!
1*
b11 6
19
1>
1C
b11 G
#601080000000
0!
0*
09
0>
0C
#601090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#601100000000
0!
0*
09
0>
0C
#601110000000
1!
1*
b101 6
19
1>
1C
b101 G
#601120000000
0!
0*
09
0>
0C
#601130000000
1!
1*
b110 6
19
1>
1C
b110 G
#601140000000
0!
0*
09
0>
0C
#601150000000
1!
1*
b111 6
19
1>
1C
b111 G
#601160000000
0!
1"
0*
1+
09
1:
0>
0C
#601170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#601180000000
0!
0*
09
0>
0C
#601190000000
1!
1*
b1 6
19
1>
1C
b1 G
#601200000000
0!
0*
09
0>
0C
#601210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#601220000000
0!
0*
09
0>
0C
#601230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#601240000000
0!
0*
09
0>
0C
#601250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#601260000000
0!
0*
09
0>
0C
#601270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#601280000000
0!
0#
0*
0,
09
0>
0?
0C
#601290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#601300000000
0!
0*
09
0>
0C
#601310000000
1!
1*
19
1>
1C
#601320000000
0!
0*
09
0>
0C
#601330000000
1!
1*
19
1>
1C
#601340000000
0!
0*
09
0>
0C
#601350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#601360000000
0!
0*
09
0>
0C
#601370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#601380000000
0!
0*
09
0>
0C
#601390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#601400000000
0!
0*
09
0>
0C
#601410000000
1!
1*
b10 6
19
1>
1C
b10 G
#601420000000
0!
0*
09
0>
0C
#601430000000
1!
1*
b11 6
19
1>
1C
b11 G
#601440000000
0!
0*
09
0>
0C
#601450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#601460000000
0!
0*
09
0>
0C
#601470000000
1!
1*
b101 6
19
1>
1C
b101 G
#601480000000
0!
0*
09
0>
0C
#601490000000
1!
1*
b110 6
19
1>
1C
b110 G
#601500000000
0!
0*
09
0>
0C
#601510000000
1!
1*
b111 6
19
1>
1C
b111 G
#601520000000
0!
0*
09
0>
0C
#601530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#601540000000
0!
0*
09
0>
0C
#601550000000
1!
1*
b1 6
19
1>
1C
b1 G
#601560000000
0!
0*
09
0>
0C
#601570000000
1!
1*
b10 6
19
1>
1C
b10 G
#601580000000
0!
0*
09
0>
0C
#601590000000
1!
1*
b11 6
19
1>
1C
b11 G
#601600000000
0!
0*
09
0>
0C
#601610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#601620000000
0!
0*
09
0>
0C
#601630000000
1!
1*
b101 6
19
1>
1C
b101 G
#601640000000
0!
0*
09
0>
0C
#601650000000
1!
1*
b110 6
19
1>
1C
b110 G
#601660000000
0!
0*
09
0>
0C
#601670000000
1!
1*
b111 6
19
1>
1C
b111 G
#601680000000
0!
0*
09
0>
0C
#601690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#601700000000
0!
0*
09
0>
0C
#601710000000
1!
1*
b1 6
19
1>
1C
b1 G
#601720000000
0!
0*
09
0>
0C
#601730000000
1!
1*
b10 6
19
1>
1C
b10 G
#601740000000
0!
0*
09
0>
0C
#601750000000
1!
1*
b11 6
19
1>
1C
b11 G
#601760000000
0!
0*
09
0>
0C
#601770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#601780000000
0!
0*
09
0>
0C
#601790000000
1!
1*
b101 6
19
1>
1C
b101 G
#601800000000
0!
0*
09
0>
0C
#601810000000
1!
1*
b110 6
19
1>
1C
b110 G
#601820000000
0!
0*
09
0>
0C
#601830000000
1!
1*
b111 6
19
1>
1C
b111 G
#601840000000
0!
1"
0*
1+
09
1:
0>
0C
#601850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#601860000000
0!
0*
09
0>
0C
#601870000000
1!
1*
b1 6
19
1>
1C
b1 G
#601880000000
0!
0*
09
0>
0C
#601890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#601900000000
0!
0*
09
0>
0C
#601910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#601920000000
0!
0*
09
0>
0C
#601930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#601940000000
0!
0*
09
0>
0C
#601950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#601960000000
0!
0#
0*
0,
09
0>
0?
0C
#601970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#601980000000
0!
0*
09
0>
0C
#601990000000
1!
1*
19
1>
1C
#602000000000
0!
0*
09
0>
0C
#602010000000
1!
1*
19
1>
1C
#602020000000
0!
0*
09
0>
0C
#602030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#602040000000
0!
0*
09
0>
0C
#602050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#602060000000
0!
0*
09
0>
0C
#602070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#602080000000
0!
0*
09
0>
0C
#602090000000
1!
1*
b10 6
19
1>
1C
b10 G
#602100000000
0!
0*
09
0>
0C
#602110000000
1!
1*
b11 6
19
1>
1C
b11 G
#602120000000
0!
0*
09
0>
0C
#602130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#602140000000
0!
0*
09
0>
0C
#602150000000
1!
1*
b101 6
19
1>
1C
b101 G
#602160000000
0!
0*
09
0>
0C
#602170000000
1!
1*
b110 6
19
1>
1C
b110 G
#602180000000
0!
0*
09
0>
0C
#602190000000
1!
1*
b111 6
19
1>
1C
b111 G
#602200000000
0!
0*
09
0>
0C
#602210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#602220000000
0!
0*
09
0>
0C
#602230000000
1!
1*
b1 6
19
1>
1C
b1 G
#602240000000
0!
0*
09
0>
0C
#602250000000
1!
1*
b10 6
19
1>
1C
b10 G
#602260000000
0!
0*
09
0>
0C
#602270000000
1!
1*
b11 6
19
1>
1C
b11 G
#602280000000
0!
0*
09
0>
0C
#602290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#602300000000
0!
0*
09
0>
0C
#602310000000
1!
1*
b101 6
19
1>
1C
b101 G
#602320000000
0!
0*
09
0>
0C
#602330000000
1!
1*
b110 6
19
1>
1C
b110 G
#602340000000
0!
0*
09
0>
0C
#602350000000
1!
1*
b111 6
19
1>
1C
b111 G
#602360000000
0!
0*
09
0>
0C
#602370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#602380000000
0!
0*
09
0>
0C
#602390000000
1!
1*
b1 6
19
1>
1C
b1 G
#602400000000
0!
0*
09
0>
0C
#602410000000
1!
1*
b10 6
19
1>
1C
b10 G
#602420000000
0!
0*
09
0>
0C
#602430000000
1!
1*
b11 6
19
1>
1C
b11 G
#602440000000
0!
0*
09
0>
0C
#602450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#602460000000
0!
0*
09
0>
0C
#602470000000
1!
1*
b101 6
19
1>
1C
b101 G
#602480000000
0!
0*
09
0>
0C
#602490000000
1!
1*
b110 6
19
1>
1C
b110 G
#602500000000
0!
0*
09
0>
0C
#602510000000
1!
1*
b111 6
19
1>
1C
b111 G
#602520000000
0!
1"
0*
1+
09
1:
0>
0C
#602530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#602540000000
0!
0*
09
0>
0C
#602550000000
1!
1*
b1 6
19
1>
1C
b1 G
#602560000000
0!
0*
09
0>
0C
#602570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#602580000000
0!
0*
09
0>
0C
#602590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#602600000000
0!
0*
09
0>
0C
#602610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#602620000000
0!
0*
09
0>
0C
#602630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#602640000000
0!
0#
0*
0,
09
0>
0?
0C
#602650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#602660000000
0!
0*
09
0>
0C
#602670000000
1!
1*
19
1>
1C
#602680000000
0!
0*
09
0>
0C
#602690000000
1!
1*
19
1>
1C
#602700000000
0!
0*
09
0>
0C
#602710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#602720000000
0!
0*
09
0>
0C
#602730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#602740000000
0!
0*
09
0>
0C
#602750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#602760000000
0!
0*
09
0>
0C
#602770000000
1!
1*
b10 6
19
1>
1C
b10 G
#602780000000
0!
0*
09
0>
0C
#602790000000
1!
1*
b11 6
19
1>
1C
b11 G
#602800000000
0!
0*
09
0>
0C
#602810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#602820000000
0!
0*
09
0>
0C
#602830000000
1!
1*
b101 6
19
1>
1C
b101 G
#602840000000
0!
0*
09
0>
0C
#602850000000
1!
1*
b110 6
19
1>
1C
b110 G
#602860000000
0!
0*
09
0>
0C
#602870000000
1!
1*
b111 6
19
1>
1C
b111 G
#602880000000
0!
0*
09
0>
0C
#602890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#602900000000
0!
0*
09
0>
0C
#602910000000
1!
1*
b1 6
19
1>
1C
b1 G
#602920000000
0!
0*
09
0>
0C
#602930000000
1!
1*
b10 6
19
1>
1C
b10 G
#602940000000
0!
0*
09
0>
0C
#602950000000
1!
1*
b11 6
19
1>
1C
b11 G
#602960000000
0!
0*
09
0>
0C
#602970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#602980000000
0!
0*
09
0>
0C
#602990000000
1!
1*
b101 6
19
1>
1C
b101 G
#603000000000
0!
0*
09
0>
0C
#603010000000
1!
1*
b110 6
19
1>
1C
b110 G
#603020000000
0!
0*
09
0>
0C
#603030000000
1!
1*
b111 6
19
1>
1C
b111 G
#603040000000
0!
0*
09
0>
0C
#603050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#603060000000
0!
0*
09
0>
0C
#603070000000
1!
1*
b1 6
19
1>
1C
b1 G
#603080000000
0!
0*
09
0>
0C
#603090000000
1!
1*
b10 6
19
1>
1C
b10 G
#603100000000
0!
0*
09
0>
0C
#603110000000
1!
1*
b11 6
19
1>
1C
b11 G
#603120000000
0!
0*
09
0>
0C
#603130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#603140000000
0!
0*
09
0>
0C
#603150000000
1!
1*
b101 6
19
1>
1C
b101 G
#603160000000
0!
0*
09
0>
0C
#603170000000
1!
1*
b110 6
19
1>
1C
b110 G
#603180000000
0!
0*
09
0>
0C
#603190000000
1!
1*
b111 6
19
1>
1C
b111 G
#603200000000
0!
1"
0*
1+
09
1:
0>
0C
#603210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#603220000000
0!
0*
09
0>
0C
#603230000000
1!
1*
b1 6
19
1>
1C
b1 G
#603240000000
0!
0*
09
0>
0C
#603250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#603260000000
0!
0*
09
0>
0C
#603270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#603280000000
0!
0*
09
0>
0C
#603290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#603300000000
0!
0*
09
0>
0C
#603310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#603320000000
0!
0#
0*
0,
09
0>
0?
0C
#603330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#603340000000
0!
0*
09
0>
0C
#603350000000
1!
1*
19
1>
1C
#603360000000
0!
0*
09
0>
0C
#603370000000
1!
1*
19
1>
1C
#603380000000
0!
0*
09
0>
0C
#603390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#603400000000
0!
0*
09
0>
0C
#603410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#603420000000
0!
0*
09
0>
0C
#603430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#603440000000
0!
0*
09
0>
0C
#603450000000
1!
1*
b10 6
19
1>
1C
b10 G
#603460000000
0!
0*
09
0>
0C
#603470000000
1!
1*
b11 6
19
1>
1C
b11 G
#603480000000
0!
0*
09
0>
0C
#603490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#603500000000
0!
0*
09
0>
0C
#603510000000
1!
1*
b101 6
19
1>
1C
b101 G
#603520000000
0!
0*
09
0>
0C
#603530000000
1!
1*
b110 6
19
1>
1C
b110 G
#603540000000
0!
0*
09
0>
0C
#603550000000
1!
1*
b111 6
19
1>
1C
b111 G
#603560000000
0!
0*
09
0>
0C
#603570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#603580000000
0!
0*
09
0>
0C
#603590000000
1!
1*
b1 6
19
1>
1C
b1 G
#603600000000
0!
0*
09
0>
0C
#603610000000
1!
1*
b10 6
19
1>
1C
b10 G
#603620000000
0!
0*
09
0>
0C
#603630000000
1!
1*
b11 6
19
1>
1C
b11 G
#603640000000
0!
0*
09
0>
0C
#603650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#603660000000
0!
0*
09
0>
0C
#603670000000
1!
1*
b101 6
19
1>
1C
b101 G
#603680000000
0!
0*
09
0>
0C
#603690000000
1!
1*
b110 6
19
1>
1C
b110 G
#603700000000
0!
0*
09
0>
0C
#603710000000
1!
1*
b111 6
19
1>
1C
b111 G
#603720000000
0!
0*
09
0>
0C
#603730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#603740000000
0!
0*
09
0>
0C
#603750000000
1!
1*
b1 6
19
1>
1C
b1 G
#603760000000
0!
0*
09
0>
0C
#603770000000
1!
1*
b10 6
19
1>
1C
b10 G
#603780000000
0!
0*
09
0>
0C
#603790000000
1!
1*
b11 6
19
1>
1C
b11 G
#603800000000
0!
0*
09
0>
0C
#603810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#603820000000
0!
0*
09
0>
0C
#603830000000
1!
1*
b101 6
19
1>
1C
b101 G
#603840000000
0!
0*
09
0>
0C
#603850000000
1!
1*
b110 6
19
1>
1C
b110 G
#603860000000
0!
0*
09
0>
0C
#603870000000
1!
1*
b111 6
19
1>
1C
b111 G
#603880000000
0!
1"
0*
1+
09
1:
0>
0C
#603890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#603900000000
0!
0*
09
0>
0C
#603910000000
1!
1*
b1 6
19
1>
1C
b1 G
#603920000000
0!
0*
09
0>
0C
#603930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#603940000000
0!
0*
09
0>
0C
#603950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#603960000000
0!
0*
09
0>
0C
#603970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#603980000000
0!
0*
09
0>
0C
#603990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#604000000000
0!
0#
0*
0,
09
0>
0?
0C
#604010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#604020000000
0!
0*
09
0>
0C
#604030000000
1!
1*
19
1>
1C
#604040000000
0!
0*
09
0>
0C
#604050000000
1!
1*
19
1>
1C
#604060000000
0!
0*
09
0>
0C
#604070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#604080000000
0!
0*
09
0>
0C
#604090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#604100000000
0!
0*
09
0>
0C
#604110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#604120000000
0!
0*
09
0>
0C
#604130000000
1!
1*
b10 6
19
1>
1C
b10 G
#604140000000
0!
0*
09
0>
0C
#604150000000
1!
1*
b11 6
19
1>
1C
b11 G
#604160000000
0!
0*
09
0>
0C
#604170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#604180000000
0!
0*
09
0>
0C
#604190000000
1!
1*
b101 6
19
1>
1C
b101 G
#604200000000
0!
0*
09
0>
0C
#604210000000
1!
1*
b110 6
19
1>
1C
b110 G
#604220000000
0!
0*
09
0>
0C
#604230000000
1!
1*
b111 6
19
1>
1C
b111 G
#604240000000
0!
0*
09
0>
0C
#604250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#604260000000
0!
0*
09
0>
0C
#604270000000
1!
1*
b1 6
19
1>
1C
b1 G
#604280000000
0!
0*
09
0>
0C
#604290000000
1!
1*
b10 6
19
1>
1C
b10 G
#604300000000
0!
0*
09
0>
0C
#604310000000
1!
1*
b11 6
19
1>
1C
b11 G
#604320000000
0!
0*
09
0>
0C
#604330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#604340000000
0!
0*
09
0>
0C
#604350000000
1!
1*
b101 6
19
1>
1C
b101 G
#604360000000
0!
0*
09
0>
0C
#604370000000
1!
1*
b110 6
19
1>
1C
b110 G
#604380000000
0!
0*
09
0>
0C
#604390000000
1!
1*
b111 6
19
1>
1C
b111 G
#604400000000
0!
0*
09
0>
0C
#604410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#604420000000
0!
0*
09
0>
0C
#604430000000
1!
1*
b1 6
19
1>
1C
b1 G
#604440000000
0!
0*
09
0>
0C
#604450000000
1!
1*
b10 6
19
1>
1C
b10 G
#604460000000
0!
0*
09
0>
0C
#604470000000
1!
1*
b11 6
19
1>
1C
b11 G
#604480000000
0!
0*
09
0>
0C
#604490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#604500000000
0!
0*
09
0>
0C
#604510000000
1!
1*
b101 6
19
1>
1C
b101 G
#604520000000
0!
0*
09
0>
0C
#604530000000
1!
1*
b110 6
19
1>
1C
b110 G
#604540000000
0!
0*
09
0>
0C
#604550000000
1!
1*
b111 6
19
1>
1C
b111 G
#604560000000
0!
1"
0*
1+
09
1:
0>
0C
#604570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#604580000000
0!
0*
09
0>
0C
#604590000000
1!
1*
b1 6
19
1>
1C
b1 G
#604600000000
0!
0*
09
0>
0C
#604610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#604620000000
0!
0*
09
0>
0C
#604630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#604640000000
0!
0*
09
0>
0C
#604650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#604660000000
0!
0*
09
0>
0C
#604670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#604680000000
0!
0#
0*
0,
09
0>
0?
0C
#604690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#604700000000
0!
0*
09
0>
0C
#604710000000
1!
1*
19
1>
1C
#604720000000
0!
0*
09
0>
0C
#604730000000
1!
1*
19
1>
1C
#604740000000
0!
0*
09
0>
0C
#604750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#604760000000
0!
0*
09
0>
0C
#604770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#604780000000
0!
0*
09
0>
0C
#604790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#604800000000
0!
0*
09
0>
0C
#604810000000
1!
1*
b10 6
19
1>
1C
b10 G
#604820000000
0!
0*
09
0>
0C
#604830000000
1!
1*
b11 6
19
1>
1C
b11 G
#604840000000
0!
0*
09
0>
0C
#604850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#604860000000
0!
0*
09
0>
0C
#604870000000
1!
1*
b101 6
19
1>
1C
b101 G
#604880000000
0!
0*
09
0>
0C
#604890000000
1!
1*
b110 6
19
1>
1C
b110 G
#604900000000
0!
0*
09
0>
0C
#604910000000
1!
1*
b111 6
19
1>
1C
b111 G
#604920000000
0!
0*
09
0>
0C
#604930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#604940000000
0!
0*
09
0>
0C
#604950000000
1!
1*
b1 6
19
1>
1C
b1 G
#604960000000
0!
0*
09
0>
0C
#604970000000
1!
1*
b10 6
19
1>
1C
b10 G
#604980000000
0!
0*
09
0>
0C
#604990000000
1!
1*
b11 6
19
1>
1C
b11 G
#605000000000
0!
0*
09
0>
0C
#605010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#605020000000
0!
0*
09
0>
0C
#605030000000
1!
1*
b101 6
19
1>
1C
b101 G
#605040000000
0!
0*
09
0>
0C
#605050000000
1!
1*
b110 6
19
1>
1C
b110 G
#605060000000
0!
0*
09
0>
0C
#605070000000
1!
1*
b111 6
19
1>
1C
b111 G
#605080000000
0!
0*
09
0>
0C
#605090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#605100000000
0!
0*
09
0>
0C
#605110000000
1!
1*
b1 6
19
1>
1C
b1 G
#605120000000
0!
0*
09
0>
0C
#605130000000
1!
1*
b10 6
19
1>
1C
b10 G
#605140000000
0!
0*
09
0>
0C
#605150000000
1!
1*
b11 6
19
1>
1C
b11 G
#605160000000
0!
0*
09
0>
0C
#605170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#605180000000
0!
0*
09
0>
0C
#605190000000
1!
1*
b101 6
19
1>
1C
b101 G
#605200000000
0!
0*
09
0>
0C
#605210000000
1!
1*
b110 6
19
1>
1C
b110 G
#605220000000
0!
0*
09
0>
0C
#605230000000
1!
1*
b111 6
19
1>
1C
b111 G
#605240000000
0!
1"
0*
1+
09
1:
0>
0C
#605250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#605260000000
0!
0*
09
0>
0C
#605270000000
1!
1*
b1 6
19
1>
1C
b1 G
#605280000000
0!
0*
09
0>
0C
#605290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#605300000000
0!
0*
09
0>
0C
#605310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#605320000000
0!
0*
09
0>
0C
#605330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#605340000000
0!
0*
09
0>
0C
#605350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#605360000000
0!
0#
0*
0,
09
0>
0?
0C
#605370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#605380000000
0!
0*
09
0>
0C
#605390000000
1!
1*
19
1>
1C
#605400000000
0!
0*
09
0>
0C
#605410000000
1!
1*
19
1>
1C
#605420000000
0!
0*
09
0>
0C
#605430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#605440000000
0!
0*
09
0>
0C
#605450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#605460000000
0!
0*
09
0>
0C
#605470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#605480000000
0!
0*
09
0>
0C
#605490000000
1!
1*
b10 6
19
1>
1C
b10 G
#605500000000
0!
0*
09
0>
0C
#605510000000
1!
1*
b11 6
19
1>
1C
b11 G
#605520000000
0!
0*
09
0>
0C
#605530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#605540000000
0!
0*
09
0>
0C
#605550000000
1!
1*
b101 6
19
1>
1C
b101 G
#605560000000
0!
0*
09
0>
0C
#605570000000
1!
1*
b110 6
19
1>
1C
b110 G
#605580000000
0!
0*
09
0>
0C
#605590000000
1!
1*
b111 6
19
1>
1C
b111 G
#605600000000
0!
0*
09
0>
0C
#605610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#605620000000
0!
0*
09
0>
0C
#605630000000
1!
1*
b1 6
19
1>
1C
b1 G
#605640000000
0!
0*
09
0>
0C
#605650000000
1!
1*
b10 6
19
1>
1C
b10 G
#605660000000
0!
0*
09
0>
0C
#605670000000
1!
1*
b11 6
19
1>
1C
b11 G
#605680000000
0!
0*
09
0>
0C
#605690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#605700000000
0!
0*
09
0>
0C
#605710000000
1!
1*
b101 6
19
1>
1C
b101 G
#605720000000
0!
0*
09
0>
0C
#605730000000
1!
1*
b110 6
19
1>
1C
b110 G
#605740000000
0!
0*
09
0>
0C
#605750000000
1!
1*
b111 6
19
1>
1C
b111 G
#605760000000
0!
0*
09
0>
0C
#605770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#605780000000
0!
0*
09
0>
0C
#605790000000
1!
1*
b1 6
19
1>
1C
b1 G
#605800000000
0!
0*
09
0>
0C
#605810000000
1!
1*
b10 6
19
1>
1C
b10 G
#605820000000
0!
0*
09
0>
0C
#605830000000
1!
1*
b11 6
19
1>
1C
b11 G
#605840000000
0!
0*
09
0>
0C
#605850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#605860000000
0!
0*
09
0>
0C
#605870000000
1!
1*
b101 6
19
1>
1C
b101 G
#605880000000
0!
0*
09
0>
0C
#605890000000
1!
1*
b110 6
19
1>
1C
b110 G
#605900000000
0!
0*
09
0>
0C
#605910000000
1!
1*
b111 6
19
1>
1C
b111 G
#605920000000
0!
1"
0*
1+
09
1:
0>
0C
#605930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#605940000000
0!
0*
09
0>
0C
#605950000000
1!
1*
b1 6
19
1>
1C
b1 G
#605960000000
0!
0*
09
0>
0C
#605970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#605980000000
0!
0*
09
0>
0C
#605990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#606000000000
0!
0*
09
0>
0C
#606010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#606020000000
0!
0*
09
0>
0C
#606030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#606040000000
0!
0#
0*
0,
09
0>
0?
0C
#606050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#606060000000
0!
0*
09
0>
0C
#606070000000
1!
1*
19
1>
1C
#606080000000
0!
0*
09
0>
0C
#606090000000
1!
1*
19
1>
1C
#606100000000
0!
0*
09
0>
0C
#606110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#606120000000
0!
0*
09
0>
0C
#606130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#606140000000
0!
0*
09
0>
0C
#606150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#606160000000
0!
0*
09
0>
0C
#606170000000
1!
1*
b10 6
19
1>
1C
b10 G
#606180000000
0!
0*
09
0>
0C
#606190000000
1!
1*
b11 6
19
1>
1C
b11 G
#606200000000
0!
0*
09
0>
0C
#606210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#606220000000
0!
0*
09
0>
0C
#606230000000
1!
1*
b101 6
19
1>
1C
b101 G
#606240000000
0!
0*
09
0>
0C
#606250000000
1!
1*
b110 6
19
1>
1C
b110 G
#606260000000
0!
0*
09
0>
0C
#606270000000
1!
1*
b111 6
19
1>
1C
b111 G
#606280000000
0!
0*
09
0>
0C
#606290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#606300000000
0!
0*
09
0>
0C
#606310000000
1!
1*
b1 6
19
1>
1C
b1 G
#606320000000
0!
0*
09
0>
0C
#606330000000
1!
1*
b10 6
19
1>
1C
b10 G
#606340000000
0!
0*
09
0>
0C
#606350000000
1!
1*
b11 6
19
1>
1C
b11 G
#606360000000
0!
0*
09
0>
0C
#606370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#606380000000
0!
0*
09
0>
0C
#606390000000
1!
1*
b101 6
19
1>
1C
b101 G
#606400000000
0!
0*
09
0>
0C
#606410000000
1!
1*
b110 6
19
1>
1C
b110 G
#606420000000
0!
0*
09
0>
0C
#606430000000
1!
1*
b111 6
19
1>
1C
b111 G
#606440000000
0!
0*
09
0>
0C
#606450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#606460000000
0!
0*
09
0>
0C
#606470000000
1!
1*
b1 6
19
1>
1C
b1 G
#606480000000
0!
0*
09
0>
0C
#606490000000
1!
1*
b10 6
19
1>
1C
b10 G
#606500000000
0!
0*
09
0>
0C
#606510000000
1!
1*
b11 6
19
1>
1C
b11 G
#606520000000
0!
0*
09
0>
0C
#606530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#606540000000
0!
0*
09
0>
0C
#606550000000
1!
1*
b101 6
19
1>
1C
b101 G
#606560000000
0!
0*
09
0>
0C
#606570000000
1!
1*
b110 6
19
1>
1C
b110 G
#606580000000
0!
0*
09
0>
0C
#606590000000
1!
1*
b111 6
19
1>
1C
b111 G
#606600000000
0!
1"
0*
1+
09
1:
0>
0C
#606610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#606620000000
0!
0*
09
0>
0C
#606630000000
1!
1*
b1 6
19
1>
1C
b1 G
#606640000000
0!
0*
09
0>
0C
#606650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#606660000000
0!
0*
09
0>
0C
#606670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#606680000000
0!
0*
09
0>
0C
#606690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#606700000000
0!
0*
09
0>
0C
#606710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#606720000000
0!
0#
0*
0,
09
0>
0?
0C
#606730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#606740000000
0!
0*
09
0>
0C
#606750000000
1!
1*
19
1>
1C
#606760000000
0!
0*
09
0>
0C
#606770000000
1!
1*
19
1>
1C
#606780000000
0!
0*
09
0>
0C
#606790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#606800000000
0!
0*
09
0>
0C
#606810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#606820000000
0!
0*
09
0>
0C
#606830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#606840000000
0!
0*
09
0>
0C
#606850000000
1!
1*
b10 6
19
1>
1C
b10 G
#606860000000
0!
0*
09
0>
0C
#606870000000
1!
1*
b11 6
19
1>
1C
b11 G
#606880000000
0!
0*
09
0>
0C
#606890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#606900000000
0!
0*
09
0>
0C
#606910000000
1!
1*
b101 6
19
1>
1C
b101 G
#606920000000
0!
0*
09
0>
0C
#606930000000
1!
1*
b110 6
19
1>
1C
b110 G
#606940000000
0!
0*
09
0>
0C
#606950000000
1!
1*
b111 6
19
1>
1C
b111 G
#606960000000
0!
0*
09
0>
0C
#606970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#606980000000
0!
0*
09
0>
0C
#606990000000
1!
1*
b1 6
19
1>
1C
b1 G
#607000000000
0!
0*
09
0>
0C
#607010000000
1!
1*
b10 6
19
1>
1C
b10 G
#607020000000
0!
0*
09
0>
0C
#607030000000
1!
1*
b11 6
19
1>
1C
b11 G
#607040000000
0!
0*
09
0>
0C
#607050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#607060000000
0!
0*
09
0>
0C
#607070000000
1!
1*
b101 6
19
1>
1C
b101 G
#607080000000
0!
0*
09
0>
0C
#607090000000
1!
1*
b110 6
19
1>
1C
b110 G
#607100000000
0!
0*
09
0>
0C
#607110000000
1!
1*
b111 6
19
1>
1C
b111 G
#607120000000
0!
0*
09
0>
0C
#607130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#607140000000
0!
0*
09
0>
0C
#607150000000
1!
1*
b1 6
19
1>
1C
b1 G
#607160000000
0!
0*
09
0>
0C
#607170000000
1!
1*
b10 6
19
1>
1C
b10 G
#607180000000
0!
0*
09
0>
0C
#607190000000
1!
1*
b11 6
19
1>
1C
b11 G
#607200000000
0!
0*
09
0>
0C
#607210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#607220000000
0!
0*
09
0>
0C
#607230000000
1!
1*
b101 6
19
1>
1C
b101 G
#607240000000
0!
0*
09
0>
0C
#607250000000
1!
1*
b110 6
19
1>
1C
b110 G
#607260000000
0!
0*
09
0>
0C
#607270000000
1!
1*
b111 6
19
1>
1C
b111 G
#607280000000
0!
1"
0*
1+
09
1:
0>
0C
#607290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#607300000000
0!
0*
09
0>
0C
#607310000000
1!
1*
b1 6
19
1>
1C
b1 G
#607320000000
0!
0*
09
0>
0C
#607330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#607340000000
0!
0*
09
0>
0C
#607350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#607360000000
0!
0*
09
0>
0C
#607370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#607380000000
0!
0*
09
0>
0C
#607390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#607400000000
0!
0#
0*
0,
09
0>
0?
0C
#607410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#607420000000
0!
0*
09
0>
0C
#607430000000
1!
1*
19
1>
1C
#607440000000
0!
0*
09
0>
0C
#607450000000
1!
1*
19
1>
1C
#607460000000
0!
0*
09
0>
0C
#607470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#607480000000
0!
0*
09
0>
0C
#607490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#607500000000
0!
0*
09
0>
0C
#607510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#607520000000
0!
0*
09
0>
0C
#607530000000
1!
1*
b10 6
19
1>
1C
b10 G
#607540000000
0!
0*
09
0>
0C
#607550000000
1!
1*
b11 6
19
1>
1C
b11 G
#607560000000
0!
0*
09
0>
0C
#607570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#607580000000
0!
0*
09
0>
0C
#607590000000
1!
1*
b101 6
19
1>
1C
b101 G
#607600000000
0!
0*
09
0>
0C
#607610000000
1!
1*
b110 6
19
1>
1C
b110 G
#607620000000
0!
0*
09
0>
0C
#607630000000
1!
1*
b111 6
19
1>
1C
b111 G
#607640000000
0!
0*
09
0>
0C
#607650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#607660000000
0!
0*
09
0>
0C
#607670000000
1!
1*
b1 6
19
1>
1C
b1 G
#607680000000
0!
0*
09
0>
0C
#607690000000
1!
1*
b10 6
19
1>
1C
b10 G
#607700000000
0!
0*
09
0>
0C
#607710000000
1!
1*
b11 6
19
1>
1C
b11 G
#607720000000
0!
0*
09
0>
0C
#607730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#607740000000
0!
0*
09
0>
0C
#607750000000
1!
1*
b101 6
19
1>
1C
b101 G
#607760000000
0!
0*
09
0>
0C
#607770000000
1!
1*
b110 6
19
1>
1C
b110 G
#607780000000
0!
0*
09
0>
0C
#607790000000
1!
1*
b111 6
19
1>
1C
b111 G
#607800000000
0!
0*
09
0>
0C
#607810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#607820000000
0!
0*
09
0>
0C
#607830000000
1!
1*
b1 6
19
1>
1C
b1 G
#607840000000
0!
0*
09
0>
0C
#607850000000
1!
1*
b10 6
19
1>
1C
b10 G
#607860000000
0!
0*
09
0>
0C
#607870000000
1!
1*
b11 6
19
1>
1C
b11 G
#607880000000
0!
0*
09
0>
0C
#607890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#607900000000
0!
0*
09
0>
0C
#607910000000
1!
1*
b101 6
19
1>
1C
b101 G
#607920000000
0!
0*
09
0>
0C
#607930000000
1!
1*
b110 6
19
1>
1C
b110 G
#607940000000
0!
0*
09
0>
0C
#607950000000
1!
1*
b111 6
19
1>
1C
b111 G
#607960000000
0!
1"
0*
1+
09
1:
0>
0C
#607970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#607980000000
0!
0*
09
0>
0C
#607990000000
1!
1*
b1 6
19
1>
1C
b1 G
#608000000000
0!
0*
09
0>
0C
#608010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#608020000000
0!
0*
09
0>
0C
#608030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#608040000000
0!
0*
09
0>
0C
#608050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#608060000000
0!
0*
09
0>
0C
#608070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#608080000000
0!
0#
0*
0,
09
0>
0?
0C
#608090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#608100000000
0!
0*
09
0>
0C
#608110000000
1!
1*
19
1>
1C
#608120000000
0!
0*
09
0>
0C
#608130000000
1!
1*
19
1>
1C
#608140000000
0!
0*
09
0>
0C
#608150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#608160000000
0!
0*
09
0>
0C
#608170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#608180000000
0!
0*
09
0>
0C
#608190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#608200000000
0!
0*
09
0>
0C
#608210000000
1!
1*
b10 6
19
1>
1C
b10 G
#608220000000
0!
0*
09
0>
0C
#608230000000
1!
1*
b11 6
19
1>
1C
b11 G
#608240000000
0!
0*
09
0>
0C
#608250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#608260000000
0!
0*
09
0>
0C
#608270000000
1!
1*
b101 6
19
1>
1C
b101 G
#608280000000
0!
0*
09
0>
0C
#608290000000
1!
1*
b110 6
19
1>
1C
b110 G
#608300000000
0!
0*
09
0>
0C
#608310000000
1!
1*
b111 6
19
1>
1C
b111 G
#608320000000
0!
0*
09
0>
0C
#608330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#608340000000
0!
0*
09
0>
0C
#608350000000
1!
1*
b1 6
19
1>
1C
b1 G
#608360000000
0!
0*
09
0>
0C
#608370000000
1!
1*
b10 6
19
1>
1C
b10 G
#608380000000
0!
0*
09
0>
0C
#608390000000
1!
1*
b11 6
19
1>
1C
b11 G
#608400000000
0!
0*
09
0>
0C
#608410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#608420000000
0!
0*
09
0>
0C
#608430000000
1!
1*
b101 6
19
1>
1C
b101 G
#608440000000
0!
0*
09
0>
0C
#608450000000
1!
1*
b110 6
19
1>
1C
b110 G
#608460000000
0!
0*
09
0>
0C
#608470000000
1!
1*
b111 6
19
1>
1C
b111 G
#608480000000
0!
0*
09
0>
0C
#608490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#608500000000
0!
0*
09
0>
0C
#608510000000
1!
1*
b1 6
19
1>
1C
b1 G
#608520000000
0!
0*
09
0>
0C
#608530000000
1!
1*
b10 6
19
1>
1C
b10 G
#608540000000
0!
0*
09
0>
0C
#608550000000
1!
1*
b11 6
19
1>
1C
b11 G
#608560000000
0!
0*
09
0>
0C
#608570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#608580000000
0!
0*
09
0>
0C
#608590000000
1!
1*
b101 6
19
1>
1C
b101 G
#608600000000
0!
0*
09
0>
0C
#608610000000
1!
1*
b110 6
19
1>
1C
b110 G
#608620000000
0!
0*
09
0>
0C
#608630000000
1!
1*
b111 6
19
1>
1C
b111 G
#608640000000
0!
1"
0*
1+
09
1:
0>
0C
#608650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#608660000000
0!
0*
09
0>
0C
#608670000000
1!
1*
b1 6
19
1>
1C
b1 G
#608680000000
0!
0*
09
0>
0C
#608690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#608700000000
0!
0*
09
0>
0C
#608710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#608720000000
0!
0*
09
0>
0C
#608730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#608740000000
0!
0*
09
0>
0C
#608750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#608760000000
0!
0#
0*
0,
09
0>
0?
0C
#608770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#608780000000
0!
0*
09
0>
0C
#608790000000
1!
1*
19
1>
1C
#608800000000
0!
0*
09
0>
0C
#608810000000
1!
1*
19
1>
1C
#608820000000
0!
0*
09
0>
0C
#608830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#608840000000
0!
0*
09
0>
0C
#608850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#608860000000
0!
0*
09
0>
0C
#608870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#608880000000
0!
0*
09
0>
0C
#608890000000
1!
1*
b10 6
19
1>
1C
b10 G
#608900000000
0!
0*
09
0>
0C
#608910000000
1!
1*
b11 6
19
1>
1C
b11 G
#608920000000
0!
0*
09
0>
0C
#608930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#608940000000
0!
0*
09
0>
0C
#608950000000
1!
1*
b101 6
19
1>
1C
b101 G
#608960000000
0!
0*
09
0>
0C
#608970000000
1!
1*
b110 6
19
1>
1C
b110 G
#608980000000
0!
0*
09
0>
0C
#608990000000
1!
1*
b111 6
19
1>
1C
b111 G
#609000000000
0!
0*
09
0>
0C
#609010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#609020000000
0!
0*
09
0>
0C
#609030000000
1!
1*
b1 6
19
1>
1C
b1 G
#609040000000
0!
0*
09
0>
0C
#609050000000
1!
1*
b10 6
19
1>
1C
b10 G
#609060000000
0!
0*
09
0>
0C
#609070000000
1!
1*
b11 6
19
1>
1C
b11 G
#609080000000
0!
0*
09
0>
0C
#609090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#609100000000
0!
0*
09
0>
0C
#609110000000
1!
1*
b101 6
19
1>
1C
b101 G
#609120000000
0!
0*
09
0>
0C
#609130000000
1!
1*
b110 6
19
1>
1C
b110 G
#609140000000
0!
0*
09
0>
0C
#609150000000
1!
1*
b111 6
19
1>
1C
b111 G
#609160000000
0!
0*
09
0>
0C
#609170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#609180000000
0!
0*
09
0>
0C
#609190000000
1!
1*
b1 6
19
1>
1C
b1 G
#609200000000
0!
0*
09
0>
0C
#609210000000
1!
1*
b10 6
19
1>
1C
b10 G
#609220000000
0!
0*
09
0>
0C
#609230000000
1!
1*
b11 6
19
1>
1C
b11 G
#609240000000
0!
0*
09
0>
0C
#609250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#609260000000
0!
0*
09
0>
0C
#609270000000
1!
1*
b101 6
19
1>
1C
b101 G
#609280000000
0!
0*
09
0>
0C
#609290000000
1!
1*
b110 6
19
1>
1C
b110 G
#609300000000
0!
0*
09
0>
0C
#609310000000
1!
1*
b111 6
19
1>
1C
b111 G
#609320000000
0!
1"
0*
1+
09
1:
0>
0C
#609330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#609340000000
0!
0*
09
0>
0C
#609350000000
1!
1*
b1 6
19
1>
1C
b1 G
#609360000000
0!
0*
09
0>
0C
#609370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#609380000000
0!
0*
09
0>
0C
#609390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#609400000000
0!
0*
09
0>
0C
#609410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#609420000000
0!
0*
09
0>
0C
#609430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#609440000000
0!
0#
0*
0,
09
0>
0?
0C
#609450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#609460000000
0!
0*
09
0>
0C
#609470000000
1!
1*
19
1>
1C
#609480000000
0!
0*
09
0>
0C
#609490000000
1!
1*
19
1>
1C
#609500000000
0!
0*
09
0>
0C
#609510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#609520000000
0!
0*
09
0>
0C
#609530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#609540000000
0!
0*
09
0>
0C
#609550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#609560000000
0!
0*
09
0>
0C
#609570000000
1!
1*
b10 6
19
1>
1C
b10 G
#609580000000
0!
0*
09
0>
0C
#609590000000
1!
1*
b11 6
19
1>
1C
b11 G
#609600000000
0!
0*
09
0>
0C
#609610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#609620000000
0!
0*
09
0>
0C
#609630000000
1!
1*
b101 6
19
1>
1C
b101 G
#609640000000
0!
0*
09
0>
0C
#609650000000
1!
1*
b110 6
19
1>
1C
b110 G
#609660000000
0!
0*
09
0>
0C
#609670000000
1!
1*
b111 6
19
1>
1C
b111 G
#609680000000
0!
0*
09
0>
0C
#609690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#609700000000
0!
0*
09
0>
0C
#609710000000
1!
1*
b1 6
19
1>
1C
b1 G
#609720000000
0!
0*
09
0>
0C
#609730000000
1!
1*
b10 6
19
1>
1C
b10 G
#609740000000
0!
0*
09
0>
0C
#609750000000
1!
1*
b11 6
19
1>
1C
b11 G
#609760000000
0!
0*
09
0>
0C
#609770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#609780000000
0!
0*
09
0>
0C
#609790000000
1!
1*
b101 6
19
1>
1C
b101 G
#609800000000
0!
0*
09
0>
0C
#609810000000
1!
1*
b110 6
19
1>
1C
b110 G
#609820000000
0!
0*
09
0>
0C
#609830000000
1!
1*
b111 6
19
1>
1C
b111 G
#609840000000
0!
0*
09
0>
0C
#609850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#609860000000
0!
0*
09
0>
0C
#609870000000
1!
1*
b1 6
19
1>
1C
b1 G
#609880000000
0!
0*
09
0>
0C
#609890000000
1!
1*
b10 6
19
1>
1C
b10 G
#609900000000
0!
0*
09
0>
0C
#609910000000
1!
1*
b11 6
19
1>
1C
b11 G
#609920000000
0!
0*
09
0>
0C
#609930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#609940000000
0!
0*
09
0>
0C
#609950000000
1!
1*
b101 6
19
1>
1C
b101 G
#609960000000
0!
0*
09
0>
0C
#609970000000
1!
1*
b110 6
19
1>
1C
b110 G
#609980000000
0!
0*
09
0>
0C
#609990000000
1!
1*
b111 6
19
1>
1C
b111 G
#610000000000
0!
1"
0*
1+
09
1:
0>
0C
#610010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#610020000000
0!
0*
09
0>
0C
#610030000000
1!
1*
b1 6
19
1>
1C
b1 G
#610040000000
0!
0*
09
0>
0C
#610050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#610060000000
0!
0*
09
0>
0C
#610070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#610080000000
0!
0*
09
0>
0C
#610090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#610100000000
0!
0*
09
0>
0C
#610110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#610120000000
0!
0#
0*
0,
09
0>
0?
0C
#610130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#610140000000
0!
0*
09
0>
0C
#610150000000
1!
1*
19
1>
1C
#610160000000
0!
0*
09
0>
0C
#610170000000
1!
1*
19
1>
1C
#610180000000
0!
0*
09
0>
0C
#610190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#610200000000
0!
0*
09
0>
0C
#610210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#610220000000
0!
0*
09
0>
0C
#610230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#610240000000
0!
0*
09
0>
0C
#610250000000
1!
1*
b10 6
19
1>
1C
b10 G
#610260000000
0!
0*
09
0>
0C
#610270000000
1!
1*
b11 6
19
1>
1C
b11 G
#610280000000
0!
0*
09
0>
0C
#610290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#610300000000
0!
0*
09
0>
0C
#610310000000
1!
1*
b101 6
19
1>
1C
b101 G
#610320000000
0!
0*
09
0>
0C
#610330000000
1!
1*
b110 6
19
1>
1C
b110 G
#610340000000
0!
0*
09
0>
0C
#610350000000
1!
1*
b111 6
19
1>
1C
b111 G
#610360000000
0!
0*
09
0>
0C
#610370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#610380000000
0!
0*
09
0>
0C
#610390000000
1!
1*
b1 6
19
1>
1C
b1 G
#610400000000
0!
0*
09
0>
0C
#610410000000
1!
1*
b10 6
19
1>
1C
b10 G
#610420000000
0!
0*
09
0>
0C
#610430000000
1!
1*
b11 6
19
1>
1C
b11 G
#610440000000
0!
0*
09
0>
0C
#610450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#610460000000
0!
0*
09
0>
0C
#610470000000
1!
1*
b101 6
19
1>
1C
b101 G
#610480000000
0!
0*
09
0>
0C
#610490000000
1!
1*
b110 6
19
1>
1C
b110 G
#610500000000
0!
0*
09
0>
0C
#610510000000
1!
1*
b111 6
19
1>
1C
b111 G
#610520000000
0!
0*
09
0>
0C
#610530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#610540000000
0!
0*
09
0>
0C
#610550000000
1!
1*
b1 6
19
1>
1C
b1 G
#610560000000
0!
0*
09
0>
0C
#610570000000
1!
1*
b10 6
19
1>
1C
b10 G
#610580000000
0!
0*
09
0>
0C
#610590000000
1!
1*
b11 6
19
1>
1C
b11 G
#610600000000
0!
0*
09
0>
0C
#610610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#610620000000
0!
0*
09
0>
0C
#610630000000
1!
1*
b101 6
19
1>
1C
b101 G
#610640000000
0!
0*
09
0>
0C
#610650000000
1!
1*
b110 6
19
1>
1C
b110 G
#610660000000
0!
0*
09
0>
0C
#610670000000
1!
1*
b111 6
19
1>
1C
b111 G
#610680000000
0!
1"
0*
1+
09
1:
0>
0C
#610690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#610700000000
0!
0*
09
0>
0C
#610710000000
1!
1*
b1 6
19
1>
1C
b1 G
#610720000000
0!
0*
09
0>
0C
#610730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#610740000000
0!
0*
09
0>
0C
#610750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#610760000000
0!
0*
09
0>
0C
#610770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#610780000000
0!
0*
09
0>
0C
#610790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#610800000000
0!
0#
0*
0,
09
0>
0?
0C
#610810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#610820000000
0!
0*
09
0>
0C
#610830000000
1!
1*
19
1>
1C
#610840000000
0!
0*
09
0>
0C
#610850000000
1!
1*
19
1>
1C
#610860000000
0!
0*
09
0>
0C
#610870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#610880000000
0!
0*
09
0>
0C
#610890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#610900000000
0!
0*
09
0>
0C
#610910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#610920000000
0!
0*
09
0>
0C
#610930000000
1!
1*
b10 6
19
1>
1C
b10 G
#610940000000
0!
0*
09
0>
0C
#610950000000
1!
1*
b11 6
19
1>
1C
b11 G
#610960000000
0!
0*
09
0>
0C
#610970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#610980000000
0!
0*
09
0>
0C
#610990000000
1!
1*
b101 6
19
1>
1C
b101 G
#611000000000
0!
0*
09
0>
0C
#611010000000
1!
1*
b110 6
19
1>
1C
b110 G
#611020000000
0!
0*
09
0>
0C
#611030000000
1!
1*
b111 6
19
1>
1C
b111 G
#611040000000
0!
0*
09
0>
0C
#611050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#611060000000
0!
0*
09
0>
0C
#611070000000
1!
1*
b1 6
19
1>
1C
b1 G
#611080000000
0!
0*
09
0>
0C
#611090000000
1!
1*
b10 6
19
1>
1C
b10 G
#611100000000
0!
0*
09
0>
0C
#611110000000
1!
1*
b11 6
19
1>
1C
b11 G
#611120000000
0!
0*
09
0>
0C
#611130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#611140000000
0!
0*
09
0>
0C
#611150000000
1!
1*
b101 6
19
1>
1C
b101 G
#611160000000
0!
0*
09
0>
0C
#611170000000
1!
1*
b110 6
19
1>
1C
b110 G
#611180000000
0!
0*
09
0>
0C
#611190000000
1!
1*
b111 6
19
1>
1C
b111 G
#611200000000
0!
0*
09
0>
0C
#611210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#611220000000
0!
0*
09
0>
0C
#611230000000
1!
1*
b1 6
19
1>
1C
b1 G
#611240000000
0!
0*
09
0>
0C
#611250000000
1!
1*
b10 6
19
1>
1C
b10 G
#611260000000
0!
0*
09
0>
0C
#611270000000
1!
1*
b11 6
19
1>
1C
b11 G
#611280000000
0!
0*
09
0>
0C
#611290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#611300000000
0!
0*
09
0>
0C
#611310000000
1!
1*
b101 6
19
1>
1C
b101 G
#611320000000
0!
0*
09
0>
0C
#611330000000
1!
1*
b110 6
19
1>
1C
b110 G
#611340000000
0!
0*
09
0>
0C
#611350000000
1!
1*
b111 6
19
1>
1C
b111 G
#611360000000
0!
1"
0*
1+
09
1:
0>
0C
#611370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#611380000000
0!
0*
09
0>
0C
#611390000000
1!
1*
b1 6
19
1>
1C
b1 G
#611400000000
0!
0*
09
0>
0C
#611410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#611420000000
0!
0*
09
0>
0C
#611430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#611440000000
0!
0*
09
0>
0C
#611450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#611460000000
0!
0*
09
0>
0C
#611470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#611480000000
0!
0#
0*
0,
09
0>
0?
0C
#611490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#611500000000
0!
0*
09
0>
0C
#611510000000
1!
1*
19
1>
1C
#611520000000
0!
0*
09
0>
0C
#611530000000
1!
1*
19
1>
1C
#611540000000
0!
0*
09
0>
0C
#611550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#611560000000
0!
0*
09
0>
0C
#611570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#611580000000
0!
0*
09
0>
0C
#611590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#611600000000
0!
0*
09
0>
0C
#611610000000
1!
1*
b10 6
19
1>
1C
b10 G
#611620000000
0!
0*
09
0>
0C
#611630000000
1!
1*
b11 6
19
1>
1C
b11 G
#611640000000
0!
0*
09
0>
0C
#611650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#611660000000
0!
0*
09
0>
0C
#611670000000
1!
1*
b101 6
19
1>
1C
b101 G
#611680000000
0!
0*
09
0>
0C
#611690000000
1!
1*
b110 6
19
1>
1C
b110 G
#611700000000
0!
0*
09
0>
0C
#611710000000
1!
1*
b111 6
19
1>
1C
b111 G
#611720000000
0!
0*
09
0>
0C
#611730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#611740000000
0!
0*
09
0>
0C
#611750000000
1!
1*
b1 6
19
1>
1C
b1 G
#611760000000
0!
0*
09
0>
0C
#611770000000
1!
1*
b10 6
19
1>
1C
b10 G
#611780000000
0!
0*
09
0>
0C
#611790000000
1!
1*
b11 6
19
1>
1C
b11 G
#611800000000
0!
0*
09
0>
0C
#611810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#611820000000
0!
0*
09
0>
0C
#611830000000
1!
1*
b101 6
19
1>
1C
b101 G
#611840000000
0!
0*
09
0>
0C
#611850000000
1!
1*
b110 6
19
1>
1C
b110 G
#611860000000
0!
0*
09
0>
0C
#611870000000
1!
1*
b111 6
19
1>
1C
b111 G
#611880000000
0!
0*
09
0>
0C
#611890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#611900000000
0!
0*
09
0>
0C
#611910000000
1!
1*
b1 6
19
1>
1C
b1 G
#611920000000
0!
0*
09
0>
0C
#611930000000
1!
1*
b10 6
19
1>
1C
b10 G
#611940000000
0!
0*
09
0>
0C
#611950000000
1!
1*
b11 6
19
1>
1C
b11 G
#611960000000
0!
0*
09
0>
0C
#611970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#611980000000
0!
0*
09
0>
0C
#611990000000
1!
1*
b101 6
19
1>
1C
b101 G
#612000000000
0!
0*
09
0>
0C
#612010000000
1!
1*
b110 6
19
1>
1C
b110 G
#612020000000
0!
0*
09
0>
0C
#612030000000
1!
1*
b111 6
19
1>
1C
b111 G
#612040000000
0!
1"
0*
1+
09
1:
0>
0C
#612050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#612060000000
0!
0*
09
0>
0C
#612070000000
1!
1*
b1 6
19
1>
1C
b1 G
#612080000000
0!
0*
09
0>
0C
#612090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#612100000000
0!
0*
09
0>
0C
#612110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#612120000000
0!
0*
09
0>
0C
#612130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#612140000000
0!
0*
09
0>
0C
#612150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#612160000000
0!
0#
0*
0,
09
0>
0?
0C
#612170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#612180000000
0!
0*
09
0>
0C
#612190000000
1!
1*
19
1>
1C
#612200000000
0!
0*
09
0>
0C
#612210000000
1!
1*
19
1>
1C
#612220000000
0!
0*
09
0>
0C
#612230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#612240000000
0!
0*
09
0>
0C
#612250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#612260000000
0!
0*
09
0>
0C
#612270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#612280000000
0!
0*
09
0>
0C
#612290000000
1!
1*
b10 6
19
1>
1C
b10 G
#612300000000
0!
0*
09
0>
0C
#612310000000
1!
1*
b11 6
19
1>
1C
b11 G
#612320000000
0!
0*
09
0>
0C
#612330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#612340000000
0!
0*
09
0>
0C
#612350000000
1!
1*
b101 6
19
1>
1C
b101 G
#612360000000
0!
0*
09
0>
0C
#612370000000
1!
1*
b110 6
19
1>
1C
b110 G
#612380000000
0!
0*
09
0>
0C
#612390000000
1!
1*
b111 6
19
1>
1C
b111 G
#612400000000
0!
0*
09
0>
0C
#612410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#612420000000
0!
0*
09
0>
0C
#612430000000
1!
1*
b1 6
19
1>
1C
b1 G
#612440000000
0!
0*
09
0>
0C
#612450000000
1!
1*
b10 6
19
1>
1C
b10 G
#612460000000
0!
0*
09
0>
0C
#612470000000
1!
1*
b11 6
19
1>
1C
b11 G
#612480000000
0!
0*
09
0>
0C
#612490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#612500000000
0!
0*
09
0>
0C
#612510000000
1!
1*
b101 6
19
1>
1C
b101 G
#612520000000
0!
0*
09
0>
0C
#612530000000
1!
1*
b110 6
19
1>
1C
b110 G
#612540000000
0!
0*
09
0>
0C
#612550000000
1!
1*
b111 6
19
1>
1C
b111 G
#612560000000
0!
0*
09
0>
0C
#612570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#612580000000
0!
0*
09
0>
0C
#612590000000
1!
1*
b1 6
19
1>
1C
b1 G
#612600000000
0!
0*
09
0>
0C
#612610000000
1!
1*
b10 6
19
1>
1C
b10 G
#612620000000
0!
0*
09
0>
0C
#612630000000
1!
1*
b11 6
19
1>
1C
b11 G
#612640000000
0!
0*
09
0>
0C
#612650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#612660000000
0!
0*
09
0>
0C
#612670000000
1!
1*
b101 6
19
1>
1C
b101 G
#612680000000
0!
0*
09
0>
0C
#612690000000
1!
1*
b110 6
19
1>
1C
b110 G
#612700000000
0!
0*
09
0>
0C
#612710000000
1!
1*
b111 6
19
1>
1C
b111 G
#612720000000
0!
1"
0*
1+
09
1:
0>
0C
#612730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#612740000000
0!
0*
09
0>
0C
#612750000000
1!
1*
b1 6
19
1>
1C
b1 G
#612760000000
0!
0*
09
0>
0C
#612770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#612780000000
0!
0*
09
0>
0C
#612790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#612800000000
0!
0*
09
0>
0C
#612810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#612820000000
0!
0*
09
0>
0C
#612830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#612840000000
0!
0#
0*
0,
09
0>
0?
0C
#612850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#612860000000
0!
0*
09
0>
0C
#612870000000
1!
1*
19
1>
1C
#612880000000
0!
0*
09
0>
0C
#612890000000
1!
1*
19
1>
1C
#612900000000
0!
0*
09
0>
0C
#612910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#612920000000
0!
0*
09
0>
0C
#612930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#612940000000
0!
0*
09
0>
0C
#612950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#612960000000
0!
0*
09
0>
0C
#612970000000
1!
1*
b10 6
19
1>
1C
b10 G
#612980000000
0!
0*
09
0>
0C
#612990000000
1!
1*
b11 6
19
1>
1C
b11 G
#613000000000
0!
0*
09
0>
0C
#613010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#613020000000
0!
0*
09
0>
0C
#613030000000
1!
1*
b101 6
19
1>
1C
b101 G
#613040000000
0!
0*
09
0>
0C
#613050000000
1!
1*
b110 6
19
1>
1C
b110 G
#613060000000
0!
0*
09
0>
0C
#613070000000
1!
1*
b111 6
19
1>
1C
b111 G
#613080000000
0!
0*
09
0>
0C
#613090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#613100000000
0!
0*
09
0>
0C
#613110000000
1!
1*
b1 6
19
1>
1C
b1 G
#613120000000
0!
0*
09
0>
0C
#613130000000
1!
1*
b10 6
19
1>
1C
b10 G
#613140000000
0!
0*
09
0>
0C
#613150000000
1!
1*
b11 6
19
1>
1C
b11 G
#613160000000
0!
0*
09
0>
0C
#613170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#613180000000
0!
0*
09
0>
0C
#613190000000
1!
1*
b101 6
19
1>
1C
b101 G
#613200000000
0!
0*
09
0>
0C
#613210000000
1!
1*
b110 6
19
1>
1C
b110 G
#613220000000
0!
0*
09
0>
0C
#613230000000
1!
1*
b111 6
19
1>
1C
b111 G
#613240000000
0!
0*
09
0>
0C
#613250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#613260000000
0!
0*
09
0>
0C
#613270000000
1!
1*
b1 6
19
1>
1C
b1 G
#613280000000
0!
0*
09
0>
0C
#613290000000
1!
1*
b10 6
19
1>
1C
b10 G
#613300000000
0!
0*
09
0>
0C
#613310000000
1!
1*
b11 6
19
1>
1C
b11 G
#613320000000
0!
0*
09
0>
0C
#613330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#613340000000
0!
0*
09
0>
0C
#613350000000
1!
1*
b101 6
19
1>
1C
b101 G
#613360000000
0!
0*
09
0>
0C
#613370000000
1!
1*
b110 6
19
1>
1C
b110 G
#613380000000
0!
0*
09
0>
0C
#613390000000
1!
1*
b111 6
19
1>
1C
b111 G
#613400000000
0!
1"
0*
1+
09
1:
0>
0C
#613410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#613420000000
0!
0*
09
0>
0C
#613430000000
1!
1*
b1 6
19
1>
1C
b1 G
#613440000000
0!
0*
09
0>
0C
#613450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#613460000000
0!
0*
09
0>
0C
#613470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#613480000000
0!
0*
09
0>
0C
#613490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#613500000000
0!
0*
09
0>
0C
#613510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#613520000000
0!
0#
0*
0,
09
0>
0?
0C
#613530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#613540000000
0!
0*
09
0>
0C
#613550000000
1!
1*
19
1>
1C
#613560000000
0!
0*
09
0>
0C
#613570000000
1!
1*
19
1>
1C
#613580000000
0!
0*
09
0>
0C
#613590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#613600000000
0!
0*
09
0>
0C
#613610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#613620000000
0!
0*
09
0>
0C
#613630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#613640000000
0!
0*
09
0>
0C
#613650000000
1!
1*
b10 6
19
1>
1C
b10 G
#613660000000
0!
0*
09
0>
0C
#613670000000
1!
1*
b11 6
19
1>
1C
b11 G
#613680000000
0!
0*
09
0>
0C
#613690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#613700000000
0!
0*
09
0>
0C
#613710000000
1!
1*
b101 6
19
1>
1C
b101 G
#613720000000
0!
0*
09
0>
0C
#613730000000
1!
1*
b110 6
19
1>
1C
b110 G
#613740000000
0!
0*
09
0>
0C
#613750000000
1!
1*
b111 6
19
1>
1C
b111 G
#613760000000
0!
0*
09
0>
0C
#613770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#613780000000
0!
0*
09
0>
0C
#613790000000
1!
1*
b1 6
19
1>
1C
b1 G
#613800000000
0!
0*
09
0>
0C
#613810000000
1!
1*
b10 6
19
1>
1C
b10 G
#613820000000
0!
0*
09
0>
0C
#613830000000
1!
1*
b11 6
19
1>
1C
b11 G
#613840000000
0!
0*
09
0>
0C
#613850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#613860000000
0!
0*
09
0>
0C
#613870000000
1!
1*
b101 6
19
1>
1C
b101 G
#613880000000
0!
0*
09
0>
0C
#613890000000
1!
1*
b110 6
19
1>
1C
b110 G
#613900000000
0!
0*
09
0>
0C
#613910000000
1!
1*
b111 6
19
1>
1C
b111 G
#613920000000
0!
0*
09
0>
0C
#613930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#613940000000
0!
0*
09
0>
0C
#613950000000
1!
1*
b1 6
19
1>
1C
b1 G
#613960000000
0!
0*
09
0>
0C
#613970000000
1!
1*
b10 6
19
1>
1C
b10 G
#613980000000
0!
0*
09
0>
0C
#613990000000
1!
1*
b11 6
19
1>
1C
b11 G
#614000000000
0!
0*
09
0>
0C
#614010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#614020000000
0!
0*
09
0>
0C
#614030000000
1!
1*
b101 6
19
1>
1C
b101 G
#614040000000
0!
0*
09
0>
0C
#614050000000
1!
1*
b110 6
19
1>
1C
b110 G
#614060000000
0!
0*
09
0>
0C
#614070000000
1!
1*
b111 6
19
1>
1C
b111 G
#614080000000
0!
1"
0*
1+
09
1:
0>
0C
#614090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#614100000000
0!
0*
09
0>
0C
#614110000000
1!
1*
b1 6
19
1>
1C
b1 G
#614120000000
0!
0*
09
0>
0C
#614130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#614140000000
0!
0*
09
0>
0C
#614150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#614160000000
0!
0*
09
0>
0C
#614170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#614180000000
0!
0*
09
0>
0C
#614190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#614200000000
0!
0#
0*
0,
09
0>
0?
0C
#614210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#614220000000
0!
0*
09
0>
0C
#614230000000
1!
1*
19
1>
1C
#614240000000
0!
0*
09
0>
0C
#614250000000
1!
1*
19
1>
1C
#614260000000
0!
0*
09
0>
0C
#614270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#614280000000
0!
0*
09
0>
0C
#614290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#614300000000
0!
0*
09
0>
0C
#614310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#614320000000
0!
0*
09
0>
0C
#614330000000
1!
1*
b10 6
19
1>
1C
b10 G
#614340000000
0!
0*
09
0>
0C
#614350000000
1!
1*
b11 6
19
1>
1C
b11 G
#614360000000
0!
0*
09
0>
0C
#614370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#614380000000
0!
0*
09
0>
0C
#614390000000
1!
1*
b101 6
19
1>
1C
b101 G
#614400000000
0!
0*
09
0>
0C
#614410000000
1!
1*
b110 6
19
1>
1C
b110 G
#614420000000
0!
0*
09
0>
0C
#614430000000
1!
1*
b111 6
19
1>
1C
b111 G
#614440000000
0!
0*
09
0>
0C
#614450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#614460000000
0!
0*
09
0>
0C
#614470000000
1!
1*
b1 6
19
1>
1C
b1 G
#614480000000
0!
0*
09
0>
0C
#614490000000
1!
1*
b10 6
19
1>
1C
b10 G
#614500000000
0!
0*
09
0>
0C
#614510000000
1!
1*
b11 6
19
1>
1C
b11 G
#614520000000
0!
0*
09
0>
0C
#614530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#614540000000
0!
0*
09
0>
0C
#614550000000
1!
1*
b101 6
19
1>
1C
b101 G
#614560000000
0!
0*
09
0>
0C
#614570000000
1!
1*
b110 6
19
1>
1C
b110 G
#614580000000
0!
0*
09
0>
0C
#614590000000
1!
1*
b111 6
19
1>
1C
b111 G
#614600000000
0!
0*
09
0>
0C
#614610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#614620000000
0!
0*
09
0>
0C
#614630000000
1!
1*
b1 6
19
1>
1C
b1 G
#614640000000
0!
0*
09
0>
0C
#614650000000
1!
1*
b10 6
19
1>
1C
b10 G
#614660000000
0!
0*
09
0>
0C
#614670000000
1!
1*
b11 6
19
1>
1C
b11 G
#614680000000
0!
0*
09
0>
0C
#614690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#614700000000
0!
0*
09
0>
0C
#614710000000
1!
1*
b101 6
19
1>
1C
b101 G
#614720000000
0!
0*
09
0>
0C
#614730000000
1!
1*
b110 6
19
1>
1C
b110 G
#614740000000
0!
0*
09
0>
0C
#614750000000
1!
1*
b111 6
19
1>
1C
b111 G
#614760000000
0!
1"
0*
1+
09
1:
0>
0C
#614770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#614780000000
0!
0*
09
0>
0C
#614790000000
1!
1*
b1 6
19
1>
1C
b1 G
#614800000000
0!
0*
09
0>
0C
#614810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#614820000000
0!
0*
09
0>
0C
#614830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#614840000000
0!
0*
09
0>
0C
#614850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#614860000000
0!
0*
09
0>
0C
#614870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#614880000000
0!
0#
0*
0,
09
0>
0?
0C
#614890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#614900000000
0!
0*
09
0>
0C
#614910000000
1!
1*
19
1>
1C
#614920000000
0!
0*
09
0>
0C
#614930000000
1!
1*
19
1>
1C
#614940000000
0!
0*
09
0>
0C
#614950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#614960000000
0!
0*
09
0>
0C
#614970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#614980000000
0!
0*
09
0>
0C
#614990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#615000000000
0!
0*
09
0>
0C
#615010000000
1!
1*
b10 6
19
1>
1C
b10 G
#615020000000
0!
0*
09
0>
0C
#615030000000
1!
1*
b11 6
19
1>
1C
b11 G
#615040000000
0!
0*
09
0>
0C
#615050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#615060000000
0!
0*
09
0>
0C
#615070000000
1!
1*
b101 6
19
1>
1C
b101 G
#615080000000
0!
0*
09
0>
0C
#615090000000
1!
1*
b110 6
19
1>
1C
b110 G
#615100000000
0!
0*
09
0>
0C
#615110000000
1!
1*
b111 6
19
1>
1C
b111 G
#615120000000
0!
0*
09
0>
0C
#615130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#615140000000
0!
0*
09
0>
0C
#615150000000
1!
1*
b1 6
19
1>
1C
b1 G
#615160000000
0!
0*
09
0>
0C
#615170000000
1!
1*
b10 6
19
1>
1C
b10 G
#615180000000
0!
0*
09
0>
0C
#615190000000
1!
1*
b11 6
19
1>
1C
b11 G
#615200000000
0!
0*
09
0>
0C
#615210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#615220000000
0!
0*
09
0>
0C
#615230000000
1!
1*
b101 6
19
1>
1C
b101 G
#615240000000
0!
0*
09
0>
0C
#615250000000
1!
1*
b110 6
19
1>
1C
b110 G
#615260000000
0!
0*
09
0>
0C
#615270000000
1!
1*
b111 6
19
1>
1C
b111 G
#615280000000
0!
0*
09
0>
0C
#615290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#615300000000
0!
0*
09
0>
0C
#615310000000
1!
1*
b1 6
19
1>
1C
b1 G
#615320000000
0!
0*
09
0>
0C
#615330000000
1!
1*
b10 6
19
1>
1C
b10 G
#615340000000
0!
0*
09
0>
0C
#615350000000
1!
1*
b11 6
19
1>
1C
b11 G
#615360000000
0!
0*
09
0>
0C
#615370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#615380000000
0!
0*
09
0>
0C
#615390000000
1!
1*
b101 6
19
1>
1C
b101 G
#615400000000
0!
0*
09
0>
0C
#615410000000
1!
1*
b110 6
19
1>
1C
b110 G
#615420000000
0!
0*
09
0>
0C
#615430000000
1!
1*
b111 6
19
1>
1C
b111 G
#615440000000
0!
1"
0*
1+
09
1:
0>
0C
#615450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#615460000000
0!
0*
09
0>
0C
#615470000000
1!
1*
b1 6
19
1>
1C
b1 G
#615480000000
0!
0*
09
0>
0C
#615490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#615500000000
0!
0*
09
0>
0C
#615510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#615520000000
0!
0*
09
0>
0C
#615530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#615540000000
0!
0*
09
0>
0C
#615550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#615560000000
0!
0#
0*
0,
09
0>
0?
0C
#615570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#615580000000
0!
0*
09
0>
0C
#615590000000
1!
1*
19
1>
1C
#615600000000
0!
0*
09
0>
0C
#615610000000
1!
1*
19
1>
1C
#615620000000
0!
0*
09
0>
0C
#615630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#615640000000
0!
0*
09
0>
0C
#615650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#615660000000
0!
0*
09
0>
0C
#615670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#615680000000
0!
0*
09
0>
0C
#615690000000
1!
1*
b10 6
19
1>
1C
b10 G
#615700000000
0!
0*
09
0>
0C
#615710000000
1!
1*
b11 6
19
1>
1C
b11 G
#615720000000
0!
0*
09
0>
0C
#615730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#615740000000
0!
0*
09
0>
0C
#615750000000
1!
1*
b101 6
19
1>
1C
b101 G
#615760000000
0!
0*
09
0>
0C
#615770000000
1!
1*
b110 6
19
1>
1C
b110 G
#615780000000
0!
0*
09
0>
0C
#615790000000
1!
1*
b111 6
19
1>
1C
b111 G
#615800000000
0!
0*
09
0>
0C
#615810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#615820000000
0!
0*
09
0>
0C
#615830000000
1!
1*
b1 6
19
1>
1C
b1 G
#615840000000
0!
0*
09
0>
0C
#615850000000
1!
1*
b10 6
19
1>
1C
b10 G
#615860000000
0!
0*
09
0>
0C
#615870000000
1!
1*
b11 6
19
1>
1C
b11 G
#615880000000
0!
0*
09
0>
0C
#615890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#615900000000
0!
0*
09
0>
0C
#615910000000
1!
1*
b101 6
19
1>
1C
b101 G
#615920000000
0!
0*
09
0>
0C
#615930000000
1!
1*
b110 6
19
1>
1C
b110 G
#615940000000
0!
0*
09
0>
0C
#615950000000
1!
1*
b111 6
19
1>
1C
b111 G
#615960000000
0!
0*
09
0>
0C
#615970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#615980000000
0!
0*
09
0>
0C
#615990000000
1!
1*
b1 6
19
1>
1C
b1 G
#616000000000
0!
0*
09
0>
0C
#616010000000
1!
1*
b10 6
19
1>
1C
b10 G
#616020000000
0!
0*
09
0>
0C
#616030000000
1!
1*
b11 6
19
1>
1C
b11 G
#616040000000
0!
0*
09
0>
0C
#616050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#616060000000
0!
0*
09
0>
0C
#616070000000
1!
1*
b101 6
19
1>
1C
b101 G
#616080000000
0!
0*
09
0>
0C
#616090000000
1!
1*
b110 6
19
1>
1C
b110 G
#616100000000
0!
0*
09
0>
0C
#616110000000
1!
1*
b111 6
19
1>
1C
b111 G
#616120000000
0!
1"
0*
1+
09
1:
0>
0C
#616130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#616140000000
0!
0*
09
0>
0C
#616150000000
1!
1*
b1 6
19
1>
1C
b1 G
#616160000000
0!
0*
09
0>
0C
#616170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#616180000000
0!
0*
09
0>
0C
#616190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#616200000000
0!
0*
09
0>
0C
#616210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#616220000000
0!
0*
09
0>
0C
#616230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#616240000000
0!
0#
0*
0,
09
0>
0?
0C
#616250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#616260000000
0!
0*
09
0>
0C
#616270000000
1!
1*
19
1>
1C
#616280000000
0!
0*
09
0>
0C
#616290000000
1!
1*
19
1>
1C
#616300000000
0!
0*
09
0>
0C
#616310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#616320000000
0!
0*
09
0>
0C
#616330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#616340000000
0!
0*
09
0>
0C
#616350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#616360000000
0!
0*
09
0>
0C
#616370000000
1!
1*
b10 6
19
1>
1C
b10 G
#616380000000
0!
0*
09
0>
0C
#616390000000
1!
1*
b11 6
19
1>
1C
b11 G
#616400000000
0!
0*
09
0>
0C
#616410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#616420000000
0!
0*
09
0>
0C
#616430000000
1!
1*
b101 6
19
1>
1C
b101 G
#616440000000
0!
0*
09
0>
0C
#616450000000
1!
1*
b110 6
19
1>
1C
b110 G
#616460000000
0!
0*
09
0>
0C
#616470000000
1!
1*
b111 6
19
1>
1C
b111 G
#616480000000
0!
0*
09
0>
0C
#616490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#616500000000
0!
0*
09
0>
0C
#616510000000
1!
1*
b1 6
19
1>
1C
b1 G
#616520000000
0!
0*
09
0>
0C
#616530000000
1!
1*
b10 6
19
1>
1C
b10 G
#616540000000
0!
0*
09
0>
0C
#616550000000
1!
1*
b11 6
19
1>
1C
b11 G
#616560000000
0!
0*
09
0>
0C
#616570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#616580000000
0!
0*
09
0>
0C
#616590000000
1!
1*
b101 6
19
1>
1C
b101 G
#616600000000
0!
0*
09
0>
0C
#616610000000
1!
1*
b110 6
19
1>
1C
b110 G
#616620000000
0!
0*
09
0>
0C
#616630000000
1!
1*
b111 6
19
1>
1C
b111 G
#616640000000
0!
0*
09
0>
0C
#616650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#616660000000
0!
0*
09
0>
0C
#616670000000
1!
1*
b1 6
19
1>
1C
b1 G
#616680000000
0!
0*
09
0>
0C
#616690000000
1!
1*
b10 6
19
1>
1C
b10 G
#616700000000
0!
0*
09
0>
0C
#616710000000
1!
1*
b11 6
19
1>
1C
b11 G
#616720000000
0!
0*
09
0>
0C
#616730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#616740000000
0!
0*
09
0>
0C
#616750000000
1!
1*
b101 6
19
1>
1C
b101 G
#616760000000
0!
0*
09
0>
0C
#616770000000
1!
1*
b110 6
19
1>
1C
b110 G
#616780000000
0!
0*
09
0>
0C
#616790000000
1!
1*
b111 6
19
1>
1C
b111 G
#616800000000
0!
1"
0*
1+
09
1:
0>
0C
#616810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#616820000000
0!
0*
09
0>
0C
#616830000000
1!
1*
b1 6
19
1>
1C
b1 G
#616840000000
0!
0*
09
0>
0C
#616850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#616860000000
0!
0*
09
0>
0C
#616870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#616880000000
0!
0*
09
0>
0C
#616890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#616900000000
0!
0*
09
0>
0C
#616910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#616920000000
0!
0#
0*
0,
09
0>
0?
0C
#616930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#616940000000
0!
0*
09
0>
0C
#616950000000
1!
1*
19
1>
1C
#616960000000
0!
0*
09
0>
0C
#616970000000
1!
1*
19
1>
1C
#616980000000
0!
0*
09
0>
0C
#616990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#617000000000
0!
0*
09
0>
0C
#617010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#617020000000
0!
0*
09
0>
0C
#617030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#617040000000
0!
0*
09
0>
0C
#617050000000
1!
1*
b10 6
19
1>
1C
b10 G
#617060000000
0!
0*
09
0>
0C
#617070000000
1!
1*
b11 6
19
1>
1C
b11 G
#617080000000
0!
0*
09
0>
0C
#617090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#617100000000
0!
0*
09
0>
0C
#617110000000
1!
1*
b101 6
19
1>
1C
b101 G
#617120000000
0!
0*
09
0>
0C
#617130000000
1!
1*
b110 6
19
1>
1C
b110 G
#617140000000
0!
0*
09
0>
0C
#617150000000
1!
1*
b111 6
19
1>
1C
b111 G
#617160000000
0!
0*
09
0>
0C
#617170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#617180000000
0!
0*
09
0>
0C
#617190000000
1!
1*
b1 6
19
1>
1C
b1 G
#617200000000
0!
0*
09
0>
0C
#617210000000
1!
1*
b10 6
19
1>
1C
b10 G
#617220000000
0!
0*
09
0>
0C
#617230000000
1!
1*
b11 6
19
1>
1C
b11 G
#617240000000
0!
0*
09
0>
0C
#617250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#617260000000
0!
0*
09
0>
0C
#617270000000
1!
1*
b101 6
19
1>
1C
b101 G
#617280000000
0!
0*
09
0>
0C
#617290000000
1!
1*
b110 6
19
1>
1C
b110 G
#617300000000
0!
0*
09
0>
0C
#617310000000
1!
1*
b111 6
19
1>
1C
b111 G
#617320000000
0!
0*
09
0>
0C
#617330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#617340000000
0!
0*
09
0>
0C
#617350000000
1!
1*
b1 6
19
1>
1C
b1 G
#617360000000
0!
0*
09
0>
0C
#617370000000
1!
1*
b10 6
19
1>
1C
b10 G
#617380000000
0!
0*
09
0>
0C
#617390000000
1!
1*
b11 6
19
1>
1C
b11 G
#617400000000
0!
0*
09
0>
0C
#617410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#617420000000
0!
0*
09
0>
0C
#617430000000
1!
1*
b101 6
19
1>
1C
b101 G
#617440000000
0!
0*
09
0>
0C
#617450000000
1!
1*
b110 6
19
1>
1C
b110 G
#617460000000
0!
0*
09
0>
0C
#617470000000
1!
1*
b111 6
19
1>
1C
b111 G
#617480000000
0!
1"
0*
1+
09
1:
0>
0C
#617490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#617500000000
0!
0*
09
0>
0C
#617510000000
1!
1*
b1 6
19
1>
1C
b1 G
#617520000000
0!
0*
09
0>
0C
#617530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#617540000000
0!
0*
09
0>
0C
#617550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#617560000000
0!
0*
09
0>
0C
#617570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#617580000000
0!
0*
09
0>
0C
#617590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#617600000000
0!
0#
0*
0,
09
0>
0?
0C
#617610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#617620000000
0!
0*
09
0>
0C
#617630000000
1!
1*
19
1>
1C
#617640000000
0!
0*
09
0>
0C
#617650000000
1!
1*
19
1>
1C
#617660000000
0!
0*
09
0>
0C
#617670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#617680000000
0!
0*
09
0>
0C
#617690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#617700000000
0!
0*
09
0>
0C
#617710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#617720000000
0!
0*
09
0>
0C
#617730000000
1!
1*
b10 6
19
1>
1C
b10 G
#617740000000
0!
0*
09
0>
0C
#617750000000
1!
1*
b11 6
19
1>
1C
b11 G
#617760000000
0!
0*
09
0>
0C
#617770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#617780000000
0!
0*
09
0>
0C
#617790000000
1!
1*
b101 6
19
1>
1C
b101 G
#617800000000
0!
0*
09
0>
0C
#617810000000
1!
1*
b110 6
19
1>
1C
b110 G
#617820000000
0!
0*
09
0>
0C
#617830000000
1!
1*
b111 6
19
1>
1C
b111 G
#617840000000
0!
0*
09
0>
0C
#617850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#617860000000
0!
0*
09
0>
0C
#617870000000
1!
1*
b1 6
19
1>
1C
b1 G
#617880000000
0!
0*
09
0>
0C
#617890000000
1!
1*
b10 6
19
1>
1C
b10 G
#617900000000
0!
0*
09
0>
0C
#617910000000
1!
1*
b11 6
19
1>
1C
b11 G
#617920000000
0!
0*
09
0>
0C
#617930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#617940000000
0!
0*
09
0>
0C
#617950000000
1!
1*
b101 6
19
1>
1C
b101 G
#617960000000
0!
0*
09
0>
0C
#617970000000
1!
1*
b110 6
19
1>
1C
b110 G
#617980000000
0!
0*
09
0>
0C
#617990000000
1!
1*
b111 6
19
1>
1C
b111 G
#618000000000
0!
0*
09
0>
0C
#618010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#618020000000
0!
0*
09
0>
0C
#618030000000
1!
1*
b1 6
19
1>
1C
b1 G
#618040000000
0!
0*
09
0>
0C
#618050000000
1!
1*
b10 6
19
1>
1C
b10 G
#618060000000
0!
0*
09
0>
0C
#618070000000
1!
1*
b11 6
19
1>
1C
b11 G
#618080000000
0!
0*
09
0>
0C
#618090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#618100000000
0!
0*
09
0>
0C
#618110000000
1!
1*
b101 6
19
1>
1C
b101 G
#618120000000
0!
0*
09
0>
0C
#618130000000
1!
1*
b110 6
19
1>
1C
b110 G
#618140000000
0!
0*
09
0>
0C
#618150000000
1!
1*
b111 6
19
1>
1C
b111 G
#618160000000
0!
1"
0*
1+
09
1:
0>
0C
#618170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#618180000000
0!
0*
09
0>
0C
#618190000000
1!
1*
b1 6
19
1>
1C
b1 G
#618200000000
0!
0*
09
0>
0C
#618210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#618220000000
0!
0*
09
0>
0C
#618230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#618240000000
0!
0*
09
0>
0C
#618250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#618260000000
0!
0*
09
0>
0C
#618270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#618280000000
0!
0#
0*
0,
09
0>
0?
0C
#618290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#618300000000
0!
0*
09
0>
0C
#618310000000
1!
1*
19
1>
1C
#618320000000
0!
0*
09
0>
0C
#618330000000
1!
1*
19
1>
1C
#618340000000
0!
0*
09
0>
0C
#618350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#618360000000
0!
0*
09
0>
0C
#618370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#618380000000
0!
0*
09
0>
0C
#618390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#618400000000
0!
0*
09
0>
0C
#618410000000
1!
1*
b10 6
19
1>
1C
b10 G
#618420000000
0!
0*
09
0>
0C
#618430000000
1!
1*
b11 6
19
1>
1C
b11 G
#618440000000
0!
0*
09
0>
0C
#618450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#618460000000
0!
0*
09
0>
0C
#618470000000
1!
1*
b101 6
19
1>
1C
b101 G
#618480000000
0!
0*
09
0>
0C
#618490000000
1!
1*
b110 6
19
1>
1C
b110 G
#618500000000
0!
0*
09
0>
0C
#618510000000
1!
1*
b111 6
19
1>
1C
b111 G
#618520000000
0!
0*
09
0>
0C
#618530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#618540000000
0!
0*
09
0>
0C
#618550000000
1!
1*
b1 6
19
1>
1C
b1 G
#618560000000
0!
0*
09
0>
0C
#618570000000
1!
1*
b10 6
19
1>
1C
b10 G
#618580000000
0!
0*
09
0>
0C
#618590000000
1!
1*
b11 6
19
1>
1C
b11 G
#618600000000
0!
0*
09
0>
0C
#618610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#618620000000
0!
0*
09
0>
0C
#618630000000
1!
1*
b101 6
19
1>
1C
b101 G
#618640000000
0!
0*
09
0>
0C
#618650000000
1!
1*
b110 6
19
1>
1C
b110 G
#618660000000
0!
0*
09
0>
0C
#618670000000
1!
1*
b111 6
19
1>
1C
b111 G
#618680000000
0!
0*
09
0>
0C
#618690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#618700000000
0!
0*
09
0>
0C
#618710000000
1!
1*
b1 6
19
1>
1C
b1 G
#618720000000
0!
0*
09
0>
0C
#618730000000
1!
1*
b10 6
19
1>
1C
b10 G
#618740000000
0!
0*
09
0>
0C
#618750000000
1!
1*
b11 6
19
1>
1C
b11 G
#618760000000
0!
0*
09
0>
0C
#618770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#618780000000
0!
0*
09
0>
0C
#618790000000
1!
1*
b101 6
19
1>
1C
b101 G
#618800000000
0!
0*
09
0>
0C
#618810000000
1!
1*
b110 6
19
1>
1C
b110 G
#618820000000
0!
0*
09
0>
0C
#618830000000
1!
1*
b111 6
19
1>
1C
b111 G
#618840000000
0!
1"
0*
1+
09
1:
0>
0C
#618850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#618860000000
0!
0*
09
0>
0C
#618870000000
1!
1*
b1 6
19
1>
1C
b1 G
#618880000000
0!
0*
09
0>
0C
#618890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#618900000000
0!
0*
09
0>
0C
#618910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#618920000000
0!
0*
09
0>
0C
#618930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#618940000000
0!
0*
09
0>
0C
#618950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#618960000000
0!
0#
0*
0,
09
0>
0?
0C
#618970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#618980000000
0!
0*
09
0>
0C
#618990000000
1!
1*
19
1>
1C
#619000000000
0!
0*
09
0>
0C
#619010000000
1!
1*
19
1>
1C
#619020000000
0!
0*
09
0>
0C
#619030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#619040000000
0!
0*
09
0>
0C
#619050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#619060000000
0!
0*
09
0>
0C
#619070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#619080000000
0!
0*
09
0>
0C
#619090000000
1!
1*
b10 6
19
1>
1C
b10 G
#619100000000
0!
0*
09
0>
0C
#619110000000
1!
1*
b11 6
19
1>
1C
b11 G
#619120000000
0!
0*
09
0>
0C
#619130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#619140000000
0!
0*
09
0>
0C
#619150000000
1!
1*
b101 6
19
1>
1C
b101 G
#619160000000
0!
0*
09
0>
0C
#619170000000
1!
1*
b110 6
19
1>
1C
b110 G
#619180000000
0!
0*
09
0>
0C
#619190000000
1!
1*
b111 6
19
1>
1C
b111 G
#619200000000
0!
0*
09
0>
0C
#619210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#619220000000
0!
0*
09
0>
0C
#619230000000
1!
1*
b1 6
19
1>
1C
b1 G
#619240000000
0!
0*
09
0>
0C
#619250000000
1!
1*
b10 6
19
1>
1C
b10 G
#619260000000
0!
0*
09
0>
0C
#619270000000
1!
1*
b11 6
19
1>
1C
b11 G
#619280000000
0!
0*
09
0>
0C
#619290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#619300000000
0!
0*
09
0>
0C
#619310000000
1!
1*
b101 6
19
1>
1C
b101 G
#619320000000
0!
0*
09
0>
0C
#619330000000
1!
1*
b110 6
19
1>
1C
b110 G
#619340000000
0!
0*
09
0>
0C
#619350000000
1!
1*
b111 6
19
1>
1C
b111 G
#619360000000
0!
0*
09
0>
0C
#619370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#619380000000
0!
0*
09
0>
0C
#619390000000
1!
1*
b1 6
19
1>
1C
b1 G
#619400000000
0!
0*
09
0>
0C
#619410000000
1!
1*
b10 6
19
1>
1C
b10 G
#619420000000
0!
0*
09
0>
0C
#619430000000
1!
1*
b11 6
19
1>
1C
b11 G
#619440000000
0!
0*
09
0>
0C
#619450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#619460000000
0!
0*
09
0>
0C
#619470000000
1!
1*
b101 6
19
1>
1C
b101 G
#619480000000
0!
0*
09
0>
0C
#619490000000
1!
1*
b110 6
19
1>
1C
b110 G
#619500000000
0!
0*
09
0>
0C
#619510000000
1!
1*
b111 6
19
1>
1C
b111 G
#619520000000
0!
1"
0*
1+
09
1:
0>
0C
#619530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#619540000000
0!
0*
09
0>
0C
#619550000000
1!
1*
b1 6
19
1>
1C
b1 G
#619560000000
0!
0*
09
0>
0C
#619570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#619580000000
0!
0*
09
0>
0C
#619590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#619600000000
0!
0*
09
0>
0C
#619610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#619620000000
0!
0*
09
0>
0C
#619630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#619640000000
0!
0#
0*
0,
09
0>
0?
0C
#619650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#619660000000
0!
0*
09
0>
0C
#619670000000
1!
1*
19
1>
1C
#619680000000
0!
0*
09
0>
0C
#619690000000
1!
1*
19
1>
1C
#619700000000
0!
0*
09
0>
0C
#619710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#619720000000
0!
0*
09
0>
0C
#619730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#619740000000
0!
0*
09
0>
0C
#619750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#619760000000
0!
0*
09
0>
0C
#619770000000
1!
1*
b10 6
19
1>
1C
b10 G
#619780000000
0!
0*
09
0>
0C
#619790000000
1!
1*
b11 6
19
1>
1C
b11 G
#619800000000
0!
0*
09
0>
0C
#619810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#619820000000
0!
0*
09
0>
0C
#619830000000
1!
1*
b101 6
19
1>
1C
b101 G
#619840000000
0!
0*
09
0>
0C
#619850000000
1!
1*
b110 6
19
1>
1C
b110 G
#619860000000
0!
0*
09
0>
0C
#619870000000
1!
1*
b111 6
19
1>
1C
b111 G
#619880000000
0!
0*
09
0>
0C
#619890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#619900000000
0!
0*
09
0>
0C
#619910000000
1!
1*
b1 6
19
1>
1C
b1 G
#619920000000
0!
0*
09
0>
0C
#619930000000
1!
1*
b10 6
19
1>
1C
b10 G
#619940000000
0!
0*
09
0>
0C
#619950000000
1!
1*
b11 6
19
1>
1C
b11 G
#619960000000
0!
0*
09
0>
0C
#619970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#619980000000
0!
0*
09
0>
0C
#619990000000
1!
1*
b101 6
19
1>
1C
b101 G
#620000000000
0!
0*
09
0>
0C
#620010000000
1!
1*
b110 6
19
1>
1C
b110 G
#620020000000
0!
0*
09
0>
0C
#620030000000
1!
1*
b111 6
19
1>
1C
b111 G
#620040000000
0!
0*
09
0>
0C
#620050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#620060000000
0!
0*
09
0>
0C
#620070000000
1!
1*
b1 6
19
1>
1C
b1 G
#620080000000
0!
0*
09
0>
0C
#620090000000
1!
1*
b10 6
19
1>
1C
b10 G
#620100000000
0!
0*
09
0>
0C
#620110000000
1!
1*
b11 6
19
1>
1C
b11 G
#620120000000
0!
0*
09
0>
0C
#620130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#620140000000
0!
0*
09
0>
0C
#620150000000
1!
1*
b101 6
19
1>
1C
b101 G
#620160000000
0!
0*
09
0>
0C
#620170000000
1!
1*
b110 6
19
1>
1C
b110 G
#620180000000
0!
0*
09
0>
0C
#620190000000
1!
1*
b111 6
19
1>
1C
b111 G
#620200000000
0!
1"
0*
1+
09
1:
0>
0C
#620210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#620220000000
0!
0*
09
0>
0C
#620230000000
1!
1*
b1 6
19
1>
1C
b1 G
#620240000000
0!
0*
09
0>
0C
#620250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#620260000000
0!
0*
09
0>
0C
#620270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#620280000000
0!
0*
09
0>
0C
#620290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#620300000000
0!
0*
09
0>
0C
#620310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#620320000000
0!
0#
0*
0,
09
0>
0?
0C
#620330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#620340000000
0!
0*
09
0>
0C
#620350000000
1!
1*
19
1>
1C
#620360000000
0!
0*
09
0>
0C
#620370000000
1!
1*
19
1>
1C
#620380000000
0!
0*
09
0>
0C
#620390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#620400000000
0!
0*
09
0>
0C
#620410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#620420000000
0!
0*
09
0>
0C
#620430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#620440000000
0!
0*
09
0>
0C
#620450000000
1!
1*
b10 6
19
1>
1C
b10 G
#620460000000
0!
0*
09
0>
0C
#620470000000
1!
1*
b11 6
19
1>
1C
b11 G
#620480000000
0!
0*
09
0>
0C
#620490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#620500000000
0!
0*
09
0>
0C
#620510000000
1!
1*
b101 6
19
1>
1C
b101 G
#620520000000
0!
0*
09
0>
0C
#620530000000
1!
1*
b110 6
19
1>
1C
b110 G
#620540000000
0!
0*
09
0>
0C
#620550000000
1!
1*
b111 6
19
1>
1C
b111 G
#620560000000
0!
0*
09
0>
0C
#620570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#620580000000
0!
0*
09
0>
0C
#620590000000
1!
1*
b1 6
19
1>
1C
b1 G
#620600000000
0!
0*
09
0>
0C
#620610000000
1!
1*
b10 6
19
1>
1C
b10 G
#620620000000
0!
0*
09
0>
0C
#620630000000
1!
1*
b11 6
19
1>
1C
b11 G
#620640000000
0!
0*
09
0>
0C
#620650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#620660000000
0!
0*
09
0>
0C
#620670000000
1!
1*
b101 6
19
1>
1C
b101 G
#620680000000
0!
0*
09
0>
0C
#620690000000
1!
1*
b110 6
19
1>
1C
b110 G
#620700000000
0!
0*
09
0>
0C
#620710000000
1!
1*
b111 6
19
1>
1C
b111 G
#620720000000
0!
0*
09
0>
0C
#620730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#620740000000
0!
0*
09
0>
0C
#620750000000
1!
1*
b1 6
19
1>
1C
b1 G
#620760000000
0!
0*
09
0>
0C
#620770000000
1!
1*
b10 6
19
1>
1C
b10 G
#620780000000
0!
0*
09
0>
0C
#620790000000
1!
1*
b11 6
19
1>
1C
b11 G
#620800000000
0!
0*
09
0>
0C
#620810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#620820000000
0!
0*
09
0>
0C
#620830000000
1!
1*
b101 6
19
1>
1C
b101 G
#620840000000
0!
0*
09
0>
0C
#620850000000
1!
1*
b110 6
19
1>
1C
b110 G
#620860000000
0!
0*
09
0>
0C
#620870000000
1!
1*
b111 6
19
1>
1C
b111 G
#620880000000
0!
1"
0*
1+
09
1:
0>
0C
#620890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#620900000000
0!
0*
09
0>
0C
#620910000000
1!
1*
b1 6
19
1>
1C
b1 G
#620920000000
0!
0*
09
0>
0C
#620930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#620940000000
0!
0*
09
0>
0C
#620950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#620960000000
0!
0*
09
0>
0C
#620970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#620980000000
0!
0*
09
0>
0C
#620990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#621000000000
0!
0#
0*
0,
09
0>
0?
0C
#621010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#621020000000
0!
0*
09
0>
0C
#621030000000
1!
1*
19
1>
1C
#621040000000
0!
0*
09
0>
0C
#621050000000
1!
1*
19
1>
1C
#621060000000
0!
0*
09
0>
0C
#621070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#621080000000
0!
0*
09
0>
0C
#621090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#621100000000
0!
0*
09
0>
0C
#621110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#621120000000
0!
0*
09
0>
0C
#621130000000
1!
1*
b10 6
19
1>
1C
b10 G
#621140000000
0!
0*
09
0>
0C
#621150000000
1!
1*
b11 6
19
1>
1C
b11 G
#621160000000
0!
0*
09
0>
0C
#621170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#621180000000
0!
0*
09
0>
0C
#621190000000
1!
1*
b101 6
19
1>
1C
b101 G
#621200000000
0!
0*
09
0>
0C
#621210000000
1!
1*
b110 6
19
1>
1C
b110 G
#621220000000
0!
0*
09
0>
0C
#621230000000
1!
1*
b111 6
19
1>
1C
b111 G
#621240000000
0!
0*
09
0>
0C
#621250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#621260000000
0!
0*
09
0>
0C
#621270000000
1!
1*
b1 6
19
1>
1C
b1 G
#621280000000
0!
0*
09
0>
0C
#621290000000
1!
1*
b10 6
19
1>
1C
b10 G
#621300000000
0!
0*
09
0>
0C
#621310000000
1!
1*
b11 6
19
1>
1C
b11 G
#621320000000
0!
0*
09
0>
0C
#621330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#621340000000
0!
0*
09
0>
0C
#621350000000
1!
1*
b101 6
19
1>
1C
b101 G
#621360000000
0!
0*
09
0>
0C
#621370000000
1!
1*
b110 6
19
1>
1C
b110 G
#621380000000
0!
0*
09
0>
0C
#621390000000
1!
1*
b111 6
19
1>
1C
b111 G
#621400000000
0!
0*
09
0>
0C
#621410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#621420000000
0!
0*
09
0>
0C
#621430000000
1!
1*
b1 6
19
1>
1C
b1 G
#621440000000
0!
0*
09
0>
0C
#621450000000
1!
1*
b10 6
19
1>
1C
b10 G
#621460000000
0!
0*
09
0>
0C
#621470000000
1!
1*
b11 6
19
1>
1C
b11 G
#621480000000
0!
0*
09
0>
0C
#621490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#621500000000
0!
0*
09
0>
0C
#621510000000
1!
1*
b101 6
19
1>
1C
b101 G
#621520000000
0!
0*
09
0>
0C
#621530000000
1!
1*
b110 6
19
1>
1C
b110 G
#621540000000
0!
0*
09
0>
0C
#621550000000
1!
1*
b111 6
19
1>
1C
b111 G
#621560000000
0!
1"
0*
1+
09
1:
0>
0C
#621570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#621580000000
0!
0*
09
0>
0C
#621590000000
1!
1*
b1 6
19
1>
1C
b1 G
#621600000000
0!
0*
09
0>
0C
#621610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#621620000000
0!
0*
09
0>
0C
#621630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#621640000000
0!
0*
09
0>
0C
#621650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#621660000000
0!
0*
09
0>
0C
#621670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#621680000000
0!
0#
0*
0,
09
0>
0?
0C
#621690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#621700000000
0!
0*
09
0>
0C
#621710000000
1!
1*
19
1>
1C
#621720000000
0!
0*
09
0>
0C
#621730000000
1!
1*
19
1>
1C
#621740000000
0!
0*
09
0>
0C
#621750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#621760000000
0!
0*
09
0>
0C
#621770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#621780000000
0!
0*
09
0>
0C
#621790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#621800000000
0!
0*
09
0>
0C
#621810000000
1!
1*
b10 6
19
1>
1C
b10 G
#621820000000
0!
0*
09
0>
0C
#621830000000
1!
1*
b11 6
19
1>
1C
b11 G
#621840000000
0!
0*
09
0>
0C
#621850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#621860000000
0!
0*
09
0>
0C
#621870000000
1!
1*
b101 6
19
1>
1C
b101 G
#621880000000
0!
0*
09
0>
0C
#621890000000
1!
1*
b110 6
19
1>
1C
b110 G
#621900000000
0!
0*
09
0>
0C
#621910000000
1!
1*
b111 6
19
1>
1C
b111 G
#621920000000
0!
0*
09
0>
0C
#621930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#621940000000
0!
0*
09
0>
0C
#621950000000
1!
1*
b1 6
19
1>
1C
b1 G
#621960000000
0!
0*
09
0>
0C
#621970000000
1!
1*
b10 6
19
1>
1C
b10 G
#621980000000
0!
0*
09
0>
0C
#621990000000
1!
1*
b11 6
19
1>
1C
b11 G
#622000000000
0!
0*
09
0>
0C
#622010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#622020000000
0!
0*
09
0>
0C
#622030000000
1!
1*
b101 6
19
1>
1C
b101 G
#622040000000
0!
0*
09
0>
0C
#622050000000
1!
1*
b110 6
19
1>
1C
b110 G
#622060000000
0!
0*
09
0>
0C
#622070000000
1!
1*
b111 6
19
1>
1C
b111 G
#622080000000
0!
0*
09
0>
0C
#622090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#622100000000
0!
0*
09
0>
0C
#622110000000
1!
1*
b1 6
19
1>
1C
b1 G
#622120000000
0!
0*
09
0>
0C
#622130000000
1!
1*
b10 6
19
1>
1C
b10 G
#622140000000
0!
0*
09
0>
0C
#622150000000
1!
1*
b11 6
19
1>
1C
b11 G
#622160000000
0!
0*
09
0>
0C
#622170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#622180000000
0!
0*
09
0>
0C
#622190000000
1!
1*
b101 6
19
1>
1C
b101 G
#622200000000
0!
0*
09
0>
0C
#622210000000
1!
1*
b110 6
19
1>
1C
b110 G
#622220000000
0!
0*
09
0>
0C
#622230000000
1!
1*
b111 6
19
1>
1C
b111 G
#622240000000
0!
1"
0*
1+
09
1:
0>
0C
#622250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#622260000000
0!
0*
09
0>
0C
#622270000000
1!
1*
b1 6
19
1>
1C
b1 G
#622280000000
0!
0*
09
0>
0C
#622290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#622300000000
0!
0*
09
0>
0C
#622310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#622320000000
0!
0*
09
0>
0C
#622330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#622340000000
0!
0*
09
0>
0C
#622350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#622360000000
0!
0#
0*
0,
09
0>
0?
0C
#622370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#622380000000
0!
0*
09
0>
0C
#622390000000
1!
1*
19
1>
1C
#622400000000
0!
0*
09
0>
0C
#622410000000
1!
1*
19
1>
1C
#622420000000
0!
0*
09
0>
0C
#622430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#622440000000
0!
0*
09
0>
0C
#622450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#622460000000
0!
0*
09
0>
0C
#622470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#622480000000
0!
0*
09
0>
0C
#622490000000
1!
1*
b10 6
19
1>
1C
b10 G
#622500000000
0!
0*
09
0>
0C
#622510000000
1!
1*
b11 6
19
1>
1C
b11 G
#622520000000
0!
0*
09
0>
0C
#622530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#622540000000
0!
0*
09
0>
0C
#622550000000
1!
1*
b101 6
19
1>
1C
b101 G
#622560000000
0!
0*
09
0>
0C
#622570000000
1!
1*
b110 6
19
1>
1C
b110 G
#622580000000
0!
0*
09
0>
0C
#622590000000
1!
1*
b111 6
19
1>
1C
b111 G
#622600000000
0!
0*
09
0>
0C
#622610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#622620000000
0!
0*
09
0>
0C
#622630000000
1!
1*
b1 6
19
1>
1C
b1 G
#622640000000
0!
0*
09
0>
0C
#622650000000
1!
1*
b10 6
19
1>
1C
b10 G
#622660000000
0!
0*
09
0>
0C
#622670000000
1!
1*
b11 6
19
1>
1C
b11 G
#622680000000
0!
0*
09
0>
0C
#622690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#622700000000
0!
0*
09
0>
0C
#622710000000
1!
1*
b101 6
19
1>
1C
b101 G
#622720000000
0!
0*
09
0>
0C
#622730000000
1!
1*
b110 6
19
1>
1C
b110 G
#622740000000
0!
0*
09
0>
0C
#622750000000
1!
1*
b111 6
19
1>
1C
b111 G
#622760000000
0!
0*
09
0>
0C
#622770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#622780000000
0!
0*
09
0>
0C
#622790000000
1!
1*
b1 6
19
1>
1C
b1 G
#622800000000
0!
0*
09
0>
0C
#622810000000
1!
1*
b10 6
19
1>
1C
b10 G
#622820000000
0!
0*
09
0>
0C
#622830000000
1!
1*
b11 6
19
1>
1C
b11 G
#622840000000
0!
0*
09
0>
0C
#622850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#622860000000
0!
0*
09
0>
0C
#622870000000
1!
1*
b101 6
19
1>
1C
b101 G
#622880000000
0!
0*
09
0>
0C
#622890000000
1!
1*
b110 6
19
1>
1C
b110 G
#622900000000
0!
0*
09
0>
0C
#622910000000
1!
1*
b111 6
19
1>
1C
b111 G
#622920000000
0!
1"
0*
1+
09
1:
0>
0C
#622930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#622940000000
0!
0*
09
0>
0C
#622950000000
1!
1*
b1 6
19
1>
1C
b1 G
#622960000000
0!
0*
09
0>
0C
#622970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#622980000000
0!
0*
09
0>
0C
#622990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#623000000000
0!
0*
09
0>
0C
#623010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#623020000000
0!
0*
09
0>
0C
#623030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#623040000000
0!
0#
0*
0,
09
0>
0?
0C
#623050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#623060000000
0!
0*
09
0>
0C
#623070000000
1!
1*
19
1>
1C
#623080000000
0!
0*
09
0>
0C
#623090000000
1!
1*
19
1>
1C
#623100000000
0!
0*
09
0>
0C
#623110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#623120000000
0!
0*
09
0>
0C
#623130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#623140000000
0!
0*
09
0>
0C
#623150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#623160000000
0!
0*
09
0>
0C
#623170000000
1!
1*
b10 6
19
1>
1C
b10 G
#623180000000
0!
0*
09
0>
0C
#623190000000
1!
1*
b11 6
19
1>
1C
b11 G
#623200000000
0!
0*
09
0>
0C
#623210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#623220000000
0!
0*
09
0>
0C
#623230000000
1!
1*
b101 6
19
1>
1C
b101 G
#623240000000
0!
0*
09
0>
0C
#623250000000
1!
1*
b110 6
19
1>
1C
b110 G
#623260000000
0!
0*
09
0>
0C
#623270000000
1!
1*
b111 6
19
1>
1C
b111 G
#623280000000
0!
0*
09
0>
0C
#623290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#623300000000
0!
0*
09
0>
0C
#623310000000
1!
1*
b1 6
19
1>
1C
b1 G
#623320000000
0!
0*
09
0>
0C
#623330000000
1!
1*
b10 6
19
1>
1C
b10 G
#623340000000
0!
0*
09
0>
0C
#623350000000
1!
1*
b11 6
19
1>
1C
b11 G
#623360000000
0!
0*
09
0>
0C
#623370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#623380000000
0!
0*
09
0>
0C
#623390000000
1!
1*
b101 6
19
1>
1C
b101 G
#623400000000
0!
0*
09
0>
0C
#623410000000
1!
1*
b110 6
19
1>
1C
b110 G
#623420000000
0!
0*
09
0>
0C
#623430000000
1!
1*
b111 6
19
1>
1C
b111 G
#623440000000
0!
0*
09
0>
0C
#623450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#623460000000
0!
0*
09
0>
0C
#623470000000
1!
1*
b1 6
19
1>
1C
b1 G
#623480000000
0!
0*
09
0>
0C
#623490000000
1!
1*
b10 6
19
1>
1C
b10 G
#623500000000
0!
0*
09
0>
0C
#623510000000
1!
1*
b11 6
19
1>
1C
b11 G
#623520000000
0!
0*
09
0>
0C
#623530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#623540000000
0!
0*
09
0>
0C
#623550000000
1!
1*
b101 6
19
1>
1C
b101 G
#623560000000
0!
0*
09
0>
0C
#623570000000
1!
1*
b110 6
19
1>
1C
b110 G
#623580000000
0!
0*
09
0>
0C
#623590000000
1!
1*
b111 6
19
1>
1C
b111 G
#623600000000
0!
1"
0*
1+
09
1:
0>
0C
#623610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#623620000000
0!
0*
09
0>
0C
#623630000000
1!
1*
b1 6
19
1>
1C
b1 G
#623640000000
0!
0*
09
0>
0C
#623650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#623660000000
0!
0*
09
0>
0C
#623670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#623680000000
0!
0*
09
0>
0C
#623690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#623700000000
0!
0*
09
0>
0C
#623710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#623720000000
0!
0#
0*
0,
09
0>
0?
0C
#623730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#623740000000
0!
0*
09
0>
0C
#623750000000
1!
1*
19
1>
1C
#623760000000
0!
0*
09
0>
0C
#623770000000
1!
1*
19
1>
1C
#623780000000
0!
0*
09
0>
0C
#623790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#623800000000
0!
0*
09
0>
0C
#623810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#623820000000
0!
0*
09
0>
0C
#623830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#623840000000
0!
0*
09
0>
0C
#623850000000
1!
1*
b10 6
19
1>
1C
b10 G
#623860000000
0!
0*
09
0>
0C
#623870000000
1!
1*
b11 6
19
1>
1C
b11 G
#623880000000
0!
0*
09
0>
0C
#623890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#623900000000
0!
0*
09
0>
0C
#623910000000
1!
1*
b101 6
19
1>
1C
b101 G
#623920000000
0!
0*
09
0>
0C
#623930000000
1!
1*
b110 6
19
1>
1C
b110 G
#623940000000
0!
0*
09
0>
0C
#623950000000
1!
1*
b111 6
19
1>
1C
b111 G
#623960000000
0!
0*
09
0>
0C
#623970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#623980000000
0!
0*
09
0>
0C
#623990000000
1!
1*
b1 6
19
1>
1C
b1 G
#624000000000
0!
0*
09
0>
0C
#624010000000
1!
1*
b10 6
19
1>
1C
b10 G
#624020000000
0!
0*
09
0>
0C
#624030000000
1!
1*
b11 6
19
1>
1C
b11 G
#624040000000
0!
0*
09
0>
0C
#624050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#624060000000
0!
0*
09
0>
0C
#624070000000
1!
1*
b101 6
19
1>
1C
b101 G
#624080000000
0!
0*
09
0>
0C
#624090000000
1!
1*
b110 6
19
1>
1C
b110 G
#624100000000
0!
0*
09
0>
0C
#624110000000
1!
1*
b111 6
19
1>
1C
b111 G
#624120000000
0!
0*
09
0>
0C
#624130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#624140000000
0!
0*
09
0>
0C
#624150000000
1!
1*
b1 6
19
1>
1C
b1 G
#624160000000
0!
0*
09
0>
0C
#624170000000
1!
1*
b10 6
19
1>
1C
b10 G
#624180000000
0!
0*
09
0>
0C
#624190000000
1!
1*
b11 6
19
1>
1C
b11 G
#624200000000
0!
0*
09
0>
0C
#624210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#624220000000
0!
0*
09
0>
0C
#624230000000
1!
1*
b101 6
19
1>
1C
b101 G
#624240000000
0!
0*
09
0>
0C
#624250000000
1!
1*
b110 6
19
1>
1C
b110 G
#624260000000
0!
0*
09
0>
0C
#624270000000
1!
1*
b111 6
19
1>
1C
b111 G
#624280000000
0!
1"
0*
1+
09
1:
0>
0C
#624290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#624300000000
0!
0*
09
0>
0C
#624310000000
1!
1*
b1 6
19
1>
1C
b1 G
#624320000000
0!
0*
09
0>
0C
#624330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#624340000000
0!
0*
09
0>
0C
#624350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#624360000000
0!
0*
09
0>
0C
#624370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#624380000000
0!
0*
09
0>
0C
#624390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#624400000000
0!
0#
0*
0,
09
0>
0?
0C
#624410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#624420000000
0!
0*
09
0>
0C
#624430000000
1!
1*
19
1>
1C
#624440000000
0!
0*
09
0>
0C
#624450000000
1!
1*
19
1>
1C
#624460000000
0!
0*
09
0>
0C
#624470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#624480000000
0!
0*
09
0>
0C
#624490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#624500000000
0!
0*
09
0>
0C
#624510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#624520000000
0!
0*
09
0>
0C
#624530000000
1!
1*
b10 6
19
1>
1C
b10 G
#624540000000
0!
0*
09
0>
0C
#624550000000
1!
1*
b11 6
19
1>
1C
b11 G
#624560000000
0!
0*
09
0>
0C
#624570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#624580000000
0!
0*
09
0>
0C
#624590000000
1!
1*
b101 6
19
1>
1C
b101 G
#624600000000
0!
0*
09
0>
0C
#624610000000
1!
1*
b110 6
19
1>
1C
b110 G
#624620000000
0!
0*
09
0>
0C
#624630000000
1!
1*
b111 6
19
1>
1C
b111 G
#624640000000
0!
0*
09
0>
0C
#624650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#624660000000
0!
0*
09
0>
0C
#624670000000
1!
1*
b1 6
19
1>
1C
b1 G
#624680000000
0!
0*
09
0>
0C
#624690000000
1!
1*
b10 6
19
1>
1C
b10 G
#624700000000
0!
0*
09
0>
0C
#624710000000
1!
1*
b11 6
19
1>
1C
b11 G
#624720000000
0!
0*
09
0>
0C
#624730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#624740000000
0!
0*
09
0>
0C
#624750000000
1!
1*
b101 6
19
1>
1C
b101 G
#624760000000
0!
0*
09
0>
0C
#624770000000
1!
1*
b110 6
19
1>
1C
b110 G
#624780000000
0!
0*
09
0>
0C
#624790000000
1!
1*
b111 6
19
1>
1C
b111 G
#624800000000
0!
0*
09
0>
0C
#624810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#624820000000
0!
0*
09
0>
0C
#624830000000
1!
1*
b1 6
19
1>
1C
b1 G
#624840000000
0!
0*
09
0>
0C
#624850000000
1!
1*
b10 6
19
1>
1C
b10 G
#624860000000
0!
0*
09
0>
0C
#624870000000
1!
1*
b11 6
19
1>
1C
b11 G
#624880000000
0!
0*
09
0>
0C
#624890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#624900000000
0!
0*
09
0>
0C
#624910000000
1!
1*
b101 6
19
1>
1C
b101 G
#624920000000
0!
0*
09
0>
0C
#624930000000
1!
1*
b110 6
19
1>
1C
b110 G
#624940000000
0!
0*
09
0>
0C
#624950000000
1!
1*
b111 6
19
1>
1C
b111 G
#624960000000
0!
1"
0*
1+
09
1:
0>
0C
#624970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#624980000000
0!
0*
09
0>
0C
#624990000000
1!
1*
b1 6
19
1>
1C
b1 G
#625000000000
0!
0*
09
0>
0C
#625010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#625020000000
0!
0*
09
0>
0C
#625030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#625040000000
0!
0*
09
0>
0C
#625050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#625060000000
0!
0*
09
0>
0C
#625070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#625080000000
0!
0#
0*
0,
09
0>
0?
0C
#625090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#625100000000
0!
0*
09
0>
0C
#625110000000
1!
1*
19
1>
1C
#625120000000
0!
0*
09
0>
0C
#625130000000
1!
1*
19
1>
1C
#625140000000
0!
0*
09
0>
0C
#625150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#625160000000
0!
0*
09
0>
0C
#625170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#625180000000
0!
0*
09
0>
0C
#625190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#625200000000
0!
0*
09
0>
0C
#625210000000
1!
1*
b10 6
19
1>
1C
b10 G
#625220000000
0!
0*
09
0>
0C
#625230000000
1!
1*
b11 6
19
1>
1C
b11 G
#625240000000
0!
0*
09
0>
0C
#625250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#625260000000
0!
0*
09
0>
0C
#625270000000
1!
1*
b101 6
19
1>
1C
b101 G
#625280000000
0!
0*
09
0>
0C
#625290000000
1!
1*
b110 6
19
1>
1C
b110 G
#625300000000
0!
0*
09
0>
0C
#625310000000
1!
1*
b111 6
19
1>
1C
b111 G
#625320000000
0!
0*
09
0>
0C
#625330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#625340000000
0!
0*
09
0>
0C
#625350000000
1!
1*
b1 6
19
1>
1C
b1 G
#625360000000
0!
0*
09
0>
0C
#625370000000
1!
1*
b10 6
19
1>
1C
b10 G
#625380000000
0!
0*
09
0>
0C
#625390000000
1!
1*
b11 6
19
1>
1C
b11 G
#625400000000
0!
0*
09
0>
0C
#625410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#625420000000
0!
0*
09
0>
0C
#625430000000
1!
1*
b101 6
19
1>
1C
b101 G
#625440000000
0!
0*
09
0>
0C
#625450000000
1!
1*
b110 6
19
1>
1C
b110 G
#625460000000
0!
0*
09
0>
0C
#625470000000
1!
1*
b111 6
19
1>
1C
b111 G
#625480000000
0!
0*
09
0>
0C
#625490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#625500000000
0!
0*
09
0>
0C
#625510000000
1!
1*
b1 6
19
1>
1C
b1 G
#625520000000
0!
0*
09
0>
0C
#625530000000
1!
1*
b10 6
19
1>
1C
b10 G
#625540000000
0!
0*
09
0>
0C
#625550000000
1!
1*
b11 6
19
1>
1C
b11 G
#625560000000
0!
0*
09
0>
0C
#625570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#625580000000
0!
0*
09
0>
0C
#625590000000
1!
1*
b101 6
19
1>
1C
b101 G
#625600000000
0!
0*
09
0>
0C
#625610000000
1!
1*
b110 6
19
1>
1C
b110 G
#625620000000
0!
0*
09
0>
0C
#625630000000
1!
1*
b111 6
19
1>
1C
b111 G
#625640000000
0!
1"
0*
1+
09
1:
0>
0C
#625650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#625660000000
0!
0*
09
0>
0C
#625670000000
1!
1*
b1 6
19
1>
1C
b1 G
#625680000000
0!
0*
09
0>
0C
#625690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#625700000000
0!
0*
09
0>
0C
#625710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#625720000000
0!
0*
09
0>
0C
#625730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#625740000000
0!
0*
09
0>
0C
#625750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#625760000000
0!
0#
0*
0,
09
0>
0?
0C
#625770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#625780000000
0!
0*
09
0>
0C
#625790000000
1!
1*
19
1>
1C
#625800000000
0!
0*
09
0>
0C
#625810000000
1!
1*
19
1>
1C
#625820000000
0!
0*
09
0>
0C
#625830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#625840000000
0!
0*
09
0>
0C
#625850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#625860000000
0!
0*
09
0>
0C
#625870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#625880000000
0!
0*
09
0>
0C
#625890000000
1!
1*
b10 6
19
1>
1C
b10 G
#625900000000
0!
0*
09
0>
0C
#625910000000
1!
1*
b11 6
19
1>
1C
b11 G
#625920000000
0!
0*
09
0>
0C
#625930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#625940000000
0!
0*
09
0>
0C
#625950000000
1!
1*
b101 6
19
1>
1C
b101 G
#625960000000
0!
0*
09
0>
0C
#625970000000
1!
1*
b110 6
19
1>
1C
b110 G
#625980000000
0!
0*
09
0>
0C
#625990000000
1!
1*
b111 6
19
1>
1C
b111 G
#626000000000
0!
0*
09
0>
0C
#626010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#626020000000
0!
0*
09
0>
0C
#626030000000
1!
1*
b1 6
19
1>
1C
b1 G
#626040000000
0!
0*
09
0>
0C
#626050000000
1!
1*
b10 6
19
1>
1C
b10 G
#626060000000
0!
0*
09
0>
0C
#626070000000
1!
1*
b11 6
19
1>
1C
b11 G
#626080000000
0!
0*
09
0>
0C
#626090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#626100000000
0!
0*
09
0>
0C
#626110000000
1!
1*
b101 6
19
1>
1C
b101 G
#626120000000
0!
0*
09
0>
0C
#626130000000
1!
1*
b110 6
19
1>
1C
b110 G
#626140000000
0!
0*
09
0>
0C
#626150000000
1!
1*
b111 6
19
1>
1C
b111 G
#626160000000
0!
0*
09
0>
0C
#626170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#626180000000
0!
0*
09
0>
0C
#626190000000
1!
1*
b1 6
19
1>
1C
b1 G
#626200000000
0!
0*
09
0>
0C
#626210000000
1!
1*
b10 6
19
1>
1C
b10 G
#626220000000
0!
0*
09
0>
0C
#626230000000
1!
1*
b11 6
19
1>
1C
b11 G
#626240000000
0!
0*
09
0>
0C
#626250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#626260000000
0!
0*
09
0>
0C
#626270000000
1!
1*
b101 6
19
1>
1C
b101 G
#626280000000
0!
0*
09
0>
0C
#626290000000
1!
1*
b110 6
19
1>
1C
b110 G
#626300000000
0!
0*
09
0>
0C
#626310000000
1!
1*
b111 6
19
1>
1C
b111 G
#626320000000
0!
1"
0*
1+
09
1:
0>
0C
#626330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#626340000000
0!
0*
09
0>
0C
#626350000000
1!
1*
b1 6
19
1>
1C
b1 G
#626360000000
0!
0*
09
0>
0C
#626370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#626380000000
0!
0*
09
0>
0C
#626390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#626400000000
0!
0*
09
0>
0C
#626410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#626420000000
0!
0*
09
0>
0C
#626430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#626440000000
0!
0#
0*
0,
09
0>
0?
0C
#626450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#626460000000
0!
0*
09
0>
0C
#626470000000
1!
1*
19
1>
1C
#626480000000
0!
0*
09
0>
0C
#626490000000
1!
1*
19
1>
1C
#626500000000
0!
0*
09
0>
0C
#626510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#626520000000
0!
0*
09
0>
0C
#626530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#626540000000
0!
0*
09
0>
0C
#626550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#626560000000
0!
0*
09
0>
0C
#626570000000
1!
1*
b10 6
19
1>
1C
b10 G
#626580000000
0!
0*
09
0>
0C
#626590000000
1!
1*
b11 6
19
1>
1C
b11 G
#626600000000
0!
0*
09
0>
0C
#626610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#626620000000
0!
0*
09
0>
0C
#626630000000
1!
1*
b101 6
19
1>
1C
b101 G
#626640000000
0!
0*
09
0>
0C
#626650000000
1!
1*
b110 6
19
1>
1C
b110 G
#626660000000
0!
0*
09
0>
0C
#626670000000
1!
1*
b111 6
19
1>
1C
b111 G
#626680000000
0!
0*
09
0>
0C
#626690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#626700000000
0!
0*
09
0>
0C
#626710000000
1!
1*
b1 6
19
1>
1C
b1 G
#626720000000
0!
0*
09
0>
0C
#626730000000
1!
1*
b10 6
19
1>
1C
b10 G
#626740000000
0!
0*
09
0>
0C
#626750000000
1!
1*
b11 6
19
1>
1C
b11 G
#626760000000
0!
0*
09
0>
0C
#626770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#626780000000
0!
0*
09
0>
0C
#626790000000
1!
1*
b101 6
19
1>
1C
b101 G
#626800000000
0!
0*
09
0>
0C
#626810000000
1!
1*
b110 6
19
1>
1C
b110 G
#626820000000
0!
0*
09
0>
0C
#626830000000
1!
1*
b111 6
19
1>
1C
b111 G
#626840000000
0!
0*
09
0>
0C
#626850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#626860000000
0!
0*
09
0>
0C
#626870000000
1!
1*
b1 6
19
1>
1C
b1 G
#626880000000
0!
0*
09
0>
0C
#626890000000
1!
1*
b10 6
19
1>
1C
b10 G
#626900000000
0!
0*
09
0>
0C
#626910000000
1!
1*
b11 6
19
1>
1C
b11 G
#626920000000
0!
0*
09
0>
0C
#626930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#626940000000
0!
0*
09
0>
0C
#626950000000
1!
1*
b101 6
19
1>
1C
b101 G
#626960000000
0!
0*
09
0>
0C
#626970000000
1!
1*
b110 6
19
1>
1C
b110 G
#626980000000
0!
0*
09
0>
0C
#626990000000
1!
1*
b111 6
19
1>
1C
b111 G
#627000000000
0!
1"
0*
1+
09
1:
0>
0C
#627010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#627020000000
0!
0*
09
0>
0C
#627030000000
1!
1*
b1 6
19
1>
1C
b1 G
#627040000000
0!
0*
09
0>
0C
#627050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#627060000000
0!
0*
09
0>
0C
#627070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#627080000000
0!
0*
09
0>
0C
#627090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#627100000000
0!
0*
09
0>
0C
#627110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#627120000000
0!
0#
0*
0,
09
0>
0?
0C
#627130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#627140000000
0!
0*
09
0>
0C
#627150000000
1!
1*
19
1>
1C
#627160000000
0!
0*
09
0>
0C
#627170000000
1!
1*
19
1>
1C
#627180000000
0!
0*
09
0>
0C
#627190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#627200000000
0!
0*
09
0>
0C
#627210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#627220000000
0!
0*
09
0>
0C
#627230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#627240000000
0!
0*
09
0>
0C
#627250000000
1!
1*
b10 6
19
1>
1C
b10 G
#627260000000
0!
0*
09
0>
0C
#627270000000
1!
1*
b11 6
19
1>
1C
b11 G
#627280000000
0!
0*
09
0>
0C
#627290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#627300000000
0!
0*
09
0>
0C
#627310000000
1!
1*
b101 6
19
1>
1C
b101 G
#627320000000
0!
0*
09
0>
0C
#627330000000
1!
1*
b110 6
19
1>
1C
b110 G
#627340000000
0!
0*
09
0>
0C
#627350000000
1!
1*
b111 6
19
1>
1C
b111 G
#627360000000
0!
0*
09
0>
0C
#627370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#627380000000
0!
0*
09
0>
0C
#627390000000
1!
1*
b1 6
19
1>
1C
b1 G
#627400000000
0!
0*
09
0>
0C
#627410000000
1!
1*
b10 6
19
1>
1C
b10 G
#627420000000
0!
0*
09
0>
0C
#627430000000
1!
1*
b11 6
19
1>
1C
b11 G
#627440000000
0!
0*
09
0>
0C
#627450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#627460000000
0!
0*
09
0>
0C
#627470000000
1!
1*
b101 6
19
1>
1C
b101 G
#627480000000
0!
0*
09
0>
0C
#627490000000
1!
1*
b110 6
19
1>
1C
b110 G
#627500000000
0!
0*
09
0>
0C
#627510000000
1!
1*
b111 6
19
1>
1C
b111 G
#627520000000
0!
0*
09
0>
0C
#627530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#627540000000
0!
0*
09
0>
0C
#627550000000
1!
1*
b1 6
19
1>
1C
b1 G
#627560000000
0!
0*
09
0>
0C
#627570000000
1!
1*
b10 6
19
1>
1C
b10 G
#627580000000
0!
0*
09
0>
0C
#627590000000
1!
1*
b11 6
19
1>
1C
b11 G
#627600000000
0!
0*
09
0>
0C
#627610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#627620000000
0!
0*
09
0>
0C
#627630000000
1!
1*
b101 6
19
1>
1C
b101 G
#627640000000
0!
0*
09
0>
0C
#627650000000
1!
1*
b110 6
19
1>
1C
b110 G
#627660000000
0!
0*
09
0>
0C
#627670000000
1!
1*
b111 6
19
1>
1C
b111 G
#627680000000
0!
1"
0*
1+
09
1:
0>
0C
#627690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#627700000000
0!
0*
09
0>
0C
#627710000000
1!
1*
b1 6
19
1>
1C
b1 G
#627720000000
0!
0*
09
0>
0C
#627730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#627740000000
0!
0*
09
0>
0C
#627750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#627760000000
0!
0*
09
0>
0C
#627770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#627780000000
0!
0*
09
0>
0C
#627790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#627800000000
0!
0#
0*
0,
09
0>
0?
0C
#627810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#627820000000
0!
0*
09
0>
0C
#627830000000
1!
1*
19
1>
1C
#627840000000
0!
0*
09
0>
0C
#627850000000
1!
1*
19
1>
1C
#627860000000
0!
0*
09
0>
0C
#627870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#627880000000
0!
0*
09
0>
0C
#627890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#627900000000
0!
0*
09
0>
0C
#627910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#627920000000
0!
0*
09
0>
0C
#627930000000
1!
1*
b10 6
19
1>
1C
b10 G
#627940000000
0!
0*
09
0>
0C
#627950000000
1!
1*
b11 6
19
1>
1C
b11 G
#627960000000
0!
0*
09
0>
0C
#627970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#627980000000
0!
0*
09
0>
0C
#627990000000
1!
1*
b101 6
19
1>
1C
b101 G
#628000000000
0!
0*
09
0>
0C
#628010000000
1!
1*
b110 6
19
1>
1C
b110 G
#628020000000
0!
0*
09
0>
0C
#628030000000
1!
1*
b111 6
19
1>
1C
b111 G
#628040000000
0!
0*
09
0>
0C
#628050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#628060000000
0!
0*
09
0>
0C
#628070000000
1!
1*
b1 6
19
1>
1C
b1 G
#628080000000
0!
0*
09
0>
0C
#628090000000
1!
1*
b10 6
19
1>
1C
b10 G
#628100000000
0!
0*
09
0>
0C
#628110000000
1!
1*
b11 6
19
1>
1C
b11 G
#628120000000
0!
0*
09
0>
0C
#628130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#628140000000
0!
0*
09
0>
0C
#628150000000
1!
1*
b101 6
19
1>
1C
b101 G
#628160000000
0!
0*
09
0>
0C
#628170000000
1!
1*
b110 6
19
1>
1C
b110 G
#628180000000
0!
0*
09
0>
0C
#628190000000
1!
1*
b111 6
19
1>
1C
b111 G
#628200000000
0!
0*
09
0>
0C
#628210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#628220000000
0!
0*
09
0>
0C
#628230000000
1!
1*
b1 6
19
1>
1C
b1 G
#628240000000
0!
0*
09
0>
0C
#628250000000
1!
1*
b10 6
19
1>
1C
b10 G
#628260000000
0!
0*
09
0>
0C
#628270000000
1!
1*
b11 6
19
1>
1C
b11 G
#628280000000
0!
0*
09
0>
0C
#628290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#628300000000
0!
0*
09
0>
0C
#628310000000
1!
1*
b101 6
19
1>
1C
b101 G
#628320000000
0!
0*
09
0>
0C
#628330000000
1!
1*
b110 6
19
1>
1C
b110 G
#628340000000
0!
0*
09
0>
0C
#628350000000
1!
1*
b111 6
19
1>
1C
b111 G
#628360000000
0!
1"
0*
1+
09
1:
0>
0C
#628370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#628380000000
0!
0*
09
0>
0C
#628390000000
1!
1*
b1 6
19
1>
1C
b1 G
#628400000000
0!
0*
09
0>
0C
#628410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#628420000000
0!
0*
09
0>
0C
#628430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#628440000000
0!
0*
09
0>
0C
#628450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#628460000000
0!
0*
09
0>
0C
#628470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#628480000000
0!
0#
0*
0,
09
0>
0?
0C
#628490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#628500000000
0!
0*
09
0>
0C
#628510000000
1!
1*
19
1>
1C
#628520000000
0!
0*
09
0>
0C
#628530000000
1!
1*
19
1>
1C
#628540000000
0!
0*
09
0>
0C
#628550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#628560000000
0!
0*
09
0>
0C
#628570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#628580000000
0!
0*
09
0>
0C
#628590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#628600000000
0!
0*
09
0>
0C
#628610000000
1!
1*
b10 6
19
1>
1C
b10 G
#628620000000
0!
0*
09
0>
0C
#628630000000
1!
1*
b11 6
19
1>
1C
b11 G
#628640000000
0!
0*
09
0>
0C
#628650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#628660000000
0!
0*
09
0>
0C
#628670000000
1!
1*
b101 6
19
1>
1C
b101 G
#628680000000
0!
0*
09
0>
0C
#628690000000
1!
1*
b110 6
19
1>
1C
b110 G
#628700000000
0!
0*
09
0>
0C
#628710000000
1!
1*
b111 6
19
1>
1C
b111 G
#628720000000
0!
0*
09
0>
0C
#628730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#628740000000
0!
0*
09
0>
0C
#628750000000
1!
1*
b1 6
19
1>
1C
b1 G
#628760000000
0!
0*
09
0>
0C
#628770000000
1!
1*
b10 6
19
1>
1C
b10 G
#628780000000
0!
0*
09
0>
0C
#628790000000
1!
1*
b11 6
19
1>
1C
b11 G
#628800000000
0!
0*
09
0>
0C
#628810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#628820000000
0!
0*
09
0>
0C
#628830000000
1!
1*
b101 6
19
1>
1C
b101 G
#628840000000
0!
0*
09
0>
0C
#628850000000
1!
1*
b110 6
19
1>
1C
b110 G
#628860000000
0!
0*
09
0>
0C
#628870000000
1!
1*
b111 6
19
1>
1C
b111 G
#628880000000
0!
0*
09
0>
0C
#628890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#628900000000
0!
0*
09
0>
0C
#628910000000
1!
1*
b1 6
19
1>
1C
b1 G
#628920000000
0!
0*
09
0>
0C
#628930000000
1!
1*
b10 6
19
1>
1C
b10 G
#628940000000
0!
0*
09
0>
0C
#628950000000
1!
1*
b11 6
19
1>
1C
b11 G
#628960000000
0!
0*
09
0>
0C
#628970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#628980000000
0!
0*
09
0>
0C
#628990000000
1!
1*
b101 6
19
1>
1C
b101 G
#629000000000
0!
0*
09
0>
0C
#629010000000
1!
1*
b110 6
19
1>
1C
b110 G
#629020000000
0!
0*
09
0>
0C
#629030000000
1!
1*
b111 6
19
1>
1C
b111 G
#629040000000
0!
1"
0*
1+
09
1:
0>
0C
#629050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#629060000000
0!
0*
09
0>
0C
#629070000000
1!
1*
b1 6
19
1>
1C
b1 G
#629080000000
0!
0*
09
0>
0C
#629090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#629100000000
0!
0*
09
0>
0C
#629110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#629120000000
0!
0*
09
0>
0C
#629130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#629140000000
0!
0*
09
0>
0C
#629150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#629160000000
0!
0#
0*
0,
09
0>
0?
0C
#629170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#629180000000
0!
0*
09
0>
0C
#629190000000
1!
1*
19
1>
1C
#629200000000
0!
0*
09
0>
0C
#629210000000
1!
1*
19
1>
1C
#629220000000
0!
0*
09
0>
0C
#629230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#629240000000
0!
0*
09
0>
0C
#629250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#629260000000
0!
0*
09
0>
0C
#629270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#629280000000
0!
0*
09
0>
0C
#629290000000
1!
1*
b10 6
19
1>
1C
b10 G
#629300000000
0!
0*
09
0>
0C
#629310000000
1!
1*
b11 6
19
1>
1C
b11 G
#629320000000
0!
0*
09
0>
0C
#629330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#629340000000
0!
0*
09
0>
0C
#629350000000
1!
1*
b101 6
19
1>
1C
b101 G
#629360000000
0!
0*
09
0>
0C
#629370000000
1!
1*
b110 6
19
1>
1C
b110 G
#629380000000
0!
0*
09
0>
0C
#629390000000
1!
1*
b111 6
19
1>
1C
b111 G
#629400000000
0!
0*
09
0>
0C
#629410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#629420000000
0!
0*
09
0>
0C
#629430000000
1!
1*
b1 6
19
1>
1C
b1 G
#629440000000
0!
0*
09
0>
0C
#629450000000
1!
1*
b10 6
19
1>
1C
b10 G
#629460000000
0!
0*
09
0>
0C
#629470000000
1!
1*
b11 6
19
1>
1C
b11 G
#629480000000
0!
0*
09
0>
0C
#629490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#629500000000
0!
0*
09
0>
0C
#629510000000
1!
1*
b101 6
19
1>
1C
b101 G
#629520000000
0!
0*
09
0>
0C
#629530000000
1!
1*
b110 6
19
1>
1C
b110 G
#629540000000
0!
0*
09
0>
0C
#629550000000
1!
1*
b111 6
19
1>
1C
b111 G
#629560000000
0!
0*
09
0>
0C
#629570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#629580000000
0!
0*
09
0>
0C
#629590000000
1!
1*
b1 6
19
1>
1C
b1 G
#629600000000
0!
0*
09
0>
0C
#629610000000
1!
1*
b10 6
19
1>
1C
b10 G
#629620000000
0!
0*
09
0>
0C
#629630000000
1!
1*
b11 6
19
1>
1C
b11 G
#629640000000
0!
0*
09
0>
0C
#629650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#629660000000
0!
0*
09
0>
0C
#629670000000
1!
1*
b101 6
19
1>
1C
b101 G
#629680000000
0!
0*
09
0>
0C
#629690000000
1!
1*
b110 6
19
1>
1C
b110 G
#629700000000
0!
0*
09
0>
0C
#629710000000
1!
1*
b111 6
19
1>
1C
b111 G
#629720000000
0!
1"
0*
1+
09
1:
0>
0C
#629730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#629740000000
0!
0*
09
0>
0C
#629750000000
1!
1*
b1 6
19
1>
1C
b1 G
#629760000000
0!
0*
09
0>
0C
#629770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#629780000000
0!
0*
09
0>
0C
#629790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#629800000000
0!
0*
09
0>
0C
#629810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#629820000000
0!
0*
09
0>
0C
#629830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#629840000000
0!
0#
0*
0,
09
0>
0?
0C
#629850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#629860000000
0!
0*
09
0>
0C
#629870000000
1!
1*
19
1>
1C
#629880000000
0!
0*
09
0>
0C
#629890000000
1!
1*
19
1>
1C
#629900000000
0!
0*
09
0>
0C
#629910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#629920000000
0!
0*
09
0>
0C
#629930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#629940000000
0!
0*
09
0>
0C
#629950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#629960000000
0!
0*
09
0>
0C
#629970000000
1!
1*
b10 6
19
1>
1C
b10 G
#629980000000
0!
0*
09
0>
0C
#629990000000
1!
1*
b11 6
19
1>
1C
b11 G
#630000000000
0!
0*
09
0>
0C
#630010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#630020000000
0!
0*
09
0>
0C
#630030000000
1!
1*
b101 6
19
1>
1C
b101 G
#630040000000
0!
0*
09
0>
0C
#630050000000
1!
1*
b110 6
19
1>
1C
b110 G
#630060000000
0!
0*
09
0>
0C
#630070000000
1!
1*
b111 6
19
1>
1C
b111 G
#630080000000
0!
0*
09
0>
0C
#630090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#630100000000
0!
0*
09
0>
0C
#630110000000
1!
1*
b1 6
19
1>
1C
b1 G
#630120000000
0!
0*
09
0>
0C
#630130000000
1!
1*
b10 6
19
1>
1C
b10 G
#630140000000
0!
0*
09
0>
0C
#630150000000
1!
1*
b11 6
19
1>
1C
b11 G
#630160000000
0!
0*
09
0>
0C
#630170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#630180000000
0!
0*
09
0>
0C
#630190000000
1!
1*
b101 6
19
1>
1C
b101 G
#630200000000
0!
0*
09
0>
0C
#630210000000
1!
1*
b110 6
19
1>
1C
b110 G
#630220000000
0!
0*
09
0>
0C
#630230000000
1!
1*
b111 6
19
1>
1C
b111 G
#630240000000
0!
0*
09
0>
0C
#630250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#630260000000
0!
0*
09
0>
0C
#630270000000
1!
1*
b1 6
19
1>
1C
b1 G
#630280000000
0!
0*
09
0>
0C
#630290000000
1!
1*
b10 6
19
1>
1C
b10 G
#630300000000
0!
0*
09
0>
0C
#630310000000
1!
1*
b11 6
19
1>
1C
b11 G
#630320000000
0!
0*
09
0>
0C
#630330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#630340000000
0!
0*
09
0>
0C
#630350000000
1!
1*
b101 6
19
1>
1C
b101 G
#630360000000
0!
0*
09
0>
0C
#630370000000
1!
1*
b110 6
19
1>
1C
b110 G
#630380000000
0!
0*
09
0>
0C
#630390000000
1!
1*
b111 6
19
1>
1C
b111 G
#630400000000
0!
1"
0*
1+
09
1:
0>
0C
#630410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#630420000000
0!
0*
09
0>
0C
#630430000000
1!
1*
b1 6
19
1>
1C
b1 G
#630440000000
0!
0*
09
0>
0C
#630450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#630460000000
0!
0*
09
0>
0C
#630470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#630480000000
0!
0*
09
0>
0C
#630490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#630500000000
0!
0*
09
0>
0C
#630510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#630520000000
0!
0#
0*
0,
09
0>
0?
0C
#630530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#630540000000
0!
0*
09
0>
0C
#630550000000
1!
1*
19
1>
1C
#630560000000
0!
0*
09
0>
0C
#630570000000
1!
1*
19
1>
1C
#630580000000
0!
0*
09
0>
0C
#630590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#630600000000
0!
0*
09
0>
0C
#630610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#630620000000
0!
0*
09
0>
0C
#630630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#630640000000
0!
0*
09
0>
0C
#630650000000
1!
1*
b10 6
19
1>
1C
b10 G
#630660000000
0!
0*
09
0>
0C
#630670000000
1!
1*
b11 6
19
1>
1C
b11 G
#630680000000
0!
0*
09
0>
0C
#630690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#630700000000
0!
0*
09
0>
0C
#630710000000
1!
1*
b101 6
19
1>
1C
b101 G
#630720000000
0!
0*
09
0>
0C
#630730000000
1!
1*
b110 6
19
1>
1C
b110 G
#630740000000
0!
0*
09
0>
0C
#630750000000
1!
1*
b111 6
19
1>
1C
b111 G
#630760000000
0!
0*
09
0>
0C
#630770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#630780000000
0!
0*
09
0>
0C
#630790000000
1!
1*
b1 6
19
1>
1C
b1 G
#630800000000
0!
0*
09
0>
0C
#630810000000
1!
1*
b10 6
19
1>
1C
b10 G
#630820000000
0!
0*
09
0>
0C
#630830000000
1!
1*
b11 6
19
1>
1C
b11 G
#630840000000
0!
0*
09
0>
0C
#630850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#630860000000
0!
0*
09
0>
0C
#630870000000
1!
1*
b101 6
19
1>
1C
b101 G
#630880000000
0!
0*
09
0>
0C
#630890000000
1!
1*
b110 6
19
1>
1C
b110 G
#630900000000
0!
0*
09
0>
0C
#630910000000
1!
1*
b111 6
19
1>
1C
b111 G
#630920000000
0!
0*
09
0>
0C
#630930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#630940000000
0!
0*
09
0>
0C
#630950000000
1!
1*
b1 6
19
1>
1C
b1 G
#630960000000
0!
0*
09
0>
0C
#630970000000
1!
1*
b10 6
19
1>
1C
b10 G
#630980000000
0!
0*
09
0>
0C
#630990000000
1!
1*
b11 6
19
1>
1C
b11 G
#631000000000
0!
0*
09
0>
0C
#631010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#631020000000
0!
0*
09
0>
0C
#631030000000
1!
1*
b101 6
19
1>
1C
b101 G
#631040000000
0!
0*
09
0>
0C
#631050000000
1!
1*
b110 6
19
1>
1C
b110 G
#631060000000
0!
0*
09
0>
0C
#631070000000
1!
1*
b111 6
19
1>
1C
b111 G
#631080000000
0!
1"
0*
1+
09
1:
0>
0C
#631090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#631100000000
0!
0*
09
0>
0C
#631110000000
1!
1*
b1 6
19
1>
1C
b1 G
#631120000000
0!
0*
09
0>
0C
#631130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#631140000000
0!
0*
09
0>
0C
#631150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#631160000000
0!
0*
09
0>
0C
#631170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#631180000000
0!
0*
09
0>
0C
#631190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#631200000000
0!
0#
0*
0,
09
0>
0?
0C
#631210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#631220000000
0!
0*
09
0>
0C
#631230000000
1!
1*
19
1>
1C
#631240000000
0!
0*
09
0>
0C
#631250000000
1!
1*
19
1>
1C
#631260000000
0!
0*
09
0>
0C
#631270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#631280000000
0!
0*
09
0>
0C
#631290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#631300000000
0!
0*
09
0>
0C
#631310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#631320000000
0!
0*
09
0>
0C
#631330000000
1!
1*
b10 6
19
1>
1C
b10 G
#631340000000
0!
0*
09
0>
0C
#631350000000
1!
1*
b11 6
19
1>
1C
b11 G
#631360000000
0!
0*
09
0>
0C
#631370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#631380000000
0!
0*
09
0>
0C
#631390000000
1!
1*
b101 6
19
1>
1C
b101 G
#631400000000
0!
0*
09
0>
0C
#631410000000
1!
1*
b110 6
19
1>
1C
b110 G
#631420000000
0!
0*
09
0>
0C
#631430000000
1!
1*
b111 6
19
1>
1C
b111 G
#631440000000
0!
0*
09
0>
0C
#631450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#631460000000
0!
0*
09
0>
0C
#631470000000
1!
1*
b1 6
19
1>
1C
b1 G
#631480000000
0!
0*
09
0>
0C
#631490000000
1!
1*
b10 6
19
1>
1C
b10 G
#631500000000
0!
0*
09
0>
0C
#631510000000
1!
1*
b11 6
19
1>
1C
b11 G
#631520000000
0!
0*
09
0>
0C
#631530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#631540000000
0!
0*
09
0>
0C
#631550000000
1!
1*
b101 6
19
1>
1C
b101 G
#631560000000
0!
0*
09
0>
0C
#631570000000
1!
1*
b110 6
19
1>
1C
b110 G
#631580000000
0!
0*
09
0>
0C
#631590000000
1!
1*
b111 6
19
1>
1C
b111 G
#631600000000
0!
0*
09
0>
0C
#631610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#631620000000
0!
0*
09
0>
0C
#631630000000
1!
1*
b1 6
19
1>
1C
b1 G
#631640000000
0!
0*
09
0>
0C
#631650000000
1!
1*
b10 6
19
1>
1C
b10 G
#631660000000
0!
0*
09
0>
0C
#631670000000
1!
1*
b11 6
19
1>
1C
b11 G
#631680000000
0!
0*
09
0>
0C
#631690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#631700000000
0!
0*
09
0>
0C
#631710000000
1!
1*
b101 6
19
1>
1C
b101 G
#631720000000
0!
0*
09
0>
0C
#631730000000
1!
1*
b110 6
19
1>
1C
b110 G
#631740000000
0!
0*
09
0>
0C
#631750000000
1!
1*
b111 6
19
1>
1C
b111 G
#631760000000
0!
1"
0*
1+
09
1:
0>
0C
#631770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#631780000000
0!
0*
09
0>
0C
#631790000000
1!
1*
b1 6
19
1>
1C
b1 G
#631800000000
0!
0*
09
0>
0C
#631810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#631820000000
0!
0*
09
0>
0C
#631830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#631840000000
0!
0*
09
0>
0C
#631850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#631860000000
0!
0*
09
0>
0C
#631870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#631880000000
0!
0#
0*
0,
09
0>
0?
0C
#631890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#631900000000
0!
0*
09
0>
0C
#631910000000
1!
1*
19
1>
1C
#631920000000
0!
0*
09
0>
0C
#631930000000
1!
1*
19
1>
1C
#631940000000
0!
0*
09
0>
0C
#631950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#631960000000
0!
0*
09
0>
0C
#631970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#631980000000
0!
0*
09
0>
0C
#631990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#632000000000
0!
0*
09
0>
0C
#632010000000
1!
1*
b10 6
19
1>
1C
b10 G
#632020000000
0!
0*
09
0>
0C
#632030000000
1!
1*
b11 6
19
1>
1C
b11 G
#632040000000
0!
0*
09
0>
0C
#632050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#632060000000
0!
0*
09
0>
0C
#632070000000
1!
1*
b101 6
19
1>
1C
b101 G
#632080000000
0!
0*
09
0>
0C
#632090000000
1!
1*
b110 6
19
1>
1C
b110 G
#632100000000
0!
0*
09
0>
0C
#632110000000
1!
1*
b111 6
19
1>
1C
b111 G
#632120000000
0!
0*
09
0>
0C
#632130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#632140000000
0!
0*
09
0>
0C
#632150000000
1!
1*
b1 6
19
1>
1C
b1 G
#632160000000
0!
0*
09
0>
0C
#632170000000
1!
1*
b10 6
19
1>
1C
b10 G
#632180000000
0!
0*
09
0>
0C
#632190000000
1!
1*
b11 6
19
1>
1C
b11 G
#632200000000
0!
0*
09
0>
0C
#632210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#632220000000
0!
0*
09
0>
0C
#632230000000
1!
1*
b101 6
19
1>
1C
b101 G
#632240000000
0!
0*
09
0>
0C
#632250000000
1!
1*
b110 6
19
1>
1C
b110 G
#632260000000
0!
0*
09
0>
0C
#632270000000
1!
1*
b111 6
19
1>
1C
b111 G
#632280000000
0!
0*
09
0>
0C
#632290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#632300000000
0!
0*
09
0>
0C
#632310000000
1!
1*
b1 6
19
1>
1C
b1 G
#632320000000
0!
0*
09
0>
0C
#632330000000
1!
1*
b10 6
19
1>
1C
b10 G
#632340000000
0!
0*
09
0>
0C
#632350000000
1!
1*
b11 6
19
1>
1C
b11 G
#632360000000
0!
0*
09
0>
0C
#632370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#632380000000
0!
0*
09
0>
0C
#632390000000
1!
1*
b101 6
19
1>
1C
b101 G
#632400000000
0!
0*
09
0>
0C
#632410000000
1!
1*
b110 6
19
1>
1C
b110 G
#632420000000
0!
0*
09
0>
0C
#632430000000
1!
1*
b111 6
19
1>
1C
b111 G
#632440000000
0!
1"
0*
1+
09
1:
0>
0C
#632450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#632460000000
0!
0*
09
0>
0C
#632470000000
1!
1*
b1 6
19
1>
1C
b1 G
#632480000000
0!
0*
09
0>
0C
#632490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#632500000000
0!
0*
09
0>
0C
#632510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#632520000000
0!
0*
09
0>
0C
#632530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#632540000000
0!
0*
09
0>
0C
#632550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#632560000000
0!
0#
0*
0,
09
0>
0?
0C
#632570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#632580000000
0!
0*
09
0>
0C
#632590000000
1!
1*
19
1>
1C
#632600000000
0!
0*
09
0>
0C
#632610000000
1!
1*
19
1>
1C
#632620000000
0!
0*
09
0>
0C
#632630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#632640000000
0!
0*
09
0>
0C
#632650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#632660000000
0!
0*
09
0>
0C
#632670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#632680000000
0!
0*
09
0>
0C
#632690000000
1!
1*
b10 6
19
1>
1C
b10 G
#632700000000
0!
0*
09
0>
0C
#632710000000
1!
1*
b11 6
19
1>
1C
b11 G
#632720000000
0!
0*
09
0>
0C
#632730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#632740000000
0!
0*
09
0>
0C
#632750000000
1!
1*
b101 6
19
1>
1C
b101 G
#632760000000
0!
0*
09
0>
0C
#632770000000
1!
1*
b110 6
19
1>
1C
b110 G
#632780000000
0!
0*
09
0>
0C
#632790000000
1!
1*
b111 6
19
1>
1C
b111 G
#632800000000
0!
0*
09
0>
0C
#632810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#632820000000
0!
0*
09
0>
0C
#632830000000
1!
1*
b1 6
19
1>
1C
b1 G
#632840000000
0!
0*
09
0>
0C
#632850000000
1!
1*
b10 6
19
1>
1C
b10 G
#632860000000
0!
0*
09
0>
0C
#632870000000
1!
1*
b11 6
19
1>
1C
b11 G
#632880000000
0!
0*
09
0>
0C
#632890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#632900000000
0!
0*
09
0>
0C
#632910000000
1!
1*
b101 6
19
1>
1C
b101 G
#632920000000
0!
0*
09
0>
0C
#632930000000
1!
1*
b110 6
19
1>
1C
b110 G
#632940000000
0!
0*
09
0>
0C
#632950000000
1!
1*
b111 6
19
1>
1C
b111 G
#632960000000
0!
0*
09
0>
0C
#632970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#632980000000
0!
0*
09
0>
0C
#632990000000
1!
1*
b1 6
19
1>
1C
b1 G
#633000000000
0!
0*
09
0>
0C
#633010000000
1!
1*
b10 6
19
1>
1C
b10 G
#633020000000
0!
0*
09
0>
0C
#633030000000
1!
1*
b11 6
19
1>
1C
b11 G
#633040000000
0!
0*
09
0>
0C
#633050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#633060000000
0!
0*
09
0>
0C
#633070000000
1!
1*
b101 6
19
1>
1C
b101 G
#633080000000
0!
0*
09
0>
0C
#633090000000
1!
1*
b110 6
19
1>
1C
b110 G
#633100000000
0!
0*
09
0>
0C
#633110000000
1!
1*
b111 6
19
1>
1C
b111 G
#633120000000
0!
1"
0*
1+
09
1:
0>
0C
#633130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#633140000000
0!
0*
09
0>
0C
#633150000000
1!
1*
b1 6
19
1>
1C
b1 G
#633160000000
0!
0*
09
0>
0C
#633170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#633180000000
0!
0*
09
0>
0C
#633190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#633200000000
0!
0*
09
0>
0C
#633210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#633220000000
0!
0*
09
0>
0C
#633230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#633240000000
0!
0#
0*
0,
09
0>
0?
0C
#633250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#633260000000
0!
0*
09
0>
0C
#633270000000
1!
1*
19
1>
1C
#633280000000
0!
0*
09
0>
0C
#633290000000
1!
1*
19
1>
1C
#633300000000
0!
0*
09
0>
0C
#633310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#633320000000
0!
0*
09
0>
0C
#633330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#633340000000
0!
0*
09
0>
0C
#633350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#633360000000
0!
0*
09
0>
0C
#633370000000
1!
1*
b10 6
19
1>
1C
b10 G
#633380000000
0!
0*
09
0>
0C
#633390000000
1!
1*
b11 6
19
1>
1C
b11 G
#633400000000
0!
0*
09
0>
0C
#633410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#633420000000
0!
0*
09
0>
0C
#633430000000
1!
1*
b101 6
19
1>
1C
b101 G
#633440000000
0!
0*
09
0>
0C
#633450000000
1!
1*
b110 6
19
1>
1C
b110 G
#633460000000
0!
0*
09
0>
0C
#633470000000
1!
1*
b111 6
19
1>
1C
b111 G
#633480000000
0!
0*
09
0>
0C
#633490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#633500000000
0!
0*
09
0>
0C
#633510000000
1!
1*
b1 6
19
1>
1C
b1 G
#633520000000
0!
0*
09
0>
0C
#633530000000
1!
1*
b10 6
19
1>
1C
b10 G
#633540000000
0!
0*
09
0>
0C
#633550000000
1!
1*
b11 6
19
1>
1C
b11 G
#633560000000
0!
0*
09
0>
0C
#633570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#633580000000
0!
0*
09
0>
0C
#633590000000
1!
1*
b101 6
19
1>
1C
b101 G
#633600000000
0!
0*
09
0>
0C
#633610000000
1!
1*
b110 6
19
1>
1C
b110 G
#633620000000
0!
0*
09
0>
0C
#633630000000
1!
1*
b111 6
19
1>
1C
b111 G
#633640000000
0!
0*
09
0>
0C
#633650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#633660000000
0!
0*
09
0>
0C
#633670000000
1!
1*
b1 6
19
1>
1C
b1 G
#633680000000
0!
0*
09
0>
0C
#633690000000
1!
1*
b10 6
19
1>
1C
b10 G
#633700000000
0!
0*
09
0>
0C
#633710000000
1!
1*
b11 6
19
1>
1C
b11 G
#633720000000
0!
0*
09
0>
0C
#633730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#633740000000
0!
0*
09
0>
0C
#633750000000
1!
1*
b101 6
19
1>
1C
b101 G
#633760000000
0!
0*
09
0>
0C
#633770000000
1!
1*
b110 6
19
1>
1C
b110 G
#633780000000
0!
0*
09
0>
0C
#633790000000
1!
1*
b111 6
19
1>
1C
b111 G
#633800000000
0!
1"
0*
1+
09
1:
0>
0C
#633810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#633820000000
0!
0*
09
0>
0C
#633830000000
1!
1*
b1 6
19
1>
1C
b1 G
#633840000000
0!
0*
09
0>
0C
#633850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#633860000000
0!
0*
09
0>
0C
#633870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#633880000000
0!
0*
09
0>
0C
#633890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#633900000000
0!
0*
09
0>
0C
#633910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#633920000000
0!
0#
0*
0,
09
0>
0?
0C
#633930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#633940000000
0!
0*
09
0>
0C
#633950000000
1!
1*
19
1>
1C
#633960000000
0!
0*
09
0>
0C
#633970000000
1!
1*
19
1>
1C
#633980000000
0!
0*
09
0>
0C
#633990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#634000000000
0!
0*
09
0>
0C
#634010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#634020000000
0!
0*
09
0>
0C
#634030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#634040000000
0!
0*
09
0>
0C
#634050000000
1!
1*
b10 6
19
1>
1C
b10 G
#634060000000
0!
0*
09
0>
0C
#634070000000
1!
1*
b11 6
19
1>
1C
b11 G
#634080000000
0!
0*
09
0>
0C
#634090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#634100000000
0!
0*
09
0>
0C
#634110000000
1!
1*
b101 6
19
1>
1C
b101 G
#634120000000
0!
0*
09
0>
0C
#634130000000
1!
1*
b110 6
19
1>
1C
b110 G
#634140000000
0!
0*
09
0>
0C
#634150000000
1!
1*
b111 6
19
1>
1C
b111 G
#634160000000
0!
0*
09
0>
0C
#634170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#634180000000
0!
0*
09
0>
0C
#634190000000
1!
1*
b1 6
19
1>
1C
b1 G
#634200000000
0!
0*
09
0>
0C
#634210000000
1!
1*
b10 6
19
1>
1C
b10 G
#634220000000
0!
0*
09
0>
0C
#634230000000
1!
1*
b11 6
19
1>
1C
b11 G
#634240000000
0!
0*
09
0>
0C
#634250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#634260000000
0!
0*
09
0>
0C
#634270000000
1!
1*
b101 6
19
1>
1C
b101 G
#634280000000
0!
0*
09
0>
0C
#634290000000
1!
1*
b110 6
19
1>
1C
b110 G
#634300000000
0!
0*
09
0>
0C
#634310000000
1!
1*
b111 6
19
1>
1C
b111 G
#634320000000
0!
0*
09
0>
0C
#634330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#634340000000
0!
0*
09
0>
0C
#634350000000
1!
1*
b1 6
19
1>
1C
b1 G
#634360000000
0!
0*
09
0>
0C
#634370000000
1!
1*
b10 6
19
1>
1C
b10 G
#634380000000
0!
0*
09
0>
0C
#634390000000
1!
1*
b11 6
19
1>
1C
b11 G
#634400000000
0!
0*
09
0>
0C
#634410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#634420000000
0!
0*
09
0>
0C
#634430000000
1!
1*
b101 6
19
1>
1C
b101 G
#634440000000
0!
0*
09
0>
0C
#634450000000
1!
1*
b110 6
19
1>
1C
b110 G
#634460000000
0!
0*
09
0>
0C
#634470000000
1!
1*
b111 6
19
1>
1C
b111 G
#634480000000
0!
1"
0*
1+
09
1:
0>
0C
#634490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#634500000000
0!
0*
09
0>
0C
#634510000000
1!
1*
b1 6
19
1>
1C
b1 G
#634520000000
0!
0*
09
0>
0C
#634530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#634540000000
0!
0*
09
0>
0C
#634550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#634560000000
0!
0*
09
0>
0C
#634570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#634580000000
0!
0*
09
0>
0C
#634590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#634600000000
0!
0#
0*
0,
09
0>
0?
0C
#634610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#634620000000
0!
0*
09
0>
0C
#634630000000
1!
1*
19
1>
1C
#634640000000
0!
0*
09
0>
0C
#634650000000
1!
1*
19
1>
1C
#634660000000
0!
0*
09
0>
0C
#634670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#634680000000
0!
0*
09
0>
0C
#634690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#634700000000
0!
0*
09
0>
0C
#634710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#634720000000
0!
0*
09
0>
0C
#634730000000
1!
1*
b10 6
19
1>
1C
b10 G
#634740000000
0!
0*
09
0>
0C
#634750000000
1!
1*
b11 6
19
1>
1C
b11 G
#634760000000
0!
0*
09
0>
0C
#634770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#634780000000
0!
0*
09
0>
0C
#634790000000
1!
1*
b101 6
19
1>
1C
b101 G
#634800000000
0!
0*
09
0>
0C
#634810000000
1!
1*
b110 6
19
1>
1C
b110 G
#634820000000
0!
0*
09
0>
0C
#634830000000
1!
1*
b111 6
19
1>
1C
b111 G
#634840000000
0!
0*
09
0>
0C
#634850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#634860000000
0!
0*
09
0>
0C
#634870000000
1!
1*
b1 6
19
1>
1C
b1 G
#634880000000
0!
0*
09
0>
0C
#634890000000
1!
1*
b10 6
19
1>
1C
b10 G
#634900000000
0!
0*
09
0>
0C
#634910000000
1!
1*
b11 6
19
1>
1C
b11 G
#634920000000
0!
0*
09
0>
0C
#634930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#634940000000
0!
0*
09
0>
0C
#634950000000
1!
1*
b101 6
19
1>
1C
b101 G
#634960000000
0!
0*
09
0>
0C
#634970000000
1!
1*
b110 6
19
1>
1C
b110 G
#634980000000
0!
0*
09
0>
0C
#634990000000
1!
1*
b111 6
19
1>
1C
b111 G
#635000000000
0!
0*
09
0>
0C
#635010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#635020000000
0!
0*
09
0>
0C
#635030000000
1!
1*
b1 6
19
1>
1C
b1 G
#635040000000
0!
0*
09
0>
0C
#635050000000
1!
1*
b10 6
19
1>
1C
b10 G
#635060000000
0!
0*
09
0>
0C
#635070000000
1!
1*
b11 6
19
1>
1C
b11 G
#635080000000
0!
0*
09
0>
0C
#635090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#635100000000
0!
0*
09
0>
0C
#635110000000
1!
1*
b101 6
19
1>
1C
b101 G
#635120000000
0!
0*
09
0>
0C
#635130000000
1!
1*
b110 6
19
1>
1C
b110 G
#635140000000
0!
0*
09
0>
0C
#635150000000
1!
1*
b111 6
19
1>
1C
b111 G
#635160000000
0!
1"
0*
1+
09
1:
0>
0C
#635170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#635180000000
0!
0*
09
0>
0C
#635190000000
1!
1*
b1 6
19
1>
1C
b1 G
#635200000000
0!
0*
09
0>
0C
#635210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#635220000000
0!
0*
09
0>
0C
#635230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#635240000000
0!
0*
09
0>
0C
#635250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#635260000000
0!
0*
09
0>
0C
#635270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#635280000000
0!
0#
0*
0,
09
0>
0?
0C
#635290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#635300000000
0!
0*
09
0>
0C
#635310000000
1!
1*
19
1>
1C
#635320000000
0!
0*
09
0>
0C
#635330000000
1!
1*
19
1>
1C
#635340000000
0!
0*
09
0>
0C
#635350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#635360000000
0!
0*
09
0>
0C
#635370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#635380000000
0!
0*
09
0>
0C
#635390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#635400000000
0!
0*
09
0>
0C
#635410000000
1!
1*
b10 6
19
1>
1C
b10 G
#635420000000
0!
0*
09
0>
0C
#635430000000
1!
1*
b11 6
19
1>
1C
b11 G
#635440000000
0!
0*
09
0>
0C
#635450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#635460000000
0!
0*
09
0>
0C
#635470000000
1!
1*
b101 6
19
1>
1C
b101 G
#635480000000
0!
0*
09
0>
0C
#635490000000
1!
1*
b110 6
19
1>
1C
b110 G
#635500000000
0!
0*
09
0>
0C
#635510000000
1!
1*
b111 6
19
1>
1C
b111 G
#635520000000
0!
0*
09
0>
0C
#635530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#635540000000
0!
0*
09
0>
0C
#635550000000
1!
1*
b1 6
19
1>
1C
b1 G
#635560000000
0!
0*
09
0>
0C
#635570000000
1!
1*
b10 6
19
1>
1C
b10 G
#635580000000
0!
0*
09
0>
0C
#635590000000
1!
1*
b11 6
19
1>
1C
b11 G
#635600000000
0!
0*
09
0>
0C
#635610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#635620000000
0!
0*
09
0>
0C
#635630000000
1!
1*
b101 6
19
1>
1C
b101 G
#635640000000
0!
0*
09
0>
0C
#635650000000
1!
1*
b110 6
19
1>
1C
b110 G
#635660000000
0!
0*
09
0>
0C
#635670000000
1!
1*
b111 6
19
1>
1C
b111 G
#635680000000
0!
0*
09
0>
0C
#635690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#635700000000
0!
0*
09
0>
0C
#635710000000
1!
1*
b1 6
19
1>
1C
b1 G
#635720000000
0!
0*
09
0>
0C
#635730000000
1!
1*
b10 6
19
1>
1C
b10 G
#635740000000
0!
0*
09
0>
0C
#635750000000
1!
1*
b11 6
19
1>
1C
b11 G
#635760000000
0!
0*
09
0>
0C
#635770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#635780000000
0!
0*
09
0>
0C
#635790000000
1!
1*
b101 6
19
1>
1C
b101 G
#635800000000
0!
0*
09
0>
0C
#635810000000
1!
1*
b110 6
19
1>
1C
b110 G
#635820000000
0!
0*
09
0>
0C
#635830000000
1!
1*
b111 6
19
1>
1C
b111 G
#635840000000
0!
1"
0*
1+
09
1:
0>
0C
#635850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#635860000000
0!
0*
09
0>
0C
#635870000000
1!
1*
b1 6
19
1>
1C
b1 G
#635880000000
0!
0*
09
0>
0C
#635890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#635900000000
0!
0*
09
0>
0C
#635910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#635920000000
0!
0*
09
0>
0C
#635930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#635940000000
0!
0*
09
0>
0C
#635950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#635960000000
0!
0#
0*
0,
09
0>
0?
0C
#635970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#635980000000
0!
0*
09
0>
0C
#635990000000
1!
1*
19
1>
1C
#636000000000
0!
0*
09
0>
0C
#636010000000
1!
1*
19
1>
1C
#636020000000
0!
0*
09
0>
0C
#636030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#636040000000
0!
0*
09
0>
0C
#636050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#636060000000
0!
0*
09
0>
0C
#636070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#636080000000
0!
0*
09
0>
0C
#636090000000
1!
1*
b10 6
19
1>
1C
b10 G
#636100000000
0!
0*
09
0>
0C
#636110000000
1!
1*
b11 6
19
1>
1C
b11 G
#636120000000
0!
0*
09
0>
0C
#636130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#636140000000
0!
0*
09
0>
0C
#636150000000
1!
1*
b101 6
19
1>
1C
b101 G
#636160000000
0!
0*
09
0>
0C
#636170000000
1!
1*
b110 6
19
1>
1C
b110 G
#636180000000
0!
0*
09
0>
0C
#636190000000
1!
1*
b111 6
19
1>
1C
b111 G
#636200000000
0!
0*
09
0>
0C
#636210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#636220000000
0!
0*
09
0>
0C
#636230000000
1!
1*
b1 6
19
1>
1C
b1 G
#636240000000
0!
0*
09
0>
0C
#636250000000
1!
1*
b10 6
19
1>
1C
b10 G
#636260000000
0!
0*
09
0>
0C
#636270000000
1!
1*
b11 6
19
1>
1C
b11 G
#636280000000
0!
0*
09
0>
0C
#636290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#636300000000
0!
0*
09
0>
0C
#636310000000
1!
1*
b101 6
19
1>
1C
b101 G
#636320000000
0!
0*
09
0>
0C
#636330000000
1!
1*
b110 6
19
1>
1C
b110 G
#636340000000
0!
0*
09
0>
0C
#636350000000
1!
1*
b111 6
19
1>
1C
b111 G
#636360000000
0!
0*
09
0>
0C
#636370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#636380000000
0!
0*
09
0>
0C
#636390000000
1!
1*
b1 6
19
1>
1C
b1 G
#636400000000
0!
0*
09
0>
0C
#636410000000
1!
1*
b10 6
19
1>
1C
b10 G
#636420000000
0!
0*
09
0>
0C
#636430000000
1!
1*
b11 6
19
1>
1C
b11 G
#636440000000
0!
0*
09
0>
0C
#636450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#636460000000
0!
0*
09
0>
0C
#636470000000
1!
1*
b101 6
19
1>
1C
b101 G
#636480000000
0!
0*
09
0>
0C
#636490000000
1!
1*
b110 6
19
1>
1C
b110 G
#636500000000
0!
0*
09
0>
0C
#636510000000
1!
1*
b111 6
19
1>
1C
b111 G
#636520000000
0!
1"
0*
1+
09
1:
0>
0C
#636530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#636540000000
0!
0*
09
0>
0C
#636550000000
1!
1*
b1 6
19
1>
1C
b1 G
#636560000000
0!
0*
09
0>
0C
#636570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#636580000000
0!
0*
09
0>
0C
#636590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#636600000000
0!
0*
09
0>
0C
#636610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#636620000000
0!
0*
09
0>
0C
#636630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#636640000000
0!
0#
0*
0,
09
0>
0?
0C
#636650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#636660000000
0!
0*
09
0>
0C
#636670000000
1!
1*
19
1>
1C
#636680000000
0!
0*
09
0>
0C
#636690000000
1!
1*
19
1>
1C
#636700000000
0!
0*
09
0>
0C
#636710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#636720000000
0!
0*
09
0>
0C
#636730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#636740000000
0!
0*
09
0>
0C
#636750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#636760000000
0!
0*
09
0>
0C
#636770000000
1!
1*
b10 6
19
1>
1C
b10 G
#636780000000
0!
0*
09
0>
0C
#636790000000
1!
1*
b11 6
19
1>
1C
b11 G
#636800000000
0!
0*
09
0>
0C
#636810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#636820000000
0!
0*
09
0>
0C
#636830000000
1!
1*
b101 6
19
1>
1C
b101 G
#636840000000
0!
0*
09
0>
0C
#636850000000
1!
1*
b110 6
19
1>
1C
b110 G
#636860000000
0!
0*
09
0>
0C
#636870000000
1!
1*
b111 6
19
1>
1C
b111 G
#636880000000
0!
0*
09
0>
0C
#636890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#636900000000
0!
0*
09
0>
0C
#636910000000
1!
1*
b1 6
19
1>
1C
b1 G
#636920000000
0!
0*
09
0>
0C
#636930000000
1!
1*
b10 6
19
1>
1C
b10 G
#636940000000
0!
0*
09
0>
0C
#636950000000
1!
1*
b11 6
19
1>
1C
b11 G
#636960000000
0!
0*
09
0>
0C
#636970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#636980000000
0!
0*
09
0>
0C
#636990000000
1!
1*
b101 6
19
1>
1C
b101 G
#637000000000
0!
0*
09
0>
0C
#637010000000
1!
1*
b110 6
19
1>
1C
b110 G
#637020000000
0!
0*
09
0>
0C
#637030000000
1!
1*
b111 6
19
1>
1C
b111 G
#637040000000
0!
0*
09
0>
0C
#637050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#637060000000
0!
0*
09
0>
0C
#637070000000
1!
1*
b1 6
19
1>
1C
b1 G
#637080000000
0!
0*
09
0>
0C
#637090000000
1!
1*
b10 6
19
1>
1C
b10 G
#637100000000
0!
0*
09
0>
0C
#637110000000
1!
1*
b11 6
19
1>
1C
b11 G
#637120000000
0!
0*
09
0>
0C
#637130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#637140000000
0!
0*
09
0>
0C
#637150000000
1!
1*
b101 6
19
1>
1C
b101 G
#637160000000
0!
0*
09
0>
0C
#637170000000
1!
1*
b110 6
19
1>
1C
b110 G
#637180000000
0!
0*
09
0>
0C
#637190000000
1!
1*
b111 6
19
1>
1C
b111 G
#637200000000
0!
1"
0*
1+
09
1:
0>
0C
#637210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#637220000000
0!
0*
09
0>
0C
#637230000000
1!
1*
b1 6
19
1>
1C
b1 G
#637240000000
0!
0*
09
0>
0C
#637250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#637260000000
0!
0*
09
0>
0C
#637270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#637280000000
0!
0*
09
0>
0C
#637290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#637300000000
0!
0*
09
0>
0C
#637310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#637320000000
0!
0#
0*
0,
09
0>
0?
0C
#637330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#637340000000
0!
0*
09
0>
0C
#637350000000
1!
1*
19
1>
1C
#637360000000
0!
0*
09
0>
0C
#637370000000
1!
1*
19
1>
1C
#637380000000
0!
0*
09
0>
0C
#637390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#637400000000
0!
0*
09
0>
0C
#637410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#637420000000
0!
0*
09
0>
0C
#637430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#637440000000
0!
0*
09
0>
0C
#637450000000
1!
1*
b10 6
19
1>
1C
b10 G
#637460000000
0!
0*
09
0>
0C
#637470000000
1!
1*
b11 6
19
1>
1C
b11 G
#637480000000
0!
0*
09
0>
0C
#637490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#637500000000
0!
0*
09
0>
0C
#637510000000
1!
1*
b101 6
19
1>
1C
b101 G
#637520000000
0!
0*
09
0>
0C
#637530000000
1!
1*
b110 6
19
1>
1C
b110 G
#637540000000
0!
0*
09
0>
0C
#637550000000
1!
1*
b111 6
19
1>
1C
b111 G
#637560000000
0!
0*
09
0>
0C
#637570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#637580000000
0!
0*
09
0>
0C
#637590000000
1!
1*
b1 6
19
1>
1C
b1 G
#637600000000
0!
0*
09
0>
0C
#637610000000
1!
1*
b10 6
19
1>
1C
b10 G
#637620000000
0!
0*
09
0>
0C
#637630000000
1!
1*
b11 6
19
1>
1C
b11 G
#637640000000
0!
0*
09
0>
0C
#637650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#637660000000
0!
0*
09
0>
0C
#637670000000
1!
1*
b101 6
19
1>
1C
b101 G
#637680000000
0!
0*
09
0>
0C
#637690000000
1!
1*
b110 6
19
1>
1C
b110 G
#637700000000
0!
0*
09
0>
0C
#637710000000
1!
1*
b111 6
19
1>
1C
b111 G
#637720000000
0!
0*
09
0>
0C
#637730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#637740000000
0!
0*
09
0>
0C
#637750000000
1!
1*
b1 6
19
1>
1C
b1 G
#637760000000
0!
0*
09
0>
0C
#637770000000
1!
1*
b10 6
19
1>
1C
b10 G
#637780000000
0!
0*
09
0>
0C
#637790000000
1!
1*
b11 6
19
1>
1C
b11 G
#637800000000
0!
0*
09
0>
0C
#637810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#637820000000
0!
0*
09
0>
0C
#637830000000
1!
1*
b101 6
19
1>
1C
b101 G
#637840000000
0!
0*
09
0>
0C
#637850000000
1!
1*
b110 6
19
1>
1C
b110 G
#637860000000
0!
0*
09
0>
0C
#637870000000
1!
1*
b111 6
19
1>
1C
b111 G
#637880000000
0!
1"
0*
1+
09
1:
0>
0C
#637890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#637900000000
0!
0*
09
0>
0C
#637910000000
1!
1*
b1 6
19
1>
1C
b1 G
#637920000000
0!
0*
09
0>
0C
#637930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#637940000000
0!
0*
09
0>
0C
#637950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#637960000000
0!
0*
09
0>
0C
#637970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#637980000000
0!
0*
09
0>
0C
#637990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#638000000000
0!
0#
0*
0,
09
0>
0?
0C
#638010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#638020000000
0!
0*
09
0>
0C
#638030000000
1!
1*
19
1>
1C
#638040000000
0!
0*
09
0>
0C
#638050000000
1!
1*
19
1>
1C
#638060000000
0!
0*
09
0>
0C
#638070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#638080000000
0!
0*
09
0>
0C
#638090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#638100000000
0!
0*
09
0>
0C
#638110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#638120000000
0!
0*
09
0>
0C
#638130000000
1!
1*
b10 6
19
1>
1C
b10 G
#638140000000
0!
0*
09
0>
0C
#638150000000
1!
1*
b11 6
19
1>
1C
b11 G
#638160000000
0!
0*
09
0>
0C
#638170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#638180000000
0!
0*
09
0>
0C
#638190000000
1!
1*
b101 6
19
1>
1C
b101 G
#638200000000
0!
0*
09
0>
0C
#638210000000
1!
1*
b110 6
19
1>
1C
b110 G
#638220000000
0!
0*
09
0>
0C
#638230000000
1!
1*
b111 6
19
1>
1C
b111 G
#638240000000
0!
0*
09
0>
0C
#638250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#638260000000
0!
0*
09
0>
0C
#638270000000
1!
1*
b1 6
19
1>
1C
b1 G
#638280000000
0!
0*
09
0>
0C
#638290000000
1!
1*
b10 6
19
1>
1C
b10 G
#638300000000
0!
0*
09
0>
0C
#638310000000
1!
1*
b11 6
19
1>
1C
b11 G
#638320000000
0!
0*
09
0>
0C
#638330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#638340000000
0!
0*
09
0>
0C
#638350000000
1!
1*
b101 6
19
1>
1C
b101 G
#638360000000
0!
0*
09
0>
0C
#638370000000
1!
1*
b110 6
19
1>
1C
b110 G
#638380000000
0!
0*
09
0>
0C
#638390000000
1!
1*
b111 6
19
1>
1C
b111 G
#638400000000
0!
0*
09
0>
0C
#638410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#638420000000
0!
0*
09
0>
0C
#638430000000
1!
1*
b1 6
19
1>
1C
b1 G
#638440000000
0!
0*
09
0>
0C
#638450000000
1!
1*
b10 6
19
1>
1C
b10 G
#638460000000
0!
0*
09
0>
0C
#638470000000
1!
1*
b11 6
19
1>
1C
b11 G
#638480000000
0!
0*
09
0>
0C
#638490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#638500000000
0!
0*
09
0>
0C
#638510000000
1!
1*
b101 6
19
1>
1C
b101 G
#638520000000
0!
0*
09
0>
0C
#638530000000
1!
1*
b110 6
19
1>
1C
b110 G
#638540000000
0!
0*
09
0>
0C
#638550000000
1!
1*
b111 6
19
1>
1C
b111 G
#638560000000
0!
1"
0*
1+
09
1:
0>
0C
#638570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#638580000000
0!
0*
09
0>
0C
#638590000000
1!
1*
b1 6
19
1>
1C
b1 G
#638600000000
0!
0*
09
0>
0C
#638610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#638620000000
0!
0*
09
0>
0C
#638630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#638640000000
0!
0*
09
0>
0C
#638650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#638660000000
0!
0*
09
0>
0C
#638670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#638680000000
0!
0#
0*
0,
09
0>
0?
0C
#638690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#638700000000
0!
0*
09
0>
0C
#638710000000
1!
1*
19
1>
1C
#638720000000
0!
0*
09
0>
0C
#638730000000
1!
1*
19
1>
1C
#638740000000
0!
0*
09
0>
0C
#638750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#638760000000
0!
0*
09
0>
0C
#638770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#638780000000
0!
0*
09
0>
0C
#638790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#638800000000
0!
0*
09
0>
0C
#638810000000
1!
1*
b10 6
19
1>
1C
b10 G
#638820000000
0!
0*
09
0>
0C
#638830000000
1!
1*
b11 6
19
1>
1C
b11 G
#638840000000
0!
0*
09
0>
0C
#638850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#638860000000
0!
0*
09
0>
0C
#638870000000
1!
1*
b101 6
19
1>
1C
b101 G
#638880000000
0!
0*
09
0>
0C
#638890000000
1!
1*
b110 6
19
1>
1C
b110 G
#638900000000
0!
0*
09
0>
0C
#638910000000
1!
1*
b111 6
19
1>
1C
b111 G
#638920000000
0!
0*
09
0>
0C
#638930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#638940000000
0!
0*
09
0>
0C
#638950000000
1!
1*
b1 6
19
1>
1C
b1 G
#638960000000
0!
0*
09
0>
0C
#638970000000
1!
1*
b10 6
19
1>
1C
b10 G
#638980000000
0!
0*
09
0>
0C
#638990000000
1!
1*
b11 6
19
1>
1C
b11 G
#639000000000
0!
0*
09
0>
0C
#639010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#639020000000
0!
0*
09
0>
0C
#639030000000
1!
1*
b101 6
19
1>
1C
b101 G
#639040000000
0!
0*
09
0>
0C
#639050000000
1!
1*
b110 6
19
1>
1C
b110 G
#639060000000
0!
0*
09
0>
0C
#639070000000
1!
1*
b111 6
19
1>
1C
b111 G
#639080000000
0!
0*
09
0>
0C
#639090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#639100000000
0!
0*
09
0>
0C
#639110000000
1!
1*
b1 6
19
1>
1C
b1 G
#639120000000
0!
0*
09
0>
0C
#639130000000
1!
1*
b10 6
19
1>
1C
b10 G
#639140000000
0!
0*
09
0>
0C
#639150000000
1!
1*
b11 6
19
1>
1C
b11 G
#639160000000
0!
0*
09
0>
0C
#639170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#639180000000
0!
0*
09
0>
0C
#639190000000
1!
1*
b101 6
19
1>
1C
b101 G
#639200000000
0!
0*
09
0>
0C
#639210000000
1!
1*
b110 6
19
1>
1C
b110 G
#639220000000
0!
0*
09
0>
0C
#639230000000
1!
1*
b111 6
19
1>
1C
b111 G
#639240000000
0!
1"
0*
1+
09
1:
0>
0C
#639250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#639260000000
0!
0*
09
0>
0C
#639270000000
1!
1*
b1 6
19
1>
1C
b1 G
#639280000000
0!
0*
09
0>
0C
#639290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#639300000000
0!
0*
09
0>
0C
#639310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#639320000000
0!
0*
09
0>
0C
#639330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#639340000000
0!
0*
09
0>
0C
#639350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#639360000000
0!
0#
0*
0,
09
0>
0?
0C
#639370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#639380000000
0!
0*
09
0>
0C
#639390000000
1!
1*
19
1>
1C
#639400000000
0!
0*
09
0>
0C
#639410000000
1!
1*
19
1>
1C
#639420000000
0!
0*
09
0>
0C
#639430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#639440000000
0!
0*
09
0>
0C
#639450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#639460000000
0!
0*
09
0>
0C
#639470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#639480000000
0!
0*
09
0>
0C
#639490000000
1!
1*
b10 6
19
1>
1C
b10 G
#639500000000
0!
0*
09
0>
0C
#639510000000
1!
1*
b11 6
19
1>
1C
b11 G
#639520000000
0!
0*
09
0>
0C
#639530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#639540000000
0!
0*
09
0>
0C
#639550000000
1!
1*
b101 6
19
1>
1C
b101 G
#639560000000
0!
0*
09
0>
0C
#639570000000
1!
1*
b110 6
19
1>
1C
b110 G
#639580000000
0!
0*
09
0>
0C
#639590000000
1!
1*
b111 6
19
1>
1C
b111 G
#639600000000
0!
0*
09
0>
0C
#639610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#639620000000
0!
0*
09
0>
0C
#639630000000
1!
1*
b1 6
19
1>
1C
b1 G
#639640000000
0!
0*
09
0>
0C
#639650000000
1!
1*
b10 6
19
1>
1C
b10 G
#639660000000
0!
0*
09
0>
0C
#639670000000
1!
1*
b11 6
19
1>
1C
b11 G
#639680000000
0!
0*
09
0>
0C
#639690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#639700000000
0!
0*
09
0>
0C
#639710000000
1!
1*
b101 6
19
1>
1C
b101 G
#639720000000
0!
0*
09
0>
0C
#639730000000
1!
1*
b110 6
19
1>
1C
b110 G
#639740000000
0!
0*
09
0>
0C
#639750000000
1!
1*
b111 6
19
1>
1C
b111 G
#639760000000
0!
0*
09
0>
0C
#639770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#639780000000
0!
0*
09
0>
0C
#639790000000
1!
1*
b1 6
19
1>
1C
b1 G
#639800000000
0!
0*
09
0>
0C
#639810000000
1!
1*
b10 6
19
1>
1C
b10 G
#639820000000
0!
0*
09
0>
0C
#639830000000
1!
1*
b11 6
19
1>
1C
b11 G
#639840000000
0!
0*
09
0>
0C
#639850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#639860000000
0!
0*
09
0>
0C
#639870000000
1!
1*
b101 6
19
1>
1C
b101 G
#639880000000
0!
0*
09
0>
0C
#639890000000
1!
1*
b110 6
19
1>
1C
b110 G
#639900000000
0!
0*
09
0>
0C
#639910000000
1!
1*
b111 6
19
1>
1C
b111 G
#639920000000
0!
1"
0*
1+
09
1:
0>
0C
#639930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#639940000000
0!
0*
09
0>
0C
#639950000000
1!
1*
b1 6
19
1>
1C
b1 G
#639960000000
0!
0*
09
0>
0C
#639970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#639980000000
0!
0*
09
0>
0C
#639990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#640000000000
0!
0*
09
0>
0C
#640010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#640020000000
0!
0*
09
0>
0C
#640030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#640040000000
0!
0#
0*
0,
09
0>
0?
0C
#640050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#640060000000
0!
0*
09
0>
0C
#640070000000
1!
1*
19
1>
1C
#640080000000
0!
0*
09
0>
0C
#640090000000
1!
1*
19
1>
1C
#640100000000
0!
0*
09
0>
0C
#640110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#640120000000
0!
0*
09
0>
0C
#640130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#640140000000
0!
0*
09
0>
0C
#640150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#640160000000
0!
0*
09
0>
0C
#640170000000
1!
1*
b10 6
19
1>
1C
b10 G
#640180000000
0!
0*
09
0>
0C
#640190000000
1!
1*
b11 6
19
1>
1C
b11 G
#640200000000
0!
0*
09
0>
0C
#640210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#640220000000
0!
0*
09
0>
0C
#640230000000
1!
1*
b101 6
19
1>
1C
b101 G
#640240000000
0!
0*
09
0>
0C
#640250000000
1!
1*
b110 6
19
1>
1C
b110 G
#640260000000
0!
0*
09
0>
0C
#640270000000
1!
1*
b111 6
19
1>
1C
b111 G
#640280000000
0!
0*
09
0>
0C
#640290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#640300000000
0!
0*
09
0>
0C
#640310000000
1!
1*
b1 6
19
1>
1C
b1 G
#640320000000
0!
0*
09
0>
0C
#640330000000
1!
1*
b10 6
19
1>
1C
b10 G
#640340000000
0!
0*
09
0>
0C
#640350000000
1!
1*
b11 6
19
1>
1C
b11 G
#640360000000
0!
0*
09
0>
0C
#640370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#640380000000
0!
0*
09
0>
0C
#640390000000
1!
1*
b101 6
19
1>
1C
b101 G
#640400000000
0!
0*
09
0>
0C
#640410000000
1!
1*
b110 6
19
1>
1C
b110 G
#640420000000
0!
0*
09
0>
0C
#640430000000
1!
1*
b111 6
19
1>
1C
b111 G
#640440000000
0!
0*
09
0>
0C
#640450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#640460000000
0!
0*
09
0>
0C
#640470000000
1!
1*
b1 6
19
1>
1C
b1 G
#640480000000
0!
0*
09
0>
0C
#640490000000
1!
1*
b10 6
19
1>
1C
b10 G
#640500000000
0!
0*
09
0>
0C
#640510000000
1!
1*
b11 6
19
1>
1C
b11 G
#640520000000
0!
0*
09
0>
0C
#640530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#640540000000
0!
0*
09
0>
0C
#640550000000
1!
1*
b101 6
19
1>
1C
b101 G
#640560000000
0!
0*
09
0>
0C
#640570000000
1!
1*
b110 6
19
1>
1C
b110 G
#640580000000
0!
0*
09
0>
0C
#640590000000
1!
1*
b111 6
19
1>
1C
b111 G
#640600000000
0!
1"
0*
1+
09
1:
0>
0C
#640610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#640620000000
0!
0*
09
0>
0C
#640630000000
1!
1*
b1 6
19
1>
1C
b1 G
#640640000000
0!
0*
09
0>
0C
#640650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#640660000000
0!
0*
09
0>
0C
#640670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#640680000000
0!
0*
09
0>
0C
#640690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#640700000000
0!
0*
09
0>
0C
#640710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#640720000000
0!
0#
0*
0,
09
0>
0?
0C
#640730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#640740000000
0!
0*
09
0>
0C
#640750000000
1!
1*
19
1>
1C
#640760000000
0!
0*
09
0>
0C
#640770000000
1!
1*
19
1>
1C
#640780000000
0!
0*
09
0>
0C
#640790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#640800000000
0!
0*
09
0>
0C
#640810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#640820000000
0!
0*
09
0>
0C
#640830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#640840000000
0!
0*
09
0>
0C
#640850000000
1!
1*
b10 6
19
1>
1C
b10 G
#640860000000
0!
0*
09
0>
0C
#640870000000
1!
1*
b11 6
19
1>
1C
b11 G
#640880000000
0!
0*
09
0>
0C
#640890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#640900000000
0!
0*
09
0>
0C
#640910000000
1!
1*
b101 6
19
1>
1C
b101 G
#640920000000
0!
0*
09
0>
0C
#640930000000
1!
1*
b110 6
19
1>
1C
b110 G
#640940000000
0!
0*
09
0>
0C
#640950000000
1!
1*
b111 6
19
1>
1C
b111 G
#640960000000
0!
0*
09
0>
0C
#640970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#640980000000
0!
0*
09
0>
0C
#640990000000
1!
1*
b1 6
19
1>
1C
b1 G
#641000000000
0!
0*
09
0>
0C
#641010000000
1!
1*
b10 6
19
1>
1C
b10 G
#641020000000
0!
0*
09
0>
0C
#641030000000
1!
1*
b11 6
19
1>
1C
b11 G
#641040000000
0!
0*
09
0>
0C
#641050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#641060000000
0!
0*
09
0>
0C
#641070000000
1!
1*
b101 6
19
1>
1C
b101 G
#641080000000
0!
0*
09
0>
0C
#641090000000
1!
1*
b110 6
19
1>
1C
b110 G
#641100000000
0!
0*
09
0>
0C
#641110000000
1!
1*
b111 6
19
1>
1C
b111 G
#641120000000
0!
0*
09
0>
0C
#641130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#641140000000
0!
0*
09
0>
0C
#641150000000
1!
1*
b1 6
19
1>
1C
b1 G
#641160000000
0!
0*
09
0>
0C
#641170000000
1!
1*
b10 6
19
1>
1C
b10 G
#641180000000
0!
0*
09
0>
0C
#641190000000
1!
1*
b11 6
19
1>
1C
b11 G
#641200000000
0!
0*
09
0>
0C
#641210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#641220000000
0!
0*
09
0>
0C
#641230000000
1!
1*
b101 6
19
1>
1C
b101 G
#641240000000
0!
0*
09
0>
0C
#641250000000
1!
1*
b110 6
19
1>
1C
b110 G
#641260000000
0!
0*
09
0>
0C
#641270000000
1!
1*
b111 6
19
1>
1C
b111 G
#641280000000
0!
1"
0*
1+
09
1:
0>
0C
#641290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#641300000000
0!
0*
09
0>
0C
#641310000000
1!
1*
b1 6
19
1>
1C
b1 G
#641320000000
0!
0*
09
0>
0C
#641330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#641340000000
0!
0*
09
0>
0C
#641350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#641360000000
0!
0*
09
0>
0C
#641370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#641380000000
0!
0*
09
0>
0C
#641390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#641400000000
0!
0#
0*
0,
09
0>
0?
0C
#641410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#641420000000
0!
0*
09
0>
0C
#641430000000
1!
1*
19
1>
1C
#641440000000
0!
0*
09
0>
0C
#641450000000
1!
1*
19
1>
1C
#641460000000
0!
0*
09
0>
0C
#641470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#641480000000
0!
0*
09
0>
0C
#641490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#641500000000
0!
0*
09
0>
0C
#641510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#641520000000
0!
0*
09
0>
0C
#641530000000
1!
1*
b10 6
19
1>
1C
b10 G
#641540000000
0!
0*
09
0>
0C
#641550000000
1!
1*
b11 6
19
1>
1C
b11 G
#641560000000
0!
0*
09
0>
0C
#641570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#641580000000
0!
0*
09
0>
0C
#641590000000
1!
1*
b101 6
19
1>
1C
b101 G
#641600000000
0!
0*
09
0>
0C
#641610000000
1!
1*
b110 6
19
1>
1C
b110 G
#641620000000
0!
0*
09
0>
0C
#641630000000
1!
1*
b111 6
19
1>
1C
b111 G
#641640000000
0!
0*
09
0>
0C
#641650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#641660000000
0!
0*
09
0>
0C
#641670000000
1!
1*
b1 6
19
1>
1C
b1 G
#641680000000
0!
0*
09
0>
0C
#641690000000
1!
1*
b10 6
19
1>
1C
b10 G
#641700000000
0!
0*
09
0>
0C
#641710000000
1!
1*
b11 6
19
1>
1C
b11 G
#641720000000
0!
0*
09
0>
0C
#641730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#641740000000
0!
0*
09
0>
0C
#641750000000
1!
1*
b101 6
19
1>
1C
b101 G
#641760000000
0!
0*
09
0>
0C
#641770000000
1!
1*
b110 6
19
1>
1C
b110 G
#641780000000
0!
0*
09
0>
0C
#641790000000
1!
1*
b111 6
19
1>
1C
b111 G
#641800000000
0!
0*
09
0>
0C
#641810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#641820000000
0!
0*
09
0>
0C
#641830000000
1!
1*
b1 6
19
1>
1C
b1 G
#641840000000
0!
0*
09
0>
0C
#641850000000
1!
1*
b10 6
19
1>
1C
b10 G
#641860000000
0!
0*
09
0>
0C
#641870000000
1!
1*
b11 6
19
1>
1C
b11 G
#641880000000
0!
0*
09
0>
0C
#641890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#641900000000
0!
0*
09
0>
0C
#641910000000
1!
1*
b101 6
19
1>
1C
b101 G
#641920000000
0!
0*
09
0>
0C
#641930000000
1!
1*
b110 6
19
1>
1C
b110 G
#641940000000
0!
0*
09
0>
0C
#641950000000
1!
1*
b111 6
19
1>
1C
b111 G
#641960000000
0!
1"
0*
1+
09
1:
0>
0C
#641970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#641980000000
0!
0*
09
0>
0C
#641990000000
1!
1*
b1 6
19
1>
1C
b1 G
#642000000000
0!
0*
09
0>
0C
#642010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#642020000000
0!
0*
09
0>
0C
#642030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#642040000000
0!
0*
09
0>
0C
#642050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#642060000000
0!
0*
09
0>
0C
#642070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#642080000000
0!
0#
0*
0,
09
0>
0?
0C
#642090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#642100000000
0!
0*
09
0>
0C
#642110000000
1!
1*
19
1>
1C
#642120000000
0!
0*
09
0>
0C
#642130000000
1!
1*
19
1>
1C
#642140000000
0!
0*
09
0>
0C
#642150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#642160000000
0!
0*
09
0>
0C
#642170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#642180000000
0!
0*
09
0>
0C
#642190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#642200000000
0!
0*
09
0>
0C
#642210000000
1!
1*
b10 6
19
1>
1C
b10 G
#642220000000
0!
0*
09
0>
0C
#642230000000
1!
1*
b11 6
19
1>
1C
b11 G
#642240000000
0!
0*
09
0>
0C
#642250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#642260000000
0!
0*
09
0>
0C
#642270000000
1!
1*
b101 6
19
1>
1C
b101 G
#642280000000
0!
0*
09
0>
0C
#642290000000
1!
1*
b110 6
19
1>
1C
b110 G
#642300000000
0!
0*
09
0>
0C
#642310000000
1!
1*
b111 6
19
1>
1C
b111 G
#642320000000
0!
0*
09
0>
0C
#642330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#642340000000
0!
0*
09
0>
0C
#642350000000
1!
1*
b1 6
19
1>
1C
b1 G
#642360000000
0!
0*
09
0>
0C
#642370000000
1!
1*
b10 6
19
1>
1C
b10 G
#642380000000
0!
0*
09
0>
0C
#642390000000
1!
1*
b11 6
19
1>
1C
b11 G
#642400000000
0!
0*
09
0>
0C
#642410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#642420000000
0!
0*
09
0>
0C
#642430000000
1!
1*
b101 6
19
1>
1C
b101 G
#642440000000
0!
0*
09
0>
0C
#642450000000
1!
1*
b110 6
19
1>
1C
b110 G
#642460000000
0!
0*
09
0>
0C
#642470000000
1!
1*
b111 6
19
1>
1C
b111 G
#642480000000
0!
0*
09
0>
0C
#642490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#642500000000
0!
0*
09
0>
0C
#642510000000
1!
1*
b1 6
19
1>
1C
b1 G
#642520000000
0!
0*
09
0>
0C
#642530000000
1!
1*
b10 6
19
1>
1C
b10 G
#642540000000
0!
0*
09
0>
0C
#642550000000
1!
1*
b11 6
19
1>
1C
b11 G
#642560000000
0!
0*
09
0>
0C
#642570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#642580000000
0!
0*
09
0>
0C
#642590000000
1!
1*
b101 6
19
1>
1C
b101 G
#642600000000
0!
0*
09
0>
0C
#642610000000
1!
1*
b110 6
19
1>
1C
b110 G
#642620000000
0!
0*
09
0>
0C
#642630000000
1!
1*
b111 6
19
1>
1C
b111 G
#642640000000
0!
1"
0*
1+
09
1:
0>
0C
#642650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#642660000000
0!
0*
09
0>
0C
#642670000000
1!
1*
b1 6
19
1>
1C
b1 G
#642680000000
0!
0*
09
0>
0C
#642690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#642700000000
0!
0*
09
0>
0C
#642710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#642720000000
0!
0*
09
0>
0C
#642730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#642740000000
0!
0*
09
0>
0C
#642750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#642760000000
0!
0#
0*
0,
09
0>
0?
0C
#642770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#642780000000
0!
0*
09
0>
0C
#642790000000
1!
1*
19
1>
1C
#642800000000
0!
0*
09
0>
0C
#642810000000
1!
1*
19
1>
1C
#642820000000
0!
0*
09
0>
0C
#642830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#642840000000
0!
0*
09
0>
0C
#642850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#642860000000
0!
0*
09
0>
0C
#642870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#642880000000
0!
0*
09
0>
0C
#642890000000
1!
1*
b10 6
19
1>
1C
b10 G
#642900000000
0!
0*
09
0>
0C
#642910000000
1!
1*
b11 6
19
1>
1C
b11 G
#642920000000
0!
0*
09
0>
0C
#642930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#642940000000
0!
0*
09
0>
0C
#642950000000
1!
1*
b101 6
19
1>
1C
b101 G
#642960000000
0!
0*
09
0>
0C
#642970000000
1!
1*
b110 6
19
1>
1C
b110 G
#642980000000
0!
0*
09
0>
0C
#642990000000
1!
1*
b111 6
19
1>
1C
b111 G
#643000000000
0!
0*
09
0>
0C
#643010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#643020000000
0!
0*
09
0>
0C
#643030000000
1!
1*
b1 6
19
1>
1C
b1 G
#643040000000
0!
0*
09
0>
0C
#643050000000
1!
1*
b10 6
19
1>
1C
b10 G
#643060000000
0!
0*
09
0>
0C
#643070000000
1!
1*
b11 6
19
1>
1C
b11 G
#643080000000
0!
0*
09
0>
0C
#643090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#643100000000
0!
0*
09
0>
0C
#643110000000
1!
1*
b101 6
19
1>
1C
b101 G
#643120000000
0!
0*
09
0>
0C
#643130000000
1!
1*
b110 6
19
1>
1C
b110 G
#643140000000
0!
0*
09
0>
0C
#643150000000
1!
1*
b111 6
19
1>
1C
b111 G
#643160000000
0!
0*
09
0>
0C
#643170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#643180000000
0!
0*
09
0>
0C
#643190000000
1!
1*
b1 6
19
1>
1C
b1 G
#643200000000
0!
0*
09
0>
0C
#643210000000
1!
1*
b10 6
19
1>
1C
b10 G
#643220000000
0!
0*
09
0>
0C
#643230000000
1!
1*
b11 6
19
1>
1C
b11 G
#643240000000
0!
0*
09
0>
0C
#643250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#643260000000
0!
0*
09
0>
0C
#643270000000
1!
1*
b101 6
19
1>
1C
b101 G
#643280000000
0!
0*
09
0>
0C
#643290000000
1!
1*
b110 6
19
1>
1C
b110 G
#643300000000
0!
0*
09
0>
0C
#643310000000
1!
1*
b111 6
19
1>
1C
b111 G
#643320000000
0!
1"
0*
1+
09
1:
0>
0C
#643330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#643340000000
0!
0*
09
0>
0C
#643350000000
1!
1*
b1 6
19
1>
1C
b1 G
#643360000000
0!
0*
09
0>
0C
#643370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#643380000000
0!
0*
09
0>
0C
#643390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#643400000000
0!
0*
09
0>
0C
#643410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#643420000000
0!
0*
09
0>
0C
#643430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#643440000000
0!
0#
0*
0,
09
0>
0?
0C
#643450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#643460000000
0!
0*
09
0>
0C
#643470000000
1!
1*
19
1>
1C
#643480000000
0!
0*
09
0>
0C
#643490000000
1!
1*
19
1>
1C
#643500000000
0!
0*
09
0>
0C
#643510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#643520000000
0!
0*
09
0>
0C
#643530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#643540000000
0!
0*
09
0>
0C
#643550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#643560000000
0!
0*
09
0>
0C
#643570000000
1!
1*
b10 6
19
1>
1C
b10 G
#643580000000
0!
0*
09
0>
0C
#643590000000
1!
1*
b11 6
19
1>
1C
b11 G
#643600000000
0!
0*
09
0>
0C
#643610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#643620000000
0!
0*
09
0>
0C
#643630000000
1!
1*
b101 6
19
1>
1C
b101 G
#643640000000
0!
0*
09
0>
0C
#643650000000
1!
1*
b110 6
19
1>
1C
b110 G
#643660000000
0!
0*
09
0>
0C
#643670000000
1!
1*
b111 6
19
1>
1C
b111 G
#643680000000
0!
0*
09
0>
0C
#643690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#643700000000
0!
0*
09
0>
0C
#643710000000
1!
1*
b1 6
19
1>
1C
b1 G
#643720000000
0!
0*
09
0>
0C
#643730000000
1!
1*
b10 6
19
1>
1C
b10 G
#643740000000
0!
0*
09
0>
0C
#643750000000
1!
1*
b11 6
19
1>
1C
b11 G
#643760000000
0!
0*
09
0>
0C
#643770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#643780000000
0!
0*
09
0>
0C
#643790000000
1!
1*
b101 6
19
1>
1C
b101 G
#643800000000
0!
0*
09
0>
0C
#643810000000
1!
1*
b110 6
19
1>
1C
b110 G
#643820000000
0!
0*
09
0>
0C
#643830000000
1!
1*
b111 6
19
1>
1C
b111 G
#643840000000
0!
0*
09
0>
0C
#643850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#643860000000
0!
0*
09
0>
0C
#643870000000
1!
1*
b1 6
19
1>
1C
b1 G
#643880000000
0!
0*
09
0>
0C
#643890000000
1!
1*
b10 6
19
1>
1C
b10 G
#643900000000
0!
0*
09
0>
0C
#643910000000
1!
1*
b11 6
19
1>
1C
b11 G
#643920000000
0!
0*
09
0>
0C
#643930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#643940000000
0!
0*
09
0>
0C
#643950000000
1!
1*
b101 6
19
1>
1C
b101 G
#643960000000
0!
0*
09
0>
0C
#643970000000
1!
1*
b110 6
19
1>
1C
b110 G
#643980000000
0!
0*
09
0>
0C
#643990000000
1!
1*
b111 6
19
1>
1C
b111 G
#644000000000
0!
1"
0*
1+
09
1:
0>
0C
#644010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#644020000000
0!
0*
09
0>
0C
#644030000000
1!
1*
b1 6
19
1>
1C
b1 G
#644040000000
0!
0*
09
0>
0C
#644050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#644060000000
0!
0*
09
0>
0C
#644070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#644080000000
0!
0*
09
0>
0C
#644090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#644100000000
0!
0*
09
0>
0C
#644110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#644120000000
0!
0#
0*
0,
09
0>
0?
0C
#644130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#644140000000
0!
0*
09
0>
0C
#644150000000
1!
1*
19
1>
1C
#644160000000
0!
0*
09
0>
0C
#644170000000
1!
1*
19
1>
1C
#644180000000
0!
0*
09
0>
0C
#644190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#644200000000
0!
0*
09
0>
0C
#644210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#644220000000
0!
0*
09
0>
0C
#644230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#644240000000
0!
0*
09
0>
0C
#644250000000
1!
1*
b10 6
19
1>
1C
b10 G
#644260000000
0!
0*
09
0>
0C
#644270000000
1!
1*
b11 6
19
1>
1C
b11 G
#644280000000
0!
0*
09
0>
0C
#644290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#644300000000
0!
0*
09
0>
0C
#644310000000
1!
1*
b101 6
19
1>
1C
b101 G
#644320000000
0!
0*
09
0>
0C
#644330000000
1!
1*
b110 6
19
1>
1C
b110 G
#644340000000
0!
0*
09
0>
0C
#644350000000
1!
1*
b111 6
19
1>
1C
b111 G
#644360000000
0!
0*
09
0>
0C
#644370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#644380000000
0!
0*
09
0>
0C
#644390000000
1!
1*
b1 6
19
1>
1C
b1 G
#644400000000
0!
0*
09
0>
0C
#644410000000
1!
1*
b10 6
19
1>
1C
b10 G
#644420000000
0!
0*
09
0>
0C
#644430000000
1!
1*
b11 6
19
1>
1C
b11 G
#644440000000
0!
0*
09
0>
0C
#644450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#644460000000
0!
0*
09
0>
0C
#644470000000
1!
1*
b101 6
19
1>
1C
b101 G
#644480000000
0!
0*
09
0>
0C
#644490000000
1!
1*
b110 6
19
1>
1C
b110 G
#644500000000
0!
0*
09
0>
0C
#644510000000
1!
1*
b111 6
19
1>
1C
b111 G
#644520000000
0!
0*
09
0>
0C
#644530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#644540000000
0!
0*
09
0>
0C
#644550000000
1!
1*
b1 6
19
1>
1C
b1 G
#644560000000
0!
0*
09
0>
0C
#644570000000
1!
1*
b10 6
19
1>
1C
b10 G
#644580000000
0!
0*
09
0>
0C
#644590000000
1!
1*
b11 6
19
1>
1C
b11 G
#644600000000
0!
0*
09
0>
0C
#644610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#644620000000
0!
0*
09
0>
0C
#644630000000
1!
1*
b101 6
19
1>
1C
b101 G
#644640000000
0!
0*
09
0>
0C
#644650000000
1!
1*
b110 6
19
1>
1C
b110 G
#644660000000
0!
0*
09
0>
0C
#644670000000
1!
1*
b111 6
19
1>
1C
b111 G
#644680000000
0!
1"
0*
1+
09
1:
0>
0C
#644690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#644700000000
0!
0*
09
0>
0C
#644710000000
1!
1*
b1 6
19
1>
1C
b1 G
#644720000000
0!
0*
09
0>
0C
#644730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#644740000000
0!
0*
09
0>
0C
#644750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#644760000000
0!
0*
09
0>
0C
#644770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#644780000000
0!
0*
09
0>
0C
#644790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#644800000000
0!
0#
0*
0,
09
0>
0?
0C
#644810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#644820000000
0!
0*
09
0>
0C
#644830000000
1!
1*
19
1>
1C
#644840000000
0!
0*
09
0>
0C
#644850000000
1!
1*
19
1>
1C
#644860000000
0!
0*
09
0>
0C
#644870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#644880000000
0!
0*
09
0>
0C
#644890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#644900000000
0!
0*
09
0>
0C
#644910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#644920000000
0!
0*
09
0>
0C
#644930000000
1!
1*
b10 6
19
1>
1C
b10 G
#644940000000
0!
0*
09
0>
0C
#644950000000
1!
1*
b11 6
19
1>
1C
b11 G
#644960000000
0!
0*
09
0>
0C
#644970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#644980000000
0!
0*
09
0>
0C
#644990000000
1!
1*
b101 6
19
1>
1C
b101 G
#645000000000
0!
0*
09
0>
0C
#645010000000
1!
1*
b110 6
19
1>
1C
b110 G
#645020000000
0!
0*
09
0>
0C
#645030000000
1!
1*
b111 6
19
1>
1C
b111 G
#645040000000
0!
0*
09
0>
0C
#645050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#645060000000
0!
0*
09
0>
0C
#645070000000
1!
1*
b1 6
19
1>
1C
b1 G
#645080000000
0!
0*
09
0>
0C
#645090000000
1!
1*
b10 6
19
1>
1C
b10 G
#645100000000
0!
0*
09
0>
0C
#645110000000
1!
1*
b11 6
19
1>
1C
b11 G
#645120000000
0!
0*
09
0>
0C
#645130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#645140000000
0!
0*
09
0>
0C
#645150000000
1!
1*
b101 6
19
1>
1C
b101 G
#645160000000
0!
0*
09
0>
0C
#645170000000
1!
1*
b110 6
19
1>
1C
b110 G
#645180000000
0!
0*
09
0>
0C
#645190000000
1!
1*
b111 6
19
1>
1C
b111 G
#645200000000
0!
0*
09
0>
0C
#645210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#645220000000
0!
0*
09
0>
0C
#645230000000
1!
1*
b1 6
19
1>
1C
b1 G
#645240000000
0!
0*
09
0>
0C
#645250000000
1!
1*
b10 6
19
1>
1C
b10 G
#645260000000
0!
0*
09
0>
0C
#645270000000
1!
1*
b11 6
19
1>
1C
b11 G
#645280000000
0!
0*
09
0>
0C
#645290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#645300000000
0!
0*
09
0>
0C
#645310000000
1!
1*
b101 6
19
1>
1C
b101 G
#645320000000
0!
0*
09
0>
0C
#645330000000
1!
1*
b110 6
19
1>
1C
b110 G
#645340000000
0!
0*
09
0>
0C
#645350000000
1!
1*
b111 6
19
1>
1C
b111 G
#645360000000
0!
1"
0*
1+
09
1:
0>
0C
#645370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#645380000000
0!
0*
09
0>
0C
#645390000000
1!
1*
b1 6
19
1>
1C
b1 G
#645400000000
0!
0*
09
0>
0C
#645410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#645420000000
0!
0*
09
0>
0C
#645430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#645440000000
0!
0*
09
0>
0C
#645450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#645460000000
0!
0*
09
0>
0C
#645470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#645480000000
0!
0#
0*
0,
09
0>
0?
0C
#645490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#645500000000
0!
0*
09
0>
0C
#645510000000
1!
1*
19
1>
1C
#645520000000
0!
0*
09
0>
0C
#645530000000
1!
1*
19
1>
1C
#645540000000
0!
0*
09
0>
0C
#645550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#645560000000
0!
0*
09
0>
0C
#645570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#645580000000
0!
0*
09
0>
0C
#645590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#645600000000
0!
0*
09
0>
0C
#645610000000
1!
1*
b10 6
19
1>
1C
b10 G
#645620000000
0!
0*
09
0>
0C
#645630000000
1!
1*
b11 6
19
1>
1C
b11 G
#645640000000
0!
0*
09
0>
0C
#645650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#645660000000
0!
0*
09
0>
0C
#645670000000
1!
1*
b101 6
19
1>
1C
b101 G
#645680000000
0!
0*
09
0>
0C
#645690000000
1!
1*
b110 6
19
1>
1C
b110 G
#645700000000
0!
0*
09
0>
0C
#645710000000
1!
1*
b111 6
19
1>
1C
b111 G
#645720000000
0!
0*
09
0>
0C
#645730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#645740000000
0!
0*
09
0>
0C
#645750000000
1!
1*
b1 6
19
1>
1C
b1 G
#645760000000
0!
0*
09
0>
0C
#645770000000
1!
1*
b10 6
19
1>
1C
b10 G
#645780000000
0!
0*
09
0>
0C
#645790000000
1!
1*
b11 6
19
1>
1C
b11 G
#645800000000
0!
0*
09
0>
0C
#645810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#645820000000
0!
0*
09
0>
0C
#645830000000
1!
1*
b101 6
19
1>
1C
b101 G
#645840000000
0!
0*
09
0>
0C
#645850000000
1!
1*
b110 6
19
1>
1C
b110 G
#645860000000
0!
0*
09
0>
0C
#645870000000
1!
1*
b111 6
19
1>
1C
b111 G
#645880000000
0!
0*
09
0>
0C
#645890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#645900000000
0!
0*
09
0>
0C
#645910000000
1!
1*
b1 6
19
1>
1C
b1 G
#645920000000
0!
0*
09
0>
0C
#645930000000
1!
1*
b10 6
19
1>
1C
b10 G
#645940000000
0!
0*
09
0>
0C
#645950000000
1!
1*
b11 6
19
1>
1C
b11 G
#645960000000
0!
0*
09
0>
0C
#645970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#645980000000
0!
0*
09
0>
0C
#645990000000
1!
1*
b101 6
19
1>
1C
b101 G
#646000000000
0!
0*
09
0>
0C
#646010000000
1!
1*
b110 6
19
1>
1C
b110 G
#646020000000
0!
0*
09
0>
0C
#646030000000
1!
1*
b111 6
19
1>
1C
b111 G
#646040000000
0!
1"
0*
1+
09
1:
0>
0C
#646050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#646060000000
0!
0*
09
0>
0C
#646070000000
1!
1*
b1 6
19
1>
1C
b1 G
#646080000000
0!
0*
09
0>
0C
#646090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#646100000000
0!
0*
09
0>
0C
#646110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#646120000000
0!
0*
09
0>
0C
#646130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#646140000000
0!
0*
09
0>
0C
#646150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#646160000000
0!
0#
0*
0,
09
0>
0?
0C
#646170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#646180000000
0!
0*
09
0>
0C
#646190000000
1!
1*
19
1>
1C
#646200000000
0!
0*
09
0>
0C
#646210000000
1!
1*
19
1>
1C
#646220000000
0!
0*
09
0>
0C
#646230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#646240000000
0!
0*
09
0>
0C
#646250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#646260000000
0!
0*
09
0>
0C
#646270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#646280000000
0!
0*
09
0>
0C
#646290000000
1!
1*
b10 6
19
1>
1C
b10 G
#646300000000
0!
0*
09
0>
0C
#646310000000
1!
1*
b11 6
19
1>
1C
b11 G
#646320000000
0!
0*
09
0>
0C
#646330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#646340000000
0!
0*
09
0>
0C
#646350000000
1!
1*
b101 6
19
1>
1C
b101 G
#646360000000
0!
0*
09
0>
0C
#646370000000
1!
1*
b110 6
19
1>
1C
b110 G
#646380000000
0!
0*
09
0>
0C
#646390000000
1!
1*
b111 6
19
1>
1C
b111 G
#646400000000
0!
0*
09
0>
0C
#646410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#646420000000
0!
0*
09
0>
0C
#646430000000
1!
1*
b1 6
19
1>
1C
b1 G
#646440000000
0!
0*
09
0>
0C
#646450000000
1!
1*
b10 6
19
1>
1C
b10 G
#646460000000
0!
0*
09
0>
0C
#646470000000
1!
1*
b11 6
19
1>
1C
b11 G
#646480000000
0!
0*
09
0>
0C
#646490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#646500000000
0!
0*
09
0>
0C
#646510000000
1!
1*
b101 6
19
1>
1C
b101 G
#646520000000
0!
0*
09
0>
0C
#646530000000
1!
1*
b110 6
19
1>
1C
b110 G
#646540000000
0!
0*
09
0>
0C
#646550000000
1!
1*
b111 6
19
1>
1C
b111 G
#646560000000
0!
0*
09
0>
0C
#646570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#646580000000
0!
0*
09
0>
0C
#646590000000
1!
1*
b1 6
19
1>
1C
b1 G
#646600000000
0!
0*
09
0>
0C
#646610000000
1!
1*
b10 6
19
1>
1C
b10 G
#646620000000
0!
0*
09
0>
0C
#646630000000
1!
1*
b11 6
19
1>
1C
b11 G
#646640000000
0!
0*
09
0>
0C
#646650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#646660000000
0!
0*
09
0>
0C
#646670000000
1!
1*
b101 6
19
1>
1C
b101 G
#646680000000
0!
0*
09
0>
0C
#646690000000
1!
1*
b110 6
19
1>
1C
b110 G
#646700000000
0!
0*
09
0>
0C
#646710000000
1!
1*
b111 6
19
1>
1C
b111 G
#646720000000
0!
1"
0*
1+
09
1:
0>
0C
#646730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#646740000000
0!
0*
09
0>
0C
#646750000000
1!
1*
b1 6
19
1>
1C
b1 G
#646760000000
0!
0*
09
0>
0C
#646770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#646780000000
0!
0*
09
0>
0C
#646790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#646800000000
0!
0*
09
0>
0C
#646810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#646820000000
0!
0*
09
0>
0C
#646830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#646840000000
0!
0#
0*
0,
09
0>
0?
0C
#646850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#646860000000
0!
0*
09
0>
0C
#646870000000
1!
1*
19
1>
1C
#646880000000
0!
0*
09
0>
0C
#646890000000
1!
1*
19
1>
1C
#646900000000
0!
0*
09
0>
0C
#646910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#646920000000
0!
0*
09
0>
0C
#646930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#646940000000
0!
0*
09
0>
0C
#646950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#646960000000
0!
0*
09
0>
0C
#646970000000
1!
1*
b10 6
19
1>
1C
b10 G
#646980000000
0!
0*
09
0>
0C
#646990000000
1!
1*
b11 6
19
1>
1C
b11 G
#647000000000
0!
0*
09
0>
0C
#647010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#647020000000
0!
0*
09
0>
0C
#647030000000
1!
1*
b101 6
19
1>
1C
b101 G
#647040000000
0!
0*
09
0>
0C
#647050000000
1!
1*
b110 6
19
1>
1C
b110 G
#647060000000
0!
0*
09
0>
0C
#647070000000
1!
1*
b111 6
19
1>
1C
b111 G
#647080000000
0!
0*
09
0>
0C
#647090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#647100000000
0!
0*
09
0>
0C
#647110000000
1!
1*
b1 6
19
1>
1C
b1 G
#647120000000
0!
0*
09
0>
0C
#647130000000
1!
1*
b10 6
19
1>
1C
b10 G
#647140000000
0!
0*
09
0>
0C
#647150000000
1!
1*
b11 6
19
1>
1C
b11 G
#647160000000
0!
0*
09
0>
0C
#647170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#647180000000
0!
0*
09
0>
0C
#647190000000
1!
1*
b101 6
19
1>
1C
b101 G
#647200000000
0!
0*
09
0>
0C
#647210000000
1!
1*
b110 6
19
1>
1C
b110 G
#647220000000
0!
0*
09
0>
0C
#647230000000
1!
1*
b111 6
19
1>
1C
b111 G
#647240000000
0!
0*
09
0>
0C
#647250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#647260000000
0!
0*
09
0>
0C
#647270000000
1!
1*
b1 6
19
1>
1C
b1 G
#647280000000
0!
0*
09
0>
0C
#647290000000
1!
1*
b10 6
19
1>
1C
b10 G
#647300000000
0!
0*
09
0>
0C
#647310000000
1!
1*
b11 6
19
1>
1C
b11 G
#647320000000
0!
0*
09
0>
0C
#647330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#647340000000
0!
0*
09
0>
0C
#647350000000
1!
1*
b101 6
19
1>
1C
b101 G
#647360000000
0!
0*
09
0>
0C
#647370000000
1!
1*
b110 6
19
1>
1C
b110 G
#647380000000
0!
0*
09
0>
0C
#647390000000
1!
1*
b111 6
19
1>
1C
b111 G
#647400000000
0!
1"
0*
1+
09
1:
0>
0C
#647410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#647420000000
0!
0*
09
0>
0C
#647430000000
1!
1*
b1 6
19
1>
1C
b1 G
#647440000000
0!
0*
09
0>
0C
#647450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#647460000000
0!
0*
09
0>
0C
#647470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#647480000000
0!
0*
09
0>
0C
#647490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#647500000000
0!
0*
09
0>
0C
#647510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#647520000000
0!
0#
0*
0,
09
0>
0?
0C
#647530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#647540000000
0!
0*
09
0>
0C
#647550000000
1!
1*
19
1>
1C
#647560000000
0!
0*
09
0>
0C
#647570000000
1!
1*
19
1>
1C
#647580000000
0!
0*
09
0>
0C
#647590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#647600000000
0!
0*
09
0>
0C
#647610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#647620000000
0!
0*
09
0>
0C
#647630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#647640000000
0!
0*
09
0>
0C
#647650000000
1!
1*
b10 6
19
1>
1C
b10 G
#647660000000
0!
0*
09
0>
0C
#647670000000
1!
1*
b11 6
19
1>
1C
b11 G
#647680000000
0!
0*
09
0>
0C
#647690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#647700000000
0!
0*
09
0>
0C
#647710000000
1!
1*
b101 6
19
1>
1C
b101 G
#647720000000
0!
0*
09
0>
0C
#647730000000
1!
1*
b110 6
19
1>
1C
b110 G
#647740000000
0!
0*
09
0>
0C
#647750000000
1!
1*
b111 6
19
1>
1C
b111 G
#647760000000
0!
0*
09
0>
0C
#647770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#647780000000
0!
0*
09
0>
0C
#647790000000
1!
1*
b1 6
19
1>
1C
b1 G
#647800000000
0!
0*
09
0>
0C
#647810000000
1!
1*
b10 6
19
1>
1C
b10 G
#647820000000
0!
0*
09
0>
0C
#647830000000
1!
1*
b11 6
19
1>
1C
b11 G
#647840000000
0!
0*
09
0>
0C
#647850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#647860000000
0!
0*
09
0>
0C
#647870000000
1!
1*
b101 6
19
1>
1C
b101 G
#647880000000
0!
0*
09
0>
0C
#647890000000
1!
1*
b110 6
19
1>
1C
b110 G
#647900000000
0!
0*
09
0>
0C
#647910000000
1!
1*
b111 6
19
1>
1C
b111 G
#647920000000
0!
0*
09
0>
0C
#647930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#647940000000
0!
0*
09
0>
0C
#647950000000
1!
1*
b1 6
19
1>
1C
b1 G
#647960000000
0!
0*
09
0>
0C
#647970000000
1!
1*
b10 6
19
1>
1C
b10 G
#647980000000
0!
0*
09
0>
0C
#647990000000
1!
1*
b11 6
19
1>
1C
b11 G
#648000000000
0!
0*
09
0>
0C
#648010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#648020000000
0!
0*
09
0>
0C
#648030000000
1!
1*
b101 6
19
1>
1C
b101 G
#648040000000
0!
0*
09
0>
0C
#648050000000
1!
1*
b110 6
19
1>
1C
b110 G
#648060000000
0!
0*
09
0>
0C
#648070000000
1!
1*
b111 6
19
1>
1C
b111 G
#648080000000
0!
1"
0*
1+
09
1:
0>
0C
#648090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#648100000000
0!
0*
09
0>
0C
#648110000000
1!
1*
b1 6
19
1>
1C
b1 G
#648120000000
0!
0*
09
0>
0C
#648130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#648140000000
0!
0*
09
0>
0C
#648150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#648160000000
0!
0*
09
0>
0C
#648170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#648180000000
0!
0*
09
0>
0C
#648190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#648200000000
0!
0#
0*
0,
09
0>
0?
0C
#648210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#648220000000
0!
0*
09
0>
0C
#648230000000
1!
1*
19
1>
1C
#648240000000
0!
0*
09
0>
0C
#648250000000
1!
1*
19
1>
1C
#648260000000
0!
0*
09
0>
0C
#648270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#648280000000
0!
0*
09
0>
0C
#648290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#648300000000
0!
0*
09
0>
0C
#648310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#648320000000
0!
0*
09
0>
0C
#648330000000
1!
1*
b10 6
19
1>
1C
b10 G
#648340000000
0!
0*
09
0>
0C
#648350000000
1!
1*
b11 6
19
1>
1C
b11 G
#648360000000
0!
0*
09
0>
0C
#648370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#648380000000
0!
0*
09
0>
0C
#648390000000
1!
1*
b101 6
19
1>
1C
b101 G
#648400000000
0!
0*
09
0>
0C
#648410000000
1!
1*
b110 6
19
1>
1C
b110 G
#648420000000
0!
0*
09
0>
0C
#648430000000
1!
1*
b111 6
19
1>
1C
b111 G
#648440000000
0!
0*
09
0>
0C
#648450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#648460000000
0!
0*
09
0>
0C
#648470000000
1!
1*
b1 6
19
1>
1C
b1 G
#648480000000
0!
0*
09
0>
0C
#648490000000
1!
1*
b10 6
19
1>
1C
b10 G
#648500000000
0!
0*
09
0>
0C
#648510000000
1!
1*
b11 6
19
1>
1C
b11 G
#648520000000
0!
0*
09
0>
0C
#648530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#648540000000
0!
0*
09
0>
0C
#648550000000
1!
1*
b101 6
19
1>
1C
b101 G
#648560000000
0!
0*
09
0>
0C
#648570000000
1!
1*
b110 6
19
1>
1C
b110 G
#648580000000
0!
0*
09
0>
0C
#648590000000
1!
1*
b111 6
19
1>
1C
b111 G
#648600000000
0!
0*
09
0>
0C
#648610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#648620000000
0!
0*
09
0>
0C
#648630000000
1!
1*
b1 6
19
1>
1C
b1 G
#648640000000
0!
0*
09
0>
0C
#648650000000
1!
1*
b10 6
19
1>
1C
b10 G
#648660000000
0!
0*
09
0>
0C
#648670000000
1!
1*
b11 6
19
1>
1C
b11 G
#648680000000
0!
0*
09
0>
0C
#648690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#648700000000
0!
0*
09
0>
0C
#648710000000
1!
1*
b101 6
19
1>
1C
b101 G
#648720000000
0!
0*
09
0>
0C
#648730000000
1!
1*
b110 6
19
1>
1C
b110 G
#648740000000
0!
0*
09
0>
0C
#648750000000
1!
1*
b111 6
19
1>
1C
b111 G
#648760000000
0!
1"
0*
1+
09
1:
0>
0C
#648770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#648780000000
0!
0*
09
0>
0C
#648790000000
1!
1*
b1 6
19
1>
1C
b1 G
#648800000000
0!
0*
09
0>
0C
#648810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#648820000000
0!
0*
09
0>
0C
#648830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#648840000000
0!
0*
09
0>
0C
#648850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#648860000000
0!
0*
09
0>
0C
#648870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#648880000000
0!
0#
0*
0,
09
0>
0?
0C
#648890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#648900000000
0!
0*
09
0>
0C
#648910000000
1!
1*
19
1>
1C
#648920000000
0!
0*
09
0>
0C
#648930000000
1!
1*
19
1>
1C
#648940000000
0!
0*
09
0>
0C
#648950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#648960000000
0!
0*
09
0>
0C
#648970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#648980000000
0!
0*
09
0>
0C
#648990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#649000000000
0!
0*
09
0>
0C
#649010000000
1!
1*
b10 6
19
1>
1C
b10 G
#649020000000
0!
0*
09
0>
0C
#649030000000
1!
1*
b11 6
19
1>
1C
b11 G
#649040000000
0!
0*
09
0>
0C
#649050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#649060000000
0!
0*
09
0>
0C
#649070000000
1!
1*
b101 6
19
1>
1C
b101 G
#649080000000
0!
0*
09
0>
0C
#649090000000
1!
1*
b110 6
19
1>
1C
b110 G
#649100000000
0!
0*
09
0>
0C
#649110000000
1!
1*
b111 6
19
1>
1C
b111 G
#649120000000
0!
0*
09
0>
0C
#649130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#649140000000
0!
0*
09
0>
0C
#649150000000
1!
1*
b1 6
19
1>
1C
b1 G
#649160000000
0!
0*
09
0>
0C
#649170000000
1!
1*
b10 6
19
1>
1C
b10 G
#649180000000
0!
0*
09
0>
0C
#649190000000
1!
1*
b11 6
19
1>
1C
b11 G
#649200000000
0!
0*
09
0>
0C
#649210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#649220000000
0!
0*
09
0>
0C
#649230000000
1!
1*
b101 6
19
1>
1C
b101 G
#649240000000
0!
0*
09
0>
0C
#649250000000
1!
1*
b110 6
19
1>
1C
b110 G
#649260000000
0!
0*
09
0>
0C
#649270000000
1!
1*
b111 6
19
1>
1C
b111 G
#649280000000
0!
0*
09
0>
0C
#649290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#649300000000
0!
0*
09
0>
0C
#649310000000
1!
1*
b1 6
19
1>
1C
b1 G
#649320000000
0!
0*
09
0>
0C
#649330000000
1!
1*
b10 6
19
1>
1C
b10 G
#649340000000
0!
0*
09
0>
0C
#649350000000
1!
1*
b11 6
19
1>
1C
b11 G
#649360000000
0!
0*
09
0>
0C
#649370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#649380000000
0!
0*
09
0>
0C
#649390000000
1!
1*
b101 6
19
1>
1C
b101 G
#649400000000
0!
0*
09
0>
0C
#649410000000
1!
1*
b110 6
19
1>
1C
b110 G
#649420000000
0!
0*
09
0>
0C
#649430000000
1!
1*
b111 6
19
1>
1C
b111 G
#649440000000
0!
1"
0*
1+
09
1:
0>
0C
#649450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#649460000000
0!
0*
09
0>
0C
#649470000000
1!
1*
b1 6
19
1>
1C
b1 G
#649480000000
0!
0*
09
0>
0C
#649490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#649500000000
0!
0*
09
0>
0C
#649510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#649520000000
0!
0*
09
0>
0C
#649530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#649540000000
0!
0*
09
0>
0C
#649550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#649560000000
0!
0#
0*
0,
09
0>
0?
0C
#649570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#649580000000
0!
0*
09
0>
0C
#649590000000
1!
1*
19
1>
1C
#649600000000
0!
0*
09
0>
0C
#649610000000
1!
1*
19
1>
1C
#649620000000
0!
0*
09
0>
0C
#649630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#649640000000
0!
0*
09
0>
0C
#649650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#649660000000
0!
0*
09
0>
0C
#649670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#649680000000
0!
0*
09
0>
0C
#649690000000
1!
1*
b10 6
19
1>
1C
b10 G
#649700000000
0!
0*
09
0>
0C
#649710000000
1!
1*
b11 6
19
1>
1C
b11 G
#649720000000
0!
0*
09
0>
0C
#649730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#649740000000
0!
0*
09
0>
0C
#649750000000
1!
1*
b101 6
19
1>
1C
b101 G
#649760000000
0!
0*
09
0>
0C
#649770000000
1!
1*
b110 6
19
1>
1C
b110 G
#649780000000
0!
0*
09
0>
0C
#649790000000
1!
1*
b111 6
19
1>
1C
b111 G
#649800000000
0!
0*
09
0>
0C
#649810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#649820000000
0!
0*
09
0>
0C
#649830000000
1!
1*
b1 6
19
1>
1C
b1 G
#649840000000
0!
0*
09
0>
0C
#649850000000
1!
1*
b10 6
19
1>
1C
b10 G
#649860000000
0!
0*
09
0>
0C
#649870000000
1!
1*
b11 6
19
1>
1C
b11 G
#649880000000
0!
0*
09
0>
0C
#649890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#649900000000
0!
0*
09
0>
0C
#649910000000
1!
1*
b101 6
19
1>
1C
b101 G
#649920000000
0!
0*
09
0>
0C
#649930000000
1!
1*
b110 6
19
1>
1C
b110 G
#649940000000
0!
0*
09
0>
0C
#649950000000
1!
1*
b111 6
19
1>
1C
b111 G
#649960000000
0!
0*
09
0>
0C
#649970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#649980000000
0!
0*
09
0>
0C
#649990000000
1!
1*
b1 6
19
1>
1C
b1 G
#650000000000
0!
0*
09
0>
0C
#650010000000
1!
1*
b10 6
19
1>
1C
b10 G
#650020000000
0!
0*
09
0>
0C
#650030000000
1!
1*
b11 6
19
1>
1C
b11 G
#650040000000
0!
0*
09
0>
0C
#650050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#650060000000
0!
0*
09
0>
0C
#650070000000
1!
1*
b101 6
19
1>
1C
b101 G
#650080000000
0!
0*
09
0>
0C
#650090000000
1!
1*
b110 6
19
1>
1C
b110 G
#650100000000
0!
0*
09
0>
0C
#650110000000
1!
1*
b111 6
19
1>
1C
b111 G
#650120000000
0!
1"
0*
1+
09
1:
0>
0C
#650130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#650140000000
0!
0*
09
0>
0C
#650150000000
1!
1*
b1 6
19
1>
1C
b1 G
#650160000000
0!
0*
09
0>
0C
#650170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#650180000000
0!
0*
09
0>
0C
#650190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#650200000000
0!
0*
09
0>
0C
#650210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#650220000000
0!
0*
09
0>
0C
#650230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#650240000000
0!
0#
0*
0,
09
0>
0?
0C
#650250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#650260000000
0!
0*
09
0>
0C
#650270000000
1!
1*
19
1>
1C
#650280000000
0!
0*
09
0>
0C
#650290000000
1!
1*
19
1>
1C
#650300000000
0!
0*
09
0>
0C
#650310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#650320000000
0!
0*
09
0>
0C
#650330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#650340000000
0!
0*
09
0>
0C
#650350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#650360000000
0!
0*
09
0>
0C
#650370000000
1!
1*
b10 6
19
1>
1C
b10 G
#650380000000
0!
0*
09
0>
0C
#650390000000
1!
1*
b11 6
19
1>
1C
b11 G
#650400000000
0!
0*
09
0>
0C
#650410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#650420000000
0!
0*
09
0>
0C
#650430000000
1!
1*
b101 6
19
1>
1C
b101 G
#650440000000
0!
0*
09
0>
0C
#650450000000
1!
1*
b110 6
19
1>
1C
b110 G
#650460000000
0!
0*
09
0>
0C
#650470000000
1!
1*
b111 6
19
1>
1C
b111 G
#650480000000
0!
0*
09
0>
0C
#650490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#650500000000
0!
0*
09
0>
0C
#650510000000
1!
1*
b1 6
19
1>
1C
b1 G
#650520000000
0!
0*
09
0>
0C
#650530000000
1!
1*
b10 6
19
1>
1C
b10 G
#650540000000
0!
0*
09
0>
0C
#650550000000
1!
1*
b11 6
19
1>
1C
b11 G
#650560000000
0!
0*
09
0>
0C
#650570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#650580000000
0!
0*
09
0>
0C
#650590000000
1!
1*
b101 6
19
1>
1C
b101 G
#650600000000
0!
0*
09
0>
0C
#650610000000
1!
1*
b110 6
19
1>
1C
b110 G
#650620000000
0!
0*
09
0>
0C
#650630000000
1!
1*
b111 6
19
1>
1C
b111 G
#650640000000
0!
0*
09
0>
0C
#650650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#650660000000
0!
0*
09
0>
0C
#650670000000
1!
1*
b1 6
19
1>
1C
b1 G
#650680000000
0!
0*
09
0>
0C
#650690000000
1!
1*
b10 6
19
1>
1C
b10 G
#650700000000
0!
0*
09
0>
0C
#650710000000
1!
1*
b11 6
19
1>
1C
b11 G
#650720000000
0!
0*
09
0>
0C
#650730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#650740000000
0!
0*
09
0>
0C
#650750000000
1!
1*
b101 6
19
1>
1C
b101 G
#650760000000
0!
0*
09
0>
0C
#650770000000
1!
1*
b110 6
19
1>
1C
b110 G
#650780000000
0!
0*
09
0>
0C
#650790000000
1!
1*
b111 6
19
1>
1C
b111 G
#650800000000
0!
1"
0*
1+
09
1:
0>
0C
#650810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#650820000000
0!
0*
09
0>
0C
#650830000000
1!
1*
b1 6
19
1>
1C
b1 G
#650840000000
0!
0*
09
0>
0C
#650850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#650860000000
0!
0*
09
0>
0C
#650870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#650880000000
0!
0*
09
0>
0C
#650890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#650900000000
0!
0*
09
0>
0C
#650910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#650920000000
0!
0#
0*
0,
09
0>
0?
0C
#650930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#650940000000
0!
0*
09
0>
0C
#650950000000
1!
1*
19
1>
1C
#650960000000
0!
0*
09
0>
0C
#650970000000
1!
1*
19
1>
1C
#650980000000
0!
0*
09
0>
0C
#650990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#651000000000
0!
0*
09
0>
0C
#651010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#651020000000
0!
0*
09
0>
0C
#651030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#651040000000
0!
0*
09
0>
0C
#651050000000
1!
1*
b10 6
19
1>
1C
b10 G
#651060000000
0!
0*
09
0>
0C
#651070000000
1!
1*
b11 6
19
1>
1C
b11 G
#651080000000
0!
0*
09
0>
0C
#651090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#651100000000
0!
0*
09
0>
0C
#651110000000
1!
1*
b101 6
19
1>
1C
b101 G
#651120000000
0!
0*
09
0>
0C
#651130000000
1!
1*
b110 6
19
1>
1C
b110 G
#651140000000
0!
0*
09
0>
0C
#651150000000
1!
1*
b111 6
19
1>
1C
b111 G
#651160000000
0!
0*
09
0>
0C
#651170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#651180000000
0!
0*
09
0>
0C
#651190000000
1!
1*
b1 6
19
1>
1C
b1 G
#651200000000
0!
0*
09
0>
0C
#651210000000
1!
1*
b10 6
19
1>
1C
b10 G
#651220000000
0!
0*
09
0>
0C
#651230000000
1!
1*
b11 6
19
1>
1C
b11 G
#651240000000
0!
0*
09
0>
0C
#651250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#651260000000
0!
0*
09
0>
0C
#651270000000
1!
1*
b101 6
19
1>
1C
b101 G
#651280000000
0!
0*
09
0>
0C
#651290000000
1!
1*
b110 6
19
1>
1C
b110 G
#651300000000
0!
0*
09
0>
0C
#651310000000
1!
1*
b111 6
19
1>
1C
b111 G
#651320000000
0!
0*
09
0>
0C
#651330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#651340000000
0!
0*
09
0>
0C
#651350000000
1!
1*
b1 6
19
1>
1C
b1 G
#651360000000
0!
0*
09
0>
0C
#651370000000
1!
1*
b10 6
19
1>
1C
b10 G
#651380000000
0!
0*
09
0>
0C
#651390000000
1!
1*
b11 6
19
1>
1C
b11 G
#651400000000
0!
0*
09
0>
0C
#651410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#651420000000
0!
0*
09
0>
0C
#651430000000
1!
1*
b101 6
19
1>
1C
b101 G
#651440000000
0!
0*
09
0>
0C
#651450000000
1!
1*
b110 6
19
1>
1C
b110 G
#651460000000
0!
0*
09
0>
0C
#651470000000
1!
1*
b111 6
19
1>
1C
b111 G
#651480000000
0!
1"
0*
1+
09
1:
0>
0C
#651490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#651500000000
0!
0*
09
0>
0C
#651510000000
1!
1*
b1 6
19
1>
1C
b1 G
#651520000000
0!
0*
09
0>
0C
#651530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#651540000000
0!
0*
09
0>
0C
#651550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#651560000000
0!
0*
09
0>
0C
#651570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#651580000000
0!
0*
09
0>
0C
#651590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#651600000000
0!
0#
0*
0,
09
0>
0?
0C
#651610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#651620000000
0!
0*
09
0>
0C
#651630000000
1!
1*
19
1>
1C
#651640000000
0!
0*
09
0>
0C
#651650000000
1!
1*
19
1>
1C
#651660000000
0!
0*
09
0>
0C
#651670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#651680000000
0!
0*
09
0>
0C
#651690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#651700000000
0!
0*
09
0>
0C
#651710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#651720000000
0!
0*
09
0>
0C
#651730000000
1!
1*
b10 6
19
1>
1C
b10 G
#651740000000
0!
0*
09
0>
0C
#651750000000
1!
1*
b11 6
19
1>
1C
b11 G
#651760000000
0!
0*
09
0>
0C
#651770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#651780000000
0!
0*
09
0>
0C
#651790000000
1!
1*
b101 6
19
1>
1C
b101 G
#651800000000
0!
0*
09
0>
0C
#651810000000
1!
1*
b110 6
19
1>
1C
b110 G
#651820000000
0!
0*
09
0>
0C
#651830000000
1!
1*
b111 6
19
1>
1C
b111 G
#651840000000
0!
0*
09
0>
0C
#651850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#651860000000
0!
0*
09
0>
0C
#651870000000
1!
1*
b1 6
19
1>
1C
b1 G
#651880000000
0!
0*
09
0>
0C
#651890000000
1!
1*
b10 6
19
1>
1C
b10 G
#651900000000
0!
0*
09
0>
0C
#651910000000
1!
1*
b11 6
19
1>
1C
b11 G
#651920000000
0!
0*
09
0>
0C
#651930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#651940000000
0!
0*
09
0>
0C
#651950000000
1!
1*
b101 6
19
1>
1C
b101 G
#651960000000
0!
0*
09
0>
0C
#651970000000
1!
1*
b110 6
19
1>
1C
b110 G
#651980000000
0!
0*
09
0>
0C
#651990000000
1!
1*
b111 6
19
1>
1C
b111 G
#652000000000
0!
0*
09
0>
0C
#652010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#652020000000
0!
0*
09
0>
0C
#652030000000
1!
1*
b1 6
19
1>
1C
b1 G
#652040000000
0!
0*
09
0>
0C
#652050000000
1!
1*
b10 6
19
1>
1C
b10 G
#652060000000
0!
0*
09
0>
0C
#652070000000
1!
1*
b11 6
19
1>
1C
b11 G
#652080000000
0!
0*
09
0>
0C
#652090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#652100000000
0!
0*
09
0>
0C
#652110000000
1!
1*
b101 6
19
1>
1C
b101 G
#652120000000
0!
0*
09
0>
0C
#652130000000
1!
1*
b110 6
19
1>
1C
b110 G
#652140000000
0!
0*
09
0>
0C
#652150000000
1!
1*
b111 6
19
1>
1C
b111 G
#652160000000
0!
1"
0*
1+
09
1:
0>
0C
#652170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#652180000000
0!
0*
09
0>
0C
#652190000000
1!
1*
b1 6
19
1>
1C
b1 G
#652200000000
0!
0*
09
0>
0C
#652210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#652220000000
0!
0*
09
0>
0C
#652230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#652240000000
0!
0*
09
0>
0C
#652250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#652260000000
0!
0*
09
0>
0C
#652270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#652280000000
0!
0#
0*
0,
09
0>
0?
0C
#652290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#652300000000
0!
0*
09
0>
0C
#652310000000
1!
1*
19
1>
1C
#652320000000
0!
0*
09
0>
0C
#652330000000
1!
1*
19
1>
1C
#652340000000
0!
0*
09
0>
0C
#652350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#652360000000
0!
0*
09
0>
0C
#652370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#652380000000
0!
0*
09
0>
0C
#652390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#652400000000
0!
0*
09
0>
0C
#652410000000
1!
1*
b10 6
19
1>
1C
b10 G
#652420000000
0!
0*
09
0>
0C
#652430000000
1!
1*
b11 6
19
1>
1C
b11 G
#652440000000
0!
0*
09
0>
0C
#652450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#652460000000
0!
0*
09
0>
0C
#652470000000
1!
1*
b101 6
19
1>
1C
b101 G
#652480000000
0!
0*
09
0>
0C
#652490000000
1!
1*
b110 6
19
1>
1C
b110 G
#652500000000
0!
0*
09
0>
0C
#652510000000
1!
1*
b111 6
19
1>
1C
b111 G
#652520000000
0!
0*
09
0>
0C
#652530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#652540000000
0!
0*
09
0>
0C
#652550000000
1!
1*
b1 6
19
1>
1C
b1 G
#652560000000
0!
0*
09
0>
0C
#652570000000
1!
1*
b10 6
19
1>
1C
b10 G
#652580000000
0!
0*
09
0>
0C
#652590000000
1!
1*
b11 6
19
1>
1C
b11 G
#652600000000
0!
0*
09
0>
0C
#652610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#652620000000
0!
0*
09
0>
0C
#652630000000
1!
1*
b101 6
19
1>
1C
b101 G
#652640000000
0!
0*
09
0>
0C
#652650000000
1!
1*
b110 6
19
1>
1C
b110 G
#652660000000
0!
0*
09
0>
0C
#652670000000
1!
1*
b111 6
19
1>
1C
b111 G
#652680000000
0!
0*
09
0>
0C
#652690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#652700000000
0!
0*
09
0>
0C
#652710000000
1!
1*
b1 6
19
1>
1C
b1 G
#652720000000
0!
0*
09
0>
0C
#652730000000
1!
1*
b10 6
19
1>
1C
b10 G
#652740000000
0!
0*
09
0>
0C
#652750000000
1!
1*
b11 6
19
1>
1C
b11 G
#652760000000
0!
0*
09
0>
0C
#652770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#652780000000
0!
0*
09
0>
0C
#652790000000
1!
1*
b101 6
19
1>
1C
b101 G
#652800000000
0!
0*
09
0>
0C
#652810000000
1!
1*
b110 6
19
1>
1C
b110 G
#652820000000
0!
0*
09
0>
0C
#652830000000
1!
1*
b111 6
19
1>
1C
b111 G
#652840000000
0!
1"
0*
1+
09
1:
0>
0C
#652850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#652860000000
0!
0*
09
0>
0C
#652870000000
1!
1*
b1 6
19
1>
1C
b1 G
#652880000000
0!
0*
09
0>
0C
#652890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#652900000000
0!
0*
09
0>
0C
#652910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#652920000000
0!
0*
09
0>
0C
#652930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#652940000000
0!
0*
09
0>
0C
#652950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#652960000000
0!
0#
0*
0,
09
0>
0?
0C
#652970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#652980000000
0!
0*
09
0>
0C
#652990000000
1!
1*
19
1>
1C
#653000000000
0!
0*
09
0>
0C
#653010000000
1!
1*
19
1>
1C
#653020000000
0!
0*
09
0>
0C
#653030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#653040000000
0!
0*
09
0>
0C
#653050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#653060000000
0!
0*
09
0>
0C
#653070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#653080000000
0!
0*
09
0>
0C
#653090000000
1!
1*
b10 6
19
1>
1C
b10 G
#653100000000
0!
0*
09
0>
0C
#653110000000
1!
1*
b11 6
19
1>
1C
b11 G
#653120000000
0!
0*
09
0>
0C
#653130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#653140000000
0!
0*
09
0>
0C
#653150000000
1!
1*
b101 6
19
1>
1C
b101 G
#653160000000
0!
0*
09
0>
0C
#653170000000
1!
1*
b110 6
19
1>
1C
b110 G
#653180000000
0!
0*
09
0>
0C
#653190000000
1!
1*
b111 6
19
1>
1C
b111 G
#653200000000
0!
0*
09
0>
0C
#653210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#653220000000
0!
0*
09
0>
0C
#653230000000
1!
1*
b1 6
19
1>
1C
b1 G
#653240000000
0!
0*
09
0>
0C
#653250000000
1!
1*
b10 6
19
1>
1C
b10 G
#653260000000
0!
0*
09
0>
0C
#653270000000
1!
1*
b11 6
19
1>
1C
b11 G
#653280000000
0!
0*
09
0>
0C
#653290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#653300000000
0!
0*
09
0>
0C
#653310000000
1!
1*
b101 6
19
1>
1C
b101 G
#653320000000
0!
0*
09
0>
0C
#653330000000
1!
1*
b110 6
19
1>
1C
b110 G
#653340000000
0!
0*
09
0>
0C
#653350000000
1!
1*
b111 6
19
1>
1C
b111 G
#653360000000
0!
0*
09
0>
0C
#653370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#653380000000
0!
0*
09
0>
0C
#653390000000
1!
1*
b1 6
19
1>
1C
b1 G
#653400000000
0!
0*
09
0>
0C
#653410000000
1!
1*
b10 6
19
1>
1C
b10 G
#653420000000
0!
0*
09
0>
0C
#653430000000
1!
1*
b11 6
19
1>
1C
b11 G
#653440000000
0!
0*
09
0>
0C
#653450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#653460000000
0!
0*
09
0>
0C
#653470000000
1!
1*
b101 6
19
1>
1C
b101 G
#653480000000
0!
0*
09
0>
0C
#653490000000
1!
1*
b110 6
19
1>
1C
b110 G
#653500000000
0!
0*
09
0>
0C
#653510000000
1!
1*
b111 6
19
1>
1C
b111 G
#653520000000
0!
1"
0*
1+
09
1:
0>
0C
#653530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#653540000000
0!
0*
09
0>
0C
#653550000000
1!
1*
b1 6
19
1>
1C
b1 G
#653560000000
0!
0*
09
0>
0C
#653570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#653580000000
0!
0*
09
0>
0C
#653590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#653600000000
0!
0*
09
0>
0C
#653610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#653620000000
0!
0*
09
0>
0C
#653630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#653640000000
0!
0#
0*
0,
09
0>
0?
0C
#653650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#653660000000
0!
0*
09
0>
0C
#653670000000
1!
1*
19
1>
1C
#653680000000
0!
0*
09
0>
0C
#653690000000
1!
1*
19
1>
1C
#653700000000
0!
0*
09
0>
0C
#653710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#653720000000
0!
0*
09
0>
0C
#653730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#653740000000
0!
0*
09
0>
0C
#653750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#653760000000
0!
0*
09
0>
0C
#653770000000
1!
1*
b10 6
19
1>
1C
b10 G
#653780000000
0!
0*
09
0>
0C
#653790000000
1!
1*
b11 6
19
1>
1C
b11 G
#653800000000
0!
0*
09
0>
0C
#653810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#653820000000
0!
0*
09
0>
0C
#653830000000
1!
1*
b101 6
19
1>
1C
b101 G
#653840000000
0!
0*
09
0>
0C
#653850000000
1!
1*
b110 6
19
1>
1C
b110 G
#653860000000
0!
0*
09
0>
0C
#653870000000
1!
1*
b111 6
19
1>
1C
b111 G
#653880000000
0!
0*
09
0>
0C
#653890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#653900000000
0!
0*
09
0>
0C
#653910000000
1!
1*
b1 6
19
1>
1C
b1 G
#653920000000
0!
0*
09
0>
0C
#653930000000
1!
1*
b10 6
19
1>
1C
b10 G
#653940000000
0!
0*
09
0>
0C
#653950000000
1!
1*
b11 6
19
1>
1C
b11 G
#653960000000
0!
0*
09
0>
0C
#653970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#653980000000
0!
0*
09
0>
0C
#653990000000
1!
1*
b101 6
19
1>
1C
b101 G
#654000000000
0!
0*
09
0>
0C
#654010000000
1!
1*
b110 6
19
1>
1C
b110 G
#654020000000
0!
0*
09
0>
0C
#654030000000
1!
1*
b111 6
19
1>
1C
b111 G
#654040000000
0!
0*
09
0>
0C
#654050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#654060000000
0!
0*
09
0>
0C
#654070000000
1!
1*
b1 6
19
1>
1C
b1 G
#654080000000
0!
0*
09
0>
0C
#654090000000
1!
1*
b10 6
19
1>
1C
b10 G
#654100000000
0!
0*
09
0>
0C
#654110000000
1!
1*
b11 6
19
1>
1C
b11 G
#654120000000
0!
0*
09
0>
0C
#654130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#654140000000
0!
0*
09
0>
0C
#654150000000
1!
1*
b101 6
19
1>
1C
b101 G
#654160000000
0!
0*
09
0>
0C
#654170000000
1!
1*
b110 6
19
1>
1C
b110 G
#654180000000
0!
0*
09
0>
0C
#654190000000
1!
1*
b111 6
19
1>
1C
b111 G
#654200000000
0!
1"
0*
1+
09
1:
0>
0C
#654210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#654220000000
0!
0*
09
0>
0C
#654230000000
1!
1*
b1 6
19
1>
1C
b1 G
#654240000000
0!
0*
09
0>
0C
#654250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#654260000000
0!
0*
09
0>
0C
#654270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#654280000000
0!
0*
09
0>
0C
#654290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#654300000000
0!
0*
09
0>
0C
#654310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#654320000000
0!
0#
0*
0,
09
0>
0?
0C
#654330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#654340000000
0!
0*
09
0>
0C
#654350000000
1!
1*
19
1>
1C
#654360000000
0!
0*
09
0>
0C
#654370000000
1!
1*
19
1>
1C
#654380000000
0!
0*
09
0>
0C
#654390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#654400000000
0!
0*
09
0>
0C
#654410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#654420000000
0!
0*
09
0>
0C
#654430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#654440000000
0!
0*
09
0>
0C
#654450000000
1!
1*
b10 6
19
1>
1C
b10 G
#654460000000
0!
0*
09
0>
0C
#654470000000
1!
1*
b11 6
19
1>
1C
b11 G
#654480000000
0!
0*
09
0>
0C
#654490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#654500000000
0!
0*
09
0>
0C
#654510000000
1!
1*
b101 6
19
1>
1C
b101 G
#654520000000
0!
0*
09
0>
0C
#654530000000
1!
1*
b110 6
19
1>
1C
b110 G
#654540000000
0!
0*
09
0>
0C
#654550000000
1!
1*
b111 6
19
1>
1C
b111 G
#654560000000
0!
0*
09
0>
0C
#654570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#654580000000
0!
0*
09
0>
0C
#654590000000
1!
1*
b1 6
19
1>
1C
b1 G
#654600000000
0!
0*
09
0>
0C
#654610000000
1!
1*
b10 6
19
1>
1C
b10 G
#654620000000
0!
0*
09
0>
0C
#654630000000
1!
1*
b11 6
19
1>
1C
b11 G
#654640000000
0!
0*
09
0>
0C
#654650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#654660000000
0!
0*
09
0>
0C
#654670000000
1!
1*
b101 6
19
1>
1C
b101 G
#654680000000
0!
0*
09
0>
0C
#654690000000
1!
1*
b110 6
19
1>
1C
b110 G
#654700000000
0!
0*
09
0>
0C
#654710000000
1!
1*
b111 6
19
1>
1C
b111 G
#654720000000
0!
0*
09
0>
0C
#654730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#654740000000
0!
0*
09
0>
0C
#654750000000
1!
1*
b1 6
19
1>
1C
b1 G
#654760000000
0!
0*
09
0>
0C
#654770000000
1!
1*
b10 6
19
1>
1C
b10 G
#654780000000
0!
0*
09
0>
0C
#654790000000
1!
1*
b11 6
19
1>
1C
b11 G
#654800000000
0!
0*
09
0>
0C
#654810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#654820000000
0!
0*
09
0>
0C
#654830000000
1!
1*
b101 6
19
1>
1C
b101 G
#654840000000
0!
0*
09
0>
0C
#654850000000
1!
1*
b110 6
19
1>
1C
b110 G
#654860000000
0!
0*
09
0>
0C
#654870000000
1!
1*
b111 6
19
1>
1C
b111 G
#654880000000
0!
1"
0*
1+
09
1:
0>
0C
#654890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#654900000000
0!
0*
09
0>
0C
#654910000000
1!
1*
b1 6
19
1>
1C
b1 G
#654920000000
0!
0*
09
0>
0C
#654930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#654940000000
0!
0*
09
0>
0C
#654950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#654960000000
0!
0*
09
0>
0C
#654970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#654980000000
0!
0*
09
0>
0C
#654990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#655000000000
0!
0#
0*
0,
09
0>
0?
0C
#655010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#655020000000
0!
0*
09
0>
0C
#655030000000
1!
1*
19
1>
1C
#655040000000
0!
0*
09
0>
0C
#655050000000
1!
1*
19
1>
1C
#655060000000
0!
0*
09
0>
0C
#655070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#655080000000
0!
0*
09
0>
0C
#655090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#655100000000
0!
0*
09
0>
0C
#655110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#655120000000
0!
0*
09
0>
0C
#655130000000
1!
1*
b10 6
19
1>
1C
b10 G
#655140000000
0!
0*
09
0>
0C
#655150000000
1!
1*
b11 6
19
1>
1C
b11 G
#655160000000
0!
0*
09
0>
0C
#655170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#655180000000
0!
0*
09
0>
0C
#655190000000
1!
1*
b101 6
19
1>
1C
b101 G
#655200000000
0!
0*
09
0>
0C
#655210000000
1!
1*
b110 6
19
1>
1C
b110 G
#655220000000
0!
0*
09
0>
0C
#655230000000
1!
1*
b111 6
19
1>
1C
b111 G
#655240000000
0!
0*
09
0>
0C
#655250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#655260000000
0!
0*
09
0>
0C
#655270000000
1!
1*
b1 6
19
1>
1C
b1 G
#655280000000
0!
0*
09
0>
0C
#655290000000
1!
1*
b10 6
19
1>
1C
b10 G
#655300000000
0!
0*
09
0>
0C
#655310000000
1!
1*
b11 6
19
1>
1C
b11 G
#655320000000
0!
0*
09
0>
0C
#655330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#655340000000
0!
0*
09
0>
0C
#655350000000
1!
1*
b101 6
19
1>
1C
b101 G
#655360000000
0!
0*
09
0>
0C
#655370000000
1!
1*
b110 6
19
1>
1C
b110 G
#655380000000
0!
0*
09
0>
0C
#655390000000
1!
1*
b111 6
19
1>
1C
b111 G
#655400000000
0!
0*
09
0>
0C
#655410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#655420000000
0!
0*
09
0>
0C
#655430000000
1!
1*
b1 6
19
1>
1C
b1 G
#655440000000
0!
0*
09
0>
0C
#655450000000
1!
1*
b10 6
19
1>
1C
b10 G
#655460000000
0!
0*
09
0>
0C
#655470000000
1!
1*
b11 6
19
1>
1C
b11 G
#655480000000
0!
0*
09
0>
0C
#655490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#655500000000
0!
0*
09
0>
0C
#655510000000
1!
1*
b101 6
19
1>
1C
b101 G
#655520000000
0!
0*
09
0>
0C
#655530000000
1!
1*
b110 6
19
1>
1C
b110 G
#655540000000
0!
0*
09
0>
0C
#655550000000
1!
1*
b111 6
19
1>
1C
b111 G
#655560000000
0!
1"
0*
1+
09
1:
0>
0C
#655570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#655580000000
0!
0*
09
0>
0C
#655590000000
1!
1*
b1 6
19
1>
1C
b1 G
#655600000000
0!
0*
09
0>
0C
#655610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#655620000000
0!
0*
09
0>
0C
#655630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#655640000000
0!
0*
09
0>
0C
#655650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#655660000000
0!
0*
09
0>
0C
#655670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#655680000000
0!
0#
0*
0,
09
0>
0?
0C
#655690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#655700000000
0!
0*
09
0>
0C
#655710000000
1!
1*
19
1>
1C
#655720000000
0!
0*
09
0>
0C
#655730000000
1!
1*
19
1>
1C
#655740000000
0!
0*
09
0>
0C
#655750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#655760000000
0!
0*
09
0>
0C
#655770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#655780000000
0!
0*
09
0>
0C
#655790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#655800000000
0!
0*
09
0>
0C
#655810000000
1!
1*
b10 6
19
1>
1C
b10 G
#655820000000
0!
0*
09
0>
0C
#655830000000
1!
1*
b11 6
19
1>
1C
b11 G
#655840000000
0!
0*
09
0>
0C
#655850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#655860000000
0!
0*
09
0>
0C
#655870000000
1!
1*
b101 6
19
1>
1C
b101 G
#655880000000
0!
0*
09
0>
0C
#655890000000
1!
1*
b110 6
19
1>
1C
b110 G
#655900000000
0!
0*
09
0>
0C
#655910000000
1!
1*
b111 6
19
1>
1C
b111 G
#655920000000
0!
0*
09
0>
0C
#655930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#655940000000
0!
0*
09
0>
0C
#655950000000
1!
1*
b1 6
19
1>
1C
b1 G
#655960000000
0!
0*
09
0>
0C
#655970000000
1!
1*
b10 6
19
1>
1C
b10 G
#655980000000
0!
0*
09
0>
0C
#655990000000
1!
1*
b11 6
19
1>
1C
b11 G
#656000000000
0!
0*
09
0>
0C
#656010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#656020000000
0!
0*
09
0>
0C
#656030000000
1!
1*
b101 6
19
1>
1C
b101 G
#656040000000
0!
0*
09
0>
0C
#656050000000
1!
1*
b110 6
19
1>
1C
b110 G
#656060000000
0!
0*
09
0>
0C
#656070000000
1!
1*
b111 6
19
1>
1C
b111 G
#656080000000
0!
0*
09
0>
0C
#656090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#656100000000
0!
0*
09
0>
0C
#656110000000
1!
1*
b1 6
19
1>
1C
b1 G
#656120000000
0!
0*
09
0>
0C
#656130000000
1!
1*
b10 6
19
1>
1C
b10 G
#656140000000
0!
0*
09
0>
0C
#656150000000
1!
1*
b11 6
19
1>
1C
b11 G
#656160000000
0!
0*
09
0>
0C
#656170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#656180000000
0!
0*
09
0>
0C
#656190000000
1!
1*
b101 6
19
1>
1C
b101 G
#656200000000
0!
0*
09
0>
0C
#656210000000
1!
1*
b110 6
19
1>
1C
b110 G
#656220000000
0!
0*
09
0>
0C
#656230000000
1!
1*
b111 6
19
1>
1C
b111 G
#656240000000
0!
1"
0*
1+
09
1:
0>
0C
#656250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#656260000000
0!
0*
09
0>
0C
#656270000000
1!
1*
b1 6
19
1>
1C
b1 G
#656280000000
0!
0*
09
0>
0C
#656290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#656300000000
0!
0*
09
0>
0C
#656310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#656320000000
0!
0*
09
0>
0C
#656330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#656340000000
0!
0*
09
0>
0C
#656350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#656360000000
0!
0#
0*
0,
09
0>
0?
0C
#656370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#656380000000
0!
0*
09
0>
0C
#656390000000
1!
1*
19
1>
1C
#656400000000
0!
0*
09
0>
0C
#656410000000
1!
1*
19
1>
1C
#656420000000
0!
0*
09
0>
0C
#656430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#656440000000
0!
0*
09
0>
0C
#656450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#656460000000
0!
0*
09
0>
0C
#656470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#656480000000
0!
0*
09
0>
0C
#656490000000
1!
1*
b10 6
19
1>
1C
b10 G
#656500000000
0!
0*
09
0>
0C
#656510000000
1!
1*
b11 6
19
1>
1C
b11 G
#656520000000
0!
0*
09
0>
0C
#656530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#656540000000
0!
0*
09
0>
0C
#656550000000
1!
1*
b101 6
19
1>
1C
b101 G
#656560000000
0!
0*
09
0>
0C
#656570000000
1!
1*
b110 6
19
1>
1C
b110 G
#656580000000
0!
0*
09
0>
0C
#656590000000
1!
1*
b111 6
19
1>
1C
b111 G
#656600000000
0!
0*
09
0>
0C
#656610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#656620000000
0!
0*
09
0>
0C
#656630000000
1!
1*
b1 6
19
1>
1C
b1 G
#656640000000
0!
0*
09
0>
0C
#656650000000
1!
1*
b10 6
19
1>
1C
b10 G
#656660000000
0!
0*
09
0>
0C
#656670000000
1!
1*
b11 6
19
1>
1C
b11 G
#656680000000
0!
0*
09
0>
0C
#656690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#656700000000
0!
0*
09
0>
0C
#656710000000
1!
1*
b101 6
19
1>
1C
b101 G
#656720000000
0!
0*
09
0>
0C
#656730000000
1!
1*
b110 6
19
1>
1C
b110 G
#656740000000
0!
0*
09
0>
0C
#656750000000
1!
1*
b111 6
19
1>
1C
b111 G
#656760000000
0!
0*
09
0>
0C
#656770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#656780000000
0!
0*
09
0>
0C
#656790000000
1!
1*
b1 6
19
1>
1C
b1 G
#656800000000
0!
0*
09
0>
0C
#656810000000
1!
1*
b10 6
19
1>
1C
b10 G
#656820000000
0!
0*
09
0>
0C
#656830000000
1!
1*
b11 6
19
1>
1C
b11 G
#656840000000
0!
0*
09
0>
0C
#656850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#656860000000
0!
0*
09
0>
0C
#656870000000
1!
1*
b101 6
19
1>
1C
b101 G
#656880000000
0!
0*
09
0>
0C
#656890000000
1!
1*
b110 6
19
1>
1C
b110 G
#656900000000
0!
0*
09
0>
0C
#656910000000
1!
1*
b111 6
19
1>
1C
b111 G
#656920000000
0!
1"
0*
1+
09
1:
0>
0C
#656930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#656940000000
0!
0*
09
0>
0C
#656950000000
1!
1*
b1 6
19
1>
1C
b1 G
#656960000000
0!
0*
09
0>
0C
#656970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#656980000000
0!
0*
09
0>
0C
#656990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#657000000000
0!
0*
09
0>
0C
#657010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#657020000000
0!
0*
09
0>
0C
#657030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#657040000000
0!
0#
0*
0,
09
0>
0?
0C
#657050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#657060000000
0!
0*
09
0>
0C
#657070000000
1!
1*
19
1>
1C
#657080000000
0!
0*
09
0>
0C
#657090000000
1!
1*
19
1>
1C
#657100000000
0!
0*
09
0>
0C
#657110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#657120000000
0!
0*
09
0>
0C
#657130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#657140000000
0!
0*
09
0>
0C
#657150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#657160000000
0!
0*
09
0>
0C
#657170000000
1!
1*
b10 6
19
1>
1C
b10 G
#657180000000
0!
0*
09
0>
0C
#657190000000
1!
1*
b11 6
19
1>
1C
b11 G
#657200000000
0!
0*
09
0>
0C
#657210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#657220000000
0!
0*
09
0>
0C
#657230000000
1!
1*
b101 6
19
1>
1C
b101 G
#657240000000
0!
0*
09
0>
0C
#657250000000
1!
1*
b110 6
19
1>
1C
b110 G
#657260000000
0!
0*
09
0>
0C
#657270000000
1!
1*
b111 6
19
1>
1C
b111 G
#657280000000
0!
0*
09
0>
0C
#657290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#657300000000
0!
0*
09
0>
0C
#657310000000
1!
1*
b1 6
19
1>
1C
b1 G
#657320000000
0!
0*
09
0>
0C
#657330000000
1!
1*
b10 6
19
1>
1C
b10 G
#657340000000
0!
0*
09
0>
0C
#657350000000
1!
1*
b11 6
19
1>
1C
b11 G
#657360000000
0!
0*
09
0>
0C
#657370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#657380000000
0!
0*
09
0>
0C
#657390000000
1!
1*
b101 6
19
1>
1C
b101 G
#657400000000
0!
0*
09
0>
0C
#657410000000
1!
1*
b110 6
19
1>
1C
b110 G
#657420000000
0!
0*
09
0>
0C
#657430000000
1!
1*
b111 6
19
1>
1C
b111 G
#657440000000
0!
0*
09
0>
0C
#657450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#657460000000
0!
0*
09
0>
0C
#657470000000
1!
1*
b1 6
19
1>
1C
b1 G
#657480000000
0!
0*
09
0>
0C
#657490000000
1!
1*
b10 6
19
1>
1C
b10 G
#657500000000
0!
0*
09
0>
0C
#657510000000
1!
1*
b11 6
19
1>
1C
b11 G
#657520000000
0!
0*
09
0>
0C
#657530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#657540000000
0!
0*
09
0>
0C
#657550000000
1!
1*
b101 6
19
1>
1C
b101 G
#657560000000
0!
0*
09
0>
0C
#657570000000
1!
1*
b110 6
19
1>
1C
b110 G
#657580000000
0!
0*
09
0>
0C
#657590000000
1!
1*
b111 6
19
1>
1C
b111 G
#657600000000
0!
1"
0*
1+
09
1:
0>
0C
#657610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#657620000000
0!
0*
09
0>
0C
#657630000000
1!
1*
b1 6
19
1>
1C
b1 G
#657640000000
0!
0*
09
0>
0C
#657650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#657660000000
0!
0*
09
0>
0C
#657670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#657680000000
0!
0*
09
0>
0C
#657690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#657700000000
0!
0*
09
0>
0C
#657710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#657720000000
0!
0#
0*
0,
09
0>
0?
0C
#657730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#657740000000
0!
0*
09
0>
0C
#657750000000
1!
1*
19
1>
1C
#657760000000
0!
0*
09
0>
0C
#657770000000
1!
1*
19
1>
1C
#657780000000
0!
0*
09
0>
0C
#657790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#657800000000
0!
0*
09
0>
0C
#657810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#657820000000
0!
0*
09
0>
0C
#657830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#657840000000
0!
0*
09
0>
0C
#657850000000
1!
1*
b10 6
19
1>
1C
b10 G
#657860000000
0!
0*
09
0>
0C
#657870000000
1!
1*
b11 6
19
1>
1C
b11 G
#657880000000
0!
0*
09
0>
0C
#657890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#657900000000
0!
0*
09
0>
0C
#657910000000
1!
1*
b101 6
19
1>
1C
b101 G
#657920000000
0!
0*
09
0>
0C
#657930000000
1!
1*
b110 6
19
1>
1C
b110 G
#657940000000
0!
0*
09
0>
0C
#657950000000
1!
1*
b111 6
19
1>
1C
b111 G
#657960000000
0!
0*
09
0>
0C
#657970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#657980000000
0!
0*
09
0>
0C
#657990000000
1!
1*
b1 6
19
1>
1C
b1 G
#658000000000
0!
0*
09
0>
0C
#658010000000
1!
1*
b10 6
19
1>
1C
b10 G
#658020000000
0!
0*
09
0>
0C
#658030000000
1!
1*
b11 6
19
1>
1C
b11 G
#658040000000
0!
0*
09
0>
0C
#658050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#658060000000
0!
0*
09
0>
0C
#658070000000
1!
1*
b101 6
19
1>
1C
b101 G
#658080000000
0!
0*
09
0>
0C
#658090000000
1!
1*
b110 6
19
1>
1C
b110 G
#658100000000
0!
0*
09
0>
0C
#658110000000
1!
1*
b111 6
19
1>
1C
b111 G
#658120000000
0!
0*
09
0>
0C
#658130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#658140000000
0!
0*
09
0>
0C
#658150000000
1!
1*
b1 6
19
1>
1C
b1 G
#658160000000
0!
0*
09
0>
0C
#658170000000
1!
1*
b10 6
19
1>
1C
b10 G
#658180000000
0!
0*
09
0>
0C
#658190000000
1!
1*
b11 6
19
1>
1C
b11 G
#658200000000
0!
0*
09
0>
0C
#658210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#658220000000
0!
0*
09
0>
0C
#658230000000
1!
1*
b101 6
19
1>
1C
b101 G
#658240000000
0!
0*
09
0>
0C
#658250000000
1!
1*
b110 6
19
1>
1C
b110 G
#658260000000
0!
0*
09
0>
0C
#658270000000
1!
1*
b111 6
19
1>
1C
b111 G
#658280000000
0!
1"
0*
1+
09
1:
0>
0C
#658290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#658300000000
0!
0*
09
0>
0C
#658310000000
1!
1*
b1 6
19
1>
1C
b1 G
#658320000000
0!
0*
09
0>
0C
#658330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#658340000000
0!
0*
09
0>
0C
#658350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#658360000000
0!
0*
09
0>
0C
#658370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#658380000000
0!
0*
09
0>
0C
#658390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#658400000000
0!
0#
0*
0,
09
0>
0?
0C
#658410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#658420000000
0!
0*
09
0>
0C
#658430000000
1!
1*
19
1>
1C
#658440000000
0!
0*
09
0>
0C
#658450000000
1!
1*
19
1>
1C
#658460000000
0!
0*
09
0>
0C
#658470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#658480000000
0!
0*
09
0>
0C
#658490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#658500000000
0!
0*
09
0>
0C
#658510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#658520000000
0!
0*
09
0>
0C
#658530000000
1!
1*
b10 6
19
1>
1C
b10 G
#658540000000
0!
0*
09
0>
0C
#658550000000
1!
1*
b11 6
19
1>
1C
b11 G
#658560000000
0!
0*
09
0>
0C
#658570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#658580000000
0!
0*
09
0>
0C
#658590000000
1!
1*
b101 6
19
1>
1C
b101 G
#658600000000
0!
0*
09
0>
0C
#658610000000
1!
1*
b110 6
19
1>
1C
b110 G
#658620000000
0!
0*
09
0>
0C
#658630000000
1!
1*
b111 6
19
1>
1C
b111 G
#658640000000
0!
0*
09
0>
0C
#658650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#658660000000
0!
0*
09
0>
0C
#658670000000
1!
1*
b1 6
19
1>
1C
b1 G
#658680000000
0!
0*
09
0>
0C
#658690000000
1!
1*
b10 6
19
1>
1C
b10 G
#658700000000
0!
0*
09
0>
0C
#658710000000
1!
1*
b11 6
19
1>
1C
b11 G
#658720000000
0!
0*
09
0>
0C
#658730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#658740000000
0!
0*
09
0>
0C
#658750000000
1!
1*
b101 6
19
1>
1C
b101 G
#658760000000
0!
0*
09
0>
0C
#658770000000
1!
1*
b110 6
19
1>
1C
b110 G
#658780000000
0!
0*
09
0>
0C
#658790000000
1!
1*
b111 6
19
1>
1C
b111 G
#658800000000
0!
0*
09
0>
0C
#658810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#658820000000
0!
0*
09
0>
0C
#658830000000
1!
1*
b1 6
19
1>
1C
b1 G
#658840000000
0!
0*
09
0>
0C
#658850000000
1!
1*
b10 6
19
1>
1C
b10 G
#658860000000
0!
0*
09
0>
0C
#658870000000
1!
1*
b11 6
19
1>
1C
b11 G
#658880000000
0!
0*
09
0>
0C
#658890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#658900000000
0!
0*
09
0>
0C
#658910000000
1!
1*
b101 6
19
1>
1C
b101 G
#658920000000
0!
0*
09
0>
0C
#658930000000
1!
1*
b110 6
19
1>
1C
b110 G
#658940000000
0!
0*
09
0>
0C
#658950000000
1!
1*
b111 6
19
1>
1C
b111 G
#658960000000
0!
1"
0*
1+
09
1:
0>
0C
#658970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#658980000000
0!
0*
09
0>
0C
#658990000000
1!
1*
b1 6
19
1>
1C
b1 G
#659000000000
0!
0*
09
0>
0C
#659010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#659020000000
0!
0*
09
0>
0C
#659030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#659040000000
0!
0*
09
0>
0C
#659050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#659060000000
0!
0*
09
0>
0C
#659070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#659080000000
0!
0#
0*
0,
09
0>
0?
0C
#659090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#659100000000
0!
0*
09
0>
0C
#659110000000
1!
1*
19
1>
1C
#659120000000
0!
0*
09
0>
0C
#659130000000
1!
1*
19
1>
1C
#659140000000
0!
0*
09
0>
0C
#659150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#659160000000
0!
0*
09
0>
0C
#659170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#659180000000
0!
0*
09
0>
0C
#659190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#659200000000
0!
0*
09
0>
0C
#659210000000
1!
1*
b10 6
19
1>
1C
b10 G
#659220000000
0!
0*
09
0>
0C
#659230000000
1!
1*
b11 6
19
1>
1C
b11 G
#659240000000
0!
0*
09
0>
0C
#659250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#659260000000
0!
0*
09
0>
0C
#659270000000
1!
1*
b101 6
19
1>
1C
b101 G
#659280000000
0!
0*
09
0>
0C
#659290000000
1!
1*
b110 6
19
1>
1C
b110 G
#659300000000
0!
0*
09
0>
0C
#659310000000
1!
1*
b111 6
19
1>
1C
b111 G
#659320000000
0!
0*
09
0>
0C
#659330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#659340000000
0!
0*
09
0>
0C
#659350000000
1!
1*
b1 6
19
1>
1C
b1 G
#659360000000
0!
0*
09
0>
0C
#659370000000
1!
1*
b10 6
19
1>
1C
b10 G
#659380000000
0!
0*
09
0>
0C
#659390000000
1!
1*
b11 6
19
1>
1C
b11 G
#659400000000
0!
0*
09
0>
0C
#659410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#659420000000
0!
0*
09
0>
0C
#659430000000
1!
1*
b101 6
19
1>
1C
b101 G
#659440000000
0!
0*
09
0>
0C
#659450000000
1!
1*
b110 6
19
1>
1C
b110 G
#659460000000
0!
0*
09
0>
0C
#659470000000
1!
1*
b111 6
19
1>
1C
b111 G
#659480000000
0!
0*
09
0>
0C
#659490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#659500000000
0!
0*
09
0>
0C
#659510000000
1!
1*
b1 6
19
1>
1C
b1 G
#659520000000
0!
0*
09
0>
0C
#659530000000
1!
1*
b10 6
19
1>
1C
b10 G
#659540000000
0!
0*
09
0>
0C
#659550000000
1!
1*
b11 6
19
1>
1C
b11 G
#659560000000
0!
0*
09
0>
0C
#659570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#659580000000
0!
0*
09
0>
0C
#659590000000
1!
1*
b101 6
19
1>
1C
b101 G
#659600000000
0!
0*
09
0>
0C
#659610000000
1!
1*
b110 6
19
1>
1C
b110 G
#659620000000
0!
0*
09
0>
0C
#659630000000
1!
1*
b111 6
19
1>
1C
b111 G
#659640000000
0!
1"
0*
1+
09
1:
0>
0C
#659650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#659660000000
0!
0*
09
0>
0C
#659670000000
1!
1*
b1 6
19
1>
1C
b1 G
#659680000000
0!
0*
09
0>
0C
#659690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#659700000000
0!
0*
09
0>
0C
#659710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#659720000000
0!
0*
09
0>
0C
#659730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#659740000000
0!
0*
09
0>
0C
#659750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#659760000000
0!
0#
0*
0,
09
0>
0?
0C
#659770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#659780000000
0!
0*
09
0>
0C
#659790000000
1!
1*
19
1>
1C
#659800000000
0!
0*
09
0>
0C
#659810000000
1!
1*
19
1>
1C
#659820000000
0!
0*
09
0>
0C
#659830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#659840000000
0!
0*
09
0>
0C
#659850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#659860000000
0!
0*
09
0>
0C
#659870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#659880000000
0!
0*
09
0>
0C
#659890000000
1!
1*
b10 6
19
1>
1C
b10 G
#659900000000
0!
0*
09
0>
0C
#659910000000
1!
1*
b11 6
19
1>
1C
b11 G
#659920000000
0!
0*
09
0>
0C
#659930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#659940000000
0!
0*
09
0>
0C
#659950000000
1!
1*
b101 6
19
1>
1C
b101 G
#659960000000
0!
0*
09
0>
0C
#659970000000
1!
1*
b110 6
19
1>
1C
b110 G
#659980000000
0!
0*
09
0>
0C
#659990000000
1!
1*
b111 6
19
1>
1C
b111 G
#660000000000
0!
0*
09
0>
0C
#660010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#660020000000
0!
0*
09
0>
0C
#660030000000
1!
1*
b1 6
19
1>
1C
b1 G
#660040000000
0!
0*
09
0>
0C
#660050000000
1!
1*
b10 6
19
1>
1C
b10 G
#660060000000
0!
0*
09
0>
0C
#660070000000
1!
1*
b11 6
19
1>
1C
b11 G
#660080000000
0!
0*
09
0>
0C
#660090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#660100000000
0!
0*
09
0>
0C
#660110000000
1!
1*
b101 6
19
1>
1C
b101 G
#660120000000
0!
0*
09
0>
0C
#660130000000
1!
1*
b110 6
19
1>
1C
b110 G
#660140000000
0!
0*
09
0>
0C
#660150000000
1!
1*
b111 6
19
1>
1C
b111 G
#660160000000
0!
0*
09
0>
0C
#660170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#660180000000
0!
0*
09
0>
0C
#660190000000
1!
1*
b1 6
19
1>
1C
b1 G
#660200000000
0!
0*
09
0>
0C
#660210000000
1!
1*
b10 6
19
1>
1C
b10 G
#660220000000
0!
0*
09
0>
0C
#660230000000
1!
1*
b11 6
19
1>
1C
b11 G
#660240000000
0!
0*
09
0>
0C
#660250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#660260000000
0!
0*
09
0>
0C
#660270000000
1!
1*
b101 6
19
1>
1C
b101 G
#660280000000
0!
0*
09
0>
0C
#660290000000
1!
1*
b110 6
19
1>
1C
b110 G
#660300000000
0!
0*
09
0>
0C
#660310000000
1!
1*
b111 6
19
1>
1C
b111 G
#660320000000
0!
1"
0*
1+
09
1:
0>
0C
#660330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#660340000000
0!
0*
09
0>
0C
#660350000000
1!
1*
b1 6
19
1>
1C
b1 G
#660360000000
0!
0*
09
0>
0C
#660370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#660380000000
0!
0*
09
0>
0C
#660390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#660400000000
0!
0*
09
0>
0C
#660410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#660420000000
0!
0*
09
0>
0C
#660430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#660440000000
0!
0#
0*
0,
09
0>
0?
0C
#660450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#660460000000
0!
0*
09
0>
0C
#660470000000
1!
1*
19
1>
1C
#660480000000
0!
0*
09
0>
0C
#660490000000
1!
1*
19
1>
1C
#660500000000
0!
0*
09
0>
0C
#660510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#660520000000
0!
0*
09
0>
0C
#660530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#660540000000
0!
0*
09
0>
0C
#660550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#660560000000
0!
0*
09
0>
0C
#660570000000
1!
1*
b10 6
19
1>
1C
b10 G
#660580000000
0!
0*
09
0>
0C
#660590000000
1!
1*
b11 6
19
1>
1C
b11 G
#660600000000
0!
0*
09
0>
0C
#660610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#660620000000
0!
0*
09
0>
0C
#660630000000
1!
1*
b101 6
19
1>
1C
b101 G
#660640000000
0!
0*
09
0>
0C
#660650000000
1!
1*
b110 6
19
1>
1C
b110 G
#660660000000
0!
0*
09
0>
0C
#660670000000
1!
1*
b111 6
19
1>
1C
b111 G
#660680000000
0!
0*
09
0>
0C
#660690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#660700000000
0!
0*
09
0>
0C
#660710000000
1!
1*
b1 6
19
1>
1C
b1 G
#660720000000
0!
0*
09
0>
0C
#660730000000
1!
1*
b10 6
19
1>
1C
b10 G
#660740000000
0!
0*
09
0>
0C
#660750000000
1!
1*
b11 6
19
1>
1C
b11 G
#660760000000
0!
0*
09
0>
0C
#660770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#660780000000
0!
0*
09
0>
0C
#660790000000
1!
1*
b101 6
19
1>
1C
b101 G
#660800000000
0!
0*
09
0>
0C
#660810000000
1!
1*
b110 6
19
1>
1C
b110 G
#660820000000
0!
0*
09
0>
0C
#660830000000
1!
1*
b111 6
19
1>
1C
b111 G
#660840000000
0!
0*
09
0>
0C
#660850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#660860000000
0!
0*
09
0>
0C
#660870000000
1!
1*
b1 6
19
1>
1C
b1 G
#660880000000
0!
0*
09
0>
0C
#660890000000
1!
1*
b10 6
19
1>
1C
b10 G
#660900000000
0!
0*
09
0>
0C
#660910000000
1!
1*
b11 6
19
1>
1C
b11 G
#660920000000
0!
0*
09
0>
0C
#660930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#660940000000
0!
0*
09
0>
0C
#660950000000
1!
1*
b101 6
19
1>
1C
b101 G
#660960000000
0!
0*
09
0>
0C
#660970000000
1!
1*
b110 6
19
1>
1C
b110 G
#660980000000
0!
0*
09
0>
0C
#660990000000
1!
1*
b111 6
19
1>
1C
b111 G
#661000000000
0!
1"
0*
1+
09
1:
0>
0C
#661010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#661020000000
0!
0*
09
0>
0C
#661030000000
1!
1*
b1 6
19
1>
1C
b1 G
#661040000000
0!
0*
09
0>
0C
#661050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#661060000000
0!
0*
09
0>
0C
#661070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#661080000000
0!
0*
09
0>
0C
#661090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#661100000000
0!
0*
09
0>
0C
#661110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#661120000000
0!
0#
0*
0,
09
0>
0?
0C
#661130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#661140000000
0!
0*
09
0>
0C
#661150000000
1!
1*
19
1>
1C
#661160000000
0!
0*
09
0>
0C
#661170000000
1!
1*
19
1>
1C
#661180000000
0!
0*
09
0>
0C
#661190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#661200000000
0!
0*
09
0>
0C
#661210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#661220000000
0!
0*
09
0>
0C
#661230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#661240000000
0!
0*
09
0>
0C
#661250000000
1!
1*
b10 6
19
1>
1C
b10 G
#661260000000
0!
0*
09
0>
0C
#661270000000
1!
1*
b11 6
19
1>
1C
b11 G
#661280000000
0!
0*
09
0>
0C
#661290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#661300000000
0!
0*
09
0>
0C
#661310000000
1!
1*
b101 6
19
1>
1C
b101 G
#661320000000
0!
0*
09
0>
0C
#661330000000
1!
1*
b110 6
19
1>
1C
b110 G
#661340000000
0!
0*
09
0>
0C
#661350000000
1!
1*
b111 6
19
1>
1C
b111 G
#661360000000
0!
0*
09
0>
0C
#661370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#661380000000
0!
0*
09
0>
0C
#661390000000
1!
1*
b1 6
19
1>
1C
b1 G
#661400000000
0!
0*
09
0>
0C
#661410000000
1!
1*
b10 6
19
1>
1C
b10 G
#661420000000
0!
0*
09
0>
0C
#661430000000
1!
1*
b11 6
19
1>
1C
b11 G
#661440000000
0!
0*
09
0>
0C
#661450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#661460000000
0!
0*
09
0>
0C
#661470000000
1!
1*
b101 6
19
1>
1C
b101 G
#661480000000
0!
0*
09
0>
0C
#661490000000
1!
1*
b110 6
19
1>
1C
b110 G
#661500000000
0!
0*
09
0>
0C
#661510000000
1!
1*
b111 6
19
1>
1C
b111 G
#661520000000
0!
0*
09
0>
0C
#661530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#661540000000
0!
0*
09
0>
0C
#661550000000
1!
1*
b1 6
19
1>
1C
b1 G
#661560000000
0!
0*
09
0>
0C
#661570000000
1!
1*
b10 6
19
1>
1C
b10 G
#661580000000
0!
0*
09
0>
0C
#661590000000
1!
1*
b11 6
19
1>
1C
b11 G
#661600000000
0!
0*
09
0>
0C
#661610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#661620000000
0!
0*
09
0>
0C
#661630000000
1!
1*
b101 6
19
1>
1C
b101 G
#661640000000
0!
0*
09
0>
0C
#661650000000
1!
1*
b110 6
19
1>
1C
b110 G
#661660000000
0!
0*
09
0>
0C
#661670000000
1!
1*
b111 6
19
1>
1C
b111 G
#661680000000
0!
1"
0*
1+
09
1:
0>
0C
#661690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#661700000000
0!
0*
09
0>
0C
#661710000000
1!
1*
b1 6
19
1>
1C
b1 G
#661720000000
0!
0*
09
0>
0C
#661730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#661740000000
0!
0*
09
0>
0C
#661750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#661760000000
0!
0*
09
0>
0C
#661770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#661780000000
0!
0*
09
0>
0C
#661790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#661800000000
0!
0#
0*
0,
09
0>
0?
0C
#661810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#661820000000
0!
0*
09
0>
0C
#661830000000
1!
1*
19
1>
1C
#661840000000
0!
0*
09
0>
0C
#661850000000
1!
1*
19
1>
1C
#661860000000
0!
0*
09
0>
0C
#661870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#661880000000
0!
0*
09
0>
0C
#661890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#661900000000
0!
0*
09
0>
0C
#661910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#661920000000
0!
0*
09
0>
0C
#661930000000
1!
1*
b10 6
19
1>
1C
b10 G
#661940000000
0!
0*
09
0>
0C
#661950000000
1!
1*
b11 6
19
1>
1C
b11 G
#661960000000
0!
0*
09
0>
0C
#661970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#661980000000
0!
0*
09
0>
0C
#661990000000
1!
1*
b101 6
19
1>
1C
b101 G
#662000000000
0!
0*
09
0>
0C
#662010000000
1!
1*
b110 6
19
1>
1C
b110 G
#662020000000
0!
0*
09
0>
0C
#662030000000
1!
1*
b111 6
19
1>
1C
b111 G
#662040000000
0!
0*
09
0>
0C
#662050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#662060000000
0!
0*
09
0>
0C
#662070000000
1!
1*
b1 6
19
1>
1C
b1 G
#662080000000
0!
0*
09
0>
0C
#662090000000
1!
1*
b10 6
19
1>
1C
b10 G
#662100000000
0!
0*
09
0>
0C
#662110000000
1!
1*
b11 6
19
1>
1C
b11 G
#662120000000
0!
0*
09
0>
0C
#662130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#662140000000
0!
0*
09
0>
0C
#662150000000
1!
1*
b101 6
19
1>
1C
b101 G
#662160000000
0!
0*
09
0>
0C
#662170000000
1!
1*
b110 6
19
1>
1C
b110 G
#662180000000
0!
0*
09
0>
0C
#662190000000
1!
1*
b111 6
19
1>
1C
b111 G
#662200000000
0!
0*
09
0>
0C
#662210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#662220000000
0!
0*
09
0>
0C
#662230000000
1!
1*
b1 6
19
1>
1C
b1 G
#662240000000
0!
0*
09
0>
0C
#662250000000
1!
1*
b10 6
19
1>
1C
b10 G
#662260000000
0!
0*
09
0>
0C
#662270000000
1!
1*
b11 6
19
1>
1C
b11 G
#662280000000
0!
0*
09
0>
0C
#662290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#662300000000
0!
0*
09
0>
0C
#662310000000
1!
1*
b101 6
19
1>
1C
b101 G
#662320000000
0!
0*
09
0>
0C
#662330000000
1!
1*
b110 6
19
1>
1C
b110 G
#662340000000
0!
0*
09
0>
0C
#662350000000
1!
1*
b111 6
19
1>
1C
b111 G
#662360000000
0!
1"
0*
1+
09
1:
0>
0C
#662370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#662380000000
0!
0*
09
0>
0C
#662390000000
1!
1*
b1 6
19
1>
1C
b1 G
#662400000000
0!
0*
09
0>
0C
#662410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#662420000000
0!
0*
09
0>
0C
#662430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#662440000000
0!
0*
09
0>
0C
#662450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#662460000000
0!
0*
09
0>
0C
#662470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#662480000000
0!
0#
0*
0,
09
0>
0?
0C
#662490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#662500000000
0!
0*
09
0>
0C
#662510000000
1!
1*
19
1>
1C
#662520000000
0!
0*
09
0>
0C
#662530000000
1!
1*
19
1>
1C
#662540000000
0!
0*
09
0>
0C
#662550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#662560000000
0!
0*
09
0>
0C
#662570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#662580000000
0!
0*
09
0>
0C
#662590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#662600000000
0!
0*
09
0>
0C
#662610000000
1!
1*
b10 6
19
1>
1C
b10 G
#662620000000
0!
0*
09
0>
0C
#662630000000
1!
1*
b11 6
19
1>
1C
b11 G
#662640000000
0!
0*
09
0>
0C
#662650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#662660000000
0!
0*
09
0>
0C
#662670000000
1!
1*
b101 6
19
1>
1C
b101 G
#662680000000
0!
0*
09
0>
0C
#662690000000
1!
1*
b110 6
19
1>
1C
b110 G
#662700000000
0!
0*
09
0>
0C
#662710000000
1!
1*
b111 6
19
1>
1C
b111 G
#662720000000
0!
0*
09
0>
0C
#662730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#662740000000
0!
0*
09
0>
0C
#662750000000
1!
1*
b1 6
19
1>
1C
b1 G
#662760000000
0!
0*
09
0>
0C
#662770000000
1!
1*
b10 6
19
1>
1C
b10 G
#662780000000
0!
0*
09
0>
0C
#662790000000
1!
1*
b11 6
19
1>
1C
b11 G
#662800000000
0!
0*
09
0>
0C
#662810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#662820000000
0!
0*
09
0>
0C
#662830000000
1!
1*
b101 6
19
1>
1C
b101 G
#662840000000
0!
0*
09
0>
0C
#662850000000
1!
1*
b110 6
19
1>
1C
b110 G
#662860000000
0!
0*
09
0>
0C
#662870000000
1!
1*
b111 6
19
1>
1C
b111 G
#662880000000
0!
0*
09
0>
0C
#662890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#662900000000
0!
0*
09
0>
0C
#662910000000
1!
1*
b1 6
19
1>
1C
b1 G
#662920000000
0!
0*
09
0>
0C
#662930000000
1!
1*
b10 6
19
1>
1C
b10 G
#662940000000
0!
0*
09
0>
0C
#662950000000
1!
1*
b11 6
19
1>
1C
b11 G
#662960000000
0!
0*
09
0>
0C
#662970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#662980000000
0!
0*
09
0>
0C
#662990000000
1!
1*
b101 6
19
1>
1C
b101 G
#663000000000
0!
0*
09
0>
0C
#663010000000
1!
1*
b110 6
19
1>
1C
b110 G
#663020000000
0!
0*
09
0>
0C
#663030000000
1!
1*
b111 6
19
1>
1C
b111 G
#663040000000
0!
1"
0*
1+
09
1:
0>
0C
#663050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#663060000000
0!
0*
09
0>
0C
#663070000000
1!
1*
b1 6
19
1>
1C
b1 G
#663080000000
0!
0*
09
0>
0C
#663090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#663100000000
0!
0*
09
0>
0C
#663110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#663120000000
0!
0*
09
0>
0C
#663130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#663140000000
0!
0*
09
0>
0C
#663150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#663160000000
0!
0#
0*
0,
09
0>
0?
0C
#663170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#663180000000
0!
0*
09
0>
0C
#663190000000
1!
1*
19
1>
1C
#663200000000
0!
0*
09
0>
0C
#663210000000
1!
1*
19
1>
1C
#663220000000
0!
0*
09
0>
0C
#663230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#663240000000
0!
0*
09
0>
0C
#663250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#663260000000
0!
0*
09
0>
0C
#663270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#663280000000
0!
0*
09
0>
0C
#663290000000
1!
1*
b10 6
19
1>
1C
b10 G
#663300000000
0!
0*
09
0>
0C
#663310000000
1!
1*
b11 6
19
1>
1C
b11 G
#663320000000
0!
0*
09
0>
0C
#663330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#663340000000
0!
0*
09
0>
0C
#663350000000
1!
1*
b101 6
19
1>
1C
b101 G
#663360000000
0!
0*
09
0>
0C
#663370000000
1!
1*
b110 6
19
1>
1C
b110 G
#663380000000
0!
0*
09
0>
0C
#663390000000
1!
1*
b111 6
19
1>
1C
b111 G
#663400000000
0!
0*
09
0>
0C
#663410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#663420000000
0!
0*
09
0>
0C
#663430000000
1!
1*
b1 6
19
1>
1C
b1 G
#663440000000
0!
0*
09
0>
0C
#663450000000
1!
1*
b10 6
19
1>
1C
b10 G
#663460000000
0!
0*
09
0>
0C
#663470000000
1!
1*
b11 6
19
1>
1C
b11 G
#663480000000
0!
0*
09
0>
0C
#663490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#663500000000
0!
0*
09
0>
0C
#663510000000
1!
1*
b101 6
19
1>
1C
b101 G
#663520000000
0!
0*
09
0>
0C
#663530000000
1!
1*
b110 6
19
1>
1C
b110 G
#663540000000
0!
0*
09
0>
0C
#663550000000
1!
1*
b111 6
19
1>
1C
b111 G
#663560000000
0!
0*
09
0>
0C
#663570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#663580000000
0!
0*
09
0>
0C
#663590000000
1!
1*
b1 6
19
1>
1C
b1 G
#663600000000
0!
0*
09
0>
0C
#663610000000
1!
1*
b10 6
19
1>
1C
b10 G
#663620000000
0!
0*
09
0>
0C
#663630000000
1!
1*
b11 6
19
1>
1C
b11 G
#663640000000
0!
0*
09
0>
0C
#663650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#663660000000
0!
0*
09
0>
0C
#663670000000
1!
1*
b101 6
19
1>
1C
b101 G
#663680000000
0!
0*
09
0>
0C
#663690000000
1!
1*
b110 6
19
1>
1C
b110 G
#663700000000
0!
0*
09
0>
0C
#663710000000
1!
1*
b111 6
19
1>
1C
b111 G
#663720000000
0!
1"
0*
1+
09
1:
0>
0C
#663730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#663740000000
0!
0*
09
0>
0C
#663750000000
1!
1*
b1 6
19
1>
1C
b1 G
#663760000000
0!
0*
09
0>
0C
#663770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#663780000000
0!
0*
09
0>
0C
#663790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#663800000000
0!
0*
09
0>
0C
#663810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#663820000000
0!
0*
09
0>
0C
#663830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#663840000000
0!
0#
0*
0,
09
0>
0?
0C
#663850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#663860000000
0!
0*
09
0>
0C
#663870000000
1!
1*
19
1>
1C
#663880000000
0!
0*
09
0>
0C
#663890000000
1!
1*
19
1>
1C
#663900000000
0!
0*
09
0>
0C
#663910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#663920000000
0!
0*
09
0>
0C
#663930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#663940000000
0!
0*
09
0>
0C
#663950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#663960000000
0!
0*
09
0>
0C
#663970000000
1!
1*
b10 6
19
1>
1C
b10 G
#663980000000
0!
0*
09
0>
0C
#663990000000
1!
1*
b11 6
19
1>
1C
b11 G
#664000000000
0!
0*
09
0>
0C
#664010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#664020000000
0!
0*
09
0>
0C
#664030000000
1!
1*
b101 6
19
1>
1C
b101 G
#664040000000
0!
0*
09
0>
0C
#664050000000
1!
1*
b110 6
19
1>
1C
b110 G
#664060000000
0!
0*
09
0>
0C
#664070000000
1!
1*
b111 6
19
1>
1C
b111 G
#664080000000
0!
0*
09
0>
0C
#664090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#664100000000
0!
0*
09
0>
0C
#664110000000
1!
1*
b1 6
19
1>
1C
b1 G
#664120000000
0!
0*
09
0>
0C
#664130000000
1!
1*
b10 6
19
1>
1C
b10 G
#664140000000
0!
0*
09
0>
0C
#664150000000
1!
1*
b11 6
19
1>
1C
b11 G
#664160000000
0!
0*
09
0>
0C
#664170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#664180000000
0!
0*
09
0>
0C
#664190000000
1!
1*
b101 6
19
1>
1C
b101 G
#664200000000
0!
0*
09
0>
0C
#664210000000
1!
1*
b110 6
19
1>
1C
b110 G
#664220000000
0!
0*
09
0>
0C
#664230000000
1!
1*
b111 6
19
1>
1C
b111 G
#664240000000
0!
0*
09
0>
0C
#664250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#664260000000
0!
0*
09
0>
0C
#664270000000
1!
1*
b1 6
19
1>
1C
b1 G
#664280000000
0!
0*
09
0>
0C
#664290000000
1!
1*
b10 6
19
1>
1C
b10 G
#664300000000
0!
0*
09
0>
0C
#664310000000
1!
1*
b11 6
19
1>
1C
b11 G
#664320000000
0!
0*
09
0>
0C
#664330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#664340000000
0!
0*
09
0>
0C
#664350000000
1!
1*
b101 6
19
1>
1C
b101 G
#664360000000
0!
0*
09
0>
0C
#664370000000
1!
1*
b110 6
19
1>
1C
b110 G
#664380000000
0!
0*
09
0>
0C
#664390000000
1!
1*
b111 6
19
1>
1C
b111 G
#664400000000
0!
1"
0*
1+
09
1:
0>
0C
#664410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#664420000000
0!
0*
09
0>
0C
#664430000000
1!
1*
b1 6
19
1>
1C
b1 G
#664440000000
0!
0*
09
0>
0C
#664450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#664460000000
0!
0*
09
0>
0C
#664470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#664480000000
0!
0*
09
0>
0C
#664490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#664500000000
0!
0*
09
0>
0C
#664510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#664520000000
0!
0#
0*
0,
09
0>
0?
0C
#664530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#664540000000
0!
0*
09
0>
0C
#664550000000
1!
1*
19
1>
1C
#664560000000
0!
0*
09
0>
0C
#664570000000
1!
1*
19
1>
1C
#664580000000
0!
0*
09
0>
0C
#664590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#664600000000
0!
0*
09
0>
0C
#664610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#664620000000
0!
0*
09
0>
0C
#664630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#664640000000
0!
0*
09
0>
0C
#664650000000
1!
1*
b10 6
19
1>
1C
b10 G
#664660000000
0!
0*
09
0>
0C
#664670000000
1!
1*
b11 6
19
1>
1C
b11 G
#664680000000
0!
0*
09
0>
0C
#664690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#664700000000
0!
0*
09
0>
0C
#664710000000
1!
1*
b101 6
19
1>
1C
b101 G
#664720000000
0!
0*
09
0>
0C
#664730000000
1!
1*
b110 6
19
1>
1C
b110 G
#664740000000
0!
0*
09
0>
0C
#664750000000
1!
1*
b111 6
19
1>
1C
b111 G
#664760000000
0!
0*
09
0>
0C
#664770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#664780000000
0!
0*
09
0>
0C
#664790000000
1!
1*
b1 6
19
1>
1C
b1 G
#664800000000
0!
0*
09
0>
0C
#664810000000
1!
1*
b10 6
19
1>
1C
b10 G
#664820000000
0!
0*
09
0>
0C
#664830000000
1!
1*
b11 6
19
1>
1C
b11 G
#664840000000
0!
0*
09
0>
0C
#664850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#664860000000
0!
0*
09
0>
0C
#664870000000
1!
1*
b101 6
19
1>
1C
b101 G
#664880000000
0!
0*
09
0>
0C
#664890000000
1!
1*
b110 6
19
1>
1C
b110 G
#664900000000
0!
0*
09
0>
0C
#664910000000
1!
1*
b111 6
19
1>
1C
b111 G
#664920000000
0!
0*
09
0>
0C
#664930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#664940000000
0!
0*
09
0>
0C
#664950000000
1!
1*
b1 6
19
1>
1C
b1 G
#664960000000
0!
0*
09
0>
0C
#664970000000
1!
1*
b10 6
19
1>
1C
b10 G
#664980000000
0!
0*
09
0>
0C
#664990000000
1!
1*
b11 6
19
1>
1C
b11 G
#665000000000
0!
0*
09
0>
0C
#665010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#665020000000
0!
0*
09
0>
0C
#665030000000
1!
1*
b101 6
19
1>
1C
b101 G
#665040000000
0!
0*
09
0>
0C
#665050000000
1!
1*
b110 6
19
1>
1C
b110 G
#665060000000
0!
0*
09
0>
0C
#665070000000
1!
1*
b111 6
19
1>
1C
b111 G
#665080000000
0!
1"
0*
1+
09
1:
0>
0C
#665090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#665100000000
0!
0*
09
0>
0C
#665110000000
1!
1*
b1 6
19
1>
1C
b1 G
#665120000000
0!
0*
09
0>
0C
#665130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#665140000000
0!
0*
09
0>
0C
#665150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#665160000000
0!
0*
09
0>
0C
#665170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#665180000000
0!
0*
09
0>
0C
#665190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#665200000000
0!
0#
0*
0,
09
0>
0?
0C
#665210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#665220000000
0!
0*
09
0>
0C
#665230000000
1!
1*
19
1>
1C
#665240000000
0!
0*
09
0>
0C
#665250000000
1!
1*
19
1>
1C
#665260000000
0!
0*
09
0>
0C
#665270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#665280000000
0!
0*
09
0>
0C
#665290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#665300000000
0!
0*
09
0>
0C
#665310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#665320000000
0!
0*
09
0>
0C
#665330000000
1!
1*
b10 6
19
1>
1C
b10 G
#665340000000
0!
0*
09
0>
0C
#665350000000
1!
1*
b11 6
19
1>
1C
b11 G
#665360000000
0!
0*
09
0>
0C
#665370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#665380000000
0!
0*
09
0>
0C
#665390000000
1!
1*
b101 6
19
1>
1C
b101 G
#665400000000
0!
0*
09
0>
0C
#665410000000
1!
1*
b110 6
19
1>
1C
b110 G
#665420000000
0!
0*
09
0>
0C
#665430000000
1!
1*
b111 6
19
1>
1C
b111 G
#665440000000
0!
0*
09
0>
0C
#665450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#665460000000
0!
0*
09
0>
0C
#665470000000
1!
1*
b1 6
19
1>
1C
b1 G
#665480000000
0!
0*
09
0>
0C
#665490000000
1!
1*
b10 6
19
1>
1C
b10 G
#665500000000
0!
0*
09
0>
0C
#665510000000
1!
1*
b11 6
19
1>
1C
b11 G
#665520000000
0!
0*
09
0>
0C
#665530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#665540000000
0!
0*
09
0>
0C
#665550000000
1!
1*
b101 6
19
1>
1C
b101 G
#665560000000
0!
0*
09
0>
0C
#665570000000
1!
1*
b110 6
19
1>
1C
b110 G
#665580000000
0!
0*
09
0>
0C
#665590000000
1!
1*
b111 6
19
1>
1C
b111 G
#665600000000
0!
0*
09
0>
0C
#665610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#665620000000
0!
0*
09
0>
0C
#665630000000
1!
1*
b1 6
19
1>
1C
b1 G
#665640000000
0!
0*
09
0>
0C
#665650000000
1!
1*
b10 6
19
1>
1C
b10 G
#665660000000
0!
0*
09
0>
0C
#665670000000
1!
1*
b11 6
19
1>
1C
b11 G
#665680000000
0!
0*
09
0>
0C
#665690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#665700000000
0!
0*
09
0>
0C
#665710000000
1!
1*
b101 6
19
1>
1C
b101 G
#665720000000
0!
0*
09
0>
0C
#665730000000
1!
1*
b110 6
19
1>
1C
b110 G
#665740000000
0!
0*
09
0>
0C
#665750000000
1!
1*
b111 6
19
1>
1C
b111 G
#665760000000
0!
1"
0*
1+
09
1:
0>
0C
#665770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#665780000000
0!
0*
09
0>
0C
#665790000000
1!
1*
b1 6
19
1>
1C
b1 G
#665800000000
0!
0*
09
0>
0C
#665810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#665820000000
0!
0*
09
0>
0C
#665830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#665840000000
0!
0*
09
0>
0C
#665850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#665860000000
0!
0*
09
0>
0C
#665870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#665880000000
0!
0#
0*
0,
09
0>
0?
0C
#665890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#665900000000
0!
0*
09
0>
0C
#665910000000
1!
1*
19
1>
1C
#665920000000
0!
0*
09
0>
0C
#665930000000
1!
1*
19
1>
1C
#665940000000
0!
0*
09
0>
0C
#665950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#665960000000
0!
0*
09
0>
0C
#665970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#665980000000
0!
0*
09
0>
0C
#665990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#666000000000
0!
0*
09
0>
0C
#666010000000
1!
1*
b10 6
19
1>
1C
b10 G
#666020000000
0!
0*
09
0>
0C
#666030000000
1!
1*
b11 6
19
1>
1C
b11 G
#666040000000
0!
0*
09
0>
0C
#666050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#666060000000
0!
0*
09
0>
0C
#666070000000
1!
1*
b101 6
19
1>
1C
b101 G
#666080000000
0!
0*
09
0>
0C
#666090000000
1!
1*
b110 6
19
1>
1C
b110 G
#666100000000
0!
0*
09
0>
0C
#666110000000
1!
1*
b111 6
19
1>
1C
b111 G
#666120000000
0!
0*
09
0>
0C
#666130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#666140000000
0!
0*
09
0>
0C
#666150000000
1!
1*
b1 6
19
1>
1C
b1 G
#666160000000
0!
0*
09
0>
0C
#666170000000
1!
1*
b10 6
19
1>
1C
b10 G
#666180000000
0!
0*
09
0>
0C
#666190000000
1!
1*
b11 6
19
1>
1C
b11 G
#666200000000
0!
0*
09
0>
0C
#666210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#666220000000
0!
0*
09
0>
0C
#666230000000
1!
1*
b101 6
19
1>
1C
b101 G
#666240000000
0!
0*
09
0>
0C
#666250000000
1!
1*
b110 6
19
1>
1C
b110 G
#666260000000
0!
0*
09
0>
0C
#666270000000
1!
1*
b111 6
19
1>
1C
b111 G
#666280000000
0!
0*
09
0>
0C
#666290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#666300000000
0!
0*
09
0>
0C
#666310000000
1!
1*
b1 6
19
1>
1C
b1 G
#666320000000
0!
0*
09
0>
0C
#666330000000
1!
1*
b10 6
19
1>
1C
b10 G
#666340000000
0!
0*
09
0>
0C
#666350000000
1!
1*
b11 6
19
1>
1C
b11 G
#666360000000
0!
0*
09
0>
0C
#666370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#666380000000
0!
0*
09
0>
0C
#666390000000
1!
1*
b101 6
19
1>
1C
b101 G
#666400000000
0!
0*
09
0>
0C
#666410000000
1!
1*
b110 6
19
1>
1C
b110 G
#666420000000
0!
0*
09
0>
0C
#666430000000
1!
1*
b111 6
19
1>
1C
b111 G
#666440000000
0!
1"
0*
1+
09
1:
0>
0C
#666450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#666460000000
0!
0*
09
0>
0C
#666470000000
1!
1*
b1 6
19
1>
1C
b1 G
#666480000000
0!
0*
09
0>
0C
#666490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#666500000000
0!
0*
09
0>
0C
#666510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#666520000000
0!
0*
09
0>
0C
#666530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#666540000000
0!
0*
09
0>
0C
#666550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#666560000000
0!
0#
0*
0,
09
0>
0?
0C
#666570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#666580000000
0!
0*
09
0>
0C
#666590000000
1!
1*
19
1>
1C
#666600000000
0!
0*
09
0>
0C
#666610000000
1!
1*
19
1>
1C
#666620000000
0!
0*
09
0>
0C
#666630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#666640000000
0!
0*
09
0>
0C
#666650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#666660000000
0!
0*
09
0>
0C
#666670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#666680000000
0!
0*
09
0>
0C
#666690000000
1!
1*
b10 6
19
1>
1C
b10 G
#666700000000
0!
0*
09
0>
0C
#666710000000
1!
1*
b11 6
19
1>
1C
b11 G
#666720000000
0!
0*
09
0>
0C
#666730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#666740000000
0!
0*
09
0>
0C
#666750000000
1!
1*
b101 6
19
1>
1C
b101 G
#666760000000
0!
0*
09
0>
0C
#666770000000
1!
1*
b110 6
19
1>
1C
b110 G
#666780000000
0!
0*
09
0>
0C
#666790000000
1!
1*
b111 6
19
1>
1C
b111 G
#666800000000
0!
0*
09
0>
0C
#666810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#666820000000
0!
0*
09
0>
0C
#666830000000
1!
1*
b1 6
19
1>
1C
b1 G
#666840000000
0!
0*
09
0>
0C
#666850000000
1!
1*
b10 6
19
1>
1C
b10 G
#666860000000
0!
0*
09
0>
0C
#666870000000
1!
1*
b11 6
19
1>
1C
b11 G
#666880000000
0!
0*
09
0>
0C
#666890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#666900000000
0!
0*
09
0>
0C
#666910000000
1!
1*
b101 6
19
1>
1C
b101 G
#666920000000
0!
0*
09
0>
0C
#666930000000
1!
1*
b110 6
19
1>
1C
b110 G
#666940000000
0!
0*
09
0>
0C
#666950000000
1!
1*
b111 6
19
1>
1C
b111 G
#666960000000
0!
0*
09
0>
0C
#666970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#666980000000
0!
0*
09
0>
0C
#666990000000
1!
1*
b1 6
19
1>
1C
b1 G
#667000000000
0!
0*
09
0>
0C
#667010000000
1!
1*
b10 6
19
1>
1C
b10 G
#667020000000
0!
0*
09
0>
0C
#667030000000
1!
1*
b11 6
19
1>
1C
b11 G
#667040000000
0!
0*
09
0>
0C
#667050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#667060000000
0!
0*
09
0>
0C
#667070000000
1!
1*
b101 6
19
1>
1C
b101 G
#667080000000
0!
0*
09
0>
0C
#667090000000
1!
1*
b110 6
19
1>
1C
b110 G
#667100000000
0!
0*
09
0>
0C
#667110000000
1!
1*
b111 6
19
1>
1C
b111 G
#667120000000
0!
1"
0*
1+
09
1:
0>
0C
#667130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#667140000000
0!
0*
09
0>
0C
#667150000000
1!
1*
b1 6
19
1>
1C
b1 G
#667160000000
0!
0*
09
0>
0C
#667170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#667180000000
0!
0*
09
0>
0C
#667190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#667200000000
0!
0*
09
0>
0C
#667210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#667220000000
0!
0*
09
0>
0C
#667230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#667240000000
0!
0#
0*
0,
09
0>
0?
0C
#667250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#667260000000
0!
0*
09
0>
0C
#667270000000
1!
1*
19
1>
1C
#667280000000
0!
0*
09
0>
0C
#667290000000
1!
1*
19
1>
1C
#667300000000
0!
0*
09
0>
0C
#667310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#667320000000
0!
0*
09
0>
0C
#667330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#667340000000
0!
0*
09
0>
0C
#667350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#667360000000
0!
0*
09
0>
0C
#667370000000
1!
1*
b10 6
19
1>
1C
b10 G
#667380000000
0!
0*
09
0>
0C
#667390000000
1!
1*
b11 6
19
1>
1C
b11 G
#667400000000
0!
0*
09
0>
0C
#667410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#667420000000
0!
0*
09
0>
0C
#667430000000
1!
1*
b101 6
19
1>
1C
b101 G
#667440000000
0!
0*
09
0>
0C
#667450000000
1!
1*
b110 6
19
1>
1C
b110 G
#667460000000
0!
0*
09
0>
0C
#667470000000
1!
1*
b111 6
19
1>
1C
b111 G
#667480000000
0!
0*
09
0>
0C
#667490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#667500000000
0!
0*
09
0>
0C
#667510000000
1!
1*
b1 6
19
1>
1C
b1 G
#667520000000
0!
0*
09
0>
0C
#667530000000
1!
1*
b10 6
19
1>
1C
b10 G
#667540000000
0!
0*
09
0>
0C
#667550000000
1!
1*
b11 6
19
1>
1C
b11 G
#667560000000
0!
0*
09
0>
0C
#667570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#667580000000
0!
0*
09
0>
0C
#667590000000
1!
1*
b101 6
19
1>
1C
b101 G
#667600000000
0!
0*
09
0>
0C
#667610000000
1!
1*
b110 6
19
1>
1C
b110 G
#667620000000
0!
0*
09
0>
0C
#667630000000
1!
1*
b111 6
19
1>
1C
b111 G
#667640000000
0!
0*
09
0>
0C
#667650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#667660000000
0!
0*
09
0>
0C
#667670000000
1!
1*
b1 6
19
1>
1C
b1 G
#667680000000
0!
0*
09
0>
0C
#667690000000
1!
1*
b10 6
19
1>
1C
b10 G
#667700000000
0!
0*
09
0>
0C
#667710000000
1!
1*
b11 6
19
1>
1C
b11 G
#667720000000
0!
0*
09
0>
0C
#667730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#667740000000
0!
0*
09
0>
0C
#667750000000
1!
1*
b101 6
19
1>
1C
b101 G
#667760000000
0!
0*
09
0>
0C
#667770000000
1!
1*
b110 6
19
1>
1C
b110 G
#667780000000
0!
0*
09
0>
0C
#667790000000
1!
1*
b111 6
19
1>
1C
b111 G
#667800000000
0!
1"
0*
1+
09
1:
0>
0C
#667810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#667820000000
0!
0*
09
0>
0C
#667830000000
1!
1*
b1 6
19
1>
1C
b1 G
#667840000000
0!
0*
09
0>
0C
#667850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#667860000000
0!
0*
09
0>
0C
#667870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#667880000000
0!
0*
09
0>
0C
#667890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#667900000000
0!
0*
09
0>
0C
#667910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#667920000000
0!
0#
0*
0,
09
0>
0?
0C
#667930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#667940000000
0!
0*
09
0>
0C
#667950000000
1!
1*
19
1>
1C
#667960000000
0!
0*
09
0>
0C
#667970000000
1!
1*
19
1>
1C
#667980000000
0!
0*
09
0>
0C
#667990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#668000000000
0!
0*
09
0>
0C
#668010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#668020000000
0!
0*
09
0>
0C
#668030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#668040000000
0!
0*
09
0>
0C
#668050000000
1!
1*
b10 6
19
1>
1C
b10 G
#668060000000
0!
0*
09
0>
0C
#668070000000
1!
1*
b11 6
19
1>
1C
b11 G
#668080000000
0!
0*
09
0>
0C
#668090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#668100000000
0!
0*
09
0>
0C
#668110000000
1!
1*
b101 6
19
1>
1C
b101 G
#668120000000
0!
0*
09
0>
0C
#668130000000
1!
1*
b110 6
19
1>
1C
b110 G
#668140000000
0!
0*
09
0>
0C
#668150000000
1!
1*
b111 6
19
1>
1C
b111 G
#668160000000
0!
0*
09
0>
0C
#668170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#668180000000
0!
0*
09
0>
0C
#668190000000
1!
1*
b1 6
19
1>
1C
b1 G
#668200000000
0!
0*
09
0>
0C
#668210000000
1!
1*
b10 6
19
1>
1C
b10 G
#668220000000
0!
0*
09
0>
0C
#668230000000
1!
1*
b11 6
19
1>
1C
b11 G
#668240000000
0!
0*
09
0>
0C
#668250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#668260000000
0!
0*
09
0>
0C
#668270000000
1!
1*
b101 6
19
1>
1C
b101 G
#668280000000
0!
0*
09
0>
0C
#668290000000
1!
1*
b110 6
19
1>
1C
b110 G
#668300000000
0!
0*
09
0>
0C
#668310000000
1!
1*
b111 6
19
1>
1C
b111 G
#668320000000
0!
0*
09
0>
0C
#668330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#668340000000
0!
0*
09
0>
0C
#668350000000
1!
1*
b1 6
19
1>
1C
b1 G
#668360000000
0!
0*
09
0>
0C
#668370000000
1!
1*
b10 6
19
1>
1C
b10 G
#668380000000
0!
0*
09
0>
0C
#668390000000
1!
1*
b11 6
19
1>
1C
b11 G
#668400000000
0!
0*
09
0>
0C
#668410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#668420000000
0!
0*
09
0>
0C
#668430000000
1!
1*
b101 6
19
1>
1C
b101 G
#668440000000
0!
0*
09
0>
0C
#668450000000
1!
1*
b110 6
19
1>
1C
b110 G
#668460000000
0!
0*
09
0>
0C
#668470000000
1!
1*
b111 6
19
1>
1C
b111 G
#668480000000
0!
1"
0*
1+
09
1:
0>
0C
#668490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#668500000000
0!
0*
09
0>
0C
#668510000000
1!
1*
b1 6
19
1>
1C
b1 G
#668520000000
0!
0*
09
0>
0C
#668530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#668540000000
0!
0*
09
0>
0C
#668550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#668560000000
0!
0*
09
0>
0C
#668570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#668580000000
0!
0*
09
0>
0C
#668590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#668600000000
0!
0#
0*
0,
09
0>
0?
0C
#668610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#668620000000
0!
0*
09
0>
0C
#668630000000
1!
1*
19
1>
1C
#668640000000
0!
0*
09
0>
0C
#668650000000
1!
1*
19
1>
1C
#668660000000
0!
0*
09
0>
0C
#668670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#668680000000
0!
0*
09
0>
0C
#668690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#668700000000
0!
0*
09
0>
0C
#668710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#668720000000
0!
0*
09
0>
0C
#668730000000
1!
1*
b10 6
19
1>
1C
b10 G
#668740000000
0!
0*
09
0>
0C
#668750000000
1!
1*
b11 6
19
1>
1C
b11 G
#668760000000
0!
0*
09
0>
0C
#668770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#668780000000
0!
0*
09
0>
0C
#668790000000
1!
1*
b101 6
19
1>
1C
b101 G
#668800000000
0!
0*
09
0>
0C
#668810000000
1!
1*
b110 6
19
1>
1C
b110 G
#668820000000
0!
0*
09
0>
0C
#668830000000
1!
1*
b111 6
19
1>
1C
b111 G
#668840000000
0!
0*
09
0>
0C
#668850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#668860000000
0!
0*
09
0>
0C
#668870000000
1!
1*
b1 6
19
1>
1C
b1 G
#668880000000
0!
0*
09
0>
0C
#668890000000
1!
1*
b10 6
19
1>
1C
b10 G
#668900000000
0!
0*
09
0>
0C
#668910000000
1!
1*
b11 6
19
1>
1C
b11 G
#668920000000
0!
0*
09
0>
0C
#668930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#668940000000
0!
0*
09
0>
0C
#668950000000
1!
1*
b101 6
19
1>
1C
b101 G
#668960000000
0!
0*
09
0>
0C
#668970000000
1!
1*
b110 6
19
1>
1C
b110 G
#668980000000
0!
0*
09
0>
0C
#668990000000
1!
1*
b111 6
19
1>
1C
b111 G
#669000000000
0!
0*
09
0>
0C
#669010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#669020000000
0!
0*
09
0>
0C
#669030000000
1!
1*
b1 6
19
1>
1C
b1 G
#669040000000
0!
0*
09
0>
0C
#669050000000
1!
1*
b10 6
19
1>
1C
b10 G
#669060000000
0!
0*
09
0>
0C
#669070000000
1!
1*
b11 6
19
1>
1C
b11 G
#669080000000
0!
0*
09
0>
0C
#669090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#669100000000
0!
0*
09
0>
0C
#669110000000
1!
1*
b101 6
19
1>
1C
b101 G
#669120000000
0!
0*
09
0>
0C
#669130000000
1!
1*
b110 6
19
1>
1C
b110 G
#669140000000
0!
0*
09
0>
0C
#669150000000
1!
1*
b111 6
19
1>
1C
b111 G
#669160000000
0!
1"
0*
1+
09
1:
0>
0C
#669170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#669180000000
0!
0*
09
0>
0C
#669190000000
1!
1*
b1 6
19
1>
1C
b1 G
#669200000000
0!
0*
09
0>
0C
#669210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#669220000000
0!
0*
09
0>
0C
#669230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#669240000000
0!
0*
09
0>
0C
#669250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#669260000000
0!
0*
09
0>
0C
#669270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#669280000000
0!
0#
0*
0,
09
0>
0?
0C
#669290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#669300000000
0!
0*
09
0>
0C
#669310000000
1!
1*
19
1>
1C
#669320000000
0!
0*
09
0>
0C
#669330000000
1!
1*
19
1>
1C
#669340000000
0!
0*
09
0>
0C
#669350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#669360000000
0!
0*
09
0>
0C
#669370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#669380000000
0!
0*
09
0>
0C
#669390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#669400000000
0!
0*
09
0>
0C
#669410000000
1!
1*
b10 6
19
1>
1C
b10 G
#669420000000
0!
0*
09
0>
0C
#669430000000
1!
1*
b11 6
19
1>
1C
b11 G
#669440000000
0!
0*
09
0>
0C
#669450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#669460000000
0!
0*
09
0>
0C
#669470000000
1!
1*
b101 6
19
1>
1C
b101 G
#669480000000
0!
0*
09
0>
0C
#669490000000
1!
1*
b110 6
19
1>
1C
b110 G
#669500000000
0!
0*
09
0>
0C
#669510000000
1!
1*
b111 6
19
1>
1C
b111 G
#669520000000
0!
0*
09
0>
0C
#669530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#669540000000
0!
0*
09
0>
0C
#669550000000
1!
1*
b1 6
19
1>
1C
b1 G
#669560000000
0!
0*
09
0>
0C
#669570000000
1!
1*
b10 6
19
1>
1C
b10 G
#669580000000
0!
0*
09
0>
0C
#669590000000
1!
1*
b11 6
19
1>
1C
b11 G
#669600000000
0!
0*
09
0>
0C
#669610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#669620000000
0!
0*
09
0>
0C
#669630000000
1!
1*
b101 6
19
1>
1C
b101 G
#669640000000
0!
0*
09
0>
0C
#669650000000
1!
1*
b110 6
19
1>
1C
b110 G
#669660000000
0!
0*
09
0>
0C
#669670000000
1!
1*
b111 6
19
1>
1C
b111 G
#669680000000
0!
0*
09
0>
0C
#669690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#669700000000
0!
0*
09
0>
0C
#669710000000
1!
1*
b1 6
19
1>
1C
b1 G
#669720000000
0!
0*
09
0>
0C
#669730000000
1!
1*
b10 6
19
1>
1C
b10 G
#669740000000
0!
0*
09
0>
0C
#669750000000
1!
1*
b11 6
19
1>
1C
b11 G
#669760000000
0!
0*
09
0>
0C
#669770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#669780000000
0!
0*
09
0>
0C
#669790000000
1!
1*
b101 6
19
1>
1C
b101 G
#669800000000
0!
0*
09
0>
0C
#669810000000
1!
1*
b110 6
19
1>
1C
b110 G
#669820000000
0!
0*
09
0>
0C
#669830000000
1!
1*
b111 6
19
1>
1C
b111 G
#669840000000
0!
1"
0*
1+
09
1:
0>
0C
#669850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#669860000000
0!
0*
09
0>
0C
#669870000000
1!
1*
b1 6
19
1>
1C
b1 G
#669880000000
0!
0*
09
0>
0C
#669890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#669900000000
0!
0*
09
0>
0C
#669910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#669920000000
0!
0*
09
0>
0C
#669930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#669940000000
0!
0*
09
0>
0C
#669950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#669960000000
0!
0#
0*
0,
09
0>
0?
0C
#669970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#669980000000
0!
0*
09
0>
0C
#669990000000
1!
1*
19
1>
1C
#670000000000
0!
0*
09
0>
0C
#670010000000
1!
1*
19
1>
1C
#670020000000
0!
0*
09
0>
0C
#670030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#670040000000
0!
0*
09
0>
0C
#670050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#670060000000
0!
0*
09
0>
0C
#670070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#670080000000
0!
0*
09
0>
0C
#670090000000
1!
1*
b10 6
19
1>
1C
b10 G
#670100000000
0!
0*
09
0>
0C
#670110000000
1!
1*
b11 6
19
1>
1C
b11 G
#670120000000
0!
0*
09
0>
0C
#670130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#670140000000
0!
0*
09
0>
0C
#670150000000
1!
1*
b101 6
19
1>
1C
b101 G
#670160000000
0!
0*
09
0>
0C
#670170000000
1!
1*
b110 6
19
1>
1C
b110 G
#670180000000
0!
0*
09
0>
0C
#670190000000
1!
1*
b111 6
19
1>
1C
b111 G
#670200000000
0!
0*
09
0>
0C
#670210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#670220000000
0!
0*
09
0>
0C
#670230000000
1!
1*
b1 6
19
1>
1C
b1 G
#670240000000
0!
0*
09
0>
0C
#670250000000
1!
1*
b10 6
19
1>
1C
b10 G
#670260000000
0!
0*
09
0>
0C
#670270000000
1!
1*
b11 6
19
1>
1C
b11 G
#670280000000
0!
0*
09
0>
0C
#670290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#670300000000
0!
0*
09
0>
0C
#670310000000
1!
1*
b101 6
19
1>
1C
b101 G
#670320000000
0!
0*
09
0>
0C
#670330000000
1!
1*
b110 6
19
1>
1C
b110 G
#670340000000
0!
0*
09
0>
0C
#670350000000
1!
1*
b111 6
19
1>
1C
b111 G
#670360000000
0!
0*
09
0>
0C
#670370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#670380000000
0!
0*
09
0>
0C
#670390000000
1!
1*
b1 6
19
1>
1C
b1 G
#670400000000
0!
0*
09
0>
0C
#670410000000
1!
1*
b10 6
19
1>
1C
b10 G
#670420000000
0!
0*
09
0>
0C
#670430000000
1!
1*
b11 6
19
1>
1C
b11 G
#670440000000
0!
0*
09
0>
0C
#670450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#670460000000
0!
0*
09
0>
0C
#670470000000
1!
1*
b101 6
19
1>
1C
b101 G
#670480000000
0!
0*
09
0>
0C
#670490000000
1!
1*
b110 6
19
1>
1C
b110 G
#670500000000
0!
0*
09
0>
0C
#670510000000
1!
1*
b111 6
19
1>
1C
b111 G
#670520000000
0!
1"
0*
1+
09
1:
0>
0C
#670530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#670540000000
0!
0*
09
0>
0C
#670550000000
1!
1*
b1 6
19
1>
1C
b1 G
#670560000000
0!
0*
09
0>
0C
#670570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#670580000000
0!
0*
09
0>
0C
#670590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#670600000000
0!
0*
09
0>
0C
#670610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#670620000000
0!
0*
09
0>
0C
#670630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#670640000000
0!
0#
0*
0,
09
0>
0?
0C
#670650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#670660000000
0!
0*
09
0>
0C
#670670000000
1!
1*
19
1>
1C
#670680000000
0!
0*
09
0>
0C
#670690000000
1!
1*
19
1>
1C
#670700000000
0!
0*
09
0>
0C
#670710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#670720000000
0!
0*
09
0>
0C
#670730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#670740000000
0!
0*
09
0>
0C
#670750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#670760000000
0!
0*
09
0>
0C
#670770000000
1!
1*
b10 6
19
1>
1C
b10 G
#670780000000
0!
0*
09
0>
0C
#670790000000
1!
1*
b11 6
19
1>
1C
b11 G
#670800000000
0!
0*
09
0>
0C
#670810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#670820000000
0!
0*
09
0>
0C
#670830000000
1!
1*
b101 6
19
1>
1C
b101 G
#670840000000
0!
0*
09
0>
0C
#670850000000
1!
1*
b110 6
19
1>
1C
b110 G
#670860000000
0!
0*
09
0>
0C
#670870000000
1!
1*
b111 6
19
1>
1C
b111 G
#670880000000
0!
0*
09
0>
0C
#670890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#670900000000
0!
0*
09
0>
0C
#670910000000
1!
1*
b1 6
19
1>
1C
b1 G
#670920000000
0!
0*
09
0>
0C
#670930000000
1!
1*
b10 6
19
1>
1C
b10 G
#670940000000
0!
0*
09
0>
0C
#670950000000
1!
1*
b11 6
19
1>
1C
b11 G
#670960000000
0!
0*
09
0>
0C
#670970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#670980000000
0!
0*
09
0>
0C
#670990000000
1!
1*
b101 6
19
1>
1C
b101 G
#671000000000
0!
0*
09
0>
0C
#671010000000
1!
1*
b110 6
19
1>
1C
b110 G
#671020000000
0!
0*
09
0>
0C
#671030000000
1!
1*
b111 6
19
1>
1C
b111 G
#671040000000
0!
0*
09
0>
0C
#671050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#671060000000
0!
0*
09
0>
0C
#671070000000
1!
1*
b1 6
19
1>
1C
b1 G
#671080000000
0!
0*
09
0>
0C
#671090000000
1!
1*
b10 6
19
1>
1C
b10 G
#671100000000
0!
0*
09
0>
0C
#671110000000
1!
1*
b11 6
19
1>
1C
b11 G
#671120000000
0!
0*
09
0>
0C
#671130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#671140000000
0!
0*
09
0>
0C
#671150000000
1!
1*
b101 6
19
1>
1C
b101 G
#671160000000
0!
0*
09
0>
0C
#671170000000
1!
1*
b110 6
19
1>
1C
b110 G
#671180000000
0!
0*
09
0>
0C
#671190000000
1!
1*
b111 6
19
1>
1C
b111 G
#671200000000
0!
1"
0*
1+
09
1:
0>
0C
#671210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#671220000000
0!
0*
09
0>
0C
#671230000000
1!
1*
b1 6
19
1>
1C
b1 G
#671240000000
0!
0*
09
0>
0C
#671250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#671260000000
0!
0*
09
0>
0C
#671270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#671280000000
0!
0*
09
0>
0C
#671290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#671300000000
0!
0*
09
0>
0C
#671310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#671320000000
0!
0#
0*
0,
09
0>
0?
0C
#671330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#671340000000
0!
0*
09
0>
0C
#671350000000
1!
1*
19
1>
1C
#671360000000
0!
0*
09
0>
0C
#671370000000
1!
1*
19
1>
1C
#671380000000
0!
0*
09
0>
0C
#671390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#671400000000
0!
0*
09
0>
0C
#671410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#671420000000
0!
0*
09
0>
0C
#671430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#671440000000
0!
0*
09
0>
0C
#671450000000
1!
1*
b10 6
19
1>
1C
b10 G
#671460000000
0!
0*
09
0>
0C
#671470000000
1!
1*
b11 6
19
1>
1C
b11 G
#671480000000
0!
0*
09
0>
0C
#671490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#671500000000
0!
0*
09
0>
0C
#671510000000
1!
1*
b101 6
19
1>
1C
b101 G
#671520000000
0!
0*
09
0>
0C
#671530000000
1!
1*
b110 6
19
1>
1C
b110 G
#671540000000
0!
0*
09
0>
0C
#671550000000
1!
1*
b111 6
19
1>
1C
b111 G
#671560000000
0!
0*
09
0>
0C
#671570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#671580000000
0!
0*
09
0>
0C
#671590000000
1!
1*
b1 6
19
1>
1C
b1 G
#671600000000
0!
0*
09
0>
0C
#671610000000
1!
1*
b10 6
19
1>
1C
b10 G
#671620000000
0!
0*
09
0>
0C
#671630000000
1!
1*
b11 6
19
1>
1C
b11 G
#671640000000
0!
0*
09
0>
0C
#671650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#671660000000
0!
0*
09
0>
0C
#671670000000
1!
1*
b101 6
19
1>
1C
b101 G
#671680000000
0!
0*
09
0>
0C
#671690000000
1!
1*
b110 6
19
1>
1C
b110 G
#671700000000
0!
0*
09
0>
0C
#671710000000
1!
1*
b111 6
19
1>
1C
b111 G
#671720000000
0!
0*
09
0>
0C
#671730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#671740000000
0!
0*
09
0>
0C
#671750000000
1!
1*
b1 6
19
1>
1C
b1 G
#671760000000
0!
0*
09
0>
0C
#671770000000
1!
1*
b10 6
19
1>
1C
b10 G
#671780000000
0!
0*
09
0>
0C
#671790000000
1!
1*
b11 6
19
1>
1C
b11 G
#671800000000
0!
0*
09
0>
0C
#671810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#671820000000
0!
0*
09
0>
0C
#671830000000
1!
1*
b101 6
19
1>
1C
b101 G
#671840000000
0!
0*
09
0>
0C
#671850000000
1!
1*
b110 6
19
1>
1C
b110 G
#671860000000
0!
0*
09
0>
0C
#671870000000
1!
1*
b111 6
19
1>
1C
b111 G
#671880000000
0!
1"
0*
1+
09
1:
0>
0C
#671890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#671900000000
0!
0*
09
0>
0C
#671910000000
1!
1*
b1 6
19
1>
1C
b1 G
#671920000000
0!
0*
09
0>
0C
#671930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#671940000000
0!
0*
09
0>
0C
#671950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#671960000000
0!
0*
09
0>
0C
#671970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#671980000000
0!
0*
09
0>
0C
#671990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#672000000000
0!
0#
0*
0,
09
0>
0?
0C
#672010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#672020000000
0!
0*
09
0>
0C
#672030000000
1!
1*
19
1>
1C
#672040000000
0!
0*
09
0>
0C
#672050000000
1!
1*
19
1>
1C
#672060000000
0!
0*
09
0>
0C
#672070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#672080000000
0!
0*
09
0>
0C
#672090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#672100000000
0!
0*
09
0>
0C
#672110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#672120000000
0!
0*
09
0>
0C
#672130000000
1!
1*
b10 6
19
1>
1C
b10 G
#672140000000
0!
0*
09
0>
0C
#672150000000
1!
1*
b11 6
19
1>
1C
b11 G
#672160000000
0!
0*
09
0>
0C
#672170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#672180000000
0!
0*
09
0>
0C
#672190000000
1!
1*
b101 6
19
1>
1C
b101 G
#672200000000
0!
0*
09
0>
0C
#672210000000
1!
1*
b110 6
19
1>
1C
b110 G
#672220000000
0!
0*
09
0>
0C
#672230000000
1!
1*
b111 6
19
1>
1C
b111 G
#672240000000
0!
0*
09
0>
0C
#672250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#672260000000
0!
0*
09
0>
0C
#672270000000
1!
1*
b1 6
19
1>
1C
b1 G
#672280000000
0!
0*
09
0>
0C
#672290000000
1!
1*
b10 6
19
1>
1C
b10 G
#672300000000
0!
0*
09
0>
0C
#672310000000
1!
1*
b11 6
19
1>
1C
b11 G
#672320000000
0!
0*
09
0>
0C
#672330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#672340000000
0!
0*
09
0>
0C
#672350000000
1!
1*
b101 6
19
1>
1C
b101 G
#672360000000
0!
0*
09
0>
0C
#672370000000
1!
1*
b110 6
19
1>
1C
b110 G
#672380000000
0!
0*
09
0>
0C
#672390000000
1!
1*
b111 6
19
1>
1C
b111 G
#672400000000
0!
0*
09
0>
0C
#672410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#672420000000
0!
0*
09
0>
0C
#672430000000
1!
1*
b1 6
19
1>
1C
b1 G
#672440000000
0!
0*
09
0>
0C
#672450000000
1!
1*
b10 6
19
1>
1C
b10 G
#672460000000
0!
0*
09
0>
0C
#672470000000
1!
1*
b11 6
19
1>
1C
b11 G
#672480000000
0!
0*
09
0>
0C
#672490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#672500000000
0!
0*
09
0>
0C
#672510000000
1!
1*
b101 6
19
1>
1C
b101 G
#672520000000
0!
0*
09
0>
0C
#672530000000
1!
1*
b110 6
19
1>
1C
b110 G
#672540000000
0!
0*
09
0>
0C
#672550000000
1!
1*
b111 6
19
1>
1C
b111 G
#672560000000
0!
1"
0*
1+
09
1:
0>
0C
#672570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#672580000000
0!
0*
09
0>
0C
#672590000000
1!
1*
b1 6
19
1>
1C
b1 G
#672600000000
0!
0*
09
0>
0C
#672610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#672620000000
0!
0*
09
0>
0C
#672630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#672640000000
0!
0*
09
0>
0C
#672650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#672660000000
0!
0*
09
0>
0C
#672670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#672680000000
0!
0#
0*
0,
09
0>
0?
0C
#672690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#672700000000
0!
0*
09
0>
0C
#672710000000
1!
1*
19
1>
1C
#672720000000
0!
0*
09
0>
0C
#672730000000
1!
1*
19
1>
1C
#672740000000
0!
0*
09
0>
0C
#672750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#672760000000
0!
0*
09
0>
0C
#672770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#672780000000
0!
0*
09
0>
0C
#672790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#672800000000
0!
0*
09
0>
0C
#672810000000
1!
1*
b10 6
19
1>
1C
b10 G
#672820000000
0!
0*
09
0>
0C
#672830000000
1!
1*
b11 6
19
1>
1C
b11 G
#672840000000
0!
0*
09
0>
0C
#672850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#672860000000
0!
0*
09
0>
0C
#672870000000
1!
1*
b101 6
19
1>
1C
b101 G
#672880000000
0!
0*
09
0>
0C
#672890000000
1!
1*
b110 6
19
1>
1C
b110 G
#672900000000
0!
0*
09
0>
0C
#672910000000
1!
1*
b111 6
19
1>
1C
b111 G
#672920000000
0!
0*
09
0>
0C
#672930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#672940000000
0!
0*
09
0>
0C
#672950000000
1!
1*
b1 6
19
1>
1C
b1 G
#672960000000
0!
0*
09
0>
0C
#672970000000
1!
1*
b10 6
19
1>
1C
b10 G
#672980000000
0!
0*
09
0>
0C
#672990000000
1!
1*
b11 6
19
1>
1C
b11 G
#673000000000
0!
0*
09
0>
0C
#673010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#673020000000
0!
0*
09
0>
0C
#673030000000
1!
1*
b101 6
19
1>
1C
b101 G
#673040000000
0!
0*
09
0>
0C
#673050000000
1!
1*
b110 6
19
1>
1C
b110 G
#673060000000
0!
0*
09
0>
0C
#673070000000
1!
1*
b111 6
19
1>
1C
b111 G
#673080000000
0!
0*
09
0>
0C
#673090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#673100000000
0!
0*
09
0>
0C
#673110000000
1!
1*
b1 6
19
1>
1C
b1 G
#673120000000
0!
0*
09
0>
0C
#673130000000
1!
1*
b10 6
19
1>
1C
b10 G
#673140000000
0!
0*
09
0>
0C
#673150000000
1!
1*
b11 6
19
1>
1C
b11 G
#673160000000
0!
0*
09
0>
0C
#673170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#673180000000
0!
0*
09
0>
0C
#673190000000
1!
1*
b101 6
19
1>
1C
b101 G
#673200000000
0!
0*
09
0>
0C
#673210000000
1!
1*
b110 6
19
1>
1C
b110 G
#673220000000
0!
0*
09
0>
0C
#673230000000
1!
1*
b111 6
19
1>
1C
b111 G
#673240000000
0!
1"
0*
1+
09
1:
0>
0C
#673250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#673260000000
0!
0*
09
0>
0C
#673270000000
1!
1*
b1 6
19
1>
1C
b1 G
#673280000000
0!
0*
09
0>
0C
#673290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#673300000000
0!
0*
09
0>
0C
#673310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#673320000000
0!
0*
09
0>
0C
#673330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#673340000000
0!
0*
09
0>
0C
#673350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#673360000000
0!
0#
0*
0,
09
0>
0?
0C
#673370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#673380000000
0!
0*
09
0>
0C
#673390000000
1!
1*
19
1>
1C
#673400000000
0!
0*
09
0>
0C
#673410000000
1!
1*
19
1>
1C
#673420000000
0!
0*
09
0>
0C
#673430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#673440000000
0!
0*
09
0>
0C
#673450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#673460000000
0!
0*
09
0>
0C
#673470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#673480000000
0!
0*
09
0>
0C
#673490000000
1!
1*
b10 6
19
1>
1C
b10 G
#673500000000
0!
0*
09
0>
0C
#673510000000
1!
1*
b11 6
19
1>
1C
b11 G
#673520000000
0!
0*
09
0>
0C
#673530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#673540000000
0!
0*
09
0>
0C
#673550000000
1!
1*
b101 6
19
1>
1C
b101 G
#673560000000
0!
0*
09
0>
0C
#673570000000
1!
1*
b110 6
19
1>
1C
b110 G
#673580000000
0!
0*
09
0>
0C
#673590000000
1!
1*
b111 6
19
1>
1C
b111 G
#673600000000
0!
0*
09
0>
0C
#673610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#673620000000
0!
0*
09
0>
0C
#673630000000
1!
1*
b1 6
19
1>
1C
b1 G
#673640000000
0!
0*
09
0>
0C
#673650000000
1!
1*
b10 6
19
1>
1C
b10 G
#673660000000
0!
0*
09
0>
0C
#673670000000
1!
1*
b11 6
19
1>
1C
b11 G
#673680000000
0!
0*
09
0>
0C
#673690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#673700000000
0!
0*
09
0>
0C
#673710000000
1!
1*
b101 6
19
1>
1C
b101 G
#673720000000
0!
0*
09
0>
0C
#673730000000
1!
1*
b110 6
19
1>
1C
b110 G
#673740000000
0!
0*
09
0>
0C
#673750000000
1!
1*
b111 6
19
1>
1C
b111 G
#673760000000
0!
0*
09
0>
0C
#673770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#673780000000
0!
0*
09
0>
0C
#673790000000
1!
1*
b1 6
19
1>
1C
b1 G
#673800000000
0!
0*
09
0>
0C
#673810000000
1!
1*
b10 6
19
1>
1C
b10 G
#673820000000
0!
0*
09
0>
0C
#673830000000
1!
1*
b11 6
19
1>
1C
b11 G
#673840000000
0!
0*
09
0>
0C
#673850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#673860000000
0!
0*
09
0>
0C
#673870000000
1!
1*
b101 6
19
1>
1C
b101 G
#673880000000
0!
0*
09
0>
0C
#673890000000
1!
1*
b110 6
19
1>
1C
b110 G
#673900000000
0!
0*
09
0>
0C
#673910000000
1!
1*
b111 6
19
1>
1C
b111 G
#673920000000
0!
1"
0*
1+
09
1:
0>
0C
#673930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#673940000000
0!
0*
09
0>
0C
#673950000000
1!
1*
b1 6
19
1>
1C
b1 G
#673960000000
0!
0*
09
0>
0C
#673970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#673980000000
0!
0*
09
0>
0C
#673990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#674000000000
0!
0*
09
0>
0C
#674010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#674020000000
0!
0*
09
0>
0C
#674030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#674040000000
0!
0#
0*
0,
09
0>
0?
0C
#674050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#674060000000
0!
0*
09
0>
0C
#674070000000
1!
1*
19
1>
1C
#674080000000
0!
0*
09
0>
0C
#674090000000
1!
1*
19
1>
1C
#674100000000
0!
0*
09
0>
0C
#674110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#674120000000
0!
0*
09
0>
0C
#674130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#674140000000
0!
0*
09
0>
0C
#674150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#674160000000
0!
0*
09
0>
0C
#674170000000
1!
1*
b10 6
19
1>
1C
b10 G
#674180000000
0!
0*
09
0>
0C
#674190000000
1!
1*
b11 6
19
1>
1C
b11 G
#674200000000
0!
0*
09
0>
0C
#674210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#674220000000
0!
0*
09
0>
0C
#674230000000
1!
1*
b101 6
19
1>
1C
b101 G
#674240000000
0!
0*
09
0>
0C
#674250000000
1!
1*
b110 6
19
1>
1C
b110 G
#674260000000
0!
0*
09
0>
0C
#674270000000
1!
1*
b111 6
19
1>
1C
b111 G
#674280000000
0!
0*
09
0>
0C
#674290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#674300000000
0!
0*
09
0>
0C
#674310000000
1!
1*
b1 6
19
1>
1C
b1 G
#674320000000
0!
0*
09
0>
0C
#674330000000
1!
1*
b10 6
19
1>
1C
b10 G
#674340000000
0!
0*
09
0>
0C
#674350000000
1!
1*
b11 6
19
1>
1C
b11 G
#674360000000
0!
0*
09
0>
0C
#674370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#674380000000
0!
0*
09
0>
0C
#674390000000
1!
1*
b101 6
19
1>
1C
b101 G
#674400000000
0!
0*
09
0>
0C
#674410000000
1!
1*
b110 6
19
1>
1C
b110 G
#674420000000
0!
0*
09
0>
0C
#674430000000
1!
1*
b111 6
19
1>
1C
b111 G
#674440000000
0!
0*
09
0>
0C
#674450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#674460000000
0!
0*
09
0>
0C
#674470000000
1!
1*
b1 6
19
1>
1C
b1 G
#674480000000
0!
0*
09
0>
0C
#674490000000
1!
1*
b10 6
19
1>
1C
b10 G
#674500000000
0!
0*
09
0>
0C
#674510000000
1!
1*
b11 6
19
1>
1C
b11 G
#674520000000
0!
0*
09
0>
0C
#674530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#674540000000
0!
0*
09
0>
0C
#674550000000
1!
1*
b101 6
19
1>
1C
b101 G
#674560000000
0!
0*
09
0>
0C
#674570000000
1!
1*
b110 6
19
1>
1C
b110 G
#674580000000
0!
0*
09
0>
0C
#674590000000
1!
1*
b111 6
19
1>
1C
b111 G
#674600000000
0!
1"
0*
1+
09
1:
0>
0C
#674610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#674620000000
0!
0*
09
0>
0C
#674630000000
1!
1*
b1 6
19
1>
1C
b1 G
#674640000000
0!
0*
09
0>
0C
#674650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#674660000000
0!
0*
09
0>
0C
#674670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#674680000000
0!
0*
09
0>
0C
#674690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#674700000000
0!
0*
09
0>
0C
#674710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#674720000000
0!
0#
0*
0,
09
0>
0?
0C
#674730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#674740000000
0!
0*
09
0>
0C
#674750000000
1!
1*
19
1>
1C
#674760000000
0!
0*
09
0>
0C
#674770000000
1!
1*
19
1>
1C
#674780000000
0!
0*
09
0>
0C
#674790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#674800000000
0!
0*
09
0>
0C
#674810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#674820000000
0!
0*
09
0>
0C
#674830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#674840000000
0!
0*
09
0>
0C
#674850000000
1!
1*
b10 6
19
1>
1C
b10 G
#674860000000
0!
0*
09
0>
0C
#674870000000
1!
1*
b11 6
19
1>
1C
b11 G
#674880000000
0!
0*
09
0>
0C
#674890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#674900000000
0!
0*
09
0>
0C
#674910000000
1!
1*
b101 6
19
1>
1C
b101 G
#674920000000
0!
0*
09
0>
0C
#674930000000
1!
1*
b110 6
19
1>
1C
b110 G
#674940000000
0!
0*
09
0>
0C
#674950000000
1!
1*
b111 6
19
1>
1C
b111 G
#674960000000
0!
0*
09
0>
0C
#674970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#674980000000
0!
0*
09
0>
0C
#674990000000
1!
1*
b1 6
19
1>
1C
b1 G
#675000000000
0!
0*
09
0>
0C
#675010000000
1!
1*
b10 6
19
1>
1C
b10 G
#675020000000
0!
0*
09
0>
0C
#675030000000
1!
1*
b11 6
19
1>
1C
b11 G
#675040000000
0!
0*
09
0>
0C
#675050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#675060000000
0!
0*
09
0>
0C
#675070000000
1!
1*
b101 6
19
1>
1C
b101 G
#675080000000
0!
0*
09
0>
0C
#675090000000
1!
1*
b110 6
19
1>
1C
b110 G
#675100000000
0!
0*
09
0>
0C
#675110000000
1!
1*
b111 6
19
1>
1C
b111 G
#675120000000
0!
0*
09
0>
0C
#675130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#675140000000
0!
0*
09
0>
0C
#675150000000
1!
1*
b1 6
19
1>
1C
b1 G
#675160000000
0!
0*
09
0>
0C
#675170000000
1!
1*
b10 6
19
1>
1C
b10 G
#675180000000
0!
0*
09
0>
0C
#675190000000
1!
1*
b11 6
19
1>
1C
b11 G
#675200000000
0!
0*
09
0>
0C
#675210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#675220000000
0!
0*
09
0>
0C
#675230000000
1!
1*
b101 6
19
1>
1C
b101 G
#675240000000
0!
0*
09
0>
0C
#675250000000
1!
1*
b110 6
19
1>
1C
b110 G
#675260000000
0!
0*
09
0>
0C
#675270000000
1!
1*
b111 6
19
1>
1C
b111 G
#675280000000
0!
1"
0*
1+
09
1:
0>
0C
#675290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#675300000000
0!
0*
09
0>
0C
#675310000000
1!
1*
b1 6
19
1>
1C
b1 G
#675320000000
0!
0*
09
0>
0C
#675330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#675340000000
0!
0*
09
0>
0C
#675350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#675360000000
0!
0*
09
0>
0C
#675370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#675380000000
0!
0*
09
0>
0C
#675390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#675400000000
0!
0#
0*
0,
09
0>
0?
0C
#675410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#675420000000
0!
0*
09
0>
0C
#675430000000
1!
1*
19
1>
1C
#675440000000
0!
0*
09
0>
0C
#675450000000
1!
1*
19
1>
1C
#675460000000
0!
0*
09
0>
0C
#675470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#675480000000
0!
0*
09
0>
0C
#675490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#675500000000
0!
0*
09
0>
0C
#675510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#675520000000
0!
0*
09
0>
0C
#675530000000
1!
1*
b10 6
19
1>
1C
b10 G
#675540000000
0!
0*
09
0>
0C
#675550000000
1!
1*
b11 6
19
1>
1C
b11 G
#675560000000
0!
0*
09
0>
0C
#675570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#675580000000
0!
0*
09
0>
0C
#675590000000
1!
1*
b101 6
19
1>
1C
b101 G
#675600000000
0!
0*
09
0>
0C
#675610000000
1!
1*
b110 6
19
1>
1C
b110 G
#675620000000
0!
0*
09
0>
0C
#675630000000
1!
1*
b111 6
19
1>
1C
b111 G
#675640000000
0!
0*
09
0>
0C
#675650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#675660000000
0!
0*
09
0>
0C
#675670000000
1!
1*
b1 6
19
1>
1C
b1 G
#675680000000
0!
0*
09
0>
0C
#675690000000
1!
1*
b10 6
19
1>
1C
b10 G
#675700000000
0!
0*
09
0>
0C
#675710000000
1!
1*
b11 6
19
1>
1C
b11 G
#675720000000
0!
0*
09
0>
0C
#675730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#675740000000
0!
0*
09
0>
0C
#675750000000
1!
1*
b101 6
19
1>
1C
b101 G
#675760000000
0!
0*
09
0>
0C
#675770000000
1!
1*
b110 6
19
1>
1C
b110 G
#675780000000
0!
0*
09
0>
0C
#675790000000
1!
1*
b111 6
19
1>
1C
b111 G
#675800000000
0!
0*
09
0>
0C
#675810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#675820000000
0!
0*
09
0>
0C
#675830000000
1!
1*
b1 6
19
1>
1C
b1 G
#675840000000
0!
0*
09
0>
0C
#675850000000
1!
1*
b10 6
19
1>
1C
b10 G
#675860000000
0!
0*
09
0>
0C
#675870000000
1!
1*
b11 6
19
1>
1C
b11 G
#675880000000
0!
0*
09
0>
0C
#675890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#675900000000
0!
0*
09
0>
0C
#675910000000
1!
1*
b101 6
19
1>
1C
b101 G
#675920000000
0!
0*
09
0>
0C
#675930000000
1!
1*
b110 6
19
1>
1C
b110 G
#675940000000
0!
0*
09
0>
0C
#675950000000
1!
1*
b111 6
19
1>
1C
b111 G
#675960000000
0!
1"
0*
1+
09
1:
0>
0C
#675970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#675980000000
0!
0*
09
0>
0C
#675990000000
1!
1*
b1 6
19
1>
1C
b1 G
#676000000000
0!
0*
09
0>
0C
#676010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#676020000000
0!
0*
09
0>
0C
#676030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#676040000000
0!
0*
09
0>
0C
#676050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#676060000000
0!
0*
09
0>
0C
#676070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#676080000000
0!
0#
0*
0,
09
0>
0?
0C
#676090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#676100000000
0!
0*
09
0>
0C
#676110000000
1!
1*
19
1>
1C
#676120000000
0!
0*
09
0>
0C
#676130000000
1!
1*
19
1>
1C
#676140000000
0!
0*
09
0>
0C
#676150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#676160000000
0!
0*
09
0>
0C
#676170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#676180000000
0!
0*
09
0>
0C
#676190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#676200000000
0!
0*
09
0>
0C
#676210000000
1!
1*
b10 6
19
1>
1C
b10 G
#676220000000
0!
0*
09
0>
0C
#676230000000
1!
1*
b11 6
19
1>
1C
b11 G
#676240000000
0!
0*
09
0>
0C
#676250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#676260000000
0!
0*
09
0>
0C
#676270000000
1!
1*
b101 6
19
1>
1C
b101 G
#676280000000
0!
0*
09
0>
0C
#676290000000
1!
1*
b110 6
19
1>
1C
b110 G
#676300000000
0!
0*
09
0>
0C
#676310000000
1!
1*
b111 6
19
1>
1C
b111 G
#676320000000
0!
0*
09
0>
0C
#676330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#676340000000
0!
0*
09
0>
0C
#676350000000
1!
1*
b1 6
19
1>
1C
b1 G
#676360000000
0!
0*
09
0>
0C
#676370000000
1!
1*
b10 6
19
1>
1C
b10 G
#676380000000
0!
0*
09
0>
0C
#676390000000
1!
1*
b11 6
19
1>
1C
b11 G
#676400000000
0!
0*
09
0>
0C
#676410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#676420000000
0!
0*
09
0>
0C
#676430000000
1!
1*
b101 6
19
1>
1C
b101 G
#676440000000
0!
0*
09
0>
0C
#676450000000
1!
1*
b110 6
19
1>
1C
b110 G
#676460000000
0!
0*
09
0>
0C
#676470000000
1!
1*
b111 6
19
1>
1C
b111 G
#676480000000
0!
0*
09
0>
0C
#676490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#676500000000
0!
0*
09
0>
0C
#676510000000
1!
1*
b1 6
19
1>
1C
b1 G
#676520000000
0!
0*
09
0>
0C
#676530000000
1!
1*
b10 6
19
1>
1C
b10 G
#676540000000
0!
0*
09
0>
0C
#676550000000
1!
1*
b11 6
19
1>
1C
b11 G
#676560000000
0!
0*
09
0>
0C
#676570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#676580000000
0!
0*
09
0>
0C
#676590000000
1!
1*
b101 6
19
1>
1C
b101 G
#676600000000
0!
0*
09
0>
0C
#676610000000
1!
1*
b110 6
19
1>
1C
b110 G
#676620000000
0!
0*
09
0>
0C
#676630000000
1!
1*
b111 6
19
1>
1C
b111 G
#676640000000
0!
1"
0*
1+
09
1:
0>
0C
#676650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#676660000000
0!
0*
09
0>
0C
#676670000000
1!
1*
b1 6
19
1>
1C
b1 G
#676680000000
0!
0*
09
0>
0C
#676690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#676700000000
0!
0*
09
0>
0C
#676710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#676720000000
0!
0*
09
0>
0C
#676730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#676740000000
0!
0*
09
0>
0C
#676750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#676760000000
0!
0#
0*
0,
09
0>
0?
0C
#676770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#676780000000
0!
0*
09
0>
0C
#676790000000
1!
1*
19
1>
1C
#676800000000
0!
0*
09
0>
0C
#676810000000
1!
1*
19
1>
1C
#676820000000
0!
0*
09
0>
0C
#676830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#676840000000
0!
0*
09
0>
0C
#676850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#676860000000
0!
0*
09
0>
0C
#676870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#676880000000
0!
0*
09
0>
0C
#676890000000
1!
1*
b10 6
19
1>
1C
b10 G
#676900000000
0!
0*
09
0>
0C
#676910000000
1!
1*
b11 6
19
1>
1C
b11 G
#676920000000
0!
0*
09
0>
0C
#676930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#676940000000
0!
0*
09
0>
0C
#676950000000
1!
1*
b101 6
19
1>
1C
b101 G
#676960000000
0!
0*
09
0>
0C
#676970000000
1!
1*
b110 6
19
1>
1C
b110 G
#676980000000
0!
0*
09
0>
0C
#676990000000
1!
1*
b111 6
19
1>
1C
b111 G
#677000000000
0!
0*
09
0>
0C
#677010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#677020000000
0!
0*
09
0>
0C
#677030000000
1!
1*
b1 6
19
1>
1C
b1 G
#677040000000
0!
0*
09
0>
0C
#677050000000
1!
1*
b10 6
19
1>
1C
b10 G
#677060000000
0!
0*
09
0>
0C
#677070000000
1!
1*
b11 6
19
1>
1C
b11 G
#677080000000
0!
0*
09
0>
0C
#677090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#677100000000
0!
0*
09
0>
0C
#677110000000
1!
1*
b101 6
19
1>
1C
b101 G
#677120000000
0!
0*
09
0>
0C
#677130000000
1!
1*
b110 6
19
1>
1C
b110 G
#677140000000
0!
0*
09
0>
0C
#677150000000
1!
1*
b111 6
19
1>
1C
b111 G
#677160000000
0!
0*
09
0>
0C
#677170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#677180000000
0!
0*
09
0>
0C
#677190000000
1!
1*
b1 6
19
1>
1C
b1 G
#677200000000
0!
0*
09
0>
0C
#677210000000
1!
1*
b10 6
19
1>
1C
b10 G
#677220000000
0!
0*
09
0>
0C
#677230000000
1!
1*
b11 6
19
1>
1C
b11 G
#677240000000
0!
0*
09
0>
0C
#677250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#677260000000
0!
0*
09
0>
0C
#677270000000
1!
1*
b101 6
19
1>
1C
b101 G
#677280000000
0!
0*
09
0>
0C
#677290000000
1!
1*
b110 6
19
1>
1C
b110 G
#677300000000
0!
0*
09
0>
0C
#677310000000
1!
1*
b111 6
19
1>
1C
b111 G
#677320000000
0!
1"
0*
1+
09
1:
0>
0C
#677330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#677340000000
0!
0*
09
0>
0C
#677350000000
1!
1*
b1 6
19
1>
1C
b1 G
#677360000000
0!
0*
09
0>
0C
#677370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#677380000000
0!
0*
09
0>
0C
#677390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#677400000000
0!
0*
09
0>
0C
#677410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#677420000000
0!
0*
09
0>
0C
#677430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#677440000000
0!
0#
0*
0,
09
0>
0?
0C
#677450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#677460000000
0!
0*
09
0>
0C
#677470000000
1!
1*
19
1>
1C
#677480000000
0!
0*
09
0>
0C
#677490000000
1!
1*
19
1>
1C
#677500000000
0!
0*
09
0>
0C
#677510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#677520000000
0!
0*
09
0>
0C
#677530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#677540000000
0!
0*
09
0>
0C
#677550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#677560000000
0!
0*
09
0>
0C
#677570000000
1!
1*
b10 6
19
1>
1C
b10 G
#677580000000
0!
0*
09
0>
0C
#677590000000
1!
1*
b11 6
19
1>
1C
b11 G
#677600000000
0!
0*
09
0>
0C
#677610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#677620000000
0!
0*
09
0>
0C
#677630000000
1!
1*
b101 6
19
1>
1C
b101 G
#677640000000
0!
0*
09
0>
0C
#677650000000
1!
1*
b110 6
19
1>
1C
b110 G
#677660000000
0!
0*
09
0>
0C
#677670000000
1!
1*
b111 6
19
1>
1C
b111 G
#677680000000
0!
0*
09
0>
0C
#677690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#677700000000
0!
0*
09
0>
0C
#677710000000
1!
1*
b1 6
19
1>
1C
b1 G
#677720000000
0!
0*
09
0>
0C
#677730000000
1!
1*
b10 6
19
1>
1C
b10 G
#677740000000
0!
0*
09
0>
0C
#677750000000
1!
1*
b11 6
19
1>
1C
b11 G
#677760000000
0!
0*
09
0>
0C
#677770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#677780000000
0!
0*
09
0>
0C
#677790000000
1!
1*
b101 6
19
1>
1C
b101 G
#677800000000
0!
0*
09
0>
0C
#677810000000
1!
1*
b110 6
19
1>
1C
b110 G
#677820000000
0!
0*
09
0>
0C
#677830000000
1!
1*
b111 6
19
1>
1C
b111 G
#677840000000
0!
0*
09
0>
0C
#677850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#677860000000
0!
0*
09
0>
0C
#677870000000
1!
1*
b1 6
19
1>
1C
b1 G
#677880000000
0!
0*
09
0>
0C
#677890000000
1!
1*
b10 6
19
1>
1C
b10 G
#677900000000
0!
0*
09
0>
0C
#677910000000
1!
1*
b11 6
19
1>
1C
b11 G
#677920000000
0!
0*
09
0>
0C
#677930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#677940000000
0!
0*
09
0>
0C
#677950000000
1!
1*
b101 6
19
1>
1C
b101 G
#677960000000
0!
0*
09
0>
0C
#677970000000
1!
1*
b110 6
19
1>
1C
b110 G
#677980000000
0!
0*
09
0>
0C
#677990000000
1!
1*
b111 6
19
1>
1C
b111 G
#678000000000
0!
1"
0*
1+
09
1:
0>
0C
#678010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#678020000000
0!
0*
09
0>
0C
#678030000000
1!
1*
b1 6
19
1>
1C
b1 G
#678040000000
0!
0*
09
0>
0C
#678050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#678060000000
0!
0*
09
0>
0C
#678070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#678080000000
0!
0*
09
0>
0C
#678090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#678100000000
0!
0*
09
0>
0C
#678110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#678120000000
0!
0#
0*
0,
09
0>
0?
0C
#678130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#678140000000
0!
0*
09
0>
0C
#678150000000
1!
1*
19
1>
1C
#678160000000
0!
0*
09
0>
0C
#678170000000
1!
1*
19
1>
1C
#678180000000
0!
0*
09
0>
0C
#678190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#678200000000
0!
0*
09
0>
0C
#678210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#678220000000
0!
0*
09
0>
0C
#678230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#678240000000
0!
0*
09
0>
0C
#678250000000
1!
1*
b10 6
19
1>
1C
b10 G
#678260000000
0!
0*
09
0>
0C
#678270000000
1!
1*
b11 6
19
1>
1C
b11 G
#678280000000
0!
0*
09
0>
0C
#678290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#678300000000
0!
0*
09
0>
0C
#678310000000
1!
1*
b101 6
19
1>
1C
b101 G
#678320000000
0!
0*
09
0>
0C
#678330000000
1!
1*
b110 6
19
1>
1C
b110 G
#678340000000
0!
0*
09
0>
0C
#678350000000
1!
1*
b111 6
19
1>
1C
b111 G
#678360000000
0!
0*
09
0>
0C
#678370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#678380000000
0!
0*
09
0>
0C
#678390000000
1!
1*
b1 6
19
1>
1C
b1 G
#678400000000
0!
0*
09
0>
0C
#678410000000
1!
1*
b10 6
19
1>
1C
b10 G
#678420000000
0!
0*
09
0>
0C
#678430000000
1!
1*
b11 6
19
1>
1C
b11 G
#678440000000
0!
0*
09
0>
0C
#678450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#678460000000
0!
0*
09
0>
0C
#678470000000
1!
1*
b101 6
19
1>
1C
b101 G
#678480000000
0!
0*
09
0>
0C
#678490000000
1!
1*
b110 6
19
1>
1C
b110 G
#678500000000
0!
0*
09
0>
0C
#678510000000
1!
1*
b111 6
19
1>
1C
b111 G
#678520000000
0!
0*
09
0>
0C
#678530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#678540000000
0!
0*
09
0>
0C
#678550000000
1!
1*
b1 6
19
1>
1C
b1 G
#678560000000
0!
0*
09
0>
0C
#678570000000
1!
1*
b10 6
19
1>
1C
b10 G
#678580000000
0!
0*
09
0>
0C
#678590000000
1!
1*
b11 6
19
1>
1C
b11 G
#678600000000
0!
0*
09
0>
0C
#678610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#678620000000
0!
0*
09
0>
0C
#678630000000
1!
1*
b101 6
19
1>
1C
b101 G
#678640000000
0!
0*
09
0>
0C
#678650000000
1!
1*
b110 6
19
1>
1C
b110 G
#678660000000
0!
0*
09
0>
0C
#678670000000
1!
1*
b111 6
19
1>
1C
b111 G
#678680000000
0!
1"
0*
1+
09
1:
0>
0C
#678690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#678700000000
0!
0*
09
0>
0C
#678710000000
1!
1*
b1 6
19
1>
1C
b1 G
#678720000000
0!
0*
09
0>
0C
#678730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#678740000000
0!
0*
09
0>
0C
#678750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#678760000000
0!
0*
09
0>
0C
#678770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#678780000000
0!
0*
09
0>
0C
#678790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#678800000000
0!
0#
0*
0,
09
0>
0?
0C
#678810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#678820000000
0!
0*
09
0>
0C
#678830000000
1!
1*
19
1>
1C
#678840000000
0!
0*
09
0>
0C
#678850000000
1!
1*
19
1>
1C
#678860000000
0!
0*
09
0>
0C
#678870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#678880000000
0!
0*
09
0>
0C
#678890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#678900000000
0!
0*
09
0>
0C
#678910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#678920000000
0!
0*
09
0>
0C
#678930000000
1!
1*
b10 6
19
1>
1C
b10 G
#678940000000
0!
0*
09
0>
0C
#678950000000
1!
1*
b11 6
19
1>
1C
b11 G
#678960000000
0!
0*
09
0>
0C
#678970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#678980000000
0!
0*
09
0>
0C
#678990000000
1!
1*
b101 6
19
1>
1C
b101 G
#679000000000
0!
0*
09
0>
0C
#679010000000
1!
1*
b110 6
19
1>
1C
b110 G
#679020000000
0!
0*
09
0>
0C
#679030000000
1!
1*
b111 6
19
1>
1C
b111 G
#679040000000
0!
0*
09
0>
0C
#679050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#679060000000
0!
0*
09
0>
0C
#679070000000
1!
1*
b1 6
19
1>
1C
b1 G
#679080000000
0!
0*
09
0>
0C
#679090000000
1!
1*
b10 6
19
1>
1C
b10 G
#679100000000
0!
0*
09
0>
0C
#679110000000
1!
1*
b11 6
19
1>
1C
b11 G
#679120000000
0!
0*
09
0>
0C
#679130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#679140000000
0!
0*
09
0>
0C
#679150000000
1!
1*
b101 6
19
1>
1C
b101 G
#679160000000
0!
0*
09
0>
0C
#679170000000
1!
1*
b110 6
19
1>
1C
b110 G
#679180000000
0!
0*
09
0>
0C
#679190000000
1!
1*
b111 6
19
1>
1C
b111 G
#679200000000
0!
0*
09
0>
0C
#679210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#679220000000
0!
0*
09
0>
0C
#679230000000
1!
1*
b1 6
19
1>
1C
b1 G
#679240000000
0!
0*
09
0>
0C
#679250000000
1!
1*
b10 6
19
1>
1C
b10 G
#679260000000
0!
0*
09
0>
0C
#679270000000
1!
1*
b11 6
19
1>
1C
b11 G
#679280000000
0!
0*
09
0>
0C
#679290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#679300000000
0!
0*
09
0>
0C
#679310000000
1!
1*
b101 6
19
1>
1C
b101 G
#679320000000
0!
0*
09
0>
0C
#679330000000
1!
1*
b110 6
19
1>
1C
b110 G
#679340000000
0!
0*
09
0>
0C
#679350000000
1!
1*
b111 6
19
1>
1C
b111 G
#679360000000
0!
1"
0*
1+
09
1:
0>
0C
#679370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#679380000000
0!
0*
09
0>
0C
#679390000000
1!
1*
b1 6
19
1>
1C
b1 G
#679400000000
0!
0*
09
0>
0C
#679410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#679420000000
0!
0*
09
0>
0C
#679430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#679440000000
0!
0*
09
0>
0C
#679450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#679460000000
0!
0*
09
0>
0C
#679470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#679480000000
0!
0#
0*
0,
09
0>
0?
0C
#679490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#679500000000
0!
0*
09
0>
0C
#679510000000
1!
1*
19
1>
1C
#679520000000
0!
0*
09
0>
0C
#679530000000
1!
1*
19
1>
1C
#679540000000
0!
0*
09
0>
0C
#679550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#679560000000
0!
0*
09
0>
0C
#679570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#679580000000
0!
0*
09
0>
0C
#679590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#679600000000
0!
0*
09
0>
0C
#679610000000
1!
1*
b10 6
19
1>
1C
b10 G
#679620000000
0!
0*
09
0>
0C
#679630000000
1!
1*
b11 6
19
1>
1C
b11 G
#679640000000
0!
0*
09
0>
0C
#679650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#679660000000
0!
0*
09
0>
0C
#679670000000
1!
1*
b101 6
19
1>
1C
b101 G
#679680000000
0!
0*
09
0>
0C
#679690000000
1!
1*
b110 6
19
1>
1C
b110 G
#679700000000
0!
0*
09
0>
0C
#679710000000
1!
1*
b111 6
19
1>
1C
b111 G
#679720000000
0!
0*
09
0>
0C
#679730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#679740000000
0!
0*
09
0>
0C
#679750000000
1!
1*
b1 6
19
1>
1C
b1 G
#679760000000
0!
0*
09
0>
0C
#679770000000
1!
1*
b10 6
19
1>
1C
b10 G
#679780000000
0!
0*
09
0>
0C
#679790000000
1!
1*
b11 6
19
1>
1C
b11 G
#679800000000
0!
0*
09
0>
0C
#679810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#679820000000
0!
0*
09
0>
0C
#679830000000
1!
1*
b101 6
19
1>
1C
b101 G
#679840000000
0!
0*
09
0>
0C
#679850000000
1!
1*
b110 6
19
1>
1C
b110 G
#679860000000
0!
0*
09
0>
0C
#679870000000
1!
1*
b111 6
19
1>
1C
b111 G
#679880000000
0!
0*
09
0>
0C
#679890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#679900000000
0!
0*
09
0>
0C
#679910000000
1!
1*
b1 6
19
1>
1C
b1 G
#679920000000
0!
0*
09
0>
0C
#679930000000
1!
1*
b10 6
19
1>
1C
b10 G
#679940000000
0!
0*
09
0>
0C
#679950000000
1!
1*
b11 6
19
1>
1C
b11 G
#679960000000
0!
0*
09
0>
0C
#679970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#679980000000
0!
0*
09
0>
0C
#679990000000
1!
1*
b101 6
19
1>
1C
b101 G
#680000000000
0!
0*
09
0>
0C
#680010000000
1!
1*
b110 6
19
1>
1C
b110 G
#680020000000
0!
0*
09
0>
0C
#680030000000
1!
1*
b111 6
19
1>
1C
b111 G
#680040000000
0!
1"
0*
1+
09
1:
0>
0C
#680050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#680060000000
0!
0*
09
0>
0C
#680070000000
1!
1*
b1 6
19
1>
1C
b1 G
#680080000000
0!
0*
09
0>
0C
#680090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#680100000000
0!
0*
09
0>
0C
#680110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#680120000000
0!
0*
09
0>
0C
#680130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#680140000000
0!
0*
09
0>
0C
#680150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#680160000000
0!
0#
0*
0,
09
0>
0?
0C
#680170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#680180000000
0!
0*
09
0>
0C
#680190000000
1!
1*
19
1>
1C
#680200000000
0!
0*
09
0>
0C
#680210000000
1!
1*
19
1>
1C
#680220000000
0!
0*
09
0>
0C
#680230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#680240000000
0!
0*
09
0>
0C
#680250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#680260000000
0!
0*
09
0>
0C
#680270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#680280000000
0!
0*
09
0>
0C
#680290000000
1!
1*
b10 6
19
1>
1C
b10 G
#680300000000
0!
0*
09
0>
0C
#680310000000
1!
1*
b11 6
19
1>
1C
b11 G
#680320000000
0!
0*
09
0>
0C
#680330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#680340000000
0!
0*
09
0>
0C
#680350000000
1!
1*
b101 6
19
1>
1C
b101 G
#680360000000
0!
0*
09
0>
0C
#680370000000
1!
1*
b110 6
19
1>
1C
b110 G
#680380000000
0!
0*
09
0>
0C
#680390000000
1!
1*
b111 6
19
1>
1C
b111 G
#680400000000
0!
0*
09
0>
0C
#680410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#680420000000
0!
0*
09
0>
0C
#680430000000
1!
1*
b1 6
19
1>
1C
b1 G
#680440000000
0!
0*
09
0>
0C
#680450000000
1!
1*
b10 6
19
1>
1C
b10 G
#680460000000
0!
0*
09
0>
0C
#680470000000
1!
1*
b11 6
19
1>
1C
b11 G
#680480000000
0!
0*
09
0>
0C
#680490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#680500000000
0!
0*
09
0>
0C
#680510000000
1!
1*
b101 6
19
1>
1C
b101 G
#680520000000
0!
0*
09
0>
0C
#680530000000
1!
1*
b110 6
19
1>
1C
b110 G
#680540000000
0!
0*
09
0>
0C
#680550000000
1!
1*
b111 6
19
1>
1C
b111 G
#680560000000
0!
0*
09
0>
0C
#680570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#680580000000
0!
0*
09
0>
0C
#680590000000
1!
1*
b1 6
19
1>
1C
b1 G
#680600000000
0!
0*
09
0>
0C
#680610000000
1!
1*
b10 6
19
1>
1C
b10 G
#680620000000
0!
0*
09
0>
0C
#680630000000
1!
1*
b11 6
19
1>
1C
b11 G
#680640000000
0!
0*
09
0>
0C
#680650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#680660000000
0!
0*
09
0>
0C
#680670000000
1!
1*
b101 6
19
1>
1C
b101 G
#680680000000
0!
0*
09
0>
0C
#680690000000
1!
1*
b110 6
19
1>
1C
b110 G
#680700000000
0!
0*
09
0>
0C
#680710000000
1!
1*
b111 6
19
1>
1C
b111 G
#680720000000
0!
1"
0*
1+
09
1:
0>
0C
#680730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#680740000000
0!
0*
09
0>
0C
#680750000000
1!
1*
b1 6
19
1>
1C
b1 G
#680760000000
0!
0*
09
0>
0C
#680770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#680780000000
0!
0*
09
0>
0C
#680790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#680800000000
0!
0*
09
0>
0C
#680810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#680820000000
0!
0*
09
0>
0C
#680830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#680840000000
0!
0#
0*
0,
09
0>
0?
0C
#680850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#680860000000
0!
0*
09
0>
0C
#680870000000
1!
1*
19
1>
1C
#680880000000
0!
0*
09
0>
0C
#680890000000
1!
1*
19
1>
1C
#680900000000
0!
0*
09
0>
0C
#680910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#680920000000
0!
0*
09
0>
0C
#680930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#680940000000
0!
0*
09
0>
0C
#680950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#680960000000
0!
0*
09
0>
0C
#680970000000
1!
1*
b10 6
19
1>
1C
b10 G
#680980000000
0!
0*
09
0>
0C
#680990000000
1!
1*
b11 6
19
1>
1C
b11 G
#681000000000
0!
0*
09
0>
0C
#681010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#681020000000
0!
0*
09
0>
0C
#681030000000
1!
1*
b101 6
19
1>
1C
b101 G
#681040000000
0!
0*
09
0>
0C
#681050000000
1!
1*
b110 6
19
1>
1C
b110 G
#681060000000
0!
0*
09
0>
0C
#681070000000
1!
1*
b111 6
19
1>
1C
b111 G
#681080000000
0!
0*
09
0>
0C
#681090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#681100000000
0!
0*
09
0>
0C
#681110000000
1!
1*
b1 6
19
1>
1C
b1 G
#681120000000
0!
0*
09
0>
0C
#681130000000
1!
1*
b10 6
19
1>
1C
b10 G
#681140000000
0!
0*
09
0>
0C
#681150000000
1!
1*
b11 6
19
1>
1C
b11 G
#681160000000
0!
0*
09
0>
0C
#681170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#681180000000
0!
0*
09
0>
0C
#681190000000
1!
1*
b101 6
19
1>
1C
b101 G
#681200000000
0!
0*
09
0>
0C
#681210000000
1!
1*
b110 6
19
1>
1C
b110 G
#681220000000
0!
0*
09
0>
0C
#681230000000
1!
1*
b111 6
19
1>
1C
b111 G
#681240000000
0!
0*
09
0>
0C
#681250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#681260000000
0!
0*
09
0>
0C
#681270000000
1!
1*
b1 6
19
1>
1C
b1 G
#681280000000
0!
0*
09
0>
0C
#681290000000
1!
1*
b10 6
19
1>
1C
b10 G
#681300000000
0!
0*
09
0>
0C
#681310000000
1!
1*
b11 6
19
1>
1C
b11 G
#681320000000
0!
0*
09
0>
0C
#681330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#681340000000
0!
0*
09
0>
0C
#681350000000
1!
1*
b101 6
19
1>
1C
b101 G
#681360000000
0!
0*
09
0>
0C
#681370000000
1!
1*
b110 6
19
1>
1C
b110 G
#681380000000
0!
0*
09
0>
0C
#681390000000
1!
1*
b111 6
19
1>
1C
b111 G
#681400000000
0!
1"
0*
1+
09
1:
0>
0C
#681410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#681420000000
0!
0*
09
0>
0C
#681430000000
1!
1*
b1 6
19
1>
1C
b1 G
#681440000000
0!
0*
09
0>
0C
#681450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#681460000000
0!
0*
09
0>
0C
#681470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#681480000000
0!
0*
09
0>
0C
#681490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#681500000000
0!
0*
09
0>
0C
#681510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#681520000000
0!
0#
0*
0,
09
0>
0?
0C
#681530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#681540000000
0!
0*
09
0>
0C
#681550000000
1!
1*
19
1>
1C
#681560000000
0!
0*
09
0>
0C
#681570000000
1!
1*
19
1>
1C
#681580000000
0!
0*
09
0>
0C
#681590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#681600000000
0!
0*
09
0>
0C
#681610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#681620000000
0!
0*
09
0>
0C
#681630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#681640000000
0!
0*
09
0>
0C
#681650000000
1!
1*
b10 6
19
1>
1C
b10 G
#681660000000
0!
0*
09
0>
0C
#681670000000
1!
1*
b11 6
19
1>
1C
b11 G
#681680000000
0!
0*
09
0>
0C
#681690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#681700000000
0!
0*
09
0>
0C
#681710000000
1!
1*
b101 6
19
1>
1C
b101 G
#681720000000
0!
0*
09
0>
0C
#681730000000
1!
1*
b110 6
19
1>
1C
b110 G
#681740000000
0!
0*
09
0>
0C
#681750000000
1!
1*
b111 6
19
1>
1C
b111 G
#681760000000
0!
0*
09
0>
0C
#681770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#681780000000
0!
0*
09
0>
0C
#681790000000
1!
1*
b1 6
19
1>
1C
b1 G
#681800000000
0!
0*
09
0>
0C
#681810000000
1!
1*
b10 6
19
1>
1C
b10 G
#681820000000
0!
0*
09
0>
0C
#681830000000
1!
1*
b11 6
19
1>
1C
b11 G
#681840000000
0!
0*
09
0>
0C
#681850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#681860000000
0!
0*
09
0>
0C
#681870000000
1!
1*
b101 6
19
1>
1C
b101 G
#681880000000
0!
0*
09
0>
0C
#681890000000
1!
1*
b110 6
19
1>
1C
b110 G
#681900000000
0!
0*
09
0>
0C
#681910000000
1!
1*
b111 6
19
1>
1C
b111 G
#681920000000
0!
0*
09
0>
0C
#681930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#681940000000
0!
0*
09
0>
0C
#681950000000
1!
1*
b1 6
19
1>
1C
b1 G
#681960000000
0!
0*
09
0>
0C
#681970000000
1!
1*
b10 6
19
1>
1C
b10 G
#681980000000
0!
0*
09
0>
0C
#681990000000
1!
1*
b11 6
19
1>
1C
b11 G
#682000000000
0!
0*
09
0>
0C
#682010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#682020000000
0!
0*
09
0>
0C
#682030000000
1!
1*
b101 6
19
1>
1C
b101 G
#682040000000
0!
0*
09
0>
0C
#682050000000
1!
1*
b110 6
19
1>
1C
b110 G
#682060000000
0!
0*
09
0>
0C
#682070000000
1!
1*
b111 6
19
1>
1C
b111 G
#682080000000
0!
1"
0*
1+
09
1:
0>
0C
#682090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#682100000000
0!
0*
09
0>
0C
#682110000000
1!
1*
b1 6
19
1>
1C
b1 G
#682120000000
0!
0*
09
0>
0C
#682130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#682140000000
0!
0*
09
0>
0C
#682150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#682160000000
0!
0*
09
0>
0C
#682170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#682180000000
0!
0*
09
0>
0C
#682190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#682200000000
0!
0#
0*
0,
09
0>
0?
0C
#682210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#682220000000
0!
0*
09
0>
0C
#682230000000
1!
1*
19
1>
1C
#682240000000
0!
0*
09
0>
0C
#682250000000
1!
1*
19
1>
1C
#682260000000
0!
0*
09
0>
0C
#682270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#682280000000
0!
0*
09
0>
0C
#682290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#682300000000
0!
0*
09
0>
0C
#682310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#682320000000
0!
0*
09
0>
0C
#682330000000
1!
1*
b10 6
19
1>
1C
b10 G
#682340000000
0!
0*
09
0>
0C
#682350000000
1!
1*
b11 6
19
1>
1C
b11 G
#682360000000
0!
0*
09
0>
0C
#682370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#682380000000
0!
0*
09
0>
0C
#682390000000
1!
1*
b101 6
19
1>
1C
b101 G
#682400000000
0!
0*
09
0>
0C
#682410000000
1!
1*
b110 6
19
1>
1C
b110 G
#682420000000
0!
0*
09
0>
0C
#682430000000
1!
1*
b111 6
19
1>
1C
b111 G
#682440000000
0!
0*
09
0>
0C
#682450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#682460000000
0!
0*
09
0>
0C
#682470000000
1!
1*
b1 6
19
1>
1C
b1 G
#682480000000
0!
0*
09
0>
0C
#682490000000
1!
1*
b10 6
19
1>
1C
b10 G
#682500000000
0!
0*
09
0>
0C
#682510000000
1!
1*
b11 6
19
1>
1C
b11 G
#682520000000
0!
0*
09
0>
0C
#682530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#682540000000
0!
0*
09
0>
0C
#682550000000
1!
1*
b101 6
19
1>
1C
b101 G
#682560000000
0!
0*
09
0>
0C
#682570000000
1!
1*
b110 6
19
1>
1C
b110 G
#682580000000
0!
0*
09
0>
0C
#682590000000
1!
1*
b111 6
19
1>
1C
b111 G
#682600000000
0!
0*
09
0>
0C
#682610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#682620000000
0!
0*
09
0>
0C
#682630000000
1!
1*
b1 6
19
1>
1C
b1 G
#682640000000
0!
0*
09
0>
0C
#682650000000
1!
1*
b10 6
19
1>
1C
b10 G
#682660000000
0!
0*
09
0>
0C
#682670000000
1!
1*
b11 6
19
1>
1C
b11 G
#682680000000
0!
0*
09
0>
0C
#682690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#682700000000
0!
0*
09
0>
0C
#682710000000
1!
1*
b101 6
19
1>
1C
b101 G
#682720000000
0!
0*
09
0>
0C
#682730000000
1!
1*
b110 6
19
1>
1C
b110 G
#682740000000
0!
0*
09
0>
0C
#682750000000
1!
1*
b111 6
19
1>
1C
b111 G
#682760000000
0!
1"
0*
1+
09
1:
0>
0C
#682770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#682780000000
0!
0*
09
0>
0C
#682790000000
1!
1*
b1 6
19
1>
1C
b1 G
#682800000000
0!
0*
09
0>
0C
#682810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#682820000000
0!
0*
09
0>
0C
#682830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#682840000000
0!
0*
09
0>
0C
#682850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#682860000000
0!
0*
09
0>
0C
#682870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#682880000000
0!
0#
0*
0,
09
0>
0?
0C
#682890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#682900000000
0!
0*
09
0>
0C
#682910000000
1!
1*
19
1>
1C
#682920000000
0!
0*
09
0>
0C
#682930000000
1!
1*
19
1>
1C
#682940000000
0!
0*
09
0>
0C
#682950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#682960000000
0!
0*
09
0>
0C
#682970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#682980000000
0!
0*
09
0>
0C
#682990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#683000000000
0!
0*
09
0>
0C
#683010000000
1!
1*
b10 6
19
1>
1C
b10 G
#683020000000
0!
0*
09
0>
0C
#683030000000
1!
1*
b11 6
19
1>
1C
b11 G
#683040000000
0!
0*
09
0>
0C
#683050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#683060000000
0!
0*
09
0>
0C
#683070000000
1!
1*
b101 6
19
1>
1C
b101 G
#683080000000
0!
0*
09
0>
0C
#683090000000
1!
1*
b110 6
19
1>
1C
b110 G
#683100000000
0!
0*
09
0>
0C
#683110000000
1!
1*
b111 6
19
1>
1C
b111 G
#683120000000
0!
0*
09
0>
0C
#683130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#683140000000
0!
0*
09
0>
0C
#683150000000
1!
1*
b1 6
19
1>
1C
b1 G
#683160000000
0!
0*
09
0>
0C
#683170000000
1!
1*
b10 6
19
1>
1C
b10 G
#683180000000
0!
0*
09
0>
0C
#683190000000
1!
1*
b11 6
19
1>
1C
b11 G
#683200000000
0!
0*
09
0>
0C
#683210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#683220000000
0!
0*
09
0>
0C
#683230000000
1!
1*
b101 6
19
1>
1C
b101 G
#683240000000
0!
0*
09
0>
0C
#683250000000
1!
1*
b110 6
19
1>
1C
b110 G
#683260000000
0!
0*
09
0>
0C
#683270000000
1!
1*
b111 6
19
1>
1C
b111 G
#683280000000
0!
0*
09
0>
0C
#683290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#683300000000
0!
0*
09
0>
0C
#683310000000
1!
1*
b1 6
19
1>
1C
b1 G
#683320000000
0!
0*
09
0>
0C
#683330000000
1!
1*
b10 6
19
1>
1C
b10 G
#683340000000
0!
0*
09
0>
0C
#683350000000
1!
1*
b11 6
19
1>
1C
b11 G
#683360000000
0!
0*
09
0>
0C
#683370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#683380000000
0!
0*
09
0>
0C
#683390000000
1!
1*
b101 6
19
1>
1C
b101 G
#683400000000
0!
0*
09
0>
0C
#683410000000
1!
1*
b110 6
19
1>
1C
b110 G
#683420000000
0!
0*
09
0>
0C
#683430000000
1!
1*
b111 6
19
1>
1C
b111 G
#683440000000
0!
1"
0*
1+
09
1:
0>
0C
#683450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#683460000000
0!
0*
09
0>
0C
#683470000000
1!
1*
b1 6
19
1>
1C
b1 G
#683480000000
0!
0*
09
0>
0C
#683490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#683500000000
0!
0*
09
0>
0C
#683510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#683520000000
0!
0*
09
0>
0C
#683530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#683540000000
0!
0*
09
0>
0C
#683550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#683560000000
0!
0#
0*
0,
09
0>
0?
0C
#683570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#683580000000
0!
0*
09
0>
0C
#683590000000
1!
1*
19
1>
1C
#683600000000
0!
0*
09
0>
0C
#683610000000
1!
1*
19
1>
1C
#683620000000
0!
0*
09
0>
0C
#683630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#683640000000
0!
0*
09
0>
0C
#683650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#683660000000
0!
0*
09
0>
0C
#683670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#683680000000
0!
0*
09
0>
0C
#683690000000
1!
1*
b10 6
19
1>
1C
b10 G
#683700000000
0!
0*
09
0>
0C
#683710000000
1!
1*
b11 6
19
1>
1C
b11 G
#683720000000
0!
0*
09
0>
0C
#683730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#683740000000
0!
0*
09
0>
0C
#683750000000
1!
1*
b101 6
19
1>
1C
b101 G
#683760000000
0!
0*
09
0>
0C
#683770000000
1!
1*
b110 6
19
1>
1C
b110 G
#683780000000
0!
0*
09
0>
0C
#683790000000
1!
1*
b111 6
19
1>
1C
b111 G
#683800000000
0!
0*
09
0>
0C
#683810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#683820000000
0!
0*
09
0>
0C
#683830000000
1!
1*
b1 6
19
1>
1C
b1 G
#683840000000
0!
0*
09
0>
0C
#683850000000
1!
1*
b10 6
19
1>
1C
b10 G
#683860000000
0!
0*
09
0>
0C
#683870000000
1!
1*
b11 6
19
1>
1C
b11 G
#683880000000
0!
0*
09
0>
0C
#683890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#683900000000
0!
0*
09
0>
0C
#683910000000
1!
1*
b101 6
19
1>
1C
b101 G
#683920000000
0!
0*
09
0>
0C
#683930000000
1!
1*
b110 6
19
1>
1C
b110 G
#683940000000
0!
0*
09
0>
0C
#683950000000
1!
1*
b111 6
19
1>
1C
b111 G
#683960000000
0!
0*
09
0>
0C
#683970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#683980000000
0!
0*
09
0>
0C
#683990000000
1!
1*
b1 6
19
1>
1C
b1 G
#684000000000
0!
0*
09
0>
0C
#684010000000
1!
1*
b10 6
19
1>
1C
b10 G
#684020000000
0!
0*
09
0>
0C
#684030000000
1!
1*
b11 6
19
1>
1C
b11 G
#684040000000
0!
0*
09
0>
0C
#684050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#684060000000
0!
0*
09
0>
0C
#684070000000
1!
1*
b101 6
19
1>
1C
b101 G
#684080000000
0!
0*
09
0>
0C
#684090000000
1!
1*
b110 6
19
1>
1C
b110 G
#684100000000
0!
0*
09
0>
0C
#684110000000
1!
1*
b111 6
19
1>
1C
b111 G
#684120000000
0!
1"
0*
1+
09
1:
0>
0C
#684130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#684140000000
0!
0*
09
0>
0C
#684150000000
1!
1*
b1 6
19
1>
1C
b1 G
#684160000000
0!
0*
09
0>
0C
#684170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#684180000000
0!
0*
09
0>
0C
#684190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#684200000000
0!
0*
09
0>
0C
#684210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#684220000000
0!
0*
09
0>
0C
#684230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#684240000000
0!
0#
0*
0,
09
0>
0?
0C
#684250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#684260000000
0!
0*
09
0>
0C
#684270000000
1!
1*
19
1>
1C
#684280000000
0!
0*
09
0>
0C
#684290000000
1!
1*
19
1>
1C
#684300000000
0!
0*
09
0>
0C
#684310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#684320000000
0!
0*
09
0>
0C
#684330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#684340000000
0!
0*
09
0>
0C
#684350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#684360000000
0!
0*
09
0>
0C
#684370000000
1!
1*
b10 6
19
1>
1C
b10 G
#684380000000
0!
0*
09
0>
0C
#684390000000
1!
1*
b11 6
19
1>
1C
b11 G
#684400000000
0!
0*
09
0>
0C
#684410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#684420000000
0!
0*
09
0>
0C
#684430000000
1!
1*
b101 6
19
1>
1C
b101 G
#684440000000
0!
0*
09
0>
0C
#684450000000
1!
1*
b110 6
19
1>
1C
b110 G
#684460000000
0!
0*
09
0>
0C
#684470000000
1!
1*
b111 6
19
1>
1C
b111 G
#684480000000
0!
0*
09
0>
0C
#684490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#684500000000
0!
0*
09
0>
0C
#684510000000
1!
1*
b1 6
19
1>
1C
b1 G
#684520000000
0!
0*
09
0>
0C
#684530000000
1!
1*
b10 6
19
1>
1C
b10 G
#684540000000
0!
0*
09
0>
0C
#684550000000
1!
1*
b11 6
19
1>
1C
b11 G
#684560000000
0!
0*
09
0>
0C
#684570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#684580000000
0!
0*
09
0>
0C
#684590000000
1!
1*
b101 6
19
1>
1C
b101 G
#684600000000
0!
0*
09
0>
0C
#684610000000
1!
1*
b110 6
19
1>
1C
b110 G
#684620000000
0!
0*
09
0>
0C
#684630000000
1!
1*
b111 6
19
1>
1C
b111 G
#684640000000
0!
0*
09
0>
0C
#684650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#684660000000
0!
0*
09
0>
0C
#684670000000
1!
1*
b1 6
19
1>
1C
b1 G
#684680000000
0!
0*
09
0>
0C
#684690000000
1!
1*
b10 6
19
1>
1C
b10 G
#684700000000
0!
0*
09
0>
0C
#684710000000
1!
1*
b11 6
19
1>
1C
b11 G
#684720000000
0!
0*
09
0>
0C
#684730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#684740000000
0!
0*
09
0>
0C
#684750000000
1!
1*
b101 6
19
1>
1C
b101 G
#684760000000
0!
0*
09
0>
0C
#684770000000
1!
1*
b110 6
19
1>
1C
b110 G
#684780000000
0!
0*
09
0>
0C
#684790000000
1!
1*
b111 6
19
1>
1C
b111 G
#684800000000
0!
1"
0*
1+
09
1:
0>
0C
#684810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#684820000000
0!
0*
09
0>
0C
#684830000000
1!
1*
b1 6
19
1>
1C
b1 G
#684840000000
0!
0*
09
0>
0C
#684850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#684860000000
0!
0*
09
0>
0C
#684870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#684880000000
0!
0*
09
0>
0C
#684890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#684900000000
0!
0*
09
0>
0C
#684910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#684920000000
0!
0#
0*
0,
09
0>
0?
0C
#684930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#684940000000
0!
0*
09
0>
0C
#684950000000
1!
1*
19
1>
1C
#684960000000
0!
0*
09
0>
0C
#684970000000
1!
1*
19
1>
1C
#684980000000
0!
0*
09
0>
0C
#684990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#685000000000
0!
0*
09
0>
0C
#685010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#685020000000
0!
0*
09
0>
0C
#685030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#685040000000
0!
0*
09
0>
0C
#685050000000
1!
1*
b10 6
19
1>
1C
b10 G
#685060000000
0!
0*
09
0>
0C
#685070000000
1!
1*
b11 6
19
1>
1C
b11 G
#685080000000
0!
0*
09
0>
0C
#685090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#685100000000
0!
0*
09
0>
0C
#685110000000
1!
1*
b101 6
19
1>
1C
b101 G
#685120000000
0!
0*
09
0>
0C
#685130000000
1!
1*
b110 6
19
1>
1C
b110 G
#685140000000
0!
0*
09
0>
0C
#685150000000
1!
1*
b111 6
19
1>
1C
b111 G
#685160000000
0!
0*
09
0>
0C
#685170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#685180000000
0!
0*
09
0>
0C
#685190000000
1!
1*
b1 6
19
1>
1C
b1 G
#685200000000
0!
0*
09
0>
0C
#685210000000
1!
1*
b10 6
19
1>
1C
b10 G
#685220000000
0!
0*
09
0>
0C
#685230000000
1!
1*
b11 6
19
1>
1C
b11 G
#685240000000
0!
0*
09
0>
0C
#685250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#685260000000
0!
0*
09
0>
0C
#685270000000
1!
1*
b101 6
19
1>
1C
b101 G
#685280000000
0!
0*
09
0>
0C
#685290000000
1!
1*
b110 6
19
1>
1C
b110 G
#685300000000
0!
0*
09
0>
0C
#685310000000
1!
1*
b111 6
19
1>
1C
b111 G
#685320000000
0!
0*
09
0>
0C
#685330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#685340000000
0!
0*
09
0>
0C
#685350000000
1!
1*
b1 6
19
1>
1C
b1 G
#685360000000
0!
0*
09
0>
0C
#685370000000
1!
1*
b10 6
19
1>
1C
b10 G
#685380000000
0!
0*
09
0>
0C
#685390000000
1!
1*
b11 6
19
1>
1C
b11 G
#685400000000
0!
0*
09
0>
0C
#685410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#685420000000
0!
0*
09
0>
0C
#685430000000
1!
1*
b101 6
19
1>
1C
b101 G
#685440000000
0!
0*
09
0>
0C
#685450000000
1!
1*
b110 6
19
1>
1C
b110 G
#685460000000
0!
0*
09
0>
0C
#685470000000
1!
1*
b111 6
19
1>
1C
b111 G
#685480000000
0!
1"
0*
1+
09
1:
0>
0C
#685490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#685500000000
0!
0*
09
0>
0C
#685510000000
1!
1*
b1 6
19
1>
1C
b1 G
#685520000000
0!
0*
09
0>
0C
#685530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#685540000000
0!
0*
09
0>
0C
#685550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#685560000000
0!
0*
09
0>
0C
#685570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#685580000000
0!
0*
09
0>
0C
#685590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#685600000000
0!
0#
0*
0,
09
0>
0?
0C
#685610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#685620000000
0!
0*
09
0>
0C
#685630000000
1!
1*
19
1>
1C
#685640000000
0!
0*
09
0>
0C
#685650000000
1!
1*
19
1>
1C
#685660000000
0!
0*
09
0>
0C
#685670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#685680000000
0!
0*
09
0>
0C
#685690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#685700000000
0!
0*
09
0>
0C
#685710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#685720000000
0!
0*
09
0>
0C
#685730000000
1!
1*
b10 6
19
1>
1C
b10 G
#685740000000
0!
0*
09
0>
0C
#685750000000
1!
1*
b11 6
19
1>
1C
b11 G
#685760000000
0!
0*
09
0>
0C
#685770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#685780000000
0!
0*
09
0>
0C
#685790000000
1!
1*
b101 6
19
1>
1C
b101 G
#685800000000
0!
0*
09
0>
0C
#685810000000
1!
1*
b110 6
19
1>
1C
b110 G
#685820000000
0!
0*
09
0>
0C
#685830000000
1!
1*
b111 6
19
1>
1C
b111 G
#685840000000
0!
0*
09
0>
0C
#685850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#685860000000
0!
0*
09
0>
0C
#685870000000
1!
1*
b1 6
19
1>
1C
b1 G
#685880000000
0!
0*
09
0>
0C
#685890000000
1!
1*
b10 6
19
1>
1C
b10 G
#685900000000
0!
0*
09
0>
0C
#685910000000
1!
1*
b11 6
19
1>
1C
b11 G
#685920000000
0!
0*
09
0>
0C
#685930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#685940000000
0!
0*
09
0>
0C
#685950000000
1!
1*
b101 6
19
1>
1C
b101 G
#685960000000
0!
0*
09
0>
0C
#685970000000
1!
1*
b110 6
19
1>
1C
b110 G
#685980000000
0!
0*
09
0>
0C
#685990000000
1!
1*
b111 6
19
1>
1C
b111 G
#686000000000
0!
0*
09
0>
0C
#686010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#686020000000
0!
0*
09
0>
0C
#686030000000
1!
1*
b1 6
19
1>
1C
b1 G
#686040000000
0!
0*
09
0>
0C
#686050000000
1!
1*
b10 6
19
1>
1C
b10 G
#686060000000
0!
0*
09
0>
0C
#686070000000
1!
1*
b11 6
19
1>
1C
b11 G
#686080000000
0!
0*
09
0>
0C
#686090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#686100000000
0!
0*
09
0>
0C
#686110000000
1!
1*
b101 6
19
1>
1C
b101 G
#686120000000
0!
0*
09
0>
0C
#686130000000
1!
1*
b110 6
19
1>
1C
b110 G
#686140000000
0!
0*
09
0>
0C
#686150000000
1!
1*
b111 6
19
1>
1C
b111 G
#686160000000
0!
1"
0*
1+
09
1:
0>
0C
#686170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#686180000000
0!
0*
09
0>
0C
#686190000000
1!
1*
b1 6
19
1>
1C
b1 G
#686200000000
0!
0*
09
0>
0C
#686210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#686220000000
0!
0*
09
0>
0C
#686230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#686240000000
0!
0*
09
0>
0C
#686250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#686260000000
0!
0*
09
0>
0C
#686270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#686280000000
0!
0#
0*
0,
09
0>
0?
0C
#686290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#686300000000
0!
0*
09
0>
0C
#686310000000
1!
1*
19
1>
1C
#686320000000
0!
0*
09
0>
0C
#686330000000
1!
1*
19
1>
1C
#686340000000
0!
0*
09
0>
0C
#686350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#686360000000
0!
0*
09
0>
0C
#686370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#686380000000
0!
0*
09
0>
0C
#686390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#686400000000
0!
0*
09
0>
0C
#686410000000
1!
1*
b10 6
19
1>
1C
b10 G
#686420000000
0!
0*
09
0>
0C
#686430000000
1!
1*
b11 6
19
1>
1C
b11 G
#686440000000
0!
0*
09
0>
0C
#686450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#686460000000
0!
0*
09
0>
0C
#686470000000
1!
1*
b101 6
19
1>
1C
b101 G
#686480000000
0!
0*
09
0>
0C
#686490000000
1!
1*
b110 6
19
1>
1C
b110 G
#686500000000
0!
0*
09
0>
0C
#686510000000
1!
1*
b111 6
19
1>
1C
b111 G
#686520000000
0!
0*
09
0>
0C
#686530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#686540000000
0!
0*
09
0>
0C
#686550000000
1!
1*
b1 6
19
1>
1C
b1 G
#686560000000
0!
0*
09
0>
0C
#686570000000
1!
1*
b10 6
19
1>
1C
b10 G
#686580000000
0!
0*
09
0>
0C
#686590000000
1!
1*
b11 6
19
1>
1C
b11 G
#686600000000
0!
0*
09
0>
0C
#686610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#686620000000
0!
0*
09
0>
0C
#686630000000
1!
1*
b101 6
19
1>
1C
b101 G
#686640000000
0!
0*
09
0>
0C
#686650000000
1!
1*
b110 6
19
1>
1C
b110 G
#686660000000
0!
0*
09
0>
0C
#686670000000
1!
1*
b111 6
19
1>
1C
b111 G
#686680000000
0!
0*
09
0>
0C
#686690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#686700000000
0!
0*
09
0>
0C
#686710000000
1!
1*
b1 6
19
1>
1C
b1 G
#686720000000
0!
0*
09
0>
0C
#686730000000
1!
1*
b10 6
19
1>
1C
b10 G
#686740000000
0!
0*
09
0>
0C
#686750000000
1!
1*
b11 6
19
1>
1C
b11 G
#686760000000
0!
0*
09
0>
0C
#686770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#686780000000
0!
0*
09
0>
0C
#686790000000
1!
1*
b101 6
19
1>
1C
b101 G
#686800000000
0!
0*
09
0>
0C
#686810000000
1!
1*
b110 6
19
1>
1C
b110 G
#686820000000
0!
0*
09
0>
0C
#686830000000
1!
1*
b111 6
19
1>
1C
b111 G
#686840000000
0!
1"
0*
1+
09
1:
0>
0C
#686850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#686860000000
0!
0*
09
0>
0C
#686870000000
1!
1*
b1 6
19
1>
1C
b1 G
#686880000000
0!
0*
09
0>
0C
#686890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#686900000000
0!
0*
09
0>
0C
#686910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#686920000000
0!
0*
09
0>
0C
#686930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#686940000000
0!
0*
09
0>
0C
#686950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#686960000000
0!
0#
0*
0,
09
0>
0?
0C
#686970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#686980000000
0!
0*
09
0>
0C
#686990000000
1!
1*
19
1>
1C
#687000000000
0!
0*
09
0>
0C
#687010000000
1!
1*
19
1>
1C
#687020000000
0!
0*
09
0>
0C
#687030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#687040000000
0!
0*
09
0>
0C
#687050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#687060000000
0!
0*
09
0>
0C
#687070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#687080000000
0!
0*
09
0>
0C
#687090000000
1!
1*
b10 6
19
1>
1C
b10 G
#687100000000
0!
0*
09
0>
0C
#687110000000
1!
1*
b11 6
19
1>
1C
b11 G
#687120000000
0!
0*
09
0>
0C
#687130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#687140000000
0!
0*
09
0>
0C
#687150000000
1!
1*
b101 6
19
1>
1C
b101 G
#687160000000
0!
0*
09
0>
0C
#687170000000
1!
1*
b110 6
19
1>
1C
b110 G
#687180000000
0!
0*
09
0>
0C
#687190000000
1!
1*
b111 6
19
1>
1C
b111 G
#687200000000
0!
0*
09
0>
0C
#687210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#687220000000
0!
0*
09
0>
0C
#687230000000
1!
1*
b1 6
19
1>
1C
b1 G
#687240000000
0!
0*
09
0>
0C
#687250000000
1!
1*
b10 6
19
1>
1C
b10 G
#687260000000
0!
0*
09
0>
0C
#687270000000
1!
1*
b11 6
19
1>
1C
b11 G
#687280000000
0!
0*
09
0>
0C
#687290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#687300000000
0!
0*
09
0>
0C
#687310000000
1!
1*
b101 6
19
1>
1C
b101 G
#687320000000
0!
0*
09
0>
0C
#687330000000
1!
1*
b110 6
19
1>
1C
b110 G
#687340000000
0!
0*
09
0>
0C
#687350000000
1!
1*
b111 6
19
1>
1C
b111 G
#687360000000
0!
0*
09
0>
0C
#687370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#687380000000
0!
0*
09
0>
0C
#687390000000
1!
1*
b1 6
19
1>
1C
b1 G
#687400000000
0!
0*
09
0>
0C
#687410000000
1!
1*
b10 6
19
1>
1C
b10 G
#687420000000
0!
0*
09
0>
0C
#687430000000
1!
1*
b11 6
19
1>
1C
b11 G
#687440000000
0!
0*
09
0>
0C
#687450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#687460000000
0!
0*
09
0>
0C
#687470000000
1!
1*
b101 6
19
1>
1C
b101 G
#687480000000
0!
0*
09
0>
0C
#687490000000
1!
1*
b110 6
19
1>
1C
b110 G
#687500000000
0!
0*
09
0>
0C
#687510000000
1!
1*
b111 6
19
1>
1C
b111 G
#687520000000
0!
1"
0*
1+
09
1:
0>
0C
#687530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#687540000000
0!
0*
09
0>
0C
#687550000000
1!
1*
b1 6
19
1>
1C
b1 G
#687560000000
0!
0*
09
0>
0C
#687570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#687580000000
0!
0*
09
0>
0C
#687590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#687600000000
0!
0*
09
0>
0C
#687610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#687620000000
0!
0*
09
0>
0C
#687630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#687640000000
0!
0#
0*
0,
09
0>
0?
0C
#687650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#687660000000
0!
0*
09
0>
0C
#687670000000
1!
1*
19
1>
1C
#687680000000
0!
0*
09
0>
0C
#687690000000
1!
1*
19
1>
1C
#687700000000
0!
0*
09
0>
0C
#687710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#687720000000
0!
0*
09
0>
0C
#687730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#687740000000
0!
0*
09
0>
0C
#687750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#687760000000
0!
0*
09
0>
0C
#687770000000
1!
1*
b10 6
19
1>
1C
b10 G
#687780000000
0!
0*
09
0>
0C
#687790000000
1!
1*
b11 6
19
1>
1C
b11 G
#687800000000
0!
0*
09
0>
0C
#687810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#687820000000
0!
0*
09
0>
0C
#687830000000
1!
1*
b101 6
19
1>
1C
b101 G
#687840000000
0!
0*
09
0>
0C
#687850000000
1!
1*
b110 6
19
1>
1C
b110 G
#687860000000
0!
0*
09
0>
0C
#687870000000
1!
1*
b111 6
19
1>
1C
b111 G
#687880000000
0!
0*
09
0>
0C
#687890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#687900000000
0!
0*
09
0>
0C
#687910000000
1!
1*
b1 6
19
1>
1C
b1 G
#687920000000
0!
0*
09
0>
0C
#687930000000
1!
1*
b10 6
19
1>
1C
b10 G
#687940000000
0!
0*
09
0>
0C
#687950000000
1!
1*
b11 6
19
1>
1C
b11 G
#687960000000
0!
0*
09
0>
0C
#687970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#687980000000
0!
0*
09
0>
0C
#687990000000
1!
1*
b101 6
19
1>
1C
b101 G
#688000000000
0!
0*
09
0>
0C
#688010000000
1!
1*
b110 6
19
1>
1C
b110 G
#688020000000
0!
0*
09
0>
0C
#688030000000
1!
1*
b111 6
19
1>
1C
b111 G
#688040000000
0!
0*
09
0>
0C
#688050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#688060000000
0!
0*
09
0>
0C
#688070000000
1!
1*
b1 6
19
1>
1C
b1 G
#688080000000
0!
0*
09
0>
0C
#688090000000
1!
1*
b10 6
19
1>
1C
b10 G
#688100000000
0!
0*
09
0>
0C
#688110000000
1!
1*
b11 6
19
1>
1C
b11 G
#688120000000
0!
0*
09
0>
0C
#688130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#688140000000
0!
0*
09
0>
0C
#688150000000
1!
1*
b101 6
19
1>
1C
b101 G
#688160000000
0!
0*
09
0>
0C
#688170000000
1!
1*
b110 6
19
1>
1C
b110 G
#688180000000
0!
0*
09
0>
0C
#688190000000
1!
1*
b111 6
19
1>
1C
b111 G
#688200000000
0!
1"
0*
1+
09
1:
0>
0C
#688210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#688220000000
0!
0*
09
0>
0C
#688230000000
1!
1*
b1 6
19
1>
1C
b1 G
#688240000000
0!
0*
09
0>
0C
#688250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#688260000000
0!
0*
09
0>
0C
#688270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#688280000000
0!
0*
09
0>
0C
#688290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#688300000000
0!
0*
09
0>
0C
#688310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#688320000000
0!
0#
0*
0,
09
0>
0?
0C
#688330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#688340000000
0!
0*
09
0>
0C
#688350000000
1!
1*
19
1>
1C
#688360000000
0!
0*
09
0>
0C
#688370000000
1!
1*
19
1>
1C
#688380000000
0!
0*
09
0>
0C
#688390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#688400000000
0!
0*
09
0>
0C
#688410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#688420000000
0!
0*
09
0>
0C
#688430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#688440000000
0!
0*
09
0>
0C
#688450000000
1!
1*
b10 6
19
1>
1C
b10 G
#688460000000
0!
0*
09
0>
0C
#688470000000
1!
1*
b11 6
19
1>
1C
b11 G
#688480000000
0!
0*
09
0>
0C
#688490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#688500000000
0!
0*
09
0>
0C
#688510000000
1!
1*
b101 6
19
1>
1C
b101 G
#688520000000
0!
0*
09
0>
0C
#688530000000
1!
1*
b110 6
19
1>
1C
b110 G
#688540000000
0!
0*
09
0>
0C
#688550000000
1!
1*
b111 6
19
1>
1C
b111 G
#688560000000
0!
0*
09
0>
0C
#688570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#688580000000
0!
0*
09
0>
0C
#688590000000
1!
1*
b1 6
19
1>
1C
b1 G
#688600000000
0!
0*
09
0>
0C
#688610000000
1!
1*
b10 6
19
1>
1C
b10 G
#688620000000
0!
0*
09
0>
0C
#688630000000
1!
1*
b11 6
19
1>
1C
b11 G
#688640000000
0!
0*
09
0>
0C
#688650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#688660000000
0!
0*
09
0>
0C
#688670000000
1!
1*
b101 6
19
1>
1C
b101 G
#688680000000
0!
0*
09
0>
0C
#688690000000
1!
1*
b110 6
19
1>
1C
b110 G
#688700000000
0!
0*
09
0>
0C
#688710000000
1!
1*
b111 6
19
1>
1C
b111 G
#688720000000
0!
0*
09
0>
0C
#688730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#688740000000
0!
0*
09
0>
0C
#688750000000
1!
1*
b1 6
19
1>
1C
b1 G
#688760000000
0!
0*
09
0>
0C
#688770000000
1!
1*
b10 6
19
1>
1C
b10 G
#688780000000
0!
0*
09
0>
0C
#688790000000
1!
1*
b11 6
19
1>
1C
b11 G
#688800000000
0!
0*
09
0>
0C
#688810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#688820000000
0!
0*
09
0>
0C
#688830000000
1!
1*
b101 6
19
1>
1C
b101 G
#688840000000
0!
0*
09
0>
0C
#688850000000
1!
1*
b110 6
19
1>
1C
b110 G
#688860000000
0!
0*
09
0>
0C
#688870000000
1!
1*
b111 6
19
1>
1C
b111 G
#688880000000
0!
1"
0*
1+
09
1:
0>
0C
#688890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#688900000000
0!
0*
09
0>
0C
#688910000000
1!
1*
b1 6
19
1>
1C
b1 G
#688920000000
0!
0*
09
0>
0C
#688930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#688940000000
0!
0*
09
0>
0C
#688950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#688960000000
0!
0*
09
0>
0C
#688970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#688980000000
0!
0*
09
0>
0C
#688990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#689000000000
0!
0#
0*
0,
09
0>
0?
0C
#689010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#689020000000
0!
0*
09
0>
0C
#689030000000
1!
1*
19
1>
1C
#689040000000
0!
0*
09
0>
0C
#689050000000
1!
1*
19
1>
1C
#689060000000
0!
0*
09
0>
0C
#689070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#689080000000
0!
0*
09
0>
0C
#689090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#689100000000
0!
0*
09
0>
0C
#689110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#689120000000
0!
0*
09
0>
0C
#689130000000
1!
1*
b10 6
19
1>
1C
b10 G
#689140000000
0!
0*
09
0>
0C
#689150000000
1!
1*
b11 6
19
1>
1C
b11 G
#689160000000
0!
0*
09
0>
0C
#689170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#689180000000
0!
0*
09
0>
0C
#689190000000
1!
1*
b101 6
19
1>
1C
b101 G
#689200000000
0!
0*
09
0>
0C
#689210000000
1!
1*
b110 6
19
1>
1C
b110 G
#689220000000
0!
0*
09
0>
0C
#689230000000
1!
1*
b111 6
19
1>
1C
b111 G
#689240000000
0!
0*
09
0>
0C
#689250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#689260000000
0!
0*
09
0>
0C
#689270000000
1!
1*
b1 6
19
1>
1C
b1 G
#689280000000
0!
0*
09
0>
0C
#689290000000
1!
1*
b10 6
19
1>
1C
b10 G
#689300000000
0!
0*
09
0>
0C
#689310000000
1!
1*
b11 6
19
1>
1C
b11 G
#689320000000
0!
0*
09
0>
0C
#689330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#689340000000
0!
0*
09
0>
0C
#689350000000
1!
1*
b101 6
19
1>
1C
b101 G
#689360000000
0!
0*
09
0>
0C
#689370000000
1!
1*
b110 6
19
1>
1C
b110 G
#689380000000
0!
0*
09
0>
0C
#689390000000
1!
1*
b111 6
19
1>
1C
b111 G
#689400000000
0!
0*
09
0>
0C
#689410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#689420000000
0!
0*
09
0>
0C
#689430000000
1!
1*
b1 6
19
1>
1C
b1 G
#689440000000
0!
0*
09
0>
0C
#689450000000
1!
1*
b10 6
19
1>
1C
b10 G
#689460000000
0!
0*
09
0>
0C
#689470000000
1!
1*
b11 6
19
1>
1C
b11 G
#689480000000
0!
0*
09
0>
0C
#689490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#689500000000
0!
0*
09
0>
0C
#689510000000
1!
1*
b101 6
19
1>
1C
b101 G
#689520000000
0!
0*
09
0>
0C
#689530000000
1!
1*
b110 6
19
1>
1C
b110 G
#689540000000
0!
0*
09
0>
0C
#689550000000
1!
1*
b111 6
19
1>
1C
b111 G
#689560000000
0!
1"
0*
1+
09
1:
0>
0C
#689570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#689580000000
0!
0*
09
0>
0C
#689590000000
1!
1*
b1 6
19
1>
1C
b1 G
#689600000000
0!
0*
09
0>
0C
#689610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#689620000000
0!
0*
09
0>
0C
#689630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#689640000000
0!
0*
09
0>
0C
#689650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#689660000000
0!
0*
09
0>
0C
#689670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#689680000000
0!
0#
0*
0,
09
0>
0?
0C
#689690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#689700000000
0!
0*
09
0>
0C
#689710000000
1!
1*
19
1>
1C
#689720000000
0!
0*
09
0>
0C
#689730000000
1!
1*
19
1>
1C
#689740000000
0!
0*
09
0>
0C
#689750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#689760000000
0!
0*
09
0>
0C
#689770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#689780000000
0!
0*
09
0>
0C
#689790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#689800000000
0!
0*
09
0>
0C
#689810000000
1!
1*
b10 6
19
1>
1C
b10 G
#689820000000
0!
0*
09
0>
0C
#689830000000
1!
1*
b11 6
19
1>
1C
b11 G
#689840000000
0!
0*
09
0>
0C
#689850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#689860000000
0!
0*
09
0>
0C
#689870000000
1!
1*
b101 6
19
1>
1C
b101 G
#689880000000
0!
0*
09
0>
0C
#689890000000
1!
1*
b110 6
19
1>
1C
b110 G
#689900000000
0!
0*
09
0>
0C
#689910000000
1!
1*
b111 6
19
1>
1C
b111 G
#689920000000
0!
0*
09
0>
0C
#689930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#689940000000
0!
0*
09
0>
0C
#689950000000
1!
1*
b1 6
19
1>
1C
b1 G
#689960000000
0!
0*
09
0>
0C
#689970000000
1!
1*
b10 6
19
1>
1C
b10 G
#689980000000
0!
0*
09
0>
0C
#689990000000
1!
1*
b11 6
19
1>
1C
b11 G
#690000000000
0!
0*
09
0>
0C
#690010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#690020000000
0!
0*
09
0>
0C
#690030000000
1!
1*
b101 6
19
1>
1C
b101 G
#690040000000
0!
0*
09
0>
0C
#690050000000
1!
1*
b110 6
19
1>
1C
b110 G
#690060000000
0!
0*
09
0>
0C
#690070000000
1!
1*
b111 6
19
1>
1C
b111 G
#690080000000
0!
0*
09
0>
0C
#690090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#690100000000
0!
0*
09
0>
0C
#690110000000
1!
1*
b1 6
19
1>
1C
b1 G
#690120000000
0!
0*
09
0>
0C
#690130000000
1!
1*
b10 6
19
1>
1C
b10 G
#690140000000
0!
0*
09
0>
0C
#690150000000
1!
1*
b11 6
19
1>
1C
b11 G
#690160000000
0!
0*
09
0>
0C
#690170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#690180000000
0!
0*
09
0>
0C
#690190000000
1!
1*
b101 6
19
1>
1C
b101 G
#690200000000
0!
0*
09
0>
0C
#690210000000
1!
1*
b110 6
19
1>
1C
b110 G
#690220000000
0!
0*
09
0>
0C
#690230000000
1!
1*
b111 6
19
1>
1C
b111 G
#690240000000
0!
1"
0*
1+
09
1:
0>
0C
#690250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#690260000000
0!
0*
09
0>
0C
#690270000000
1!
1*
b1 6
19
1>
1C
b1 G
#690280000000
0!
0*
09
0>
0C
#690290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#690300000000
0!
0*
09
0>
0C
#690310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#690320000000
0!
0*
09
0>
0C
#690330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#690340000000
0!
0*
09
0>
0C
#690350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#690360000000
0!
0#
0*
0,
09
0>
0?
0C
#690370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#690380000000
0!
0*
09
0>
0C
#690390000000
1!
1*
19
1>
1C
#690400000000
0!
0*
09
0>
0C
#690410000000
1!
1*
19
1>
1C
#690420000000
0!
0*
09
0>
0C
#690430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#690440000000
0!
0*
09
0>
0C
#690450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#690460000000
0!
0*
09
0>
0C
#690470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#690480000000
0!
0*
09
0>
0C
#690490000000
1!
1*
b10 6
19
1>
1C
b10 G
#690500000000
0!
0*
09
0>
0C
#690510000000
1!
1*
b11 6
19
1>
1C
b11 G
#690520000000
0!
0*
09
0>
0C
#690530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#690540000000
0!
0*
09
0>
0C
#690550000000
1!
1*
b101 6
19
1>
1C
b101 G
#690560000000
0!
0*
09
0>
0C
#690570000000
1!
1*
b110 6
19
1>
1C
b110 G
#690580000000
0!
0*
09
0>
0C
#690590000000
1!
1*
b111 6
19
1>
1C
b111 G
#690600000000
0!
0*
09
0>
0C
#690610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#690620000000
0!
0*
09
0>
0C
#690630000000
1!
1*
b1 6
19
1>
1C
b1 G
#690640000000
0!
0*
09
0>
0C
#690650000000
1!
1*
b10 6
19
1>
1C
b10 G
#690660000000
0!
0*
09
0>
0C
#690670000000
1!
1*
b11 6
19
1>
1C
b11 G
#690680000000
0!
0*
09
0>
0C
#690690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#690700000000
0!
0*
09
0>
0C
#690710000000
1!
1*
b101 6
19
1>
1C
b101 G
#690720000000
0!
0*
09
0>
0C
#690730000000
1!
1*
b110 6
19
1>
1C
b110 G
#690740000000
0!
0*
09
0>
0C
#690750000000
1!
1*
b111 6
19
1>
1C
b111 G
#690760000000
0!
0*
09
0>
0C
#690770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#690780000000
0!
0*
09
0>
0C
#690790000000
1!
1*
b1 6
19
1>
1C
b1 G
#690800000000
0!
0*
09
0>
0C
#690810000000
1!
1*
b10 6
19
1>
1C
b10 G
#690820000000
0!
0*
09
0>
0C
#690830000000
1!
1*
b11 6
19
1>
1C
b11 G
#690840000000
0!
0*
09
0>
0C
#690850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#690860000000
0!
0*
09
0>
0C
#690870000000
1!
1*
b101 6
19
1>
1C
b101 G
#690880000000
0!
0*
09
0>
0C
#690890000000
1!
1*
b110 6
19
1>
1C
b110 G
#690900000000
0!
0*
09
0>
0C
#690910000000
1!
1*
b111 6
19
1>
1C
b111 G
#690920000000
0!
1"
0*
1+
09
1:
0>
0C
#690930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#690940000000
0!
0*
09
0>
0C
#690950000000
1!
1*
b1 6
19
1>
1C
b1 G
#690960000000
0!
0*
09
0>
0C
#690970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#690980000000
0!
0*
09
0>
0C
#690990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#691000000000
0!
0*
09
0>
0C
#691010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#691020000000
0!
0*
09
0>
0C
#691030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#691040000000
0!
0#
0*
0,
09
0>
0?
0C
#691050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#691060000000
0!
0*
09
0>
0C
#691070000000
1!
1*
19
1>
1C
#691080000000
0!
0*
09
0>
0C
#691090000000
1!
1*
19
1>
1C
#691100000000
0!
0*
09
0>
0C
#691110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#691120000000
0!
0*
09
0>
0C
#691130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#691140000000
0!
0*
09
0>
0C
#691150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#691160000000
0!
0*
09
0>
0C
#691170000000
1!
1*
b10 6
19
1>
1C
b10 G
#691180000000
0!
0*
09
0>
0C
#691190000000
1!
1*
b11 6
19
1>
1C
b11 G
#691200000000
0!
0*
09
0>
0C
#691210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#691220000000
0!
0*
09
0>
0C
#691230000000
1!
1*
b101 6
19
1>
1C
b101 G
#691240000000
0!
0*
09
0>
0C
#691250000000
1!
1*
b110 6
19
1>
1C
b110 G
#691260000000
0!
0*
09
0>
0C
#691270000000
1!
1*
b111 6
19
1>
1C
b111 G
#691280000000
0!
0*
09
0>
0C
#691290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#691300000000
0!
0*
09
0>
0C
#691310000000
1!
1*
b1 6
19
1>
1C
b1 G
#691320000000
0!
0*
09
0>
0C
#691330000000
1!
1*
b10 6
19
1>
1C
b10 G
#691340000000
0!
0*
09
0>
0C
#691350000000
1!
1*
b11 6
19
1>
1C
b11 G
#691360000000
0!
0*
09
0>
0C
#691370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#691380000000
0!
0*
09
0>
0C
#691390000000
1!
1*
b101 6
19
1>
1C
b101 G
#691400000000
0!
0*
09
0>
0C
#691410000000
1!
1*
b110 6
19
1>
1C
b110 G
#691420000000
0!
0*
09
0>
0C
#691430000000
1!
1*
b111 6
19
1>
1C
b111 G
#691440000000
0!
0*
09
0>
0C
#691450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#691460000000
0!
0*
09
0>
0C
#691470000000
1!
1*
b1 6
19
1>
1C
b1 G
#691480000000
0!
0*
09
0>
0C
#691490000000
1!
1*
b10 6
19
1>
1C
b10 G
#691500000000
0!
0*
09
0>
0C
#691510000000
1!
1*
b11 6
19
1>
1C
b11 G
#691520000000
0!
0*
09
0>
0C
#691530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#691540000000
0!
0*
09
0>
0C
#691550000000
1!
1*
b101 6
19
1>
1C
b101 G
#691560000000
0!
0*
09
0>
0C
#691570000000
1!
1*
b110 6
19
1>
1C
b110 G
#691580000000
0!
0*
09
0>
0C
#691590000000
1!
1*
b111 6
19
1>
1C
b111 G
#691600000000
0!
1"
0*
1+
09
1:
0>
0C
#691610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#691620000000
0!
0*
09
0>
0C
#691630000000
1!
1*
b1 6
19
1>
1C
b1 G
#691640000000
0!
0*
09
0>
0C
#691650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#691660000000
0!
0*
09
0>
0C
#691670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#691680000000
0!
0*
09
0>
0C
#691690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#691700000000
0!
0*
09
0>
0C
#691710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#691720000000
0!
0#
0*
0,
09
0>
0?
0C
#691730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#691740000000
0!
0*
09
0>
0C
#691750000000
1!
1*
19
1>
1C
#691760000000
0!
0*
09
0>
0C
#691770000000
1!
1*
19
1>
1C
#691780000000
0!
0*
09
0>
0C
#691790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#691800000000
0!
0*
09
0>
0C
#691810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#691820000000
0!
0*
09
0>
0C
#691830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#691840000000
0!
0*
09
0>
0C
#691850000000
1!
1*
b10 6
19
1>
1C
b10 G
#691860000000
0!
0*
09
0>
0C
#691870000000
1!
1*
b11 6
19
1>
1C
b11 G
#691880000000
0!
0*
09
0>
0C
#691890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#691900000000
0!
0*
09
0>
0C
#691910000000
1!
1*
b101 6
19
1>
1C
b101 G
#691920000000
0!
0*
09
0>
0C
#691930000000
1!
1*
b110 6
19
1>
1C
b110 G
#691940000000
0!
0*
09
0>
0C
#691950000000
1!
1*
b111 6
19
1>
1C
b111 G
#691960000000
0!
0*
09
0>
0C
#691970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#691980000000
0!
0*
09
0>
0C
#691990000000
1!
1*
b1 6
19
1>
1C
b1 G
#692000000000
0!
0*
09
0>
0C
#692010000000
1!
1*
b10 6
19
1>
1C
b10 G
#692020000000
0!
0*
09
0>
0C
#692030000000
1!
1*
b11 6
19
1>
1C
b11 G
#692040000000
0!
0*
09
0>
0C
#692050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#692060000000
0!
0*
09
0>
0C
#692070000000
1!
1*
b101 6
19
1>
1C
b101 G
#692080000000
0!
0*
09
0>
0C
#692090000000
1!
1*
b110 6
19
1>
1C
b110 G
#692100000000
0!
0*
09
0>
0C
#692110000000
1!
1*
b111 6
19
1>
1C
b111 G
#692120000000
0!
0*
09
0>
0C
#692130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#692140000000
0!
0*
09
0>
0C
#692150000000
1!
1*
b1 6
19
1>
1C
b1 G
#692160000000
0!
0*
09
0>
0C
#692170000000
1!
1*
b10 6
19
1>
1C
b10 G
#692180000000
0!
0*
09
0>
0C
#692190000000
1!
1*
b11 6
19
1>
1C
b11 G
#692200000000
0!
0*
09
0>
0C
#692210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#692220000000
0!
0*
09
0>
0C
#692230000000
1!
1*
b101 6
19
1>
1C
b101 G
#692240000000
0!
0*
09
0>
0C
#692250000000
1!
1*
b110 6
19
1>
1C
b110 G
#692260000000
0!
0*
09
0>
0C
#692270000000
1!
1*
b111 6
19
1>
1C
b111 G
#692280000000
0!
1"
0*
1+
09
1:
0>
0C
#692290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#692300000000
0!
0*
09
0>
0C
#692310000000
1!
1*
b1 6
19
1>
1C
b1 G
#692320000000
0!
0*
09
0>
0C
#692330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#692340000000
0!
0*
09
0>
0C
#692350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#692360000000
0!
0*
09
0>
0C
#692370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#692380000000
0!
0*
09
0>
0C
#692390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#692400000000
0!
0#
0*
0,
09
0>
0?
0C
#692410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#692420000000
0!
0*
09
0>
0C
#692430000000
1!
1*
19
1>
1C
#692440000000
0!
0*
09
0>
0C
#692450000000
1!
1*
19
1>
1C
#692460000000
0!
0*
09
0>
0C
#692470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#692480000000
0!
0*
09
0>
0C
#692490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#692500000000
0!
0*
09
0>
0C
#692510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#692520000000
0!
0*
09
0>
0C
#692530000000
1!
1*
b10 6
19
1>
1C
b10 G
#692540000000
0!
0*
09
0>
0C
#692550000000
1!
1*
b11 6
19
1>
1C
b11 G
#692560000000
0!
0*
09
0>
0C
#692570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#692580000000
0!
0*
09
0>
0C
#692590000000
1!
1*
b101 6
19
1>
1C
b101 G
#692600000000
0!
0*
09
0>
0C
#692610000000
1!
1*
b110 6
19
1>
1C
b110 G
#692620000000
0!
0*
09
0>
0C
#692630000000
1!
1*
b111 6
19
1>
1C
b111 G
#692640000000
0!
0*
09
0>
0C
#692650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#692660000000
0!
0*
09
0>
0C
#692670000000
1!
1*
b1 6
19
1>
1C
b1 G
#692680000000
0!
0*
09
0>
0C
#692690000000
1!
1*
b10 6
19
1>
1C
b10 G
#692700000000
0!
0*
09
0>
0C
#692710000000
1!
1*
b11 6
19
1>
1C
b11 G
#692720000000
0!
0*
09
0>
0C
#692730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#692740000000
0!
0*
09
0>
0C
#692750000000
1!
1*
b101 6
19
1>
1C
b101 G
#692760000000
0!
0*
09
0>
0C
#692770000000
1!
1*
b110 6
19
1>
1C
b110 G
#692780000000
0!
0*
09
0>
0C
#692790000000
1!
1*
b111 6
19
1>
1C
b111 G
#692800000000
0!
0*
09
0>
0C
#692810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#692820000000
0!
0*
09
0>
0C
#692830000000
1!
1*
b1 6
19
1>
1C
b1 G
#692840000000
0!
0*
09
0>
0C
#692850000000
1!
1*
b10 6
19
1>
1C
b10 G
#692860000000
0!
0*
09
0>
0C
#692870000000
1!
1*
b11 6
19
1>
1C
b11 G
#692880000000
0!
0*
09
0>
0C
#692890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#692900000000
0!
0*
09
0>
0C
#692910000000
1!
1*
b101 6
19
1>
1C
b101 G
#692920000000
0!
0*
09
0>
0C
#692930000000
1!
1*
b110 6
19
1>
1C
b110 G
#692940000000
0!
0*
09
0>
0C
#692950000000
1!
1*
b111 6
19
1>
1C
b111 G
#692960000000
0!
1"
0*
1+
09
1:
0>
0C
#692970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#692980000000
0!
0*
09
0>
0C
#692990000000
1!
1*
b1 6
19
1>
1C
b1 G
#693000000000
0!
0*
09
0>
0C
#693010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#693020000000
0!
0*
09
0>
0C
#693030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#693040000000
0!
0*
09
0>
0C
#693050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#693060000000
0!
0*
09
0>
0C
#693070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#693080000000
0!
0#
0*
0,
09
0>
0?
0C
#693090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#693100000000
0!
0*
09
0>
0C
#693110000000
1!
1*
19
1>
1C
#693120000000
0!
0*
09
0>
0C
#693130000000
1!
1*
19
1>
1C
#693140000000
0!
0*
09
0>
0C
#693150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#693160000000
0!
0*
09
0>
0C
#693170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#693180000000
0!
0*
09
0>
0C
#693190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#693200000000
0!
0*
09
0>
0C
#693210000000
1!
1*
b10 6
19
1>
1C
b10 G
#693220000000
0!
0*
09
0>
0C
#693230000000
1!
1*
b11 6
19
1>
1C
b11 G
#693240000000
0!
0*
09
0>
0C
#693250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#693260000000
0!
0*
09
0>
0C
#693270000000
1!
1*
b101 6
19
1>
1C
b101 G
#693280000000
0!
0*
09
0>
0C
#693290000000
1!
1*
b110 6
19
1>
1C
b110 G
#693300000000
0!
0*
09
0>
0C
#693310000000
1!
1*
b111 6
19
1>
1C
b111 G
#693320000000
0!
0*
09
0>
0C
#693330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#693340000000
0!
0*
09
0>
0C
#693350000000
1!
1*
b1 6
19
1>
1C
b1 G
#693360000000
0!
0*
09
0>
0C
#693370000000
1!
1*
b10 6
19
1>
1C
b10 G
#693380000000
0!
0*
09
0>
0C
#693390000000
1!
1*
b11 6
19
1>
1C
b11 G
#693400000000
0!
0*
09
0>
0C
#693410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#693420000000
0!
0*
09
0>
0C
#693430000000
1!
1*
b101 6
19
1>
1C
b101 G
#693440000000
0!
0*
09
0>
0C
#693450000000
1!
1*
b110 6
19
1>
1C
b110 G
#693460000000
0!
0*
09
0>
0C
#693470000000
1!
1*
b111 6
19
1>
1C
b111 G
#693480000000
0!
0*
09
0>
0C
#693490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#693500000000
0!
0*
09
0>
0C
#693510000000
1!
1*
b1 6
19
1>
1C
b1 G
#693520000000
0!
0*
09
0>
0C
#693530000000
1!
1*
b10 6
19
1>
1C
b10 G
#693540000000
0!
0*
09
0>
0C
#693550000000
1!
1*
b11 6
19
1>
1C
b11 G
#693560000000
0!
0*
09
0>
0C
#693570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#693580000000
0!
0*
09
0>
0C
#693590000000
1!
1*
b101 6
19
1>
1C
b101 G
#693600000000
0!
0*
09
0>
0C
#693610000000
1!
1*
b110 6
19
1>
1C
b110 G
#693620000000
0!
0*
09
0>
0C
#693630000000
1!
1*
b111 6
19
1>
1C
b111 G
#693640000000
0!
1"
0*
1+
09
1:
0>
0C
#693650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#693660000000
0!
0*
09
0>
0C
#693670000000
1!
1*
b1 6
19
1>
1C
b1 G
#693680000000
0!
0*
09
0>
0C
#693690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#693700000000
0!
0*
09
0>
0C
#693710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#693720000000
0!
0*
09
0>
0C
#693730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#693740000000
0!
0*
09
0>
0C
#693750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#693760000000
0!
0#
0*
0,
09
0>
0?
0C
#693770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#693780000000
0!
0*
09
0>
0C
#693790000000
1!
1*
19
1>
1C
#693800000000
0!
0*
09
0>
0C
#693810000000
1!
1*
19
1>
1C
#693820000000
0!
0*
09
0>
0C
#693830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#693840000000
0!
0*
09
0>
0C
#693850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#693860000000
0!
0*
09
0>
0C
#693870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#693880000000
0!
0*
09
0>
0C
#693890000000
1!
1*
b10 6
19
1>
1C
b10 G
#693900000000
0!
0*
09
0>
0C
#693910000000
1!
1*
b11 6
19
1>
1C
b11 G
#693920000000
0!
0*
09
0>
0C
#693930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#693940000000
0!
0*
09
0>
0C
#693950000000
1!
1*
b101 6
19
1>
1C
b101 G
#693960000000
0!
0*
09
0>
0C
#693970000000
1!
1*
b110 6
19
1>
1C
b110 G
#693980000000
0!
0*
09
0>
0C
#693990000000
1!
1*
b111 6
19
1>
1C
b111 G
#694000000000
0!
0*
09
0>
0C
#694010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#694020000000
0!
0*
09
0>
0C
#694030000000
1!
1*
b1 6
19
1>
1C
b1 G
#694040000000
0!
0*
09
0>
0C
#694050000000
1!
1*
b10 6
19
1>
1C
b10 G
#694060000000
0!
0*
09
0>
0C
#694070000000
1!
1*
b11 6
19
1>
1C
b11 G
#694080000000
0!
0*
09
0>
0C
#694090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#694100000000
0!
0*
09
0>
0C
#694110000000
1!
1*
b101 6
19
1>
1C
b101 G
#694120000000
0!
0*
09
0>
0C
#694130000000
1!
1*
b110 6
19
1>
1C
b110 G
#694140000000
0!
0*
09
0>
0C
#694150000000
1!
1*
b111 6
19
1>
1C
b111 G
#694160000000
0!
0*
09
0>
0C
#694170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#694180000000
0!
0*
09
0>
0C
#694190000000
1!
1*
b1 6
19
1>
1C
b1 G
#694200000000
0!
0*
09
0>
0C
#694210000000
1!
1*
b10 6
19
1>
1C
b10 G
#694220000000
0!
0*
09
0>
0C
#694230000000
1!
1*
b11 6
19
1>
1C
b11 G
#694240000000
0!
0*
09
0>
0C
#694250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#694260000000
0!
0*
09
0>
0C
#694270000000
1!
1*
b101 6
19
1>
1C
b101 G
#694280000000
0!
0*
09
0>
0C
#694290000000
1!
1*
b110 6
19
1>
1C
b110 G
#694300000000
0!
0*
09
0>
0C
#694310000000
1!
1*
b111 6
19
1>
1C
b111 G
#694320000000
0!
1"
0*
1+
09
1:
0>
0C
#694330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#694340000000
0!
0*
09
0>
0C
#694350000000
1!
1*
b1 6
19
1>
1C
b1 G
#694360000000
0!
0*
09
0>
0C
#694370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#694380000000
0!
0*
09
0>
0C
#694390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#694400000000
0!
0*
09
0>
0C
#694410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#694420000000
0!
0*
09
0>
0C
#694430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#694440000000
0!
0#
0*
0,
09
0>
0?
0C
#694450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#694460000000
0!
0*
09
0>
0C
#694470000000
1!
1*
19
1>
1C
#694480000000
0!
0*
09
0>
0C
#694490000000
1!
1*
19
1>
1C
#694500000000
0!
0*
09
0>
0C
#694510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#694520000000
0!
0*
09
0>
0C
#694530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#694540000000
0!
0*
09
0>
0C
#694550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#694560000000
0!
0*
09
0>
0C
#694570000000
1!
1*
b10 6
19
1>
1C
b10 G
#694580000000
0!
0*
09
0>
0C
#694590000000
1!
1*
b11 6
19
1>
1C
b11 G
#694600000000
0!
0*
09
0>
0C
#694610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#694620000000
0!
0*
09
0>
0C
#694630000000
1!
1*
b101 6
19
1>
1C
b101 G
#694640000000
0!
0*
09
0>
0C
#694650000000
1!
1*
b110 6
19
1>
1C
b110 G
#694660000000
0!
0*
09
0>
0C
#694670000000
1!
1*
b111 6
19
1>
1C
b111 G
#694680000000
0!
0*
09
0>
0C
#694690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#694700000000
0!
0*
09
0>
0C
#694710000000
1!
1*
b1 6
19
1>
1C
b1 G
#694720000000
0!
0*
09
0>
0C
#694730000000
1!
1*
b10 6
19
1>
1C
b10 G
#694740000000
0!
0*
09
0>
0C
#694750000000
1!
1*
b11 6
19
1>
1C
b11 G
#694760000000
0!
0*
09
0>
0C
#694770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#694780000000
0!
0*
09
0>
0C
#694790000000
1!
1*
b101 6
19
1>
1C
b101 G
#694800000000
0!
0*
09
0>
0C
#694810000000
1!
1*
b110 6
19
1>
1C
b110 G
#694820000000
0!
0*
09
0>
0C
#694830000000
1!
1*
b111 6
19
1>
1C
b111 G
#694840000000
0!
0*
09
0>
0C
#694850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#694860000000
0!
0*
09
0>
0C
#694870000000
1!
1*
b1 6
19
1>
1C
b1 G
#694880000000
0!
0*
09
0>
0C
#694890000000
1!
1*
b10 6
19
1>
1C
b10 G
#694900000000
0!
0*
09
0>
0C
#694910000000
1!
1*
b11 6
19
1>
1C
b11 G
#694920000000
0!
0*
09
0>
0C
#694930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#694940000000
0!
0*
09
0>
0C
#694950000000
1!
1*
b101 6
19
1>
1C
b101 G
#694960000000
0!
0*
09
0>
0C
#694970000000
1!
1*
b110 6
19
1>
1C
b110 G
#694980000000
0!
0*
09
0>
0C
#694990000000
1!
1*
b111 6
19
1>
1C
b111 G
#695000000000
0!
1"
0*
1+
09
1:
0>
0C
#695010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#695020000000
0!
0*
09
0>
0C
#695030000000
1!
1*
b1 6
19
1>
1C
b1 G
#695040000000
0!
0*
09
0>
0C
#695050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#695060000000
0!
0*
09
0>
0C
#695070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#695080000000
0!
0*
09
0>
0C
#695090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#695100000000
0!
0*
09
0>
0C
#695110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#695120000000
0!
0#
0*
0,
09
0>
0?
0C
#695130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#695140000000
0!
0*
09
0>
0C
#695150000000
1!
1*
19
1>
1C
#695160000000
0!
0*
09
0>
0C
#695170000000
1!
1*
19
1>
1C
#695180000000
0!
0*
09
0>
0C
#695190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#695200000000
0!
0*
09
0>
0C
#695210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#695220000000
0!
0*
09
0>
0C
#695230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#695240000000
0!
0*
09
0>
0C
#695250000000
1!
1*
b10 6
19
1>
1C
b10 G
#695260000000
0!
0*
09
0>
0C
#695270000000
1!
1*
b11 6
19
1>
1C
b11 G
#695280000000
0!
0*
09
0>
0C
#695290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#695300000000
0!
0*
09
0>
0C
#695310000000
1!
1*
b101 6
19
1>
1C
b101 G
#695320000000
0!
0*
09
0>
0C
#695330000000
1!
1*
b110 6
19
1>
1C
b110 G
#695340000000
0!
0*
09
0>
0C
#695350000000
1!
1*
b111 6
19
1>
1C
b111 G
#695360000000
0!
0*
09
0>
0C
#695370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#695380000000
0!
0*
09
0>
0C
#695390000000
1!
1*
b1 6
19
1>
1C
b1 G
#695400000000
0!
0*
09
0>
0C
#695410000000
1!
1*
b10 6
19
1>
1C
b10 G
#695420000000
0!
0*
09
0>
0C
#695430000000
1!
1*
b11 6
19
1>
1C
b11 G
#695440000000
0!
0*
09
0>
0C
#695450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#695460000000
0!
0*
09
0>
0C
#695470000000
1!
1*
b101 6
19
1>
1C
b101 G
#695480000000
0!
0*
09
0>
0C
#695490000000
1!
1*
b110 6
19
1>
1C
b110 G
#695500000000
0!
0*
09
0>
0C
#695510000000
1!
1*
b111 6
19
1>
1C
b111 G
#695520000000
0!
0*
09
0>
0C
#695530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#695540000000
0!
0*
09
0>
0C
#695550000000
1!
1*
b1 6
19
1>
1C
b1 G
#695560000000
0!
0*
09
0>
0C
#695570000000
1!
1*
b10 6
19
1>
1C
b10 G
#695580000000
0!
0*
09
0>
0C
#695590000000
1!
1*
b11 6
19
1>
1C
b11 G
#695600000000
0!
0*
09
0>
0C
#695610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#695620000000
0!
0*
09
0>
0C
#695630000000
1!
1*
b101 6
19
1>
1C
b101 G
#695640000000
0!
0*
09
0>
0C
#695650000000
1!
1*
b110 6
19
1>
1C
b110 G
#695660000000
0!
0*
09
0>
0C
#695670000000
1!
1*
b111 6
19
1>
1C
b111 G
#695680000000
0!
1"
0*
1+
09
1:
0>
0C
#695690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#695700000000
0!
0*
09
0>
0C
#695710000000
1!
1*
b1 6
19
1>
1C
b1 G
#695720000000
0!
0*
09
0>
0C
#695730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#695740000000
0!
0*
09
0>
0C
#695750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#695760000000
0!
0*
09
0>
0C
#695770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#695780000000
0!
0*
09
0>
0C
#695790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#695800000000
0!
0#
0*
0,
09
0>
0?
0C
#695810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#695820000000
0!
0*
09
0>
0C
#695830000000
1!
1*
19
1>
1C
#695840000000
0!
0*
09
0>
0C
#695850000000
1!
1*
19
1>
1C
#695860000000
0!
0*
09
0>
0C
#695870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#695880000000
0!
0*
09
0>
0C
#695890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#695900000000
0!
0*
09
0>
0C
#695910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#695920000000
0!
0*
09
0>
0C
#695930000000
1!
1*
b10 6
19
1>
1C
b10 G
#695940000000
0!
0*
09
0>
0C
#695950000000
1!
1*
b11 6
19
1>
1C
b11 G
#695960000000
0!
0*
09
0>
0C
#695970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#695980000000
0!
0*
09
0>
0C
#695990000000
1!
1*
b101 6
19
1>
1C
b101 G
#696000000000
0!
0*
09
0>
0C
#696010000000
1!
1*
b110 6
19
1>
1C
b110 G
#696020000000
0!
0*
09
0>
0C
#696030000000
1!
1*
b111 6
19
1>
1C
b111 G
#696040000000
0!
0*
09
0>
0C
#696050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#696060000000
0!
0*
09
0>
0C
#696070000000
1!
1*
b1 6
19
1>
1C
b1 G
#696080000000
0!
0*
09
0>
0C
#696090000000
1!
1*
b10 6
19
1>
1C
b10 G
#696100000000
0!
0*
09
0>
0C
#696110000000
1!
1*
b11 6
19
1>
1C
b11 G
#696120000000
0!
0*
09
0>
0C
#696130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#696140000000
0!
0*
09
0>
0C
#696150000000
1!
1*
b101 6
19
1>
1C
b101 G
#696160000000
0!
0*
09
0>
0C
#696170000000
1!
1*
b110 6
19
1>
1C
b110 G
#696180000000
0!
0*
09
0>
0C
#696190000000
1!
1*
b111 6
19
1>
1C
b111 G
#696200000000
0!
0*
09
0>
0C
#696210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#696220000000
0!
0*
09
0>
0C
#696230000000
1!
1*
b1 6
19
1>
1C
b1 G
#696240000000
0!
0*
09
0>
0C
#696250000000
1!
1*
b10 6
19
1>
1C
b10 G
#696260000000
0!
0*
09
0>
0C
#696270000000
1!
1*
b11 6
19
1>
1C
b11 G
#696280000000
0!
0*
09
0>
0C
#696290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#696300000000
0!
0*
09
0>
0C
#696310000000
1!
1*
b101 6
19
1>
1C
b101 G
#696320000000
0!
0*
09
0>
0C
#696330000000
1!
1*
b110 6
19
1>
1C
b110 G
#696340000000
0!
0*
09
0>
0C
#696350000000
1!
1*
b111 6
19
1>
1C
b111 G
#696360000000
0!
1"
0*
1+
09
1:
0>
0C
#696370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#696380000000
0!
0*
09
0>
0C
#696390000000
1!
1*
b1 6
19
1>
1C
b1 G
#696400000000
0!
0*
09
0>
0C
#696410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#696420000000
0!
0*
09
0>
0C
#696430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#696440000000
0!
0*
09
0>
0C
#696450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#696460000000
0!
0*
09
0>
0C
#696470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#696480000000
0!
0#
0*
0,
09
0>
0?
0C
#696490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#696500000000
0!
0*
09
0>
0C
#696510000000
1!
1*
19
1>
1C
#696520000000
0!
0*
09
0>
0C
#696530000000
1!
1*
19
1>
1C
#696540000000
0!
0*
09
0>
0C
#696550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#696560000000
0!
0*
09
0>
0C
#696570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#696580000000
0!
0*
09
0>
0C
#696590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#696600000000
0!
0*
09
0>
0C
#696610000000
1!
1*
b10 6
19
1>
1C
b10 G
#696620000000
0!
0*
09
0>
0C
#696630000000
1!
1*
b11 6
19
1>
1C
b11 G
#696640000000
0!
0*
09
0>
0C
#696650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#696660000000
0!
0*
09
0>
0C
#696670000000
1!
1*
b101 6
19
1>
1C
b101 G
#696680000000
0!
0*
09
0>
0C
#696690000000
1!
1*
b110 6
19
1>
1C
b110 G
#696700000000
0!
0*
09
0>
0C
#696710000000
1!
1*
b111 6
19
1>
1C
b111 G
#696720000000
0!
0*
09
0>
0C
#696730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#696740000000
0!
0*
09
0>
0C
#696750000000
1!
1*
b1 6
19
1>
1C
b1 G
#696760000000
0!
0*
09
0>
0C
#696770000000
1!
1*
b10 6
19
1>
1C
b10 G
#696780000000
0!
0*
09
0>
0C
#696790000000
1!
1*
b11 6
19
1>
1C
b11 G
#696800000000
0!
0*
09
0>
0C
#696810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#696820000000
0!
0*
09
0>
0C
#696830000000
1!
1*
b101 6
19
1>
1C
b101 G
#696840000000
0!
0*
09
0>
0C
#696850000000
1!
1*
b110 6
19
1>
1C
b110 G
#696860000000
0!
0*
09
0>
0C
#696870000000
1!
1*
b111 6
19
1>
1C
b111 G
#696880000000
0!
0*
09
0>
0C
#696890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#696900000000
0!
0*
09
0>
0C
#696910000000
1!
1*
b1 6
19
1>
1C
b1 G
#696920000000
0!
0*
09
0>
0C
#696930000000
1!
1*
b10 6
19
1>
1C
b10 G
#696940000000
0!
0*
09
0>
0C
#696950000000
1!
1*
b11 6
19
1>
1C
b11 G
#696960000000
0!
0*
09
0>
0C
#696970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#696980000000
0!
0*
09
0>
0C
#696990000000
1!
1*
b101 6
19
1>
1C
b101 G
#697000000000
0!
0*
09
0>
0C
#697010000000
1!
1*
b110 6
19
1>
1C
b110 G
#697020000000
0!
0*
09
0>
0C
#697030000000
1!
1*
b111 6
19
1>
1C
b111 G
#697040000000
0!
1"
0*
1+
09
1:
0>
0C
#697050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#697060000000
0!
0*
09
0>
0C
#697070000000
1!
1*
b1 6
19
1>
1C
b1 G
#697080000000
0!
0*
09
0>
0C
#697090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#697100000000
0!
0*
09
0>
0C
#697110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#697120000000
0!
0*
09
0>
0C
#697130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#697140000000
0!
0*
09
0>
0C
#697150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#697160000000
0!
0#
0*
0,
09
0>
0?
0C
#697170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#697180000000
0!
0*
09
0>
0C
#697190000000
1!
1*
19
1>
1C
#697200000000
0!
0*
09
0>
0C
#697210000000
1!
1*
19
1>
1C
#697220000000
0!
0*
09
0>
0C
#697230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#697240000000
0!
0*
09
0>
0C
#697250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#697260000000
0!
0*
09
0>
0C
#697270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#697280000000
0!
0*
09
0>
0C
#697290000000
1!
1*
b10 6
19
1>
1C
b10 G
#697300000000
0!
0*
09
0>
0C
#697310000000
1!
1*
b11 6
19
1>
1C
b11 G
#697320000000
0!
0*
09
0>
0C
#697330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#697340000000
0!
0*
09
0>
0C
#697350000000
1!
1*
b101 6
19
1>
1C
b101 G
#697360000000
0!
0*
09
0>
0C
#697370000000
1!
1*
b110 6
19
1>
1C
b110 G
#697380000000
0!
0*
09
0>
0C
#697390000000
1!
1*
b111 6
19
1>
1C
b111 G
#697400000000
0!
0*
09
0>
0C
#697410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#697420000000
0!
0*
09
0>
0C
#697430000000
1!
1*
b1 6
19
1>
1C
b1 G
#697440000000
0!
0*
09
0>
0C
#697450000000
1!
1*
b10 6
19
1>
1C
b10 G
#697460000000
0!
0*
09
0>
0C
#697470000000
1!
1*
b11 6
19
1>
1C
b11 G
#697480000000
0!
0*
09
0>
0C
#697490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#697500000000
0!
0*
09
0>
0C
#697510000000
1!
1*
b101 6
19
1>
1C
b101 G
#697520000000
0!
0*
09
0>
0C
#697530000000
1!
1*
b110 6
19
1>
1C
b110 G
#697540000000
0!
0*
09
0>
0C
#697550000000
1!
1*
b111 6
19
1>
1C
b111 G
#697560000000
0!
0*
09
0>
0C
#697570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#697580000000
0!
0*
09
0>
0C
#697590000000
1!
1*
b1 6
19
1>
1C
b1 G
#697600000000
0!
0*
09
0>
0C
#697610000000
1!
1*
b10 6
19
1>
1C
b10 G
#697620000000
0!
0*
09
0>
0C
#697630000000
1!
1*
b11 6
19
1>
1C
b11 G
#697640000000
0!
0*
09
0>
0C
#697650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#697660000000
0!
0*
09
0>
0C
#697670000000
1!
1*
b101 6
19
1>
1C
b101 G
#697680000000
0!
0*
09
0>
0C
#697690000000
1!
1*
b110 6
19
1>
1C
b110 G
#697700000000
0!
0*
09
0>
0C
#697710000000
1!
1*
b111 6
19
1>
1C
b111 G
#697720000000
0!
1"
0*
1+
09
1:
0>
0C
#697730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#697740000000
0!
0*
09
0>
0C
#697750000000
1!
1*
b1 6
19
1>
1C
b1 G
#697760000000
0!
0*
09
0>
0C
#697770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#697780000000
0!
0*
09
0>
0C
#697790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#697800000000
0!
0*
09
0>
0C
#697810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#697820000000
0!
0*
09
0>
0C
#697830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#697840000000
0!
0#
0*
0,
09
0>
0?
0C
#697850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#697860000000
0!
0*
09
0>
0C
#697870000000
1!
1*
19
1>
1C
#697880000000
0!
0*
09
0>
0C
#697890000000
1!
1*
19
1>
1C
#697900000000
0!
0*
09
0>
0C
#697910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#697920000000
0!
0*
09
0>
0C
#697930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#697940000000
0!
0*
09
0>
0C
#697950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#697960000000
0!
0*
09
0>
0C
#697970000000
1!
1*
b10 6
19
1>
1C
b10 G
#697980000000
0!
0*
09
0>
0C
#697990000000
1!
1*
b11 6
19
1>
1C
b11 G
#698000000000
0!
0*
09
0>
0C
#698010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#698020000000
0!
0*
09
0>
0C
#698030000000
1!
1*
b101 6
19
1>
1C
b101 G
#698040000000
0!
0*
09
0>
0C
#698050000000
1!
1*
b110 6
19
1>
1C
b110 G
#698060000000
0!
0*
09
0>
0C
#698070000000
1!
1*
b111 6
19
1>
1C
b111 G
#698080000000
0!
0*
09
0>
0C
#698090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#698100000000
0!
0*
09
0>
0C
#698110000000
1!
1*
b1 6
19
1>
1C
b1 G
#698120000000
0!
0*
09
0>
0C
#698130000000
1!
1*
b10 6
19
1>
1C
b10 G
#698140000000
0!
0*
09
0>
0C
#698150000000
1!
1*
b11 6
19
1>
1C
b11 G
#698160000000
0!
0*
09
0>
0C
#698170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#698180000000
0!
0*
09
0>
0C
#698190000000
1!
1*
b101 6
19
1>
1C
b101 G
#698200000000
0!
0*
09
0>
0C
#698210000000
1!
1*
b110 6
19
1>
1C
b110 G
#698220000000
0!
0*
09
0>
0C
#698230000000
1!
1*
b111 6
19
1>
1C
b111 G
#698240000000
0!
0*
09
0>
0C
#698250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#698260000000
0!
0*
09
0>
0C
#698270000000
1!
1*
b1 6
19
1>
1C
b1 G
#698280000000
0!
0*
09
0>
0C
#698290000000
1!
1*
b10 6
19
1>
1C
b10 G
#698300000000
0!
0*
09
0>
0C
#698310000000
1!
1*
b11 6
19
1>
1C
b11 G
#698320000000
0!
0*
09
0>
0C
#698330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#698340000000
0!
0*
09
0>
0C
#698350000000
1!
1*
b101 6
19
1>
1C
b101 G
#698360000000
0!
0*
09
0>
0C
#698370000000
1!
1*
b110 6
19
1>
1C
b110 G
#698380000000
0!
0*
09
0>
0C
#698390000000
1!
1*
b111 6
19
1>
1C
b111 G
#698400000000
0!
1"
0*
1+
09
1:
0>
0C
#698410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#698420000000
0!
0*
09
0>
0C
#698430000000
1!
1*
b1 6
19
1>
1C
b1 G
#698440000000
0!
0*
09
0>
0C
#698450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#698460000000
0!
0*
09
0>
0C
#698470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#698480000000
0!
0*
09
0>
0C
#698490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#698500000000
0!
0*
09
0>
0C
#698510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#698520000000
0!
0#
0*
0,
09
0>
0?
0C
#698530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#698540000000
0!
0*
09
0>
0C
#698550000000
1!
1*
19
1>
1C
#698560000000
0!
0*
09
0>
0C
#698570000000
1!
1*
19
1>
1C
#698580000000
0!
0*
09
0>
0C
#698590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#698600000000
0!
0*
09
0>
0C
#698610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#698620000000
0!
0*
09
0>
0C
#698630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#698640000000
0!
0*
09
0>
0C
#698650000000
1!
1*
b10 6
19
1>
1C
b10 G
#698660000000
0!
0*
09
0>
0C
#698670000000
1!
1*
b11 6
19
1>
1C
b11 G
#698680000000
0!
0*
09
0>
0C
#698690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#698700000000
0!
0*
09
0>
0C
#698710000000
1!
1*
b101 6
19
1>
1C
b101 G
#698720000000
0!
0*
09
0>
0C
#698730000000
1!
1*
b110 6
19
1>
1C
b110 G
#698740000000
0!
0*
09
0>
0C
#698750000000
1!
1*
b111 6
19
1>
1C
b111 G
#698760000000
0!
0*
09
0>
0C
#698770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#698780000000
0!
0*
09
0>
0C
#698790000000
1!
1*
b1 6
19
1>
1C
b1 G
#698800000000
0!
0*
09
0>
0C
#698810000000
1!
1*
b10 6
19
1>
1C
b10 G
#698820000000
0!
0*
09
0>
0C
#698830000000
1!
1*
b11 6
19
1>
1C
b11 G
#698840000000
0!
0*
09
0>
0C
#698850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#698860000000
0!
0*
09
0>
0C
#698870000000
1!
1*
b101 6
19
1>
1C
b101 G
#698880000000
0!
0*
09
0>
0C
#698890000000
1!
1*
b110 6
19
1>
1C
b110 G
#698900000000
0!
0*
09
0>
0C
#698910000000
1!
1*
b111 6
19
1>
1C
b111 G
#698920000000
0!
0*
09
0>
0C
#698930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#698940000000
0!
0*
09
0>
0C
#698950000000
1!
1*
b1 6
19
1>
1C
b1 G
#698960000000
0!
0*
09
0>
0C
#698970000000
1!
1*
b10 6
19
1>
1C
b10 G
#698980000000
0!
0*
09
0>
0C
#698990000000
1!
1*
b11 6
19
1>
1C
b11 G
#699000000000
0!
0*
09
0>
0C
#699010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#699020000000
0!
0*
09
0>
0C
#699030000000
1!
1*
b101 6
19
1>
1C
b101 G
#699040000000
0!
0*
09
0>
0C
#699050000000
1!
1*
b110 6
19
1>
1C
b110 G
#699060000000
0!
0*
09
0>
0C
#699070000000
1!
1*
b111 6
19
1>
1C
b111 G
#699080000000
0!
1"
0*
1+
09
1:
0>
0C
#699090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#699100000000
0!
0*
09
0>
0C
#699110000000
1!
1*
b1 6
19
1>
1C
b1 G
#699120000000
0!
0*
09
0>
0C
#699130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#699140000000
0!
0*
09
0>
0C
#699150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#699160000000
0!
0*
09
0>
0C
#699170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#699180000000
0!
0*
09
0>
0C
#699190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#699200000000
0!
0#
0*
0,
09
0>
0?
0C
#699210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#699220000000
0!
0*
09
0>
0C
#699230000000
1!
1*
19
1>
1C
#699240000000
0!
0*
09
0>
0C
#699250000000
1!
1*
19
1>
1C
#699260000000
0!
0*
09
0>
0C
#699270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#699280000000
0!
0*
09
0>
0C
#699290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#699300000000
0!
0*
09
0>
0C
#699310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#699320000000
0!
0*
09
0>
0C
#699330000000
1!
1*
b10 6
19
1>
1C
b10 G
#699340000000
0!
0*
09
0>
0C
#699350000000
1!
1*
b11 6
19
1>
1C
b11 G
#699360000000
0!
0*
09
0>
0C
#699370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#699380000000
0!
0*
09
0>
0C
#699390000000
1!
1*
b101 6
19
1>
1C
b101 G
#699400000000
0!
0*
09
0>
0C
#699410000000
1!
1*
b110 6
19
1>
1C
b110 G
#699420000000
0!
0*
09
0>
0C
#699430000000
1!
1*
b111 6
19
1>
1C
b111 G
#699440000000
0!
0*
09
0>
0C
#699450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#699460000000
0!
0*
09
0>
0C
#699470000000
1!
1*
b1 6
19
1>
1C
b1 G
#699480000000
0!
0*
09
0>
0C
#699490000000
1!
1*
b10 6
19
1>
1C
b10 G
#699500000000
0!
0*
09
0>
0C
#699510000000
1!
1*
b11 6
19
1>
1C
b11 G
#699520000000
0!
0*
09
0>
0C
#699530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#699540000000
0!
0*
09
0>
0C
#699550000000
1!
1*
b101 6
19
1>
1C
b101 G
#699560000000
0!
0*
09
0>
0C
#699570000000
1!
1*
b110 6
19
1>
1C
b110 G
#699580000000
0!
0*
09
0>
0C
#699590000000
1!
1*
b111 6
19
1>
1C
b111 G
#699600000000
0!
0*
09
0>
0C
#699610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#699620000000
0!
0*
09
0>
0C
#699630000000
1!
1*
b1 6
19
1>
1C
b1 G
#699640000000
0!
0*
09
0>
0C
#699650000000
1!
1*
b10 6
19
1>
1C
b10 G
#699660000000
0!
0*
09
0>
0C
#699670000000
1!
1*
b11 6
19
1>
1C
b11 G
#699680000000
0!
0*
09
0>
0C
#699690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#699700000000
0!
0*
09
0>
0C
#699710000000
1!
1*
b101 6
19
1>
1C
b101 G
#699720000000
0!
0*
09
0>
0C
#699730000000
1!
1*
b110 6
19
1>
1C
b110 G
#699740000000
0!
0*
09
0>
0C
#699750000000
1!
1*
b111 6
19
1>
1C
b111 G
#699760000000
0!
1"
0*
1+
09
1:
0>
0C
#699770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#699780000000
0!
0*
09
0>
0C
#699790000000
1!
1*
b1 6
19
1>
1C
b1 G
#699800000000
0!
0*
09
0>
0C
#699810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#699820000000
0!
0*
09
0>
0C
#699830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#699840000000
0!
0*
09
0>
0C
#699850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#699860000000
0!
0*
09
0>
0C
#699870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#699880000000
0!
0#
0*
0,
09
0>
0?
0C
#699890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#699900000000
0!
0*
09
0>
0C
#699910000000
1!
1*
19
1>
1C
#699920000000
0!
0*
09
0>
0C
#699930000000
1!
1*
19
1>
1C
#699940000000
0!
0*
09
0>
0C
#699950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#699960000000
0!
0*
09
0>
0C
#699970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#699980000000
0!
0*
09
0>
0C
#699990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#700000000000
0!
0*
09
0>
0C
#700010000000
1!
1*
b10 6
19
1>
1C
b10 G
#700020000000
0!
0*
09
0>
0C
#700030000000
1!
1*
b11 6
19
1>
1C
b11 G
#700040000000
0!
0*
09
0>
0C
#700050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#700060000000
0!
0*
09
0>
0C
#700070000000
1!
1*
b101 6
19
1>
1C
b101 G
#700080000000
0!
0*
09
0>
0C
#700090000000
1!
1*
b110 6
19
1>
1C
b110 G
#700100000000
0!
0*
09
0>
0C
#700110000000
1!
1*
b111 6
19
1>
1C
b111 G
#700120000000
0!
0*
09
0>
0C
#700130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#700140000000
0!
0*
09
0>
0C
#700150000000
1!
1*
b1 6
19
1>
1C
b1 G
#700160000000
0!
0*
09
0>
0C
#700170000000
1!
1*
b10 6
19
1>
1C
b10 G
#700180000000
0!
0*
09
0>
0C
#700190000000
1!
1*
b11 6
19
1>
1C
b11 G
#700200000000
0!
0*
09
0>
0C
#700210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#700220000000
0!
0*
09
0>
0C
#700230000000
1!
1*
b101 6
19
1>
1C
b101 G
#700240000000
0!
0*
09
0>
0C
#700250000000
1!
1*
b110 6
19
1>
1C
b110 G
#700260000000
0!
0*
09
0>
0C
#700270000000
1!
1*
b111 6
19
1>
1C
b111 G
#700280000000
0!
0*
09
0>
0C
#700290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#700300000000
0!
0*
09
0>
0C
#700310000000
1!
1*
b1 6
19
1>
1C
b1 G
#700320000000
0!
0*
09
0>
0C
#700330000000
1!
1*
b10 6
19
1>
1C
b10 G
#700340000000
0!
0*
09
0>
0C
#700350000000
1!
1*
b11 6
19
1>
1C
b11 G
#700360000000
0!
0*
09
0>
0C
#700370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#700380000000
0!
0*
09
0>
0C
#700390000000
1!
1*
b101 6
19
1>
1C
b101 G
#700400000000
0!
0*
09
0>
0C
#700410000000
1!
1*
b110 6
19
1>
1C
b110 G
#700420000000
0!
0*
09
0>
0C
#700430000000
1!
1*
b111 6
19
1>
1C
b111 G
#700440000000
0!
1"
0*
1+
09
1:
0>
0C
#700450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#700460000000
0!
0*
09
0>
0C
#700470000000
1!
1*
b1 6
19
1>
1C
b1 G
#700480000000
0!
0*
09
0>
0C
#700490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#700500000000
0!
0*
09
0>
0C
#700510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#700520000000
0!
0*
09
0>
0C
#700530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#700540000000
0!
0*
09
0>
0C
#700550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#700560000000
0!
0#
0*
0,
09
0>
0?
0C
#700570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#700580000000
0!
0*
09
0>
0C
#700590000000
1!
1*
19
1>
1C
#700600000000
0!
0*
09
0>
0C
#700610000000
1!
1*
19
1>
1C
#700620000000
0!
0*
09
0>
0C
#700630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#700640000000
0!
0*
09
0>
0C
#700650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#700660000000
0!
0*
09
0>
0C
#700670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#700680000000
0!
0*
09
0>
0C
#700690000000
1!
1*
b10 6
19
1>
1C
b10 G
#700700000000
0!
0*
09
0>
0C
#700710000000
1!
1*
b11 6
19
1>
1C
b11 G
#700720000000
0!
0*
09
0>
0C
#700730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#700740000000
0!
0*
09
0>
0C
#700750000000
1!
1*
b101 6
19
1>
1C
b101 G
#700760000000
0!
0*
09
0>
0C
#700770000000
1!
1*
b110 6
19
1>
1C
b110 G
#700780000000
0!
0*
09
0>
0C
#700790000000
1!
1*
b111 6
19
1>
1C
b111 G
#700800000000
0!
0*
09
0>
0C
#700810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#700820000000
0!
0*
09
0>
0C
#700830000000
1!
1*
b1 6
19
1>
1C
b1 G
#700840000000
0!
0*
09
0>
0C
#700850000000
1!
1*
b10 6
19
1>
1C
b10 G
#700860000000
0!
0*
09
0>
0C
#700870000000
1!
1*
b11 6
19
1>
1C
b11 G
#700880000000
0!
0*
09
0>
0C
#700890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#700900000000
0!
0*
09
0>
0C
#700910000000
1!
1*
b101 6
19
1>
1C
b101 G
#700920000000
0!
0*
09
0>
0C
#700930000000
1!
1*
b110 6
19
1>
1C
b110 G
#700940000000
0!
0*
09
0>
0C
#700950000000
1!
1*
b111 6
19
1>
1C
b111 G
#700960000000
0!
0*
09
0>
0C
#700970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#700980000000
0!
0*
09
0>
0C
#700990000000
1!
1*
b1 6
19
1>
1C
b1 G
#701000000000
0!
0*
09
0>
0C
#701010000000
1!
1*
b10 6
19
1>
1C
b10 G
#701020000000
0!
0*
09
0>
0C
#701030000000
1!
1*
b11 6
19
1>
1C
b11 G
#701040000000
0!
0*
09
0>
0C
#701050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#701060000000
0!
0*
09
0>
0C
#701070000000
1!
1*
b101 6
19
1>
1C
b101 G
#701080000000
0!
0*
09
0>
0C
#701090000000
1!
1*
b110 6
19
1>
1C
b110 G
#701100000000
0!
0*
09
0>
0C
#701110000000
1!
1*
b111 6
19
1>
1C
b111 G
#701120000000
0!
1"
0*
1+
09
1:
0>
0C
#701130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#701140000000
0!
0*
09
0>
0C
#701150000000
1!
1*
b1 6
19
1>
1C
b1 G
#701160000000
0!
0*
09
0>
0C
#701170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#701180000000
0!
0*
09
0>
0C
#701190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#701200000000
0!
0*
09
0>
0C
#701210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#701220000000
0!
0*
09
0>
0C
#701230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#701240000000
0!
0#
0*
0,
09
0>
0?
0C
#701250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#701260000000
0!
0*
09
0>
0C
#701270000000
1!
1*
19
1>
1C
#701280000000
0!
0*
09
0>
0C
#701290000000
1!
1*
19
1>
1C
#701300000000
0!
0*
09
0>
0C
#701310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#701320000000
0!
0*
09
0>
0C
#701330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#701340000000
0!
0*
09
0>
0C
#701350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#701360000000
0!
0*
09
0>
0C
#701370000000
1!
1*
b10 6
19
1>
1C
b10 G
#701380000000
0!
0*
09
0>
0C
#701390000000
1!
1*
b11 6
19
1>
1C
b11 G
#701400000000
0!
0*
09
0>
0C
#701410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#701420000000
0!
0*
09
0>
0C
#701430000000
1!
1*
b101 6
19
1>
1C
b101 G
#701440000000
0!
0*
09
0>
0C
#701450000000
1!
1*
b110 6
19
1>
1C
b110 G
#701460000000
0!
0*
09
0>
0C
#701470000000
1!
1*
b111 6
19
1>
1C
b111 G
#701480000000
0!
0*
09
0>
0C
#701490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#701500000000
0!
0*
09
0>
0C
#701510000000
1!
1*
b1 6
19
1>
1C
b1 G
#701520000000
0!
0*
09
0>
0C
#701530000000
1!
1*
b10 6
19
1>
1C
b10 G
#701540000000
0!
0*
09
0>
0C
#701550000000
1!
1*
b11 6
19
1>
1C
b11 G
#701560000000
0!
0*
09
0>
0C
#701570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#701580000000
0!
0*
09
0>
0C
#701590000000
1!
1*
b101 6
19
1>
1C
b101 G
#701600000000
0!
0*
09
0>
0C
#701610000000
1!
1*
b110 6
19
1>
1C
b110 G
#701620000000
0!
0*
09
0>
0C
#701630000000
1!
1*
b111 6
19
1>
1C
b111 G
#701640000000
0!
0*
09
0>
0C
#701650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#701660000000
0!
0*
09
0>
0C
#701670000000
1!
1*
b1 6
19
1>
1C
b1 G
#701680000000
0!
0*
09
0>
0C
#701690000000
1!
1*
b10 6
19
1>
1C
b10 G
#701700000000
0!
0*
09
0>
0C
#701710000000
1!
1*
b11 6
19
1>
1C
b11 G
#701720000000
0!
0*
09
0>
0C
#701730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#701740000000
0!
0*
09
0>
0C
#701750000000
1!
1*
b101 6
19
1>
1C
b101 G
#701760000000
0!
0*
09
0>
0C
#701770000000
1!
1*
b110 6
19
1>
1C
b110 G
#701780000000
0!
0*
09
0>
0C
#701790000000
1!
1*
b111 6
19
1>
1C
b111 G
#701800000000
0!
1"
0*
1+
09
1:
0>
0C
#701810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#701820000000
0!
0*
09
0>
0C
#701830000000
1!
1*
b1 6
19
1>
1C
b1 G
#701840000000
0!
0*
09
0>
0C
#701850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#701860000000
0!
0*
09
0>
0C
#701870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#701880000000
0!
0*
09
0>
0C
#701890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#701900000000
0!
0*
09
0>
0C
#701910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#701920000000
0!
0#
0*
0,
09
0>
0?
0C
#701930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#701940000000
0!
0*
09
0>
0C
#701950000000
1!
1*
19
1>
1C
#701960000000
0!
0*
09
0>
0C
#701970000000
1!
1*
19
1>
1C
#701980000000
0!
0*
09
0>
0C
#701990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#702000000000
0!
0*
09
0>
0C
#702010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#702020000000
0!
0*
09
0>
0C
#702030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#702040000000
0!
0*
09
0>
0C
#702050000000
1!
1*
b10 6
19
1>
1C
b10 G
#702060000000
0!
0*
09
0>
0C
#702070000000
1!
1*
b11 6
19
1>
1C
b11 G
#702080000000
0!
0*
09
0>
0C
#702090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#702100000000
0!
0*
09
0>
0C
#702110000000
1!
1*
b101 6
19
1>
1C
b101 G
#702120000000
0!
0*
09
0>
0C
#702130000000
1!
1*
b110 6
19
1>
1C
b110 G
#702140000000
0!
0*
09
0>
0C
#702150000000
1!
1*
b111 6
19
1>
1C
b111 G
#702160000000
0!
0*
09
0>
0C
#702170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#702180000000
0!
0*
09
0>
0C
#702190000000
1!
1*
b1 6
19
1>
1C
b1 G
#702200000000
0!
0*
09
0>
0C
#702210000000
1!
1*
b10 6
19
1>
1C
b10 G
#702220000000
0!
0*
09
0>
0C
#702230000000
1!
1*
b11 6
19
1>
1C
b11 G
#702240000000
0!
0*
09
0>
0C
#702250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#702260000000
0!
0*
09
0>
0C
#702270000000
1!
1*
b101 6
19
1>
1C
b101 G
#702280000000
0!
0*
09
0>
0C
#702290000000
1!
1*
b110 6
19
1>
1C
b110 G
#702300000000
0!
0*
09
0>
0C
#702310000000
1!
1*
b111 6
19
1>
1C
b111 G
#702320000000
0!
0*
09
0>
0C
#702330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#702340000000
0!
0*
09
0>
0C
#702350000000
1!
1*
b1 6
19
1>
1C
b1 G
#702360000000
0!
0*
09
0>
0C
#702370000000
1!
1*
b10 6
19
1>
1C
b10 G
#702380000000
0!
0*
09
0>
0C
#702390000000
1!
1*
b11 6
19
1>
1C
b11 G
#702400000000
0!
0*
09
0>
0C
#702410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#702420000000
0!
0*
09
0>
0C
#702430000000
1!
1*
b101 6
19
1>
1C
b101 G
#702440000000
0!
0*
09
0>
0C
#702450000000
1!
1*
b110 6
19
1>
1C
b110 G
#702460000000
0!
0*
09
0>
0C
#702470000000
1!
1*
b111 6
19
1>
1C
b111 G
#702480000000
0!
1"
0*
1+
09
1:
0>
0C
#702490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#702500000000
0!
0*
09
0>
0C
#702510000000
1!
1*
b1 6
19
1>
1C
b1 G
#702520000000
0!
0*
09
0>
0C
#702530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#702540000000
0!
0*
09
0>
0C
#702550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#702560000000
0!
0*
09
0>
0C
#702570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#702580000000
0!
0*
09
0>
0C
#702590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#702600000000
0!
0#
0*
0,
09
0>
0?
0C
#702610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#702620000000
0!
0*
09
0>
0C
#702630000000
1!
1*
19
1>
1C
#702640000000
0!
0*
09
0>
0C
#702650000000
1!
1*
19
1>
1C
#702660000000
0!
0*
09
0>
0C
#702670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#702680000000
0!
0*
09
0>
0C
#702690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#702700000000
0!
0*
09
0>
0C
#702710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#702720000000
0!
0*
09
0>
0C
#702730000000
1!
1*
b10 6
19
1>
1C
b10 G
#702740000000
0!
0*
09
0>
0C
#702750000000
1!
1*
b11 6
19
1>
1C
b11 G
#702760000000
0!
0*
09
0>
0C
#702770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#702780000000
0!
0*
09
0>
0C
#702790000000
1!
1*
b101 6
19
1>
1C
b101 G
#702800000000
0!
0*
09
0>
0C
#702810000000
1!
1*
b110 6
19
1>
1C
b110 G
#702820000000
0!
0*
09
0>
0C
#702830000000
1!
1*
b111 6
19
1>
1C
b111 G
#702840000000
0!
0*
09
0>
0C
#702850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#702860000000
0!
0*
09
0>
0C
#702870000000
1!
1*
b1 6
19
1>
1C
b1 G
#702880000000
0!
0*
09
0>
0C
#702890000000
1!
1*
b10 6
19
1>
1C
b10 G
#702900000000
0!
0*
09
0>
0C
#702910000000
1!
1*
b11 6
19
1>
1C
b11 G
#702920000000
0!
0*
09
0>
0C
#702930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#702940000000
0!
0*
09
0>
0C
#702950000000
1!
1*
b101 6
19
1>
1C
b101 G
#702960000000
0!
0*
09
0>
0C
#702970000000
1!
1*
b110 6
19
1>
1C
b110 G
#702980000000
0!
0*
09
0>
0C
#702990000000
1!
1*
b111 6
19
1>
1C
b111 G
#703000000000
0!
0*
09
0>
0C
#703010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#703020000000
0!
0*
09
0>
0C
#703030000000
1!
1*
b1 6
19
1>
1C
b1 G
#703040000000
0!
0*
09
0>
0C
#703050000000
1!
1*
b10 6
19
1>
1C
b10 G
#703060000000
0!
0*
09
0>
0C
#703070000000
1!
1*
b11 6
19
1>
1C
b11 G
#703080000000
0!
0*
09
0>
0C
#703090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#703100000000
0!
0*
09
0>
0C
#703110000000
1!
1*
b101 6
19
1>
1C
b101 G
#703120000000
0!
0*
09
0>
0C
#703130000000
1!
1*
b110 6
19
1>
1C
b110 G
#703140000000
0!
0*
09
0>
0C
#703150000000
1!
1*
b111 6
19
1>
1C
b111 G
#703160000000
0!
1"
0*
1+
09
1:
0>
0C
#703170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#703180000000
0!
0*
09
0>
0C
#703190000000
1!
1*
b1 6
19
1>
1C
b1 G
#703200000000
0!
0*
09
0>
0C
#703210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#703220000000
0!
0*
09
0>
0C
#703230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#703240000000
0!
0*
09
0>
0C
#703250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#703260000000
0!
0*
09
0>
0C
#703270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#703280000000
0!
0#
0*
0,
09
0>
0?
0C
#703290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#703300000000
0!
0*
09
0>
0C
#703310000000
1!
1*
19
1>
1C
#703320000000
0!
0*
09
0>
0C
#703330000000
1!
1*
19
1>
1C
#703340000000
0!
0*
09
0>
0C
#703350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#703360000000
0!
0*
09
0>
0C
#703370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#703380000000
0!
0*
09
0>
0C
#703390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#703400000000
0!
0*
09
0>
0C
#703410000000
1!
1*
b10 6
19
1>
1C
b10 G
#703420000000
0!
0*
09
0>
0C
#703430000000
1!
1*
b11 6
19
1>
1C
b11 G
#703440000000
0!
0*
09
0>
0C
#703450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#703460000000
0!
0*
09
0>
0C
#703470000000
1!
1*
b101 6
19
1>
1C
b101 G
#703480000000
0!
0*
09
0>
0C
#703490000000
1!
1*
b110 6
19
1>
1C
b110 G
#703500000000
0!
0*
09
0>
0C
#703510000000
1!
1*
b111 6
19
1>
1C
b111 G
#703520000000
0!
0*
09
0>
0C
#703530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#703540000000
0!
0*
09
0>
0C
#703550000000
1!
1*
b1 6
19
1>
1C
b1 G
#703560000000
0!
0*
09
0>
0C
#703570000000
1!
1*
b10 6
19
1>
1C
b10 G
#703580000000
0!
0*
09
0>
0C
#703590000000
1!
1*
b11 6
19
1>
1C
b11 G
#703600000000
0!
0*
09
0>
0C
#703610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#703620000000
0!
0*
09
0>
0C
#703630000000
1!
1*
b101 6
19
1>
1C
b101 G
#703640000000
0!
0*
09
0>
0C
#703650000000
1!
1*
b110 6
19
1>
1C
b110 G
#703660000000
0!
0*
09
0>
0C
#703670000000
1!
1*
b111 6
19
1>
1C
b111 G
#703680000000
0!
0*
09
0>
0C
#703690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#703700000000
0!
0*
09
0>
0C
#703710000000
1!
1*
b1 6
19
1>
1C
b1 G
#703720000000
0!
0*
09
0>
0C
#703730000000
1!
1*
b10 6
19
1>
1C
b10 G
#703740000000
0!
0*
09
0>
0C
#703750000000
1!
1*
b11 6
19
1>
1C
b11 G
#703760000000
0!
0*
09
0>
0C
#703770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#703780000000
0!
0*
09
0>
0C
#703790000000
1!
1*
b101 6
19
1>
1C
b101 G
#703800000000
0!
0*
09
0>
0C
#703810000000
1!
1*
b110 6
19
1>
1C
b110 G
#703820000000
0!
0*
09
0>
0C
#703830000000
1!
1*
b111 6
19
1>
1C
b111 G
#703840000000
0!
1"
0*
1+
09
1:
0>
0C
#703850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#703860000000
0!
0*
09
0>
0C
#703870000000
1!
1*
b1 6
19
1>
1C
b1 G
#703880000000
0!
0*
09
0>
0C
#703890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#703900000000
0!
0*
09
0>
0C
#703910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#703920000000
0!
0*
09
0>
0C
#703930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#703940000000
0!
0*
09
0>
0C
#703950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#703960000000
0!
0#
0*
0,
09
0>
0?
0C
#703970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#703980000000
0!
0*
09
0>
0C
#703990000000
1!
1*
19
1>
1C
#704000000000
0!
0*
09
0>
0C
#704010000000
1!
1*
19
1>
1C
#704020000000
0!
0*
09
0>
0C
#704030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#704040000000
0!
0*
09
0>
0C
#704050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#704060000000
0!
0*
09
0>
0C
#704070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#704080000000
0!
0*
09
0>
0C
#704090000000
1!
1*
b10 6
19
1>
1C
b10 G
#704100000000
0!
0*
09
0>
0C
#704110000000
1!
1*
b11 6
19
1>
1C
b11 G
#704120000000
0!
0*
09
0>
0C
#704130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#704140000000
0!
0*
09
0>
0C
#704150000000
1!
1*
b101 6
19
1>
1C
b101 G
#704160000000
0!
0*
09
0>
0C
#704170000000
1!
1*
b110 6
19
1>
1C
b110 G
#704180000000
0!
0*
09
0>
0C
#704190000000
1!
1*
b111 6
19
1>
1C
b111 G
#704200000000
0!
0*
09
0>
0C
#704210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#704220000000
0!
0*
09
0>
0C
#704230000000
1!
1*
b1 6
19
1>
1C
b1 G
#704240000000
0!
0*
09
0>
0C
#704250000000
1!
1*
b10 6
19
1>
1C
b10 G
#704260000000
0!
0*
09
0>
0C
#704270000000
1!
1*
b11 6
19
1>
1C
b11 G
#704280000000
0!
0*
09
0>
0C
#704290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#704300000000
0!
0*
09
0>
0C
#704310000000
1!
1*
b101 6
19
1>
1C
b101 G
#704320000000
0!
0*
09
0>
0C
#704330000000
1!
1*
b110 6
19
1>
1C
b110 G
#704340000000
0!
0*
09
0>
0C
#704350000000
1!
1*
b111 6
19
1>
1C
b111 G
#704360000000
0!
0*
09
0>
0C
#704370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#704380000000
0!
0*
09
0>
0C
#704390000000
1!
1*
b1 6
19
1>
1C
b1 G
#704400000000
0!
0*
09
0>
0C
#704410000000
1!
1*
b10 6
19
1>
1C
b10 G
#704420000000
0!
0*
09
0>
0C
#704430000000
1!
1*
b11 6
19
1>
1C
b11 G
#704440000000
0!
0*
09
0>
0C
#704450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#704460000000
0!
0*
09
0>
0C
#704470000000
1!
1*
b101 6
19
1>
1C
b101 G
#704480000000
0!
0*
09
0>
0C
#704490000000
1!
1*
b110 6
19
1>
1C
b110 G
#704500000000
0!
0*
09
0>
0C
#704510000000
1!
1*
b111 6
19
1>
1C
b111 G
#704520000000
0!
1"
0*
1+
09
1:
0>
0C
#704530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#704540000000
0!
0*
09
0>
0C
#704550000000
1!
1*
b1 6
19
1>
1C
b1 G
#704560000000
0!
0*
09
0>
0C
#704570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#704580000000
0!
0*
09
0>
0C
#704590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#704600000000
0!
0*
09
0>
0C
#704610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#704620000000
0!
0*
09
0>
0C
#704630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#704640000000
0!
0#
0*
0,
09
0>
0?
0C
#704650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#704660000000
0!
0*
09
0>
0C
#704670000000
1!
1*
19
1>
1C
#704680000000
0!
0*
09
0>
0C
#704690000000
1!
1*
19
1>
1C
#704700000000
0!
0*
09
0>
0C
#704710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#704720000000
0!
0*
09
0>
0C
#704730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#704740000000
0!
0*
09
0>
0C
#704750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#704760000000
0!
0*
09
0>
0C
#704770000000
1!
1*
b10 6
19
1>
1C
b10 G
#704780000000
0!
0*
09
0>
0C
#704790000000
1!
1*
b11 6
19
1>
1C
b11 G
#704800000000
0!
0*
09
0>
0C
#704810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#704820000000
0!
0*
09
0>
0C
#704830000000
1!
1*
b101 6
19
1>
1C
b101 G
#704840000000
0!
0*
09
0>
0C
#704850000000
1!
1*
b110 6
19
1>
1C
b110 G
#704860000000
0!
0*
09
0>
0C
#704870000000
1!
1*
b111 6
19
1>
1C
b111 G
#704880000000
0!
0*
09
0>
0C
#704890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#704900000000
0!
0*
09
0>
0C
#704910000000
1!
1*
b1 6
19
1>
1C
b1 G
#704920000000
0!
0*
09
0>
0C
#704930000000
1!
1*
b10 6
19
1>
1C
b10 G
#704940000000
0!
0*
09
0>
0C
#704950000000
1!
1*
b11 6
19
1>
1C
b11 G
#704960000000
0!
0*
09
0>
0C
#704970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#704980000000
0!
0*
09
0>
0C
#704990000000
1!
1*
b101 6
19
1>
1C
b101 G
#705000000000
0!
0*
09
0>
0C
#705010000000
1!
1*
b110 6
19
1>
1C
b110 G
#705020000000
0!
0*
09
0>
0C
#705030000000
1!
1*
b111 6
19
1>
1C
b111 G
#705040000000
0!
0*
09
0>
0C
#705050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#705060000000
0!
0*
09
0>
0C
#705070000000
1!
1*
b1 6
19
1>
1C
b1 G
#705080000000
0!
0*
09
0>
0C
#705090000000
1!
1*
b10 6
19
1>
1C
b10 G
#705100000000
0!
0*
09
0>
0C
#705110000000
1!
1*
b11 6
19
1>
1C
b11 G
#705120000000
0!
0*
09
0>
0C
#705130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#705140000000
0!
0*
09
0>
0C
#705150000000
1!
1*
b101 6
19
1>
1C
b101 G
#705160000000
0!
0*
09
0>
0C
#705170000000
1!
1*
b110 6
19
1>
1C
b110 G
#705180000000
0!
0*
09
0>
0C
#705190000000
1!
1*
b111 6
19
1>
1C
b111 G
#705200000000
0!
1"
0*
1+
09
1:
0>
0C
#705210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#705220000000
0!
0*
09
0>
0C
#705230000000
1!
1*
b1 6
19
1>
1C
b1 G
#705240000000
0!
0*
09
0>
0C
#705250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#705260000000
0!
0*
09
0>
0C
#705270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#705280000000
0!
0*
09
0>
0C
#705290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#705300000000
0!
0*
09
0>
0C
#705310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#705320000000
0!
0#
0*
0,
09
0>
0?
0C
#705330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#705340000000
0!
0*
09
0>
0C
#705350000000
1!
1*
19
1>
1C
#705360000000
0!
0*
09
0>
0C
#705370000000
1!
1*
19
1>
1C
#705380000000
0!
0*
09
0>
0C
#705390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#705400000000
0!
0*
09
0>
0C
#705410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#705420000000
0!
0*
09
0>
0C
#705430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#705440000000
0!
0*
09
0>
0C
#705450000000
1!
1*
b10 6
19
1>
1C
b10 G
#705460000000
0!
0*
09
0>
0C
#705470000000
1!
1*
b11 6
19
1>
1C
b11 G
#705480000000
0!
0*
09
0>
0C
#705490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#705500000000
0!
0*
09
0>
0C
#705510000000
1!
1*
b101 6
19
1>
1C
b101 G
#705520000000
0!
0*
09
0>
0C
#705530000000
1!
1*
b110 6
19
1>
1C
b110 G
#705540000000
0!
0*
09
0>
0C
#705550000000
1!
1*
b111 6
19
1>
1C
b111 G
#705560000000
0!
0*
09
0>
0C
#705570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#705580000000
0!
0*
09
0>
0C
#705590000000
1!
1*
b1 6
19
1>
1C
b1 G
#705600000000
0!
0*
09
0>
0C
#705610000000
1!
1*
b10 6
19
1>
1C
b10 G
#705620000000
0!
0*
09
0>
0C
#705630000000
1!
1*
b11 6
19
1>
1C
b11 G
#705640000000
0!
0*
09
0>
0C
#705650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#705660000000
0!
0*
09
0>
0C
#705670000000
1!
1*
b101 6
19
1>
1C
b101 G
#705680000000
0!
0*
09
0>
0C
#705690000000
1!
1*
b110 6
19
1>
1C
b110 G
#705700000000
0!
0*
09
0>
0C
#705710000000
1!
1*
b111 6
19
1>
1C
b111 G
#705720000000
0!
0*
09
0>
0C
#705730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#705740000000
0!
0*
09
0>
0C
#705750000000
1!
1*
b1 6
19
1>
1C
b1 G
#705760000000
0!
0*
09
0>
0C
#705770000000
1!
1*
b10 6
19
1>
1C
b10 G
#705780000000
0!
0*
09
0>
0C
#705790000000
1!
1*
b11 6
19
1>
1C
b11 G
#705800000000
0!
0*
09
0>
0C
#705810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#705820000000
0!
0*
09
0>
0C
#705830000000
1!
1*
b101 6
19
1>
1C
b101 G
#705840000000
0!
0*
09
0>
0C
#705850000000
1!
1*
b110 6
19
1>
1C
b110 G
#705860000000
0!
0*
09
0>
0C
#705870000000
1!
1*
b111 6
19
1>
1C
b111 G
#705880000000
0!
1"
0*
1+
09
1:
0>
0C
#705890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#705900000000
0!
0*
09
0>
0C
#705910000000
1!
1*
b1 6
19
1>
1C
b1 G
#705920000000
0!
0*
09
0>
0C
#705930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#705940000000
0!
0*
09
0>
0C
#705950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#705960000000
0!
0*
09
0>
0C
#705970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#705980000000
0!
0*
09
0>
0C
#705990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#706000000000
0!
0#
0*
0,
09
0>
0?
0C
#706010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#706020000000
0!
0*
09
0>
0C
#706030000000
1!
1*
19
1>
1C
#706040000000
0!
0*
09
0>
0C
#706050000000
1!
1*
19
1>
1C
#706060000000
0!
0*
09
0>
0C
#706070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#706080000000
0!
0*
09
0>
0C
#706090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#706100000000
0!
0*
09
0>
0C
#706110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#706120000000
0!
0*
09
0>
0C
#706130000000
1!
1*
b10 6
19
1>
1C
b10 G
#706140000000
0!
0*
09
0>
0C
#706150000000
1!
1*
b11 6
19
1>
1C
b11 G
#706160000000
0!
0*
09
0>
0C
#706170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#706180000000
0!
0*
09
0>
0C
#706190000000
1!
1*
b101 6
19
1>
1C
b101 G
#706200000000
0!
0*
09
0>
0C
#706210000000
1!
1*
b110 6
19
1>
1C
b110 G
#706220000000
0!
0*
09
0>
0C
#706230000000
1!
1*
b111 6
19
1>
1C
b111 G
#706240000000
0!
0*
09
0>
0C
#706250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#706260000000
0!
0*
09
0>
0C
#706270000000
1!
1*
b1 6
19
1>
1C
b1 G
#706280000000
0!
0*
09
0>
0C
#706290000000
1!
1*
b10 6
19
1>
1C
b10 G
#706300000000
0!
0*
09
0>
0C
#706310000000
1!
1*
b11 6
19
1>
1C
b11 G
#706320000000
0!
0*
09
0>
0C
#706330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#706340000000
0!
0*
09
0>
0C
#706350000000
1!
1*
b101 6
19
1>
1C
b101 G
#706360000000
0!
0*
09
0>
0C
#706370000000
1!
1*
b110 6
19
1>
1C
b110 G
#706380000000
0!
0*
09
0>
0C
#706390000000
1!
1*
b111 6
19
1>
1C
b111 G
#706400000000
0!
0*
09
0>
0C
#706410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#706420000000
0!
0*
09
0>
0C
#706430000000
1!
1*
b1 6
19
1>
1C
b1 G
#706440000000
0!
0*
09
0>
0C
#706450000000
1!
1*
b10 6
19
1>
1C
b10 G
#706460000000
0!
0*
09
0>
0C
#706470000000
1!
1*
b11 6
19
1>
1C
b11 G
#706480000000
0!
0*
09
0>
0C
#706490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#706500000000
0!
0*
09
0>
0C
#706510000000
1!
1*
b101 6
19
1>
1C
b101 G
#706520000000
0!
0*
09
0>
0C
#706530000000
1!
1*
b110 6
19
1>
1C
b110 G
#706540000000
0!
0*
09
0>
0C
#706550000000
1!
1*
b111 6
19
1>
1C
b111 G
#706560000000
0!
1"
0*
1+
09
1:
0>
0C
#706570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#706580000000
0!
0*
09
0>
0C
#706590000000
1!
1*
b1 6
19
1>
1C
b1 G
#706600000000
0!
0*
09
0>
0C
#706610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#706620000000
0!
0*
09
0>
0C
#706630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#706640000000
0!
0*
09
0>
0C
#706650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#706660000000
0!
0*
09
0>
0C
#706670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#706680000000
0!
0#
0*
0,
09
0>
0?
0C
#706690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#706700000000
0!
0*
09
0>
0C
#706710000000
1!
1*
19
1>
1C
#706720000000
0!
0*
09
0>
0C
#706730000000
1!
1*
19
1>
1C
#706740000000
0!
0*
09
0>
0C
#706750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#706760000000
0!
0*
09
0>
0C
#706770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#706780000000
0!
0*
09
0>
0C
#706790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#706800000000
0!
0*
09
0>
0C
#706810000000
1!
1*
b10 6
19
1>
1C
b10 G
#706820000000
0!
0*
09
0>
0C
#706830000000
1!
1*
b11 6
19
1>
1C
b11 G
#706840000000
0!
0*
09
0>
0C
#706850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#706860000000
0!
0*
09
0>
0C
#706870000000
1!
1*
b101 6
19
1>
1C
b101 G
#706880000000
0!
0*
09
0>
0C
#706890000000
1!
1*
b110 6
19
1>
1C
b110 G
#706900000000
0!
0*
09
0>
0C
#706910000000
1!
1*
b111 6
19
1>
1C
b111 G
#706920000000
0!
0*
09
0>
0C
#706930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#706940000000
0!
0*
09
0>
0C
#706950000000
1!
1*
b1 6
19
1>
1C
b1 G
#706960000000
0!
0*
09
0>
0C
#706970000000
1!
1*
b10 6
19
1>
1C
b10 G
#706980000000
0!
0*
09
0>
0C
#706990000000
1!
1*
b11 6
19
1>
1C
b11 G
#707000000000
0!
0*
09
0>
0C
#707010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#707020000000
0!
0*
09
0>
0C
#707030000000
1!
1*
b101 6
19
1>
1C
b101 G
#707040000000
0!
0*
09
0>
0C
#707050000000
1!
1*
b110 6
19
1>
1C
b110 G
#707060000000
0!
0*
09
0>
0C
#707070000000
1!
1*
b111 6
19
1>
1C
b111 G
#707080000000
0!
0*
09
0>
0C
#707090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#707100000000
0!
0*
09
0>
0C
#707110000000
1!
1*
b1 6
19
1>
1C
b1 G
#707120000000
0!
0*
09
0>
0C
#707130000000
1!
1*
b10 6
19
1>
1C
b10 G
#707140000000
0!
0*
09
0>
0C
#707150000000
1!
1*
b11 6
19
1>
1C
b11 G
#707160000000
0!
0*
09
0>
0C
#707170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#707180000000
0!
0*
09
0>
0C
#707190000000
1!
1*
b101 6
19
1>
1C
b101 G
#707200000000
0!
0*
09
0>
0C
#707210000000
1!
1*
b110 6
19
1>
1C
b110 G
#707220000000
0!
0*
09
0>
0C
#707230000000
1!
1*
b111 6
19
1>
1C
b111 G
#707240000000
0!
1"
0*
1+
09
1:
0>
0C
#707250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#707260000000
0!
0*
09
0>
0C
#707270000000
1!
1*
b1 6
19
1>
1C
b1 G
#707280000000
0!
0*
09
0>
0C
#707290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#707300000000
0!
0*
09
0>
0C
#707310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#707320000000
0!
0*
09
0>
0C
#707330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#707340000000
0!
0*
09
0>
0C
#707350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#707360000000
0!
0#
0*
0,
09
0>
0?
0C
#707370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#707380000000
0!
0*
09
0>
0C
#707390000000
1!
1*
19
1>
1C
#707400000000
0!
0*
09
0>
0C
#707410000000
1!
1*
19
1>
1C
#707420000000
0!
0*
09
0>
0C
#707430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#707440000000
0!
0*
09
0>
0C
#707450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#707460000000
0!
0*
09
0>
0C
#707470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#707480000000
0!
0*
09
0>
0C
#707490000000
1!
1*
b10 6
19
1>
1C
b10 G
#707500000000
0!
0*
09
0>
0C
#707510000000
1!
1*
b11 6
19
1>
1C
b11 G
#707520000000
0!
0*
09
0>
0C
#707530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#707540000000
0!
0*
09
0>
0C
#707550000000
1!
1*
b101 6
19
1>
1C
b101 G
#707560000000
0!
0*
09
0>
0C
#707570000000
1!
1*
b110 6
19
1>
1C
b110 G
#707580000000
0!
0*
09
0>
0C
#707590000000
1!
1*
b111 6
19
1>
1C
b111 G
#707600000000
0!
0*
09
0>
0C
#707610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#707620000000
0!
0*
09
0>
0C
#707630000000
1!
1*
b1 6
19
1>
1C
b1 G
#707640000000
0!
0*
09
0>
0C
#707650000000
1!
1*
b10 6
19
1>
1C
b10 G
#707660000000
0!
0*
09
0>
0C
#707670000000
1!
1*
b11 6
19
1>
1C
b11 G
#707680000000
0!
0*
09
0>
0C
#707690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#707700000000
0!
0*
09
0>
0C
#707710000000
1!
1*
b101 6
19
1>
1C
b101 G
#707720000000
0!
0*
09
0>
0C
#707730000000
1!
1*
b110 6
19
1>
1C
b110 G
#707740000000
0!
0*
09
0>
0C
#707750000000
1!
1*
b111 6
19
1>
1C
b111 G
#707760000000
0!
0*
09
0>
0C
#707770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#707780000000
0!
0*
09
0>
0C
#707790000000
1!
1*
b1 6
19
1>
1C
b1 G
#707800000000
0!
0*
09
0>
0C
#707810000000
1!
1*
b10 6
19
1>
1C
b10 G
#707820000000
0!
0*
09
0>
0C
#707830000000
1!
1*
b11 6
19
1>
1C
b11 G
#707840000000
0!
0*
09
0>
0C
#707850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#707860000000
0!
0*
09
0>
0C
#707870000000
1!
1*
b101 6
19
1>
1C
b101 G
#707880000000
0!
0*
09
0>
0C
#707890000000
1!
1*
b110 6
19
1>
1C
b110 G
#707900000000
0!
0*
09
0>
0C
#707910000000
1!
1*
b111 6
19
1>
1C
b111 G
#707920000000
0!
1"
0*
1+
09
1:
0>
0C
#707930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#707940000000
0!
0*
09
0>
0C
#707950000000
1!
1*
b1 6
19
1>
1C
b1 G
#707960000000
0!
0*
09
0>
0C
#707970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#707980000000
0!
0*
09
0>
0C
#707990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#708000000000
0!
0*
09
0>
0C
#708010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#708020000000
0!
0*
09
0>
0C
#708030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#708040000000
0!
0#
0*
0,
09
0>
0?
0C
#708050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#708060000000
0!
0*
09
0>
0C
#708070000000
1!
1*
19
1>
1C
#708080000000
0!
0*
09
0>
0C
#708090000000
1!
1*
19
1>
1C
#708100000000
0!
0*
09
0>
0C
#708110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#708120000000
0!
0*
09
0>
0C
#708130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#708140000000
0!
0*
09
0>
0C
#708150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#708160000000
0!
0*
09
0>
0C
#708170000000
1!
1*
b10 6
19
1>
1C
b10 G
#708180000000
0!
0*
09
0>
0C
#708190000000
1!
1*
b11 6
19
1>
1C
b11 G
#708200000000
0!
0*
09
0>
0C
#708210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#708220000000
0!
0*
09
0>
0C
#708230000000
1!
1*
b101 6
19
1>
1C
b101 G
#708240000000
0!
0*
09
0>
0C
#708250000000
1!
1*
b110 6
19
1>
1C
b110 G
#708260000000
0!
0*
09
0>
0C
#708270000000
1!
1*
b111 6
19
1>
1C
b111 G
#708280000000
0!
0*
09
0>
0C
#708290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#708300000000
0!
0*
09
0>
0C
#708310000000
1!
1*
b1 6
19
1>
1C
b1 G
#708320000000
0!
0*
09
0>
0C
#708330000000
1!
1*
b10 6
19
1>
1C
b10 G
#708340000000
0!
0*
09
0>
0C
#708350000000
1!
1*
b11 6
19
1>
1C
b11 G
#708360000000
0!
0*
09
0>
0C
#708370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#708380000000
0!
0*
09
0>
0C
#708390000000
1!
1*
b101 6
19
1>
1C
b101 G
#708400000000
0!
0*
09
0>
0C
#708410000000
1!
1*
b110 6
19
1>
1C
b110 G
#708420000000
0!
0*
09
0>
0C
#708430000000
1!
1*
b111 6
19
1>
1C
b111 G
#708440000000
0!
0*
09
0>
0C
#708450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#708460000000
0!
0*
09
0>
0C
#708470000000
1!
1*
b1 6
19
1>
1C
b1 G
#708480000000
0!
0*
09
0>
0C
#708490000000
1!
1*
b10 6
19
1>
1C
b10 G
#708500000000
0!
0*
09
0>
0C
#708510000000
1!
1*
b11 6
19
1>
1C
b11 G
#708520000000
0!
0*
09
0>
0C
#708530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#708540000000
0!
0*
09
0>
0C
#708550000000
1!
1*
b101 6
19
1>
1C
b101 G
#708560000000
0!
0*
09
0>
0C
#708570000000
1!
1*
b110 6
19
1>
1C
b110 G
#708580000000
0!
0*
09
0>
0C
#708590000000
1!
1*
b111 6
19
1>
1C
b111 G
#708600000000
0!
1"
0*
1+
09
1:
0>
0C
#708610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#708620000000
0!
0*
09
0>
0C
#708630000000
1!
1*
b1 6
19
1>
1C
b1 G
#708640000000
0!
0*
09
0>
0C
#708650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#708660000000
0!
0*
09
0>
0C
#708670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#708680000000
0!
0*
09
0>
0C
#708690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#708700000000
0!
0*
09
0>
0C
#708710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#708720000000
0!
0#
0*
0,
09
0>
0?
0C
#708730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#708740000000
0!
0*
09
0>
0C
#708750000000
1!
1*
19
1>
1C
#708760000000
0!
0*
09
0>
0C
#708770000000
1!
1*
19
1>
1C
#708780000000
0!
0*
09
0>
0C
#708790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#708800000000
0!
0*
09
0>
0C
#708810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#708820000000
0!
0*
09
0>
0C
#708830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#708840000000
0!
0*
09
0>
0C
#708850000000
1!
1*
b10 6
19
1>
1C
b10 G
#708860000000
0!
0*
09
0>
0C
#708870000000
1!
1*
b11 6
19
1>
1C
b11 G
#708880000000
0!
0*
09
0>
0C
#708890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#708900000000
0!
0*
09
0>
0C
#708910000000
1!
1*
b101 6
19
1>
1C
b101 G
#708920000000
0!
0*
09
0>
0C
#708930000000
1!
1*
b110 6
19
1>
1C
b110 G
#708940000000
0!
0*
09
0>
0C
#708950000000
1!
1*
b111 6
19
1>
1C
b111 G
#708960000000
0!
0*
09
0>
0C
#708970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#708980000000
0!
0*
09
0>
0C
#708990000000
1!
1*
b1 6
19
1>
1C
b1 G
#709000000000
0!
0*
09
0>
0C
#709010000000
1!
1*
b10 6
19
1>
1C
b10 G
#709020000000
0!
0*
09
0>
0C
#709030000000
1!
1*
b11 6
19
1>
1C
b11 G
#709040000000
0!
0*
09
0>
0C
#709050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#709060000000
0!
0*
09
0>
0C
#709070000000
1!
1*
b101 6
19
1>
1C
b101 G
#709080000000
0!
0*
09
0>
0C
#709090000000
1!
1*
b110 6
19
1>
1C
b110 G
#709100000000
0!
0*
09
0>
0C
#709110000000
1!
1*
b111 6
19
1>
1C
b111 G
#709120000000
0!
0*
09
0>
0C
#709130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#709140000000
0!
0*
09
0>
0C
#709150000000
1!
1*
b1 6
19
1>
1C
b1 G
#709160000000
0!
0*
09
0>
0C
#709170000000
1!
1*
b10 6
19
1>
1C
b10 G
#709180000000
0!
0*
09
0>
0C
#709190000000
1!
1*
b11 6
19
1>
1C
b11 G
#709200000000
0!
0*
09
0>
0C
#709210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#709220000000
0!
0*
09
0>
0C
#709230000000
1!
1*
b101 6
19
1>
1C
b101 G
#709240000000
0!
0*
09
0>
0C
#709250000000
1!
1*
b110 6
19
1>
1C
b110 G
#709260000000
0!
0*
09
0>
0C
#709270000000
1!
1*
b111 6
19
1>
1C
b111 G
#709280000000
0!
1"
0*
1+
09
1:
0>
0C
#709290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#709300000000
0!
0*
09
0>
0C
#709310000000
1!
1*
b1 6
19
1>
1C
b1 G
#709320000000
0!
0*
09
0>
0C
#709330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#709340000000
0!
0*
09
0>
0C
#709350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#709360000000
0!
0*
09
0>
0C
#709370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#709380000000
0!
0*
09
0>
0C
#709390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#709400000000
0!
0#
0*
0,
09
0>
0?
0C
#709410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#709420000000
0!
0*
09
0>
0C
#709430000000
1!
1*
19
1>
1C
#709440000000
0!
0*
09
0>
0C
#709450000000
1!
1*
19
1>
1C
#709460000000
0!
0*
09
0>
0C
#709470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#709480000000
0!
0*
09
0>
0C
#709490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#709500000000
0!
0*
09
0>
0C
#709510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#709520000000
0!
0*
09
0>
0C
#709530000000
1!
1*
b10 6
19
1>
1C
b10 G
#709540000000
0!
0*
09
0>
0C
#709550000000
1!
1*
b11 6
19
1>
1C
b11 G
#709560000000
0!
0*
09
0>
0C
#709570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#709580000000
0!
0*
09
0>
0C
#709590000000
1!
1*
b101 6
19
1>
1C
b101 G
#709600000000
0!
0*
09
0>
0C
#709610000000
1!
1*
b110 6
19
1>
1C
b110 G
#709620000000
0!
0*
09
0>
0C
#709630000000
1!
1*
b111 6
19
1>
1C
b111 G
#709640000000
0!
0*
09
0>
0C
#709650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#709660000000
0!
0*
09
0>
0C
#709670000000
1!
1*
b1 6
19
1>
1C
b1 G
#709680000000
0!
0*
09
0>
0C
#709690000000
1!
1*
b10 6
19
1>
1C
b10 G
#709700000000
0!
0*
09
0>
0C
#709710000000
1!
1*
b11 6
19
1>
1C
b11 G
#709720000000
0!
0*
09
0>
0C
#709730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#709740000000
0!
0*
09
0>
0C
#709750000000
1!
1*
b101 6
19
1>
1C
b101 G
#709760000000
0!
0*
09
0>
0C
#709770000000
1!
1*
b110 6
19
1>
1C
b110 G
#709780000000
0!
0*
09
0>
0C
#709790000000
1!
1*
b111 6
19
1>
1C
b111 G
#709800000000
0!
0*
09
0>
0C
#709810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#709820000000
0!
0*
09
0>
0C
#709830000000
1!
1*
b1 6
19
1>
1C
b1 G
#709840000000
0!
0*
09
0>
0C
#709850000000
1!
1*
b10 6
19
1>
1C
b10 G
#709860000000
0!
0*
09
0>
0C
#709870000000
1!
1*
b11 6
19
1>
1C
b11 G
#709880000000
0!
0*
09
0>
0C
#709890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#709900000000
0!
0*
09
0>
0C
#709910000000
1!
1*
b101 6
19
1>
1C
b101 G
#709920000000
0!
0*
09
0>
0C
#709930000000
1!
1*
b110 6
19
1>
1C
b110 G
#709940000000
0!
0*
09
0>
0C
#709950000000
1!
1*
b111 6
19
1>
1C
b111 G
#709960000000
0!
1"
0*
1+
09
1:
0>
0C
#709970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#709980000000
0!
0*
09
0>
0C
#709990000000
1!
1*
b1 6
19
1>
1C
b1 G
#710000000000
0!
0*
09
0>
0C
#710010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#710020000000
0!
0*
09
0>
0C
#710030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#710040000000
0!
0*
09
0>
0C
#710050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#710060000000
0!
0*
09
0>
0C
#710070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#710080000000
0!
0#
0*
0,
09
0>
0?
0C
#710090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#710100000000
0!
0*
09
0>
0C
#710110000000
1!
1*
19
1>
1C
#710120000000
0!
0*
09
0>
0C
#710130000000
1!
1*
19
1>
1C
#710140000000
0!
0*
09
0>
0C
#710150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#710160000000
0!
0*
09
0>
0C
#710170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#710180000000
0!
0*
09
0>
0C
#710190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#710200000000
0!
0*
09
0>
0C
#710210000000
1!
1*
b10 6
19
1>
1C
b10 G
#710220000000
0!
0*
09
0>
0C
#710230000000
1!
1*
b11 6
19
1>
1C
b11 G
#710240000000
0!
0*
09
0>
0C
#710250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#710260000000
0!
0*
09
0>
0C
#710270000000
1!
1*
b101 6
19
1>
1C
b101 G
#710280000000
0!
0*
09
0>
0C
#710290000000
1!
1*
b110 6
19
1>
1C
b110 G
#710300000000
0!
0*
09
0>
0C
#710310000000
1!
1*
b111 6
19
1>
1C
b111 G
#710320000000
0!
0*
09
0>
0C
#710330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#710340000000
0!
0*
09
0>
0C
#710350000000
1!
1*
b1 6
19
1>
1C
b1 G
#710360000000
0!
0*
09
0>
0C
#710370000000
1!
1*
b10 6
19
1>
1C
b10 G
#710380000000
0!
0*
09
0>
0C
#710390000000
1!
1*
b11 6
19
1>
1C
b11 G
#710400000000
0!
0*
09
0>
0C
#710410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#710420000000
0!
0*
09
0>
0C
#710430000000
1!
1*
b101 6
19
1>
1C
b101 G
#710440000000
0!
0*
09
0>
0C
#710450000000
1!
1*
b110 6
19
1>
1C
b110 G
#710460000000
0!
0*
09
0>
0C
#710470000000
1!
1*
b111 6
19
1>
1C
b111 G
#710480000000
0!
0*
09
0>
0C
#710490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#710500000000
0!
0*
09
0>
0C
#710510000000
1!
1*
b1 6
19
1>
1C
b1 G
#710520000000
0!
0*
09
0>
0C
#710530000000
1!
1*
b10 6
19
1>
1C
b10 G
#710540000000
0!
0*
09
0>
0C
#710550000000
1!
1*
b11 6
19
1>
1C
b11 G
#710560000000
0!
0*
09
0>
0C
#710570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#710580000000
0!
0*
09
0>
0C
#710590000000
1!
1*
b101 6
19
1>
1C
b101 G
#710600000000
0!
0*
09
0>
0C
#710610000000
1!
1*
b110 6
19
1>
1C
b110 G
#710620000000
0!
0*
09
0>
0C
#710630000000
1!
1*
b111 6
19
1>
1C
b111 G
#710640000000
0!
1"
0*
1+
09
1:
0>
0C
#710650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#710660000000
0!
0*
09
0>
0C
#710670000000
1!
1*
b1 6
19
1>
1C
b1 G
#710680000000
0!
0*
09
0>
0C
#710690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#710700000000
0!
0*
09
0>
0C
#710710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#710720000000
0!
0*
09
0>
0C
#710730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#710740000000
0!
0*
09
0>
0C
#710750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#710760000000
0!
0#
0*
0,
09
0>
0?
0C
#710770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#710780000000
0!
0*
09
0>
0C
#710790000000
1!
1*
19
1>
1C
#710800000000
0!
0*
09
0>
0C
#710810000000
1!
1*
19
1>
1C
#710820000000
0!
0*
09
0>
0C
#710830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#710840000000
0!
0*
09
0>
0C
#710850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#710860000000
0!
0*
09
0>
0C
#710870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#710880000000
0!
0*
09
0>
0C
#710890000000
1!
1*
b10 6
19
1>
1C
b10 G
#710900000000
0!
0*
09
0>
0C
#710910000000
1!
1*
b11 6
19
1>
1C
b11 G
#710920000000
0!
0*
09
0>
0C
#710930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#710940000000
0!
0*
09
0>
0C
#710950000000
1!
1*
b101 6
19
1>
1C
b101 G
#710960000000
0!
0*
09
0>
0C
#710970000000
1!
1*
b110 6
19
1>
1C
b110 G
#710980000000
0!
0*
09
0>
0C
#710990000000
1!
1*
b111 6
19
1>
1C
b111 G
#711000000000
0!
0*
09
0>
0C
#711010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#711020000000
0!
0*
09
0>
0C
#711030000000
1!
1*
b1 6
19
1>
1C
b1 G
#711040000000
0!
0*
09
0>
0C
#711050000000
1!
1*
b10 6
19
1>
1C
b10 G
#711060000000
0!
0*
09
0>
0C
#711070000000
1!
1*
b11 6
19
1>
1C
b11 G
#711080000000
0!
0*
09
0>
0C
#711090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#711100000000
0!
0*
09
0>
0C
#711110000000
1!
1*
b101 6
19
1>
1C
b101 G
#711120000000
0!
0*
09
0>
0C
#711130000000
1!
1*
b110 6
19
1>
1C
b110 G
#711140000000
0!
0*
09
0>
0C
#711150000000
1!
1*
b111 6
19
1>
1C
b111 G
#711160000000
0!
0*
09
0>
0C
#711170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#711180000000
0!
0*
09
0>
0C
#711190000000
1!
1*
b1 6
19
1>
1C
b1 G
#711200000000
0!
0*
09
0>
0C
#711210000000
1!
1*
b10 6
19
1>
1C
b10 G
#711220000000
0!
0*
09
0>
0C
#711230000000
1!
1*
b11 6
19
1>
1C
b11 G
#711240000000
0!
0*
09
0>
0C
#711250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#711260000000
0!
0*
09
0>
0C
#711270000000
1!
1*
b101 6
19
1>
1C
b101 G
#711280000000
0!
0*
09
0>
0C
#711290000000
1!
1*
b110 6
19
1>
1C
b110 G
#711300000000
0!
0*
09
0>
0C
#711310000000
1!
1*
b111 6
19
1>
1C
b111 G
#711320000000
0!
1"
0*
1+
09
1:
0>
0C
#711330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#711340000000
0!
0*
09
0>
0C
#711350000000
1!
1*
b1 6
19
1>
1C
b1 G
#711360000000
0!
0*
09
0>
0C
#711370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#711380000000
0!
0*
09
0>
0C
#711390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#711400000000
0!
0*
09
0>
0C
#711410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#711420000000
0!
0*
09
0>
0C
#711430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#711440000000
0!
0#
0*
0,
09
0>
0?
0C
#711450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#711460000000
0!
0*
09
0>
0C
#711470000000
1!
1*
19
1>
1C
#711480000000
0!
0*
09
0>
0C
#711490000000
1!
1*
19
1>
1C
#711500000000
0!
0*
09
0>
0C
#711510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#711520000000
0!
0*
09
0>
0C
#711530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#711540000000
0!
0*
09
0>
0C
#711550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#711560000000
0!
0*
09
0>
0C
#711570000000
1!
1*
b10 6
19
1>
1C
b10 G
#711580000000
0!
0*
09
0>
0C
#711590000000
1!
1*
b11 6
19
1>
1C
b11 G
#711600000000
0!
0*
09
0>
0C
#711610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#711620000000
0!
0*
09
0>
0C
#711630000000
1!
1*
b101 6
19
1>
1C
b101 G
#711640000000
0!
0*
09
0>
0C
#711650000000
1!
1*
b110 6
19
1>
1C
b110 G
#711660000000
0!
0*
09
0>
0C
#711670000000
1!
1*
b111 6
19
1>
1C
b111 G
#711680000000
0!
0*
09
0>
0C
#711690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#711700000000
0!
0*
09
0>
0C
#711710000000
1!
1*
b1 6
19
1>
1C
b1 G
#711720000000
0!
0*
09
0>
0C
#711730000000
1!
1*
b10 6
19
1>
1C
b10 G
#711740000000
0!
0*
09
0>
0C
#711750000000
1!
1*
b11 6
19
1>
1C
b11 G
#711760000000
0!
0*
09
0>
0C
#711770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#711780000000
0!
0*
09
0>
0C
#711790000000
1!
1*
b101 6
19
1>
1C
b101 G
#711800000000
0!
0*
09
0>
0C
#711810000000
1!
1*
b110 6
19
1>
1C
b110 G
#711820000000
0!
0*
09
0>
0C
#711830000000
1!
1*
b111 6
19
1>
1C
b111 G
#711840000000
0!
0*
09
0>
0C
#711850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#711860000000
0!
0*
09
0>
0C
#711870000000
1!
1*
b1 6
19
1>
1C
b1 G
#711880000000
0!
0*
09
0>
0C
#711890000000
1!
1*
b10 6
19
1>
1C
b10 G
#711900000000
0!
0*
09
0>
0C
#711910000000
1!
1*
b11 6
19
1>
1C
b11 G
#711920000000
0!
0*
09
0>
0C
#711930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#711940000000
0!
0*
09
0>
0C
#711950000000
1!
1*
b101 6
19
1>
1C
b101 G
#711960000000
0!
0*
09
0>
0C
#711970000000
1!
1*
b110 6
19
1>
1C
b110 G
#711980000000
0!
0*
09
0>
0C
#711990000000
1!
1*
b111 6
19
1>
1C
b111 G
#712000000000
0!
1"
0*
1+
09
1:
0>
0C
#712010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#712020000000
0!
0*
09
0>
0C
#712030000000
1!
1*
b1 6
19
1>
1C
b1 G
#712040000000
0!
0*
09
0>
0C
#712050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#712060000000
0!
0*
09
0>
0C
#712070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#712080000000
0!
0*
09
0>
0C
#712090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#712100000000
0!
0*
09
0>
0C
#712110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#712120000000
0!
0#
0*
0,
09
0>
0?
0C
#712130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#712140000000
0!
0*
09
0>
0C
#712150000000
1!
1*
19
1>
1C
#712160000000
0!
0*
09
0>
0C
#712170000000
1!
1*
19
1>
1C
#712180000000
0!
0*
09
0>
0C
#712190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#712200000000
0!
0*
09
0>
0C
#712210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#712220000000
0!
0*
09
0>
0C
#712230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#712240000000
0!
0*
09
0>
0C
#712250000000
1!
1*
b10 6
19
1>
1C
b10 G
#712260000000
0!
0*
09
0>
0C
#712270000000
1!
1*
b11 6
19
1>
1C
b11 G
#712280000000
0!
0*
09
0>
0C
#712290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#712300000000
0!
0*
09
0>
0C
#712310000000
1!
1*
b101 6
19
1>
1C
b101 G
#712320000000
0!
0*
09
0>
0C
#712330000000
1!
1*
b110 6
19
1>
1C
b110 G
#712340000000
0!
0*
09
0>
0C
#712350000000
1!
1*
b111 6
19
1>
1C
b111 G
#712360000000
0!
0*
09
0>
0C
#712370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#712380000000
0!
0*
09
0>
0C
#712390000000
1!
1*
b1 6
19
1>
1C
b1 G
#712400000000
0!
0*
09
0>
0C
#712410000000
1!
1*
b10 6
19
1>
1C
b10 G
#712420000000
0!
0*
09
0>
0C
#712430000000
1!
1*
b11 6
19
1>
1C
b11 G
#712440000000
0!
0*
09
0>
0C
#712450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#712460000000
0!
0*
09
0>
0C
#712470000000
1!
1*
b101 6
19
1>
1C
b101 G
#712480000000
0!
0*
09
0>
0C
#712490000000
1!
1*
b110 6
19
1>
1C
b110 G
#712500000000
0!
0*
09
0>
0C
#712510000000
1!
1*
b111 6
19
1>
1C
b111 G
#712520000000
0!
0*
09
0>
0C
#712530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#712540000000
0!
0*
09
0>
0C
#712550000000
1!
1*
b1 6
19
1>
1C
b1 G
#712560000000
0!
0*
09
0>
0C
#712570000000
1!
1*
b10 6
19
1>
1C
b10 G
#712580000000
0!
0*
09
0>
0C
#712590000000
1!
1*
b11 6
19
1>
1C
b11 G
#712600000000
0!
0*
09
0>
0C
#712610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#712620000000
0!
0*
09
0>
0C
#712630000000
1!
1*
b101 6
19
1>
1C
b101 G
#712640000000
0!
0*
09
0>
0C
#712650000000
1!
1*
b110 6
19
1>
1C
b110 G
#712660000000
0!
0*
09
0>
0C
#712670000000
1!
1*
b111 6
19
1>
1C
b111 G
#712680000000
0!
1"
0*
1+
09
1:
0>
0C
#712690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#712700000000
0!
0*
09
0>
0C
#712710000000
1!
1*
b1 6
19
1>
1C
b1 G
#712720000000
0!
0*
09
0>
0C
#712730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#712740000000
0!
0*
09
0>
0C
#712750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#712760000000
0!
0*
09
0>
0C
#712770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#712780000000
0!
0*
09
0>
0C
#712790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#712800000000
0!
0#
0*
0,
09
0>
0?
0C
#712810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#712820000000
0!
0*
09
0>
0C
#712830000000
1!
1*
19
1>
1C
#712840000000
0!
0*
09
0>
0C
#712850000000
1!
1*
19
1>
1C
#712860000000
0!
0*
09
0>
0C
#712870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#712880000000
0!
0*
09
0>
0C
#712890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#712900000000
0!
0*
09
0>
0C
#712910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#712920000000
0!
0*
09
0>
0C
#712930000000
1!
1*
b10 6
19
1>
1C
b10 G
#712940000000
0!
0*
09
0>
0C
#712950000000
1!
1*
b11 6
19
1>
1C
b11 G
#712960000000
0!
0*
09
0>
0C
#712970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#712980000000
0!
0*
09
0>
0C
#712990000000
1!
1*
b101 6
19
1>
1C
b101 G
#713000000000
0!
0*
09
0>
0C
#713010000000
1!
1*
b110 6
19
1>
1C
b110 G
#713020000000
0!
0*
09
0>
0C
#713030000000
1!
1*
b111 6
19
1>
1C
b111 G
#713040000000
0!
0*
09
0>
0C
#713050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#713060000000
0!
0*
09
0>
0C
#713070000000
1!
1*
b1 6
19
1>
1C
b1 G
#713080000000
0!
0*
09
0>
0C
#713090000000
1!
1*
b10 6
19
1>
1C
b10 G
#713100000000
0!
0*
09
0>
0C
#713110000000
1!
1*
b11 6
19
1>
1C
b11 G
#713120000000
0!
0*
09
0>
0C
#713130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#713140000000
0!
0*
09
0>
0C
#713150000000
1!
1*
b101 6
19
1>
1C
b101 G
#713160000000
0!
0*
09
0>
0C
#713170000000
1!
1*
b110 6
19
1>
1C
b110 G
#713180000000
0!
0*
09
0>
0C
#713190000000
1!
1*
b111 6
19
1>
1C
b111 G
#713200000000
0!
0*
09
0>
0C
#713210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#713220000000
0!
0*
09
0>
0C
#713230000000
1!
1*
b1 6
19
1>
1C
b1 G
#713240000000
0!
0*
09
0>
0C
#713250000000
1!
1*
b10 6
19
1>
1C
b10 G
#713260000000
0!
0*
09
0>
0C
#713270000000
1!
1*
b11 6
19
1>
1C
b11 G
#713280000000
0!
0*
09
0>
0C
#713290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#713300000000
0!
0*
09
0>
0C
#713310000000
1!
1*
b101 6
19
1>
1C
b101 G
#713320000000
0!
0*
09
0>
0C
#713330000000
1!
1*
b110 6
19
1>
1C
b110 G
#713340000000
0!
0*
09
0>
0C
#713350000000
1!
1*
b111 6
19
1>
1C
b111 G
#713360000000
0!
1"
0*
1+
09
1:
0>
0C
#713370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#713380000000
0!
0*
09
0>
0C
#713390000000
1!
1*
b1 6
19
1>
1C
b1 G
#713400000000
0!
0*
09
0>
0C
#713410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#713420000000
0!
0*
09
0>
0C
#713430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#713440000000
0!
0*
09
0>
0C
#713450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#713460000000
0!
0*
09
0>
0C
#713470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#713480000000
0!
0#
0*
0,
09
0>
0?
0C
#713490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#713500000000
0!
0*
09
0>
0C
#713510000000
1!
1*
19
1>
1C
#713520000000
0!
0*
09
0>
0C
#713530000000
1!
1*
19
1>
1C
#713540000000
0!
0*
09
0>
0C
#713550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#713560000000
0!
0*
09
0>
0C
#713570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#713580000000
0!
0*
09
0>
0C
#713590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#713600000000
0!
0*
09
0>
0C
#713610000000
1!
1*
b10 6
19
1>
1C
b10 G
#713620000000
0!
0*
09
0>
0C
#713630000000
1!
1*
b11 6
19
1>
1C
b11 G
#713640000000
0!
0*
09
0>
0C
#713650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#713660000000
0!
0*
09
0>
0C
#713670000000
1!
1*
b101 6
19
1>
1C
b101 G
#713680000000
0!
0*
09
0>
0C
#713690000000
1!
1*
b110 6
19
1>
1C
b110 G
#713700000000
0!
0*
09
0>
0C
#713710000000
1!
1*
b111 6
19
1>
1C
b111 G
#713720000000
0!
0*
09
0>
0C
#713730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#713740000000
0!
0*
09
0>
0C
#713750000000
1!
1*
b1 6
19
1>
1C
b1 G
#713760000000
0!
0*
09
0>
0C
#713770000000
1!
1*
b10 6
19
1>
1C
b10 G
#713780000000
0!
0*
09
0>
0C
#713790000000
1!
1*
b11 6
19
1>
1C
b11 G
#713800000000
0!
0*
09
0>
0C
#713810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#713820000000
0!
0*
09
0>
0C
#713830000000
1!
1*
b101 6
19
1>
1C
b101 G
#713840000000
0!
0*
09
0>
0C
#713850000000
1!
1*
b110 6
19
1>
1C
b110 G
#713860000000
0!
0*
09
0>
0C
#713870000000
1!
1*
b111 6
19
1>
1C
b111 G
#713880000000
0!
0*
09
0>
0C
#713890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#713900000000
0!
0*
09
0>
0C
#713910000000
1!
1*
b1 6
19
1>
1C
b1 G
#713920000000
0!
0*
09
0>
0C
#713930000000
1!
1*
b10 6
19
1>
1C
b10 G
#713940000000
0!
0*
09
0>
0C
#713950000000
1!
1*
b11 6
19
1>
1C
b11 G
#713960000000
0!
0*
09
0>
0C
#713970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#713980000000
0!
0*
09
0>
0C
#713990000000
1!
1*
b101 6
19
1>
1C
b101 G
#714000000000
0!
0*
09
0>
0C
#714010000000
1!
1*
b110 6
19
1>
1C
b110 G
#714020000000
0!
0*
09
0>
0C
#714030000000
1!
1*
b111 6
19
1>
1C
b111 G
#714040000000
0!
1"
0*
1+
09
1:
0>
0C
#714050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#714060000000
0!
0*
09
0>
0C
#714070000000
1!
1*
b1 6
19
1>
1C
b1 G
#714080000000
0!
0*
09
0>
0C
#714090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#714100000000
0!
0*
09
0>
0C
#714110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#714120000000
0!
0*
09
0>
0C
#714130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#714140000000
0!
0*
09
0>
0C
#714150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#714160000000
0!
0#
0*
0,
09
0>
0?
0C
#714170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#714180000000
0!
0*
09
0>
0C
#714190000000
1!
1*
19
1>
1C
#714200000000
0!
0*
09
0>
0C
#714210000000
1!
1*
19
1>
1C
#714220000000
0!
0*
09
0>
0C
#714230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#714240000000
0!
0*
09
0>
0C
#714250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#714260000000
0!
0*
09
0>
0C
#714270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#714280000000
0!
0*
09
0>
0C
#714290000000
1!
1*
b10 6
19
1>
1C
b10 G
#714300000000
0!
0*
09
0>
0C
#714310000000
1!
1*
b11 6
19
1>
1C
b11 G
#714320000000
0!
0*
09
0>
0C
#714330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#714340000000
0!
0*
09
0>
0C
#714350000000
1!
1*
b101 6
19
1>
1C
b101 G
#714360000000
0!
0*
09
0>
0C
#714370000000
1!
1*
b110 6
19
1>
1C
b110 G
#714380000000
0!
0*
09
0>
0C
#714390000000
1!
1*
b111 6
19
1>
1C
b111 G
#714400000000
0!
0*
09
0>
0C
#714410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#714420000000
0!
0*
09
0>
0C
#714430000000
1!
1*
b1 6
19
1>
1C
b1 G
#714440000000
0!
0*
09
0>
0C
#714450000000
1!
1*
b10 6
19
1>
1C
b10 G
#714460000000
0!
0*
09
0>
0C
#714470000000
1!
1*
b11 6
19
1>
1C
b11 G
#714480000000
0!
0*
09
0>
0C
#714490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#714500000000
0!
0*
09
0>
0C
#714510000000
1!
1*
b101 6
19
1>
1C
b101 G
#714520000000
0!
0*
09
0>
0C
#714530000000
1!
1*
b110 6
19
1>
1C
b110 G
#714540000000
0!
0*
09
0>
0C
#714550000000
1!
1*
b111 6
19
1>
1C
b111 G
#714560000000
0!
0*
09
0>
0C
#714570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#714580000000
0!
0*
09
0>
0C
#714590000000
1!
1*
b1 6
19
1>
1C
b1 G
#714600000000
0!
0*
09
0>
0C
#714610000000
1!
1*
b10 6
19
1>
1C
b10 G
#714620000000
0!
0*
09
0>
0C
#714630000000
1!
1*
b11 6
19
1>
1C
b11 G
#714640000000
0!
0*
09
0>
0C
#714650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#714660000000
0!
0*
09
0>
0C
#714670000000
1!
1*
b101 6
19
1>
1C
b101 G
#714680000000
0!
0*
09
0>
0C
#714690000000
1!
1*
b110 6
19
1>
1C
b110 G
#714700000000
0!
0*
09
0>
0C
#714710000000
1!
1*
b111 6
19
1>
1C
b111 G
#714720000000
0!
1"
0*
1+
09
1:
0>
0C
#714730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#714740000000
0!
0*
09
0>
0C
#714750000000
1!
1*
b1 6
19
1>
1C
b1 G
#714760000000
0!
0*
09
0>
0C
#714770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#714780000000
0!
0*
09
0>
0C
#714790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#714800000000
0!
0*
09
0>
0C
#714810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#714820000000
0!
0*
09
0>
0C
#714830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#714840000000
0!
0#
0*
0,
09
0>
0?
0C
#714850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#714860000000
0!
0*
09
0>
0C
#714870000000
1!
1*
19
1>
1C
#714880000000
0!
0*
09
0>
0C
#714890000000
1!
1*
19
1>
1C
#714900000000
0!
0*
09
0>
0C
#714910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#714920000000
0!
0*
09
0>
0C
#714930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#714940000000
0!
0*
09
0>
0C
#714950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#714960000000
0!
0*
09
0>
0C
#714970000000
1!
1*
b10 6
19
1>
1C
b10 G
#714980000000
0!
0*
09
0>
0C
#714990000000
1!
1*
b11 6
19
1>
1C
b11 G
#715000000000
0!
0*
09
0>
0C
#715010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#715020000000
0!
0*
09
0>
0C
#715030000000
1!
1*
b101 6
19
1>
1C
b101 G
#715040000000
0!
0*
09
0>
0C
#715050000000
1!
1*
b110 6
19
1>
1C
b110 G
#715060000000
0!
0*
09
0>
0C
#715070000000
1!
1*
b111 6
19
1>
1C
b111 G
#715080000000
0!
0*
09
0>
0C
#715090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#715100000000
0!
0*
09
0>
0C
#715110000000
1!
1*
b1 6
19
1>
1C
b1 G
#715120000000
0!
0*
09
0>
0C
#715130000000
1!
1*
b10 6
19
1>
1C
b10 G
#715140000000
0!
0*
09
0>
0C
#715150000000
1!
1*
b11 6
19
1>
1C
b11 G
#715160000000
0!
0*
09
0>
0C
#715170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#715180000000
0!
0*
09
0>
0C
#715190000000
1!
1*
b101 6
19
1>
1C
b101 G
#715200000000
0!
0*
09
0>
0C
#715210000000
1!
1*
b110 6
19
1>
1C
b110 G
#715220000000
0!
0*
09
0>
0C
#715230000000
1!
1*
b111 6
19
1>
1C
b111 G
#715240000000
0!
0*
09
0>
0C
#715250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#715260000000
0!
0*
09
0>
0C
#715270000000
1!
1*
b1 6
19
1>
1C
b1 G
#715280000000
0!
0*
09
0>
0C
#715290000000
1!
1*
b10 6
19
1>
1C
b10 G
#715300000000
0!
0*
09
0>
0C
#715310000000
1!
1*
b11 6
19
1>
1C
b11 G
#715320000000
0!
0*
09
0>
0C
#715330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#715340000000
0!
0*
09
0>
0C
#715350000000
1!
1*
b101 6
19
1>
1C
b101 G
#715360000000
0!
0*
09
0>
0C
#715370000000
1!
1*
b110 6
19
1>
1C
b110 G
#715380000000
0!
0*
09
0>
0C
#715390000000
1!
1*
b111 6
19
1>
1C
b111 G
#715400000000
0!
1"
0*
1+
09
1:
0>
0C
#715410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#715420000000
0!
0*
09
0>
0C
#715430000000
1!
1*
b1 6
19
1>
1C
b1 G
#715440000000
0!
0*
09
0>
0C
#715450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#715460000000
0!
0*
09
0>
0C
#715470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#715480000000
0!
0*
09
0>
0C
#715490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#715500000000
0!
0*
09
0>
0C
#715510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#715520000000
0!
0#
0*
0,
09
0>
0?
0C
#715530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#715540000000
0!
0*
09
0>
0C
#715550000000
1!
1*
19
1>
1C
#715560000000
0!
0*
09
0>
0C
#715570000000
1!
1*
19
1>
1C
#715580000000
0!
0*
09
0>
0C
#715590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#715600000000
0!
0*
09
0>
0C
#715610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#715620000000
0!
0*
09
0>
0C
#715630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#715640000000
0!
0*
09
0>
0C
#715650000000
1!
1*
b10 6
19
1>
1C
b10 G
#715660000000
0!
0*
09
0>
0C
#715670000000
1!
1*
b11 6
19
1>
1C
b11 G
#715680000000
0!
0*
09
0>
0C
#715690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#715700000000
0!
0*
09
0>
0C
#715710000000
1!
1*
b101 6
19
1>
1C
b101 G
#715720000000
0!
0*
09
0>
0C
#715730000000
1!
1*
b110 6
19
1>
1C
b110 G
#715740000000
0!
0*
09
0>
0C
#715750000000
1!
1*
b111 6
19
1>
1C
b111 G
#715760000000
0!
0*
09
0>
0C
#715770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#715780000000
0!
0*
09
0>
0C
#715790000000
1!
1*
b1 6
19
1>
1C
b1 G
#715800000000
0!
0*
09
0>
0C
#715810000000
1!
1*
b10 6
19
1>
1C
b10 G
#715820000000
0!
0*
09
0>
0C
#715830000000
1!
1*
b11 6
19
1>
1C
b11 G
#715840000000
0!
0*
09
0>
0C
#715850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#715860000000
0!
0*
09
0>
0C
#715870000000
1!
1*
b101 6
19
1>
1C
b101 G
#715880000000
0!
0*
09
0>
0C
#715890000000
1!
1*
b110 6
19
1>
1C
b110 G
#715900000000
0!
0*
09
0>
0C
#715910000000
1!
1*
b111 6
19
1>
1C
b111 G
#715920000000
0!
0*
09
0>
0C
#715930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#715940000000
0!
0*
09
0>
0C
#715950000000
1!
1*
b1 6
19
1>
1C
b1 G
#715960000000
0!
0*
09
0>
0C
#715970000000
1!
1*
b10 6
19
1>
1C
b10 G
#715980000000
0!
0*
09
0>
0C
#715990000000
1!
1*
b11 6
19
1>
1C
b11 G
#716000000000
0!
0*
09
0>
0C
#716010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#716020000000
0!
0*
09
0>
0C
#716030000000
1!
1*
b101 6
19
1>
1C
b101 G
#716040000000
0!
0*
09
0>
0C
#716050000000
1!
1*
b110 6
19
1>
1C
b110 G
#716060000000
0!
0*
09
0>
0C
#716070000000
1!
1*
b111 6
19
1>
1C
b111 G
#716080000000
0!
1"
0*
1+
09
1:
0>
0C
#716090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#716100000000
0!
0*
09
0>
0C
#716110000000
1!
1*
b1 6
19
1>
1C
b1 G
#716120000000
0!
0*
09
0>
0C
#716130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#716140000000
0!
0*
09
0>
0C
#716150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#716160000000
0!
0*
09
0>
0C
#716170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#716180000000
0!
0*
09
0>
0C
#716190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#716200000000
0!
0#
0*
0,
09
0>
0?
0C
#716210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#716220000000
0!
0*
09
0>
0C
#716230000000
1!
1*
19
1>
1C
#716240000000
0!
0*
09
0>
0C
#716250000000
1!
1*
19
1>
1C
#716260000000
0!
0*
09
0>
0C
#716270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#716280000000
0!
0*
09
0>
0C
#716290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#716300000000
0!
0*
09
0>
0C
#716310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#716320000000
0!
0*
09
0>
0C
#716330000000
1!
1*
b10 6
19
1>
1C
b10 G
#716340000000
0!
0*
09
0>
0C
#716350000000
1!
1*
b11 6
19
1>
1C
b11 G
#716360000000
0!
0*
09
0>
0C
#716370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#716380000000
0!
0*
09
0>
0C
#716390000000
1!
1*
b101 6
19
1>
1C
b101 G
#716400000000
0!
0*
09
0>
0C
#716410000000
1!
1*
b110 6
19
1>
1C
b110 G
#716420000000
0!
0*
09
0>
0C
#716430000000
1!
1*
b111 6
19
1>
1C
b111 G
#716440000000
0!
0*
09
0>
0C
#716450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#716460000000
0!
0*
09
0>
0C
#716470000000
1!
1*
b1 6
19
1>
1C
b1 G
#716480000000
0!
0*
09
0>
0C
#716490000000
1!
1*
b10 6
19
1>
1C
b10 G
#716500000000
0!
0*
09
0>
0C
#716510000000
1!
1*
b11 6
19
1>
1C
b11 G
#716520000000
0!
0*
09
0>
0C
#716530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#716540000000
0!
0*
09
0>
0C
#716550000000
1!
1*
b101 6
19
1>
1C
b101 G
#716560000000
0!
0*
09
0>
0C
#716570000000
1!
1*
b110 6
19
1>
1C
b110 G
#716580000000
0!
0*
09
0>
0C
#716590000000
1!
1*
b111 6
19
1>
1C
b111 G
#716600000000
0!
0*
09
0>
0C
#716610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#716620000000
0!
0*
09
0>
0C
#716630000000
1!
1*
b1 6
19
1>
1C
b1 G
#716640000000
0!
0*
09
0>
0C
#716650000000
1!
1*
b10 6
19
1>
1C
b10 G
#716660000000
0!
0*
09
0>
0C
#716670000000
1!
1*
b11 6
19
1>
1C
b11 G
#716680000000
0!
0*
09
0>
0C
#716690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#716700000000
0!
0*
09
0>
0C
#716710000000
1!
1*
b101 6
19
1>
1C
b101 G
#716720000000
0!
0*
09
0>
0C
#716730000000
1!
1*
b110 6
19
1>
1C
b110 G
#716740000000
0!
0*
09
0>
0C
#716750000000
1!
1*
b111 6
19
1>
1C
b111 G
#716760000000
0!
1"
0*
1+
09
1:
0>
0C
#716770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#716780000000
0!
0*
09
0>
0C
#716790000000
1!
1*
b1 6
19
1>
1C
b1 G
#716800000000
0!
0*
09
0>
0C
#716810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#716820000000
0!
0*
09
0>
0C
#716830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#716840000000
0!
0*
09
0>
0C
#716850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#716860000000
0!
0*
09
0>
0C
#716870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#716880000000
0!
0#
0*
0,
09
0>
0?
0C
#716890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#716900000000
0!
0*
09
0>
0C
#716910000000
1!
1*
19
1>
1C
#716920000000
0!
0*
09
0>
0C
#716930000000
1!
1*
19
1>
1C
#716940000000
0!
0*
09
0>
0C
#716950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#716960000000
0!
0*
09
0>
0C
#716970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#716980000000
0!
0*
09
0>
0C
#716990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#717000000000
0!
0*
09
0>
0C
#717010000000
1!
1*
b10 6
19
1>
1C
b10 G
#717020000000
0!
0*
09
0>
0C
#717030000000
1!
1*
b11 6
19
1>
1C
b11 G
#717040000000
0!
0*
09
0>
0C
#717050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#717060000000
0!
0*
09
0>
0C
#717070000000
1!
1*
b101 6
19
1>
1C
b101 G
#717080000000
0!
0*
09
0>
0C
#717090000000
1!
1*
b110 6
19
1>
1C
b110 G
#717100000000
0!
0*
09
0>
0C
#717110000000
1!
1*
b111 6
19
1>
1C
b111 G
#717120000000
0!
0*
09
0>
0C
#717130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#717140000000
0!
0*
09
0>
0C
#717150000000
1!
1*
b1 6
19
1>
1C
b1 G
#717160000000
0!
0*
09
0>
0C
#717170000000
1!
1*
b10 6
19
1>
1C
b10 G
#717180000000
0!
0*
09
0>
0C
#717190000000
1!
1*
b11 6
19
1>
1C
b11 G
#717200000000
0!
0*
09
0>
0C
#717210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#717220000000
0!
0*
09
0>
0C
#717230000000
1!
1*
b101 6
19
1>
1C
b101 G
#717240000000
0!
0*
09
0>
0C
#717250000000
1!
1*
b110 6
19
1>
1C
b110 G
#717260000000
0!
0*
09
0>
0C
#717270000000
1!
1*
b111 6
19
1>
1C
b111 G
#717280000000
0!
0*
09
0>
0C
#717290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#717300000000
0!
0*
09
0>
0C
#717310000000
1!
1*
b1 6
19
1>
1C
b1 G
#717320000000
0!
0*
09
0>
0C
#717330000000
1!
1*
b10 6
19
1>
1C
b10 G
#717340000000
0!
0*
09
0>
0C
#717350000000
1!
1*
b11 6
19
1>
1C
b11 G
#717360000000
0!
0*
09
0>
0C
#717370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#717380000000
0!
0*
09
0>
0C
#717390000000
1!
1*
b101 6
19
1>
1C
b101 G
#717400000000
0!
0*
09
0>
0C
#717410000000
1!
1*
b110 6
19
1>
1C
b110 G
#717420000000
0!
0*
09
0>
0C
#717430000000
1!
1*
b111 6
19
1>
1C
b111 G
#717440000000
0!
1"
0*
1+
09
1:
0>
0C
#717450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#717460000000
0!
0*
09
0>
0C
#717470000000
1!
1*
b1 6
19
1>
1C
b1 G
#717480000000
0!
0*
09
0>
0C
#717490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#717500000000
0!
0*
09
0>
0C
#717510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#717520000000
0!
0*
09
0>
0C
#717530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#717540000000
0!
0*
09
0>
0C
#717550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#717560000000
0!
0#
0*
0,
09
0>
0?
0C
#717570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#717580000000
0!
0*
09
0>
0C
#717590000000
1!
1*
19
1>
1C
#717600000000
0!
0*
09
0>
0C
#717610000000
1!
1*
19
1>
1C
#717620000000
0!
0*
09
0>
0C
#717630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#717640000000
0!
0*
09
0>
0C
#717650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#717660000000
0!
0*
09
0>
0C
#717670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#717680000000
0!
0*
09
0>
0C
#717690000000
1!
1*
b10 6
19
1>
1C
b10 G
#717700000000
0!
0*
09
0>
0C
#717710000000
1!
1*
b11 6
19
1>
1C
b11 G
#717720000000
0!
0*
09
0>
0C
#717730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#717740000000
0!
0*
09
0>
0C
#717750000000
1!
1*
b101 6
19
1>
1C
b101 G
#717760000000
0!
0*
09
0>
0C
#717770000000
1!
1*
b110 6
19
1>
1C
b110 G
#717780000000
0!
0*
09
0>
0C
#717790000000
1!
1*
b111 6
19
1>
1C
b111 G
#717800000000
0!
0*
09
0>
0C
#717810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#717820000000
0!
0*
09
0>
0C
#717830000000
1!
1*
b1 6
19
1>
1C
b1 G
#717840000000
0!
0*
09
0>
0C
#717850000000
1!
1*
b10 6
19
1>
1C
b10 G
#717860000000
0!
0*
09
0>
0C
#717870000000
1!
1*
b11 6
19
1>
1C
b11 G
#717880000000
0!
0*
09
0>
0C
#717890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#717900000000
0!
0*
09
0>
0C
#717910000000
1!
1*
b101 6
19
1>
1C
b101 G
#717920000000
0!
0*
09
0>
0C
#717930000000
1!
1*
b110 6
19
1>
1C
b110 G
#717940000000
0!
0*
09
0>
0C
#717950000000
1!
1*
b111 6
19
1>
1C
b111 G
#717960000000
0!
0*
09
0>
0C
#717970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#717980000000
0!
0*
09
0>
0C
#717990000000
1!
1*
b1 6
19
1>
1C
b1 G
#718000000000
0!
0*
09
0>
0C
#718010000000
1!
1*
b10 6
19
1>
1C
b10 G
#718020000000
0!
0*
09
0>
0C
#718030000000
1!
1*
b11 6
19
1>
1C
b11 G
#718040000000
0!
0*
09
0>
0C
#718050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#718060000000
0!
0*
09
0>
0C
#718070000000
1!
1*
b101 6
19
1>
1C
b101 G
#718080000000
0!
0*
09
0>
0C
#718090000000
1!
1*
b110 6
19
1>
1C
b110 G
#718100000000
0!
0*
09
0>
0C
#718110000000
1!
1*
b111 6
19
1>
1C
b111 G
#718120000000
0!
1"
0*
1+
09
1:
0>
0C
#718130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#718140000000
0!
0*
09
0>
0C
#718150000000
1!
1*
b1 6
19
1>
1C
b1 G
#718160000000
0!
0*
09
0>
0C
#718170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#718180000000
0!
0*
09
0>
0C
#718190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#718200000000
0!
0*
09
0>
0C
#718210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#718220000000
0!
0*
09
0>
0C
#718230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#718240000000
0!
0#
0*
0,
09
0>
0?
0C
#718250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#718260000000
0!
0*
09
0>
0C
#718270000000
1!
1*
19
1>
1C
#718280000000
0!
0*
09
0>
0C
#718290000000
1!
1*
19
1>
1C
#718300000000
0!
0*
09
0>
0C
#718310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#718320000000
0!
0*
09
0>
0C
#718330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#718340000000
0!
0*
09
0>
0C
#718350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#718360000000
0!
0*
09
0>
0C
#718370000000
1!
1*
b10 6
19
1>
1C
b10 G
#718380000000
0!
0*
09
0>
0C
#718390000000
1!
1*
b11 6
19
1>
1C
b11 G
#718400000000
0!
0*
09
0>
0C
#718410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#718420000000
0!
0*
09
0>
0C
#718430000000
1!
1*
b101 6
19
1>
1C
b101 G
#718440000000
0!
0*
09
0>
0C
#718450000000
1!
1*
b110 6
19
1>
1C
b110 G
#718460000000
0!
0*
09
0>
0C
#718470000000
1!
1*
b111 6
19
1>
1C
b111 G
#718480000000
0!
0*
09
0>
0C
#718490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#718500000000
0!
0*
09
0>
0C
#718510000000
1!
1*
b1 6
19
1>
1C
b1 G
#718520000000
0!
0*
09
0>
0C
#718530000000
1!
1*
b10 6
19
1>
1C
b10 G
#718540000000
0!
0*
09
0>
0C
#718550000000
1!
1*
b11 6
19
1>
1C
b11 G
#718560000000
0!
0*
09
0>
0C
#718570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#718580000000
0!
0*
09
0>
0C
#718590000000
1!
1*
b101 6
19
1>
1C
b101 G
#718600000000
0!
0*
09
0>
0C
#718610000000
1!
1*
b110 6
19
1>
1C
b110 G
#718620000000
0!
0*
09
0>
0C
#718630000000
1!
1*
b111 6
19
1>
1C
b111 G
#718640000000
0!
0*
09
0>
0C
#718650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#718660000000
0!
0*
09
0>
0C
#718670000000
1!
1*
b1 6
19
1>
1C
b1 G
#718680000000
0!
0*
09
0>
0C
#718690000000
1!
1*
b10 6
19
1>
1C
b10 G
#718700000000
0!
0*
09
0>
0C
#718710000000
1!
1*
b11 6
19
1>
1C
b11 G
#718720000000
0!
0*
09
0>
0C
#718730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#718740000000
0!
0*
09
0>
0C
#718750000000
1!
1*
b101 6
19
1>
1C
b101 G
#718760000000
0!
0*
09
0>
0C
#718770000000
1!
1*
b110 6
19
1>
1C
b110 G
#718780000000
0!
0*
09
0>
0C
#718790000000
1!
1*
b111 6
19
1>
1C
b111 G
#718800000000
0!
1"
0*
1+
09
1:
0>
0C
#718810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#718820000000
0!
0*
09
0>
0C
#718830000000
1!
1*
b1 6
19
1>
1C
b1 G
#718840000000
0!
0*
09
0>
0C
#718850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#718860000000
0!
0*
09
0>
0C
#718870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#718880000000
0!
0*
09
0>
0C
#718890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#718900000000
0!
0*
09
0>
0C
#718910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#718920000000
0!
0#
0*
0,
09
0>
0?
0C
#718930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#718940000000
0!
0*
09
0>
0C
#718950000000
1!
1*
19
1>
1C
#718960000000
0!
0*
09
0>
0C
#718970000000
1!
1*
19
1>
1C
#718980000000
0!
0*
09
0>
0C
#718990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#719000000000
0!
0*
09
0>
0C
#719010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#719020000000
0!
0*
09
0>
0C
#719030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#719040000000
0!
0*
09
0>
0C
#719050000000
1!
1*
b10 6
19
1>
1C
b10 G
#719060000000
0!
0*
09
0>
0C
#719070000000
1!
1*
b11 6
19
1>
1C
b11 G
#719080000000
0!
0*
09
0>
0C
#719090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#719100000000
0!
0*
09
0>
0C
#719110000000
1!
1*
b101 6
19
1>
1C
b101 G
#719120000000
0!
0*
09
0>
0C
#719130000000
1!
1*
b110 6
19
1>
1C
b110 G
#719140000000
0!
0*
09
0>
0C
#719150000000
1!
1*
b111 6
19
1>
1C
b111 G
#719160000000
0!
0*
09
0>
0C
#719170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#719180000000
0!
0*
09
0>
0C
#719190000000
1!
1*
b1 6
19
1>
1C
b1 G
#719200000000
0!
0*
09
0>
0C
#719210000000
1!
1*
b10 6
19
1>
1C
b10 G
#719220000000
0!
0*
09
0>
0C
#719230000000
1!
1*
b11 6
19
1>
1C
b11 G
#719240000000
0!
0*
09
0>
0C
#719250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#719260000000
0!
0*
09
0>
0C
#719270000000
1!
1*
b101 6
19
1>
1C
b101 G
#719280000000
0!
0*
09
0>
0C
#719290000000
1!
1*
b110 6
19
1>
1C
b110 G
#719300000000
0!
0*
09
0>
0C
#719310000000
1!
1*
b111 6
19
1>
1C
b111 G
#719320000000
0!
0*
09
0>
0C
#719330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#719340000000
0!
0*
09
0>
0C
#719350000000
1!
1*
b1 6
19
1>
1C
b1 G
#719360000000
0!
0*
09
0>
0C
#719370000000
1!
1*
b10 6
19
1>
1C
b10 G
#719380000000
0!
0*
09
0>
0C
#719390000000
1!
1*
b11 6
19
1>
1C
b11 G
#719400000000
0!
0*
09
0>
0C
#719410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#719420000000
0!
0*
09
0>
0C
#719430000000
1!
1*
b101 6
19
1>
1C
b101 G
#719440000000
0!
0*
09
0>
0C
#719450000000
1!
1*
b110 6
19
1>
1C
b110 G
#719460000000
0!
0*
09
0>
0C
#719470000000
1!
1*
b111 6
19
1>
1C
b111 G
#719480000000
0!
1"
0*
1+
09
1:
0>
0C
#719490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#719500000000
0!
0*
09
0>
0C
#719510000000
1!
1*
b1 6
19
1>
1C
b1 G
#719520000000
0!
0*
09
0>
0C
#719530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#719540000000
0!
0*
09
0>
0C
#719550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#719560000000
0!
0*
09
0>
0C
#719570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#719580000000
0!
0*
09
0>
0C
#719590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#719600000000
0!
0#
0*
0,
09
0>
0?
0C
#719610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#719620000000
0!
0*
09
0>
0C
#719630000000
1!
1*
19
1>
1C
#719640000000
0!
0*
09
0>
0C
#719650000000
1!
1*
19
1>
1C
#719660000000
0!
0*
09
0>
0C
#719670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#719680000000
0!
0*
09
0>
0C
#719690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#719700000000
0!
0*
09
0>
0C
#719710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#719720000000
0!
0*
09
0>
0C
#719730000000
1!
1*
b10 6
19
1>
1C
b10 G
#719740000000
0!
0*
09
0>
0C
#719750000000
1!
1*
b11 6
19
1>
1C
b11 G
#719760000000
0!
0*
09
0>
0C
#719770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#719780000000
0!
0*
09
0>
0C
#719790000000
1!
1*
b101 6
19
1>
1C
b101 G
#719800000000
0!
0*
09
0>
0C
#719810000000
1!
1*
b110 6
19
1>
1C
b110 G
#719820000000
0!
0*
09
0>
0C
#719830000000
1!
1*
b111 6
19
1>
1C
b111 G
#719840000000
0!
0*
09
0>
0C
#719850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#719860000000
0!
0*
09
0>
0C
#719870000000
1!
1*
b1 6
19
1>
1C
b1 G
#719880000000
0!
0*
09
0>
0C
#719890000000
1!
1*
b10 6
19
1>
1C
b10 G
#719900000000
0!
0*
09
0>
0C
#719910000000
1!
1*
b11 6
19
1>
1C
b11 G
#719920000000
0!
0*
09
0>
0C
#719930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#719940000000
0!
0*
09
0>
0C
#719950000000
1!
1*
b101 6
19
1>
1C
b101 G
#719960000000
0!
0*
09
0>
0C
#719970000000
1!
1*
b110 6
19
1>
1C
b110 G
#719980000000
0!
0*
09
0>
0C
#719990000000
1!
1*
b111 6
19
1>
1C
b111 G
#720000000000
0!
0*
09
0>
0C
#720010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#720020000000
0!
0*
09
0>
0C
#720030000000
1!
1*
b1 6
19
1>
1C
b1 G
#720040000000
0!
0*
09
0>
0C
#720050000000
1!
1*
b10 6
19
1>
1C
b10 G
#720060000000
0!
0*
09
0>
0C
#720070000000
1!
1*
b11 6
19
1>
1C
b11 G
#720080000000
0!
0*
09
0>
0C
#720090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#720100000000
0!
0*
09
0>
0C
#720110000000
1!
1*
b101 6
19
1>
1C
b101 G
#720120000000
0!
0*
09
0>
0C
#720130000000
1!
1*
b110 6
19
1>
1C
b110 G
#720140000000
0!
0*
09
0>
0C
#720150000000
1!
1*
b111 6
19
1>
1C
b111 G
#720160000000
0!
1"
0*
1+
09
1:
0>
0C
#720170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#720180000000
0!
0*
09
0>
0C
#720190000000
1!
1*
b1 6
19
1>
1C
b1 G
#720200000000
0!
0*
09
0>
0C
#720210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#720220000000
0!
0*
09
0>
0C
#720230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#720240000000
0!
0*
09
0>
0C
#720250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#720260000000
0!
0*
09
0>
0C
#720270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#720280000000
0!
0#
0*
0,
09
0>
0?
0C
#720290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#720300000000
0!
0*
09
0>
0C
#720310000000
1!
1*
19
1>
1C
#720320000000
0!
0*
09
0>
0C
#720330000000
1!
1*
19
1>
1C
#720340000000
0!
0*
09
0>
0C
#720350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#720360000000
0!
0*
09
0>
0C
#720370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#720380000000
0!
0*
09
0>
0C
#720390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#720400000000
0!
0*
09
0>
0C
#720410000000
1!
1*
b10 6
19
1>
1C
b10 G
#720420000000
0!
0*
09
0>
0C
#720430000000
1!
1*
b11 6
19
1>
1C
b11 G
#720440000000
0!
0*
09
0>
0C
#720450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#720460000000
0!
0*
09
0>
0C
#720470000000
1!
1*
b101 6
19
1>
1C
b101 G
#720480000000
0!
0*
09
0>
0C
#720490000000
1!
1*
b110 6
19
1>
1C
b110 G
#720500000000
0!
0*
09
0>
0C
#720510000000
1!
1*
b111 6
19
1>
1C
b111 G
#720520000000
0!
0*
09
0>
0C
#720530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#720540000000
0!
0*
09
0>
0C
#720550000000
1!
1*
b1 6
19
1>
1C
b1 G
#720560000000
0!
0*
09
0>
0C
#720570000000
1!
1*
b10 6
19
1>
1C
b10 G
#720580000000
0!
0*
09
0>
0C
#720590000000
1!
1*
b11 6
19
1>
1C
b11 G
#720600000000
0!
0*
09
0>
0C
#720610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#720620000000
0!
0*
09
0>
0C
#720630000000
1!
1*
b101 6
19
1>
1C
b101 G
#720640000000
0!
0*
09
0>
0C
#720650000000
1!
1*
b110 6
19
1>
1C
b110 G
#720660000000
0!
0*
09
0>
0C
#720670000000
1!
1*
b111 6
19
1>
1C
b111 G
#720680000000
0!
0*
09
0>
0C
#720690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#720700000000
0!
0*
09
0>
0C
#720710000000
1!
1*
b1 6
19
1>
1C
b1 G
#720720000000
0!
0*
09
0>
0C
#720730000000
1!
1*
b10 6
19
1>
1C
b10 G
#720740000000
0!
0*
09
0>
0C
#720750000000
1!
1*
b11 6
19
1>
1C
b11 G
#720760000000
0!
0*
09
0>
0C
#720770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#720780000000
0!
0*
09
0>
0C
#720790000000
1!
1*
b101 6
19
1>
1C
b101 G
#720800000000
0!
0*
09
0>
0C
#720810000000
1!
1*
b110 6
19
1>
1C
b110 G
#720820000000
0!
0*
09
0>
0C
#720830000000
1!
1*
b111 6
19
1>
1C
b111 G
#720840000000
0!
1"
0*
1+
09
1:
0>
0C
#720850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#720860000000
0!
0*
09
0>
0C
#720870000000
1!
1*
b1 6
19
1>
1C
b1 G
#720880000000
0!
0*
09
0>
0C
#720890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#720900000000
0!
0*
09
0>
0C
#720910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#720920000000
0!
0*
09
0>
0C
#720930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#720940000000
0!
0*
09
0>
0C
#720950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#720960000000
0!
0#
0*
0,
09
0>
0?
0C
#720970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#720980000000
0!
0*
09
0>
0C
#720990000000
1!
1*
19
1>
1C
#721000000000
0!
0*
09
0>
0C
#721010000000
1!
1*
19
1>
1C
#721020000000
0!
0*
09
0>
0C
#721030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#721040000000
0!
0*
09
0>
0C
#721050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#721060000000
0!
0*
09
0>
0C
#721070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#721080000000
0!
0*
09
0>
0C
#721090000000
1!
1*
b10 6
19
1>
1C
b10 G
#721100000000
0!
0*
09
0>
0C
#721110000000
1!
1*
b11 6
19
1>
1C
b11 G
#721120000000
0!
0*
09
0>
0C
#721130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#721140000000
0!
0*
09
0>
0C
#721150000000
1!
1*
b101 6
19
1>
1C
b101 G
#721160000000
0!
0*
09
0>
0C
#721170000000
1!
1*
b110 6
19
1>
1C
b110 G
#721180000000
0!
0*
09
0>
0C
#721190000000
1!
1*
b111 6
19
1>
1C
b111 G
#721200000000
0!
0*
09
0>
0C
#721210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#721220000000
0!
0*
09
0>
0C
#721230000000
1!
1*
b1 6
19
1>
1C
b1 G
#721240000000
0!
0*
09
0>
0C
#721250000000
1!
1*
b10 6
19
1>
1C
b10 G
#721260000000
0!
0*
09
0>
0C
#721270000000
1!
1*
b11 6
19
1>
1C
b11 G
#721280000000
0!
0*
09
0>
0C
#721290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#721300000000
0!
0*
09
0>
0C
#721310000000
1!
1*
b101 6
19
1>
1C
b101 G
#721320000000
0!
0*
09
0>
0C
#721330000000
1!
1*
b110 6
19
1>
1C
b110 G
#721340000000
0!
0*
09
0>
0C
#721350000000
1!
1*
b111 6
19
1>
1C
b111 G
#721360000000
0!
0*
09
0>
0C
#721370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#721380000000
0!
0*
09
0>
0C
#721390000000
1!
1*
b1 6
19
1>
1C
b1 G
#721400000000
0!
0*
09
0>
0C
#721410000000
1!
1*
b10 6
19
1>
1C
b10 G
#721420000000
0!
0*
09
0>
0C
#721430000000
1!
1*
b11 6
19
1>
1C
b11 G
#721440000000
0!
0*
09
0>
0C
#721450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#721460000000
0!
0*
09
0>
0C
#721470000000
1!
1*
b101 6
19
1>
1C
b101 G
#721480000000
0!
0*
09
0>
0C
#721490000000
1!
1*
b110 6
19
1>
1C
b110 G
#721500000000
0!
0*
09
0>
0C
#721510000000
1!
1*
b111 6
19
1>
1C
b111 G
#721520000000
0!
1"
0*
1+
09
1:
0>
0C
#721530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#721540000000
0!
0*
09
0>
0C
#721550000000
1!
1*
b1 6
19
1>
1C
b1 G
#721560000000
0!
0*
09
0>
0C
#721570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#721580000000
0!
0*
09
0>
0C
#721590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#721600000000
0!
0*
09
0>
0C
#721610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#721620000000
0!
0*
09
0>
0C
#721630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#721640000000
0!
0#
0*
0,
09
0>
0?
0C
#721650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#721660000000
0!
0*
09
0>
0C
#721670000000
1!
1*
19
1>
1C
#721680000000
0!
0*
09
0>
0C
#721690000000
1!
1*
19
1>
1C
#721700000000
0!
0*
09
0>
0C
#721710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#721720000000
0!
0*
09
0>
0C
#721730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#721740000000
0!
0*
09
0>
0C
#721750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#721760000000
0!
0*
09
0>
0C
#721770000000
1!
1*
b10 6
19
1>
1C
b10 G
#721780000000
0!
0*
09
0>
0C
#721790000000
1!
1*
b11 6
19
1>
1C
b11 G
#721800000000
0!
0*
09
0>
0C
#721810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#721820000000
0!
0*
09
0>
0C
#721830000000
1!
1*
b101 6
19
1>
1C
b101 G
#721840000000
0!
0*
09
0>
0C
#721850000000
1!
1*
b110 6
19
1>
1C
b110 G
#721860000000
0!
0*
09
0>
0C
#721870000000
1!
1*
b111 6
19
1>
1C
b111 G
#721880000000
0!
0*
09
0>
0C
#721890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#721900000000
0!
0*
09
0>
0C
#721910000000
1!
1*
b1 6
19
1>
1C
b1 G
#721920000000
0!
0*
09
0>
0C
#721930000000
1!
1*
b10 6
19
1>
1C
b10 G
#721940000000
0!
0*
09
0>
0C
#721950000000
1!
1*
b11 6
19
1>
1C
b11 G
#721960000000
0!
0*
09
0>
0C
#721970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#721980000000
0!
0*
09
0>
0C
#721990000000
1!
1*
b101 6
19
1>
1C
b101 G
#722000000000
0!
0*
09
0>
0C
#722010000000
1!
1*
b110 6
19
1>
1C
b110 G
#722020000000
0!
0*
09
0>
0C
#722030000000
1!
1*
b111 6
19
1>
1C
b111 G
#722040000000
0!
0*
09
0>
0C
#722050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#722060000000
0!
0*
09
0>
0C
#722070000000
1!
1*
b1 6
19
1>
1C
b1 G
#722080000000
0!
0*
09
0>
0C
#722090000000
1!
1*
b10 6
19
1>
1C
b10 G
#722100000000
0!
0*
09
0>
0C
#722110000000
1!
1*
b11 6
19
1>
1C
b11 G
#722120000000
0!
0*
09
0>
0C
#722130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#722140000000
0!
0*
09
0>
0C
#722150000000
1!
1*
b101 6
19
1>
1C
b101 G
#722160000000
0!
0*
09
0>
0C
#722170000000
1!
1*
b110 6
19
1>
1C
b110 G
#722180000000
0!
0*
09
0>
0C
#722190000000
1!
1*
b111 6
19
1>
1C
b111 G
#722200000000
0!
1"
0*
1+
09
1:
0>
0C
#722210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#722220000000
0!
0*
09
0>
0C
#722230000000
1!
1*
b1 6
19
1>
1C
b1 G
#722240000000
0!
0*
09
0>
0C
#722250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#722260000000
0!
0*
09
0>
0C
#722270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#722280000000
0!
0*
09
0>
0C
#722290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#722300000000
0!
0*
09
0>
0C
#722310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#722320000000
0!
0#
0*
0,
09
0>
0?
0C
#722330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#722340000000
0!
0*
09
0>
0C
#722350000000
1!
1*
19
1>
1C
#722360000000
0!
0*
09
0>
0C
#722370000000
1!
1*
19
1>
1C
#722380000000
0!
0*
09
0>
0C
#722390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#722400000000
0!
0*
09
0>
0C
#722410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#722420000000
0!
0*
09
0>
0C
#722430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#722440000000
0!
0*
09
0>
0C
#722450000000
1!
1*
b10 6
19
1>
1C
b10 G
#722460000000
0!
0*
09
0>
0C
#722470000000
1!
1*
b11 6
19
1>
1C
b11 G
#722480000000
0!
0*
09
0>
0C
#722490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#722500000000
0!
0*
09
0>
0C
#722510000000
1!
1*
b101 6
19
1>
1C
b101 G
#722520000000
0!
0*
09
0>
0C
#722530000000
1!
1*
b110 6
19
1>
1C
b110 G
#722540000000
0!
0*
09
0>
0C
#722550000000
1!
1*
b111 6
19
1>
1C
b111 G
#722560000000
0!
0*
09
0>
0C
#722570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#722580000000
0!
0*
09
0>
0C
#722590000000
1!
1*
b1 6
19
1>
1C
b1 G
#722600000000
0!
0*
09
0>
0C
#722610000000
1!
1*
b10 6
19
1>
1C
b10 G
#722620000000
0!
0*
09
0>
0C
#722630000000
1!
1*
b11 6
19
1>
1C
b11 G
#722640000000
0!
0*
09
0>
0C
#722650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#722660000000
0!
0*
09
0>
0C
#722670000000
1!
1*
b101 6
19
1>
1C
b101 G
#722680000000
0!
0*
09
0>
0C
#722690000000
1!
1*
b110 6
19
1>
1C
b110 G
#722700000000
0!
0*
09
0>
0C
#722710000000
1!
1*
b111 6
19
1>
1C
b111 G
#722720000000
0!
0*
09
0>
0C
#722730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#722740000000
0!
0*
09
0>
0C
#722750000000
1!
1*
b1 6
19
1>
1C
b1 G
#722760000000
0!
0*
09
0>
0C
#722770000000
1!
1*
b10 6
19
1>
1C
b10 G
#722780000000
0!
0*
09
0>
0C
#722790000000
1!
1*
b11 6
19
1>
1C
b11 G
#722800000000
0!
0*
09
0>
0C
#722810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#722820000000
0!
0*
09
0>
0C
#722830000000
1!
1*
b101 6
19
1>
1C
b101 G
#722840000000
0!
0*
09
0>
0C
#722850000000
1!
1*
b110 6
19
1>
1C
b110 G
#722860000000
0!
0*
09
0>
0C
#722870000000
1!
1*
b111 6
19
1>
1C
b111 G
#722880000000
0!
1"
0*
1+
09
1:
0>
0C
#722890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#722900000000
0!
0*
09
0>
0C
#722910000000
1!
1*
b1 6
19
1>
1C
b1 G
#722920000000
0!
0*
09
0>
0C
#722930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#722940000000
0!
0*
09
0>
0C
#722950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#722960000000
0!
0*
09
0>
0C
#722970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#722980000000
0!
0*
09
0>
0C
#722990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#723000000000
0!
0#
0*
0,
09
0>
0?
0C
#723010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#723020000000
0!
0*
09
0>
0C
#723030000000
1!
1*
19
1>
1C
#723040000000
0!
0*
09
0>
0C
#723050000000
1!
1*
19
1>
1C
#723060000000
0!
0*
09
0>
0C
#723070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#723080000000
0!
0*
09
0>
0C
#723090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#723100000000
0!
0*
09
0>
0C
#723110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#723120000000
0!
0*
09
0>
0C
#723130000000
1!
1*
b10 6
19
1>
1C
b10 G
#723140000000
0!
0*
09
0>
0C
#723150000000
1!
1*
b11 6
19
1>
1C
b11 G
#723160000000
0!
0*
09
0>
0C
#723170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#723180000000
0!
0*
09
0>
0C
#723190000000
1!
1*
b101 6
19
1>
1C
b101 G
#723200000000
0!
0*
09
0>
0C
#723210000000
1!
1*
b110 6
19
1>
1C
b110 G
#723220000000
0!
0*
09
0>
0C
#723230000000
1!
1*
b111 6
19
1>
1C
b111 G
#723240000000
0!
0*
09
0>
0C
#723250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#723260000000
0!
0*
09
0>
0C
#723270000000
1!
1*
b1 6
19
1>
1C
b1 G
#723280000000
0!
0*
09
0>
0C
#723290000000
1!
1*
b10 6
19
1>
1C
b10 G
#723300000000
0!
0*
09
0>
0C
#723310000000
1!
1*
b11 6
19
1>
1C
b11 G
#723320000000
0!
0*
09
0>
0C
#723330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#723340000000
0!
0*
09
0>
0C
#723350000000
1!
1*
b101 6
19
1>
1C
b101 G
#723360000000
0!
0*
09
0>
0C
#723370000000
1!
1*
b110 6
19
1>
1C
b110 G
#723380000000
0!
0*
09
0>
0C
#723390000000
1!
1*
b111 6
19
1>
1C
b111 G
#723400000000
0!
0*
09
0>
0C
#723410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#723420000000
0!
0*
09
0>
0C
#723430000000
1!
1*
b1 6
19
1>
1C
b1 G
#723440000000
0!
0*
09
0>
0C
#723450000000
1!
1*
b10 6
19
1>
1C
b10 G
#723460000000
0!
0*
09
0>
0C
#723470000000
1!
1*
b11 6
19
1>
1C
b11 G
#723480000000
0!
0*
09
0>
0C
#723490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#723500000000
0!
0*
09
0>
0C
#723510000000
1!
1*
b101 6
19
1>
1C
b101 G
#723520000000
0!
0*
09
0>
0C
#723530000000
1!
1*
b110 6
19
1>
1C
b110 G
#723540000000
0!
0*
09
0>
0C
#723550000000
1!
1*
b111 6
19
1>
1C
b111 G
#723560000000
0!
1"
0*
1+
09
1:
0>
0C
#723570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#723580000000
0!
0*
09
0>
0C
#723590000000
1!
1*
b1 6
19
1>
1C
b1 G
#723600000000
0!
0*
09
0>
0C
#723610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#723620000000
0!
0*
09
0>
0C
#723630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#723640000000
0!
0*
09
0>
0C
#723650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#723660000000
0!
0*
09
0>
0C
#723670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#723680000000
0!
0#
0*
0,
09
0>
0?
0C
#723690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#723700000000
0!
0*
09
0>
0C
#723710000000
1!
1*
19
1>
1C
#723720000000
0!
0*
09
0>
0C
#723730000000
1!
1*
19
1>
1C
#723740000000
0!
0*
09
0>
0C
#723750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#723760000000
0!
0*
09
0>
0C
#723770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#723780000000
0!
0*
09
0>
0C
#723790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#723800000000
0!
0*
09
0>
0C
#723810000000
1!
1*
b10 6
19
1>
1C
b10 G
#723820000000
0!
0*
09
0>
0C
#723830000000
1!
1*
b11 6
19
1>
1C
b11 G
#723840000000
0!
0*
09
0>
0C
#723850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#723860000000
0!
0*
09
0>
0C
#723870000000
1!
1*
b101 6
19
1>
1C
b101 G
#723880000000
0!
0*
09
0>
0C
#723890000000
1!
1*
b110 6
19
1>
1C
b110 G
#723900000000
0!
0*
09
0>
0C
#723910000000
1!
1*
b111 6
19
1>
1C
b111 G
#723920000000
0!
0*
09
0>
0C
#723930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#723940000000
0!
0*
09
0>
0C
#723950000000
1!
1*
b1 6
19
1>
1C
b1 G
#723960000000
0!
0*
09
0>
0C
#723970000000
1!
1*
b10 6
19
1>
1C
b10 G
#723980000000
0!
0*
09
0>
0C
#723990000000
1!
1*
b11 6
19
1>
1C
b11 G
#724000000000
0!
0*
09
0>
0C
#724010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#724020000000
0!
0*
09
0>
0C
#724030000000
1!
1*
b101 6
19
1>
1C
b101 G
#724040000000
0!
0*
09
0>
0C
#724050000000
1!
1*
b110 6
19
1>
1C
b110 G
#724060000000
0!
0*
09
0>
0C
#724070000000
1!
1*
b111 6
19
1>
1C
b111 G
#724080000000
0!
0*
09
0>
0C
#724090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#724100000000
0!
0*
09
0>
0C
#724110000000
1!
1*
b1 6
19
1>
1C
b1 G
#724120000000
0!
0*
09
0>
0C
#724130000000
1!
1*
b10 6
19
1>
1C
b10 G
#724140000000
0!
0*
09
0>
0C
#724150000000
1!
1*
b11 6
19
1>
1C
b11 G
#724160000000
0!
0*
09
0>
0C
#724170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#724180000000
0!
0*
09
0>
0C
#724190000000
1!
1*
b101 6
19
1>
1C
b101 G
#724200000000
0!
0*
09
0>
0C
#724210000000
1!
1*
b110 6
19
1>
1C
b110 G
#724220000000
0!
0*
09
0>
0C
#724230000000
1!
1*
b111 6
19
1>
1C
b111 G
#724240000000
0!
1"
0*
1+
09
1:
0>
0C
#724250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#724260000000
0!
0*
09
0>
0C
#724270000000
1!
1*
b1 6
19
1>
1C
b1 G
#724280000000
0!
0*
09
0>
0C
#724290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#724300000000
0!
0*
09
0>
0C
#724310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#724320000000
0!
0*
09
0>
0C
#724330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#724340000000
0!
0*
09
0>
0C
#724350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#724360000000
0!
0#
0*
0,
09
0>
0?
0C
#724370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#724380000000
0!
0*
09
0>
0C
#724390000000
1!
1*
19
1>
1C
#724400000000
0!
0*
09
0>
0C
#724410000000
1!
1*
19
1>
1C
#724420000000
0!
0*
09
0>
0C
#724430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#724440000000
0!
0*
09
0>
0C
#724450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#724460000000
0!
0*
09
0>
0C
#724470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#724480000000
0!
0*
09
0>
0C
#724490000000
1!
1*
b10 6
19
1>
1C
b10 G
#724500000000
0!
0*
09
0>
0C
#724510000000
1!
1*
b11 6
19
1>
1C
b11 G
#724520000000
0!
0*
09
0>
0C
#724530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#724540000000
0!
0*
09
0>
0C
#724550000000
1!
1*
b101 6
19
1>
1C
b101 G
#724560000000
0!
0*
09
0>
0C
#724570000000
1!
1*
b110 6
19
1>
1C
b110 G
#724580000000
0!
0*
09
0>
0C
#724590000000
1!
1*
b111 6
19
1>
1C
b111 G
#724600000000
0!
0*
09
0>
0C
#724610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#724620000000
0!
0*
09
0>
0C
#724630000000
1!
1*
b1 6
19
1>
1C
b1 G
#724640000000
0!
0*
09
0>
0C
#724650000000
1!
1*
b10 6
19
1>
1C
b10 G
#724660000000
0!
0*
09
0>
0C
#724670000000
1!
1*
b11 6
19
1>
1C
b11 G
#724680000000
0!
0*
09
0>
0C
#724690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#724700000000
0!
0*
09
0>
0C
#724710000000
1!
1*
b101 6
19
1>
1C
b101 G
#724720000000
0!
0*
09
0>
0C
#724730000000
1!
1*
b110 6
19
1>
1C
b110 G
#724740000000
0!
0*
09
0>
0C
#724750000000
1!
1*
b111 6
19
1>
1C
b111 G
#724760000000
0!
0*
09
0>
0C
#724770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#724780000000
0!
0*
09
0>
0C
#724790000000
1!
1*
b1 6
19
1>
1C
b1 G
#724800000000
0!
0*
09
0>
0C
#724810000000
1!
1*
b10 6
19
1>
1C
b10 G
#724820000000
0!
0*
09
0>
0C
#724830000000
1!
1*
b11 6
19
1>
1C
b11 G
#724840000000
0!
0*
09
0>
0C
#724850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#724860000000
0!
0*
09
0>
0C
#724870000000
1!
1*
b101 6
19
1>
1C
b101 G
#724880000000
0!
0*
09
0>
0C
#724890000000
1!
1*
b110 6
19
1>
1C
b110 G
#724900000000
0!
0*
09
0>
0C
#724910000000
1!
1*
b111 6
19
1>
1C
b111 G
#724920000000
0!
1"
0*
1+
09
1:
0>
0C
#724930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#724940000000
0!
0*
09
0>
0C
#724950000000
1!
1*
b1 6
19
1>
1C
b1 G
#724960000000
0!
0*
09
0>
0C
#724970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#724980000000
0!
0*
09
0>
0C
#724990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#725000000000
0!
0*
09
0>
0C
#725010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#725020000000
0!
0*
09
0>
0C
#725030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#725040000000
0!
0#
0*
0,
09
0>
0?
0C
#725050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#725060000000
0!
0*
09
0>
0C
#725070000000
1!
1*
19
1>
1C
#725080000000
0!
0*
09
0>
0C
#725090000000
1!
1*
19
1>
1C
#725100000000
0!
0*
09
0>
0C
#725110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#725120000000
0!
0*
09
0>
0C
#725130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#725140000000
0!
0*
09
0>
0C
#725150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#725160000000
0!
0*
09
0>
0C
#725170000000
1!
1*
b10 6
19
1>
1C
b10 G
#725180000000
0!
0*
09
0>
0C
#725190000000
1!
1*
b11 6
19
1>
1C
b11 G
#725200000000
0!
0*
09
0>
0C
#725210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#725220000000
0!
0*
09
0>
0C
#725230000000
1!
1*
b101 6
19
1>
1C
b101 G
#725240000000
0!
0*
09
0>
0C
#725250000000
1!
1*
b110 6
19
1>
1C
b110 G
#725260000000
0!
0*
09
0>
0C
#725270000000
1!
1*
b111 6
19
1>
1C
b111 G
#725280000000
0!
0*
09
0>
0C
#725290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#725300000000
0!
0*
09
0>
0C
#725310000000
1!
1*
b1 6
19
1>
1C
b1 G
#725320000000
0!
0*
09
0>
0C
#725330000000
1!
1*
b10 6
19
1>
1C
b10 G
#725340000000
0!
0*
09
0>
0C
#725350000000
1!
1*
b11 6
19
1>
1C
b11 G
#725360000000
0!
0*
09
0>
0C
#725370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#725380000000
0!
0*
09
0>
0C
#725390000000
1!
1*
b101 6
19
1>
1C
b101 G
#725400000000
0!
0*
09
0>
0C
#725410000000
1!
1*
b110 6
19
1>
1C
b110 G
#725420000000
0!
0*
09
0>
0C
#725430000000
1!
1*
b111 6
19
1>
1C
b111 G
#725440000000
0!
0*
09
0>
0C
#725450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#725460000000
0!
0*
09
0>
0C
#725470000000
1!
1*
b1 6
19
1>
1C
b1 G
#725480000000
0!
0*
09
0>
0C
#725490000000
1!
1*
b10 6
19
1>
1C
b10 G
#725500000000
0!
0*
09
0>
0C
#725510000000
1!
1*
b11 6
19
1>
1C
b11 G
#725520000000
0!
0*
09
0>
0C
#725530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#725540000000
0!
0*
09
0>
0C
#725550000000
1!
1*
b101 6
19
1>
1C
b101 G
#725560000000
0!
0*
09
0>
0C
#725570000000
1!
1*
b110 6
19
1>
1C
b110 G
#725580000000
0!
0*
09
0>
0C
#725590000000
1!
1*
b111 6
19
1>
1C
b111 G
#725600000000
0!
1"
0*
1+
09
1:
0>
0C
#725610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#725620000000
0!
0*
09
0>
0C
#725630000000
1!
1*
b1 6
19
1>
1C
b1 G
#725640000000
0!
0*
09
0>
0C
#725650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#725660000000
0!
0*
09
0>
0C
#725670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#725680000000
0!
0*
09
0>
0C
#725690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#725700000000
0!
0*
09
0>
0C
#725710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#725720000000
0!
0#
0*
0,
09
0>
0?
0C
#725730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#725740000000
0!
0*
09
0>
0C
#725750000000
1!
1*
19
1>
1C
#725760000000
0!
0*
09
0>
0C
#725770000000
1!
1*
19
1>
1C
#725780000000
0!
0*
09
0>
0C
#725790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#725800000000
0!
0*
09
0>
0C
#725810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#725820000000
0!
0*
09
0>
0C
#725830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#725840000000
0!
0*
09
0>
0C
#725850000000
1!
1*
b10 6
19
1>
1C
b10 G
#725860000000
0!
0*
09
0>
0C
#725870000000
1!
1*
b11 6
19
1>
1C
b11 G
#725880000000
0!
0*
09
0>
0C
#725890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#725900000000
0!
0*
09
0>
0C
#725910000000
1!
1*
b101 6
19
1>
1C
b101 G
#725920000000
0!
0*
09
0>
0C
#725930000000
1!
1*
b110 6
19
1>
1C
b110 G
#725940000000
0!
0*
09
0>
0C
#725950000000
1!
1*
b111 6
19
1>
1C
b111 G
#725960000000
0!
0*
09
0>
0C
#725970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#725980000000
0!
0*
09
0>
0C
#725990000000
1!
1*
b1 6
19
1>
1C
b1 G
#726000000000
0!
0*
09
0>
0C
#726010000000
1!
1*
b10 6
19
1>
1C
b10 G
#726020000000
0!
0*
09
0>
0C
#726030000000
1!
1*
b11 6
19
1>
1C
b11 G
#726040000000
0!
0*
09
0>
0C
#726050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#726060000000
0!
0*
09
0>
0C
#726070000000
1!
1*
b101 6
19
1>
1C
b101 G
#726080000000
0!
0*
09
0>
0C
#726090000000
1!
1*
b110 6
19
1>
1C
b110 G
#726100000000
0!
0*
09
0>
0C
#726110000000
1!
1*
b111 6
19
1>
1C
b111 G
#726120000000
0!
0*
09
0>
0C
#726130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#726140000000
0!
0*
09
0>
0C
#726150000000
1!
1*
b1 6
19
1>
1C
b1 G
#726160000000
0!
0*
09
0>
0C
#726170000000
1!
1*
b10 6
19
1>
1C
b10 G
#726180000000
0!
0*
09
0>
0C
#726190000000
1!
1*
b11 6
19
1>
1C
b11 G
#726200000000
0!
0*
09
0>
0C
#726210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#726220000000
0!
0*
09
0>
0C
#726230000000
1!
1*
b101 6
19
1>
1C
b101 G
#726240000000
0!
0*
09
0>
0C
#726250000000
1!
1*
b110 6
19
1>
1C
b110 G
#726260000000
0!
0*
09
0>
0C
#726270000000
1!
1*
b111 6
19
1>
1C
b111 G
#726280000000
0!
1"
0*
1+
09
1:
0>
0C
#726290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#726300000000
0!
0*
09
0>
0C
#726310000000
1!
1*
b1 6
19
1>
1C
b1 G
#726320000000
0!
0*
09
0>
0C
#726330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#726340000000
0!
0*
09
0>
0C
#726350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#726360000000
0!
0*
09
0>
0C
#726370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#726380000000
0!
0*
09
0>
0C
#726390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#726400000000
0!
0#
0*
0,
09
0>
0?
0C
#726410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#726420000000
0!
0*
09
0>
0C
#726430000000
1!
1*
19
1>
1C
#726440000000
0!
0*
09
0>
0C
#726450000000
1!
1*
19
1>
1C
#726460000000
0!
0*
09
0>
0C
#726470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#726480000000
0!
0*
09
0>
0C
#726490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#726500000000
0!
0*
09
0>
0C
#726510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#726520000000
0!
0*
09
0>
0C
#726530000000
1!
1*
b10 6
19
1>
1C
b10 G
#726540000000
0!
0*
09
0>
0C
#726550000000
1!
1*
b11 6
19
1>
1C
b11 G
#726560000000
0!
0*
09
0>
0C
#726570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#726580000000
0!
0*
09
0>
0C
#726590000000
1!
1*
b101 6
19
1>
1C
b101 G
#726600000000
0!
0*
09
0>
0C
#726610000000
1!
1*
b110 6
19
1>
1C
b110 G
#726620000000
0!
0*
09
0>
0C
#726630000000
1!
1*
b111 6
19
1>
1C
b111 G
#726640000000
0!
0*
09
0>
0C
#726650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#726660000000
0!
0*
09
0>
0C
#726670000000
1!
1*
b1 6
19
1>
1C
b1 G
#726680000000
0!
0*
09
0>
0C
#726690000000
1!
1*
b10 6
19
1>
1C
b10 G
#726700000000
0!
0*
09
0>
0C
#726710000000
1!
1*
b11 6
19
1>
1C
b11 G
#726720000000
0!
0*
09
0>
0C
#726730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#726740000000
0!
0*
09
0>
0C
#726750000000
1!
1*
b101 6
19
1>
1C
b101 G
#726760000000
0!
0*
09
0>
0C
#726770000000
1!
1*
b110 6
19
1>
1C
b110 G
#726780000000
0!
0*
09
0>
0C
#726790000000
1!
1*
b111 6
19
1>
1C
b111 G
#726800000000
0!
0*
09
0>
0C
#726810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#726820000000
0!
0*
09
0>
0C
#726830000000
1!
1*
b1 6
19
1>
1C
b1 G
#726840000000
0!
0*
09
0>
0C
#726850000000
1!
1*
b10 6
19
1>
1C
b10 G
#726860000000
0!
0*
09
0>
0C
#726870000000
1!
1*
b11 6
19
1>
1C
b11 G
#726880000000
0!
0*
09
0>
0C
#726890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#726900000000
0!
0*
09
0>
0C
#726910000000
1!
1*
b101 6
19
1>
1C
b101 G
#726920000000
0!
0*
09
0>
0C
#726930000000
1!
1*
b110 6
19
1>
1C
b110 G
#726940000000
0!
0*
09
0>
0C
#726950000000
1!
1*
b111 6
19
1>
1C
b111 G
#726960000000
0!
1"
0*
1+
09
1:
0>
0C
#726970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#726980000000
0!
0*
09
0>
0C
#726990000000
1!
1*
b1 6
19
1>
1C
b1 G
#727000000000
0!
0*
09
0>
0C
#727010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#727020000000
0!
0*
09
0>
0C
#727030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#727040000000
0!
0*
09
0>
0C
#727050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#727060000000
0!
0*
09
0>
0C
#727070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#727080000000
0!
0#
0*
0,
09
0>
0?
0C
#727090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#727100000000
0!
0*
09
0>
0C
#727110000000
1!
1*
19
1>
1C
#727120000000
0!
0*
09
0>
0C
#727130000000
1!
1*
19
1>
1C
#727140000000
0!
0*
09
0>
0C
#727150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#727160000000
0!
0*
09
0>
0C
#727170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#727180000000
0!
0*
09
0>
0C
#727190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#727200000000
0!
0*
09
0>
0C
#727210000000
1!
1*
b10 6
19
1>
1C
b10 G
#727220000000
0!
0*
09
0>
0C
#727230000000
1!
1*
b11 6
19
1>
1C
b11 G
#727240000000
0!
0*
09
0>
0C
#727250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#727260000000
0!
0*
09
0>
0C
#727270000000
1!
1*
b101 6
19
1>
1C
b101 G
#727280000000
0!
0*
09
0>
0C
#727290000000
1!
1*
b110 6
19
1>
1C
b110 G
#727300000000
0!
0*
09
0>
0C
#727310000000
1!
1*
b111 6
19
1>
1C
b111 G
#727320000000
0!
0*
09
0>
0C
#727330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#727340000000
0!
0*
09
0>
0C
#727350000000
1!
1*
b1 6
19
1>
1C
b1 G
#727360000000
0!
0*
09
0>
0C
#727370000000
1!
1*
b10 6
19
1>
1C
b10 G
#727380000000
0!
0*
09
0>
0C
#727390000000
1!
1*
b11 6
19
1>
1C
b11 G
#727400000000
0!
0*
09
0>
0C
#727410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#727420000000
0!
0*
09
0>
0C
#727430000000
1!
1*
b101 6
19
1>
1C
b101 G
#727440000000
0!
0*
09
0>
0C
#727450000000
1!
1*
b110 6
19
1>
1C
b110 G
#727460000000
0!
0*
09
0>
0C
#727470000000
1!
1*
b111 6
19
1>
1C
b111 G
#727480000000
0!
0*
09
0>
0C
#727490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#727500000000
0!
0*
09
0>
0C
#727510000000
1!
1*
b1 6
19
1>
1C
b1 G
#727520000000
0!
0*
09
0>
0C
#727530000000
1!
1*
b10 6
19
1>
1C
b10 G
#727540000000
0!
0*
09
0>
0C
#727550000000
1!
1*
b11 6
19
1>
1C
b11 G
#727560000000
0!
0*
09
0>
0C
#727570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#727580000000
0!
0*
09
0>
0C
#727590000000
1!
1*
b101 6
19
1>
1C
b101 G
#727600000000
0!
0*
09
0>
0C
#727610000000
1!
1*
b110 6
19
1>
1C
b110 G
#727620000000
0!
0*
09
0>
0C
#727630000000
1!
1*
b111 6
19
1>
1C
b111 G
#727640000000
0!
1"
0*
1+
09
1:
0>
0C
#727650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#727660000000
0!
0*
09
0>
0C
#727670000000
1!
1*
b1 6
19
1>
1C
b1 G
#727680000000
0!
0*
09
0>
0C
#727690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#727700000000
0!
0*
09
0>
0C
#727710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#727720000000
0!
0*
09
0>
0C
#727730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#727740000000
0!
0*
09
0>
0C
#727750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#727760000000
0!
0#
0*
0,
09
0>
0?
0C
#727770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#727780000000
0!
0*
09
0>
0C
#727790000000
1!
1*
19
1>
1C
#727800000000
0!
0*
09
0>
0C
#727810000000
1!
1*
19
1>
1C
#727820000000
0!
0*
09
0>
0C
#727830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#727840000000
0!
0*
09
0>
0C
#727850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#727860000000
0!
0*
09
0>
0C
#727870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#727880000000
0!
0*
09
0>
0C
#727890000000
1!
1*
b10 6
19
1>
1C
b10 G
#727900000000
0!
0*
09
0>
0C
#727910000000
1!
1*
b11 6
19
1>
1C
b11 G
#727920000000
0!
0*
09
0>
0C
#727930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#727940000000
0!
0*
09
0>
0C
#727950000000
1!
1*
b101 6
19
1>
1C
b101 G
#727960000000
0!
0*
09
0>
0C
#727970000000
1!
1*
b110 6
19
1>
1C
b110 G
#727980000000
0!
0*
09
0>
0C
#727990000000
1!
1*
b111 6
19
1>
1C
b111 G
#728000000000
0!
0*
09
0>
0C
#728010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#728020000000
0!
0*
09
0>
0C
#728030000000
1!
1*
b1 6
19
1>
1C
b1 G
#728040000000
0!
0*
09
0>
0C
#728050000000
1!
1*
b10 6
19
1>
1C
b10 G
#728060000000
0!
0*
09
0>
0C
#728070000000
1!
1*
b11 6
19
1>
1C
b11 G
#728080000000
0!
0*
09
0>
0C
#728090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#728100000000
0!
0*
09
0>
0C
#728110000000
1!
1*
b101 6
19
1>
1C
b101 G
#728120000000
0!
0*
09
0>
0C
#728130000000
1!
1*
b110 6
19
1>
1C
b110 G
#728140000000
0!
0*
09
0>
0C
#728150000000
1!
1*
b111 6
19
1>
1C
b111 G
#728160000000
0!
0*
09
0>
0C
#728170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#728180000000
0!
0*
09
0>
0C
#728190000000
1!
1*
b1 6
19
1>
1C
b1 G
#728200000000
0!
0*
09
0>
0C
#728210000000
1!
1*
b10 6
19
1>
1C
b10 G
#728220000000
0!
0*
09
0>
0C
#728230000000
1!
1*
b11 6
19
1>
1C
b11 G
#728240000000
0!
0*
09
0>
0C
#728250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#728260000000
0!
0*
09
0>
0C
#728270000000
1!
1*
b101 6
19
1>
1C
b101 G
#728280000000
0!
0*
09
0>
0C
#728290000000
1!
1*
b110 6
19
1>
1C
b110 G
#728300000000
0!
0*
09
0>
0C
#728310000000
1!
1*
b111 6
19
1>
1C
b111 G
#728320000000
0!
1"
0*
1+
09
1:
0>
0C
#728330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#728340000000
0!
0*
09
0>
0C
#728350000000
1!
1*
b1 6
19
1>
1C
b1 G
#728360000000
0!
0*
09
0>
0C
#728370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#728380000000
0!
0*
09
0>
0C
#728390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#728400000000
0!
0*
09
0>
0C
#728410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#728420000000
0!
0*
09
0>
0C
#728430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#728440000000
0!
0#
0*
0,
09
0>
0?
0C
#728450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#728460000000
0!
0*
09
0>
0C
#728470000000
1!
1*
19
1>
1C
#728480000000
0!
0*
09
0>
0C
#728490000000
1!
1*
19
1>
1C
#728500000000
0!
0*
09
0>
0C
#728510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#728520000000
0!
0*
09
0>
0C
#728530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#728540000000
0!
0*
09
0>
0C
#728550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#728560000000
0!
0*
09
0>
0C
#728570000000
1!
1*
b10 6
19
1>
1C
b10 G
#728580000000
0!
0*
09
0>
0C
#728590000000
1!
1*
b11 6
19
1>
1C
b11 G
#728600000000
0!
0*
09
0>
0C
#728610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#728620000000
0!
0*
09
0>
0C
#728630000000
1!
1*
b101 6
19
1>
1C
b101 G
#728640000000
0!
0*
09
0>
0C
#728650000000
1!
1*
b110 6
19
1>
1C
b110 G
#728660000000
0!
0*
09
0>
0C
#728670000000
1!
1*
b111 6
19
1>
1C
b111 G
#728680000000
0!
0*
09
0>
0C
#728690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#728700000000
0!
0*
09
0>
0C
#728710000000
1!
1*
b1 6
19
1>
1C
b1 G
#728720000000
0!
0*
09
0>
0C
#728730000000
1!
1*
b10 6
19
1>
1C
b10 G
#728740000000
0!
0*
09
0>
0C
#728750000000
1!
1*
b11 6
19
1>
1C
b11 G
#728760000000
0!
0*
09
0>
0C
#728770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#728780000000
0!
0*
09
0>
0C
#728790000000
1!
1*
b101 6
19
1>
1C
b101 G
#728800000000
0!
0*
09
0>
0C
#728810000000
1!
1*
b110 6
19
1>
1C
b110 G
#728820000000
0!
0*
09
0>
0C
#728830000000
1!
1*
b111 6
19
1>
1C
b111 G
#728840000000
0!
0*
09
0>
0C
#728850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#728860000000
0!
0*
09
0>
0C
#728870000000
1!
1*
b1 6
19
1>
1C
b1 G
#728880000000
0!
0*
09
0>
0C
#728890000000
1!
1*
b10 6
19
1>
1C
b10 G
#728900000000
0!
0*
09
0>
0C
#728910000000
1!
1*
b11 6
19
1>
1C
b11 G
#728920000000
0!
0*
09
0>
0C
#728930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#728940000000
0!
0*
09
0>
0C
#728950000000
1!
1*
b101 6
19
1>
1C
b101 G
#728960000000
0!
0*
09
0>
0C
#728970000000
1!
1*
b110 6
19
1>
1C
b110 G
#728980000000
0!
0*
09
0>
0C
#728990000000
1!
1*
b111 6
19
1>
1C
b111 G
#729000000000
0!
1"
0*
1+
09
1:
0>
0C
#729010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#729020000000
0!
0*
09
0>
0C
#729030000000
1!
1*
b1 6
19
1>
1C
b1 G
#729040000000
0!
0*
09
0>
0C
#729050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#729060000000
0!
0*
09
0>
0C
#729070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#729080000000
0!
0*
09
0>
0C
#729090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#729100000000
0!
0*
09
0>
0C
#729110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#729120000000
0!
0#
0*
0,
09
0>
0?
0C
#729130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#729140000000
0!
0*
09
0>
0C
#729150000000
1!
1*
19
1>
1C
#729160000000
0!
0*
09
0>
0C
#729170000000
1!
1*
19
1>
1C
#729180000000
0!
0*
09
0>
0C
#729190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#729200000000
0!
0*
09
0>
0C
#729210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#729220000000
0!
0*
09
0>
0C
#729230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#729240000000
0!
0*
09
0>
0C
#729250000000
1!
1*
b10 6
19
1>
1C
b10 G
#729260000000
0!
0*
09
0>
0C
#729270000000
1!
1*
b11 6
19
1>
1C
b11 G
#729280000000
0!
0*
09
0>
0C
#729290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#729300000000
0!
0*
09
0>
0C
#729310000000
1!
1*
b101 6
19
1>
1C
b101 G
#729320000000
0!
0*
09
0>
0C
#729330000000
1!
1*
b110 6
19
1>
1C
b110 G
#729340000000
0!
0*
09
0>
0C
#729350000000
1!
1*
b111 6
19
1>
1C
b111 G
#729360000000
0!
0*
09
0>
0C
#729370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#729380000000
0!
0*
09
0>
0C
#729390000000
1!
1*
b1 6
19
1>
1C
b1 G
#729400000000
0!
0*
09
0>
0C
#729410000000
1!
1*
b10 6
19
1>
1C
b10 G
#729420000000
0!
0*
09
0>
0C
#729430000000
1!
1*
b11 6
19
1>
1C
b11 G
#729440000000
0!
0*
09
0>
0C
#729450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#729460000000
0!
0*
09
0>
0C
#729470000000
1!
1*
b101 6
19
1>
1C
b101 G
#729480000000
0!
0*
09
0>
0C
#729490000000
1!
1*
b110 6
19
1>
1C
b110 G
#729500000000
0!
0*
09
0>
0C
#729510000000
1!
1*
b111 6
19
1>
1C
b111 G
#729520000000
0!
0*
09
0>
0C
#729530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#729540000000
0!
0*
09
0>
0C
#729550000000
1!
1*
b1 6
19
1>
1C
b1 G
#729560000000
0!
0*
09
0>
0C
#729570000000
1!
1*
b10 6
19
1>
1C
b10 G
#729580000000
0!
0*
09
0>
0C
#729590000000
1!
1*
b11 6
19
1>
1C
b11 G
#729600000000
0!
0*
09
0>
0C
#729610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#729620000000
0!
0*
09
0>
0C
#729630000000
1!
1*
b101 6
19
1>
1C
b101 G
#729640000000
0!
0*
09
0>
0C
#729650000000
1!
1*
b110 6
19
1>
1C
b110 G
#729660000000
0!
0*
09
0>
0C
#729670000000
1!
1*
b111 6
19
1>
1C
b111 G
#729680000000
0!
1"
0*
1+
09
1:
0>
0C
#729690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#729700000000
0!
0*
09
0>
0C
#729710000000
1!
1*
b1 6
19
1>
1C
b1 G
#729720000000
0!
0*
09
0>
0C
#729730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#729740000000
0!
0*
09
0>
0C
#729750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#729760000000
0!
0*
09
0>
0C
#729770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#729780000000
0!
0*
09
0>
0C
#729790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#729800000000
0!
0#
0*
0,
09
0>
0?
0C
#729810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#729820000000
0!
0*
09
0>
0C
#729830000000
1!
1*
19
1>
1C
#729840000000
0!
0*
09
0>
0C
#729850000000
1!
1*
19
1>
1C
#729860000000
0!
0*
09
0>
0C
#729870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#729880000000
0!
0*
09
0>
0C
#729890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#729900000000
0!
0*
09
0>
0C
#729910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#729920000000
0!
0*
09
0>
0C
#729930000000
1!
1*
b10 6
19
1>
1C
b10 G
#729940000000
0!
0*
09
0>
0C
#729950000000
1!
1*
b11 6
19
1>
1C
b11 G
#729960000000
0!
0*
09
0>
0C
#729970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#729980000000
0!
0*
09
0>
0C
#729990000000
1!
1*
b101 6
19
1>
1C
b101 G
#730000000000
0!
0*
09
0>
0C
#730010000000
1!
1*
b110 6
19
1>
1C
b110 G
#730020000000
0!
0*
09
0>
0C
#730030000000
1!
1*
b111 6
19
1>
1C
b111 G
#730040000000
0!
0*
09
0>
0C
#730050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#730060000000
0!
0*
09
0>
0C
#730070000000
1!
1*
b1 6
19
1>
1C
b1 G
#730080000000
0!
0*
09
0>
0C
#730090000000
1!
1*
b10 6
19
1>
1C
b10 G
#730100000000
0!
0*
09
0>
0C
#730110000000
1!
1*
b11 6
19
1>
1C
b11 G
#730120000000
0!
0*
09
0>
0C
#730130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#730140000000
0!
0*
09
0>
0C
#730150000000
1!
1*
b101 6
19
1>
1C
b101 G
#730160000000
0!
0*
09
0>
0C
#730170000000
1!
1*
b110 6
19
1>
1C
b110 G
#730180000000
0!
0*
09
0>
0C
#730190000000
1!
1*
b111 6
19
1>
1C
b111 G
#730200000000
0!
0*
09
0>
0C
#730210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#730220000000
0!
0*
09
0>
0C
#730230000000
1!
1*
b1 6
19
1>
1C
b1 G
#730240000000
0!
0*
09
0>
0C
#730250000000
1!
1*
b10 6
19
1>
1C
b10 G
#730260000000
0!
0*
09
0>
0C
#730270000000
1!
1*
b11 6
19
1>
1C
b11 G
#730280000000
0!
0*
09
0>
0C
#730290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#730300000000
0!
0*
09
0>
0C
#730310000000
1!
1*
b101 6
19
1>
1C
b101 G
#730320000000
0!
0*
09
0>
0C
#730330000000
1!
1*
b110 6
19
1>
1C
b110 G
#730340000000
0!
0*
09
0>
0C
#730350000000
1!
1*
b111 6
19
1>
1C
b111 G
#730360000000
0!
1"
0*
1+
09
1:
0>
0C
#730370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#730380000000
0!
0*
09
0>
0C
#730390000000
1!
1*
b1 6
19
1>
1C
b1 G
#730400000000
0!
0*
09
0>
0C
#730410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#730420000000
0!
0*
09
0>
0C
#730430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#730440000000
0!
0*
09
0>
0C
#730450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#730460000000
0!
0*
09
0>
0C
#730470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#730480000000
0!
0#
0*
0,
09
0>
0?
0C
#730490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#730500000000
0!
0*
09
0>
0C
#730510000000
1!
1*
19
1>
1C
#730520000000
0!
0*
09
0>
0C
#730530000000
1!
1*
19
1>
1C
#730540000000
0!
0*
09
0>
0C
#730550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#730560000000
0!
0*
09
0>
0C
#730570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#730580000000
0!
0*
09
0>
0C
#730590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#730600000000
0!
0*
09
0>
0C
#730610000000
1!
1*
b10 6
19
1>
1C
b10 G
#730620000000
0!
0*
09
0>
0C
#730630000000
1!
1*
b11 6
19
1>
1C
b11 G
#730640000000
0!
0*
09
0>
0C
#730650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#730660000000
0!
0*
09
0>
0C
#730670000000
1!
1*
b101 6
19
1>
1C
b101 G
#730680000000
0!
0*
09
0>
0C
#730690000000
1!
1*
b110 6
19
1>
1C
b110 G
#730700000000
0!
0*
09
0>
0C
#730710000000
1!
1*
b111 6
19
1>
1C
b111 G
#730720000000
0!
0*
09
0>
0C
#730730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#730740000000
0!
0*
09
0>
0C
#730750000000
1!
1*
b1 6
19
1>
1C
b1 G
#730760000000
0!
0*
09
0>
0C
#730770000000
1!
1*
b10 6
19
1>
1C
b10 G
#730780000000
0!
0*
09
0>
0C
#730790000000
1!
1*
b11 6
19
1>
1C
b11 G
#730800000000
0!
0*
09
0>
0C
#730810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#730820000000
0!
0*
09
0>
0C
#730830000000
1!
1*
b101 6
19
1>
1C
b101 G
#730840000000
0!
0*
09
0>
0C
#730850000000
1!
1*
b110 6
19
1>
1C
b110 G
#730860000000
0!
0*
09
0>
0C
#730870000000
1!
1*
b111 6
19
1>
1C
b111 G
#730880000000
0!
0*
09
0>
0C
#730890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#730900000000
0!
0*
09
0>
0C
#730910000000
1!
1*
b1 6
19
1>
1C
b1 G
#730920000000
0!
0*
09
0>
0C
#730930000000
1!
1*
b10 6
19
1>
1C
b10 G
#730940000000
0!
0*
09
0>
0C
#730950000000
1!
1*
b11 6
19
1>
1C
b11 G
#730960000000
0!
0*
09
0>
0C
#730970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#730980000000
0!
0*
09
0>
0C
#730990000000
1!
1*
b101 6
19
1>
1C
b101 G
#731000000000
0!
0*
09
0>
0C
#731010000000
1!
1*
b110 6
19
1>
1C
b110 G
#731020000000
0!
0*
09
0>
0C
#731030000000
1!
1*
b111 6
19
1>
1C
b111 G
#731040000000
0!
1"
0*
1+
09
1:
0>
0C
#731050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#731060000000
0!
0*
09
0>
0C
#731070000000
1!
1*
b1 6
19
1>
1C
b1 G
#731080000000
0!
0*
09
0>
0C
#731090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#731100000000
0!
0*
09
0>
0C
#731110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#731120000000
0!
0*
09
0>
0C
#731130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#731140000000
0!
0*
09
0>
0C
#731150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#731160000000
0!
0#
0*
0,
09
0>
0?
0C
#731170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#731180000000
0!
0*
09
0>
0C
#731190000000
1!
1*
19
1>
1C
#731200000000
0!
0*
09
0>
0C
#731210000000
1!
1*
19
1>
1C
#731220000000
0!
0*
09
0>
0C
#731230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#731240000000
0!
0*
09
0>
0C
#731250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#731260000000
0!
0*
09
0>
0C
#731270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#731280000000
0!
0*
09
0>
0C
#731290000000
1!
1*
b10 6
19
1>
1C
b10 G
#731300000000
0!
0*
09
0>
0C
#731310000000
1!
1*
b11 6
19
1>
1C
b11 G
#731320000000
0!
0*
09
0>
0C
#731330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#731340000000
0!
0*
09
0>
0C
#731350000000
1!
1*
b101 6
19
1>
1C
b101 G
#731360000000
0!
0*
09
0>
0C
#731370000000
1!
1*
b110 6
19
1>
1C
b110 G
#731380000000
0!
0*
09
0>
0C
#731390000000
1!
1*
b111 6
19
1>
1C
b111 G
#731400000000
0!
0*
09
0>
0C
#731410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#731420000000
0!
0*
09
0>
0C
#731430000000
1!
1*
b1 6
19
1>
1C
b1 G
#731440000000
0!
0*
09
0>
0C
#731450000000
1!
1*
b10 6
19
1>
1C
b10 G
#731460000000
0!
0*
09
0>
0C
#731470000000
1!
1*
b11 6
19
1>
1C
b11 G
#731480000000
0!
0*
09
0>
0C
#731490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#731500000000
0!
0*
09
0>
0C
#731510000000
1!
1*
b101 6
19
1>
1C
b101 G
#731520000000
0!
0*
09
0>
0C
#731530000000
1!
1*
b110 6
19
1>
1C
b110 G
#731540000000
0!
0*
09
0>
0C
#731550000000
1!
1*
b111 6
19
1>
1C
b111 G
#731560000000
0!
0*
09
0>
0C
#731570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#731580000000
0!
0*
09
0>
0C
#731590000000
1!
1*
b1 6
19
1>
1C
b1 G
#731600000000
0!
0*
09
0>
0C
#731610000000
1!
1*
b10 6
19
1>
1C
b10 G
#731620000000
0!
0*
09
0>
0C
#731630000000
1!
1*
b11 6
19
1>
1C
b11 G
#731640000000
0!
0*
09
0>
0C
#731650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#731660000000
0!
0*
09
0>
0C
#731670000000
1!
1*
b101 6
19
1>
1C
b101 G
#731680000000
0!
0*
09
0>
0C
#731690000000
1!
1*
b110 6
19
1>
1C
b110 G
#731700000000
0!
0*
09
0>
0C
#731710000000
1!
1*
b111 6
19
1>
1C
b111 G
#731720000000
0!
1"
0*
1+
09
1:
0>
0C
#731730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#731740000000
0!
0*
09
0>
0C
#731750000000
1!
1*
b1 6
19
1>
1C
b1 G
#731760000000
0!
0*
09
0>
0C
#731770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#731780000000
0!
0*
09
0>
0C
#731790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#731800000000
0!
0*
09
0>
0C
#731810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#731820000000
0!
0*
09
0>
0C
#731830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#731840000000
0!
0#
0*
0,
09
0>
0?
0C
#731850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#731860000000
0!
0*
09
0>
0C
#731870000000
1!
1*
19
1>
1C
#731880000000
0!
0*
09
0>
0C
#731890000000
1!
1*
19
1>
1C
#731900000000
0!
0*
09
0>
0C
#731910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#731920000000
0!
0*
09
0>
0C
#731930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#731940000000
0!
0*
09
0>
0C
#731950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#731960000000
0!
0*
09
0>
0C
#731970000000
1!
1*
b10 6
19
1>
1C
b10 G
#731980000000
0!
0*
09
0>
0C
#731990000000
1!
1*
b11 6
19
1>
1C
b11 G
#732000000000
0!
0*
09
0>
0C
#732010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#732020000000
0!
0*
09
0>
0C
#732030000000
1!
1*
b101 6
19
1>
1C
b101 G
#732040000000
0!
0*
09
0>
0C
#732050000000
1!
1*
b110 6
19
1>
1C
b110 G
#732060000000
0!
0*
09
0>
0C
#732070000000
1!
1*
b111 6
19
1>
1C
b111 G
#732080000000
0!
0*
09
0>
0C
#732090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#732100000000
0!
0*
09
0>
0C
#732110000000
1!
1*
b1 6
19
1>
1C
b1 G
#732120000000
0!
0*
09
0>
0C
#732130000000
1!
1*
b10 6
19
1>
1C
b10 G
#732140000000
0!
0*
09
0>
0C
#732150000000
1!
1*
b11 6
19
1>
1C
b11 G
#732160000000
0!
0*
09
0>
0C
#732170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#732180000000
0!
0*
09
0>
0C
#732190000000
1!
1*
b101 6
19
1>
1C
b101 G
#732200000000
0!
0*
09
0>
0C
#732210000000
1!
1*
b110 6
19
1>
1C
b110 G
#732220000000
0!
0*
09
0>
0C
#732230000000
1!
1*
b111 6
19
1>
1C
b111 G
#732240000000
0!
0*
09
0>
0C
#732250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#732260000000
0!
0*
09
0>
0C
#732270000000
1!
1*
b1 6
19
1>
1C
b1 G
#732280000000
0!
0*
09
0>
0C
#732290000000
1!
1*
b10 6
19
1>
1C
b10 G
#732300000000
0!
0*
09
0>
0C
#732310000000
1!
1*
b11 6
19
1>
1C
b11 G
#732320000000
0!
0*
09
0>
0C
#732330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#732340000000
0!
0*
09
0>
0C
#732350000000
1!
1*
b101 6
19
1>
1C
b101 G
#732360000000
0!
0*
09
0>
0C
#732370000000
1!
1*
b110 6
19
1>
1C
b110 G
#732380000000
0!
0*
09
0>
0C
#732390000000
1!
1*
b111 6
19
1>
1C
b111 G
#732400000000
0!
1"
0*
1+
09
1:
0>
0C
#732410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#732420000000
0!
0*
09
0>
0C
#732430000000
1!
1*
b1 6
19
1>
1C
b1 G
#732440000000
0!
0*
09
0>
0C
#732450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#732460000000
0!
0*
09
0>
0C
#732470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#732480000000
0!
0*
09
0>
0C
#732490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#732500000000
0!
0*
09
0>
0C
#732510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#732520000000
0!
0#
0*
0,
09
0>
0?
0C
#732530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#732540000000
0!
0*
09
0>
0C
#732550000000
1!
1*
19
1>
1C
#732560000000
0!
0*
09
0>
0C
#732570000000
1!
1*
19
1>
1C
#732580000000
0!
0*
09
0>
0C
#732590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#732600000000
0!
0*
09
0>
0C
#732610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#732620000000
0!
0*
09
0>
0C
#732630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#732640000000
0!
0*
09
0>
0C
#732650000000
1!
1*
b10 6
19
1>
1C
b10 G
#732660000000
0!
0*
09
0>
0C
#732670000000
1!
1*
b11 6
19
1>
1C
b11 G
#732680000000
0!
0*
09
0>
0C
#732690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#732700000000
0!
0*
09
0>
0C
#732710000000
1!
1*
b101 6
19
1>
1C
b101 G
#732720000000
0!
0*
09
0>
0C
#732730000000
1!
1*
b110 6
19
1>
1C
b110 G
#732740000000
0!
0*
09
0>
0C
#732750000000
1!
1*
b111 6
19
1>
1C
b111 G
#732760000000
0!
0*
09
0>
0C
#732770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#732780000000
0!
0*
09
0>
0C
#732790000000
1!
1*
b1 6
19
1>
1C
b1 G
#732800000000
0!
0*
09
0>
0C
#732810000000
1!
1*
b10 6
19
1>
1C
b10 G
#732820000000
0!
0*
09
0>
0C
#732830000000
1!
1*
b11 6
19
1>
1C
b11 G
#732840000000
0!
0*
09
0>
0C
#732850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#732860000000
0!
0*
09
0>
0C
#732870000000
1!
1*
b101 6
19
1>
1C
b101 G
#732880000000
0!
0*
09
0>
0C
#732890000000
1!
1*
b110 6
19
1>
1C
b110 G
#732900000000
0!
0*
09
0>
0C
#732910000000
1!
1*
b111 6
19
1>
1C
b111 G
#732920000000
0!
0*
09
0>
0C
#732930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#732940000000
0!
0*
09
0>
0C
#732950000000
1!
1*
b1 6
19
1>
1C
b1 G
#732960000000
0!
0*
09
0>
0C
#732970000000
1!
1*
b10 6
19
1>
1C
b10 G
#732980000000
0!
0*
09
0>
0C
#732990000000
1!
1*
b11 6
19
1>
1C
b11 G
#733000000000
0!
0*
09
0>
0C
#733010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#733020000000
0!
0*
09
0>
0C
#733030000000
1!
1*
b101 6
19
1>
1C
b101 G
#733040000000
0!
0*
09
0>
0C
#733050000000
1!
1*
b110 6
19
1>
1C
b110 G
#733060000000
0!
0*
09
0>
0C
#733070000000
1!
1*
b111 6
19
1>
1C
b111 G
#733080000000
0!
1"
0*
1+
09
1:
0>
0C
#733090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#733100000000
0!
0*
09
0>
0C
#733110000000
1!
1*
b1 6
19
1>
1C
b1 G
#733120000000
0!
0*
09
0>
0C
#733130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#733140000000
0!
0*
09
0>
0C
#733150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#733160000000
0!
0*
09
0>
0C
#733170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#733180000000
0!
0*
09
0>
0C
#733190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#733200000000
0!
0#
0*
0,
09
0>
0?
0C
#733210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#733220000000
0!
0*
09
0>
0C
#733230000000
1!
1*
19
1>
1C
#733240000000
0!
0*
09
0>
0C
#733250000000
1!
1*
19
1>
1C
#733260000000
0!
0*
09
0>
0C
#733270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#733280000000
0!
0*
09
0>
0C
#733290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#733300000000
0!
0*
09
0>
0C
#733310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#733320000000
0!
0*
09
0>
0C
#733330000000
1!
1*
b10 6
19
1>
1C
b10 G
#733340000000
0!
0*
09
0>
0C
#733350000000
1!
1*
b11 6
19
1>
1C
b11 G
#733360000000
0!
0*
09
0>
0C
#733370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#733380000000
0!
0*
09
0>
0C
#733390000000
1!
1*
b101 6
19
1>
1C
b101 G
#733400000000
0!
0*
09
0>
0C
#733410000000
1!
1*
b110 6
19
1>
1C
b110 G
#733420000000
0!
0*
09
0>
0C
#733430000000
1!
1*
b111 6
19
1>
1C
b111 G
#733440000000
0!
0*
09
0>
0C
#733450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#733460000000
0!
0*
09
0>
0C
#733470000000
1!
1*
b1 6
19
1>
1C
b1 G
#733480000000
0!
0*
09
0>
0C
#733490000000
1!
1*
b10 6
19
1>
1C
b10 G
#733500000000
0!
0*
09
0>
0C
#733510000000
1!
1*
b11 6
19
1>
1C
b11 G
#733520000000
0!
0*
09
0>
0C
#733530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#733540000000
0!
0*
09
0>
0C
#733550000000
1!
1*
b101 6
19
1>
1C
b101 G
#733560000000
0!
0*
09
0>
0C
#733570000000
1!
1*
b110 6
19
1>
1C
b110 G
#733580000000
0!
0*
09
0>
0C
#733590000000
1!
1*
b111 6
19
1>
1C
b111 G
#733600000000
0!
0*
09
0>
0C
#733610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#733620000000
0!
0*
09
0>
0C
#733630000000
1!
1*
b1 6
19
1>
1C
b1 G
#733640000000
0!
0*
09
0>
0C
#733650000000
1!
1*
b10 6
19
1>
1C
b10 G
#733660000000
0!
0*
09
0>
0C
#733670000000
1!
1*
b11 6
19
1>
1C
b11 G
#733680000000
0!
0*
09
0>
0C
#733690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#733700000000
0!
0*
09
0>
0C
#733710000000
1!
1*
b101 6
19
1>
1C
b101 G
#733720000000
0!
0*
09
0>
0C
#733730000000
1!
1*
b110 6
19
1>
1C
b110 G
#733740000000
0!
0*
09
0>
0C
#733750000000
1!
1*
b111 6
19
1>
1C
b111 G
#733760000000
0!
1"
0*
1+
09
1:
0>
0C
#733770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#733780000000
0!
0*
09
0>
0C
#733790000000
1!
1*
b1 6
19
1>
1C
b1 G
#733800000000
0!
0*
09
0>
0C
#733810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#733820000000
0!
0*
09
0>
0C
#733830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#733840000000
0!
0*
09
0>
0C
#733850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#733860000000
0!
0*
09
0>
0C
#733870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#733880000000
0!
0#
0*
0,
09
0>
0?
0C
#733890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#733900000000
0!
0*
09
0>
0C
#733910000000
1!
1*
19
1>
1C
#733920000000
0!
0*
09
0>
0C
#733930000000
1!
1*
19
1>
1C
#733940000000
0!
0*
09
0>
0C
#733950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#733960000000
0!
0*
09
0>
0C
#733970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#733980000000
0!
0*
09
0>
0C
#733990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#734000000000
0!
0*
09
0>
0C
#734010000000
1!
1*
b10 6
19
1>
1C
b10 G
#734020000000
0!
0*
09
0>
0C
#734030000000
1!
1*
b11 6
19
1>
1C
b11 G
#734040000000
0!
0*
09
0>
0C
#734050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#734060000000
0!
0*
09
0>
0C
#734070000000
1!
1*
b101 6
19
1>
1C
b101 G
#734080000000
0!
0*
09
0>
0C
#734090000000
1!
1*
b110 6
19
1>
1C
b110 G
#734100000000
0!
0*
09
0>
0C
#734110000000
1!
1*
b111 6
19
1>
1C
b111 G
#734120000000
0!
0*
09
0>
0C
#734130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#734140000000
0!
0*
09
0>
0C
#734150000000
1!
1*
b1 6
19
1>
1C
b1 G
#734160000000
0!
0*
09
0>
0C
#734170000000
1!
1*
b10 6
19
1>
1C
b10 G
#734180000000
0!
0*
09
0>
0C
#734190000000
1!
1*
b11 6
19
1>
1C
b11 G
#734200000000
0!
0*
09
0>
0C
#734210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#734220000000
0!
0*
09
0>
0C
#734230000000
1!
1*
b101 6
19
1>
1C
b101 G
#734240000000
0!
0*
09
0>
0C
#734250000000
1!
1*
b110 6
19
1>
1C
b110 G
#734260000000
0!
0*
09
0>
0C
#734270000000
1!
1*
b111 6
19
1>
1C
b111 G
#734280000000
0!
0*
09
0>
0C
#734290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#734300000000
0!
0*
09
0>
0C
#734310000000
1!
1*
b1 6
19
1>
1C
b1 G
#734320000000
0!
0*
09
0>
0C
#734330000000
1!
1*
b10 6
19
1>
1C
b10 G
#734340000000
0!
0*
09
0>
0C
#734350000000
1!
1*
b11 6
19
1>
1C
b11 G
#734360000000
0!
0*
09
0>
0C
#734370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#734380000000
0!
0*
09
0>
0C
#734390000000
1!
1*
b101 6
19
1>
1C
b101 G
#734400000000
0!
0*
09
0>
0C
#734410000000
1!
1*
b110 6
19
1>
1C
b110 G
#734420000000
0!
0*
09
0>
0C
#734430000000
1!
1*
b111 6
19
1>
1C
b111 G
#734440000000
0!
1"
0*
1+
09
1:
0>
0C
#734450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#734460000000
0!
0*
09
0>
0C
#734470000000
1!
1*
b1 6
19
1>
1C
b1 G
#734480000000
0!
0*
09
0>
0C
#734490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#734500000000
0!
0*
09
0>
0C
#734510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#734520000000
0!
0*
09
0>
0C
#734530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#734540000000
0!
0*
09
0>
0C
#734550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#734560000000
0!
0#
0*
0,
09
0>
0?
0C
#734570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#734580000000
0!
0*
09
0>
0C
#734590000000
1!
1*
19
1>
1C
#734600000000
0!
0*
09
0>
0C
#734610000000
1!
1*
19
1>
1C
#734620000000
0!
0*
09
0>
0C
#734630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#734640000000
0!
0*
09
0>
0C
#734650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#734660000000
0!
0*
09
0>
0C
#734670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#734680000000
0!
0*
09
0>
0C
#734690000000
1!
1*
b10 6
19
1>
1C
b10 G
#734700000000
0!
0*
09
0>
0C
#734710000000
1!
1*
b11 6
19
1>
1C
b11 G
#734720000000
0!
0*
09
0>
0C
#734730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#734740000000
0!
0*
09
0>
0C
#734750000000
1!
1*
b101 6
19
1>
1C
b101 G
#734760000000
0!
0*
09
0>
0C
#734770000000
1!
1*
b110 6
19
1>
1C
b110 G
#734780000000
0!
0*
09
0>
0C
#734790000000
1!
1*
b111 6
19
1>
1C
b111 G
#734800000000
0!
0*
09
0>
0C
#734810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#734820000000
0!
0*
09
0>
0C
#734830000000
1!
1*
b1 6
19
1>
1C
b1 G
#734840000000
0!
0*
09
0>
0C
#734850000000
1!
1*
b10 6
19
1>
1C
b10 G
#734860000000
0!
0*
09
0>
0C
#734870000000
1!
1*
b11 6
19
1>
1C
b11 G
#734880000000
0!
0*
09
0>
0C
#734890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#734900000000
0!
0*
09
0>
0C
#734910000000
1!
1*
b101 6
19
1>
1C
b101 G
#734920000000
0!
0*
09
0>
0C
#734930000000
1!
1*
b110 6
19
1>
1C
b110 G
#734940000000
0!
0*
09
0>
0C
#734950000000
1!
1*
b111 6
19
1>
1C
b111 G
#734960000000
0!
0*
09
0>
0C
#734970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#734980000000
0!
0*
09
0>
0C
#734990000000
1!
1*
b1 6
19
1>
1C
b1 G
#735000000000
0!
0*
09
0>
0C
#735010000000
1!
1*
b10 6
19
1>
1C
b10 G
#735020000000
0!
0*
09
0>
0C
#735030000000
1!
1*
b11 6
19
1>
1C
b11 G
#735040000000
0!
0*
09
0>
0C
#735050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#735060000000
0!
0*
09
0>
0C
#735070000000
1!
1*
b101 6
19
1>
1C
b101 G
#735080000000
0!
0*
09
0>
0C
#735090000000
1!
1*
b110 6
19
1>
1C
b110 G
#735100000000
0!
0*
09
0>
0C
#735110000000
1!
1*
b111 6
19
1>
1C
b111 G
#735120000000
0!
1"
0*
1+
09
1:
0>
0C
#735130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#735140000000
0!
0*
09
0>
0C
#735150000000
1!
1*
b1 6
19
1>
1C
b1 G
#735160000000
0!
0*
09
0>
0C
#735170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#735180000000
0!
0*
09
0>
0C
#735190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#735200000000
0!
0*
09
0>
0C
#735210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#735220000000
0!
0*
09
0>
0C
#735230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#735240000000
0!
0#
0*
0,
09
0>
0?
0C
#735250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#735260000000
0!
0*
09
0>
0C
#735270000000
1!
1*
19
1>
1C
#735280000000
0!
0*
09
0>
0C
#735290000000
1!
1*
19
1>
1C
#735300000000
0!
0*
09
0>
0C
#735310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#735320000000
0!
0*
09
0>
0C
#735330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#735340000000
0!
0*
09
0>
0C
#735350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#735360000000
0!
0*
09
0>
0C
#735370000000
1!
1*
b10 6
19
1>
1C
b10 G
#735380000000
0!
0*
09
0>
0C
#735390000000
1!
1*
b11 6
19
1>
1C
b11 G
#735400000000
0!
0*
09
0>
0C
#735410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#735420000000
0!
0*
09
0>
0C
#735430000000
1!
1*
b101 6
19
1>
1C
b101 G
#735440000000
0!
0*
09
0>
0C
#735450000000
1!
1*
b110 6
19
1>
1C
b110 G
#735460000000
0!
0*
09
0>
0C
#735470000000
1!
1*
b111 6
19
1>
1C
b111 G
#735480000000
0!
0*
09
0>
0C
#735490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#735500000000
0!
0*
09
0>
0C
#735510000000
1!
1*
b1 6
19
1>
1C
b1 G
#735520000000
0!
0*
09
0>
0C
#735530000000
1!
1*
b10 6
19
1>
1C
b10 G
#735540000000
0!
0*
09
0>
0C
#735550000000
1!
1*
b11 6
19
1>
1C
b11 G
#735560000000
0!
0*
09
0>
0C
#735570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#735580000000
0!
0*
09
0>
0C
#735590000000
1!
1*
b101 6
19
1>
1C
b101 G
#735600000000
0!
0*
09
0>
0C
#735610000000
1!
1*
b110 6
19
1>
1C
b110 G
#735620000000
0!
0*
09
0>
0C
#735630000000
1!
1*
b111 6
19
1>
1C
b111 G
#735640000000
0!
0*
09
0>
0C
#735650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#735660000000
0!
0*
09
0>
0C
#735670000000
1!
1*
b1 6
19
1>
1C
b1 G
#735680000000
0!
0*
09
0>
0C
#735690000000
1!
1*
b10 6
19
1>
1C
b10 G
#735700000000
0!
0*
09
0>
0C
#735710000000
1!
1*
b11 6
19
1>
1C
b11 G
#735720000000
0!
0*
09
0>
0C
#735730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#735740000000
0!
0*
09
0>
0C
#735750000000
1!
1*
b101 6
19
1>
1C
b101 G
#735760000000
0!
0*
09
0>
0C
#735770000000
1!
1*
b110 6
19
1>
1C
b110 G
#735780000000
0!
0*
09
0>
0C
#735790000000
1!
1*
b111 6
19
1>
1C
b111 G
#735800000000
0!
1"
0*
1+
09
1:
0>
0C
#735810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#735820000000
0!
0*
09
0>
0C
#735830000000
1!
1*
b1 6
19
1>
1C
b1 G
#735840000000
0!
0*
09
0>
0C
#735850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#735860000000
0!
0*
09
0>
0C
#735870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#735880000000
0!
0*
09
0>
0C
#735890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#735900000000
0!
0*
09
0>
0C
#735910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#735920000000
0!
0#
0*
0,
09
0>
0?
0C
#735930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#735940000000
0!
0*
09
0>
0C
#735950000000
1!
1*
19
1>
1C
#735960000000
0!
0*
09
0>
0C
#735970000000
1!
1*
19
1>
1C
#735980000000
0!
0*
09
0>
0C
#735990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#736000000000
0!
0*
09
0>
0C
#736010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#736020000000
0!
0*
09
0>
0C
#736030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#736040000000
0!
0*
09
0>
0C
#736050000000
1!
1*
b10 6
19
1>
1C
b10 G
#736060000000
0!
0*
09
0>
0C
#736070000000
1!
1*
b11 6
19
1>
1C
b11 G
#736080000000
0!
0*
09
0>
0C
#736090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#736100000000
0!
0*
09
0>
0C
#736110000000
1!
1*
b101 6
19
1>
1C
b101 G
#736120000000
0!
0*
09
0>
0C
#736130000000
1!
1*
b110 6
19
1>
1C
b110 G
#736140000000
0!
0*
09
0>
0C
#736150000000
1!
1*
b111 6
19
1>
1C
b111 G
#736160000000
0!
0*
09
0>
0C
#736170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#736180000000
0!
0*
09
0>
0C
#736190000000
1!
1*
b1 6
19
1>
1C
b1 G
#736200000000
0!
0*
09
0>
0C
#736210000000
1!
1*
b10 6
19
1>
1C
b10 G
#736220000000
0!
0*
09
0>
0C
#736230000000
1!
1*
b11 6
19
1>
1C
b11 G
#736240000000
0!
0*
09
0>
0C
#736250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#736260000000
0!
0*
09
0>
0C
#736270000000
1!
1*
b101 6
19
1>
1C
b101 G
#736280000000
0!
0*
09
0>
0C
#736290000000
1!
1*
b110 6
19
1>
1C
b110 G
#736300000000
0!
0*
09
0>
0C
#736310000000
1!
1*
b111 6
19
1>
1C
b111 G
#736320000000
0!
0*
09
0>
0C
#736330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#736340000000
0!
0*
09
0>
0C
#736350000000
1!
1*
b1 6
19
1>
1C
b1 G
#736360000000
0!
0*
09
0>
0C
#736370000000
1!
1*
b10 6
19
1>
1C
b10 G
#736380000000
0!
0*
09
0>
0C
#736390000000
1!
1*
b11 6
19
1>
1C
b11 G
#736400000000
0!
0*
09
0>
0C
#736410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#736420000000
0!
0*
09
0>
0C
#736430000000
1!
1*
b101 6
19
1>
1C
b101 G
#736440000000
0!
0*
09
0>
0C
#736450000000
1!
1*
b110 6
19
1>
1C
b110 G
#736460000000
0!
0*
09
0>
0C
#736470000000
1!
1*
b111 6
19
1>
1C
b111 G
#736480000000
0!
1"
0*
1+
09
1:
0>
0C
#736490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#736500000000
0!
0*
09
0>
0C
#736510000000
1!
1*
b1 6
19
1>
1C
b1 G
#736520000000
0!
0*
09
0>
0C
#736530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#736540000000
0!
0*
09
0>
0C
#736550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#736560000000
0!
0*
09
0>
0C
#736570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#736580000000
0!
0*
09
0>
0C
#736590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#736600000000
0!
0#
0*
0,
09
0>
0?
0C
#736610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#736620000000
0!
0*
09
0>
0C
#736630000000
1!
1*
19
1>
1C
#736640000000
0!
0*
09
0>
0C
#736650000000
1!
1*
19
1>
1C
#736660000000
0!
0*
09
0>
0C
#736670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#736680000000
0!
0*
09
0>
0C
#736690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#736700000000
0!
0*
09
0>
0C
#736710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#736720000000
0!
0*
09
0>
0C
#736730000000
1!
1*
b10 6
19
1>
1C
b10 G
#736740000000
0!
0*
09
0>
0C
#736750000000
1!
1*
b11 6
19
1>
1C
b11 G
#736760000000
0!
0*
09
0>
0C
#736770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#736780000000
0!
0*
09
0>
0C
#736790000000
1!
1*
b101 6
19
1>
1C
b101 G
#736800000000
0!
0*
09
0>
0C
#736810000000
1!
1*
b110 6
19
1>
1C
b110 G
#736820000000
0!
0*
09
0>
0C
#736830000000
1!
1*
b111 6
19
1>
1C
b111 G
#736840000000
0!
0*
09
0>
0C
#736850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#736860000000
0!
0*
09
0>
0C
#736870000000
1!
1*
b1 6
19
1>
1C
b1 G
#736880000000
0!
0*
09
0>
0C
#736890000000
1!
1*
b10 6
19
1>
1C
b10 G
#736900000000
0!
0*
09
0>
0C
#736910000000
1!
1*
b11 6
19
1>
1C
b11 G
#736920000000
0!
0*
09
0>
0C
#736930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#736940000000
0!
0*
09
0>
0C
#736950000000
1!
1*
b101 6
19
1>
1C
b101 G
#736960000000
0!
0*
09
0>
0C
#736970000000
1!
1*
b110 6
19
1>
1C
b110 G
#736980000000
0!
0*
09
0>
0C
#736990000000
1!
1*
b111 6
19
1>
1C
b111 G
#737000000000
0!
0*
09
0>
0C
#737010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#737020000000
0!
0*
09
0>
0C
#737030000000
1!
1*
b1 6
19
1>
1C
b1 G
#737040000000
0!
0*
09
0>
0C
#737050000000
1!
1*
b10 6
19
1>
1C
b10 G
#737060000000
0!
0*
09
0>
0C
#737070000000
1!
1*
b11 6
19
1>
1C
b11 G
#737080000000
0!
0*
09
0>
0C
#737090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#737100000000
0!
0*
09
0>
0C
#737110000000
1!
1*
b101 6
19
1>
1C
b101 G
#737120000000
0!
0*
09
0>
0C
#737130000000
1!
1*
b110 6
19
1>
1C
b110 G
#737140000000
0!
0*
09
0>
0C
#737150000000
1!
1*
b111 6
19
1>
1C
b111 G
#737160000000
0!
1"
0*
1+
09
1:
0>
0C
#737170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#737180000000
0!
0*
09
0>
0C
#737190000000
1!
1*
b1 6
19
1>
1C
b1 G
#737200000000
0!
0*
09
0>
0C
#737210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#737220000000
0!
0*
09
0>
0C
#737230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#737240000000
0!
0*
09
0>
0C
#737250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#737260000000
0!
0*
09
0>
0C
#737270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#737280000000
0!
0#
0*
0,
09
0>
0?
0C
#737290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#737300000000
0!
0*
09
0>
0C
#737310000000
1!
1*
19
1>
1C
#737320000000
0!
0*
09
0>
0C
#737330000000
1!
1*
19
1>
1C
#737340000000
0!
0*
09
0>
0C
#737350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#737360000000
0!
0*
09
0>
0C
#737370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#737380000000
0!
0*
09
0>
0C
#737390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#737400000000
0!
0*
09
0>
0C
#737410000000
1!
1*
b10 6
19
1>
1C
b10 G
#737420000000
0!
0*
09
0>
0C
#737430000000
1!
1*
b11 6
19
1>
1C
b11 G
#737440000000
0!
0*
09
0>
0C
#737450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#737460000000
0!
0*
09
0>
0C
#737470000000
1!
1*
b101 6
19
1>
1C
b101 G
#737480000000
0!
0*
09
0>
0C
#737490000000
1!
1*
b110 6
19
1>
1C
b110 G
#737500000000
0!
0*
09
0>
0C
#737510000000
1!
1*
b111 6
19
1>
1C
b111 G
#737520000000
0!
0*
09
0>
0C
#737530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#737540000000
0!
0*
09
0>
0C
#737550000000
1!
1*
b1 6
19
1>
1C
b1 G
#737560000000
0!
0*
09
0>
0C
#737570000000
1!
1*
b10 6
19
1>
1C
b10 G
#737580000000
0!
0*
09
0>
0C
#737590000000
1!
1*
b11 6
19
1>
1C
b11 G
#737600000000
0!
0*
09
0>
0C
#737610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#737620000000
0!
0*
09
0>
0C
#737630000000
1!
1*
b101 6
19
1>
1C
b101 G
#737640000000
0!
0*
09
0>
0C
#737650000000
1!
1*
b110 6
19
1>
1C
b110 G
#737660000000
0!
0*
09
0>
0C
#737670000000
1!
1*
b111 6
19
1>
1C
b111 G
#737680000000
0!
0*
09
0>
0C
#737690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#737700000000
0!
0*
09
0>
0C
#737710000000
1!
1*
b1 6
19
1>
1C
b1 G
#737720000000
0!
0*
09
0>
0C
#737730000000
1!
1*
b10 6
19
1>
1C
b10 G
#737740000000
0!
0*
09
0>
0C
#737750000000
1!
1*
b11 6
19
1>
1C
b11 G
#737760000000
0!
0*
09
0>
0C
#737770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#737780000000
0!
0*
09
0>
0C
#737790000000
1!
1*
b101 6
19
1>
1C
b101 G
#737800000000
0!
0*
09
0>
0C
#737810000000
1!
1*
b110 6
19
1>
1C
b110 G
#737820000000
0!
0*
09
0>
0C
#737830000000
1!
1*
b111 6
19
1>
1C
b111 G
#737840000000
0!
1"
0*
1+
09
1:
0>
0C
#737850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#737860000000
0!
0*
09
0>
0C
#737870000000
1!
1*
b1 6
19
1>
1C
b1 G
#737880000000
0!
0*
09
0>
0C
#737890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#737900000000
0!
0*
09
0>
0C
#737910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#737920000000
0!
0*
09
0>
0C
#737930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#737940000000
0!
0*
09
0>
0C
#737950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#737960000000
0!
0#
0*
0,
09
0>
0?
0C
#737970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#737980000000
0!
0*
09
0>
0C
#737990000000
1!
1*
19
1>
1C
#738000000000
0!
0*
09
0>
0C
#738010000000
1!
1*
19
1>
1C
#738020000000
0!
0*
09
0>
0C
#738030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#738040000000
0!
0*
09
0>
0C
#738050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#738060000000
0!
0*
09
0>
0C
#738070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#738080000000
0!
0*
09
0>
0C
#738090000000
1!
1*
b10 6
19
1>
1C
b10 G
#738100000000
0!
0*
09
0>
0C
#738110000000
1!
1*
b11 6
19
1>
1C
b11 G
#738120000000
0!
0*
09
0>
0C
#738130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#738140000000
0!
0*
09
0>
0C
#738150000000
1!
1*
b101 6
19
1>
1C
b101 G
#738160000000
0!
0*
09
0>
0C
#738170000000
1!
1*
b110 6
19
1>
1C
b110 G
#738180000000
0!
0*
09
0>
0C
#738190000000
1!
1*
b111 6
19
1>
1C
b111 G
#738200000000
0!
0*
09
0>
0C
#738210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#738220000000
0!
0*
09
0>
0C
#738230000000
1!
1*
b1 6
19
1>
1C
b1 G
#738240000000
0!
0*
09
0>
0C
#738250000000
1!
1*
b10 6
19
1>
1C
b10 G
#738260000000
0!
0*
09
0>
0C
#738270000000
1!
1*
b11 6
19
1>
1C
b11 G
#738280000000
0!
0*
09
0>
0C
#738290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#738300000000
0!
0*
09
0>
0C
#738310000000
1!
1*
b101 6
19
1>
1C
b101 G
#738320000000
0!
0*
09
0>
0C
#738330000000
1!
1*
b110 6
19
1>
1C
b110 G
#738340000000
0!
0*
09
0>
0C
#738350000000
1!
1*
b111 6
19
1>
1C
b111 G
#738360000000
0!
0*
09
0>
0C
#738370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#738380000000
0!
0*
09
0>
0C
#738390000000
1!
1*
b1 6
19
1>
1C
b1 G
#738400000000
0!
0*
09
0>
0C
#738410000000
1!
1*
b10 6
19
1>
1C
b10 G
#738420000000
0!
0*
09
0>
0C
#738430000000
1!
1*
b11 6
19
1>
1C
b11 G
#738440000000
0!
0*
09
0>
0C
#738450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#738460000000
0!
0*
09
0>
0C
#738470000000
1!
1*
b101 6
19
1>
1C
b101 G
#738480000000
0!
0*
09
0>
0C
#738490000000
1!
1*
b110 6
19
1>
1C
b110 G
#738500000000
0!
0*
09
0>
0C
#738510000000
1!
1*
b111 6
19
1>
1C
b111 G
#738520000000
0!
1"
0*
1+
09
1:
0>
0C
#738530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#738540000000
0!
0*
09
0>
0C
#738550000000
1!
1*
b1 6
19
1>
1C
b1 G
#738560000000
0!
0*
09
0>
0C
#738570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#738580000000
0!
0*
09
0>
0C
#738590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#738600000000
0!
0*
09
0>
0C
#738610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#738620000000
0!
0*
09
0>
0C
#738630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#738640000000
0!
0#
0*
0,
09
0>
0?
0C
#738650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#738660000000
0!
0*
09
0>
0C
#738670000000
1!
1*
19
1>
1C
#738680000000
0!
0*
09
0>
0C
#738690000000
1!
1*
19
1>
1C
#738700000000
0!
0*
09
0>
0C
#738710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#738720000000
0!
0*
09
0>
0C
#738730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#738740000000
0!
0*
09
0>
0C
#738750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#738760000000
0!
0*
09
0>
0C
#738770000000
1!
1*
b10 6
19
1>
1C
b10 G
#738780000000
0!
0*
09
0>
0C
#738790000000
1!
1*
b11 6
19
1>
1C
b11 G
#738800000000
0!
0*
09
0>
0C
#738810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#738820000000
0!
0*
09
0>
0C
#738830000000
1!
1*
b101 6
19
1>
1C
b101 G
#738840000000
0!
0*
09
0>
0C
#738850000000
1!
1*
b110 6
19
1>
1C
b110 G
#738860000000
0!
0*
09
0>
0C
#738870000000
1!
1*
b111 6
19
1>
1C
b111 G
#738880000000
0!
0*
09
0>
0C
#738890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#738900000000
0!
0*
09
0>
0C
#738910000000
1!
1*
b1 6
19
1>
1C
b1 G
#738920000000
0!
0*
09
0>
0C
#738930000000
1!
1*
b10 6
19
1>
1C
b10 G
#738940000000
0!
0*
09
0>
0C
#738950000000
1!
1*
b11 6
19
1>
1C
b11 G
#738960000000
0!
0*
09
0>
0C
#738970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#738980000000
0!
0*
09
0>
0C
#738990000000
1!
1*
b101 6
19
1>
1C
b101 G
#739000000000
0!
0*
09
0>
0C
#739010000000
1!
1*
b110 6
19
1>
1C
b110 G
#739020000000
0!
0*
09
0>
0C
#739030000000
1!
1*
b111 6
19
1>
1C
b111 G
#739040000000
0!
0*
09
0>
0C
#739050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#739060000000
0!
0*
09
0>
0C
#739070000000
1!
1*
b1 6
19
1>
1C
b1 G
#739080000000
0!
0*
09
0>
0C
#739090000000
1!
1*
b10 6
19
1>
1C
b10 G
#739100000000
0!
0*
09
0>
0C
#739110000000
1!
1*
b11 6
19
1>
1C
b11 G
#739120000000
0!
0*
09
0>
0C
#739130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#739140000000
0!
0*
09
0>
0C
#739150000000
1!
1*
b101 6
19
1>
1C
b101 G
#739160000000
0!
0*
09
0>
0C
#739170000000
1!
1*
b110 6
19
1>
1C
b110 G
#739180000000
0!
0*
09
0>
0C
#739190000000
1!
1*
b111 6
19
1>
1C
b111 G
#739200000000
0!
1"
0*
1+
09
1:
0>
0C
#739210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#739220000000
0!
0*
09
0>
0C
#739230000000
1!
1*
b1 6
19
1>
1C
b1 G
#739240000000
0!
0*
09
0>
0C
#739250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#739260000000
0!
0*
09
0>
0C
#739270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#739280000000
0!
0*
09
0>
0C
#739290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#739300000000
0!
0*
09
0>
0C
#739310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#739320000000
0!
0#
0*
0,
09
0>
0?
0C
#739330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#739340000000
0!
0*
09
0>
0C
#739350000000
1!
1*
19
1>
1C
#739360000000
0!
0*
09
0>
0C
#739370000000
1!
1*
19
1>
1C
#739380000000
0!
0*
09
0>
0C
#739390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#739400000000
0!
0*
09
0>
0C
#739410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#739420000000
0!
0*
09
0>
0C
#739430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#739440000000
0!
0*
09
0>
0C
#739450000000
1!
1*
b10 6
19
1>
1C
b10 G
#739460000000
0!
0*
09
0>
0C
#739470000000
1!
1*
b11 6
19
1>
1C
b11 G
#739480000000
0!
0*
09
0>
0C
#739490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#739500000000
0!
0*
09
0>
0C
#739510000000
1!
1*
b101 6
19
1>
1C
b101 G
#739520000000
0!
0*
09
0>
0C
#739530000000
1!
1*
b110 6
19
1>
1C
b110 G
#739540000000
0!
0*
09
0>
0C
#739550000000
1!
1*
b111 6
19
1>
1C
b111 G
#739560000000
0!
0*
09
0>
0C
#739570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#739580000000
0!
0*
09
0>
0C
#739590000000
1!
1*
b1 6
19
1>
1C
b1 G
#739600000000
0!
0*
09
0>
0C
#739610000000
1!
1*
b10 6
19
1>
1C
b10 G
#739620000000
0!
0*
09
0>
0C
#739630000000
1!
1*
b11 6
19
1>
1C
b11 G
#739640000000
0!
0*
09
0>
0C
#739650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#739660000000
0!
0*
09
0>
0C
#739670000000
1!
1*
b101 6
19
1>
1C
b101 G
#739680000000
0!
0*
09
0>
0C
#739690000000
1!
1*
b110 6
19
1>
1C
b110 G
#739700000000
0!
0*
09
0>
0C
#739710000000
1!
1*
b111 6
19
1>
1C
b111 G
#739720000000
0!
0*
09
0>
0C
#739730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#739740000000
0!
0*
09
0>
0C
#739750000000
1!
1*
b1 6
19
1>
1C
b1 G
#739760000000
0!
0*
09
0>
0C
#739770000000
1!
1*
b10 6
19
1>
1C
b10 G
#739780000000
0!
0*
09
0>
0C
#739790000000
1!
1*
b11 6
19
1>
1C
b11 G
#739800000000
0!
0*
09
0>
0C
#739810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#739820000000
0!
0*
09
0>
0C
#739830000000
1!
1*
b101 6
19
1>
1C
b101 G
#739840000000
0!
0*
09
0>
0C
#739850000000
1!
1*
b110 6
19
1>
1C
b110 G
#739860000000
0!
0*
09
0>
0C
#739870000000
1!
1*
b111 6
19
1>
1C
b111 G
#739880000000
0!
1"
0*
1+
09
1:
0>
0C
#739890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#739900000000
0!
0*
09
0>
0C
#739910000000
1!
1*
b1 6
19
1>
1C
b1 G
#739920000000
0!
0*
09
0>
0C
#739930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#739940000000
0!
0*
09
0>
0C
#739950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#739960000000
0!
0*
09
0>
0C
#739970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#739980000000
0!
0*
09
0>
0C
#739990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#740000000000
0!
0#
0*
0,
09
0>
0?
0C
#740010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#740020000000
0!
0*
09
0>
0C
#740030000000
1!
1*
19
1>
1C
#740040000000
0!
0*
09
0>
0C
#740050000000
1!
1*
19
1>
1C
#740060000000
0!
0*
09
0>
0C
#740070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#740080000000
0!
0*
09
0>
0C
#740090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#740100000000
0!
0*
09
0>
0C
#740110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#740120000000
0!
0*
09
0>
0C
#740130000000
1!
1*
b10 6
19
1>
1C
b10 G
#740140000000
0!
0*
09
0>
0C
#740150000000
1!
1*
b11 6
19
1>
1C
b11 G
#740160000000
0!
0*
09
0>
0C
#740170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#740180000000
0!
0*
09
0>
0C
#740190000000
1!
1*
b101 6
19
1>
1C
b101 G
#740200000000
0!
0*
09
0>
0C
#740210000000
1!
1*
b110 6
19
1>
1C
b110 G
#740220000000
0!
0*
09
0>
0C
#740230000000
1!
1*
b111 6
19
1>
1C
b111 G
#740240000000
0!
0*
09
0>
0C
#740250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#740260000000
0!
0*
09
0>
0C
#740270000000
1!
1*
b1 6
19
1>
1C
b1 G
#740280000000
0!
0*
09
0>
0C
#740290000000
1!
1*
b10 6
19
1>
1C
b10 G
#740300000000
0!
0*
09
0>
0C
#740310000000
1!
1*
b11 6
19
1>
1C
b11 G
#740320000000
0!
0*
09
0>
0C
#740330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#740340000000
0!
0*
09
0>
0C
#740350000000
1!
1*
b101 6
19
1>
1C
b101 G
#740360000000
0!
0*
09
0>
0C
#740370000000
1!
1*
b110 6
19
1>
1C
b110 G
#740380000000
0!
0*
09
0>
0C
#740390000000
1!
1*
b111 6
19
1>
1C
b111 G
#740400000000
0!
0*
09
0>
0C
#740410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#740420000000
0!
0*
09
0>
0C
#740430000000
1!
1*
b1 6
19
1>
1C
b1 G
#740440000000
0!
0*
09
0>
0C
#740450000000
1!
1*
b10 6
19
1>
1C
b10 G
#740460000000
0!
0*
09
0>
0C
#740470000000
1!
1*
b11 6
19
1>
1C
b11 G
#740480000000
0!
0*
09
0>
0C
#740490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#740500000000
0!
0*
09
0>
0C
#740510000000
1!
1*
b101 6
19
1>
1C
b101 G
#740520000000
0!
0*
09
0>
0C
#740530000000
1!
1*
b110 6
19
1>
1C
b110 G
#740540000000
0!
0*
09
0>
0C
#740550000000
1!
1*
b111 6
19
1>
1C
b111 G
#740560000000
0!
1"
0*
1+
09
1:
0>
0C
#740570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#740580000000
0!
0*
09
0>
0C
#740590000000
1!
1*
b1 6
19
1>
1C
b1 G
#740600000000
0!
0*
09
0>
0C
#740610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#740620000000
0!
0*
09
0>
0C
#740630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#740640000000
0!
0*
09
0>
0C
#740650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#740660000000
0!
0*
09
0>
0C
#740670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#740680000000
0!
0#
0*
0,
09
0>
0?
0C
#740690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#740700000000
0!
0*
09
0>
0C
#740710000000
1!
1*
19
1>
1C
#740720000000
0!
0*
09
0>
0C
#740730000000
1!
1*
19
1>
1C
#740740000000
0!
0*
09
0>
0C
#740750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#740760000000
0!
0*
09
0>
0C
#740770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#740780000000
0!
0*
09
0>
0C
#740790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#740800000000
0!
0*
09
0>
0C
#740810000000
1!
1*
b10 6
19
1>
1C
b10 G
#740820000000
0!
0*
09
0>
0C
#740830000000
1!
1*
b11 6
19
1>
1C
b11 G
#740840000000
0!
0*
09
0>
0C
#740850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#740860000000
0!
0*
09
0>
0C
#740870000000
1!
1*
b101 6
19
1>
1C
b101 G
#740880000000
0!
0*
09
0>
0C
#740890000000
1!
1*
b110 6
19
1>
1C
b110 G
#740900000000
0!
0*
09
0>
0C
#740910000000
1!
1*
b111 6
19
1>
1C
b111 G
#740920000000
0!
0*
09
0>
0C
#740930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#740940000000
0!
0*
09
0>
0C
#740950000000
1!
1*
b1 6
19
1>
1C
b1 G
#740960000000
0!
0*
09
0>
0C
#740970000000
1!
1*
b10 6
19
1>
1C
b10 G
#740980000000
0!
0*
09
0>
0C
#740990000000
1!
1*
b11 6
19
1>
1C
b11 G
#741000000000
0!
0*
09
0>
0C
#741010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#741020000000
0!
0*
09
0>
0C
#741030000000
1!
1*
b101 6
19
1>
1C
b101 G
#741040000000
0!
0*
09
0>
0C
#741050000000
1!
1*
b110 6
19
1>
1C
b110 G
#741060000000
0!
0*
09
0>
0C
#741070000000
1!
1*
b111 6
19
1>
1C
b111 G
#741080000000
0!
0*
09
0>
0C
#741090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#741100000000
0!
0*
09
0>
0C
#741110000000
1!
1*
b1 6
19
1>
1C
b1 G
#741120000000
0!
0*
09
0>
0C
#741130000000
1!
1*
b10 6
19
1>
1C
b10 G
#741140000000
0!
0*
09
0>
0C
#741150000000
1!
1*
b11 6
19
1>
1C
b11 G
#741160000000
0!
0*
09
0>
0C
#741170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#741180000000
0!
0*
09
0>
0C
#741190000000
1!
1*
b101 6
19
1>
1C
b101 G
#741200000000
0!
0*
09
0>
0C
#741210000000
1!
1*
b110 6
19
1>
1C
b110 G
#741220000000
0!
0*
09
0>
0C
#741230000000
1!
1*
b111 6
19
1>
1C
b111 G
#741240000000
0!
1"
0*
1+
09
1:
0>
0C
#741250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#741260000000
0!
0*
09
0>
0C
#741270000000
1!
1*
b1 6
19
1>
1C
b1 G
#741280000000
0!
0*
09
0>
0C
#741290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#741300000000
0!
0*
09
0>
0C
#741310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#741320000000
0!
0*
09
0>
0C
#741330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#741340000000
0!
0*
09
0>
0C
#741350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#741360000000
0!
0#
0*
0,
09
0>
0?
0C
#741370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#741380000000
0!
0*
09
0>
0C
#741390000000
1!
1*
19
1>
1C
#741400000000
0!
0*
09
0>
0C
#741410000000
1!
1*
19
1>
1C
#741420000000
0!
0*
09
0>
0C
#741430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#741440000000
0!
0*
09
0>
0C
#741450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#741460000000
0!
0*
09
0>
0C
#741470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#741480000000
0!
0*
09
0>
0C
#741490000000
1!
1*
b10 6
19
1>
1C
b10 G
#741500000000
0!
0*
09
0>
0C
#741510000000
1!
1*
b11 6
19
1>
1C
b11 G
#741520000000
0!
0*
09
0>
0C
#741530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#741540000000
0!
0*
09
0>
0C
#741550000000
1!
1*
b101 6
19
1>
1C
b101 G
#741560000000
0!
0*
09
0>
0C
#741570000000
1!
1*
b110 6
19
1>
1C
b110 G
#741580000000
0!
0*
09
0>
0C
#741590000000
1!
1*
b111 6
19
1>
1C
b111 G
#741600000000
0!
0*
09
0>
0C
#741610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#741620000000
0!
0*
09
0>
0C
#741630000000
1!
1*
b1 6
19
1>
1C
b1 G
#741640000000
0!
0*
09
0>
0C
#741650000000
1!
1*
b10 6
19
1>
1C
b10 G
#741660000000
0!
0*
09
0>
0C
#741670000000
1!
1*
b11 6
19
1>
1C
b11 G
#741680000000
0!
0*
09
0>
0C
#741690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#741700000000
0!
0*
09
0>
0C
#741710000000
1!
1*
b101 6
19
1>
1C
b101 G
#741720000000
0!
0*
09
0>
0C
#741730000000
1!
1*
b110 6
19
1>
1C
b110 G
#741740000000
0!
0*
09
0>
0C
#741750000000
1!
1*
b111 6
19
1>
1C
b111 G
#741760000000
0!
0*
09
0>
0C
#741770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#741780000000
0!
0*
09
0>
0C
#741790000000
1!
1*
b1 6
19
1>
1C
b1 G
#741800000000
0!
0*
09
0>
0C
#741810000000
1!
1*
b10 6
19
1>
1C
b10 G
#741820000000
0!
0*
09
0>
0C
#741830000000
1!
1*
b11 6
19
1>
1C
b11 G
#741840000000
0!
0*
09
0>
0C
#741850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#741860000000
0!
0*
09
0>
0C
#741870000000
1!
1*
b101 6
19
1>
1C
b101 G
#741880000000
0!
0*
09
0>
0C
#741890000000
1!
1*
b110 6
19
1>
1C
b110 G
#741900000000
0!
0*
09
0>
0C
#741910000000
1!
1*
b111 6
19
1>
1C
b111 G
#741920000000
0!
1"
0*
1+
09
1:
0>
0C
#741930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#741940000000
0!
0*
09
0>
0C
#741950000000
1!
1*
b1 6
19
1>
1C
b1 G
#741960000000
0!
0*
09
0>
0C
#741970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#741980000000
0!
0*
09
0>
0C
#741990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#742000000000
0!
0*
09
0>
0C
#742010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#742020000000
0!
0*
09
0>
0C
#742030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#742040000000
0!
0#
0*
0,
09
0>
0?
0C
#742050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#742060000000
0!
0*
09
0>
0C
#742070000000
1!
1*
19
1>
1C
#742080000000
0!
0*
09
0>
0C
#742090000000
1!
1*
19
1>
1C
#742100000000
0!
0*
09
0>
0C
#742110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#742120000000
0!
0*
09
0>
0C
#742130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#742140000000
0!
0*
09
0>
0C
#742150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#742160000000
0!
0*
09
0>
0C
#742170000000
1!
1*
b10 6
19
1>
1C
b10 G
#742180000000
0!
0*
09
0>
0C
#742190000000
1!
1*
b11 6
19
1>
1C
b11 G
#742200000000
0!
0*
09
0>
0C
#742210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#742220000000
0!
0*
09
0>
0C
#742230000000
1!
1*
b101 6
19
1>
1C
b101 G
#742240000000
0!
0*
09
0>
0C
#742250000000
1!
1*
b110 6
19
1>
1C
b110 G
#742260000000
0!
0*
09
0>
0C
#742270000000
1!
1*
b111 6
19
1>
1C
b111 G
#742280000000
0!
0*
09
0>
0C
#742290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#742300000000
0!
0*
09
0>
0C
#742310000000
1!
1*
b1 6
19
1>
1C
b1 G
#742320000000
0!
0*
09
0>
0C
#742330000000
1!
1*
b10 6
19
1>
1C
b10 G
#742340000000
0!
0*
09
0>
0C
#742350000000
1!
1*
b11 6
19
1>
1C
b11 G
#742360000000
0!
0*
09
0>
0C
#742370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#742380000000
0!
0*
09
0>
0C
#742390000000
1!
1*
b101 6
19
1>
1C
b101 G
#742400000000
0!
0*
09
0>
0C
#742410000000
1!
1*
b110 6
19
1>
1C
b110 G
#742420000000
0!
0*
09
0>
0C
#742430000000
1!
1*
b111 6
19
1>
1C
b111 G
#742440000000
0!
0*
09
0>
0C
#742450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#742460000000
0!
0*
09
0>
0C
#742470000000
1!
1*
b1 6
19
1>
1C
b1 G
#742480000000
0!
0*
09
0>
0C
#742490000000
1!
1*
b10 6
19
1>
1C
b10 G
#742500000000
0!
0*
09
0>
0C
#742510000000
1!
1*
b11 6
19
1>
1C
b11 G
#742520000000
0!
0*
09
0>
0C
#742530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#742540000000
0!
0*
09
0>
0C
#742550000000
1!
1*
b101 6
19
1>
1C
b101 G
#742560000000
0!
0*
09
0>
0C
#742570000000
1!
1*
b110 6
19
1>
1C
b110 G
#742580000000
0!
0*
09
0>
0C
#742590000000
1!
1*
b111 6
19
1>
1C
b111 G
#742600000000
0!
1"
0*
1+
09
1:
0>
0C
#742610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#742620000000
0!
0*
09
0>
0C
#742630000000
1!
1*
b1 6
19
1>
1C
b1 G
#742640000000
0!
0*
09
0>
0C
#742650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#742660000000
0!
0*
09
0>
0C
#742670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#742680000000
0!
0*
09
0>
0C
#742690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#742700000000
0!
0*
09
0>
0C
#742710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#742720000000
0!
0#
0*
0,
09
0>
0?
0C
#742730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#742740000000
0!
0*
09
0>
0C
#742750000000
1!
1*
19
1>
1C
#742760000000
0!
0*
09
0>
0C
#742770000000
1!
1*
19
1>
1C
#742780000000
0!
0*
09
0>
0C
#742790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#742800000000
0!
0*
09
0>
0C
#742810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#742820000000
0!
0*
09
0>
0C
#742830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#742840000000
0!
0*
09
0>
0C
#742850000000
1!
1*
b10 6
19
1>
1C
b10 G
#742860000000
0!
0*
09
0>
0C
#742870000000
1!
1*
b11 6
19
1>
1C
b11 G
#742880000000
0!
0*
09
0>
0C
#742890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#742900000000
0!
0*
09
0>
0C
#742910000000
1!
1*
b101 6
19
1>
1C
b101 G
#742920000000
0!
0*
09
0>
0C
#742930000000
1!
1*
b110 6
19
1>
1C
b110 G
#742940000000
0!
0*
09
0>
0C
#742950000000
1!
1*
b111 6
19
1>
1C
b111 G
#742960000000
0!
0*
09
0>
0C
#742970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#742980000000
0!
0*
09
0>
0C
#742990000000
1!
1*
b1 6
19
1>
1C
b1 G
#743000000000
0!
0*
09
0>
0C
#743010000000
1!
1*
b10 6
19
1>
1C
b10 G
#743020000000
0!
0*
09
0>
0C
#743030000000
1!
1*
b11 6
19
1>
1C
b11 G
#743040000000
0!
0*
09
0>
0C
#743050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#743060000000
0!
0*
09
0>
0C
#743070000000
1!
1*
b101 6
19
1>
1C
b101 G
#743080000000
0!
0*
09
0>
0C
#743090000000
1!
1*
b110 6
19
1>
1C
b110 G
#743100000000
0!
0*
09
0>
0C
#743110000000
1!
1*
b111 6
19
1>
1C
b111 G
#743120000000
0!
0*
09
0>
0C
#743130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#743140000000
0!
0*
09
0>
0C
#743150000000
1!
1*
b1 6
19
1>
1C
b1 G
#743160000000
0!
0*
09
0>
0C
#743170000000
1!
1*
b10 6
19
1>
1C
b10 G
#743180000000
0!
0*
09
0>
0C
#743190000000
1!
1*
b11 6
19
1>
1C
b11 G
#743200000000
0!
0*
09
0>
0C
#743210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#743220000000
0!
0*
09
0>
0C
#743230000000
1!
1*
b101 6
19
1>
1C
b101 G
#743240000000
0!
0*
09
0>
0C
#743250000000
1!
1*
b110 6
19
1>
1C
b110 G
#743260000000
0!
0*
09
0>
0C
#743270000000
1!
1*
b111 6
19
1>
1C
b111 G
#743280000000
0!
1"
0*
1+
09
1:
0>
0C
#743290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#743300000000
0!
0*
09
0>
0C
#743310000000
1!
1*
b1 6
19
1>
1C
b1 G
#743320000000
0!
0*
09
0>
0C
#743330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#743340000000
0!
0*
09
0>
0C
#743350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#743360000000
0!
0*
09
0>
0C
#743370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#743380000000
0!
0*
09
0>
0C
#743390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#743400000000
0!
0#
0*
0,
09
0>
0?
0C
#743410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#743420000000
0!
0*
09
0>
0C
#743430000000
1!
1*
19
1>
1C
#743440000000
0!
0*
09
0>
0C
#743450000000
1!
1*
19
1>
1C
#743460000000
0!
0*
09
0>
0C
#743470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#743480000000
0!
0*
09
0>
0C
#743490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#743500000000
0!
0*
09
0>
0C
#743510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#743520000000
0!
0*
09
0>
0C
#743530000000
1!
1*
b10 6
19
1>
1C
b10 G
#743540000000
0!
0*
09
0>
0C
#743550000000
1!
1*
b11 6
19
1>
1C
b11 G
#743560000000
0!
0*
09
0>
0C
#743570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#743580000000
0!
0*
09
0>
0C
#743590000000
1!
1*
b101 6
19
1>
1C
b101 G
#743600000000
0!
0*
09
0>
0C
#743610000000
1!
1*
b110 6
19
1>
1C
b110 G
#743620000000
0!
0*
09
0>
0C
#743630000000
1!
1*
b111 6
19
1>
1C
b111 G
#743640000000
0!
0*
09
0>
0C
#743650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#743660000000
0!
0*
09
0>
0C
#743670000000
1!
1*
b1 6
19
1>
1C
b1 G
#743680000000
0!
0*
09
0>
0C
#743690000000
1!
1*
b10 6
19
1>
1C
b10 G
#743700000000
0!
0*
09
0>
0C
#743710000000
1!
1*
b11 6
19
1>
1C
b11 G
#743720000000
0!
0*
09
0>
0C
#743730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#743740000000
0!
0*
09
0>
0C
#743750000000
1!
1*
b101 6
19
1>
1C
b101 G
#743760000000
0!
0*
09
0>
0C
#743770000000
1!
1*
b110 6
19
1>
1C
b110 G
#743780000000
0!
0*
09
0>
0C
#743790000000
1!
1*
b111 6
19
1>
1C
b111 G
#743800000000
0!
0*
09
0>
0C
#743810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#743820000000
0!
0*
09
0>
0C
#743830000000
1!
1*
b1 6
19
1>
1C
b1 G
#743840000000
0!
0*
09
0>
0C
#743850000000
1!
1*
b10 6
19
1>
1C
b10 G
#743860000000
0!
0*
09
0>
0C
#743870000000
1!
1*
b11 6
19
1>
1C
b11 G
#743880000000
0!
0*
09
0>
0C
#743890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#743900000000
0!
0*
09
0>
0C
#743910000000
1!
1*
b101 6
19
1>
1C
b101 G
#743920000000
0!
0*
09
0>
0C
#743930000000
1!
1*
b110 6
19
1>
1C
b110 G
#743940000000
0!
0*
09
0>
0C
#743950000000
1!
1*
b111 6
19
1>
1C
b111 G
#743960000000
0!
1"
0*
1+
09
1:
0>
0C
#743970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#743980000000
0!
0*
09
0>
0C
#743990000000
1!
1*
b1 6
19
1>
1C
b1 G
#744000000000
0!
0*
09
0>
0C
#744010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#744020000000
0!
0*
09
0>
0C
#744030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#744040000000
0!
0*
09
0>
0C
#744050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#744060000000
0!
0*
09
0>
0C
#744070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#744080000000
0!
0#
0*
0,
09
0>
0?
0C
#744090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#744100000000
0!
0*
09
0>
0C
#744110000000
1!
1*
19
1>
1C
#744120000000
0!
0*
09
0>
0C
#744130000000
1!
1*
19
1>
1C
#744140000000
0!
0*
09
0>
0C
#744150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#744160000000
0!
0*
09
0>
0C
#744170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#744180000000
0!
0*
09
0>
0C
#744190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#744200000000
0!
0*
09
0>
0C
#744210000000
1!
1*
b10 6
19
1>
1C
b10 G
#744220000000
0!
0*
09
0>
0C
#744230000000
1!
1*
b11 6
19
1>
1C
b11 G
#744240000000
0!
0*
09
0>
0C
#744250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#744260000000
0!
0*
09
0>
0C
#744270000000
1!
1*
b101 6
19
1>
1C
b101 G
#744280000000
0!
0*
09
0>
0C
#744290000000
1!
1*
b110 6
19
1>
1C
b110 G
#744300000000
0!
0*
09
0>
0C
#744310000000
1!
1*
b111 6
19
1>
1C
b111 G
#744320000000
0!
0*
09
0>
0C
#744330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#744340000000
0!
0*
09
0>
0C
#744350000000
1!
1*
b1 6
19
1>
1C
b1 G
#744360000000
0!
0*
09
0>
0C
#744370000000
1!
1*
b10 6
19
1>
1C
b10 G
#744380000000
0!
0*
09
0>
0C
#744390000000
1!
1*
b11 6
19
1>
1C
b11 G
#744400000000
0!
0*
09
0>
0C
#744410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#744420000000
0!
0*
09
0>
0C
#744430000000
1!
1*
b101 6
19
1>
1C
b101 G
#744440000000
0!
0*
09
0>
0C
#744450000000
1!
1*
b110 6
19
1>
1C
b110 G
#744460000000
0!
0*
09
0>
0C
#744470000000
1!
1*
b111 6
19
1>
1C
b111 G
#744480000000
0!
0*
09
0>
0C
#744490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#744500000000
0!
0*
09
0>
0C
#744510000000
1!
1*
b1 6
19
1>
1C
b1 G
#744520000000
0!
0*
09
0>
0C
#744530000000
1!
1*
b10 6
19
1>
1C
b10 G
#744540000000
0!
0*
09
0>
0C
#744550000000
1!
1*
b11 6
19
1>
1C
b11 G
#744560000000
0!
0*
09
0>
0C
#744570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#744580000000
0!
0*
09
0>
0C
#744590000000
1!
1*
b101 6
19
1>
1C
b101 G
#744600000000
0!
0*
09
0>
0C
#744610000000
1!
1*
b110 6
19
1>
1C
b110 G
#744620000000
0!
0*
09
0>
0C
#744630000000
1!
1*
b111 6
19
1>
1C
b111 G
#744640000000
0!
1"
0*
1+
09
1:
0>
0C
#744650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#744660000000
0!
0*
09
0>
0C
#744670000000
1!
1*
b1 6
19
1>
1C
b1 G
#744680000000
0!
0*
09
0>
0C
#744690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#744700000000
0!
0*
09
0>
0C
#744710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#744720000000
0!
0*
09
0>
0C
#744730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#744740000000
0!
0*
09
0>
0C
#744750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#744760000000
0!
0#
0*
0,
09
0>
0?
0C
#744770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#744780000000
0!
0*
09
0>
0C
#744790000000
1!
1*
19
1>
1C
#744800000000
0!
0*
09
0>
0C
#744810000000
1!
1*
19
1>
1C
#744820000000
0!
0*
09
0>
0C
#744830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#744840000000
0!
0*
09
0>
0C
#744850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#744860000000
0!
0*
09
0>
0C
#744870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#744880000000
0!
0*
09
0>
0C
#744890000000
1!
1*
b10 6
19
1>
1C
b10 G
#744900000000
0!
0*
09
0>
0C
#744910000000
1!
1*
b11 6
19
1>
1C
b11 G
#744920000000
0!
0*
09
0>
0C
#744930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#744940000000
0!
0*
09
0>
0C
#744950000000
1!
1*
b101 6
19
1>
1C
b101 G
#744960000000
0!
0*
09
0>
0C
#744970000000
1!
1*
b110 6
19
1>
1C
b110 G
#744980000000
0!
0*
09
0>
0C
#744990000000
1!
1*
b111 6
19
1>
1C
b111 G
#745000000000
0!
0*
09
0>
0C
#745010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#745020000000
0!
0*
09
0>
0C
#745030000000
1!
1*
b1 6
19
1>
1C
b1 G
#745040000000
0!
0*
09
0>
0C
#745050000000
1!
1*
b10 6
19
1>
1C
b10 G
#745060000000
0!
0*
09
0>
0C
#745070000000
1!
1*
b11 6
19
1>
1C
b11 G
#745080000000
0!
0*
09
0>
0C
#745090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#745100000000
0!
0*
09
0>
0C
#745110000000
1!
1*
b101 6
19
1>
1C
b101 G
#745120000000
0!
0*
09
0>
0C
#745130000000
1!
1*
b110 6
19
1>
1C
b110 G
#745140000000
0!
0*
09
0>
0C
#745150000000
1!
1*
b111 6
19
1>
1C
b111 G
#745160000000
0!
0*
09
0>
0C
#745170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#745180000000
0!
0*
09
0>
0C
#745190000000
1!
1*
b1 6
19
1>
1C
b1 G
#745200000000
0!
0*
09
0>
0C
#745210000000
1!
1*
b10 6
19
1>
1C
b10 G
#745220000000
0!
0*
09
0>
0C
#745230000000
1!
1*
b11 6
19
1>
1C
b11 G
#745240000000
0!
0*
09
0>
0C
#745250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#745260000000
0!
0*
09
0>
0C
#745270000000
1!
1*
b101 6
19
1>
1C
b101 G
#745280000000
0!
0*
09
0>
0C
#745290000000
1!
1*
b110 6
19
1>
1C
b110 G
#745300000000
0!
0*
09
0>
0C
#745310000000
1!
1*
b111 6
19
1>
1C
b111 G
#745320000000
0!
1"
0*
1+
09
1:
0>
0C
#745330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#745340000000
0!
0*
09
0>
0C
#745350000000
1!
1*
b1 6
19
1>
1C
b1 G
#745360000000
0!
0*
09
0>
0C
#745370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#745380000000
0!
0*
09
0>
0C
#745390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#745400000000
0!
0*
09
0>
0C
#745410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#745420000000
0!
0*
09
0>
0C
#745430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#745440000000
0!
0#
0*
0,
09
0>
0?
0C
#745450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#745460000000
0!
0*
09
0>
0C
#745470000000
1!
1*
19
1>
1C
#745480000000
0!
0*
09
0>
0C
#745490000000
1!
1*
19
1>
1C
#745500000000
0!
0*
09
0>
0C
#745510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#745520000000
0!
0*
09
0>
0C
#745530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#745540000000
0!
0*
09
0>
0C
#745550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#745560000000
0!
0*
09
0>
0C
#745570000000
1!
1*
b10 6
19
1>
1C
b10 G
#745580000000
0!
0*
09
0>
0C
#745590000000
1!
1*
b11 6
19
1>
1C
b11 G
#745600000000
0!
0*
09
0>
0C
#745610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#745620000000
0!
0*
09
0>
0C
#745630000000
1!
1*
b101 6
19
1>
1C
b101 G
#745640000000
0!
0*
09
0>
0C
#745650000000
1!
1*
b110 6
19
1>
1C
b110 G
#745660000000
0!
0*
09
0>
0C
#745670000000
1!
1*
b111 6
19
1>
1C
b111 G
#745680000000
0!
0*
09
0>
0C
#745690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#745700000000
0!
0*
09
0>
0C
#745710000000
1!
1*
b1 6
19
1>
1C
b1 G
#745720000000
0!
0*
09
0>
0C
#745730000000
1!
1*
b10 6
19
1>
1C
b10 G
#745740000000
0!
0*
09
0>
0C
#745750000000
1!
1*
b11 6
19
1>
1C
b11 G
#745760000000
0!
0*
09
0>
0C
#745770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#745780000000
0!
0*
09
0>
0C
#745790000000
1!
1*
b101 6
19
1>
1C
b101 G
#745800000000
0!
0*
09
0>
0C
#745810000000
1!
1*
b110 6
19
1>
1C
b110 G
#745820000000
0!
0*
09
0>
0C
#745830000000
1!
1*
b111 6
19
1>
1C
b111 G
#745840000000
0!
0*
09
0>
0C
#745850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#745860000000
0!
0*
09
0>
0C
#745870000000
1!
1*
b1 6
19
1>
1C
b1 G
#745880000000
0!
0*
09
0>
0C
#745890000000
1!
1*
b10 6
19
1>
1C
b10 G
#745900000000
0!
0*
09
0>
0C
#745910000000
1!
1*
b11 6
19
1>
1C
b11 G
#745920000000
0!
0*
09
0>
0C
#745930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#745940000000
0!
0*
09
0>
0C
#745950000000
1!
1*
b101 6
19
1>
1C
b101 G
#745960000000
0!
0*
09
0>
0C
#745970000000
1!
1*
b110 6
19
1>
1C
b110 G
#745980000000
0!
0*
09
0>
0C
#745990000000
1!
1*
b111 6
19
1>
1C
b111 G
#746000000000
0!
1"
0*
1+
09
1:
0>
0C
#746010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#746020000000
0!
0*
09
0>
0C
#746030000000
1!
1*
b1 6
19
1>
1C
b1 G
#746040000000
0!
0*
09
0>
0C
#746050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#746060000000
0!
0*
09
0>
0C
#746070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#746080000000
0!
0*
09
0>
0C
#746090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#746100000000
0!
0*
09
0>
0C
#746110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#746120000000
0!
0#
0*
0,
09
0>
0?
0C
#746130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#746140000000
0!
0*
09
0>
0C
#746150000000
1!
1*
19
1>
1C
#746160000000
0!
0*
09
0>
0C
#746170000000
1!
1*
19
1>
1C
#746180000000
0!
0*
09
0>
0C
#746190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#746200000000
0!
0*
09
0>
0C
#746210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#746220000000
0!
0*
09
0>
0C
#746230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#746240000000
0!
0*
09
0>
0C
#746250000000
1!
1*
b10 6
19
1>
1C
b10 G
#746260000000
0!
0*
09
0>
0C
#746270000000
1!
1*
b11 6
19
1>
1C
b11 G
#746280000000
0!
0*
09
0>
0C
#746290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#746300000000
0!
0*
09
0>
0C
#746310000000
1!
1*
b101 6
19
1>
1C
b101 G
#746320000000
0!
0*
09
0>
0C
#746330000000
1!
1*
b110 6
19
1>
1C
b110 G
#746340000000
0!
0*
09
0>
0C
#746350000000
1!
1*
b111 6
19
1>
1C
b111 G
#746360000000
0!
0*
09
0>
0C
#746370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#746380000000
0!
0*
09
0>
0C
#746390000000
1!
1*
b1 6
19
1>
1C
b1 G
#746400000000
0!
0*
09
0>
0C
#746410000000
1!
1*
b10 6
19
1>
1C
b10 G
#746420000000
0!
0*
09
0>
0C
#746430000000
1!
1*
b11 6
19
1>
1C
b11 G
#746440000000
0!
0*
09
0>
0C
#746450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#746460000000
0!
0*
09
0>
0C
#746470000000
1!
1*
b101 6
19
1>
1C
b101 G
#746480000000
0!
0*
09
0>
0C
#746490000000
1!
1*
b110 6
19
1>
1C
b110 G
#746500000000
0!
0*
09
0>
0C
#746510000000
1!
1*
b111 6
19
1>
1C
b111 G
#746520000000
0!
0*
09
0>
0C
#746530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#746540000000
0!
0*
09
0>
0C
#746550000000
1!
1*
b1 6
19
1>
1C
b1 G
#746560000000
0!
0*
09
0>
0C
#746570000000
1!
1*
b10 6
19
1>
1C
b10 G
#746580000000
0!
0*
09
0>
0C
#746590000000
1!
1*
b11 6
19
1>
1C
b11 G
#746600000000
0!
0*
09
0>
0C
#746610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#746620000000
0!
0*
09
0>
0C
#746630000000
1!
1*
b101 6
19
1>
1C
b101 G
#746640000000
0!
0*
09
0>
0C
#746650000000
1!
1*
b110 6
19
1>
1C
b110 G
#746660000000
0!
0*
09
0>
0C
#746670000000
1!
1*
b111 6
19
1>
1C
b111 G
#746680000000
0!
1"
0*
1+
09
1:
0>
0C
#746690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#746700000000
0!
0*
09
0>
0C
#746710000000
1!
1*
b1 6
19
1>
1C
b1 G
#746720000000
0!
0*
09
0>
0C
#746730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#746740000000
0!
0*
09
0>
0C
#746750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#746760000000
0!
0*
09
0>
0C
#746770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#746780000000
0!
0*
09
0>
0C
#746790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#746800000000
0!
0#
0*
0,
09
0>
0?
0C
#746810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#746820000000
0!
0*
09
0>
0C
#746830000000
1!
1*
19
1>
1C
#746840000000
0!
0*
09
0>
0C
#746850000000
1!
1*
19
1>
1C
#746860000000
0!
0*
09
0>
0C
#746870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#746880000000
0!
0*
09
0>
0C
#746890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#746900000000
0!
0*
09
0>
0C
#746910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#746920000000
0!
0*
09
0>
0C
#746930000000
1!
1*
b10 6
19
1>
1C
b10 G
#746940000000
0!
0*
09
0>
0C
#746950000000
1!
1*
b11 6
19
1>
1C
b11 G
#746960000000
0!
0*
09
0>
0C
#746970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#746980000000
0!
0*
09
0>
0C
#746990000000
1!
1*
b101 6
19
1>
1C
b101 G
#747000000000
0!
0*
09
0>
0C
#747010000000
1!
1*
b110 6
19
1>
1C
b110 G
#747020000000
0!
0*
09
0>
0C
#747030000000
1!
1*
b111 6
19
1>
1C
b111 G
#747040000000
0!
0*
09
0>
0C
#747050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#747060000000
0!
0*
09
0>
0C
#747070000000
1!
1*
b1 6
19
1>
1C
b1 G
#747080000000
0!
0*
09
0>
0C
#747090000000
1!
1*
b10 6
19
1>
1C
b10 G
#747100000000
0!
0*
09
0>
0C
#747110000000
1!
1*
b11 6
19
1>
1C
b11 G
#747120000000
0!
0*
09
0>
0C
#747130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#747140000000
0!
0*
09
0>
0C
#747150000000
1!
1*
b101 6
19
1>
1C
b101 G
#747160000000
0!
0*
09
0>
0C
#747170000000
1!
1*
b110 6
19
1>
1C
b110 G
#747180000000
0!
0*
09
0>
0C
#747190000000
1!
1*
b111 6
19
1>
1C
b111 G
#747200000000
0!
0*
09
0>
0C
#747210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#747220000000
0!
0*
09
0>
0C
#747230000000
1!
1*
b1 6
19
1>
1C
b1 G
#747240000000
0!
0*
09
0>
0C
#747250000000
1!
1*
b10 6
19
1>
1C
b10 G
#747260000000
0!
0*
09
0>
0C
#747270000000
1!
1*
b11 6
19
1>
1C
b11 G
#747280000000
0!
0*
09
0>
0C
#747290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#747300000000
0!
0*
09
0>
0C
#747310000000
1!
1*
b101 6
19
1>
1C
b101 G
#747320000000
0!
0*
09
0>
0C
#747330000000
1!
1*
b110 6
19
1>
1C
b110 G
#747340000000
0!
0*
09
0>
0C
#747350000000
1!
1*
b111 6
19
1>
1C
b111 G
#747360000000
0!
1"
0*
1+
09
1:
0>
0C
#747370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#747380000000
0!
0*
09
0>
0C
#747390000000
1!
1*
b1 6
19
1>
1C
b1 G
#747400000000
0!
0*
09
0>
0C
#747410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#747420000000
0!
0*
09
0>
0C
#747430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#747440000000
0!
0*
09
0>
0C
#747450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#747460000000
0!
0*
09
0>
0C
#747470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#747480000000
0!
0#
0*
0,
09
0>
0?
0C
#747490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#747500000000
0!
0*
09
0>
0C
#747510000000
1!
1*
19
1>
1C
#747520000000
0!
0*
09
0>
0C
#747530000000
1!
1*
19
1>
1C
#747540000000
0!
0*
09
0>
0C
#747550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#747560000000
0!
0*
09
0>
0C
#747570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#747580000000
0!
0*
09
0>
0C
#747590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#747600000000
0!
0*
09
0>
0C
#747610000000
1!
1*
b10 6
19
1>
1C
b10 G
#747620000000
0!
0*
09
0>
0C
#747630000000
1!
1*
b11 6
19
1>
1C
b11 G
#747640000000
0!
0*
09
0>
0C
#747650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#747660000000
0!
0*
09
0>
0C
#747670000000
1!
1*
b101 6
19
1>
1C
b101 G
#747680000000
0!
0*
09
0>
0C
#747690000000
1!
1*
b110 6
19
1>
1C
b110 G
#747700000000
0!
0*
09
0>
0C
#747710000000
1!
1*
b111 6
19
1>
1C
b111 G
#747720000000
0!
0*
09
0>
0C
#747730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#747740000000
0!
0*
09
0>
0C
#747750000000
1!
1*
b1 6
19
1>
1C
b1 G
#747760000000
0!
0*
09
0>
0C
#747770000000
1!
1*
b10 6
19
1>
1C
b10 G
#747780000000
0!
0*
09
0>
0C
#747790000000
1!
1*
b11 6
19
1>
1C
b11 G
#747800000000
0!
0*
09
0>
0C
#747810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#747820000000
0!
0*
09
0>
0C
#747830000000
1!
1*
b101 6
19
1>
1C
b101 G
#747840000000
0!
0*
09
0>
0C
#747850000000
1!
1*
b110 6
19
1>
1C
b110 G
#747860000000
0!
0*
09
0>
0C
#747870000000
1!
1*
b111 6
19
1>
1C
b111 G
#747880000000
0!
0*
09
0>
0C
#747890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#747900000000
0!
0*
09
0>
0C
#747910000000
1!
1*
b1 6
19
1>
1C
b1 G
#747920000000
0!
0*
09
0>
0C
#747930000000
1!
1*
b10 6
19
1>
1C
b10 G
#747940000000
0!
0*
09
0>
0C
#747950000000
1!
1*
b11 6
19
1>
1C
b11 G
#747960000000
0!
0*
09
0>
0C
#747970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#747980000000
0!
0*
09
0>
0C
#747990000000
1!
1*
b101 6
19
1>
1C
b101 G
#748000000000
0!
0*
09
0>
0C
#748010000000
1!
1*
b110 6
19
1>
1C
b110 G
#748020000000
0!
0*
09
0>
0C
#748030000000
1!
1*
b111 6
19
1>
1C
b111 G
#748040000000
0!
1"
0*
1+
09
1:
0>
0C
#748050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#748060000000
0!
0*
09
0>
0C
#748070000000
1!
1*
b1 6
19
1>
1C
b1 G
#748080000000
0!
0*
09
0>
0C
#748090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#748100000000
0!
0*
09
0>
0C
#748110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#748120000000
0!
0*
09
0>
0C
#748130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#748140000000
0!
0*
09
0>
0C
#748150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#748160000000
0!
0#
0*
0,
09
0>
0?
0C
#748170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#748180000000
0!
0*
09
0>
0C
#748190000000
1!
1*
19
1>
1C
#748200000000
0!
0*
09
0>
0C
#748210000000
1!
1*
19
1>
1C
#748220000000
0!
0*
09
0>
0C
#748230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#748240000000
0!
0*
09
0>
0C
#748250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#748260000000
0!
0*
09
0>
0C
#748270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#748280000000
0!
0*
09
0>
0C
#748290000000
1!
1*
b10 6
19
1>
1C
b10 G
#748300000000
0!
0*
09
0>
0C
#748310000000
1!
1*
b11 6
19
1>
1C
b11 G
#748320000000
0!
0*
09
0>
0C
#748330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#748340000000
0!
0*
09
0>
0C
#748350000000
1!
1*
b101 6
19
1>
1C
b101 G
#748360000000
0!
0*
09
0>
0C
#748370000000
1!
1*
b110 6
19
1>
1C
b110 G
#748380000000
0!
0*
09
0>
0C
#748390000000
1!
1*
b111 6
19
1>
1C
b111 G
#748400000000
0!
0*
09
0>
0C
#748410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#748420000000
0!
0*
09
0>
0C
#748430000000
1!
1*
b1 6
19
1>
1C
b1 G
#748440000000
0!
0*
09
0>
0C
#748450000000
1!
1*
b10 6
19
1>
1C
b10 G
#748460000000
0!
0*
09
0>
0C
#748470000000
1!
1*
b11 6
19
1>
1C
b11 G
#748480000000
0!
0*
09
0>
0C
#748490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#748500000000
0!
0*
09
0>
0C
#748510000000
1!
1*
b101 6
19
1>
1C
b101 G
#748520000000
0!
0*
09
0>
0C
#748530000000
1!
1*
b110 6
19
1>
1C
b110 G
#748540000000
0!
0*
09
0>
0C
#748550000000
1!
1*
b111 6
19
1>
1C
b111 G
#748560000000
0!
0*
09
0>
0C
#748570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#748580000000
0!
0*
09
0>
0C
#748590000000
1!
1*
b1 6
19
1>
1C
b1 G
#748600000000
0!
0*
09
0>
0C
#748610000000
1!
1*
b10 6
19
1>
1C
b10 G
#748620000000
0!
0*
09
0>
0C
#748630000000
1!
1*
b11 6
19
1>
1C
b11 G
#748640000000
0!
0*
09
0>
0C
#748650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#748660000000
0!
0*
09
0>
0C
#748670000000
1!
1*
b101 6
19
1>
1C
b101 G
#748680000000
0!
0*
09
0>
0C
#748690000000
1!
1*
b110 6
19
1>
1C
b110 G
#748700000000
0!
0*
09
0>
0C
#748710000000
1!
1*
b111 6
19
1>
1C
b111 G
#748720000000
0!
1"
0*
1+
09
1:
0>
0C
#748730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#748740000000
0!
0*
09
0>
0C
#748750000000
1!
1*
b1 6
19
1>
1C
b1 G
#748760000000
0!
0*
09
0>
0C
#748770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#748780000000
0!
0*
09
0>
0C
#748790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#748800000000
0!
0*
09
0>
0C
#748810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#748820000000
0!
0*
09
0>
0C
#748830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#748840000000
0!
0#
0*
0,
09
0>
0?
0C
#748850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#748860000000
0!
0*
09
0>
0C
#748870000000
1!
1*
19
1>
1C
#748880000000
0!
0*
09
0>
0C
#748890000000
1!
1*
19
1>
1C
#748900000000
0!
0*
09
0>
0C
#748910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#748920000000
0!
0*
09
0>
0C
#748930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#748940000000
0!
0*
09
0>
0C
#748950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#748960000000
0!
0*
09
0>
0C
#748970000000
1!
1*
b10 6
19
1>
1C
b10 G
#748980000000
0!
0*
09
0>
0C
#748990000000
1!
1*
b11 6
19
1>
1C
b11 G
#749000000000
0!
0*
09
0>
0C
#749010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#749020000000
0!
0*
09
0>
0C
#749030000000
1!
1*
b101 6
19
1>
1C
b101 G
#749040000000
0!
0*
09
0>
0C
#749050000000
1!
1*
b110 6
19
1>
1C
b110 G
#749060000000
0!
0*
09
0>
0C
#749070000000
1!
1*
b111 6
19
1>
1C
b111 G
#749080000000
0!
0*
09
0>
0C
#749090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#749100000000
0!
0*
09
0>
0C
#749110000000
1!
1*
b1 6
19
1>
1C
b1 G
#749120000000
0!
0*
09
0>
0C
#749130000000
1!
1*
b10 6
19
1>
1C
b10 G
#749140000000
0!
0*
09
0>
0C
#749150000000
1!
1*
b11 6
19
1>
1C
b11 G
#749160000000
0!
0*
09
0>
0C
#749170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#749180000000
0!
0*
09
0>
0C
#749190000000
1!
1*
b101 6
19
1>
1C
b101 G
#749200000000
0!
0*
09
0>
0C
#749210000000
1!
1*
b110 6
19
1>
1C
b110 G
#749220000000
0!
0*
09
0>
0C
#749230000000
1!
1*
b111 6
19
1>
1C
b111 G
#749240000000
0!
0*
09
0>
0C
#749250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#749260000000
0!
0*
09
0>
0C
#749270000000
1!
1*
b1 6
19
1>
1C
b1 G
#749280000000
0!
0*
09
0>
0C
#749290000000
1!
1*
b10 6
19
1>
1C
b10 G
#749300000000
0!
0*
09
0>
0C
#749310000000
1!
1*
b11 6
19
1>
1C
b11 G
#749320000000
0!
0*
09
0>
0C
#749330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#749340000000
0!
0*
09
0>
0C
#749350000000
1!
1*
b101 6
19
1>
1C
b101 G
#749360000000
0!
0*
09
0>
0C
#749370000000
1!
1*
b110 6
19
1>
1C
b110 G
#749380000000
0!
0*
09
0>
0C
#749390000000
1!
1*
b111 6
19
1>
1C
b111 G
#749400000000
0!
1"
0*
1+
09
1:
0>
0C
#749410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#749420000000
0!
0*
09
0>
0C
#749430000000
1!
1*
b1 6
19
1>
1C
b1 G
#749440000000
0!
0*
09
0>
0C
#749450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#749460000000
0!
0*
09
0>
0C
#749470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#749480000000
0!
0*
09
0>
0C
#749490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#749500000000
0!
0*
09
0>
0C
#749510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#749520000000
0!
0#
0*
0,
09
0>
0?
0C
#749530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#749540000000
0!
0*
09
0>
0C
#749550000000
1!
1*
19
1>
1C
#749560000000
0!
0*
09
0>
0C
#749570000000
1!
1*
19
1>
1C
#749580000000
0!
0*
09
0>
0C
#749590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#749600000000
0!
0*
09
0>
0C
#749610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#749620000000
0!
0*
09
0>
0C
#749630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#749640000000
0!
0*
09
0>
0C
#749650000000
1!
1*
b10 6
19
1>
1C
b10 G
#749660000000
0!
0*
09
0>
0C
#749670000000
1!
1*
b11 6
19
1>
1C
b11 G
#749680000000
0!
0*
09
0>
0C
#749690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#749700000000
0!
0*
09
0>
0C
#749710000000
1!
1*
b101 6
19
1>
1C
b101 G
#749720000000
0!
0*
09
0>
0C
#749730000000
1!
1*
b110 6
19
1>
1C
b110 G
#749740000000
0!
0*
09
0>
0C
#749750000000
1!
1*
b111 6
19
1>
1C
b111 G
#749760000000
0!
0*
09
0>
0C
#749770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#749780000000
0!
0*
09
0>
0C
#749790000000
1!
1*
b1 6
19
1>
1C
b1 G
#749800000000
0!
0*
09
0>
0C
#749810000000
1!
1*
b10 6
19
1>
1C
b10 G
#749820000000
0!
0*
09
0>
0C
#749830000000
1!
1*
b11 6
19
1>
1C
b11 G
#749840000000
0!
0*
09
0>
0C
#749850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#749860000000
0!
0*
09
0>
0C
#749870000000
1!
1*
b101 6
19
1>
1C
b101 G
#749880000000
0!
0*
09
0>
0C
#749890000000
1!
1*
b110 6
19
1>
1C
b110 G
#749900000000
0!
0*
09
0>
0C
#749910000000
1!
1*
b111 6
19
1>
1C
b111 G
#749920000000
0!
0*
09
0>
0C
#749930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#749940000000
0!
0*
09
0>
0C
#749950000000
1!
1*
b1 6
19
1>
1C
b1 G
#749960000000
0!
0*
09
0>
0C
#749970000000
1!
1*
b10 6
19
1>
1C
b10 G
#749980000000
0!
0*
09
0>
0C
#749990000000
1!
1*
b11 6
19
1>
1C
b11 G
#750000000000
0!
0*
09
0>
0C
#750010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#750020000000
0!
0*
09
0>
0C
#750030000000
1!
1*
b101 6
19
1>
1C
b101 G
#750040000000
0!
0*
09
0>
0C
#750050000000
1!
1*
b110 6
19
1>
1C
b110 G
#750060000000
0!
0*
09
0>
0C
#750070000000
1!
1*
b111 6
19
1>
1C
b111 G
#750080000000
0!
1"
0*
1+
09
1:
0>
0C
#750090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#750100000000
0!
0*
09
0>
0C
#750110000000
1!
1*
b1 6
19
1>
1C
b1 G
#750120000000
0!
0*
09
0>
0C
#750130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#750140000000
0!
0*
09
0>
0C
#750150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#750160000000
0!
0*
09
0>
0C
#750170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#750180000000
0!
0*
09
0>
0C
#750190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#750200000000
0!
0#
0*
0,
09
0>
0?
0C
#750210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#750220000000
0!
0*
09
0>
0C
#750230000000
1!
1*
19
1>
1C
#750240000000
0!
0*
09
0>
0C
#750250000000
1!
1*
19
1>
1C
#750260000000
0!
0*
09
0>
0C
#750270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#750280000000
0!
0*
09
0>
0C
#750290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#750300000000
0!
0*
09
0>
0C
#750310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#750320000000
0!
0*
09
0>
0C
#750330000000
1!
1*
b10 6
19
1>
1C
b10 G
#750340000000
0!
0*
09
0>
0C
#750350000000
1!
1*
b11 6
19
1>
1C
b11 G
#750360000000
0!
0*
09
0>
0C
#750370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#750380000000
0!
0*
09
0>
0C
#750390000000
1!
1*
b101 6
19
1>
1C
b101 G
#750400000000
0!
0*
09
0>
0C
#750410000000
1!
1*
b110 6
19
1>
1C
b110 G
#750420000000
0!
0*
09
0>
0C
#750430000000
1!
1*
b111 6
19
1>
1C
b111 G
#750440000000
0!
0*
09
0>
0C
#750450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#750460000000
0!
0*
09
0>
0C
#750470000000
1!
1*
b1 6
19
1>
1C
b1 G
#750480000000
0!
0*
09
0>
0C
#750490000000
1!
1*
b10 6
19
1>
1C
b10 G
#750500000000
0!
0*
09
0>
0C
#750510000000
1!
1*
b11 6
19
1>
1C
b11 G
#750520000000
0!
0*
09
0>
0C
#750530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#750540000000
0!
0*
09
0>
0C
#750550000000
1!
1*
b101 6
19
1>
1C
b101 G
#750560000000
0!
0*
09
0>
0C
#750570000000
1!
1*
b110 6
19
1>
1C
b110 G
#750580000000
0!
0*
09
0>
0C
#750590000000
1!
1*
b111 6
19
1>
1C
b111 G
#750600000000
0!
0*
09
0>
0C
#750610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#750620000000
0!
0*
09
0>
0C
#750630000000
1!
1*
b1 6
19
1>
1C
b1 G
#750640000000
0!
0*
09
0>
0C
#750650000000
1!
1*
b10 6
19
1>
1C
b10 G
#750660000000
0!
0*
09
0>
0C
#750670000000
1!
1*
b11 6
19
1>
1C
b11 G
#750680000000
0!
0*
09
0>
0C
#750690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#750700000000
0!
0*
09
0>
0C
#750710000000
1!
1*
b101 6
19
1>
1C
b101 G
#750720000000
0!
0*
09
0>
0C
#750730000000
1!
1*
b110 6
19
1>
1C
b110 G
#750740000000
0!
0*
09
0>
0C
#750750000000
1!
1*
b111 6
19
1>
1C
b111 G
#750760000000
0!
1"
0*
1+
09
1:
0>
0C
#750770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#750780000000
0!
0*
09
0>
0C
#750790000000
1!
1*
b1 6
19
1>
1C
b1 G
#750800000000
0!
0*
09
0>
0C
#750810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#750820000000
0!
0*
09
0>
0C
#750830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#750840000000
0!
0*
09
0>
0C
#750850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#750860000000
0!
0*
09
0>
0C
#750870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#750880000000
0!
0#
0*
0,
09
0>
0?
0C
#750890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#750900000000
0!
0*
09
0>
0C
#750910000000
1!
1*
19
1>
1C
#750920000000
0!
0*
09
0>
0C
#750930000000
1!
1*
19
1>
1C
#750940000000
0!
0*
09
0>
0C
#750950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#750960000000
0!
0*
09
0>
0C
#750970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#750980000000
0!
0*
09
0>
0C
#750990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#751000000000
0!
0*
09
0>
0C
#751010000000
1!
1*
b10 6
19
1>
1C
b10 G
#751020000000
0!
0*
09
0>
0C
#751030000000
1!
1*
b11 6
19
1>
1C
b11 G
#751040000000
0!
0*
09
0>
0C
#751050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#751060000000
0!
0*
09
0>
0C
#751070000000
1!
1*
b101 6
19
1>
1C
b101 G
#751080000000
0!
0*
09
0>
0C
#751090000000
1!
1*
b110 6
19
1>
1C
b110 G
#751100000000
0!
0*
09
0>
0C
#751110000000
1!
1*
b111 6
19
1>
1C
b111 G
#751120000000
0!
0*
09
0>
0C
#751130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#751140000000
0!
0*
09
0>
0C
#751150000000
1!
1*
b1 6
19
1>
1C
b1 G
#751160000000
0!
0*
09
0>
0C
#751170000000
1!
1*
b10 6
19
1>
1C
b10 G
#751180000000
0!
0*
09
0>
0C
#751190000000
1!
1*
b11 6
19
1>
1C
b11 G
#751200000000
0!
0*
09
0>
0C
#751210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#751220000000
0!
0*
09
0>
0C
#751230000000
1!
1*
b101 6
19
1>
1C
b101 G
#751240000000
0!
0*
09
0>
0C
#751250000000
1!
1*
b110 6
19
1>
1C
b110 G
#751260000000
0!
0*
09
0>
0C
#751270000000
1!
1*
b111 6
19
1>
1C
b111 G
#751280000000
0!
0*
09
0>
0C
#751290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#751300000000
0!
0*
09
0>
0C
#751310000000
1!
1*
b1 6
19
1>
1C
b1 G
#751320000000
0!
0*
09
0>
0C
#751330000000
1!
1*
b10 6
19
1>
1C
b10 G
#751340000000
0!
0*
09
0>
0C
#751350000000
1!
1*
b11 6
19
1>
1C
b11 G
#751360000000
0!
0*
09
0>
0C
#751370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#751380000000
0!
0*
09
0>
0C
#751390000000
1!
1*
b101 6
19
1>
1C
b101 G
#751400000000
0!
0*
09
0>
0C
#751410000000
1!
1*
b110 6
19
1>
1C
b110 G
#751420000000
0!
0*
09
0>
0C
#751430000000
1!
1*
b111 6
19
1>
1C
b111 G
#751440000000
0!
1"
0*
1+
09
1:
0>
0C
#751450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#751460000000
0!
0*
09
0>
0C
#751470000000
1!
1*
b1 6
19
1>
1C
b1 G
#751480000000
0!
0*
09
0>
0C
#751490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#751500000000
0!
0*
09
0>
0C
#751510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#751520000000
0!
0*
09
0>
0C
#751530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#751540000000
0!
0*
09
0>
0C
#751550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#751560000000
0!
0#
0*
0,
09
0>
0?
0C
#751570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#751580000000
0!
0*
09
0>
0C
#751590000000
1!
1*
19
1>
1C
#751600000000
0!
0*
09
0>
0C
#751610000000
1!
1*
19
1>
1C
#751620000000
0!
0*
09
0>
0C
#751630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#751640000000
0!
0*
09
0>
0C
#751650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#751660000000
0!
0*
09
0>
0C
#751670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#751680000000
0!
0*
09
0>
0C
#751690000000
1!
1*
b10 6
19
1>
1C
b10 G
#751700000000
0!
0*
09
0>
0C
#751710000000
1!
1*
b11 6
19
1>
1C
b11 G
#751720000000
0!
0*
09
0>
0C
#751730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#751740000000
0!
0*
09
0>
0C
#751750000000
1!
1*
b101 6
19
1>
1C
b101 G
#751760000000
0!
0*
09
0>
0C
#751770000000
1!
1*
b110 6
19
1>
1C
b110 G
#751780000000
0!
0*
09
0>
0C
#751790000000
1!
1*
b111 6
19
1>
1C
b111 G
#751800000000
0!
0*
09
0>
0C
#751810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#751820000000
0!
0*
09
0>
0C
#751830000000
1!
1*
b1 6
19
1>
1C
b1 G
#751840000000
0!
0*
09
0>
0C
#751850000000
1!
1*
b10 6
19
1>
1C
b10 G
#751860000000
0!
0*
09
0>
0C
#751870000000
1!
1*
b11 6
19
1>
1C
b11 G
#751880000000
0!
0*
09
0>
0C
#751890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#751900000000
0!
0*
09
0>
0C
#751910000000
1!
1*
b101 6
19
1>
1C
b101 G
#751920000000
0!
0*
09
0>
0C
#751930000000
1!
1*
b110 6
19
1>
1C
b110 G
#751940000000
0!
0*
09
0>
0C
#751950000000
1!
1*
b111 6
19
1>
1C
b111 G
#751960000000
0!
0*
09
0>
0C
#751970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#751980000000
0!
0*
09
0>
0C
#751990000000
1!
1*
b1 6
19
1>
1C
b1 G
#752000000000
0!
0*
09
0>
0C
#752010000000
1!
1*
b10 6
19
1>
1C
b10 G
#752020000000
0!
0*
09
0>
0C
#752030000000
1!
1*
b11 6
19
1>
1C
b11 G
#752040000000
0!
0*
09
0>
0C
#752050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#752060000000
0!
0*
09
0>
0C
#752070000000
1!
1*
b101 6
19
1>
1C
b101 G
#752080000000
0!
0*
09
0>
0C
#752090000000
1!
1*
b110 6
19
1>
1C
b110 G
#752100000000
0!
0*
09
0>
0C
#752110000000
1!
1*
b111 6
19
1>
1C
b111 G
#752120000000
0!
1"
0*
1+
09
1:
0>
0C
#752130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#752140000000
0!
0*
09
0>
0C
#752150000000
1!
1*
b1 6
19
1>
1C
b1 G
#752160000000
0!
0*
09
0>
0C
#752170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#752180000000
0!
0*
09
0>
0C
#752190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#752200000000
0!
0*
09
0>
0C
#752210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#752220000000
0!
0*
09
0>
0C
#752230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#752240000000
0!
0#
0*
0,
09
0>
0?
0C
#752250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#752260000000
0!
0*
09
0>
0C
#752270000000
1!
1*
19
1>
1C
#752280000000
0!
0*
09
0>
0C
#752290000000
1!
1*
19
1>
1C
#752300000000
0!
0*
09
0>
0C
#752310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#752320000000
0!
0*
09
0>
0C
#752330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#752340000000
0!
0*
09
0>
0C
#752350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#752360000000
0!
0*
09
0>
0C
#752370000000
1!
1*
b10 6
19
1>
1C
b10 G
#752380000000
0!
0*
09
0>
0C
#752390000000
1!
1*
b11 6
19
1>
1C
b11 G
#752400000000
0!
0*
09
0>
0C
#752410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#752420000000
0!
0*
09
0>
0C
#752430000000
1!
1*
b101 6
19
1>
1C
b101 G
#752440000000
0!
0*
09
0>
0C
#752450000000
1!
1*
b110 6
19
1>
1C
b110 G
#752460000000
0!
0*
09
0>
0C
#752470000000
1!
1*
b111 6
19
1>
1C
b111 G
#752480000000
0!
0*
09
0>
0C
#752490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#752500000000
0!
0*
09
0>
0C
#752510000000
1!
1*
b1 6
19
1>
1C
b1 G
#752520000000
0!
0*
09
0>
0C
#752530000000
1!
1*
b10 6
19
1>
1C
b10 G
#752540000000
0!
0*
09
0>
0C
#752550000000
1!
1*
b11 6
19
1>
1C
b11 G
#752560000000
0!
0*
09
0>
0C
#752570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#752580000000
0!
0*
09
0>
0C
#752590000000
1!
1*
b101 6
19
1>
1C
b101 G
#752600000000
0!
0*
09
0>
0C
#752610000000
1!
1*
b110 6
19
1>
1C
b110 G
#752620000000
0!
0*
09
0>
0C
#752630000000
1!
1*
b111 6
19
1>
1C
b111 G
#752640000000
0!
0*
09
0>
0C
#752650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#752660000000
0!
0*
09
0>
0C
#752670000000
1!
1*
b1 6
19
1>
1C
b1 G
#752680000000
0!
0*
09
0>
0C
#752690000000
1!
1*
b10 6
19
1>
1C
b10 G
#752700000000
0!
0*
09
0>
0C
#752710000000
1!
1*
b11 6
19
1>
1C
b11 G
#752720000000
0!
0*
09
0>
0C
#752730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#752740000000
0!
0*
09
0>
0C
#752750000000
1!
1*
b101 6
19
1>
1C
b101 G
#752760000000
0!
0*
09
0>
0C
#752770000000
1!
1*
b110 6
19
1>
1C
b110 G
#752780000000
0!
0*
09
0>
0C
#752790000000
1!
1*
b111 6
19
1>
1C
b111 G
#752800000000
0!
1"
0*
1+
09
1:
0>
0C
#752810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#752820000000
0!
0*
09
0>
0C
#752830000000
1!
1*
b1 6
19
1>
1C
b1 G
#752840000000
0!
0*
09
0>
0C
#752850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#752860000000
0!
0*
09
0>
0C
#752870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#752880000000
0!
0*
09
0>
0C
#752890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#752900000000
0!
0*
09
0>
0C
#752910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#752920000000
0!
0#
0*
0,
09
0>
0?
0C
#752930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#752940000000
0!
0*
09
0>
0C
#752950000000
1!
1*
19
1>
1C
#752960000000
0!
0*
09
0>
0C
#752970000000
1!
1*
19
1>
1C
#752980000000
0!
0*
09
0>
0C
#752990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#753000000000
0!
0*
09
0>
0C
#753010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#753020000000
0!
0*
09
0>
0C
#753030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#753040000000
0!
0*
09
0>
0C
#753050000000
1!
1*
b10 6
19
1>
1C
b10 G
#753060000000
0!
0*
09
0>
0C
#753070000000
1!
1*
b11 6
19
1>
1C
b11 G
#753080000000
0!
0*
09
0>
0C
#753090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#753100000000
0!
0*
09
0>
0C
#753110000000
1!
1*
b101 6
19
1>
1C
b101 G
#753120000000
0!
0*
09
0>
0C
#753130000000
1!
1*
b110 6
19
1>
1C
b110 G
#753140000000
0!
0*
09
0>
0C
#753150000000
1!
1*
b111 6
19
1>
1C
b111 G
#753160000000
0!
0*
09
0>
0C
#753170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#753180000000
0!
0*
09
0>
0C
#753190000000
1!
1*
b1 6
19
1>
1C
b1 G
#753200000000
0!
0*
09
0>
0C
#753210000000
1!
1*
b10 6
19
1>
1C
b10 G
#753220000000
0!
0*
09
0>
0C
#753230000000
1!
1*
b11 6
19
1>
1C
b11 G
#753240000000
0!
0*
09
0>
0C
#753250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#753260000000
0!
0*
09
0>
0C
#753270000000
1!
1*
b101 6
19
1>
1C
b101 G
#753280000000
0!
0*
09
0>
0C
#753290000000
1!
1*
b110 6
19
1>
1C
b110 G
#753300000000
0!
0*
09
0>
0C
#753310000000
1!
1*
b111 6
19
1>
1C
b111 G
#753320000000
0!
0*
09
0>
0C
#753330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#753340000000
0!
0*
09
0>
0C
#753350000000
1!
1*
b1 6
19
1>
1C
b1 G
#753360000000
0!
0*
09
0>
0C
#753370000000
1!
1*
b10 6
19
1>
1C
b10 G
#753380000000
0!
0*
09
0>
0C
#753390000000
1!
1*
b11 6
19
1>
1C
b11 G
#753400000000
0!
0*
09
0>
0C
#753410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#753420000000
0!
0*
09
0>
0C
#753430000000
1!
1*
b101 6
19
1>
1C
b101 G
#753440000000
0!
0*
09
0>
0C
#753450000000
1!
1*
b110 6
19
1>
1C
b110 G
#753460000000
0!
0*
09
0>
0C
#753470000000
1!
1*
b111 6
19
1>
1C
b111 G
#753480000000
0!
1"
0*
1+
09
1:
0>
0C
#753490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#753500000000
0!
0*
09
0>
0C
#753510000000
1!
1*
b1 6
19
1>
1C
b1 G
#753520000000
0!
0*
09
0>
0C
#753530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#753540000000
0!
0*
09
0>
0C
#753550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#753560000000
0!
0*
09
0>
0C
#753570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#753580000000
0!
0*
09
0>
0C
#753590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#753600000000
0!
0#
0*
0,
09
0>
0?
0C
#753610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#753620000000
0!
0*
09
0>
0C
#753630000000
1!
1*
19
1>
1C
#753640000000
0!
0*
09
0>
0C
#753650000000
1!
1*
19
1>
1C
#753660000000
0!
0*
09
0>
0C
#753670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#753680000000
0!
0*
09
0>
0C
#753690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#753700000000
0!
0*
09
0>
0C
#753710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#753720000000
0!
0*
09
0>
0C
#753730000000
1!
1*
b10 6
19
1>
1C
b10 G
#753740000000
0!
0*
09
0>
0C
#753750000000
1!
1*
b11 6
19
1>
1C
b11 G
#753760000000
0!
0*
09
0>
0C
#753770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#753780000000
0!
0*
09
0>
0C
#753790000000
1!
1*
b101 6
19
1>
1C
b101 G
#753800000000
0!
0*
09
0>
0C
#753810000000
1!
1*
b110 6
19
1>
1C
b110 G
#753820000000
0!
0*
09
0>
0C
#753830000000
1!
1*
b111 6
19
1>
1C
b111 G
#753840000000
0!
0*
09
0>
0C
#753850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#753860000000
0!
0*
09
0>
0C
#753870000000
1!
1*
b1 6
19
1>
1C
b1 G
#753880000000
0!
0*
09
0>
0C
#753890000000
1!
1*
b10 6
19
1>
1C
b10 G
#753900000000
0!
0*
09
0>
0C
#753910000000
1!
1*
b11 6
19
1>
1C
b11 G
#753920000000
0!
0*
09
0>
0C
#753930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#753940000000
0!
0*
09
0>
0C
#753950000000
1!
1*
b101 6
19
1>
1C
b101 G
#753960000000
0!
0*
09
0>
0C
#753970000000
1!
1*
b110 6
19
1>
1C
b110 G
#753980000000
0!
0*
09
0>
0C
#753990000000
1!
1*
b111 6
19
1>
1C
b111 G
#754000000000
0!
0*
09
0>
0C
#754010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#754020000000
0!
0*
09
0>
0C
#754030000000
1!
1*
b1 6
19
1>
1C
b1 G
#754040000000
0!
0*
09
0>
0C
#754050000000
1!
1*
b10 6
19
1>
1C
b10 G
#754060000000
0!
0*
09
0>
0C
#754070000000
1!
1*
b11 6
19
1>
1C
b11 G
#754080000000
0!
0*
09
0>
0C
#754090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#754100000000
0!
0*
09
0>
0C
#754110000000
1!
1*
b101 6
19
1>
1C
b101 G
#754120000000
0!
0*
09
0>
0C
#754130000000
1!
1*
b110 6
19
1>
1C
b110 G
#754140000000
0!
0*
09
0>
0C
#754150000000
1!
1*
b111 6
19
1>
1C
b111 G
#754160000000
0!
1"
0*
1+
09
1:
0>
0C
#754170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#754180000000
0!
0*
09
0>
0C
#754190000000
1!
1*
b1 6
19
1>
1C
b1 G
#754200000000
0!
0*
09
0>
0C
#754210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#754220000000
0!
0*
09
0>
0C
#754230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#754240000000
0!
0*
09
0>
0C
#754250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#754260000000
0!
0*
09
0>
0C
#754270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#754280000000
0!
0#
0*
0,
09
0>
0?
0C
#754290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#754300000000
0!
0*
09
0>
0C
#754310000000
1!
1*
19
1>
1C
#754320000000
0!
0*
09
0>
0C
#754330000000
1!
1*
19
1>
1C
#754340000000
0!
0*
09
0>
0C
#754350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#754360000000
0!
0*
09
0>
0C
#754370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#754380000000
0!
0*
09
0>
0C
#754390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#754400000000
0!
0*
09
0>
0C
#754410000000
1!
1*
b10 6
19
1>
1C
b10 G
#754420000000
0!
0*
09
0>
0C
#754430000000
1!
1*
b11 6
19
1>
1C
b11 G
#754440000000
0!
0*
09
0>
0C
#754450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#754460000000
0!
0*
09
0>
0C
#754470000000
1!
1*
b101 6
19
1>
1C
b101 G
#754480000000
0!
0*
09
0>
0C
#754490000000
1!
1*
b110 6
19
1>
1C
b110 G
#754500000000
0!
0*
09
0>
0C
#754510000000
1!
1*
b111 6
19
1>
1C
b111 G
#754520000000
0!
0*
09
0>
0C
#754530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#754540000000
0!
0*
09
0>
0C
#754550000000
1!
1*
b1 6
19
1>
1C
b1 G
#754560000000
0!
0*
09
0>
0C
#754570000000
1!
1*
b10 6
19
1>
1C
b10 G
#754580000000
0!
0*
09
0>
0C
#754590000000
1!
1*
b11 6
19
1>
1C
b11 G
#754600000000
0!
0*
09
0>
0C
#754610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#754620000000
0!
0*
09
0>
0C
#754630000000
1!
1*
b101 6
19
1>
1C
b101 G
#754640000000
0!
0*
09
0>
0C
#754650000000
1!
1*
b110 6
19
1>
1C
b110 G
#754660000000
0!
0*
09
0>
0C
#754670000000
1!
1*
b111 6
19
1>
1C
b111 G
#754680000000
0!
0*
09
0>
0C
#754690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#754700000000
0!
0*
09
0>
0C
#754710000000
1!
1*
b1 6
19
1>
1C
b1 G
#754720000000
0!
0*
09
0>
0C
#754730000000
1!
1*
b10 6
19
1>
1C
b10 G
#754740000000
0!
0*
09
0>
0C
#754750000000
1!
1*
b11 6
19
1>
1C
b11 G
#754760000000
0!
0*
09
0>
0C
#754770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#754780000000
0!
0*
09
0>
0C
#754790000000
1!
1*
b101 6
19
1>
1C
b101 G
#754800000000
0!
0*
09
0>
0C
#754810000000
1!
1*
b110 6
19
1>
1C
b110 G
#754820000000
0!
0*
09
0>
0C
#754830000000
1!
1*
b111 6
19
1>
1C
b111 G
#754840000000
0!
1"
0*
1+
09
1:
0>
0C
#754850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#754860000000
0!
0*
09
0>
0C
#754870000000
1!
1*
b1 6
19
1>
1C
b1 G
#754880000000
0!
0*
09
0>
0C
#754890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#754900000000
0!
0*
09
0>
0C
#754910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#754920000000
0!
0*
09
0>
0C
#754930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#754940000000
0!
0*
09
0>
0C
#754950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#754960000000
0!
0#
0*
0,
09
0>
0?
0C
#754970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#754980000000
0!
0*
09
0>
0C
#754990000000
1!
1*
19
1>
1C
#755000000000
0!
0*
09
0>
0C
#755010000000
1!
1*
19
1>
1C
#755020000000
0!
0*
09
0>
0C
#755030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#755040000000
0!
0*
09
0>
0C
#755050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#755060000000
0!
0*
09
0>
0C
#755070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#755080000000
0!
0*
09
0>
0C
#755090000000
1!
1*
b10 6
19
1>
1C
b10 G
#755100000000
0!
0*
09
0>
0C
#755110000000
1!
1*
b11 6
19
1>
1C
b11 G
#755120000000
0!
0*
09
0>
0C
#755130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#755140000000
0!
0*
09
0>
0C
#755150000000
1!
1*
b101 6
19
1>
1C
b101 G
#755160000000
0!
0*
09
0>
0C
#755170000000
1!
1*
b110 6
19
1>
1C
b110 G
#755180000000
0!
0*
09
0>
0C
#755190000000
1!
1*
b111 6
19
1>
1C
b111 G
#755200000000
0!
0*
09
0>
0C
#755210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#755220000000
0!
0*
09
0>
0C
#755230000000
1!
1*
b1 6
19
1>
1C
b1 G
#755240000000
0!
0*
09
0>
0C
#755250000000
1!
1*
b10 6
19
1>
1C
b10 G
#755260000000
0!
0*
09
0>
0C
#755270000000
1!
1*
b11 6
19
1>
1C
b11 G
#755280000000
0!
0*
09
0>
0C
#755290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#755300000000
0!
0*
09
0>
0C
#755310000000
1!
1*
b101 6
19
1>
1C
b101 G
#755320000000
0!
0*
09
0>
0C
#755330000000
1!
1*
b110 6
19
1>
1C
b110 G
#755340000000
0!
0*
09
0>
0C
#755350000000
1!
1*
b111 6
19
1>
1C
b111 G
#755360000000
0!
0*
09
0>
0C
#755370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#755380000000
0!
0*
09
0>
0C
#755390000000
1!
1*
b1 6
19
1>
1C
b1 G
#755400000000
0!
0*
09
0>
0C
#755410000000
1!
1*
b10 6
19
1>
1C
b10 G
#755420000000
0!
0*
09
0>
0C
#755430000000
1!
1*
b11 6
19
1>
1C
b11 G
#755440000000
0!
0*
09
0>
0C
#755450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#755460000000
0!
0*
09
0>
0C
#755470000000
1!
1*
b101 6
19
1>
1C
b101 G
#755480000000
0!
0*
09
0>
0C
#755490000000
1!
1*
b110 6
19
1>
1C
b110 G
#755500000000
0!
0*
09
0>
0C
#755510000000
1!
1*
b111 6
19
1>
1C
b111 G
#755520000000
0!
1"
0*
1+
09
1:
0>
0C
#755530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#755540000000
0!
0*
09
0>
0C
#755550000000
1!
1*
b1 6
19
1>
1C
b1 G
#755560000000
0!
0*
09
0>
0C
#755570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#755580000000
0!
0*
09
0>
0C
#755590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#755600000000
0!
0*
09
0>
0C
#755610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#755620000000
0!
0*
09
0>
0C
#755630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#755640000000
0!
0#
0*
0,
09
0>
0?
0C
#755650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#755660000000
0!
0*
09
0>
0C
#755670000000
1!
1*
19
1>
1C
#755680000000
0!
0*
09
0>
0C
#755690000000
1!
1*
19
1>
1C
#755700000000
0!
0*
09
0>
0C
#755710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#755720000000
0!
0*
09
0>
0C
#755730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#755740000000
0!
0*
09
0>
0C
#755750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#755760000000
0!
0*
09
0>
0C
#755770000000
1!
1*
b10 6
19
1>
1C
b10 G
#755780000000
0!
0*
09
0>
0C
#755790000000
1!
1*
b11 6
19
1>
1C
b11 G
#755800000000
0!
0*
09
0>
0C
#755810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#755820000000
0!
0*
09
0>
0C
#755830000000
1!
1*
b101 6
19
1>
1C
b101 G
#755840000000
0!
0*
09
0>
0C
#755850000000
1!
1*
b110 6
19
1>
1C
b110 G
#755860000000
0!
0*
09
0>
0C
#755870000000
1!
1*
b111 6
19
1>
1C
b111 G
#755880000000
0!
0*
09
0>
0C
#755890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#755900000000
0!
0*
09
0>
0C
#755910000000
1!
1*
b1 6
19
1>
1C
b1 G
#755920000000
0!
0*
09
0>
0C
#755930000000
1!
1*
b10 6
19
1>
1C
b10 G
#755940000000
0!
0*
09
0>
0C
#755950000000
1!
1*
b11 6
19
1>
1C
b11 G
#755960000000
0!
0*
09
0>
0C
#755970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#755980000000
0!
0*
09
0>
0C
#755990000000
1!
1*
b101 6
19
1>
1C
b101 G
#756000000000
0!
0*
09
0>
0C
#756010000000
1!
1*
b110 6
19
1>
1C
b110 G
#756020000000
0!
0*
09
0>
0C
#756030000000
1!
1*
b111 6
19
1>
1C
b111 G
#756040000000
0!
0*
09
0>
0C
#756050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#756060000000
0!
0*
09
0>
0C
#756070000000
1!
1*
b1 6
19
1>
1C
b1 G
#756080000000
0!
0*
09
0>
0C
#756090000000
1!
1*
b10 6
19
1>
1C
b10 G
#756100000000
0!
0*
09
0>
0C
#756110000000
1!
1*
b11 6
19
1>
1C
b11 G
#756120000000
0!
0*
09
0>
0C
#756130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#756140000000
0!
0*
09
0>
0C
#756150000000
1!
1*
b101 6
19
1>
1C
b101 G
#756160000000
0!
0*
09
0>
0C
#756170000000
1!
1*
b110 6
19
1>
1C
b110 G
#756180000000
0!
0*
09
0>
0C
#756190000000
1!
1*
b111 6
19
1>
1C
b111 G
#756200000000
0!
1"
0*
1+
09
1:
0>
0C
#756210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#756220000000
0!
0*
09
0>
0C
#756230000000
1!
1*
b1 6
19
1>
1C
b1 G
#756240000000
0!
0*
09
0>
0C
#756250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#756260000000
0!
0*
09
0>
0C
#756270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#756280000000
0!
0*
09
0>
0C
#756290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#756300000000
0!
0*
09
0>
0C
#756310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#756320000000
0!
0#
0*
0,
09
0>
0?
0C
#756330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#756340000000
0!
0*
09
0>
0C
#756350000000
1!
1*
19
1>
1C
#756360000000
0!
0*
09
0>
0C
#756370000000
1!
1*
19
1>
1C
#756380000000
0!
0*
09
0>
0C
#756390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#756400000000
0!
0*
09
0>
0C
#756410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#756420000000
0!
0*
09
0>
0C
#756430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#756440000000
0!
0*
09
0>
0C
#756450000000
1!
1*
b10 6
19
1>
1C
b10 G
#756460000000
0!
0*
09
0>
0C
#756470000000
1!
1*
b11 6
19
1>
1C
b11 G
#756480000000
0!
0*
09
0>
0C
#756490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#756500000000
0!
0*
09
0>
0C
#756510000000
1!
1*
b101 6
19
1>
1C
b101 G
#756520000000
0!
0*
09
0>
0C
#756530000000
1!
1*
b110 6
19
1>
1C
b110 G
#756540000000
0!
0*
09
0>
0C
#756550000000
1!
1*
b111 6
19
1>
1C
b111 G
#756560000000
0!
0*
09
0>
0C
#756570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#756580000000
0!
0*
09
0>
0C
#756590000000
1!
1*
b1 6
19
1>
1C
b1 G
#756600000000
0!
0*
09
0>
0C
#756610000000
1!
1*
b10 6
19
1>
1C
b10 G
#756620000000
0!
0*
09
0>
0C
#756630000000
1!
1*
b11 6
19
1>
1C
b11 G
#756640000000
0!
0*
09
0>
0C
#756650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#756660000000
0!
0*
09
0>
0C
#756670000000
1!
1*
b101 6
19
1>
1C
b101 G
#756680000000
0!
0*
09
0>
0C
#756690000000
1!
1*
b110 6
19
1>
1C
b110 G
#756700000000
0!
0*
09
0>
0C
#756710000000
1!
1*
b111 6
19
1>
1C
b111 G
#756720000000
0!
0*
09
0>
0C
#756730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#756740000000
0!
0*
09
0>
0C
#756750000000
1!
1*
b1 6
19
1>
1C
b1 G
#756760000000
0!
0*
09
0>
0C
#756770000000
1!
1*
b10 6
19
1>
1C
b10 G
#756780000000
0!
0*
09
0>
0C
#756790000000
1!
1*
b11 6
19
1>
1C
b11 G
#756800000000
0!
0*
09
0>
0C
#756810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#756820000000
0!
0*
09
0>
0C
#756830000000
1!
1*
b101 6
19
1>
1C
b101 G
#756840000000
0!
0*
09
0>
0C
#756850000000
1!
1*
b110 6
19
1>
1C
b110 G
#756860000000
0!
0*
09
0>
0C
#756870000000
1!
1*
b111 6
19
1>
1C
b111 G
#756880000000
0!
1"
0*
1+
09
1:
0>
0C
#756890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#756900000000
0!
0*
09
0>
0C
#756910000000
1!
1*
b1 6
19
1>
1C
b1 G
#756920000000
0!
0*
09
0>
0C
#756930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#756940000000
0!
0*
09
0>
0C
#756950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#756960000000
0!
0*
09
0>
0C
#756970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#756980000000
0!
0*
09
0>
0C
#756990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#757000000000
0!
0#
0*
0,
09
0>
0?
0C
#757010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#757020000000
0!
0*
09
0>
0C
#757030000000
1!
1*
19
1>
1C
#757040000000
0!
0*
09
0>
0C
#757050000000
1!
1*
19
1>
1C
#757060000000
0!
0*
09
0>
0C
#757070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#757080000000
0!
0*
09
0>
0C
#757090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#757100000000
0!
0*
09
0>
0C
#757110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#757120000000
0!
0*
09
0>
0C
#757130000000
1!
1*
b10 6
19
1>
1C
b10 G
#757140000000
0!
0*
09
0>
0C
#757150000000
1!
1*
b11 6
19
1>
1C
b11 G
#757160000000
0!
0*
09
0>
0C
#757170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#757180000000
0!
0*
09
0>
0C
#757190000000
1!
1*
b101 6
19
1>
1C
b101 G
#757200000000
0!
0*
09
0>
0C
#757210000000
1!
1*
b110 6
19
1>
1C
b110 G
#757220000000
0!
0*
09
0>
0C
#757230000000
1!
1*
b111 6
19
1>
1C
b111 G
#757240000000
0!
0*
09
0>
0C
#757250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#757260000000
0!
0*
09
0>
0C
#757270000000
1!
1*
b1 6
19
1>
1C
b1 G
#757280000000
0!
0*
09
0>
0C
#757290000000
1!
1*
b10 6
19
1>
1C
b10 G
#757300000000
0!
0*
09
0>
0C
#757310000000
1!
1*
b11 6
19
1>
1C
b11 G
#757320000000
0!
0*
09
0>
0C
#757330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#757340000000
0!
0*
09
0>
0C
#757350000000
1!
1*
b101 6
19
1>
1C
b101 G
#757360000000
0!
0*
09
0>
0C
#757370000000
1!
1*
b110 6
19
1>
1C
b110 G
#757380000000
0!
0*
09
0>
0C
#757390000000
1!
1*
b111 6
19
1>
1C
b111 G
#757400000000
0!
0*
09
0>
0C
#757410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#757420000000
0!
0*
09
0>
0C
#757430000000
1!
1*
b1 6
19
1>
1C
b1 G
#757440000000
0!
0*
09
0>
0C
#757450000000
1!
1*
b10 6
19
1>
1C
b10 G
#757460000000
0!
0*
09
0>
0C
#757470000000
1!
1*
b11 6
19
1>
1C
b11 G
#757480000000
0!
0*
09
0>
0C
#757490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#757500000000
0!
0*
09
0>
0C
#757510000000
1!
1*
b101 6
19
1>
1C
b101 G
#757520000000
0!
0*
09
0>
0C
#757530000000
1!
1*
b110 6
19
1>
1C
b110 G
#757540000000
0!
0*
09
0>
0C
#757550000000
1!
1*
b111 6
19
1>
1C
b111 G
#757560000000
0!
1"
0*
1+
09
1:
0>
0C
#757570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#757580000000
0!
0*
09
0>
0C
#757590000000
1!
1*
b1 6
19
1>
1C
b1 G
#757600000000
0!
0*
09
0>
0C
#757610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#757620000000
0!
0*
09
0>
0C
#757630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#757640000000
0!
0*
09
0>
0C
#757650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#757660000000
0!
0*
09
0>
0C
#757670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#757680000000
0!
0#
0*
0,
09
0>
0?
0C
#757690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#757700000000
0!
0*
09
0>
0C
#757710000000
1!
1*
19
1>
1C
#757720000000
0!
0*
09
0>
0C
#757730000000
1!
1*
19
1>
1C
#757740000000
0!
0*
09
0>
0C
#757750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#757760000000
0!
0*
09
0>
0C
#757770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#757780000000
0!
0*
09
0>
0C
#757790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#757800000000
0!
0*
09
0>
0C
#757810000000
1!
1*
b10 6
19
1>
1C
b10 G
#757820000000
0!
0*
09
0>
0C
#757830000000
1!
1*
b11 6
19
1>
1C
b11 G
#757840000000
0!
0*
09
0>
0C
#757850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#757860000000
0!
0*
09
0>
0C
#757870000000
1!
1*
b101 6
19
1>
1C
b101 G
#757880000000
0!
0*
09
0>
0C
#757890000000
1!
1*
b110 6
19
1>
1C
b110 G
#757900000000
0!
0*
09
0>
0C
#757910000000
1!
1*
b111 6
19
1>
1C
b111 G
#757920000000
0!
0*
09
0>
0C
#757930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#757940000000
0!
0*
09
0>
0C
#757950000000
1!
1*
b1 6
19
1>
1C
b1 G
#757960000000
0!
0*
09
0>
0C
#757970000000
1!
1*
b10 6
19
1>
1C
b10 G
#757980000000
0!
0*
09
0>
0C
#757990000000
1!
1*
b11 6
19
1>
1C
b11 G
#758000000000
0!
0*
09
0>
0C
#758010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#758020000000
0!
0*
09
0>
0C
#758030000000
1!
1*
b101 6
19
1>
1C
b101 G
#758040000000
0!
0*
09
0>
0C
#758050000000
1!
1*
b110 6
19
1>
1C
b110 G
#758060000000
0!
0*
09
0>
0C
#758070000000
1!
1*
b111 6
19
1>
1C
b111 G
#758080000000
0!
0*
09
0>
0C
#758090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#758100000000
0!
0*
09
0>
0C
#758110000000
1!
1*
b1 6
19
1>
1C
b1 G
#758120000000
0!
0*
09
0>
0C
#758130000000
1!
1*
b10 6
19
1>
1C
b10 G
#758140000000
0!
0*
09
0>
0C
#758150000000
1!
1*
b11 6
19
1>
1C
b11 G
#758160000000
0!
0*
09
0>
0C
#758170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#758180000000
0!
0*
09
0>
0C
#758190000000
1!
1*
b101 6
19
1>
1C
b101 G
#758200000000
0!
0*
09
0>
0C
#758210000000
1!
1*
b110 6
19
1>
1C
b110 G
#758220000000
0!
0*
09
0>
0C
#758230000000
1!
1*
b111 6
19
1>
1C
b111 G
#758240000000
0!
1"
0*
1+
09
1:
0>
0C
#758250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#758260000000
0!
0*
09
0>
0C
#758270000000
1!
1*
b1 6
19
1>
1C
b1 G
#758280000000
0!
0*
09
0>
0C
#758290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#758300000000
0!
0*
09
0>
0C
#758310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#758320000000
0!
0*
09
0>
0C
#758330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#758340000000
0!
0*
09
0>
0C
#758350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#758360000000
0!
0#
0*
0,
09
0>
0?
0C
#758370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#758380000000
0!
0*
09
0>
0C
#758390000000
1!
1*
19
1>
1C
#758400000000
0!
0*
09
0>
0C
#758410000000
1!
1*
19
1>
1C
#758420000000
0!
0*
09
0>
0C
#758430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#758440000000
0!
0*
09
0>
0C
#758450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#758460000000
0!
0*
09
0>
0C
#758470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#758480000000
0!
0*
09
0>
0C
#758490000000
1!
1*
b10 6
19
1>
1C
b10 G
#758500000000
0!
0*
09
0>
0C
#758510000000
1!
1*
b11 6
19
1>
1C
b11 G
#758520000000
0!
0*
09
0>
0C
#758530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#758540000000
0!
0*
09
0>
0C
#758550000000
1!
1*
b101 6
19
1>
1C
b101 G
#758560000000
0!
0*
09
0>
0C
#758570000000
1!
1*
b110 6
19
1>
1C
b110 G
#758580000000
0!
0*
09
0>
0C
#758590000000
1!
1*
b111 6
19
1>
1C
b111 G
#758600000000
0!
0*
09
0>
0C
#758610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#758620000000
0!
0*
09
0>
0C
#758630000000
1!
1*
b1 6
19
1>
1C
b1 G
#758640000000
0!
0*
09
0>
0C
#758650000000
1!
1*
b10 6
19
1>
1C
b10 G
#758660000000
0!
0*
09
0>
0C
#758670000000
1!
1*
b11 6
19
1>
1C
b11 G
#758680000000
0!
0*
09
0>
0C
#758690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#758700000000
0!
0*
09
0>
0C
#758710000000
1!
1*
b101 6
19
1>
1C
b101 G
#758720000000
0!
0*
09
0>
0C
#758730000000
1!
1*
b110 6
19
1>
1C
b110 G
#758740000000
0!
0*
09
0>
0C
#758750000000
1!
1*
b111 6
19
1>
1C
b111 G
#758760000000
0!
0*
09
0>
0C
#758770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#758780000000
0!
0*
09
0>
0C
#758790000000
1!
1*
b1 6
19
1>
1C
b1 G
#758800000000
0!
0*
09
0>
0C
#758810000000
1!
1*
b10 6
19
1>
1C
b10 G
#758820000000
0!
0*
09
0>
0C
#758830000000
1!
1*
b11 6
19
1>
1C
b11 G
#758840000000
0!
0*
09
0>
0C
#758850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#758860000000
0!
0*
09
0>
0C
#758870000000
1!
1*
b101 6
19
1>
1C
b101 G
#758880000000
0!
0*
09
0>
0C
#758890000000
1!
1*
b110 6
19
1>
1C
b110 G
#758900000000
0!
0*
09
0>
0C
#758910000000
1!
1*
b111 6
19
1>
1C
b111 G
#758920000000
0!
1"
0*
1+
09
1:
0>
0C
#758930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#758940000000
0!
0*
09
0>
0C
#758950000000
1!
1*
b1 6
19
1>
1C
b1 G
#758960000000
0!
0*
09
0>
0C
#758970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#758980000000
0!
0*
09
0>
0C
#758990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#759000000000
0!
0*
09
0>
0C
#759010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#759020000000
0!
0*
09
0>
0C
#759030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#759040000000
0!
0#
0*
0,
09
0>
0?
0C
#759050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#759060000000
0!
0*
09
0>
0C
#759070000000
1!
1*
19
1>
1C
#759080000000
0!
0*
09
0>
0C
#759090000000
1!
1*
19
1>
1C
#759100000000
0!
0*
09
0>
0C
#759110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#759120000000
0!
0*
09
0>
0C
#759130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#759140000000
0!
0*
09
0>
0C
#759150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#759160000000
0!
0*
09
0>
0C
#759170000000
1!
1*
b10 6
19
1>
1C
b10 G
#759180000000
0!
0*
09
0>
0C
#759190000000
1!
1*
b11 6
19
1>
1C
b11 G
#759200000000
0!
0*
09
0>
0C
#759210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#759220000000
0!
0*
09
0>
0C
#759230000000
1!
1*
b101 6
19
1>
1C
b101 G
#759240000000
0!
0*
09
0>
0C
#759250000000
1!
1*
b110 6
19
1>
1C
b110 G
#759260000000
0!
0*
09
0>
0C
#759270000000
1!
1*
b111 6
19
1>
1C
b111 G
#759280000000
0!
0*
09
0>
0C
#759290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#759300000000
0!
0*
09
0>
0C
#759310000000
1!
1*
b1 6
19
1>
1C
b1 G
#759320000000
0!
0*
09
0>
0C
#759330000000
1!
1*
b10 6
19
1>
1C
b10 G
#759340000000
0!
0*
09
0>
0C
#759350000000
1!
1*
b11 6
19
1>
1C
b11 G
#759360000000
0!
0*
09
0>
0C
#759370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#759380000000
0!
0*
09
0>
0C
#759390000000
1!
1*
b101 6
19
1>
1C
b101 G
#759400000000
0!
0*
09
0>
0C
#759410000000
1!
1*
b110 6
19
1>
1C
b110 G
#759420000000
0!
0*
09
0>
0C
#759430000000
1!
1*
b111 6
19
1>
1C
b111 G
#759440000000
0!
0*
09
0>
0C
#759450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#759460000000
0!
0*
09
0>
0C
#759470000000
1!
1*
b1 6
19
1>
1C
b1 G
#759480000000
0!
0*
09
0>
0C
#759490000000
1!
1*
b10 6
19
1>
1C
b10 G
#759500000000
0!
0*
09
0>
0C
#759510000000
1!
1*
b11 6
19
1>
1C
b11 G
#759520000000
0!
0*
09
0>
0C
#759530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#759540000000
0!
0*
09
0>
0C
#759550000000
1!
1*
b101 6
19
1>
1C
b101 G
#759560000000
0!
0*
09
0>
0C
#759570000000
1!
1*
b110 6
19
1>
1C
b110 G
#759580000000
0!
0*
09
0>
0C
#759590000000
1!
1*
b111 6
19
1>
1C
b111 G
#759600000000
0!
1"
0*
1+
09
1:
0>
0C
#759610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#759620000000
0!
0*
09
0>
0C
#759630000000
1!
1*
b1 6
19
1>
1C
b1 G
#759640000000
0!
0*
09
0>
0C
#759650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#759660000000
0!
0*
09
0>
0C
#759670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#759680000000
0!
0*
09
0>
0C
#759690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#759700000000
0!
0*
09
0>
0C
#759710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#759720000000
0!
0#
0*
0,
09
0>
0?
0C
#759730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#759740000000
0!
0*
09
0>
0C
#759750000000
1!
1*
19
1>
1C
#759760000000
0!
0*
09
0>
0C
#759770000000
1!
1*
19
1>
1C
#759780000000
0!
0*
09
0>
0C
#759790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#759800000000
0!
0*
09
0>
0C
#759810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#759820000000
0!
0*
09
0>
0C
#759830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#759840000000
0!
0*
09
0>
0C
#759850000000
1!
1*
b10 6
19
1>
1C
b10 G
#759860000000
0!
0*
09
0>
0C
#759870000000
1!
1*
b11 6
19
1>
1C
b11 G
#759880000000
0!
0*
09
0>
0C
#759890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#759900000000
0!
0*
09
0>
0C
#759910000000
1!
1*
b101 6
19
1>
1C
b101 G
#759920000000
0!
0*
09
0>
0C
#759930000000
1!
1*
b110 6
19
1>
1C
b110 G
#759940000000
0!
0*
09
0>
0C
#759950000000
1!
1*
b111 6
19
1>
1C
b111 G
#759960000000
0!
0*
09
0>
0C
#759970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#759980000000
0!
0*
09
0>
0C
#759990000000
1!
1*
b1 6
19
1>
1C
b1 G
#760000000000
0!
0*
09
0>
0C
#760010000000
1!
1*
b10 6
19
1>
1C
b10 G
#760020000000
0!
0*
09
0>
0C
#760030000000
1!
1*
b11 6
19
1>
1C
b11 G
#760040000000
0!
0*
09
0>
0C
#760050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#760060000000
0!
0*
09
0>
0C
#760070000000
1!
1*
b101 6
19
1>
1C
b101 G
#760080000000
0!
0*
09
0>
0C
#760090000000
1!
1*
b110 6
19
1>
1C
b110 G
#760100000000
0!
0*
09
0>
0C
#760110000000
1!
1*
b111 6
19
1>
1C
b111 G
#760120000000
0!
0*
09
0>
0C
#760130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#760140000000
0!
0*
09
0>
0C
#760150000000
1!
1*
b1 6
19
1>
1C
b1 G
#760160000000
0!
0*
09
0>
0C
#760170000000
1!
1*
b10 6
19
1>
1C
b10 G
#760180000000
0!
0*
09
0>
0C
#760190000000
1!
1*
b11 6
19
1>
1C
b11 G
#760200000000
0!
0*
09
0>
0C
#760210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#760220000000
0!
0*
09
0>
0C
#760230000000
1!
1*
b101 6
19
1>
1C
b101 G
#760240000000
0!
0*
09
0>
0C
#760250000000
1!
1*
b110 6
19
1>
1C
b110 G
#760260000000
0!
0*
09
0>
0C
#760270000000
1!
1*
b111 6
19
1>
1C
b111 G
#760280000000
0!
1"
0*
1+
09
1:
0>
0C
#760290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#760300000000
0!
0*
09
0>
0C
#760310000000
1!
1*
b1 6
19
1>
1C
b1 G
#760320000000
0!
0*
09
0>
0C
#760330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#760340000000
0!
0*
09
0>
0C
#760350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#760360000000
0!
0*
09
0>
0C
#760370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#760380000000
0!
0*
09
0>
0C
#760390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#760400000000
0!
0#
0*
0,
09
0>
0?
0C
#760410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#760420000000
0!
0*
09
0>
0C
#760430000000
1!
1*
19
1>
1C
#760440000000
0!
0*
09
0>
0C
#760450000000
1!
1*
19
1>
1C
#760460000000
0!
0*
09
0>
0C
#760470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#760480000000
0!
0*
09
0>
0C
#760490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#760500000000
0!
0*
09
0>
0C
#760510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#760520000000
0!
0*
09
0>
0C
#760530000000
1!
1*
b10 6
19
1>
1C
b10 G
#760540000000
0!
0*
09
0>
0C
#760550000000
1!
1*
b11 6
19
1>
1C
b11 G
#760560000000
0!
0*
09
0>
0C
#760570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#760580000000
0!
0*
09
0>
0C
#760590000000
1!
1*
b101 6
19
1>
1C
b101 G
#760600000000
0!
0*
09
0>
0C
#760610000000
1!
1*
b110 6
19
1>
1C
b110 G
#760620000000
0!
0*
09
0>
0C
#760630000000
1!
1*
b111 6
19
1>
1C
b111 G
#760640000000
0!
0*
09
0>
0C
#760650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#760660000000
0!
0*
09
0>
0C
#760670000000
1!
1*
b1 6
19
1>
1C
b1 G
#760680000000
0!
0*
09
0>
0C
#760690000000
1!
1*
b10 6
19
1>
1C
b10 G
#760700000000
0!
0*
09
0>
0C
#760710000000
1!
1*
b11 6
19
1>
1C
b11 G
#760720000000
0!
0*
09
0>
0C
#760730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#760740000000
0!
0*
09
0>
0C
#760750000000
1!
1*
b101 6
19
1>
1C
b101 G
#760760000000
0!
0*
09
0>
0C
#760770000000
1!
1*
b110 6
19
1>
1C
b110 G
#760780000000
0!
0*
09
0>
0C
#760790000000
1!
1*
b111 6
19
1>
1C
b111 G
#760800000000
0!
0*
09
0>
0C
#760810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#760820000000
0!
0*
09
0>
0C
#760830000000
1!
1*
b1 6
19
1>
1C
b1 G
#760840000000
0!
0*
09
0>
0C
#760850000000
1!
1*
b10 6
19
1>
1C
b10 G
#760860000000
0!
0*
09
0>
0C
#760870000000
1!
1*
b11 6
19
1>
1C
b11 G
#760880000000
0!
0*
09
0>
0C
#760890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#760900000000
0!
0*
09
0>
0C
#760910000000
1!
1*
b101 6
19
1>
1C
b101 G
#760920000000
0!
0*
09
0>
0C
#760930000000
1!
1*
b110 6
19
1>
1C
b110 G
#760940000000
0!
0*
09
0>
0C
#760950000000
1!
1*
b111 6
19
1>
1C
b111 G
#760960000000
0!
1"
0*
1+
09
1:
0>
0C
#760970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#760980000000
0!
0*
09
0>
0C
#760990000000
1!
1*
b1 6
19
1>
1C
b1 G
#761000000000
0!
0*
09
0>
0C
#761010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#761020000000
0!
0*
09
0>
0C
#761030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#761040000000
0!
0*
09
0>
0C
#761050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#761060000000
0!
0*
09
0>
0C
#761070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#761080000000
0!
0#
0*
0,
09
0>
0?
0C
#761090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#761100000000
0!
0*
09
0>
0C
#761110000000
1!
1*
19
1>
1C
#761120000000
0!
0*
09
0>
0C
#761130000000
1!
1*
19
1>
1C
#761140000000
0!
0*
09
0>
0C
#761150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#761160000000
0!
0*
09
0>
0C
#761170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#761180000000
0!
0*
09
0>
0C
#761190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#761200000000
0!
0*
09
0>
0C
#761210000000
1!
1*
b10 6
19
1>
1C
b10 G
#761220000000
0!
0*
09
0>
0C
#761230000000
1!
1*
b11 6
19
1>
1C
b11 G
#761240000000
0!
0*
09
0>
0C
#761250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#761260000000
0!
0*
09
0>
0C
#761270000000
1!
1*
b101 6
19
1>
1C
b101 G
#761280000000
0!
0*
09
0>
0C
#761290000000
1!
1*
b110 6
19
1>
1C
b110 G
#761300000000
0!
0*
09
0>
0C
#761310000000
1!
1*
b111 6
19
1>
1C
b111 G
#761320000000
0!
0*
09
0>
0C
#761330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#761340000000
0!
0*
09
0>
0C
#761350000000
1!
1*
b1 6
19
1>
1C
b1 G
#761360000000
0!
0*
09
0>
0C
#761370000000
1!
1*
b10 6
19
1>
1C
b10 G
#761380000000
0!
0*
09
0>
0C
#761390000000
1!
1*
b11 6
19
1>
1C
b11 G
#761400000000
0!
0*
09
0>
0C
#761410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#761420000000
0!
0*
09
0>
0C
#761430000000
1!
1*
b101 6
19
1>
1C
b101 G
#761440000000
0!
0*
09
0>
0C
#761450000000
1!
1*
b110 6
19
1>
1C
b110 G
#761460000000
0!
0*
09
0>
0C
#761470000000
1!
1*
b111 6
19
1>
1C
b111 G
#761480000000
0!
0*
09
0>
0C
#761490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#761500000000
0!
0*
09
0>
0C
#761510000000
1!
1*
b1 6
19
1>
1C
b1 G
#761520000000
0!
0*
09
0>
0C
#761530000000
1!
1*
b10 6
19
1>
1C
b10 G
#761540000000
0!
0*
09
0>
0C
#761550000000
1!
1*
b11 6
19
1>
1C
b11 G
#761560000000
0!
0*
09
0>
0C
#761570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#761580000000
0!
0*
09
0>
0C
#761590000000
1!
1*
b101 6
19
1>
1C
b101 G
#761600000000
0!
0*
09
0>
0C
#761610000000
1!
1*
b110 6
19
1>
1C
b110 G
#761620000000
0!
0*
09
0>
0C
#761630000000
1!
1*
b111 6
19
1>
1C
b111 G
#761640000000
0!
1"
0*
1+
09
1:
0>
0C
#761650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#761660000000
0!
0*
09
0>
0C
#761670000000
1!
1*
b1 6
19
1>
1C
b1 G
#761680000000
0!
0*
09
0>
0C
#761690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#761700000000
0!
0*
09
0>
0C
#761710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#761720000000
0!
0*
09
0>
0C
#761730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#761740000000
0!
0*
09
0>
0C
#761750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#761760000000
0!
0#
0*
0,
09
0>
0?
0C
#761770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#761780000000
0!
0*
09
0>
0C
#761790000000
1!
1*
19
1>
1C
#761800000000
0!
0*
09
0>
0C
#761810000000
1!
1*
19
1>
1C
#761820000000
0!
0*
09
0>
0C
#761830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#761840000000
0!
0*
09
0>
0C
#761850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#761860000000
0!
0*
09
0>
0C
#761870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#761880000000
0!
0*
09
0>
0C
#761890000000
1!
1*
b10 6
19
1>
1C
b10 G
#761900000000
0!
0*
09
0>
0C
#761910000000
1!
1*
b11 6
19
1>
1C
b11 G
#761920000000
0!
0*
09
0>
0C
#761930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#761940000000
0!
0*
09
0>
0C
#761950000000
1!
1*
b101 6
19
1>
1C
b101 G
#761960000000
0!
0*
09
0>
0C
#761970000000
1!
1*
b110 6
19
1>
1C
b110 G
#761980000000
0!
0*
09
0>
0C
#761990000000
1!
1*
b111 6
19
1>
1C
b111 G
#762000000000
0!
0*
09
0>
0C
#762010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#762020000000
0!
0*
09
0>
0C
#762030000000
1!
1*
b1 6
19
1>
1C
b1 G
#762040000000
0!
0*
09
0>
0C
#762050000000
1!
1*
b10 6
19
1>
1C
b10 G
#762060000000
0!
0*
09
0>
0C
#762070000000
1!
1*
b11 6
19
1>
1C
b11 G
#762080000000
0!
0*
09
0>
0C
#762090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#762100000000
0!
0*
09
0>
0C
#762110000000
1!
1*
b101 6
19
1>
1C
b101 G
#762120000000
0!
0*
09
0>
0C
#762130000000
1!
1*
b110 6
19
1>
1C
b110 G
#762140000000
0!
0*
09
0>
0C
#762150000000
1!
1*
b111 6
19
1>
1C
b111 G
#762160000000
0!
0*
09
0>
0C
#762170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#762180000000
0!
0*
09
0>
0C
#762190000000
1!
1*
b1 6
19
1>
1C
b1 G
#762200000000
0!
0*
09
0>
0C
#762210000000
1!
1*
b10 6
19
1>
1C
b10 G
#762220000000
0!
0*
09
0>
0C
#762230000000
1!
1*
b11 6
19
1>
1C
b11 G
#762240000000
0!
0*
09
0>
0C
#762250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#762260000000
0!
0*
09
0>
0C
#762270000000
1!
1*
b101 6
19
1>
1C
b101 G
#762280000000
0!
0*
09
0>
0C
#762290000000
1!
1*
b110 6
19
1>
1C
b110 G
#762300000000
0!
0*
09
0>
0C
#762310000000
1!
1*
b111 6
19
1>
1C
b111 G
#762320000000
0!
1"
0*
1+
09
1:
0>
0C
#762330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#762340000000
0!
0*
09
0>
0C
#762350000000
1!
1*
b1 6
19
1>
1C
b1 G
#762360000000
0!
0*
09
0>
0C
#762370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#762380000000
0!
0*
09
0>
0C
#762390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#762400000000
0!
0*
09
0>
0C
#762410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#762420000000
0!
0*
09
0>
0C
#762430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#762440000000
0!
0#
0*
0,
09
0>
0?
0C
#762450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#762460000000
0!
0*
09
0>
0C
#762470000000
1!
1*
19
1>
1C
#762480000000
0!
0*
09
0>
0C
#762490000000
1!
1*
19
1>
1C
#762500000000
0!
0*
09
0>
0C
#762510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#762520000000
0!
0*
09
0>
0C
#762530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#762540000000
0!
0*
09
0>
0C
#762550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#762560000000
0!
0*
09
0>
0C
#762570000000
1!
1*
b10 6
19
1>
1C
b10 G
#762580000000
0!
0*
09
0>
0C
#762590000000
1!
1*
b11 6
19
1>
1C
b11 G
#762600000000
0!
0*
09
0>
0C
#762610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#762620000000
0!
0*
09
0>
0C
#762630000000
1!
1*
b101 6
19
1>
1C
b101 G
#762640000000
0!
0*
09
0>
0C
#762650000000
1!
1*
b110 6
19
1>
1C
b110 G
#762660000000
0!
0*
09
0>
0C
#762670000000
1!
1*
b111 6
19
1>
1C
b111 G
#762680000000
0!
0*
09
0>
0C
#762690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#762700000000
0!
0*
09
0>
0C
#762710000000
1!
1*
b1 6
19
1>
1C
b1 G
#762720000000
0!
0*
09
0>
0C
#762730000000
1!
1*
b10 6
19
1>
1C
b10 G
#762740000000
0!
0*
09
0>
0C
#762750000000
1!
1*
b11 6
19
1>
1C
b11 G
#762760000000
0!
0*
09
0>
0C
#762770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#762780000000
0!
0*
09
0>
0C
#762790000000
1!
1*
b101 6
19
1>
1C
b101 G
#762800000000
0!
0*
09
0>
0C
#762810000000
1!
1*
b110 6
19
1>
1C
b110 G
#762820000000
0!
0*
09
0>
0C
#762830000000
1!
1*
b111 6
19
1>
1C
b111 G
#762840000000
0!
0*
09
0>
0C
#762850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#762860000000
0!
0*
09
0>
0C
#762870000000
1!
1*
b1 6
19
1>
1C
b1 G
#762880000000
0!
0*
09
0>
0C
#762890000000
1!
1*
b10 6
19
1>
1C
b10 G
#762900000000
0!
0*
09
0>
0C
#762910000000
1!
1*
b11 6
19
1>
1C
b11 G
#762920000000
0!
0*
09
0>
0C
#762930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#762940000000
0!
0*
09
0>
0C
#762950000000
1!
1*
b101 6
19
1>
1C
b101 G
#762960000000
0!
0*
09
0>
0C
#762970000000
1!
1*
b110 6
19
1>
1C
b110 G
#762980000000
0!
0*
09
0>
0C
#762990000000
1!
1*
b111 6
19
1>
1C
b111 G
#763000000000
0!
1"
0*
1+
09
1:
0>
0C
#763010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#763020000000
0!
0*
09
0>
0C
#763030000000
1!
1*
b1 6
19
1>
1C
b1 G
#763040000000
0!
0*
09
0>
0C
#763050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#763060000000
0!
0*
09
0>
0C
#763070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#763080000000
0!
0*
09
0>
0C
#763090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#763100000000
0!
0*
09
0>
0C
#763110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#763120000000
0!
0#
0*
0,
09
0>
0?
0C
#763130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#763140000000
0!
0*
09
0>
0C
#763150000000
1!
1*
19
1>
1C
#763160000000
0!
0*
09
0>
0C
#763170000000
1!
1*
19
1>
1C
#763180000000
0!
0*
09
0>
0C
#763190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#763200000000
0!
0*
09
0>
0C
#763210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#763220000000
0!
0*
09
0>
0C
#763230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#763240000000
0!
0*
09
0>
0C
#763250000000
1!
1*
b10 6
19
1>
1C
b10 G
#763260000000
0!
0*
09
0>
0C
#763270000000
1!
1*
b11 6
19
1>
1C
b11 G
#763280000000
0!
0*
09
0>
0C
#763290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#763300000000
0!
0*
09
0>
0C
#763310000000
1!
1*
b101 6
19
1>
1C
b101 G
#763320000000
0!
0*
09
0>
0C
#763330000000
1!
1*
b110 6
19
1>
1C
b110 G
#763340000000
0!
0*
09
0>
0C
#763350000000
1!
1*
b111 6
19
1>
1C
b111 G
#763360000000
0!
0*
09
0>
0C
#763370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#763380000000
0!
0*
09
0>
0C
#763390000000
1!
1*
b1 6
19
1>
1C
b1 G
#763400000000
0!
0*
09
0>
0C
#763410000000
1!
1*
b10 6
19
1>
1C
b10 G
#763420000000
0!
0*
09
0>
0C
#763430000000
1!
1*
b11 6
19
1>
1C
b11 G
#763440000000
0!
0*
09
0>
0C
#763450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#763460000000
0!
0*
09
0>
0C
#763470000000
1!
1*
b101 6
19
1>
1C
b101 G
#763480000000
0!
0*
09
0>
0C
#763490000000
1!
1*
b110 6
19
1>
1C
b110 G
#763500000000
0!
0*
09
0>
0C
#763510000000
1!
1*
b111 6
19
1>
1C
b111 G
#763520000000
0!
0*
09
0>
0C
#763530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#763540000000
0!
0*
09
0>
0C
#763550000000
1!
1*
b1 6
19
1>
1C
b1 G
#763560000000
0!
0*
09
0>
0C
#763570000000
1!
1*
b10 6
19
1>
1C
b10 G
#763580000000
0!
0*
09
0>
0C
#763590000000
1!
1*
b11 6
19
1>
1C
b11 G
#763600000000
0!
0*
09
0>
0C
#763610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#763620000000
0!
0*
09
0>
0C
#763630000000
1!
1*
b101 6
19
1>
1C
b101 G
#763640000000
0!
0*
09
0>
0C
#763650000000
1!
1*
b110 6
19
1>
1C
b110 G
#763660000000
0!
0*
09
0>
0C
#763670000000
1!
1*
b111 6
19
1>
1C
b111 G
#763680000000
0!
1"
0*
1+
09
1:
0>
0C
#763690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#763700000000
0!
0*
09
0>
0C
#763710000000
1!
1*
b1 6
19
1>
1C
b1 G
#763720000000
0!
0*
09
0>
0C
#763730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#763740000000
0!
0*
09
0>
0C
#763750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#763760000000
0!
0*
09
0>
0C
#763770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#763780000000
0!
0*
09
0>
0C
#763790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#763800000000
0!
0#
0*
0,
09
0>
0?
0C
#763810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#763820000000
0!
0*
09
0>
0C
#763830000000
1!
1*
19
1>
1C
#763840000000
0!
0*
09
0>
0C
#763850000000
1!
1*
19
1>
1C
#763860000000
0!
0*
09
0>
0C
#763870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#763880000000
0!
0*
09
0>
0C
#763890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#763900000000
0!
0*
09
0>
0C
#763910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#763920000000
0!
0*
09
0>
0C
#763930000000
1!
1*
b10 6
19
1>
1C
b10 G
#763940000000
0!
0*
09
0>
0C
#763950000000
1!
1*
b11 6
19
1>
1C
b11 G
#763960000000
0!
0*
09
0>
0C
#763970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#763980000000
0!
0*
09
0>
0C
#763990000000
1!
1*
b101 6
19
1>
1C
b101 G
#764000000000
0!
0*
09
0>
0C
#764010000000
1!
1*
b110 6
19
1>
1C
b110 G
#764020000000
0!
0*
09
0>
0C
#764030000000
1!
1*
b111 6
19
1>
1C
b111 G
#764040000000
0!
0*
09
0>
0C
#764050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#764060000000
0!
0*
09
0>
0C
#764070000000
1!
1*
b1 6
19
1>
1C
b1 G
#764080000000
0!
0*
09
0>
0C
#764090000000
1!
1*
b10 6
19
1>
1C
b10 G
#764100000000
0!
0*
09
0>
0C
#764110000000
1!
1*
b11 6
19
1>
1C
b11 G
#764120000000
0!
0*
09
0>
0C
#764130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#764140000000
0!
0*
09
0>
0C
#764150000000
1!
1*
b101 6
19
1>
1C
b101 G
#764160000000
0!
0*
09
0>
0C
#764170000000
1!
1*
b110 6
19
1>
1C
b110 G
#764180000000
0!
0*
09
0>
0C
#764190000000
1!
1*
b111 6
19
1>
1C
b111 G
#764200000000
0!
0*
09
0>
0C
#764210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#764220000000
0!
0*
09
0>
0C
#764230000000
1!
1*
b1 6
19
1>
1C
b1 G
#764240000000
0!
0*
09
0>
0C
#764250000000
1!
1*
b10 6
19
1>
1C
b10 G
#764260000000
0!
0*
09
0>
0C
#764270000000
1!
1*
b11 6
19
1>
1C
b11 G
#764280000000
0!
0*
09
0>
0C
#764290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#764300000000
0!
0*
09
0>
0C
#764310000000
1!
1*
b101 6
19
1>
1C
b101 G
#764320000000
0!
0*
09
0>
0C
#764330000000
1!
1*
b110 6
19
1>
1C
b110 G
#764340000000
0!
0*
09
0>
0C
#764350000000
1!
1*
b111 6
19
1>
1C
b111 G
#764360000000
0!
1"
0*
1+
09
1:
0>
0C
#764370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#764380000000
0!
0*
09
0>
0C
#764390000000
1!
1*
b1 6
19
1>
1C
b1 G
#764400000000
0!
0*
09
0>
0C
#764410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#764420000000
0!
0*
09
0>
0C
#764430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#764440000000
0!
0*
09
0>
0C
#764450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#764460000000
0!
0*
09
0>
0C
#764470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#764480000000
0!
0#
0*
0,
09
0>
0?
0C
#764490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#764500000000
0!
0*
09
0>
0C
#764510000000
1!
1*
19
1>
1C
#764520000000
0!
0*
09
0>
0C
#764530000000
1!
1*
19
1>
1C
#764540000000
0!
0*
09
0>
0C
#764550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#764560000000
0!
0*
09
0>
0C
#764570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#764580000000
0!
0*
09
0>
0C
#764590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#764600000000
0!
0*
09
0>
0C
#764610000000
1!
1*
b10 6
19
1>
1C
b10 G
#764620000000
0!
0*
09
0>
0C
#764630000000
1!
1*
b11 6
19
1>
1C
b11 G
#764640000000
0!
0*
09
0>
0C
#764650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#764660000000
0!
0*
09
0>
0C
#764670000000
1!
1*
b101 6
19
1>
1C
b101 G
#764680000000
0!
0*
09
0>
0C
#764690000000
1!
1*
b110 6
19
1>
1C
b110 G
#764700000000
0!
0*
09
0>
0C
#764710000000
1!
1*
b111 6
19
1>
1C
b111 G
#764720000000
0!
0*
09
0>
0C
#764730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#764740000000
0!
0*
09
0>
0C
#764750000000
1!
1*
b1 6
19
1>
1C
b1 G
#764760000000
0!
0*
09
0>
0C
#764770000000
1!
1*
b10 6
19
1>
1C
b10 G
#764780000000
0!
0*
09
0>
0C
#764790000000
1!
1*
b11 6
19
1>
1C
b11 G
#764800000000
0!
0*
09
0>
0C
#764810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#764820000000
0!
0*
09
0>
0C
#764830000000
1!
1*
b101 6
19
1>
1C
b101 G
#764840000000
0!
0*
09
0>
0C
#764850000000
1!
1*
b110 6
19
1>
1C
b110 G
#764860000000
0!
0*
09
0>
0C
#764870000000
1!
1*
b111 6
19
1>
1C
b111 G
#764880000000
0!
0*
09
0>
0C
#764890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#764900000000
0!
0*
09
0>
0C
#764910000000
1!
1*
b1 6
19
1>
1C
b1 G
#764920000000
0!
0*
09
0>
0C
#764930000000
1!
1*
b10 6
19
1>
1C
b10 G
#764940000000
0!
0*
09
0>
0C
#764950000000
1!
1*
b11 6
19
1>
1C
b11 G
#764960000000
0!
0*
09
0>
0C
#764970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#764980000000
0!
0*
09
0>
0C
#764990000000
1!
1*
b101 6
19
1>
1C
b101 G
#765000000000
0!
0*
09
0>
0C
#765010000000
1!
1*
b110 6
19
1>
1C
b110 G
#765020000000
0!
0*
09
0>
0C
#765030000000
1!
1*
b111 6
19
1>
1C
b111 G
#765040000000
0!
1"
0*
1+
09
1:
0>
0C
#765050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#765060000000
0!
0*
09
0>
0C
#765070000000
1!
1*
b1 6
19
1>
1C
b1 G
#765080000000
0!
0*
09
0>
0C
#765090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#765100000000
0!
0*
09
0>
0C
#765110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#765120000000
0!
0*
09
0>
0C
#765130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#765140000000
0!
0*
09
0>
0C
#765150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#765160000000
0!
0#
0*
0,
09
0>
0?
0C
#765170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#765180000000
0!
0*
09
0>
0C
#765190000000
1!
1*
19
1>
1C
#765200000000
0!
0*
09
0>
0C
#765210000000
1!
1*
19
1>
1C
#765220000000
0!
0*
09
0>
0C
#765230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#765240000000
0!
0*
09
0>
0C
#765250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#765260000000
0!
0*
09
0>
0C
#765270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#765280000000
0!
0*
09
0>
0C
#765290000000
1!
1*
b10 6
19
1>
1C
b10 G
#765300000000
0!
0*
09
0>
0C
#765310000000
1!
1*
b11 6
19
1>
1C
b11 G
#765320000000
0!
0*
09
0>
0C
#765330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#765340000000
0!
0*
09
0>
0C
#765350000000
1!
1*
b101 6
19
1>
1C
b101 G
#765360000000
0!
0*
09
0>
0C
#765370000000
1!
1*
b110 6
19
1>
1C
b110 G
#765380000000
0!
0*
09
0>
0C
#765390000000
1!
1*
b111 6
19
1>
1C
b111 G
#765400000000
0!
0*
09
0>
0C
#765410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#765420000000
0!
0*
09
0>
0C
#765430000000
1!
1*
b1 6
19
1>
1C
b1 G
#765440000000
0!
0*
09
0>
0C
#765450000000
1!
1*
b10 6
19
1>
1C
b10 G
#765460000000
0!
0*
09
0>
0C
#765470000000
1!
1*
b11 6
19
1>
1C
b11 G
#765480000000
0!
0*
09
0>
0C
#765490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#765500000000
0!
0*
09
0>
0C
#765510000000
1!
1*
b101 6
19
1>
1C
b101 G
#765520000000
0!
0*
09
0>
0C
#765530000000
1!
1*
b110 6
19
1>
1C
b110 G
#765540000000
0!
0*
09
0>
0C
#765550000000
1!
1*
b111 6
19
1>
1C
b111 G
#765560000000
0!
0*
09
0>
0C
#765570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#765580000000
0!
0*
09
0>
0C
#765590000000
1!
1*
b1 6
19
1>
1C
b1 G
#765600000000
0!
0*
09
0>
0C
#765610000000
1!
1*
b10 6
19
1>
1C
b10 G
#765620000000
0!
0*
09
0>
0C
#765630000000
1!
1*
b11 6
19
1>
1C
b11 G
#765640000000
0!
0*
09
0>
0C
#765650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#765660000000
0!
0*
09
0>
0C
#765670000000
1!
1*
b101 6
19
1>
1C
b101 G
#765680000000
0!
0*
09
0>
0C
#765690000000
1!
1*
b110 6
19
1>
1C
b110 G
#765700000000
0!
0*
09
0>
0C
#765710000000
1!
1*
b111 6
19
1>
1C
b111 G
#765720000000
0!
1"
0*
1+
09
1:
0>
0C
#765730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#765740000000
0!
0*
09
0>
0C
#765750000000
1!
1*
b1 6
19
1>
1C
b1 G
#765760000000
0!
0*
09
0>
0C
#765770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#765780000000
0!
0*
09
0>
0C
#765790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#765800000000
0!
0*
09
0>
0C
#765810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#765820000000
0!
0*
09
0>
0C
#765830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#765840000000
0!
0#
0*
0,
09
0>
0?
0C
#765850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#765860000000
0!
0*
09
0>
0C
#765870000000
1!
1*
19
1>
1C
#765880000000
0!
0*
09
0>
0C
#765890000000
1!
1*
19
1>
1C
#765900000000
0!
0*
09
0>
0C
#765910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#765920000000
0!
0*
09
0>
0C
#765930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#765940000000
0!
0*
09
0>
0C
#765950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#765960000000
0!
0*
09
0>
0C
#765970000000
1!
1*
b10 6
19
1>
1C
b10 G
#765980000000
0!
0*
09
0>
0C
#765990000000
1!
1*
b11 6
19
1>
1C
b11 G
#766000000000
0!
0*
09
0>
0C
#766010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#766020000000
0!
0*
09
0>
0C
#766030000000
1!
1*
b101 6
19
1>
1C
b101 G
#766040000000
0!
0*
09
0>
0C
#766050000000
1!
1*
b110 6
19
1>
1C
b110 G
#766060000000
0!
0*
09
0>
0C
#766070000000
1!
1*
b111 6
19
1>
1C
b111 G
#766080000000
0!
0*
09
0>
0C
#766090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#766100000000
0!
0*
09
0>
0C
#766110000000
1!
1*
b1 6
19
1>
1C
b1 G
#766120000000
0!
0*
09
0>
0C
#766130000000
1!
1*
b10 6
19
1>
1C
b10 G
#766140000000
0!
0*
09
0>
0C
#766150000000
1!
1*
b11 6
19
1>
1C
b11 G
#766160000000
0!
0*
09
0>
0C
#766170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#766180000000
0!
0*
09
0>
0C
#766190000000
1!
1*
b101 6
19
1>
1C
b101 G
#766200000000
0!
0*
09
0>
0C
#766210000000
1!
1*
b110 6
19
1>
1C
b110 G
#766220000000
0!
0*
09
0>
0C
#766230000000
1!
1*
b111 6
19
1>
1C
b111 G
#766240000000
0!
0*
09
0>
0C
#766250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#766260000000
0!
0*
09
0>
0C
#766270000000
1!
1*
b1 6
19
1>
1C
b1 G
#766280000000
0!
0*
09
0>
0C
#766290000000
1!
1*
b10 6
19
1>
1C
b10 G
#766300000000
0!
0*
09
0>
0C
#766310000000
1!
1*
b11 6
19
1>
1C
b11 G
#766320000000
0!
0*
09
0>
0C
#766330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#766340000000
0!
0*
09
0>
0C
#766350000000
1!
1*
b101 6
19
1>
1C
b101 G
#766360000000
0!
0*
09
0>
0C
#766370000000
1!
1*
b110 6
19
1>
1C
b110 G
#766380000000
0!
0*
09
0>
0C
#766390000000
1!
1*
b111 6
19
1>
1C
b111 G
#766400000000
0!
1"
0*
1+
09
1:
0>
0C
#766410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#766420000000
0!
0*
09
0>
0C
#766430000000
1!
1*
b1 6
19
1>
1C
b1 G
#766440000000
0!
0*
09
0>
0C
#766450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#766460000000
0!
0*
09
0>
0C
#766470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#766480000000
0!
0*
09
0>
0C
#766490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#766500000000
0!
0*
09
0>
0C
#766510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#766520000000
0!
0#
0*
0,
09
0>
0?
0C
#766530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#766540000000
0!
0*
09
0>
0C
#766550000000
1!
1*
19
1>
1C
#766560000000
0!
0*
09
0>
0C
#766570000000
1!
1*
19
1>
1C
#766580000000
0!
0*
09
0>
0C
#766590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#766600000000
0!
0*
09
0>
0C
#766610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#766620000000
0!
0*
09
0>
0C
#766630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#766640000000
0!
0*
09
0>
0C
#766650000000
1!
1*
b10 6
19
1>
1C
b10 G
#766660000000
0!
0*
09
0>
0C
#766670000000
1!
1*
b11 6
19
1>
1C
b11 G
#766680000000
0!
0*
09
0>
0C
#766690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#766700000000
0!
0*
09
0>
0C
#766710000000
1!
1*
b101 6
19
1>
1C
b101 G
#766720000000
0!
0*
09
0>
0C
#766730000000
1!
1*
b110 6
19
1>
1C
b110 G
#766740000000
0!
0*
09
0>
0C
#766750000000
1!
1*
b111 6
19
1>
1C
b111 G
#766760000000
0!
0*
09
0>
0C
#766770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#766780000000
0!
0*
09
0>
0C
#766790000000
1!
1*
b1 6
19
1>
1C
b1 G
#766800000000
0!
0*
09
0>
0C
#766810000000
1!
1*
b10 6
19
1>
1C
b10 G
#766820000000
0!
0*
09
0>
0C
#766830000000
1!
1*
b11 6
19
1>
1C
b11 G
#766840000000
0!
0*
09
0>
0C
#766850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#766860000000
0!
0*
09
0>
0C
#766870000000
1!
1*
b101 6
19
1>
1C
b101 G
#766880000000
0!
0*
09
0>
0C
#766890000000
1!
1*
b110 6
19
1>
1C
b110 G
#766900000000
0!
0*
09
0>
0C
#766910000000
1!
1*
b111 6
19
1>
1C
b111 G
#766920000000
0!
0*
09
0>
0C
#766930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#766940000000
0!
0*
09
0>
0C
#766950000000
1!
1*
b1 6
19
1>
1C
b1 G
#766960000000
0!
0*
09
0>
0C
#766970000000
1!
1*
b10 6
19
1>
1C
b10 G
#766980000000
0!
0*
09
0>
0C
#766990000000
1!
1*
b11 6
19
1>
1C
b11 G
#767000000000
0!
0*
09
0>
0C
#767010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#767020000000
0!
0*
09
0>
0C
#767030000000
1!
1*
b101 6
19
1>
1C
b101 G
#767040000000
0!
0*
09
0>
0C
#767050000000
1!
1*
b110 6
19
1>
1C
b110 G
#767060000000
0!
0*
09
0>
0C
#767070000000
1!
1*
b111 6
19
1>
1C
b111 G
#767080000000
0!
1"
0*
1+
09
1:
0>
0C
#767090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#767100000000
0!
0*
09
0>
0C
#767110000000
1!
1*
b1 6
19
1>
1C
b1 G
#767120000000
0!
0*
09
0>
0C
#767130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#767140000000
0!
0*
09
0>
0C
#767150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#767160000000
0!
0*
09
0>
0C
#767170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#767180000000
0!
0*
09
0>
0C
#767190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#767200000000
0!
0#
0*
0,
09
0>
0?
0C
#767210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#767220000000
0!
0*
09
0>
0C
#767230000000
1!
1*
19
1>
1C
#767240000000
0!
0*
09
0>
0C
#767250000000
1!
1*
19
1>
1C
#767260000000
0!
0*
09
0>
0C
#767270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#767280000000
0!
0*
09
0>
0C
#767290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#767300000000
0!
0*
09
0>
0C
#767310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#767320000000
0!
0*
09
0>
0C
#767330000000
1!
1*
b10 6
19
1>
1C
b10 G
#767340000000
0!
0*
09
0>
0C
#767350000000
1!
1*
b11 6
19
1>
1C
b11 G
#767360000000
0!
0*
09
0>
0C
#767370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#767380000000
0!
0*
09
0>
0C
#767390000000
1!
1*
b101 6
19
1>
1C
b101 G
#767400000000
0!
0*
09
0>
0C
#767410000000
1!
1*
b110 6
19
1>
1C
b110 G
#767420000000
0!
0*
09
0>
0C
#767430000000
1!
1*
b111 6
19
1>
1C
b111 G
#767440000000
0!
0*
09
0>
0C
#767450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#767460000000
0!
0*
09
0>
0C
#767470000000
1!
1*
b1 6
19
1>
1C
b1 G
#767480000000
0!
0*
09
0>
0C
#767490000000
1!
1*
b10 6
19
1>
1C
b10 G
#767500000000
0!
0*
09
0>
0C
#767510000000
1!
1*
b11 6
19
1>
1C
b11 G
#767520000000
0!
0*
09
0>
0C
#767530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#767540000000
0!
0*
09
0>
0C
#767550000000
1!
1*
b101 6
19
1>
1C
b101 G
#767560000000
0!
0*
09
0>
0C
#767570000000
1!
1*
b110 6
19
1>
1C
b110 G
#767580000000
0!
0*
09
0>
0C
#767590000000
1!
1*
b111 6
19
1>
1C
b111 G
#767600000000
0!
0*
09
0>
0C
#767610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#767620000000
0!
0*
09
0>
0C
#767630000000
1!
1*
b1 6
19
1>
1C
b1 G
#767640000000
0!
0*
09
0>
0C
#767650000000
1!
1*
b10 6
19
1>
1C
b10 G
#767660000000
0!
0*
09
0>
0C
#767670000000
1!
1*
b11 6
19
1>
1C
b11 G
#767680000000
0!
0*
09
0>
0C
#767690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#767700000000
0!
0*
09
0>
0C
#767710000000
1!
1*
b101 6
19
1>
1C
b101 G
#767720000000
0!
0*
09
0>
0C
#767730000000
1!
1*
b110 6
19
1>
1C
b110 G
#767740000000
0!
0*
09
0>
0C
#767750000000
1!
1*
b111 6
19
1>
1C
b111 G
#767760000000
0!
1"
0*
1+
09
1:
0>
0C
#767770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#767780000000
0!
0*
09
0>
0C
#767790000000
1!
1*
b1 6
19
1>
1C
b1 G
#767800000000
0!
0*
09
0>
0C
#767810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#767820000000
0!
0*
09
0>
0C
#767830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#767840000000
0!
0*
09
0>
0C
#767850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#767860000000
0!
0*
09
0>
0C
#767870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#767880000000
0!
0#
0*
0,
09
0>
0?
0C
#767890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#767900000000
0!
0*
09
0>
0C
#767910000000
1!
1*
19
1>
1C
#767920000000
0!
0*
09
0>
0C
#767930000000
1!
1*
19
1>
1C
#767940000000
0!
0*
09
0>
0C
#767950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#767960000000
0!
0*
09
0>
0C
#767970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#767980000000
0!
0*
09
0>
0C
#767990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#768000000000
0!
0*
09
0>
0C
#768010000000
1!
1*
b10 6
19
1>
1C
b10 G
#768020000000
0!
0*
09
0>
0C
#768030000000
1!
1*
b11 6
19
1>
1C
b11 G
#768040000000
0!
0*
09
0>
0C
#768050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#768060000000
0!
0*
09
0>
0C
#768070000000
1!
1*
b101 6
19
1>
1C
b101 G
#768080000000
0!
0*
09
0>
0C
#768090000000
1!
1*
b110 6
19
1>
1C
b110 G
#768100000000
0!
0*
09
0>
0C
#768110000000
1!
1*
b111 6
19
1>
1C
b111 G
#768120000000
0!
0*
09
0>
0C
#768130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#768140000000
0!
0*
09
0>
0C
#768150000000
1!
1*
b1 6
19
1>
1C
b1 G
#768160000000
0!
0*
09
0>
0C
#768170000000
1!
1*
b10 6
19
1>
1C
b10 G
#768180000000
0!
0*
09
0>
0C
#768190000000
1!
1*
b11 6
19
1>
1C
b11 G
#768200000000
0!
0*
09
0>
0C
#768210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#768220000000
0!
0*
09
0>
0C
#768230000000
1!
1*
b101 6
19
1>
1C
b101 G
#768240000000
0!
0*
09
0>
0C
#768250000000
1!
1*
b110 6
19
1>
1C
b110 G
#768260000000
0!
0*
09
0>
0C
#768270000000
1!
1*
b111 6
19
1>
1C
b111 G
#768280000000
0!
0*
09
0>
0C
#768290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#768300000000
0!
0*
09
0>
0C
#768310000000
1!
1*
b1 6
19
1>
1C
b1 G
#768320000000
0!
0*
09
0>
0C
#768330000000
1!
1*
b10 6
19
1>
1C
b10 G
#768340000000
0!
0*
09
0>
0C
#768350000000
1!
1*
b11 6
19
1>
1C
b11 G
#768360000000
0!
0*
09
0>
0C
#768370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#768380000000
0!
0*
09
0>
0C
#768390000000
1!
1*
b101 6
19
1>
1C
b101 G
#768400000000
0!
0*
09
0>
0C
#768410000000
1!
1*
b110 6
19
1>
1C
b110 G
#768420000000
0!
0*
09
0>
0C
#768430000000
1!
1*
b111 6
19
1>
1C
b111 G
#768440000000
0!
1"
0*
1+
09
1:
0>
0C
#768450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#768460000000
0!
0*
09
0>
0C
#768470000000
1!
1*
b1 6
19
1>
1C
b1 G
#768480000000
0!
0*
09
0>
0C
#768490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#768500000000
0!
0*
09
0>
0C
#768510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#768520000000
0!
0*
09
0>
0C
#768530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#768540000000
0!
0*
09
0>
0C
#768550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#768560000000
0!
0#
0*
0,
09
0>
0?
0C
#768570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#768580000000
0!
0*
09
0>
0C
#768590000000
1!
1*
19
1>
1C
#768600000000
0!
0*
09
0>
0C
#768610000000
1!
1*
19
1>
1C
#768620000000
0!
0*
09
0>
0C
#768630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#768640000000
0!
0*
09
0>
0C
#768650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#768660000000
0!
0*
09
0>
0C
#768670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#768680000000
0!
0*
09
0>
0C
#768690000000
1!
1*
b10 6
19
1>
1C
b10 G
#768700000000
0!
0*
09
0>
0C
#768710000000
1!
1*
b11 6
19
1>
1C
b11 G
#768720000000
0!
0*
09
0>
0C
#768730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#768740000000
0!
0*
09
0>
0C
#768750000000
1!
1*
b101 6
19
1>
1C
b101 G
#768760000000
0!
0*
09
0>
0C
#768770000000
1!
1*
b110 6
19
1>
1C
b110 G
#768780000000
0!
0*
09
0>
0C
#768790000000
1!
1*
b111 6
19
1>
1C
b111 G
#768800000000
0!
0*
09
0>
0C
#768810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#768820000000
0!
0*
09
0>
0C
#768830000000
1!
1*
b1 6
19
1>
1C
b1 G
#768840000000
0!
0*
09
0>
0C
#768850000000
1!
1*
b10 6
19
1>
1C
b10 G
#768860000000
0!
0*
09
0>
0C
#768870000000
1!
1*
b11 6
19
1>
1C
b11 G
#768880000000
0!
0*
09
0>
0C
#768890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#768900000000
0!
0*
09
0>
0C
#768910000000
1!
1*
b101 6
19
1>
1C
b101 G
#768920000000
0!
0*
09
0>
0C
#768930000000
1!
1*
b110 6
19
1>
1C
b110 G
#768940000000
0!
0*
09
0>
0C
#768950000000
1!
1*
b111 6
19
1>
1C
b111 G
#768960000000
0!
0*
09
0>
0C
#768970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#768980000000
0!
0*
09
0>
0C
#768990000000
1!
1*
b1 6
19
1>
1C
b1 G
#769000000000
0!
0*
09
0>
0C
#769010000000
1!
1*
b10 6
19
1>
1C
b10 G
#769020000000
0!
0*
09
0>
0C
#769030000000
1!
1*
b11 6
19
1>
1C
b11 G
#769040000000
0!
0*
09
0>
0C
#769050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#769060000000
0!
0*
09
0>
0C
#769070000000
1!
1*
b101 6
19
1>
1C
b101 G
#769080000000
0!
0*
09
0>
0C
#769090000000
1!
1*
b110 6
19
1>
1C
b110 G
#769100000000
0!
0*
09
0>
0C
#769110000000
1!
1*
b111 6
19
1>
1C
b111 G
#769120000000
0!
1"
0*
1+
09
1:
0>
0C
#769130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#769140000000
0!
0*
09
0>
0C
#769150000000
1!
1*
b1 6
19
1>
1C
b1 G
#769160000000
0!
0*
09
0>
0C
#769170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#769180000000
0!
0*
09
0>
0C
#769190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#769200000000
0!
0*
09
0>
0C
#769210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#769220000000
0!
0*
09
0>
0C
#769230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#769240000000
0!
0#
0*
0,
09
0>
0?
0C
#769250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#769260000000
0!
0*
09
0>
0C
#769270000000
1!
1*
19
1>
1C
#769280000000
0!
0*
09
0>
0C
#769290000000
1!
1*
19
1>
1C
#769300000000
0!
0*
09
0>
0C
#769310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#769320000000
0!
0*
09
0>
0C
#769330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#769340000000
0!
0*
09
0>
0C
#769350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#769360000000
0!
0*
09
0>
0C
#769370000000
1!
1*
b10 6
19
1>
1C
b10 G
#769380000000
0!
0*
09
0>
0C
#769390000000
1!
1*
b11 6
19
1>
1C
b11 G
#769400000000
0!
0*
09
0>
0C
#769410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#769420000000
0!
0*
09
0>
0C
#769430000000
1!
1*
b101 6
19
1>
1C
b101 G
#769440000000
0!
0*
09
0>
0C
#769450000000
1!
1*
b110 6
19
1>
1C
b110 G
#769460000000
0!
0*
09
0>
0C
#769470000000
1!
1*
b111 6
19
1>
1C
b111 G
#769480000000
0!
0*
09
0>
0C
#769490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#769500000000
0!
0*
09
0>
0C
#769510000000
1!
1*
b1 6
19
1>
1C
b1 G
#769520000000
0!
0*
09
0>
0C
#769530000000
1!
1*
b10 6
19
1>
1C
b10 G
#769540000000
0!
0*
09
0>
0C
#769550000000
1!
1*
b11 6
19
1>
1C
b11 G
#769560000000
0!
0*
09
0>
0C
#769570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#769580000000
0!
0*
09
0>
0C
#769590000000
1!
1*
b101 6
19
1>
1C
b101 G
#769600000000
0!
0*
09
0>
0C
#769610000000
1!
1*
b110 6
19
1>
1C
b110 G
#769620000000
0!
0*
09
0>
0C
#769630000000
1!
1*
b111 6
19
1>
1C
b111 G
#769640000000
0!
0*
09
0>
0C
#769650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#769660000000
0!
0*
09
0>
0C
#769670000000
1!
1*
b1 6
19
1>
1C
b1 G
#769680000000
0!
0*
09
0>
0C
#769690000000
1!
1*
b10 6
19
1>
1C
b10 G
#769700000000
0!
0*
09
0>
0C
#769710000000
1!
1*
b11 6
19
1>
1C
b11 G
#769720000000
0!
0*
09
0>
0C
#769730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#769740000000
0!
0*
09
0>
0C
#769750000000
1!
1*
b101 6
19
1>
1C
b101 G
#769760000000
0!
0*
09
0>
0C
#769770000000
1!
1*
b110 6
19
1>
1C
b110 G
#769780000000
0!
0*
09
0>
0C
#769790000000
1!
1*
b111 6
19
1>
1C
b111 G
#769800000000
0!
1"
0*
1+
09
1:
0>
0C
#769810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#769820000000
0!
0*
09
0>
0C
#769830000000
1!
1*
b1 6
19
1>
1C
b1 G
#769840000000
0!
0*
09
0>
0C
#769850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#769860000000
0!
0*
09
0>
0C
#769870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#769880000000
0!
0*
09
0>
0C
#769890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#769900000000
0!
0*
09
0>
0C
#769910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#769920000000
0!
0#
0*
0,
09
0>
0?
0C
#769930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#769940000000
0!
0*
09
0>
0C
#769950000000
1!
1*
19
1>
1C
#769960000000
0!
0*
09
0>
0C
#769970000000
1!
1*
19
1>
1C
#769980000000
0!
0*
09
0>
0C
#769990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#770000000000
0!
0*
09
0>
0C
#770010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#770020000000
0!
0*
09
0>
0C
#770030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#770040000000
0!
0*
09
0>
0C
#770050000000
1!
1*
b10 6
19
1>
1C
b10 G
#770060000000
0!
0*
09
0>
0C
#770070000000
1!
1*
b11 6
19
1>
1C
b11 G
#770080000000
0!
0*
09
0>
0C
#770090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#770100000000
0!
0*
09
0>
0C
#770110000000
1!
1*
b101 6
19
1>
1C
b101 G
#770120000000
0!
0*
09
0>
0C
#770130000000
1!
1*
b110 6
19
1>
1C
b110 G
#770140000000
0!
0*
09
0>
0C
#770150000000
1!
1*
b111 6
19
1>
1C
b111 G
#770160000000
0!
0*
09
0>
0C
#770170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#770180000000
0!
0*
09
0>
0C
#770190000000
1!
1*
b1 6
19
1>
1C
b1 G
#770200000000
0!
0*
09
0>
0C
#770210000000
1!
1*
b10 6
19
1>
1C
b10 G
#770220000000
0!
0*
09
0>
0C
#770230000000
1!
1*
b11 6
19
1>
1C
b11 G
#770240000000
0!
0*
09
0>
0C
#770250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#770260000000
0!
0*
09
0>
0C
#770270000000
1!
1*
b101 6
19
1>
1C
b101 G
#770280000000
0!
0*
09
0>
0C
#770290000000
1!
1*
b110 6
19
1>
1C
b110 G
#770300000000
0!
0*
09
0>
0C
#770310000000
1!
1*
b111 6
19
1>
1C
b111 G
#770320000000
0!
0*
09
0>
0C
#770330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#770340000000
0!
0*
09
0>
0C
#770350000000
1!
1*
b1 6
19
1>
1C
b1 G
#770360000000
0!
0*
09
0>
0C
#770370000000
1!
1*
b10 6
19
1>
1C
b10 G
#770380000000
0!
0*
09
0>
0C
#770390000000
1!
1*
b11 6
19
1>
1C
b11 G
#770400000000
0!
0*
09
0>
0C
#770410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#770420000000
0!
0*
09
0>
0C
#770430000000
1!
1*
b101 6
19
1>
1C
b101 G
#770440000000
0!
0*
09
0>
0C
#770450000000
1!
1*
b110 6
19
1>
1C
b110 G
#770460000000
0!
0*
09
0>
0C
#770470000000
1!
1*
b111 6
19
1>
1C
b111 G
#770480000000
0!
1"
0*
1+
09
1:
0>
0C
#770490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#770500000000
0!
0*
09
0>
0C
#770510000000
1!
1*
b1 6
19
1>
1C
b1 G
#770520000000
0!
0*
09
0>
0C
#770530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#770540000000
0!
0*
09
0>
0C
#770550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#770560000000
0!
0*
09
0>
0C
#770570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#770580000000
0!
0*
09
0>
0C
#770590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#770600000000
0!
0#
0*
0,
09
0>
0?
0C
#770610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#770620000000
0!
0*
09
0>
0C
#770630000000
1!
1*
19
1>
1C
#770640000000
0!
0*
09
0>
0C
#770650000000
1!
1*
19
1>
1C
#770660000000
0!
0*
09
0>
0C
#770670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#770680000000
0!
0*
09
0>
0C
#770690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#770700000000
0!
0*
09
0>
0C
#770710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#770720000000
0!
0*
09
0>
0C
#770730000000
1!
1*
b10 6
19
1>
1C
b10 G
#770740000000
0!
0*
09
0>
0C
#770750000000
1!
1*
b11 6
19
1>
1C
b11 G
#770760000000
0!
0*
09
0>
0C
#770770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#770780000000
0!
0*
09
0>
0C
#770790000000
1!
1*
b101 6
19
1>
1C
b101 G
#770800000000
0!
0*
09
0>
0C
#770810000000
1!
1*
b110 6
19
1>
1C
b110 G
#770820000000
0!
0*
09
0>
0C
#770830000000
1!
1*
b111 6
19
1>
1C
b111 G
#770840000000
0!
0*
09
0>
0C
#770850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#770860000000
0!
0*
09
0>
0C
#770870000000
1!
1*
b1 6
19
1>
1C
b1 G
#770880000000
0!
0*
09
0>
0C
#770890000000
1!
1*
b10 6
19
1>
1C
b10 G
#770900000000
0!
0*
09
0>
0C
#770910000000
1!
1*
b11 6
19
1>
1C
b11 G
#770920000000
0!
0*
09
0>
0C
#770930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#770940000000
0!
0*
09
0>
0C
#770950000000
1!
1*
b101 6
19
1>
1C
b101 G
#770960000000
0!
0*
09
0>
0C
#770970000000
1!
1*
b110 6
19
1>
1C
b110 G
#770980000000
0!
0*
09
0>
0C
#770990000000
1!
1*
b111 6
19
1>
1C
b111 G
#771000000000
0!
0*
09
0>
0C
#771010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#771020000000
0!
0*
09
0>
0C
#771030000000
1!
1*
b1 6
19
1>
1C
b1 G
#771040000000
0!
0*
09
0>
0C
#771050000000
1!
1*
b10 6
19
1>
1C
b10 G
#771060000000
0!
0*
09
0>
0C
#771070000000
1!
1*
b11 6
19
1>
1C
b11 G
#771080000000
0!
0*
09
0>
0C
#771090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#771100000000
0!
0*
09
0>
0C
#771110000000
1!
1*
b101 6
19
1>
1C
b101 G
#771120000000
0!
0*
09
0>
0C
#771130000000
1!
1*
b110 6
19
1>
1C
b110 G
#771140000000
0!
0*
09
0>
0C
#771150000000
1!
1*
b111 6
19
1>
1C
b111 G
#771160000000
0!
1"
0*
1+
09
1:
0>
0C
#771170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#771180000000
0!
0*
09
0>
0C
#771190000000
1!
1*
b1 6
19
1>
1C
b1 G
#771200000000
0!
0*
09
0>
0C
#771210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#771220000000
0!
0*
09
0>
0C
#771230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#771240000000
0!
0*
09
0>
0C
#771250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#771260000000
0!
0*
09
0>
0C
#771270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#771280000000
0!
0#
0*
0,
09
0>
0?
0C
#771290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#771300000000
0!
0*
09
0>
0C
#771310000000
1!
1*
19
1>
1C
#771320000000
0!
0*
09
0>
0C
#771330000000
1!
1*
19
1>
1C
#771340000000
0!
0*
09
0>
0C
#771350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#771360000000
0!
0*
09
0>
0C
#771370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#771380000000
0!
0*
09
0>
0C
#771390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#771400000000
0!
0*
09
0>
0C
#771410000000
1!
1*
b10 6
19
1>
1C
b10 G
#771420000000
0!
0*
09
0>
0C
#771430000000
1!
1*
b11 6
19
1>
1C
b11 G
#771440000000
0!
0*
09
0>
0C
#771450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#771460000000
0!
0*
09
0>
0C
#771470000000
1!
1*
b101 6
19
1>
1C
b101 G
#771480000000
0!
0*
09
0>
0C
#771490000000
1!
1*
b110 6
19
1>
1C
b110 G
#771500000000
0!
0*
09
0>
0C
#771510000000
1!
1*
b111 6
19
1>
1C
b111 G
#771520000000
0!
0*
09
0>
0C
#771530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#771540000000
0!
0*
09
0>
0C
#771550000000
1!
1*
b1 6
19
1>
1C
b1 G
#771560000000
0!
0*
09
0>
0C
#771570000000
1!
1*
b10 6
19
1>
1C
b10 G
#771580000000
0!
0*
09
0>
0C
#771590000000
1!
1*
b11 6
19
1>
1C
b11 G
#771600000000
0!
0*
09
0>
0C
#771610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#771620000000
0!
0*
09
0>
0C
#771630000000
1!
1*
b101 6
19
1>
1C
b101 G
#771640000000
0!
0*
09
0>
0C
#771650000000
1!
1*
b110 6
19
1>
1C
b110 G
#771660000000
0!
0*
09
0>
0C
#771670000000
1!
1*
b111 6
19
1>
1C
b111 G
#771680000000
0!
0*
09
0>
0C
#771690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#771700000000
0!
0*
09
0>
0C
#771710000000
1!
1*
b1 6
19
1>
1C
b1 G
#771720000000
0!
0*
09
0>
0C
#771730000000
1!
1*
b10 6
19
1>
1C
b10 G
#771740000000
0!
0*
09
0>
0C
#771750000000
1!
1*
b11 6
19
1>
1C
b11 G
#771760000000
0!
0*
09
0>
0C
#771770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#771780000000
0!
0*
09
0>
0C
#771790000000
1!
1*
b101 6
19
1>
1C
b101 G
#771800000000
0!
0*
09
0>
0C
#771810000000
1!
1*
b110 6
19
1>
1C
b110 G
#771820000000
0!
0*
09
0>
0C
#771830000000
1!
1*
b111 6
19
1>
1C
b111 G
#771840000000
0!
1"
0*
1+
09
1:
0>
0C
#771850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#771860000000
0!
0*
09
0>
0C
#771870000000
1!
1*
b1 6
19
1>
1C
b1 G
#771880000000
0!
0*
09
0>
0C
#771890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#771900000000
0!
0*
09
0>
0C
#771910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#771920000000
0!
0*
09
0>
0C
#771930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#771940000000
0!
0*
09
0>
0C
#771950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#771960000000
0!
0#
0*
0,
09
0>
0?
0C
#771970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#771980000000
0!
0*
09
0>
0C
#771990000000
1!
1*
19
1>
1C
#772000000000
0!
0*
09
0>
0C
#772010000000
1!
1*
19
1>
1C
#772020000000
0!
0*
09
0>
0C
#772030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#772040000000
0!
0*
09
0>
0C
#772050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#772060000000
0!
0*
09
0>
0C
#772070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#772080000000
0!
0*
09
0>
0C
#772090000000
1!
1*
b10 6
19
1>
1C
b10 G
#772100000000
0!
0*
09
0>
0C
#772110000000
1!
1*
b11 6
19
1>
1C
b11 G
#772120000000
0!
0*
09
0>
0C
#772130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#772140000000
0!
0*
09
0>
0C
#772150000000
1!
1*
b101 6
19
1>
1C
b101 G
#772160000000
0!
0*
09
0>
0C
#772170000000
1!
1*
b110 6
19
1>
1C
b110 G
#772180000000
0!
0*
09
0>
0C
#772190000000
1!
1*
b111 6
19
1>
1C
b111 G
#772200000000
0!
0*
09
0>
0C
#772210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#772220000000
0!
0*
09
0>
0C
#772230000000
1!
1*
b1 6
19
1>
1C
b1 G
#772240000000
0!
0*
09
0>
0C
#772250000000
1!
1*
b10 6
19
1>
1C
b10 G
#772260000000
0!
0*
09
0>
0C
#772270000000
1!
1*
b11 6
19
1>
1C
b11 G
#772280000000
0!
0*
09
0>
0C
#772290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#772300000000
0!
0*
09
0>
0C
#772310000000
1!
1*
b101 6
19
1>
1C
b101 G
#772320000000
0!
0*
09
0>
0C
#772330000000
1!
1*
b110 6
19
1>
1C
b110 G
#772340000000
0!
0*
09
0>
0C
#772350000000
1!
1*
b111 6
19
1>
1C
b111 G
#772360000000
0!
0*
09
0>
0C
#772370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#772380000000
0!
0*
09
0>
0C
#772390000000
1!
1*
b1 6
19
1>
1C
b1 G
#772400000000
0!
0*
09
0>
0C
#772410000000
1!
1*
b10 6
19
1>
1C
b10 G
#772420000000
0!
0*
09
0>
0C
#772430000000
1!
1*
b11 6
19
1>
1C
b11 G
#772440000000
0!
0*
09
0>
0C
#772450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#772460000000
0!
0*
09
0>
0C
#772470000000
1!
1*
b101 6
19
1>
1C
b101 G
#772480000000
0!
0*
09
0>
0C
#772490000000
1!
1*
b110 6
19
1>
1C
b110 G
#772500000000
0!
0*
09
0>
0C
#772510000000
1!
1*
b111 6
19
1>
1C
b111 G
#772520000000
0!
1"
0*
1+
09
1:
0>
0C
#772530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#772540000000
0!
0*
09
0>
0C
#772550000000
1!
1*
b1 6
19
1>
1C
b1 G
#772560000000
0!
0*
09
0>
0C
#772570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#772580000000
0!
0*
09
0>
0C
#772590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#772600000000
0!
0*
09
0>
0C
#772610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#772620000000
0!
0*
09
0>
0C
#772630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#772640000000
0!
0#
0*
0,
09
0>
0?
0C
#772650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#772660000000
0!
0*
09
0>
0C
#772670000000
1!
1*
19
1>
1C
#772680000000
0!
0*
09
0>
0C
#772690000000
1!
1*
19
1>
1C
#772700000000
0!
0*
09
0>
0C
#772710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#772720000000
0!
0*
09
0>
0C
#772730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#772740000000
0!
0*
09
0>
0C
#772750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#772760000000
0!
0*
09
0>
0C
#772770000000
1!
1*
b10 6
19
1>
1C
b10 G
#772780000000
0!
0*
09
0>
0C
#772790000000
1!
1*
b11 6
19
1>
1C
b11 G
#772800000000
0!
0*
09
0>
0C
#772810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#772820000000
0!
0*
09
0>
0C
#772830000000
1!
1*
b101 6
19
1>
1C
b101 G
#772840000000
0!
0*
09
0>
0C
#772850000000
1!
1*
b110 6
19
1>
1C
b110 G
#772860000000
0!
0*
09
0>
0C
#772870000000
1!
1*
b111 6
19
1>
1C
b111 G
#772880000000
0!
0*
09
0>
0C
#772890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#772900000000
0!
0*
09
0>
0C
#772910000000
1!
1*
b1 6
19
1>
1C
b1 G
#772920000000
0!
0*
09
0>
0C
#772930000000
1!
1*
b10 6
19
1>
1C
b10 G
#772940000000
0!
0*
09
0>
0C
#772950000000
1!
1*
b11 6
19
1>
1C
b11 G
#772960000000
0!
0*
09
0>
0C
#772970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#772980000000
0!
0*
09
0>
0C
#772990000000
1!
1*
b101 6
19
1>
1C
b101 G
#773000000000
0!
0*
09
0>
0C
#773010000000
1!
1*
b110 6
19
1>
1C
b110 G
#773020000000
0!
0*
09
0>
0C
#773030000000
1!
1*
b111 6
19
1>
1C
b111 G
#773040000000
0!
0*
09
0>
0C
#773050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#773060000000
0!
0*
09
0>
0C
#773070000000
1!
1*
b1 6
19
1>
1C
b1 G
#773080000000
0!
0*
09
0>
0C
#773090000000
1!
1*
b10 6
19
1>
1C
b10 G
#773100000000
0!
0*
09
0>
0C
#773110000000
1!
1*
b11 6
19
1>
1C
b11 G
#773120000000
0!
0*
09
0>
0C
#773130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#773140000000
0!
0*
09
0>
0C
#773150000000
1!
1*
b101 6
19
1>
1C
b101 G
#773160000000
0!
0*
09
0>
0C
#773170000000
1!
1*
b110 6
19
1>
1C
b110 G
#773180000000
0!
0*
09
0>
0C
#773190000000
1!
1*
b111 6
19
1>
1C
b111 G
#773200000000
0!
1"
0*
1+
09
1:
0>
0C
#773210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#773220000000
0!
0*
09
0>
0C
#773230000000
1!
1*
b1 6
19
1>
1C
b1 G
#773240000000
0!
0*
09
0>
0C
#773250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#773260000000
0!
0*
09
0>
0C
#773270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#773280000000
0!
0*
09
0>
0C
#773290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#773300000000
0!
0*
09
0>
0C
#773310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#773320000000
0!
0#
0*
0,
09
0>
0?
0C
#773330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#773340000000
0!
0*
09
0>
0C
#773350000000
1!
1*
19
1>
1C
#773360000000
0!
0*
09
0>
0C
#773370000000
1!
1*
19
1>
1C
#773380000000
0!
0*
09
0>
0C
#773390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#773400000000
0!
0*
09
0>
0C
#773410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#773420000000
0!
0*
09
0>
0C
#773430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#773440000000
0!
0*
09
0>
0C
#773450000000
1!
1*
b10 6
19
1>
1C
b10 G
#773460000000
0!
0*
09
0>
0C
#773470000000
1!
1*
b11 6
19
1>
1C
b11 G
#773480000000
0!
0*
09
0>
0C
#773490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#773500000000
0!
0*
09
0>
0C
#773510000000
1!
1*
b101 6
19
1>
1C
b101 G
#773520000000
0!
0*
09
0>
0C
#773530000000
1!
1*
b110 6
19
1>
1C
b110 G
#773540000000
0!
0*
09
0>
0C
#773550000000
1!
1*
b111 6
19
1>
1C
b111 G
#773560000000
0!
0*
09
0>
0C
#773570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#773580000000
0!
0*
09
0>
0C
#773590000000
1!
1*
b1 6
19
1>
1C
b1 G
#773600000000
0!
0*
09
0>
0C
#773610000000
1!
1*
b10 6
19
1>
1C
b10 G
#773620000000
0!
0*
09
0>
0C
#773630000000
1!
1*
b11 6
19
1>
1C
b11 G
#773640000000
0!
0*
09
0>
0C
#773650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#773660000000
0!
0*
09
0>
0C
#773670000000
1!
1*
b101 6
19
1>
1C
b101 G
#773680000000
0!
0*
09
0>
0C
#773690000000
1!
1*
b110 6
19
1>
1C
b110 G
#773700000000
0!
0*
09
0>
0C
#773710000000
1!
1*
b111 6
19
1>
1C
b111 G
#773720000000
0!
0*
09
0>
0C
#773730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#773740000000
0!
0*
09
0>
0C
#773750000000
1!
1*
b1 6
19
1>
1C
b1 G
#773760000000
0!
0*
09
0>
0C
#773770000000
1!
1*
b10 6
19
1>
1C
b10 G
#773780000000
0!
0*
09
0>
0C
#773790000000
1!
1*
b11 6
19
1>
1C
b11 G
#773800000000
0!
0*
09
0>
0C
#773810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#773820000000
0!
0*
09
0>
0C
#773830000000
1!
1*
b101 6
19
1>
1C
b101 G
#773840000000
0!
0*
09
0>
0C
#773850000000
1!
1*
b110 6
19
1>
1C
b110 G
#773860000000
0!
0*
09
0>
0C
#773870000000
1!
1*
b111 6
19
1>
1C
b111 G
#773880000000
0!
1"
0*
1+
09
1:
0>
0C
#773890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#773900000000
0!
0*
09
0>
0C
#773910000000
1!
1*
b1 6
19
1>
1C
b1 G
#773920000000
0!
0*
09
0>
0C
#773930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#773940000000
0!
0*
09
0>
0C
#773950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#773960000000
0!
0*
09
0>
0C
#773970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#773980000000
0!
0*
09
0>
0C
#773990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#774000000000
0!
0#
0*
0,
09
0>
0?
0C
#774010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#774020000000
0!
0*
09
0>
0C
#774030000000
1!
1*
19
1>
1C
#774040000000
0!
0*
09
0>
0C
#774050000000
1!
1*
19
1>
1C
#774060000000
0!
0*
09
0>
0C
#774070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#774080000000
0!
0*
09
0>
0C
#774090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#774100000000
0!
0*
09
0>
0C
#774110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#774120000000
0!
0*
09
0>
0C
#774130000000
1!
1*
b10 6
19
1>
1C
b10 G
#774140000000
0!
0*
09
0>
0C
#774150000000
1!
1*
b11 6
19
1>
1C
b11 G
#774160000000
0!
0*
09
0>
0C
#774170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#774180000000
0!
0*
09
0>
0C
#774190000000
1!
1*
b101 6
19
1>
1C
b101 G
#774200000000
0!
0*
09
0>
0C
#774210000000
1!
1*
b110 6
19
1>
1C
b110 G
#774220000000
0!
0*
09
0>
0C
#774230000000
1!
1*
b111 6
19
1>
1C
b111 G
#774240000000
0!
0*
09
0>
0C
#774250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#774260000000
0!
0*
09
0>
0C
#774270000000
1!
1*
b1 6
19
1>
1C
b1 G
#774280000000
0!
0*
09
0>
0C
#774290000000
1!
1*
b10 6
19
1>
1C
b10 G
#774300000000
0!
0*
09
0>
0C
#774310000000
1!
1*
b11 6
19
1>
1C
b11 G
#774320000000
0!
0*
09
0>
0C
#774330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#774340000000
0!
0*
09
0>
0C
#774350000000
1!
1*
b101 6
19
1>
1C
b101 G
#774360000000
0!
0*
09
0>
0C
#774370000000
1!
1*
b110 6
19
1>
1C
b110 G
#774380000000
0!
0*
09
0>
0C
#774390000000
1!
1*
b111 6
19
1>
1C
b111 G
#774400000000
0!
0*
09
0>
0C
#774410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#774420000000
0!
0*
09
0>
0C
#774430000000
1!
1*
b1 6
19
1>
1C
b1 G
#774440000000
0!
0*
09
0>
0C
#774450000000
1!
1*
b10 6
19
1>
1C
b10 G
#774460000000
0!
0*
09
0>
0C
#774470000000
1!
1*
b11 6
19
1>
1C
b11 G
#774480000000
0!
0*
09
0>
0C
#774490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#774500000000
0!
0*
09
0>
0C
#774510000000
1!
1*
b101 6
19
1>
1C
b101 G
#774520000000
0!
0*
09
0>
0C
#774530000000
1!
1*
b110 6
19
1>
1C
b110 G
#774540000000
0!
0*
09
0>
0C
#774550000000
1!
1*
b111 6
19
1>
1C
b111 G
#774560000000
0!
1"
0*
1+
09
1:
0>
0C
#774570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#774580000000
0!
0*
09
0>
0C
#774590000000
1!
1*
b1 6
19
1>
1C
b1 G
#774600000000
0!
0*
09
0>
0C
#774610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#774620000000
0!
0*
09
0>
0C
#774630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#774640000000
0!
0*
09
0>
0C
#774650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#774660000000
0!
0*
09
0>
0C
#774670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#774680000000
0!
0#
0*
0,
09
0>
0?
0C
#774690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#774700000000
0!
0*
09
0>
0C
#774710000000
1!
1*
19
1>
1C
#774720000000
0!
0*
09
0>
0C
#774730000000
1!
1*
19
1>
1C
#774740000000
0!
0*
09
0>
0C
#774750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#774760000000
0!
0*
09
0>
0C
#774770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#774780000000
0!
0*
09
0>
0C
#774790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#774800000000
0!
0*
09
0>
0C
#774810000000
1!
1*
b10 6
19
1>
1C
b10 G
#774820000000
0!
0*
09
0>
0C
#774830000000
1!
1*
b11 6
19
1>
1C
b11 G
#774840000000
0!
0*
09
0>
0C
#774850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#774860000000
0!
0*
09
0>
0C
#774870000000
1!
1*
b101 6
19
1>
1C
b101 G
#774880000000
0!
0*
09
0>
0C
#774890000000
1!
1*
b110 6
19
1>
1C
b110 G
#774900000000
0!
0*
09
0>
0C
#774910000000
1!
1*
b111 6
19
1>
1C
b111 G
#774920000000
0!
0*
09
0>
0C
#774930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#774940000000
0!
0*
09
0>
0C
#774950000000
1!
1*
b1 6
19
1>
1C
b1 G
#774960000000
0!
0*
09
0>
0C
#774970000000
1!
1*
b10 6
19
1>
1C
b10 G
#774980000000
0!
0*
09
0>
0C
#774990000000
1!
1*
b11 6
19
1>
1C
b11 G
#775000000000
0!
0*
09
0>
0C
#775010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#775020000000
0!
0*
09
0>
0C
#775030000000
1!
1*
b101 6
19
1>
1C
b101 G
#775040000000
0!
0*
09
0>
0C
#775050000000
1!
1*
b110 6
19
1>
1C
b110 G
#775060000000
0!
0*
09
0>
0C
#775070000000
1!
1*
b111 6
19
1>
1C
b111 G
#775080000000
0!
0*
09
0>
0C
#775090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#775100000000
0!
0*
09
0>
0C
#775110000000
1!
1*
b1 6
19
1>
1C
b1 G
#775120000000
0!
0*
09
0>
0C
#775130000000
1!
1*
b10 6
19
1>
1C
b10 G
#775140000000
0!
0*
09
0>
0C
#775150000000
1!
1*
b11 6
19
1>
1C
b11 G
#775160000000
0!
0*
09
0>
0C
#775170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#775180000000
0!
0*
09
0>
0C
#775190000000
1!
1*
b101 6
19
1>
1C
b101 G
#775200000000
0!
0*
09
0>
0C
#775210000000
1!
1*
b110 6
19
1>
1C
b110 G
#775220000000
0!
0*
09
0>
0C
#775230000000
1!
1*
b111 6
19
1>
1C
b111 G
#775240000000
0!
1"
0*
1+
09
1:
0>
0C
#775250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#775260000000
0!
0*
09
0>
0C
#775270000000
1!
1*
b1 6
19
1>
1C
b1 G
#775280000000
0!
0*
09
0>
0C
#775290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#775300000000
0!
0*
09
0>
0C
#775310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#775320000000
0!
0*
09
0>
0C
#775330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#775340000000
0!
0*
09
0>
0C
#775350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#775360000000
0!
0#
0*
0,
09
0>
0?
0C
#775370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#775380000000
0!
0*
09
0>
0C
#775390000000
1!
1*
19
1>
1C
#775400000000
0!
0*
09
0>
0C
#775410000000
1!
1*
19
1>
1C
#775420000000
0!
0*
09
0>
0C
#775430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#775440000000
0!
0*
09
0>
0C
#775450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#775460000000
0!
0*
09
0>
0C
#775470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#775480000000
0!
0*
09
0>
0C
#775490000000
1!
1*
b10 6
19
1>
1C
b10 G
#775500000000
0!
0*
09
0>
0C
#775510000000
1!
1*
b11 6
19
1>
1C
b11 G
#775520000000
0!
0*
09
0>
0C
#775530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#775540000000
0!
0*
09
0>
0C
#775550000000
1!
1*
b101 6
19
1>
1C
b101 G
#775560000000
0!
0*
09
0>
0C
#775570000000
1!
1*
b110 6
19
1>
1C
b110 G
#775580000000
0!
0*
09
0>
0C
#775590000000
1!
1*
b111 6
19
1>
1C
b111 G
#775600000000
0!
0*
09
0>
0C
#775610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#775620000000
0!
0*
09
0>
0C
#775630000000
1!
1*
b1 6
19
1>
1C
b1 G
#775640000000
0!
0*
09
0>
0C
#775650000000
1!
1*
b10 6
19
1>
1C
b10 G
#775660000000
0!
0*
09
0>
0C
#775670000000
1!
1*
b11 6
19
1>
1C
b11 G
#775680000000
0!
0*
09
0>
0C
#775690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#775700000000
0!
0*
09
0>
0C
#775710000000
1!
1*
b101 6
19
1>
1C
b101 G
#775720000000
0!
0*
09
0>
0C
#775730000000
1!
1*
b110 6
19
1>
1C
b110 G
#775740000000
0!
0*
09
0>
0C
#775750000000
1!
1*
b111 6
19
1>
1C
b111 G
#775760000000
0!
0*
09
0>
0C
#775770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#775780000000
0!
0*
09
0>
0C
#775790000000
1!
1*
b1 6
19
1>
1C
b1 G
#775800000000
0!
0*
09
0>
0C
#775810000000
1!
1*
b10 6
19
1>
1C
b10 G
#775820000000
0!
0*
09
0>
0C
#775830000000
1!
1*
b11 6
19
1>
1C
b11 G
#775840000000
0!
0*
09
0>
0C
#775850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#775860000000
0!
0*
09
0>
0C
#775870000000
1!
1*
b101 6
19
1>
1C
b101 G
#775880000000
0!
0*
09
0>
0C
#775890000000
1!
1*
b110 6
19
1>
1C
b110 G
#775900000000
0!
0*
09
0>
0C
#775910000000
1!
1*
b111 6
19
1>
1C
b111 G
#775920000000
0!
1"
0*
1+
09
1:
0>
0C
#775930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#775940000000
0!
0*
09
0>
0C
#775950000000
1!
1*
b1 6
19
1>
1C
b1 G
#775960000000
0!
0*
09
0>
0C
#775970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#775980000000
0!
0*
09
0>
0C
#775990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#776000000000
0!
0*
09
0>
0C
#776010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#776020000000
0!
0*
09
0>
0C
#776030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#776040000000
0!
0#
0*
0,
09
0>
0?
0C
#776050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#776060000000
0!
0*
09
0>
0C
#776070000000
1!
1*
19
1>
1C
#776080000000
0!
0*
09
0>
0C
#776090000000
1!
1*
19
1>
1C
#776100000000
0!
0*
09
0>
0C
#776110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#776120000000
0!
0*
09
0>
0C
#776130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#776140000000
0!
0*
09
0>
0C
#776150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#776160000000
0!
0*
09
0>
0C
#776170000000
1!
1*
b10 6
19
1>
1C
b10 G
#776180000000
0!
0*
09
0>
0C
#776190000000
1!
1*
b11 6
19
1>
1C
b11 G
#776200000000
0!
0*
09
0>
0C
#776210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#776220000000
0!
0*
09
0>
0C
#776230000000
1!
1*
b101 6
19
1>
1C
b101 G
#776240000000
0!
0*
09
0>
0C
#776250000000
1!
1*
b110 6
19
1>
1C
b110 G
#776260000000
0!
0*
09
0>
0C
#776270000000
1!
1*
b111 6
19
1>
1C
b111 G
#776280000000
0!
0*
09
0>
0C
#776290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#776300000000
0!
0*
09
0>
0C
#776310000000
1!
1*
b1 6
19
1>
1C
b1 G
#776320000000
0!
0*
09
0>
0C
#776330000000
1!
1*
b10 6
19
1>
1C
b10 G
#776340000000
0!
0*
09
0>
0C
#776350000000
1!
1*
b11 6
19
1>
1C
b11 G
#776360000000
0!
0*
09
0>
0C
#776370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#776380000000
0!
0*
09
0>
0C
#776390000000
1!
1*
b101 6
19
1>
1C
b101 G
#776400000000
0!
0*
09
0>
0C
#776410000000
1!
1*
b110 6
19
1>
1C
b110 G
#776420000000
0!
0*
09
0>
0C
#776430000000
1!
1*
b111 6
19
1>
1C
b111 G
#776440000000
0!
0*
09
0>
0C
#776450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#776460000000
0!
0*
09
0>
0C
#776470000000
1!
1*
b1 6
19
1>
1C
b1 G
#776480000000
0!
0*
09
0>
0C
#776490000000
1!
1*
b10 6
19
1>
1C
b10 G
#776500000000
0!
0*
09
0>
0C
#776510000000
1!
1*
b11 6
19
1>
1C
b11 G
#776520000000
0!
0*
09
0>
0C
#776530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#776540000000
0!
0*
09
0>
0C
#776550000000
1!
1*
b101 6
19
1>
1C
b101 G
#776560000000
0!
0*
09
0>
0C
#776570000000
1!
1*
b110 6
19
1>
1C
b110 G
#776580000000
0!
0*
09
0>
0C
#776590000000
1!
1*
b111 6
19
1>
1C
b111 G
#776600000000
0!
1"
0*
1+
09
1:
0>
0C
#776610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#776620000000
0!
0*
09
0>
0C
#776630000000
1!
1*
b1 6
19
1>
1C
b1 G
#776640000000
0!
0*
09
0>
0C
#776650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#776660000000
0!
0*
09
0>
0C
#776670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#776680000000
0!
0*
09
0>
0C
#776690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#776700000000
0!
0*
09
0>
0C
#776710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#776720000000
0!
0#
0*
0,
09
0>
0?
0C
#776730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#776740000000
0!
0*
09
0>
0C
#776750000000
1!
1*
19
1>
1C
#776760000000
0!
0*
09
0>
0C
#776770000000
1!
1*
19
1>
1C
#776780000000
0!
0*
09
0>
0C
#776790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#776800000000
0!
0*
09
0>
0C
#776810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#776820000000
0!
0*
09
0>
0C
#776830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#776840000000
0!
0*
09
0>
0C
#776850000000
1!
1*
b10 6
19
1>
1C
b10 G
#776860000000
0!
0*
09
0>
0C
#776870000000
1!
1*
b11 6
19
1>
1C
b11 G
#776880000000
0!
0*
09
0>
0C
#776890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#776900000000
0!
0*
09
0>
0C
#776910000000
1!
1*
b101 6
19
1>
1C
b101 G
#776920000000
0!
0*
09
0>
0C
#776930000000
1!
1*
b110 6
19
1>
1C
b110 G
#776940000000
0!
0*
09
0>
0C
#776950000000
1!
1*
b111 6
19
1>
1C
b111 G
#776960000000
0!
0*
09
0>
0C
#776970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#776980000000
0!
0*
09
0>
0C
#776990000000
1!
1*
b1 6
19
1>
1C
b1 G
#777000000000
0!
0*
09
0>
0C
#777010000000
1!
1*
b10 6
19
1>
1C
b10 G
#777020000000
0!
0*
09
0>
0C
#777030000000
1!
1*
b11 6
19
1>
1C
b11 G
#777040000000
0!
0*
09
0>
0C
#777050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#777060000000
0!
0*
09
0>
0C
#777070000000
1!
1*
b101 6
19
1>
1C
b101 G
#777080000000
0!
0*
09
0>
0C
#777090000000
1!
1*
b110 6
19
1>
1C
b110 G
#777100000000
0!
0*
09
0>
0C
#777110000000
1!
1*
b111 6
19
1>
1C
b111 G
#777120000000
0!
0*
09
0>
0C
#777130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#777140000000
0!
0*
09
0>
0C
#777150000000
1!
1*
b1 6
19
1>
1C
b1 G
#777160000000
0!
0*
09
0>
0C
#777170000000
1!
1*
b10 6
19
1>
1C
b10 G
#777180000000
0!
0*
09
0>
0C
#777190000000
1!
1*
b11 6
19
1>
1C
b11 G
#777200000000
0!
0*
09
0>
0C
#777210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#777220000000
0!
0*
09
0>
0C
#777230000000
1!
1*
b101 6
19
1>
1C
b101 G
#777240000000
0!
0*
09
0>
0C
#777250000000
1!
1*
b110 6
19
1>
1C
b110 G
#777260000000
0!
0*
09
0>
0C
#777270000000
1!
1*
b111 6
19
1>
1C
b111 G
#777280000000
0!
1"
0*
1+
09
1:
0>
0C
#777290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#777300000000
0!
0*
09
0>
0C
#777310000000
1!
1*
b1 6
19
1>
1C
b1 G
#777320000000
0!
0*
09
0>
0C
#777330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#777340000000
0!
0*
09
0>
0C
#777350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#777360000000
0!
0*
09
0>
0C
#777370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#777380000000
0!
0*
09
0>
0C
#777390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#777400000000
0!
0#
0*
0,
09
0>
0?
0C
#777410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#777420000000
0!
0*
09
0>
0C
#777430000000
1!
1*
19
1>
1C
#777440000000
0!
0*
09
0>
0C
#777450000000
1!
1*
19
1>
1C
#777460000000
0!
0*
09
0>
0C
#777470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#777480000000
0!
0*
09
0>
0C
#777490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#777500000000
0!
0*
09
0>
0C
#777510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#777520000000
0!
0*
09
0>
0C
#777530000000
1!
1*
b10 6
19
1>
1C
b10 G
#777540000000
0!
0*
09
0>
0C
#777550000000
1!
1*
b11 6
19
1>
1C
b11 G
#777560000000
0!
0*
09
0>
0C
#777570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#777580000000
0!
0*
09
0>
0C
#777590000000
1!
1*
b101 6
19
1>
1C
b101 G
#777600000000
0!
0*
09
0>
0C
#777610000000
1!
1*
b110 6
19
1>
1C
b110 G
#777620000000
0!
0*
09
0>
0C
#777630000000
1!
1*
b111 6
19
1>
1C
b111 G
#777640000000
0!
0*
09
0>
0C
#777650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#777660000000
0!
0*
09
0>
0C
#777670000000
1!
1*
b1 6
19
1>
1C
b1 G
#777680000000
0!
0*
09
0>
0C
#777690000000
1!
1*
b10 6
19
1>
1C
b10 G
#777700000000
0!
0*
09
0>
0C
#777710000000
1!
1*
b11 6
19
1>
1C
b11 G
#777720000000
0!
0*
09
0>
0C
#777730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#777740000000
0!
0*
09
0>
0C
#777750000000
1!
1*
b101 6
19
1>
1C
b101 G
#777760000000
0!
0*
09
0>
0C
#777770000000
1!
1*
b110 6
19
1>
1C
b110 G
#777780000000
0!
0*
09
0>
0C
#777790000000
1!
1*
b111 6
19
1>
1C
b111 G
#777800000000
0!
0*
09
0>
0C
#777810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#777820000000
0!
0*
09
0>
0C
#777830000000
1!
1*
b1 6
19
1>
1C
b1 G
#777840000000
0!
0*
09
0>
0C
#777850000000
1!
1*
b10 6
19
1>
1C
b10 G
#777860000000
0!
0*
09
0>
0C
#777870000000
1!
1*
b11 6
19
1>
1C
b11 G
#777880000000
0!
0*
09
0>
0C
#777890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#777900000000
0!
0*
09
0>
0C
#777910000000
1!
1*
b101 6
19
1>
1C
b101 G
#777920000000
0!
0*
09
0>
0C
#777930000000
1!
1*
b110 6
19
1>
1C
b110 G
#777940000000
0!
0*
09
0>
0C
#777950000000
1!
1*
b111 6
19
1>
1C
b111 G
#777960000000
0!
1"
0*
1+
09
1:
0>
0C
#777970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#777980000000
0!
0*
09
0>
0C
#777990000000
1!
1*
b1 6
19
1>
1C
b1 G
#778000000000
0!
0*
09
0>
0C
#778010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#778020000000
0!
0*
09
0>
0C
#778030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#778040000000
0!
0*
09
0>
0C
#778050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#778060000000
0!
0*
09
0>
0C
#778070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#778080000000
0!
0#
0*
0,
09
0>
0?
0C
#778090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#778100000000
0!
0*
09
0>
0C
#778110000000
1!
1*
19
1>
1C
#778120000000
0!
0*
09
0>
0C
#778130000000
1!
1*
19
1>
1C
#778140000000
0!
0*
09
0>
0C
#778150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#778160000000
0!
0*
09
0>
0C
#778170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#778180000000
0!
0*
09
0>
0C
#778190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#778200000000
0!
0*
09
0>
0C
#778210000000
1!
1*
b10 6
19
1>
1C
b10 G
#778220000000
0!
0*
09
0>
0C
#778230000000
1!
1*
b11 6
19
1>
1C
b11 G
#778240000000
0!
0*
09
0>
0C
#778250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#778260000000
0!
0*
09
0>
0C
#778270000000
1!
1*
b101 6
19
1>
1C
b101 G
#778280000000
0!
0*
09
0>
0C
#778290000000
1!
1*
b110 6
19
1>
1C
b110 G
#778300000000
0!
0*
09
0>
0C
#778310000000
1!
1*
b111 6
19
1>
1C
b111 G
#778320000000
0!
0*
09
0>
0C
#778330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#778340000000
0!
0*
09
0>
0C
#778350000000
1!
1*
b1 6
19
1>
1C
b1 G
#778360000000
0!
0*
09
0>
0C
#778370000000
1!
1*
b10 6
19
1>
1C
b10 G
#778380000000
0!
0*
09
0>
0C
#778390000000
1!
1*
b11 6
19
1>
1C
b11 G
#778400000000
0!
0*
09
0>
0C
#778410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#778420000000
0!
0*
09
0>
0C
#778430000000
1!
1*
b101 6
19
1>
1C
b101 G
#778440000000
0!
0*
09
0>
0C
#778450000000
1!
1*
b110 6
19
1>
1C
b110 G
#778460000000
0!
0*
09
0>
0C
#778470000000
1!
1*
b111 6
19
1>
1C
b111 G
#778480000000
0!
0*
09
0>
0C
#778490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#778500000000
0!
0*
09
0>
0C
#778510000000
1!
1*
b1 6
19
1>
1C
b1 G
#778520000000
0!
0*
09
0>
0C
#778530000000
1!
1*
b10 6
19
1>
1C
b10 G
#778540000000
0!
0*
09
0>
0C
#778550000000
1!
1*
b11 6
19
1>
1C
b11 G
#778560000000
0!
0*
09
0>
0C
#778570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#778580000000
0!
0*
09
0>
0C
#778590000000
1!
1*
b101 6
19
1>
1C
b101 G
#778600000000
0!
0*
09
0>
0C
#778610000000
1!
1*
b110 6
19
1>
1C
b110 G
#778620000000
0!
0*
09
0>
0C
#778630000000
1!
1*
b111 6
19
1>
1C
b111 G
#778640000000
0!
1"
0*
1+
09
1:
0>
0C
#778650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#778660000000
0!
0*
09
0>
0C
#778670000000
1!
1*
b1 6
19
1>
1C
b1 G
#778680000000
0!
0*
09
0>
0C
#778690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#778700000000
0!
0*
09
0>
0C
#778710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#778720000000
0!
0*
09
0>
0C
#778730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#778740000000
0!
0*
09
0>
0C
#778750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#778760000000
0!
0#
0*
0,
09
0>
0?
0C
#778770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#778780000000
0!
0*
09
0>
0C
#778790000000
1!
1*
19
1>
1C
#778800000000
0!
0*
09
0>
0C
#778810000000
1!
1*
19
1>
1C
#778820000000
0!
0*
09
0>
0C
#778830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#778840000000
0!
0*
09
0>
0C
#778850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#778860000000
0!
0*
09
0>
0C
#778870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#778880000000
0!
0*
09
0>
0C
#778890000000
1!
1*
b10 6
19
1>
1C
b10 G
#778900000000
0!
0*
09
0>
0C
#778910000000
1!
1*
b11 6
19
1>
1C
b11 G
#778920000000
0!
0*
09
0>
0C
#778930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#778940000000
0!
0*
09
0>
0C
#778950000000
1!
1*
b101 6
19
1>
1C
b101 G
#778960000000
0!
0*
09
0>
0C
#778970000000
1!
1*
b110 6
19
1>
1C
b110 G
#778980000000
0!
0*
09
0>
0C
#778990000000
1!
1*
b111 6
19
1>
1C
b111 G
#779000000000
0!
0*
09
0>
0C
#779010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#779020000000
0!
0*
09
0>
0C
#779030000000
1!
1*
b1 6
19
1>
1C
b1 G
#779040000000
0!
0*
09
0>
0C
#779050000000
1!
1*
b10 6
19
1>
1C
b10 G
#779060000000
0!
0*
09
0>
0C
#779070000000
1!
1*
b11 6
19
1>
1C
b11 G
#779080000000
0!
0*
09
0>
0C
#779090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#779100000000
0!
0*
09
0>
0C
#779110000000
1!
1*
b101 6
19
1>
1C
b101 G
#779120000000
0!
0*
09
0>
0C
#779130000000
1!
1*
b110 6
19
1>
1C
b110 G
#779140000000
0!
0*
09
0>
0C
#779150000000
1!
1*
b111 6
19
1>
1C
b111 G
#779160000000
0!
0*
09
0>
0C
#779170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#779180000000
0!
0*
09
0>
0C
#779190000000
1!
1*
b1 6
19
1>
1C
b1 G
#779200000000
0!
0*
09
0>
0C
#779210000000
1!
1*
b10 6
19
1>
1C
b10 G
#779220000000
0!
0*
09
0>
0C
#779230000000
1!
1*
b11 6
19
1>
1C
b11 G
#779240000000
0!
0*
09
0>
0C
#779250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#779260000000
0!
0*
09
0>
0C
#779270000000
1!
1*
b101 6
19
1>
1C
b101 G
#779280000000
0!
0*
09
0>
0C
#779290000000
1!
1*
b110 6
19
1>
1C
b110 G
#779300000000
0!
0*
09
0>
0C
#779310000000
1!
1*
b111 6
19
1>
1C
b111 G
#779320000000
0!
1"
0*
1+
09
1:
0>
0C
#779330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#779340000000
0!
0*
09
0>
0C
#779350000000
1!
1*
b1 6
19
1>
1C
b1 G
#779360000000
0!
0*
09
0>
0C
#779370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#779380000000
0!
0*
09
0>
0C
#779390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#779400000000
0!
0*
09
0>
0C
#779410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#779420000000
0!
0*
09
0>
0C
#779430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#779440000000
0!
0#
0*
0,
09
0>
0?
0C
#779450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#779460000000
0!
0*
09
0>
0C
#779470000000
1!
1*
19
1>
1C
#779480000000
0!
0*
09
0>
0C
#779490000000
1!
1*
19
1>
1C
#779500000000
0!
0*
09
0>
0C
#779510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#779520000000
0!
0*
09
0>
0C
#779530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#779540000000
0!
0*
09
0>
0C
#779550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#779560000000
0!
0*
09
0>
0C
#779570000000
1!
1*
b10 6
19
1>
1C
b10 G
#779580000000
0!
0*
09
0>
0C
#779590000000
1!
1*
b11 6
19
1>
1C
b11 G
#779600000000
0!
0*
09
0>
0C
#779610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#779620000000
0!
0*
09
0>
0C
#779630000000
1!
1*
b101 6
19
1>
1C
b101 G
#779640000000
0!
0*
09
0>
0C
#779650000000
1!
1*
b110 6
19
1>
1C
b110 G
#779660000000
0!
0*
09
0>
0C
#779670000000
1!
1*
b111 6
19
1>
1C
b111 G
#779680000000
0!
0*
09
0>
0C
#779690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#779700000000
0!
0*
09
0>
0C
#779710000000
1!
1*
b1 6
19
1>
1C
b1 G
#779720000000
0!
0*
09
0>
0C
#779730000000
1!
1*
b10 6
19
1>
1C
b10 G
#779740000000
0!
0*
09
0>
0C
#779750000000
1!
1*
b11 6
19
1>
1C
b11 G
#779760000000
0!
0*
09
0>
0C
#779770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#779780000000
0!
0*
09
0>
0C
#779790000000
1!
1*
b101 6
19
1>
1C
b101 G
#779800000000
0!
0*
09
0>
0C
#779810000000
1!
1*
b110 6
19
1>
1C
b110 G
#779820000000
0!
0*
09
0>
0C
#779830000000
1!
1*
b111 6
19
1>
1C
b111 G
#779840000000
0!
0*
09
0>
0C
#779850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#779860000000
0!
0*
09
0>
0C
#779870000000
1!
1*
b1 6
19
1>
1C
b1 G
#779880000000
0!
0*
09
0>
0C
#779890000000
1!
1*
b10 6
19
1>
1C
b10 G
#779900000000
0!
0*
09
0>
0C
#779910000000
1!
1*
b11 6
19
1>
1C
b11 G
#779920000000
0!
0*
09
0>
0C
#779930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#779940000000
0!
0*
09
0>
0C
#779950000000
1!
1*
b101 6
19
1>
1C
b101 G
#779960000000
0!
0*
09
0>
0C
#779970000000
1!
1*
b110 6
19
1>
1C
b110 G
#779980000000
0!
0*
09
0>
0C
#779990000000
1!
1*
b111 6
19
1>
1C
b111 G
#780000000000
0!
1"
0*
1+
09
1:
0>
0C
#780010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#780020000000
0!
0*
09
0>
0C
#780030000000
1!
1*
b1 6
19
1>
1C
b1 G
#780040000000
0!
0*
09
0>
0C
#780050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#780060000000
0!
0*
09
0>
0C
#780070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#780080000000
0!
0*
09
0>
0C
#780090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#780100000000
0!
0*
09
0>
0C
#780110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#780120000000
0!
0#
0*
0,
09
0>
0?
0C
#780130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#780140000000
0!
0*
09
0>
0C
#780150000000
1!
1*
19
1>
1C
#780160000000
0!
0*
09
0>
0C
#780170000000
1!
1*
19
1>
1C
#780180000000
0!
0*
09
0>
0C
#780190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#780200000000
0!
0*
09
0>
0C
#780210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#780220000000
0!
0*
09
0>
0C
#780230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#780240000000
0!
0*
09
0>
0C
#780250000000
1!
1*
b10 6
19
1>
1C
b10 G
#780260000000
0!
0*
09
0>
0C
#780270000000
1!
1*
b11 6
19
1>
1C
b11 G
#780280000000
0!
0*
09
0>
0C
#780290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#780300000000
0!
0*
09
0>
0C
#780310000000
1!
1*
b101 6
19
1>
1C
b101 G
#780320000000
0!
0*
09
0>
0C
#780330000000
1!
1*
b110 6
19
1>
1C
b110 G
#780340000000
0!
0*
09
0>
0C
#780350000000
1!
1*
b111 6
19
1>
1C
b111 G
#780360000000
0!
0*
09
0>
0C
#780370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#780380000000
0!
0*
09
0>
0C
#780390000000
1!
1*
b1 6
19
1>
1C
b1 G
#780400000000
0!
0*
09
0>
0C
#780410000000
1!
1*
b10 6
19
1>
1C
b10 G
#780420000000
0!
0*
09
0>
0C
#780430000000
1!
1*
b11 6
19
1>
1C
b11 G
#780440000000
0!
0*
09
0>
0C
#780450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#780460000000
0!
0*
09
0>
0C
#780470000000
1!
1*
b101 6
19
1>
1C
b101 G
#780480000000
0!
0*
09
0>
0C
#780490000000
1!
1*
b110 6
19
1>
1C
b110 G
#780500000000
0!
0*
09
0>
0C
#780510000000
1!
1*
b111 6
19
1>
1C
b111 G
#780520000000
0!
0*
09
0>
0C
#780530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#780540000000
0!
0*
09
0>
0C
#780550000000
1!
1*
b1 6
19
1>
1C
b1 G
#780560000000
0!
0*
09
0>
0C
#780570000000
1!
1*
b10 6
19
1>
1C
b10 G
#780580000000
0!
0*
09
0>
0C
#780590000000
1!
1*
b11 6
19
1>
1C
b11 G
#780600000000
0!
0*
09
0>
0C
#780610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#780620000000
0!
0*
09
0>
0C
#780630000000
1!
1*
b101 6
19
1>
1C
b101 G
#780640000000
0!
0*
09
0>
0C
#780650000000
1!
1*
b110 6
19
1>
1C
b110 G
#780660000000
0!
0*
09
0>
0C
#780670000000
1!
1*
b111 6
19
1>
1C
b111 G
#780680000000
0!
1"
0*
1+
09
1:
0>
0C
#780690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#780700000000
0!
0*
09
0>
0C
#780710000000
1!
1*
b1 6
19
1>
1C
b1 G
#780720000000
0!
0*
09
0>
0C
#780730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#780740000000
0!
0*
09
0>
0C
#780750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#780760000000
0!
0*
09
0>
0C
#780770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#780780000000
0!
0*
09
0>
0C
#780790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#780800000000
0!
0#
0*
0,
09
0>
0?
0C
#780810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#780820000000
0!
0*
09
0>
0C
#780830000000
1!
1*
19
1>
1C
#780840000000
0!
0*
09
0>
0C
#780850000000
1!
1*
19
1>
1C
#780860000000
0!
0*
09
0>
0C
#780870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#780880000000
0!
0*
09
0>
0C
#780890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#780900000000
0!
0*
09
0>
0C
#780910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#780920000000
0!
0*
09
0>
0C
#780930000000
1!
1*
b10 6
19
1>
1C
b10 G
#780940000000
0!
0*
09
0>
0C
#780950000000
1!
1*
b11 6
19
1>
1C
b11 G
#780960000000
0!
0*
09
0>
0C
#780970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#780980000000
0!
0*
09
0>
0C
#780990000000
1!
1*
b101 6
19
1>
1C
b101 G
#781000000000
0!
0*
09
0>
0C
#781010000000
1!
1*
b110 6
19
1>
1C
b110 G
#781020000000
0!
0*
09
0>
0C
#781030000000
1!
1*
b111 6
19
1>
1C
b111 G
#781040000000
0!
0*
09
0>
0C
#781050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#781060000000
0!
0*
09
0>
0C
#781070000000
1!
1*
b1 6
19
1>
1C
b1 G
#781080000000
0!
0*
09
0>
0C
#781090000000
1!
1*
b10 6
19
1>
1C
b10 G
#781100000000
0!
0*
09
0>
0C
#781110000000
1!
1*
b11 6
19
1>
1C
b11 G
#781120000000
0!
0*
09
0>
0C
#781130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#781140000000
0!
0*
09
0>
0C
#781150000000
1!
1*
b101 6
19
1>
1C
b101 G
#781160000000
0!
0*
09
0>
0C
#781170000000
1!
1*
b110 6
19
1>
1C
b110 G
#781180000000
0!
0*
09
0>
0C
#781190000000
1!
1*
b111 6
19
1>
1C
b111 G
#781200000000
0!
0*
09
0>
0C
#781210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#781220000000
0!
0*
09
0>
0C
#781230000000
1!
1*
b1 6
19
1>
1C
b1 G
#781240000000
0!
0*
09
0>
0C
#781250000000
1!
1*
b10 6
19
1>
1C
b10 G
#781260000000
0!
0*
09
0>
0C
#781270000000
1!
1*
b11 6
19
1>
1C
b11 G
#781280000000
0!
0*
09
0>
0C
#781290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#781300000000
0!
0*
09
0>
0C
#781310000000
1!
1*
b101 6
19
1>
1C
b101 G
#781320000000
0!
0*
09
0>
0C
#781330000000
1!
1*
b110 6
19
1>
1C
b110 G
#781340000000
0!
0*
09
0>
0C
#781350000000
1!
1*
b111 6
19
1>
1C
b111 G
#781360000000
0!
1"
0*
1+
09
1:
0>
0C
#781370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#781380000000
0!
0*
09
0>
0C
#781390000000
1!
1*
b1 6
19
1>
1C
b1 G
#781400000000
0!
0*
09
0>
0C
#781410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#781420000000
0!
0*
09
0>
0C
#781430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#781440000000
0!
0*
09
0>
0C
#781450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#781460000000
0!
0*
09
0>
0C
#781470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#781480000000
0!
0#
0*
0,
09
0>
0?
0C
#781490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#781500000000
0!
0*
09
0>
0C
#781510000000
1!
1*
19
1>
1C
#781520000000
0!
0*
09
0>
0C
#781530000000
1!
1*
19
1>
1C
#781540000000
0!
0*
09
0>
0C
#781550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#781560000000
0!
0*
09
0>
0C
#781570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#781580000000
0!
0*
09
0>
0C
#781590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#781600000000
0!
0*
09
0>
0C
#781610000000
1!
1*
b10 6
19
1>
1C
b10 G
#781620000000
0!
0*
09
0>
0C
#781630000000
1!
1*
b11 6
19
1>
1C
b11 G
#781640000000
0!
0*
09
0>
0C
#781650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#781660000000
0!
0*
09
0>
0C
#781670000000
1!
1*
b101 6
19
1>
1C
b101 G
#781680000000
0!
0*
09
0>
0C
#781690000000
1!
1*
b110 6
19
1>
1C
b110 G
#781700000000
0!
0*
09
0>
0C
#781710000000
1!
1*
b111 6
19
1>
1C
b111 G
#781720000000
0!
0*
09
0>
0C
#781730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#781740000000
0!
0*
09
0>
0C
#781750000000
1!
1*
b1 6
19
1>
1C
b1 G
#781760000000
0!
0*
09
0>
0C
#781770000000
1!
1*
b10 6
19
1>
1C
b10 G
#781780000000
0!
0*
09
0>
0C
#781790000000
1!
1*
b11 6
19
1>
1C
b11 G
#781800000000
0!
0*
09
0>
0C
#781810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#781820000000
0!
0*
09
0>
0C
#781830000000
1!
1*
b101 6
19
1>
1C
b101 G
#781840000000
0!
0*
09
0>
0C
#781850000000
1!
1*
b110 6
19
1>
1C
b110 G
#781860000000
0!
0*
09
0>
0C
#781870000000
1!
1*
b111 6
19
1>
1C
b111 G
#781880000000
0!
0*
09
0>
0C
#781890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#781900000000
0!
0*
09
0>
0C
#781910000000
1!
1*
b1 6
19
1>
1C
b1 G
#781920000000
0!
0*
09
0>
0C
#781930000000
1!
1*
b10 6
19
1>
1C
b10 G
#781940000000
0!
0*
09
0>
0C
#781950000000
1!
1*
b11 6
19
1>
1C
b11 G
#781960000000
0!
0*
09
0>
0C
#781970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#781980000000
0!
0*
09
0>
0C
#781990000000
1!
1*
b101 6
19
1>
1C
b101 G
#782000000000
0!
0*
09
0>
0C
#782010000000
1!
1*
b110 6
19
1>
1C
b110 G
#782020000000
0!
0*
09
0>
0C
#782030000000
1!
1*
b111 6
19
1>
1C
b111 G
#782040000000
0!
1"
0*
1+
09
1:
0>
0C
#782050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#782060000000
0!
0*
09
0>
0C
#782070000000
1!
1*
b1 6
19
1>
1C
b1 G
#782080000000
0!
0*
09
0>
0C
#782090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#782100000000
0!
0*
09
0>
0C
#782110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#782120000000
0!
0*
09
0>
0C
#782130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#782140000000
0!
0*
09
0>
0C
#782150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#782160000000
0!
0#
0*
0,
09
0>
0?
0C
#782170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#782180000000
0!
0*
09
0>
0C
#782190000000
1!
1*
19
1>
1C
#782200000000
0!
0*
09
0>
0C
#782210000000
1!
1*
19
1>
1C
#782220000000
0!
0*
09
0>
0C
#782230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#782240000000
0!
0*
09
0>
0C
#782250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#782260000000
0!
0*
09
0>
0C
#782270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#782280000000
0!
0*
09
0>
0C
#782290000000
1!
1*
b10 6
19
1>
1C
b10 G
#782300000000
0!
0*
09
0>
0C
#782310000000
1!
1*
b11 6
19
1>
1C
b11 G
#782320000000
0!
0*
09
0>
0C
#782330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#782340000000
0!
0*
09
0>
0C
#782350000000
1!
1*
b101 6
19
1>
1C
b101 G
#782360000000
0!
0*
09
0>
0C
#782370000000
1!
1*
b110 6
19
1>
1C
b110 G
#782380000000
0!
0*
09
0>
0C
#782390000000
1!
1*
b111 6
19
1>
1C
b111 G
#782400000000
0!
0*
09
0>
0C
#782410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#782420000000
0!
0*
09
0>
0C
#782430000000
1!
1*
b1 6
19
1>
1C
b1 G
#782440000000
0!
0*
09
0>
0C
#782450000000
1!
1*
b10 6
19
1>
1C
b10 G
#782460000000
0!
0*
09
0>
0C
#782470000000
1!
1*
b11 6
19
1>
1C
b11 G
#782480000000
0!
0*
09
0>
0C
#782490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#782500000000
0!
0*
09
0>
0C
#782510000000
1!
1*
b101 6
19
1>
1C
b101 G
#782520000000
0!
0*
09
0>
0C
#782530000000
1!
1*
b110 6
19
1>
1C
b110 G
#782540000000
0!
0*
09
0>
0C
#782550000000
1!
1*
b111 6
19
1>
1C
b111 G
#782560000000
0!
0*
09
0>
0C
#782570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#782580000000
0!
0*
09
0>
0C
#782590000000
1!
1*
b1 6
19
1>
1C
b1 G
#782600000000
0!
0*
09
0>
0C
#782610000000
1!
1*
b10 6
19
1>
1C
b10 G
#782620000000
0!
0*
09
0>
0C
#782630000000
1!
1*
b11 6
19
1>
1C
b11 G
#782640000000
0!
0*
09
0>
0C
#782650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#782660000000
0!
0*
09
0>
0C
#782670000000
1!
1*
b101 6
19
1>
1C
b101 G
#782680000000
0!
0*
09
0>
0C
#782690000000
1!
1*
b110 6
19
1>
1C
b110 G
#782700000000
0!
0*
09
0>
0C
#782710000000
1!
1*
b111 6
19
1>
1C
b111 G
#782720000000
0!
1"
0*
1+
09
1:
0>
0C
#782730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#782740000000
0!
0*
09
0>
0C
#782750000000
1!
1*
b1 6
19
1>
1C
b1 G
#782760000000
0!
0*
09
0>
0C
#782770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#782780000000
0!
0*
09
0>
0C
#782790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#782800000000
0!
0*
09
0>
0C
#782810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#782820000000
0!
0*
09
0>
0C
#782830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#782840000000
0!
0#
0*
0,
09
0>
0?
0C
#782850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#782860000000
0!
0*
09
0>
0C
#782870000000
1!
1*
19
1>
1C
#782880000000
0!
0*
09
0>
0C
#782890000000
1!
1*
19
1>
1C
#782900000000
0!
0*
09
0>
0C
#782910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#782920000000
0!
0*
09
0>
0C
#782930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#782940000000
0!
0*
09
0>
0C
#782950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#782960000000
0!
0*
09
0>
0C
#782970000000
1!
1*
b10 6
19
1>
1C
b10 G
#782980000000
0!
0*
09
0>
0C
#782990000000
1!
1*
b11 6
19
1>
1C
b11 G
#783000000000
0!
0*
09
0>
0C
#783010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#783020000000
0!
0*
09
0>
0C
#783030000000
1!
1*
b101 6
19
1>
1C
b101 G
#783040000000
0!
0*
09
0>
0C
#783050000000
1!
1*
b110 6
19
1>
1C
b110 G
#783060000000
0!
0*
09
0>
0C
#783070000000
1!
1*
b111 6
19
1>
1C
b111 G
#783080000000
0!
0*
09
0>
0C
#783090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#783100000000
0!
0*
09
0>
0C
#783110000000
1!
1*
b1 6
19
1>
1C
b1 G
#783120000000
0!
0*
09
0>
0C
#783130000000
1!
1*
b10 6
19
1>
1C
b10 G
#783140000000
0!
0*
09
0>
0C
#783150000000
1!
1*
b11 6
19
1>
1C
b11 G
#783160000000
0!
0*
09
0>
0C
#783170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#783180000000
0!
0*
09
0>
0C
#783190000000
1!
1*
b101 6
19
1>
1C
b101 G
#783200000000
0!
0*
09
0>
0C
#783210000000
1!
1*
b110 6
19
1>
1C
b110 G
#783220000000
0!
0*
09
0>
0C
#783230000000
1!
1*
b111 6
19
1>
1C
b111 G
#783240000000
0!
0*
09
0>
0C
#783250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#783260000000
0!
0*
09
0>
0C
#783270000000
1!
1*
b1 6
19
1>
1C
b1 G
#783280000000
0!
0*
09
0>
0C
#783290000000
1!
1*
b10 6
19
1>
1C
b10 G
#783300000000
0!
0*
09
0>
0C
#783310000000
1!
1*
b11 6
19
1>
1C
b11 G
#783320000000
0!
0*
09
0>
0C
#783330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#783340000000
0!
0*
09
0>
0C
#783350000000
1!
1*
b101 6
19
1>
1C
b101 G
#783360000000
0!
0*
09
0>
0C
#783370000000
1!
1*
b110 6
19
1>
1C
b110 G
#783380000000
0!
0*
09
0>
0C
#783390000000
1!
1*
b111 6
19
1>
1C
b111 G
#783400000000
0!
1"
0*
1+
09
1:
0>
0C
#783410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#783420000000
0!
0*
09
0>
0C
#783430000000
1!
1*
b1 6
19
1>
1C
b1 G
#783440000000
0!
0*
09
0>
0C
#783450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#783460000000
0!
0*
09
0>
0C
#783470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#783480000000
0!
0*
09
0>
0C
#783490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#783500000000
0!
0*
09
0>
0C
#783510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#783520000000
0!
0#
0*
0,
09
0>
0?
0C
#783530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#783540000000
0!
0*
09
0>
0C
#783550000000
1!
1*
19
1>
1C
#783560000000
0!
0*
09
0>
0C
#783570000000
1!
1*
19
1>
1C
#783580000000
0!
0*
09
0>
0C
#783590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#783600000000
0!
0*
09
0>
0C
#783610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#783620000000
0!
0*
09
0>
0C
#783630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#783640000000
0!
0*
09
0>
0C
#783650000000
1!
1*
b10 6
19
1>
1C
b10 G
#783660000000
0!
0*
09
0>
0C
#783670000000
1!
1*
b11 6
19
1>
1C
b11 G
#783680000000
0!
0*
09
0>
0C
#783690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#783700000000
0!
0*
09
0>
0C
#783710000000
1!
1*
b101 6
19
1>
1C
b101 G
#783720000000
0!
0*
09
0>
0C
#783730000000
1!
1*
b110 6
19
1>
1C
b110 G
#783740000000
0!
0*
09
0>
0C
#783750000000
1!
1*
b111 6
19
1>
1C
b111 G
#783760000000
0!
0*
09
0>
0C
#783770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#783780000000
0!
0*
09
0>
0C
#783790000000
1!
1*
b1 6
19
1>
1C
b1 G
#783800000000
0!
0*
09
0>
0C
#783810000000
1!
1*
b10 6
19
1>
1C
b10 G
#783820000000
0!
0*
09
0>
0C
#783830000000
1!
1*
b11 6
19
1>
1C
b11 G
#783840000000
0!
0*
09
0>
0C
#783850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#783860000000
0!
0*
09
0>
0C
#783870000000
1!
1*
b101 6
19
1>
1C
b101 G
#783880000000
0!
0*
09
0>
0C
#783890000000
1!
1*
b110 6
19
1>
1C
b110 G
#783900000000
0!
0*
09
0>
0C
#783910000000
1!
1*
b111 6
19
1>
1C
b111 G
#783920000000
0!
0*
09
0>
0C
#783930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#783940000000
0!
0*
09
0>
0C
#783950000000
1!
1*
b1 6
19
1>
1C
b1 G
#783960000000
0!
0*
09
0>
0C
#783970000000
1!
1*
b10 6
19
1>
1C
b10 G
#783980000000
0!
0*
09
0>
0C
#783990000000
1!
1*
b11 6
19
1>
1C
b11 G
#784000000000
0!
0*
09
0>
0C
#784010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#784020000000
0!
0*
09
0>
0C
#784030000000
1!
1*
b101 6
19
1>
1C
b101 G
#784040000000
0!
0*
09
0>
0C
#784050000000
1!
1*
b110 6
19
1>
1C
b110 G
#784060000000
0!
0*
09
0>
0C
#784070000000
1!
1*
b111 6
19
1>
1C
b111 G
#784080000000
0!
1"
0*
1+
09
1:
0>
0C
#784090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#784100000000
0!
0*
09
0>
0C
#784110000000
1!
1*
b1 6
19
1>
1C
b1 G
#784120000000
0!
0*
09
0>
0C
#784130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#784140000000
0!
0*
09
0>
0C
#784150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#784160000000
0!
0*
09
0>
0C
#784170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#784180000000
0!
0*
09
0>
0C
#784190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#784200000000
0!
0#
0*
0,
09
0>
0?
0C
#784210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#784220000000
0!
0*
09
0>
0C
#784230000000
1!
1*
19
1>
1C
#784240000000
0!
0*
09
0>
0C
#784250000000
1!
1*
19
1>
1C
#784260000000
0!
0*
09
0>
0C
#784270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#784280000000
0!
0*
09
0>
0C
#784290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#784300000000
0!
0*
09
0>
0C
#784310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#784320000000
0!
0*
09
0>
0C
#784330000000
1!
1*
b10 6
19
1>
1C
b10 G
#784340000000
0!
0*
09
0>
0C
#784350000000
1!
1*
b11 6
19
1>
1C
b11 G
#784360000000
0!
0*
09
0>
0C
#784370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#784380000000
0!
0*
09
0>
0C
#784390000000
1!
1*
b101 6
19
1>
1C
b101 G
#784400000000
0!
0*
09
0>
0C
#784410000000
1!
1*
b110 6
19
1>
1C
b110 G
#784420000000
0!
0*
09
0>
0C
#784430000000
1!
1*
b111 6
19
1>
1C
b111 G
#784440000000
0!
0*
09
0>
0C
#784450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#784460000000
0!
0*
09
0>
0C
#784470000000
1!
1*
b1 6
19
1>
1C
b1 G
#784480000000
0!
0*
09
0>
0C
#784490000000
1!
1*
b10 6
19
1>
1C
b10 G
#784500000000
0!
0*
09
0>
0C
#784510000000
1!
1*
b11 6
19
1>
1C
b11 G
#784520000000
0!
0*
09
0>
0C
#784530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#784540000000
0!
0*
09
0>
0C
#784550000000
1!
1*
b101 6
19
1>
1C
b101 G
#784560000000
0!
0*
09
0>
0C
#784570000000
1!
1*
b110 6
19
1>
1C
b110 G
#784580000000
0!
0*
09
0>
0C
#784590000000
1!
1*
b111 6
19
1>
1C
b111 G
#784600000000
0!
0*
09
0>
0C
#784610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#784620000000
0!
0*
09
0>
0C
#784630000000
1!
1*
b1 6
19
1>
1C
b1 G
#784640000000
0!
0*
09
0>
0C
#784650000000
1!
1*
b10 6
19
1>
1C
b10 G
#784660000000
0!
0*
09
0>
0C
#784670000000
1!
1*
b11 6
19
1>
1C
b11 G
#784680000000
0!
0*
09
0>
0C
#784690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#784700000000
0!
0*
09
0>
0C
#784710000000
1!
1*
b101 6
19
1>
1C
b101 G
#784720000000
0!
0*
09
0>
0C
#784730000000
1!
1*
b110 6
19
1>
1C
b110 G
#784740000000
0!
0*
09
0>
0C
#784750000000
1!
1*
b111 6
19
1>
1C
b111 G
#784760000000
0!
1"
0*
1+
09
1:
0>
0C
#784770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#784780000000
0!
0*
09
0>
0C
#784790000000
1!
1*
b1 6
19
1>
1C
b1 G
#784800000000
0!
0*
09
0>
0C
#784810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#784820000000
0!
0*
09
0>
0C
#784830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#784840000000
0!
0*
09
0>
0C
#784850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#784860000000
0!
0*
09
0>
0C
#784870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#784880000000
0!
0#
0*
0,
09
0>
0?
0C
#784890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#784900000000
0!
0*
09
0>
0C
#784910000000
1!
1*
19
1>
1C
#784920000000
0!
0*
09
0>
0C
#784930000000
1!
1*
19
1>
1C
#784940000000
0!
0*
09
0>
0C
#784950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#784960000000
0!
0*
09
0>
0C
#784970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#784980000000
0!
0*
09
0>
0C
#784990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#785000000000
0!
0*
09
0>
0C
#785010000000
1!
1*
b10 6
19
1>
1C
b10 G
#785020000000
0!
0*
09
0>
0C
#785030000000
1!
1*
b11 6
19
1>
1C
b11 G
#785040000000
0!
0*
09
0>
0C
#785050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#785060000000
0!
0*
09
0>
0C
#785070000000
1!
1*
b101 6
19
1>
1C
b101 G
#785080000000
0!
0*
09
0>
0C
#785090000000
1!
1*
b110 6
19
1>
1C
b110 G
#785100000000
0!
0*
09
0>
0C
#785110000000
1!
1*
b111 6
19
1>
1C
b111 G
#785120000000
0!
0*
09
0>
0C
#785130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#785140000000
0!
0*
09
0>
0C
#785150000000
1!
1*
b1 6
19
1>
1C
b1 G
#785160000000
0!
0*
09
0>
0C
#785170000000
1!
1*
b10 6
19
1>
1C
b10 G
#785180000000
0!
0*
09
0>
0C
#785190000000
1!
1*
b11 6
19
1>
1C
b11 G
#785200000000
0!
0*
09
0>
0C
#785210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#785220000000
0!
0*
09
0>
0C
#785230000000
1!
1*
b101 6
19
1>
1C
b101 G
#785240000000
0!
0*
09
0>
0C
#785250000000
1!
1*
b110 6
19
1>
1C
b110 G
#785260000000
0!
0*
09
0>
0C
#785270000000
1!
1*
b111 6
19
1>
1C
b111 G
#785280000000
0!
0*
09
0>
0C
#785290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#785300000000
0!
0*
09
0>
0C
#785310000000
1!
1*
b1 6
19
1>
1C
b1 G
#785320000000
0!
0*
09
0>
0C
#785330000000
1!
1*
b10 6
19
1>
1C
b10 G
#785340000000
0!
0*
09
0>
0C
#785350000000
1!
1*
b11 6
19
1>
1C
b11 G
#785360000000
0!
0*
09
0>
0C
#785370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#785380000000
0!
0*
09
0>
0C
#785390000000
1!
1*
b101 6
19
1>
1C
b101 G
#785400000000
0!
0*
09
0>
0C
#785410000000
1!
1*
b110 6
19
1>
1C
b110 G
#785420000000
0!
0*
09
0>
0C
#785430000000
1!
1*
b111 6
19
1>
1C
b111 G
#785440000000
0!
1"
0*
1+
09
1:
0>
0C
#785450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#785460000000
0!
0*
09
0>
0C
#785470000000
1!
1*
b1 6
19
1>
1C
b1 G
#785480000000
0!
0*
09
0>
0C
#785490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#785500000000
0!
0*
09
0>
0C
#785510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#785520000000
0!
0*
09
0>
0C
#785530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#785540000000
0!
0*
09
0>
0C
#785550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#785560000000
0!
0#
0*
0,
09
0>
0?
0C
#785570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#785580000000
0!
0*
09
0>
0C
#785590000000
1!
1*
19
1>
1C
#785600000000
0!
0*
09
0>
0C
#785610000000
1!
1*
19
1>
1C
#785620000000
0!
0*
09
0>
0C
#785630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#785640000000
0!
0*
09
0>
0C
#785650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#785660000000
0!
0*
09
0>
0C
#785670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#785680000000
0!
0*
09
0>
0C
#785690000000
1!
1*
b10 6
19
1>
1C
b10 G
#785700000000
0!
0*
09
0>
0C
#785710000000
1!
1*
b11 6
19
1>
1C
b11 G
#785720000000
0!
0*
09
0>
0C
#785730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#785740000000
0!
0*
09
0>
0C
#785750000000
1!
1*
b101 6
19
1>
1C
b101 G
#785760000000
0!
0*
09
0>
0C
#785770000000
1!
1*
b110 6
19
1>
1C
b110 G
#785780000000
0!
0*
09
0>
0C
#785790000000
1!
1*
b111 6
19
1>
1C
b111 G
#785800000000
0!
0*
09
0>
0C
#785810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#785820000000
0!
0*
09
0>
0C
#785830000000
1!
1*
b1 6
19
1>
1C
b1 G
#785840000000
0!
0*
09
0>
0C
#785850000000
1!
1*
b10 6
19
1>
1C
b10 G
#785860000000
0!
0*
09
0>
0C
#785870000000
1!
1*
b11 6
19
1>
1C
b11 G
#785880000000
0!
0*
09
0>
0C
#785890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#785900000000
0!
0*
09
0>
0C
#785910000000
1!
1*
b101 6
19
1>
1C
b101 G
#785920000000
0!
0*
09
0>
0C
#785930000000
1!
1*
b110 6
19
1>
1C
b110 G
#785940000000
0!
0*
09
0>
0C
#785950000000
1!
1*
b111 6
19
1>
1C
b111 G
#785960000000
0!
0*
09
0>
0C
#785970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#785980000000
0!
0*
09
0>
0C
#785990000000
1!
1*
b1 6
19
1>
1C
b1 G
#786000000000
0!
0*
09
0>
0C
#786010000000
1!
1*
b10 6
19
1>
1C
b10 G
#786020000000
0!
0*
09
0>
0C
#786030000000
1!
1*
b11 6
19
1>
1C
b11 G
#786040000000
0!
0*
09
0>
0C
#786050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#786060000000
0!
0*
09
0>
0C
#786070000000
1!
1*
b101 6
19
1>
1C
b101 G
#786080000000
0!
0*
09
0>
0C
#786090000000
1!
1*
b110 6
19
1>
1C
b110 G
#786100000000
0!
0*
09
0>
0C
#786110000000
1!
1*
b111 6
19
1>
1C
b111 G
#786120000000
0!
1"
0*
1+
09
1:
0>
0C
#786130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#786140000000
0!
0*
09
0>
0C
#786150000000
1!
1*
b1 6
19
1>
1C
b1 G
#786160000000
0!
0*
09
0>
0C
#786170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#786180000000
0!
0*
09
0>
0C
#786190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#786200000000
0!
0*
09
0>
0C
#786210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#786220000000
0!
0*
09
0>
0C
#786230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#786240000000
0!
0#
0*
0,
09
0>
0?
0C
#786250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#786260000000
0!
0*
09
0>
0C
#786270000000
1!
1*
19
1>
1C
#786280000000
0!
0*
09
0>
0C
#786290000000
1!
1*
19
1>
1C
#786300000000
0!
0*
09
0>
0C
#786310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#786320000000
0!
0*
09
0>
0C
#786330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#786340000000
0!
0*
09
0>
0C
#786350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#786360000000
0!
0*
09
0>
0C
#786370000000
1!
1*
b10 6
19
1>
1C
b10 G
#786380000000
0!
0*
09
0>
0C
#786390000000
1!
1*
b11 6
19
1>
1C
b11 G
#786400000000
0!
0*
09
0>
0C
#786410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#786420000000
0!
0*
09
0>
0C
#786430000000
1!
1*
b101 6
19
1>
1C
b101 G
#786440000000
0!
0*
09
0>
0C
#786450000000
1!
1*
b110 6
19
1>
1C
b110 G
#786460000000
0!
0*
09
0>
0C
#786470000000
1!
1*
b111 6
19
1>
1C
b111 G
#786480000000
0!
0*
09
0>
0C
#786490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#786500000000
0!
0*
09
0>
0C
#786510000000
1!
1*
b1 6
19
1>
1C
b1 G
#786520000000
0!
0*
09
0>
0C
#786530000000
1!
1*
b10 6
19
1>
1C
b10 G
#786540000000
0!
0*
09
0>
0C
#786550000000
1!
1*
b11 6
19
1>
1C
b11 G
#786560000000
0!
0*
09
0>
0C
#786570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#786580000000
0!
0*
09
0>
0C
#786590000000
1!
1*
b101 6
19
1>
1C
b101 G
#786600000000
0!
0*
09
0>
0C
#786610000000
1!
1*
b110 6
19
1>
1C
b110 G
#786620000000
0!
0*
09
0>
0C
#786630000000
1!
1*
b111 6
19
1>
1C
b111 G
#786640000000
0!
0*
09
0>
0C
#786650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#786660000000
0!
0*
09
0>
0C
#786670000000
1!
1*
b1 6
19
1>
1C
b1 G
#786680000000
0!
0*
09
0>
0C
#786690000000
1!
1*
b10 6
19
1>
1C
b10 G
#786700000000
0!
0*
09
0>
0C
#786710000000
1!
1*
b11 6
19
1>
1C
b11 G
#786720000000
0!
0*
09
0>
0C
#786730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#786740000000
0!
0*
09
0>
0C
#786750000000
1!
1*
b101 6
19
1>
1C
b101 G
#786760000000
0!
0*
09
0>
0C
#786770000000
1!
1*
b110 6
19
1>
1C
b110 G
#786780000000
0!
0*
09
0>
0C
#786790000000
1!
1*
b111 6
19
1>
1C
b111 G
#786800000000
0!
1"
0*
1+
09
1:
0>
0C
#786810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#786820000000
0!
0*
09
0>
0C
#786830000000
1!
1*
b1 6
19
1>
1C
b1 G
#786840000000
0!
0*
09
0>
0C
#786850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#786860000000
0!
0*
09
0>
0C
#786870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#786880000000
0!
0*
09
0>
0C
#786890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#786900000000
0!
0*
09
0>
0C
#786910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#786920000000
0!
0#
0*
0,
09
0>
0?
0C
#786930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#786940000000
0!
0*
09
0>
0C
#786950000000
1!
1*
19
1>
1C
#786960000000
0!
0*
09
0>
0C
#786970000000
1!
1*
19
1>
1C
#786980000000
0!
0*
09
0>
0C
#786990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#787000000000
0!
0*
09
0>
0C
#787010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#787020000000
0!
0*
09
0>
0C
#787030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#787040000000
0!
0*
09
0>
0C
#787050000000
1!
1*
b10 6
19
1>
1C
b10 G
#787060000000
0!
0*
09
0>
0C
#787070000000
1!
1*
b11 6
19
1>
1C
b11 G
#787080000000
0!
0*
09
0>
0C
#787090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#787100000000
0!
0*
09
0>
0C
#787110000000
1!
1*
b101 6
19
1>
1C
b101 G
#787120000000
0!
0*
09
0>
0C
#787130000000
1!
1*
b110 6
19
1>
1C
b110 G
#787140000000
0!
0*
09
0>
0C
#787150000000
1!
1*
b111 6
19
1>
1C
b111 G
#787160000000
0!
0*
09
0>
0C
#787170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#787180000000
0!
0*
09
0>
0C
#787190000000
1!
1*
b1 6
19
1>
1C
b1 G
#787200000000
0!
0*
09
0>
0C
#787210000000
1!
1*
b10 6
19
1>
1C
b10 G
#787220000000
0!
0*
09
0>
0C
#787230000000
1!
1*
b11 6
19
1>
1C
b11 G
#787240000000
0!
0*
09
0>
0C
#787250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#787260000000
0!
0*
09
0>
0C
#787270000000
1!
1*
b101 6
19
1>
1C
b101 G
#787280000000
0!
0*
09
0>
0C
#787290000000
1!
1*
b110 6
19
1>
1C
b110 G
#787300000000
0!
0*
09
0>
0C
#787310000000
1!
1*
b111 6
19
1>
1C
b111 G
#787320000000
0!
0*
09
0>
0C
#787330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#787340000000
0!
0*
09
0>
0C
#787350000000
1!
1*
b1 6
19
1>
1C
b1 G
#787360000000
0!
0*
09
0>
0C
#787370000000
1!
1*
b10 6
19
1>
1C
b10 G
#787380000000
0!
0*
09
0>
0C
#787390000000
1!
1*
b11 6
19
1>
1C
b11 G
#787400000000
0!
0*
09
0>
0C
#787410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#787420000000
0!
0*
09
0>
0C
#787430000000
1!
1*
b101 6
19
1>
1C
b101 G
#787440000000
0!
0*
09
0>
0C
#787450000000
1!
1*
b110 6
19
1>
1C
b110 G
#787460000000
0!
0*
09
0>
0C
#787470000000
1!
1*
b111 6
19
1>
1C
b111 G
#787480000000
0!
1"
0*
1+
09
1:
0>
0C
#787490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#787500000000
0!
0*
09
0>
0C
#787510000000
1!
1*
b1 6
19
1>
1C
b1 G
#787520000000
0!
0*
09
0>
0C
#787530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#787540000000
0!
0*
09
0>
0C
#787550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#787560000000
0!
0*
09
0>
0C
#787570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#787580000000
0!
0*
09
0>
0C
#787590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#787600000000
0!
0#
0*
0,
09
0>
0?
0C
#787610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#787620000000
0!
0*
09
0>
0C
#787630000000
1!
1*
19
1>
1C
#787640000000
0!
0*
09
0>
0C
#787650000000
1!
1*
19
1>
1C
#787660000000
0!
0*
09
0>
0C
#787670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#787680000000
0!
0*
09
0>
0C
#787690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#787700000000
0!
0*
09
0>
0C
#787710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#787720000000
0!
0*
09
0>
0C
#787730000000
1!
1*
b10 6
19
1>
1C
b10 G
#787740000000
0!
0*
09
0>
0C
#787750000000
1!
1*
b11 6
19
1>
1C
b11 G
#787760000000
0!
0*
09
0>
0C
#787770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#787780000000
0!
0*
09
0>
0C
#787790000000
1!
1*
b101 6
19
1>
1C
b101 G
#787800000000
0!
0*
09
0>
0C
#787810000000
1!
1*
b110 6
19
1>
1C
b110 G
#787820000000
0!
0*
09
0>
0C
#787830000000
1!
1*
b111 6
19
1>
1C
b111 G
#787840000000
0!
0*
09
0>
0C
#787850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#787860000000
0!
0*
09
0>
0C
#787870000000
1!
1*
b1 6
19
1>
1C
b1 G
#787880000000
0!
0*
09
0>
0C
#787890000000
1!
1*
b10 6
19
1>
1C
b10 G
#787900000000
0!
0*
09
0>
0C
#787910000000
1!
1*
b11 6
19
1>
1C
b11 G
#787920000000
0!
0*
09
0>
0C
#787930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#787940000000
0!
0*
09
0>
0C
#787950000000
1!
1*
b101 6
19
1>
1C
b101 G
#787960000000
0!
0*
09
0>
0C
#787970000000
1!
1*
b110 6
19
1>
1C
b110 G
#787980000000
0!
0*
09
0>
0C
#787990000000
1!
1*
b111 6
19
1>
1C
b111 G
#788000000000
0!
0*
09
0>
0C
#788010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#788020000000
0!
0*
09
0>
0C
#788030000000
1!
1*
b1 6
19
1>
1C
b1 G
#788040000000
0!
0*
09
0>
0C
#788050000000
1!
1*
b10 6
19
1>
1C
b10 G
#788060000000
0!
0*
09
0>
0C
#788070000000
1!
1*
b11 6
19
1>
1C
b11 G
#788080000000
0!
0*
09
0>
0C
#788090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#788100000000
0!
0*
09
0>
0C
#788110000000
1!
1*
b101 6
19
1>
1C
b101 G
#788120000000
0!
0*
09
0>
0C
#788130000000
1!
1*
b110 6
19
1>
1C
b110 G
#788140000000
0!
0*
09
0>
0C
#788150000000
1!
1*
b111 6
19
1>
1C
b111 G
#788160000000
0!
1"
0*
1+
09
1:
0>
0C
#788170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#788180000000
0!
0*
09
0>
0C
#788190000000
1!
1*
b1 6
19
1>
1C
b1 G
#788200000000
0!
0*
09
0>
0C
#788210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#788220000000
0!
0*
09
0>
0C
#788230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#788240000000
0!
0*
09
0>
0C
#788250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#788260000000
0!
0*
09
0>
0C
#788270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#788280000000
0!
0#
0*
0,
09
0>
0?
0C
#788290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#788300000000
0!
0*
09
0>
0C
#788310000000
1!
1*
19
1>
1C
#788320000000
0!
0*
09
0>
0C
#788330000000
1!
1*
19
1>
1C
#788340000000
0!
0*
09
0>
0C
#788350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#788360000000
0!
0*
09
0>
0C
#788370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#788380000000
0!
0*
09
0>
0C
#788390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#788400000000
0!
0*
09
0>
0C
#788410000000
1!
1*
b10 6
19
1>
1C
b10 G
#788420000000
0!
0*
09
0>
0C
#788430000000
1!
1*
b11 6
19
1>
1C
b11 G
#788440000000
0!
0*
09
0>
0C
#788450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#788460000000
0!
0*
09
0>
0C
#788470000000
1!
1*
b101 6
19
1>
1C
b101 G
#788480000000
0!
0*
09
0>
0C
#788490000000
1!
1*
b110 6
19
1>
1C
b110 G
#788500000000
0!
0*
09
0>
0C
#788510000000
1!
1*
b111 6
19
1>
1C
b111 G
#788520000000
0!
0*
09
0>
0C
#788530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#788540000000
0!
0*
09
0>
0C
#788550000000
1!
1*
b1 6
19
1>
1C
b1 G
#788560000000
0!
0*
09
0>
0C
#788570000000
1!
1*
b10 6
19
1>
1C
b10 G
#788580000000
0!
0*
09
0>
0C
#788590000000
1!
1*
b11 6
19
1>
1C
b11 G
#788600000000
0!
0*
09
0>
0C
#788610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#788620000000
0!
0*
09
0>
0C
#788630000000
1!
1*
b101 6
19
1>
1C
b101 G
#788640000000
0!
0*
09
0>
0C
#788650000000
1!
1*
b110 6
19
1>
1C
b110 G
#788660000000
0!
0*
09
0>
0C
#788670000000
1!
1*
b111 6
19
1>
1C
b111 G
#788680000000
0!
0*
09
0>
0C
#788690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#788700000000
0!
0*
09
0>
0C
#788710000000
1!
1*
b1 6
19
1>
1C
b1 G
#788720000000
0!
0*
09
0>
0C
#788730000000
1!
1*
b10 6
19
1>
1C
b10 G
#788740000000
0!
0*
09
0>
0C
#788750000000
1!
1*
b11 6
19
1>
1C
b11 G
#788760000000
0!
0*
09
0>
0C
#788770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#788780000000
0!
0*
09
0>
0C
#788790000000
1!
1*
b101 6
19
1>
1C
b101 G
#788800000000
0!
0*
09
0>
0C
#788810000000
1!
1*
b110 6
19
1>
1C
b110 G
#788820000000
0!
0*
09
0>
0C
#788830000000
1!
1*
b111 6
19
1>
1C
b111 G
#788840000000
0!
1"
0*
1+
09
1:
0>
0C
#788850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#788860000000
0!
0*
09
0>
0C
#788870000000
1!
1*
b1 6
19
1>
1C
b1 G
#788880000000
0!
0*
09
0>
0C
#788890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#788900000000
0!
0*
09
0>
0C
#788910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#788920000000
0!
0*
09
0>
0C
#788930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#788940000000
0!
0*
09
0>
0C
#788950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#788960000000
0!
0#
0*
0,
09
0>
0?
0C
#788970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#788980000000
0!
0*
09
0>
0C
#788990000000
1!
1*
19
1>
1C
#789000000000
0!
0*
09
0>
0C
#789010000000
1!
1*
19
1>
1C
#789020000000
0!
0*
09
0>
0C
#789030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#789040000000
0!
0*
09
0>
0C
#789050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#789060000000
0!
0*
09
0>
0C
#789070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#789080000000
0!
0*
09
0>
0C
#789090000000
1!
1*
b10 6
19
1>
1C
b10 G
#789100000000
0!
0*
09
0>
0C
#789110000000
1!
1*
b11 6
19
1>
1C
b11 G
#789120000000
0!
0*
09
0>
0C
#789130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#789140000000
0!
0*
09
0>
0C
#789150000000
1!
1*
b101 6
19
1>
1C
b101 G
#789160000000
0!
0*
09
0>
0C
#789170000000
1!
1*
b110 6
19
1>
1C
b110 G
#789180000000
0!
0*
09
0>
0C
#789190000000
1!
1*
b111 6
19
1>
1C
b111 G
#789200000000
0!
0*
09
0>
0C
#789210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#789220000000
0!
0*
09
0>
0C
#789230000000
1!
1*
b1 6
19
1>
1C
b1 G
#789240000000
0!
0*
09
0>
0C
#789250000000
1!
1*
b10 6
19
1>
1C
b10 G
#789260000000
0!
0*
09
0>
0C
#789270000000
1!
1*
b11 6
19
1>
1C
b11 G
#789280000000
0!
0*
09
0>
0C
#789290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#789300000000
0!
0*
09
0>
0C
#789310000000
1!
1*
b101 6
19
1>
1C
b101 G
#789320000000
0!
0*
09
0>
0C
#789330000000
1!
1*
b110 6
19
1>
1C
b110 G
#789340000000
0!
0*
09
0>
0C
#789350000000
1!
1*
b111 6
19
1>
1C
b111 G
#789360000000
0!
0*
09
0>
0C
#789370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#789380000000
0!
0*
09
0>
0C
#789390000000
1!
1*
b1 6
19
1>
1C
b1 G
#789400000000
0!
0*
09
0>
0C
#789410000000
1!
1*
b10 6
19
1>
1C
b10 G
#789420000000
0!
0*
09
0>
0C
#789430000000
1!
1*
b11 6
19
1>
1C
b11 G
#789440000000
0!
0*
09
0>
0C
#789450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#789460000000
0!
0*
09
0>
0C
#789470000000
1!
1*
b101 6
19
1>
1C
b101 G
#789480000000
0!
0*
09
0>
0C
#789490000000
1!
1*
b110 6
19
1>
1C
b110 G
#789500000000
0!
0*
09
0>
0C
#789510000000
1!
1*
b111 6
19
1>
1C
b111 G
#789520000000
0!
1"
0*
1+
09
1:
0>
0C
#789530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#789540000000
0!
0*
09
0>
0C
#789550000000
1!
1*
b1 6
19
1>
1C
b1 G
#789560000000
0!
0*
09
0>
0C
#789570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#789580000000
0!
0*
09
0>
0C
#789590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#789600000000
0!
0*
09
0>
0C
#789610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#789620000000
0!
0*
09
0>
0C
#789630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#789640000000
0!
0#
0*
0,
09
0>
0?
0C
#789650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#789660000000
0!
0*
09
0>
0C
#789670000000
1!
1*
19
1>
1C
#789680000000
0!
0*
09
0>
0C
#789690000000
1!
1*
19
1>
1C
#789700000000
0!
0*
09
0>
0C
#789710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#789720000000
0!
0*
09
0>
0C
#789730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#789740000000
0!
0*
09
0>
0C
#789750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#789760000000
0!
0*
09
0>
0C
#789770000000
1!
1*
b10 6
19
1>
1C
b10 G
#789780000000
0!
0*
09
0>
0C
#789790000000
1!
1*
b11 6
19
1>
1C
b11 G
#789800000000
0!
0*
09
0>
0C
#789810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#789820000000
0!
0*
09
0>
0C
#789830000000
1!
1*
b101 6
19
1>
1C
b101 G
#789840000000
0!
0*
09
0>
0C
#789850000000
1!
1*
b110 6
19
1>
1C
b110 G
#789860000000
0!
0*
09
0>
0C
#789870000000
1!
1*
b111 6
19
1>
1C
b111 G
#789880000000
0!
0*
09
0>
0C
#789890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#789900000000
0!
0*
09
0>
0C
#789910000000
1!
1*
b1 6
19
1>
1C
b1 G
#789920000000
0!
0*
09
0>
0C
#789930000000
1!
1*
b10 6
19
1>
1C
b10 G
#789940000000
0!
0*
09
0>
0C
#789950000000
1!
1*
b11 6
19
1>
1C
b11 G
#789960000000
0!
0*
09
0>
0C
#789970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#789980000000
0!
0*
09
0>
0C
#789990000000
1!
1*
b101 6
19
1>
1C
b101 G
#790000000000
0!
0*
09
0>
0C
#790010000000
1!
1*
b110 6
19
1>
1C
b110 G
#790020000000
0!
0*
09
0>
0C
#790030000000
1!
1*
b111 6
19
1>
1C
b111 G
#790040000000
0!
0*
09
0>
0C
#790050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#790060000000
0!
0*
09
0>
0C
#790070000000
1!
1*
b1 6
19
1>
1C
b1 G
#790080000000
0!
0*
09
0>
0C
#790090000000
1!
1*
b10 6
19
1>
1C
b10 G
#790100000000
0!
0*
09
0>
0C
#790110000000
1!
1*
b11 6
19
1>
1C
b11 G
#790120000000
0!
0*
09
0>
0C
#790130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#790140000000
0!
0*
09
0>
0C
#790150000000
1!
1*
b101 6
19
1>
1C
b101 G
#790160000000
0!
0*
09
0>
0C
#790170000000
1!
1*
b110 6
19
1>
1C
b110 G
#790180000000
0!
0*
09
0>
0C
#790190000000
1!
1*
b111 6
19
1>
1C
b111 G
#790200000000
0!
1"
0*
1+
09
1:
0>
0C
#790210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#790220000000
0!
0*
09
0>
0C
#790230000000
1!
1*
b1 6
19
1>
1C
b1 G
#790240000000
0!
0*
09
0>
0C
#790250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#790260000000
0!
0*
09
0>
0C
#790270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#790280000000
0!
0*
09
0>
0C
#790290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#790300000000
0!
0*
09
0>
0C
#790310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#790320000000
0!
0#
0*
0,
09
0>
0?
0C
#790330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#790340000000
0!
0*
09
0>
0C
#790350000000
1!
1*
19
1>
1C
#790360000000
0!
0*
09
0>
0C
#790370000000
1!
1*
19
1>
1C
#790380000000
0!
0*
09
0>
0C
#790390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#790400000000
0!
0*
09
0>
0C
#790410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#790420000000
0!
0*
09
0>
0C
#790430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#790440000000
0!
0*
09
0>
0C
#790450000000
1!
1*
b10 6
19
1>
1C
b10 G
#790460000000
0!
0*
09
0>
0C
#790470000000
1!
1*
b11 6
19
1>
1C
b11 G
#790480000000
0!
0*
09
0>
0C
#790490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#790500000000
0!
0*
09
0>
0C
#790510000000
1!
1*
b101 6
19
1>
1C
b101 G
#790520000000
0!
0*
09
0>
0C
#790530000000
1!
1*
b110 6
19
1>
1C
b110 G
#790540000000
0!
0*
09
0>
0C
#790550000000
1!
1*
b111 6
19
1>
1C
b111 G
#790560000000
0!
0*
09
0>
0C
#790570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#790580000000
0!
0*
09
0>
0C
#790590000000
1!
1*
b1 6
19
1>
1C
b1 G
#790600000000
0!
0*
09
0>
0C
#790610000000
1!
1*
b10 6
19
1>
1C
b10 G
#790620000000
0!
0*
09
0>
0C
#790630000000
1!
1*
b11 6
19
1>
1C
b11 G
#790640000000
0!
0*
09
0>
0C
#790650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#790660000000
0!
0*
09
0>
0C
#790670000000
1!
1*
b101 6
19
1>
1C
b101 G
#790680000000
0!
0*
09
0>
0C
#790690000000
1!
1*
b110 6
19
1>
1C
b110 G
#790700000000
0!
0*
09
0>
0C
#790710000000
1!
1*
b111 6
19
1>
1C
b111 G
#790720000000
0!
0*
09
0>
0C
#790730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#790740000000
0!
0*
09
0>
0C
#790750000000
1!
1*
b1 6
19
1>
1C
b1 G
#790760000000
0!
0*
09
0>
0C
#790770000000
1!
1*
b10 6
19
1>
1C
b10 G
#790780000000
0!
0*
09
0>
0C
#790790000000
1!
1*
b11 6
19
1>
1C
b11 G
#790800000000
0!
0*
09
0>
0C
#790810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#790820000000
0!
0*
09
0>
0C
#790830000000
1!
1*
b101 6
19
1>
1C
b101 G
#790840000000
0!
0*
09
0>
0C
#790850000000
1!
1*
b110 6
19
1>
1C
b110 G
#790860000000
0!
0*
09
0>
0C
#790870000000
1!
1*
b111 6
19
1>
1C
b111 G
#790880000000
0!
1"
0*
1+
09
1:
0>
0C
#790890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#790900000000
0!
0*
09
0>
0C
#790910000000
1!
1*
b1 6
19
1>
1C
b1 G
#790920000000
0!
0*
09
0>
0C
#790930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#790940000000
0!
0*
09
0>
0C
#790950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#790960000000
0!
0*
09
0>
0C
#790970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#790980000000
0!
0*
09
0>
0C
#790990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#791000000000
0!
0#
0*
0,
09
0>
0?
0C
#791010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#791020000000
0!
0*
09
0>
0C
#791030000000
1!
1*
19
1>
1C
#791040000000
0!
0*
09
0>
0C
#791050000000
1!
1*
19
1>
1C
#791060000000
0!
0*
09
0>
0C
#791070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#791080000000
0!
0*
09
0>
0C
#791090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#791100000000
0!
0*
09
0>
0C
#791110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#791120000000
0!
0*
09
0>
0C
#791130000000
1!
1*
b10 6
19
1>
1C
b10 G
#791140000000
0!
0*
09
0>
0C
#791150000000
1!
1*
b11 6
19
1>
1C
b11 G
#791160000000
0!
0*
09
0>
0C
#791170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#791180000000
0!
0*
09
0>
0C
#791190000000
1!
1*
b101 6
19
1>
1C
b101 G
#791200000000
0!
0*
09
0>
0C
#791210000000
1!
1*
b110 6
19
1>
1C
b110 G
#791220000000
0!
0*
09
0>
0C
#791230000000
1!
1*
b111 6
19
1>
1C
b111 G
#791240000000
0!
0*
09
0>
0C
#791250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#791260000000
0!
0*
09
0>
0C
#791270000000
1!
1*
b1 6
19
1>
1C
b1 G
#791280000000
0!
0*
09
0>
0C
#791290000000
1!
1*
b10 6
19
1>
1C
b10 G
#791300000000
0!
0*
09
0>
0C
#791310000000
1!
1*
b11 6
19
1>
1C
b11 G
#791320000000
0!
0*
09
0>
0C
#791330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#791340000000
0!
0*
09
0>
0C
#791350000000
1!
1*
b101 6
19
1>
1C
b101 G
#791360000000
0!
0*
09
0>
0C
#791370000000
1!
1*
b110 6
19
1>
1C
b110 G
#791380000000
0!
0*
09
0>
0C
#791390000000
1!
1*
b111 6
19
1>
1C
b111 G
#791400000000
0!
0*
09
0>
0C
#791410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#791420000000
0!
0*
09
0>
0C
#791430000000
1!
1*
b1 6
19
1>
1C
b1 G
#791440000000
0!
0*
09
0>
0C
#791450000000
1!
1*
b10 6
19
1>
1C
b10 G
#791460000000
0!
0*
09
0>
0C
#791470000000
1!
1*
b11 6
19
1>
1C
b11 G
#791480000000
0!
0*
09
0>
0C
#791490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#791500000000
0!
0*
09
0>
0C
#791510000000
1!
1*
b101 6
19
1>
1C
b101 G
#791520000000
0!
0*
09
0>
0C
#791530000000
1!
1*
b110 6
19
1>
1C
b110 G
#791540000000
0!
0*
09
0>
0C
#791550000000
1!
1*
b111 6
19
1>
1C
b111 G
#791560000000
0!
1"
0*
1+
09
1:
0>
0C
#791570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#791580000000
0!
0*
09
0>
0C
#791590000000
1!
1*
b1 6
19
1>
1C
b1 G
#791600000000
0!
0*
09
0>
0C
#791610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#791620000000
0!
0*
09
0>
0C
#791630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#791640000000
0!
0*
09
0>
0C
#791650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#791660000000
0!
0*
09
0>
0C
#791670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#791680000000
0!
0#
0*
0,
09
0>
0?
0C
#791690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#791700000000
0!
0*
09
0>
0C
#791710000000
1!
1*
19
1>
1C
#791720000000
0!
0*
09
0>
0C
#791730000000
1!
1*
19
1>
1C
#791740000000
0!
0*
09
0>
0C
#791750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#791760000000
0!
0*
09
0>
0C
#791770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#791780000000
0!
0*
09
0>
0C
#791790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#791800000000
0!
0*
09
0>
0C
#791810000000
1!
1*
b10 6
19
1>
1C
b10 G
#791820000000
0!
0*
09
0>
0C
#791830000000
1!
1*
b11 6
19
1>
1C
b11 G
#791840000000
0!
0*
09
0>
0C
#791850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#791860000000
0!
0*
09
0>
0C
#791870000000
1!
1*
b101 6
19
1>
1C
b101 G
#791880000000
0!
0*
09
0>
0C
#791890000000
1!
1*
b110 6
19
1>
1C
b110 G
#791900000000
0!
0*
09
0>
0C
#791910000000
1!
1*
b111 6
19
1>
1C
b111 G
#791920000000
0!
0*
09
0>
0C
#791930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#791940000000
0!
0*
09
0>
0C
#791950000000
1!
1*
b1 6
19
1>
1C
b1 G
#791960000000
0!
0*
09
0>
0C
#791970000000
1!
1*
b10 6
19
1>
1C
b10 G
#791980000000
0!
0*
09
0>
0C
#791990000000
1!
1*
b11 6
19
1>
1C
b11 G
#792000000000
0!
0*
09
0>
0C
#792010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#792020000000
0!
0*
09
0>
0C
#792030000000
1!
1*
b101 6
19
1>
1C
b101 G
#792040000000
0!
0*
09
0>
0C
#792050000000
1!
1*
b110 6
19
1>
1C
b110 G
#792060000000
0!
0*
09
0>
0C
#792070000000
1!
1*
b111 6
19
1>
1C
b111 G
#792080000000
0!
0*
09
0>
0C
#792090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#792100000000
0!
0*
09
0>
0C
#792110000000
1!
1*
b1 6
19
1>
1C
b1 G
#792120000000
0!
0*
09
0>
0C
#792130000000
1!
1*
b10 6
19
1>
1C
b10 G
#792140000000
0!
0*
09
0>
0C
#792150000000
1!
1*
b11 6
19
1>
1C
b11 G
#792160000000
0!
0*
09
0>
0C
#792170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#792180000000
0!
0*
09
0>
0C
#792190000000
1!
1*
b101 6
19
1>
1C
b101 G
#792200000000
0!
0*
09
0>
0C
#792210000000
1!
1*
b110 6
19
1>
1C
b110 G
#792220000000
0!
0*
09
0>
0C
#792230000000
1!
1*
b111 6
19
1>
1C
b111 G
#792240000000
0!
1"
0*
1+
09
1:
0>
0C
#792250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#792260000000
0!
0*
09
0>
0C
#792270000000
1!
1*
b1 6
19
1>
1C
b1 G
#792280000000
0!
0*
09
0>
0C
#792290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#792300000000
0!
0*
09
0>
0C
#792310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#792320000000
0!
0*
09
0>
0C
#792330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#792340000000
0!
0*
09
0>
0C
#792350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#792360000000
0!
0#
0*
0,
09
0>
0?
0C
#792370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#792380000000
0!
0*
09
0>
0C
#792390000000
1!
1*
19
1>
1C
#792400000000
0!
0*
09
0>
0C
#792410000000
1!
1*
19
1>
1C
#792420000000
0!
0*
09
0>
0C
#792430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#792440000000
0!
0*
09
0>
0C
#792450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#792460000000
0!
0*
09
0>
0C
#792470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#792480000000
0!
0*
09
0>
0C
#792490000000
1!
1*
b10 6
19
1>
1C
b10 G
#792500000000
0!
0*
09
0>
0C
#792510000000
1!
1*
b11 6
19
1>
1C
b11 G
#792520000000
0!
0*
09
0>
0C
#792530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#792540000000
0!
0*
09
0>
0C
#792550000000
1!
1*
b101 6
19
1>
1C
b101 G
#792560000000
0!
0*
09
0>
0C
#792570000000
1!
1*
b110 6
19
1>
1C
b110 G
#792580000000
0!
0*
09
0>
0C
#792590000000
1!
1*
b111 6
19
1>
1C
b111 G
#792600000000
0!
0*
09
0>
0C
#792610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#792620000000
0!
0*
09
0>
0C
#792630000000
1!
1*
b1 6
19
1>
1C
b1 G
#792640000000
0!
0*
09
0>
0C
#792650000000
1!
1*
b10 6
19
1>
1C
b10 G
#792660000000
0!
0*
09
0>
0C
#792670000000
1!
1*
b11 6
19
1>
1C
b11 G
#792680000000
0!
0*
09
0>
0C
#792690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#792700000000
0!
0*
09
0>
0C
#792710000000
1!
1*
b101 6
19
1>
1C
b101 G
#792720000000
0!
0*
09
0>
0C
#792730000000
1!
1*
b110 6
19
1>
1C
b110 G
#792740000000
0!
0*
09
0>
0C
#792750000000
1!
1*
b111 6
19
1>
1C
b111 G
#792760000000
0!
0*
09
0>
0C
#792770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#792780000000
0!
0*
09
0>
0C
#792790000000
1!
1*
b1 6
19
1>
1C
b1 G
#792800000000
0!
0*
09
0>
0C
#792810000000
1!
1*
b10 6
19
1>
1C
b10 G
#792820000000
0!
0*
09
0>
0C
#792830000000
1!
1*
b11 6
19
1>
1C
b11 G
#792840000000
0!
0*
09
0>
0C
#792850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#792860000000
0!
0*
09
0>
0C
#792870000000
1!
1*
b101 6
19
1>
1C
b101 G
#792880000000
0!
0*
09
0>
0C
#792890000000
1!
1*
b110 6
19
1>
1C
b110 G
#792900000000
0!
0*
09
0>
0C
#792910000000
1!
1*
b111 6
19
1>
1C
b111 G
#792920000000
0!
1"
0*
1+
09
1:
0>
0C
#792930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#792940000000
0!
0*
09
0>
0C
#792950000000
1!
1*
b1 6
19
1>
1C
b1 G
#792960000000
0!
0*
09
0>
0C
#792970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#792980000000
0!
0*
09
0>
0C
#792990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#793000000000
0!
0*
09
0>
0C
#793010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#793020000000
0!
0*
09
0>
0C
#793030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#793040000000
0!
0#
0*
0,
09
0>
0?
0C
#793050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#793060000000
0!
0*
09
0>
0C
#793070000000
1!
1*
19
1>
1C
#793080000000
0!
0*
09
0>
0C
#793090000000
1!
1*
19
1>
1C
#793100000000
0!
0*
09
0>
0C
#793110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#793120000000
0!
0*
09
0>
0C
#793130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#793140000000
0!
0*
09
0>
0C
#793150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#793160000000
0!
0*
09
0>
0C
#793170000000
1!
1*
b10 6
19
1>
1C
b10 G
#793180000000
0!
0*
09
0>
0C
#793190000000
1!
1*
b11 6
19
1>
1C
b11 G
#793200000000
0!
0*
09
0>
0C
#793210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#793220000000
0!
0*
09
0>
0C
#793230000000
1!
1*
b101 6
19
1>
1C
b101 G
#793240000000
0!
0*
09
0>
0C
#793250000000
1!
1*
b110 6
19
1>
1C
b110 G
#793260000000
0!
0*
09
0>
0C
#793270000000
1!
1*
b111 6
19
1>
1C
b111 G
#793280000000
0!
0*
09
0>
0C
#793290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#793300000000
0!
0*
09
0>
0C
#793310000000
1!
1*
b1 6
19
1>
1C
b1 G
#793320000000
0!
0*
09
0>
0C
#793330000000
1!
1*
b10 6
19
1>
1C
b10 G
#793340000000
0!
0*
09
0>
0C
#793350000000
1!
1*
b11 6
19
1>
1C
b11 G
#793360000000
0!
0*
09
0>
0C
#793370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#793380000000
0!
0*
09
0>
0C
#793390000000
1!
1*
b101 6
19
1>
1C
b101 G
#793400000000
0!
0*
09
0>
0C
#793410000000
1!
1*
b110 6
19
1>
1C
b110 G
#793420000000
0!
0*
09
0>
0C
#793430000000
1!
1*
b111 6
19
1>
1C
b111 G
#793440000000
0!
0*
09
0>
0C
#793450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#793460000000
0!
0*
09
0>
0C
#793470000000
1!
1*
b1 6
19
1>
1C
b1 G
#793480000000
0!
0*
09
0>
0C
#793490000000
1!
1*
b10 6
19
1>
1C
b10 G
#793500000000
0!
0*
09
0>
0C
#793510000000
1!
1*
b11 6
19
1>
1C
b11 G
#793520000000
0!
0*
09
0>
0C
#793530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#793540000000
0!
0*
09
0>
0C
#793550000000
1!
1*
b101 6
19
1>
1C
b101 G
#793560000000
0!
0*
09
0>
0C
#793570000000
1!
1*
b110 6
19
1>
1C
b110 G
#793580000000
0!
0*
09
0>
0C
#793590000000
1!
1*
b111 6
19
1>
1C
b111 G
#793600000000
0!
1"
0*
1+
09
1:
0>
0C
#793610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#793620000000
0!
0*
09
0>
0C
#793630000000
1!
1*
b1 6
19
1>
1C
b1 G
#793640000000
0!
0*
09
0>
0C
#793650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#793660000000
0!
0*
09
0>
0C
#793670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#793680000000
0!
0*
09
0>
0C
#793690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#793700000000
0!
0*
09
0>
0C
#793710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#793720000000
0!
0#
0*
0,
09
0>
0?
0C
#793730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#793740000000
0!
0*
09
0>
0C
#793750000000
1!
1*
19
1>
1C
#793760000000
0!
0*
09
0>
0C
#793770000000
1!
1*
19
1>
1C
#793780000000
0!
0*
09
0>
0C
#793790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#793800000000
0!
0*
09
0>
0C
#793810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#793820000000
0!
0*
09
0>
0C
#793830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#793840000000
0!
0*
09
0>
0C
#793850000000
1!
1*
b10 6
19
1>
1C
b10 G
#793860000000
0!
0*
09
0>
0C
#793870000000
1!
1*
b11 6
19
1>
1C
b11 G
#793880000000
0!
0*
09
0>
0C
#793890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#793900000000
0!
0*
09
0>
0C
#793910000000
1!
1*
b101 6
19
1>
1C
b101 G
#793920000000
0!
0*
09
0>
0C
#793930000000
1!
1*
b110 6
19
1>
1C
b110 G
#793940000000
0!
0*
09
0>
0C
#793950000000
1!
1*
b111 6
19
1>
1C
b111 G
#793960000000
0!
0*
09
0>
0C
#793970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#793980000000
0!
0*
09
0>
0C
#793990000000
1!
1*
b1 6
19
1>
1C
b1 G
#794000000000
0!
0*
09
0>
0C
#794010000000
1!
1*
b10 6
19
1>
1C
b10 G
#794020000000
0!
0*
09
0>
0C
#794030000000
1!
1*
b11 6
19
1>
1C
b11 G
#794040000000
0!
0*
09
0>
0C
#794050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#794060000000
0!
0*
09
0>
0C
#794070000000
1!
1*
b101 6
19
1>
1C
b101 G
#794080000000
0!
0*
09
0>
0C
#794090000000
1!
1*
b110 6
19
1>
1C
b110 G
#794100000000
0!
0*
09
0>
0C
#794110000000
1!
1*
b111 6
19
1>
1C
b111 G
#794120000000
0!
0*
09
0>
0C
#794130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#794140000000
0!
0*
09
0>
0C
#794150000000
1!
1*
b1 6
19
1>
1C
b1 G
#794160000000
0!
0*
09
0>
0C
#794170000000
1!
1*
b10 6
19
1>
1C
b10 G
#794180000000
0!
0*
09
0>
0C
#794190000000
1!
1*
b11 6
19
1>
1C
b11 G
#794200000000
0!
0*
09
0>
0C
#794210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#794220000000
0!
0*
09
0>
0C
#794230000000
1!
1*
b101 6
19
1>
1C
b101 G
#794240000000
0!
0*
09
0>
0C
#794250000000
1!
1*
b110 6
19
1>
1C
b110 G
#794260000000
0!
0*
09
0>
0C
#794270000000
1!
1*
b111 6
19
1>
1C
b111 G
#794280000000
0!
1"
0*
1+
09
1:
0>
0C
#794290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#794300000000
0!
0*
09
0>
0C
#794310000000
1!
1*
b1 6
19
1>
1C
b1 G
#794320000000
0!
0*
09
0>
0C
#794330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#794340000000
0!
0*
09
0>
0C
#794350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#794360000000
0!
0*
09
0>
0C
#794370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#794380000000
0!
0*
09
0>
0C
#794390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#794400000000
0!
0#
0*
0,
09
0>
0?
0C
#794410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#794420000000
0!
0*
09
0>
0C
#794430000000
1!
1*
19
1>
1C
#794440000000
0!
0*
09
0>
0C
#794450000000
1!
1*
19
1>
1C
#794460000000
0!
0*
09
0>
0C
#794470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#794480000000
0!
0*
09
0>
0C
#794490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#794500000000
0!
0*
09
0>
0C
#794510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#794520000000
0!
0*
09
0>
0C
#794530000000
1!
1*
b10 6
19
1>
1C
b10 G
#794540000000
0!
0*
09
0>
0C
#794550000000
1!
1*
b11 6
19
1>
1C
b11 G
#794560000000
0!
0*
09
0>
0C
#794570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#794580000000
0!
0*
09
0>
0C
#794590000000
1!
1*
b101 6
19
1>
1C
b101 G
#794600000000
0!
0*
09
0>
0C
#794610000000
1!
1*
b110 6
19
1>
1C
b110 G
#794620000000
0!
0*
09
0>
0C
#794630000000
1!
1*
b111 6
19
1>
1C
b111 G
#794640000000
0!
0*
09
0>
0C
#794650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#794660000000
0!
0*
09
0>
0C
#794670000000
1!
1*
b1 6
19
1>
1C
b1 G
#794680000000
0!
0*
09
0>
0C
#794690000000
1!
1*
b10 6
19
1>
1C
b10 G
#794700000000
0!
0*
09
0>
0C
#794710000000
1!
1*
b11 6
19
1>
1C
b11 G
#794720000000
0!
0*
09
0>
0C
#794730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#794740000000
0!
0*
09
0>
0C
#794750000000
1!
1*
b101 6
19
1>
1C
b101 G
#794760000000
0!
0*
09
0>
0C
#794770000000
1!
1*
b110 6
19
1>
1C
b110 G
#794780000000
0!
0*
09
0>
0C
#794790000000
1!
1*
b111 6
19
1>
1C
b111 G
#794800000000
0!
0*
09
0>
0C
#794810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#794820000000
0!
0*
09
0>
0C
#794830000000
1!
1*
b1 6
19
1>
1C
b1 G
#794840000000
0!
0*
09
0>
0C
#794850000000
1!
1*
b10 6
19
1>
1C
b10 G
#794860000000
0!
0*
09
0>
0C
#794870000000
1!
1*
b11 6
19
1>
1C
b11 G
#794880000000
0!
0*
09
0>
0C
#794890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#794900000000
0!
0*
09
0>
0C
#794910000000
1!
1*
b101 6
19
1>
1C
b101 G
#794920000000
0!
0*
09
0>
0C
#794930000000
1!
1*
b110 6
19
1>
1C
b110 G
#794940000000
0!
0*
09
0>
0C
#794950000000
1!
1*
b111 6
19
1>
1C
b111 G
#794960000000
0!
1"
0*
1+
09
1:
0>
0C
#794970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#794980000000
0!
0*
09
0>
0C
#794990000000
1!
1*
b1 6
19
1>
1C
b1 G
#795000000000
0!
0*
09
0>
0C
#795010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#795020000000
0!
0*
09
0>
0C
#795030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#795040000000
0!
0*
09
0>
0C
#795050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#795060000000
0!
0*
09
0>
0C
#795070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#795080000000
0!
0#
0*
0,
09
0>
0?
0C
#795090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#795100000000
0!
0*
09
0>
0C
#795110000000
1!
1*
19
1>
1C
#795120000000
0!
0*
09
0>
0C
#795130000000
1!
1*
19
1>
1C
#795140000000
0!
0*
09
0>
0C
#795150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#795160000000
0!
0*
09
0>
0C
#795170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#795180000000
0!
0*
09
0>
0C
#795190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#795200000000
0!
0*
09
0>
0C
#795210000000
1!
1*
b10 6
19
1>
1C
b10 G
#795220000000
0!
0*
09
0>
0C
#795230000000
1!
1*
b11 6
19
1>
1C
b11 G
#795240000000
0!
0*
09
0>
0C
#795250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#795260000000
0!
0*
09
0>
0C
#795270000000
1!
1*
b101 6
19
1>
1C
b101 G
#795280000000
0!
0*
09
0>
0C
#795290000000
1!
1*
b110 6
19
1>
1C
b110 G
#795300000000
0!
0*
09
0>
0C
#795310000000
1!
1*
b111 6
19
1>
1C
b111 G
#795320000000
0!
0*
09
0>
0C
#795330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#795340000000
0!
0*
09
0>
0C
#795350000000
1!
1*
b1 6
19
1>
1C
b1 G
#795360000000
0!
0*
09
0>
0C
#795370000000
1!
1*
b10 6
19
1>
1C
b10 G
#795380000000
0!
0*
09
0>
0C
#795390000000
1!
1*
b11 6
19
1>
1C
b11 G
#795400000000
0!
0*
09
0>
0C
#795410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#795420000000
0!
0*
09
0>
0C
#795430000000
1!
1*
b101 6
19
1>
1C
b101 G
#795440000000
0!
0*
09
0>
0C
#795450000000
1!
1*
b110 6
19
1>
1C
b110 G
#795460000000
0!
0*
09
0>
0C
#795470000000
1!
1*
b111 6
19
1>
1C
b111 G
#795480000000
0!
0*
09
0>
0C
#795490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#795500000000
0!
0*
09
0>
0C
#795510000000
1!
1*
b1 6
19
1>
1C
b1 G
#795520000000
0!
0*
09
0>
0C
#795530000000
1!
1*
b10 6
19
1>
1C
b10 G
#795540000000
0!
0*
09
0>
0C
#795550000000
1!
1*
b11 6
19
1>
1C
b11 G
#795560000000
0!
0*
09
0>
0C
#795570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#795580000000
0!
0*
09
0>
0C
#795590000000
1!
1*
b101 6
19
1>
1C
b101 G
#795600000000
0!
0*
09
0>
0C
#795610000000
1!
1*
b110 6
19
1>
1C
b110 G
#795620000000
0!
0*
09
0>
0C
#795630000000
1!
1*
b111 6
19
1>
1C
b111 G
#795640000000
0!
1"
0*
1+
09
1:
0>
0C
#795650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#795660000000
0!
0*
09
0>
0C
#795670000000
1!
1*
b1 6
19
1>
1C
b1 G
#795680000000
0!
0*
09
0>
0C
#795690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#795700000000
0!
0*
09
0>
0C
#795710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#795720000000
0!
0*
09
0>
0C
#795730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#795740000000
0!
0*
09
0>
0C
#795750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#795760000000
0!
0#
0*
0,
09
0>
0?
0C
#795770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#795780000000
0!
0*
09
0>
0C
#795790000000
1!
1*
19
1>
1C
#795800000000
0!
0*
09
0>
0C
#795810000000
1!
1*
19
1>
1C
#795820000000
0!
0*
09
0>
0C
#795830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#795840000000
0!
0*
09
0>
0C
#795850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#795860000000
0!
0*
09
0>
0C
#795870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#795880000000
0!
0*
09
0>
0C
#795890000000
1!
1*
b10 6
19
1>
1C
b10 G
#795900000000
0!
0*
09
0>
0C
#795910000000
1!
1*
b11 6
19
1>
1C
b11 G
#795920000000
0!
0*
09
0>
0C
#795930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#795940000000
0!
0*
09
0>
0C
#795950000000
1!
1*
b101 6
19
1>
1C
b101 G
#795960000000
0!
0*
09
0>
0C
#795970000000
1!
1*
b110 6
19
1>
1C
b110 G
#795980000000
0!
0*
09
0>
0C
#795990000000
1!
1*
b111 6
19
1>
1C
b111 G
#796000000000
0!
0*
09
0>
0C
#796010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#796020000000
0!
0*
09
0>
0C
#796030000000
1!
1*
b1 6
19
1>
1C
b1 G
#796040000000
0!
0*
09
0>
0C
#796050000000
1!
1*
b10 6
19
1>
1C
b10 G
#796060000000
0!
0*
09
0>
0C
#796070000000
1!
1*
b11 6
19
1>
1C
b11 G
#796080000000
0!
0*
09
0>
0C
#796090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#796100000000
0!
0*
09
0>
0C
#796110000000
1!
1*
b101 6
19
1>
1C
b101 G
#796120000000
0!
0*
09
0>
0C
#796130000000
1!
1*
b110 6
19
1>
1C
b110 G
#796140000000
0!
0*
09
0>
0C
#796150000000
1!
1*
b111 6
19
1>
1C
b111 G
#796160000000
0!
0*
09
0>
0C
#796170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#796180000000
0!
0*
09
0>
0C
#796190000000
1!
1*
b1 6
19
1>
1C
b1 G
#796200000000
0!
0*
09
0>
0C
#796210000000
1!
1*
b10 6
19
1>
1C
b10 G
#796220000000
0!
0*
09
0>
0C
#796230000000
1!
1*
b11 6
19
1>
1C
b11 G
#796240000000
0!
0*
09
0>
0C
#796250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#796260000000
0!
0*
09
0>
0C
#796270000000
1!
1*
b101 6
19
1>
1C
b101 G
#796280000000
0!
0*
09
0>
0C
#796290000000
1!
1*
b110 6
19
1>
1C
b110 G
#796300000000
0!
0*
09
0>
0C
#796310000000
1!
1*
b111 6
19
1>
1C
b111 G
#796320000000
0!
1"
0*
1+
09
1:
0>
0C
#796330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#796340000000
0!
0*
09
0>
0C
#796350000000
1!
1*
b1 6
19
1>
1C
b1 G
#796360000000
0!
0*
09
0>
0C
#796370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#796380000000
0!
0*
09
0>
0C
#796390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#796400000000
0!
0*
09
0>
0C
#796410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#796420000000
0!
0*
09
0>
0C
#796430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#796440000000
0!
0#
0*
0,
09
0>
0?
0C
#796450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#796460000000
0!
0*
09
0>
0C
#796470000000
1!
1*
19
1>
1C
#796480000000
0!
0*
09
0>
0C
#796490000000
1!
1*
19
1>
1C
#796500000000
0!
0*
09
0>
0C
#796510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#796520000000
0!
0*
09
0>
0C
#796530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#796540000000
0!
0*
09
0>
0C
#796550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#796560000000
0!
0*
09
0>
0C
#796570000000
1!
1*
b10 6
19
1>
1C
b10 G
#796580000000
0!
0*
09
0>
0C
#796590000000
1!
1*
b11 6
19
1>
1C
b11 G
#796600000000
0!
0*
09
0>
0C
#796610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#796620000000
0!
0*
09
0>
0C
#796630000000
1!
1*
b101 6
19
1>
1C
b101 G
#796640000000
0!
0*
09
0>
0C
#796650000000
1!
1*
b110 6
19
1>
1C
b110 G
#796660000000
0!
0*
09
0>
0C
#796670000000
1!
1*
b111 6
19
1>
1C
b111 G
#796680000000
0!
0*
09
0>
0C
#796690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#796700000000
0!
0*
09
0>
0C
#796710000000
1!
1*
b1 6
19
1>
1C
b1 G
#796720000000
0!
0*
09
0>
0C
#796730000000
1!
1*
b10 6
19
1>
1C
b10 G
#796740000000
0!
0*
09
0>
0C
#796750000000
1!
1*
b11 6
19
1>
1C
b11 G
#796760000000
0!
0*
09
0>
0C
#796770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#796780000000
0!
0*
09
0>
0C
#796790000000
1!
1*
b101 6
19
1>
1C
b101 G
#796800000000
0!
0*
09
0>
0C
#796810000000
1!
1*
b110 6
19
1>
1C
b110 G
#796820000000
0!
0*
09
0>
0C
#796830000000
1!
1*
b111 6
19
1>
1C
b111 G
#796840000000
0!
0*
09
0>
0C
#796850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#796860000000
0!
0*
09
0>
0C
#796870000000
1!
1*
b1 6
19
1>
1C
b1 G
#796880000000
0!
0*
09
0>
0C
#796890000000
1!
1*
b10 6
19
1>
1C
b10 G
#796900000000
0!
0*
09
0>
0C
#796910000000
1!
1*
b11 6
19
1>
1C
b11 G
#796920000000
0!
0*
09
0>
0C
#796930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#796940000000
0!
0*
09
0>
0C
#796950000000
1!
1*
b101 6
19
1>
1C
b101 G
#796960000000
0!
0*
09
0>
0C
#796970000000
1!
1*
b110 6
19
1>
1C
b110 G
#796980000000
0!
0*
09
0>
0C
#796990000000
1!
1*
b111 6
19
1>
1C
b111 G
#797000000000
0!
1"
0*
1+
09
1:
0>
0C
#797010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#797020000000
0!
0*
09
0>
0C
#797030000000
1!
1*
b1 6
19
1>
1C
b1 G
#797040000000
0!
0*
09
0>
0C
#797050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#797060000000
0!
0*
09
0>
0C
#797070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#797080000000
0!
0*
09
0>
0C
#797090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#797100000000
0!
0*
09
0>
0C
#797110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#797120000000
0!
0#
0*
0,
09
0>
0?
0C
#797130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#797140000000
0!
0*
09
0>
0C
#797150000000
1!
1*
19
1>
1C
#797160000000
0!
0*
09
0>
0C
#797170000000
1!
1*
19
1>
1C
#797180000000
0!
0*
09
0>
0C
#797190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#797200000000
0!
0*
09
0>
0C
#797210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#797220000000
0!
0*
09
0>
0C
#797230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#797240000000
0!
0*
09
0>
0C
#797250000000
1!
1*
b10 6
19
1>
1C
b10 G
#797260000000
0!
0*
09
0>
0C
#797270000000
1!
1*
b11 6
19
1>
1C
b11 G
#797280000000
0!
0*
09
0>
0C
#797290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#797300000000
0!
0*
09
0>
0C
#797310000000
1!
1*
b101 6
19
1>
1C
b101 G
#797320000000
0!
0*
09
0>
0C
#797330000000
1!
1*
b110 6
19
1>
1C
b110 G
#797340000000
0!
0*
09
0>
0C
#797350000000
1!
1*
b111 6
19
1>
1C
b111 G
#797360000000
0!
0*
09
0>
0C
#797370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#797380000000
0!
0*
09
0>
0C
#797390000000
1!
1*
b1 6
19
1>
1C
b1 G
#797400000000
0!
0*
09
0>
0C
#797410000000
1!
1*
b10 6
19
1>
1C
b10 G
#797420000000
0!
0*
09
0>
0C
#797430000000
1!
1*
b11 6
19
1>
1C
b11 G
#797440000000
0!
0*
09
0>
0C
#797450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#797460000000
0!
0*
09
0>
0C
#797470000000
1!
1*
b101 6
19
1>
1C
b101 G
#797480000000
0!
0*
09
0>
0C
#797490000000
1!
1*
b110 6
19
1>
1C
b110 G
#797500000000
0!
0*
09
0>
0C
#797510000000
1!
1*
b111 6
19
1>
1C
b111 G
#797520000000
0!
0*
09
0>
0C
#797530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#797540000000
0!
0*
09
0>
0C
#797550000000
1!
1*
b1 6
19
1>
1C
b1 G
#797560000000
0!
0*
09
0>
0C
#797570000000
1!
1*
b10 6
19
1>
1C
b10 G
#797580000000
0!
0*
09
0>
0C
#797590000000
1!
1*
b11 6
19
1>
1C
b11 G
#797600000000
0!
0*
09
0>
0C
#797610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#797620000000
0!
0*
09
0>
0C
#797630000000
1!
1*
b101 6
19
1>
1C
b101 G
#797640000000
0!
0*
09
0>
0C
#797650000000
1!
1*
b110 6
19
1>
1C
b110 G
#797660000000
0!
0*
09
0>
0C
#797670000000
1!
1*
b111 6
19
1>
1C
b111 G
#797680000000
0!
1"
0*
1+
09
1:
0>
0C
#797690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#797700000000
0!
0*
09
0>
0C
#797710000000
1!
1*
b1 6
19
1>
1C
b1 G
#797720000000
0!
0*
09
0>
0C
#797730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#797740000000
0!
0*
09
0>
0C
#797750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#797760000000
0!
0*
09
0>
0C
#797770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#797780000000
0!
0*
09
0>
0C
#797790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#797800000000
0!
0#
0*
0,
09
0>
0?
0C
#797810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#797820000000
0!
0*
09
0>
0C
#797830000000
1!
1*
19
1>
1C
#797840000000
0!
0*
09
0>
0C
#797850000000
1!
1*
19
1>
1C
#797860000000
0!
0*
09
0>
0C
#797870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#797880000000
0!
0*
09
0>
0C
#797890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#797900000000
0!
0*
09
0>
0C
#797910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#797920000000
0!
0*
09
0>
0C
#797930000000
1!
1*
b10 6
19
1>
1C
b10 G
#797940000000
0!
0*
09
0>
0C
#797950000000
1!
1*
b11 6
19
1>
1C
b11 G
#797960000000
0!
0*
09
0>
0C
#797970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#797980000000
0!
0*
09
0>
0C
#797990000000
1!
1*
b101 6
19
1>
1C
b101 G
#798000000000
0!
0*
09
0>
0C
#798010000000
1!
1*
b110 6
19
1>
1C
b110 G
#798020000000
0!
0*
09
0>
0C
#798030000000
1!
1*
b111 6
19
1>
1C
b111 G
#798040000000
0!
0*
09
0>
0C
#798050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#798060000000
0!
0*
09
0>
0C
#798070000000
1!
1*
b1 6
19
1>
1C
b1 G
#798080000000
0!
0*
09
0>
0C
#798090000000
1!
1*
b10 6
19
1>
1C
b10 G
#798100000000
0!
0*
09
0>
0C
#798110000000
1!
1*
b11 6
19
1>
1C
b11 G
#798120000000
0!
0*
09
0>
0C
#798130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#798140000000
0!
0*
09
0>
0C
#798150000000
1!
1*
b101 6
19
1>
1C
b101 G
#798160000000
0!
0*
09
0>
0C
#798170000000
1!
1*
b110 6
19
1>
1C
b110 G
#798180000000
0!
0*
09
0>
0C
#798190000000
1!
1*
b111 6
19
1>
1C
b111 G
#798200000000
0!
0*
09
0>
0C
#798210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#798220000000
0!
0*
09
0>
0C
#798230000000
1!
1*
b1 6
19
1>
1C
b1 G
#798240000000
0!
0*
09
0>
0C
#798250000000
1!
1*
b10 6
19
1>
1C
b10 G
#798260000000
0!
0*
09
0>
0C
#798270000000
1!
1*
b11 6
19
1>
1C
b11 G
#798280000000
0!
0*
09
0>
0C
#798290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#798300000000
0!
0*
09
0>
0C
#798310000000
1!
1*
b101 6
19
1>
1C
b101 G
#798320000000
0!
0*
09
0>
0C
#798330000000
1!
1*
b110 6
19
1>
1C
b110 G
#798340000000
0!
0*
09
0>
0C
#798350000000
1!
1*
b111 6
19
1>
1C
b111 G
#798360000000
0!
1"
0*
1+
09
1:
0>
0C
#798370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#798380000000
0!
0*
09
0>
0C
#798390000000
1!
1*
b1 6
19
1>
1C
b1 G
#798400000000
0!
0*
09
0>
0C
#798410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#798420000000
0!
0*
09
0>
0C
#798430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#798440000000
0!
0*
09
0>
0C
#798450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#798460000000
0!
0*
09
0>
0C
#798470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#798480000000
0!
0#
0*
0,
09
0>
0?
0C
#798490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#798500000000
0!
0*
09
0>
0C
#798510000000
1!
1*
19
1>
1C
#798520000000
0!
0*
09
0>
0C
#798530000000
1!
1*
19
1>
1C
#798540000000
0!
0*
09
0>
0C
#798550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#798560000000
0!
0*
09
0>
0C
#798570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#798580000000
0!
0*
09
0>
0C
#798590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#798600000000
0!
0*
09
0>
0C
#798610000000
1!
1*
b10 6
19
1>
1C
b10 G
#798620000000
0!
0*
09
0>
0C
#798630000000
1!
1*
b11 6
19
1>
1C
b11 G
#798640000000
0!
0*
09
0>
0C
#798650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#798660000000
0!
0*
09
0>
0C
#798670000000
1!
1*
b101 6
19
1>
1C
b101 G
#798680000000
0!
0*
09
0>
0C
#798690000000
1!
1*
b110 6
19
1>
1C
b110 G
#798700000000
0!
0*
09
0>
0C
#798710000000
1!
1*
b111 6
19
1>
1C
b111 G
#798720000000
0!
0*
09
0>
0C
#798730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#798740000000
0!
0*
09
0>
0C
#798750000000
1!
1*
b1 6
19
1>
1C
b1 G
#798760000000
0!
0*
09
0>
0C
#798770000000
1!
1*
b10 6
19
1>
1C
b10 G
#798780000000
0!
0*
09
0>
0C
#798790000000
1!
1*
b11 6
19
1>
1C
b11 G
#798800000000
0!
0*
09
0>
0C
#798810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#798820000000
0!
0*
09
0>
0C
#798830000000
1!
1*
b101 6
19
1>
1C
b101 G
#798840000000
0!
0*
09
0>
0C
#798850000000
1!
1*
b110 6
19
1>
1C
b110 G
#798860000000
0!
0*
09
0>
0C
#798870000000
1!
1*
b111 6
19
1>
1C
b111 G
#798880000000
0!
0*
09
0>
0C
#798890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#798900000000
0!
0*
09
0>
0C
#798910000000
1!
1*
b1 6
19
1>
1C
b1 G
#798920000000
0!
0*
09
0>
0C
#798930000000
1!
1*
b10 6
19
1>
1C
b10 G
#798940000000
0!
0*
09
0>
0C
#798950000000
1!
1*
b11 6
19
1>
1C
b11 G
#798960000000
0!
0*
09
0>
0C
#798970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#798980000000
0!
0*
09
0>
0C
#798990000000
1!
1*
b101 6
19
1>
1C
b101 G
#799000000000
0!
0*
09
0>
0C
#799010000000
1!
1*
b110 6
19
1>
1C
b110 G
#799020000000
0!
0*
09
0>
0C
#799030000000
1!
1*
b111 6
19
1>
1C
b111 G
#799040000000
0!
1"
0*
1+
09
1:
0>
0C
#799050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#799060000000
0!
0*
09
0>
0C
#799070000000
1!
1*
b1 6
19
1>
1C
b1 G
#799080000000
0!
0*
09
0>
0C
#799090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#799100000000
0!
0*
09
0>
0C
#799110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#799120000000
0!
0*
09
0>
0C
#799130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#799140000000
0!
0*
09
0>
0C
#799150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#799160000000
0!
0#
0*
0,
09
0>
0?
0C
#799170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#799180000000
0!
0*
09
0>
0C
#799190000000
1!
1*
19
1>
1C
#799200000000
0!
0*
09
0>
0C
#799210000000
1!
1*
19
1>
1C
#799220000000
0!
0*
09
0>
0C
#799230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#799240000000
0!
0*
09
0>
0C
#799250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#799260000000
0!
0*
09
0>
0C
#799270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#799280000000
0!
0*
09
0>
0C
#799290000000
1!
1*
b10 6
19
1>
1C
b10 G
#799300000000
0!
0*
09
0>
0C
#799310000000
1!
1*
b11 6
19
1>
1C
b11 G
#799320000000
0!
0*
09
0>
0C
#799330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#799340000000
0!
0*
09
0>
0C
#799350000000
1!
1*
b101 6
19
1>
1C
b101 G
#799360000000
0!
0*
09
0>
0C
#799370000000
1!
1*
b110 6
19
1>
1C
b110 G
#799380000000
0!
0*
09
0>
0C
#799390000000
1!
1*
b111 6
19
1>
1C
b111 G
#799400000000
0!
0*
09
0>
0C
#799410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#799420000000
0!
0*
09
0>
0C
#799430000000
1!
1*
b1 6
19
1>
1C
b1 G
#799440000000
0!
0*
09
0>
0C
#799450000000
1!
1*
b10 6
19
1>
1C
b10 G
#799460000000
0!
0*
09
0>
0C
#799470000000
1!
1*
b11 6
19
1>
1C
b11 G
#799480000000
0!
0*
09
0>
0C
#799490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#799500000000
0!
0*
09
0>
0C
#799510000000
1!
1*
b101 6
19
1>
1C
b101 G
#799520000000
0!
0*
09
0>
0C
#799530000000
1!
1*
b110 6
19
1>
1C
b110 G
#799540000000
0!
0*
09
0>
0C
#799550000000
1!
1*
b111 6
19
1>
1C
b111 G
#799560000000
0!
0*
09
0>
0C
#799570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#799580000000
0!
0*
09
0>
0C
#799590000000
1!
1*
b1 6
19
1>
1C
b1 G
#799600000000
0!
0*
09
0>
0C
#799610000000
1!
1*
b10 6
19
1>
1C
b10 G
#799620000000
0!
0*
09
0>
0C
#799630000000
1!
1*
b11 6
19
1>
1C
b11 G
#799640000000
0!
0*
09
0>
0C
#799650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#799660000000
0!
0*
09
0>
0C
#799670000000
1!
1*
b101 6
19
1>
1C
b101 G
#799680000000
0!
0*
09
0>
0C
#799690000000
1!
1*
b110 6
19
1>
1C
b110 G
#799700000000
0!
0*
09
0>
0C
#799710000000
1!
1*
b111 6
19
1>
1C
b111 G
#799720000000
0!
1"
0*
1+
09
1:
0>
0C
#799730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#799740000000
0!
0*
09
0>
0C
#799750000000
1!
1*
b1 6
19
1>
1C
b1 G
#799760000000
0!
0*
09
0>
0C
#799770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#799780000000
0!
0*
09
0>
0C
#799790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#799800000000
0!
0*
09
0>
0C
#799810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#799820000000
0!
0*
09
0>
0C
#799830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#799840000000
0!
0#
0*
0,
09
0>
0?
0C
#799850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#799860000000
0!
0*
09
0>
0C
#799870000000
1!
1*
19
1>
1C
#799880000000
0!
0*
09
0>
0C
#799890000000
1!
1*
19
1>
1C
#799900000000
0!
0*
09
0>
0C
#799910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#799920000000
0!
0*
09
0>
0C
#799930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#799940000000
0!
0*
09
0>
0C
#799950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#799960000000
0!
0*
09
0>
0C
#799970000000
1!
1*
b10 6
19
1>
1C
b10 G
#799980000000
0!
0*
09
0>
0C
#799990000000
1!
1*
b11 6
19
1>
1C
b11 G
#800000000000
0!
0*
09
0>
0C
#800010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#800020000000
0!
0*
09
0>
0C
#800030000000
1!
1*
b101 6
19
1>
1C
b101 G
#800040000000
0!
0*
09
0>
0C
#800050000000
1!
1*
b110 6
19
1>
1C
b110 G
#800060000000
0!
0*
09
0>
0C
#800070000000
1!
1*
b111 6
19
1>
1C
b111 G
#800080000000
0!
0*
09
0>
0C
#800090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#800100000000
0!
0*
09
0>
0C
#800110000000
1!
1*
b1 6
19
1>
1C
b1 G
#800120000000
0!
0*
09
0>
0C
#800130000000
1!
1*
b10 6
19
1>
1C
b10 G
#800140000000
0!
0*
09
0>
0C
#800150000000
1!
1*
b11 6
19
1>
1C
b11 G
#800160000000
0!
0*
09
0>
0C
#800170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#800180000000
0!
0*
09
0>
0C
#800190000000
1!
1*
b101 6
19
1>
1C
b101 G
#800200000000
0!
0*
09
0>
0C
#800210000000
1!
1*
b110 6
19
1>
1C
b110 G
#800220000000
0!
0*
09
0>
0C
#800230000000
1!
1*
b111 6
19
1>
1C
b111 G
#800240000000
0!
0*
09
0>
0C
#800250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#800260000000
0!
0*
09
0>
0C
#800270000000
1!
1*
b1 6
19
1>
1C
b1 G
#800280000000
0!
0*
09
0>
0C
#800290000000
1!
1*
b10 6
19
1>
1C
b10 G
#800300000000
0!
0*
09
0>
0C
#800310000000
1!
1*
b11 6
19
1>
1C
b11 G
#800320000000
0!
0*
09
0>
0C
#800330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#800340000000
0!
0*
09
0>
0C
#800350000000
1!
1*
b101 6
19
1>
1C
b101 G
#800360000000
0!
0*
09
0>
0C
#800370000000
1!
1*
b110 6
19
1>
1C
b110 G
#800380000000
0!
0*
09
0>
0C
#800390000000
1!
1*
b111 6
19
1>
1C
b111 G
#800400000000
0!
1"
0*
1+
09
1:
0>
0C
#800410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#800420000000
0!
0*
09
0>
0C
#800430000000
1!
1*
b1 6
19
1>
1C
b1 G
#800440000000
0!
0*
09
0>
0C
#800450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#800460000000
0!
0*
09
0>
0C
#800470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#800480000000
0!
0*
09
0>
0C
#800490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#800500000000
0!
0*
09
0>
0C
#800510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#800520000000
0!
0#
0*
0,
09
0>
0?
0C
#800530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#800540000000
0!
0*
09
0>
0C
#800550000000
1!
1*
19
1>
1C
#800560000000
0!
0*
09
0>
0C
#800570000000
1!
1*
19
1>
1C
#800580000000
0!
0*
09
0>
0C
#800590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#800600000000
0!
0*
09
0>
0C
#800610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#800620000000
0!
0*
09
0>
0C
#800630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#800640000000
0!
0*
09
0>
0C
#800650000000
1!
1*
b10 6
19
1>
1C
b10 G
#800660000000
0!
0*
09
0>
0C
#800670000000
1!
1*
b11 6
19
1>
1C
b11 G
#800680000000
0!
0*
09
0>
0C
#800690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#800700000000
0!
0*
09
0>
0C
#800710000000
1!
1*
b101 6
19
1>
1C
b101 G
#800720000000
0!
0*
09
0>
0C
#800730000000
1!
1*
b110 6
19
1>
1C
b110 G
#800740000000
0!
0*
09
0>
0C
#800750000000
1!
1*
b111 6
19
1>
1C
b111 G
#800760000000
0!
0*
09
0>
0C
#800770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#800780000000
0!
0*
09
0>
0C
#800790000000
1!
1*
b1 6
19
1>
1C
b1 G
#800800000000
0!
0*
09
0>
0C
#800810000000
1!
1*
b10 6
19
1>
1C
b10 G
#800820000000
0!
0*
09
0>
0C
#800830000000
1!
1*
b11 6
19
1>
1C
b11 G
#800840000000
0!
0*
09
0>
0C
#800850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#800860000000
0!
0*
09
0>
0C
#800870000000
1!
1*
b101 6
19
1>
1C
b101 G
#800880000000
0!
0*
09
0>
0C
#800890000000
1!
1*
b110 6
19
1>
1C
b110 G
#800900000000
0!
0*
09
0>
0C
#800910000000
1!
1*
b111 6
19
1>
1C
b111 G
#800920000000
0!
0*
09
0>
0C
#800930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#800940000000
0!
0*
09
0>
0C
#800950000000
1!
1*
b1 6
19
1>
1C
b1 G
#800960000000
0!
0*
09
0>
0C
#800970000000
1!
1*
b10 6
19
1>
1C
b10 G
#800980000000
0!
0*
09
0>
0C
#800990000000
1!
1*
b11 6
19
1>
1C
b11 G
#801000000000
0!
0*
09
0>
0C
#801010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#801020000000
0!
0*
09
0>
0C
#801030000000
1!
1*
b101 6
19
1>
1C
b101 G
#801040000000
0!
0*
09
0>
0C
#801050000000
1!
1*
b110 6
19
1>
1C
b110 G
#801060000000
0!
0*
09
0>
0C
#801070000000
1!
1*
b111 6
19
1>
1C
b111 G
#801080000000
0!
1"
0*
1+
09
1:
0>
0C
#801090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#801100000000
0!
0*
09
0>
0C
#801110000000
1!
1*
b1 6
19
1>
1C
b1 G
#801120000000
0!
0*
09
0>
0C
#801130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#801140000000
0!
0*
09
0>
0C
#801150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#801160000000
0!
0*
09
0>
0C
#801170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#801180000000
0!
0*
09
0>
0C
#801190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#801200000000
0!
0#
0*
0,
09
0>
0?
0C
#801210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#801220000000
0!
0*
09
0>
0C
#801230000000
1!
1*
19
1>
1C
#801240000000
0!
0*
09
0>
0C
#801250000000
1!
1*
19
1>
1C
#801260000000
0!
0*
09
0>
0C
#801270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#801280000000
0!
0*
09
0>
0C
#801290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#801300000000
0!
0*
09
0>
0C
#801310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#801320000000
0!
0*
09
0>
0C
#801330000000
1!
1*
b10 6
19
1>
1C
b10 G
#801340000000
0!
0*
09
0>
0C
#801350000000
1!
1*
b11 6
19
1>
1C
b11 G
#801360000000
0!
0*
09
0>
0C
#801370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#801380000000
0!
0*
09
0>
0C
#801390000000
1!
1*
b101 6
19
1>
1C
b101 G
#801400000000
0!
0*
09
0>
0C
#801410000000
1!
1*
b110 6
19
1>
1C
b110 G
#801420000000
0!
0*
09
0>
0C
#801430000000
1!
1*
b111 6
19
1>
1C
b111 G
#801440000000
0!
0*
09
0>
0C
#801450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#801460000000
0!
0*
09
0>
0C
#801470000000
1!
1*
b1 6
19
1>
1C
b1 G
#801480000000
0!
0*
09
0>
0C
#801490000000
1!
1*
b10 6
19
1>
1C
b10 G
#801500000000
0!
0*
09
0>
0C
#801510000000
1!
1*
b11 6
19
1>
1C
b11 G
#801520000000
0!
0*
09
0>
0C
#801530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#801540000000
0!
0*
09
0>
0C
#801550000000
1!
1*
b101 6
19
1>
1C
b101 G
#801560000000
0!
0*
09
0>
0C
#801570000000
1!
1*
b110 6
19
1>
1C
b110 G
#801580000000
0!
0*
09
0>
0C
#801590000000
1!
1*
b111 6
19
1>
1C
b111 G
#801600000000
0!
0*
09
0>
0C
#801610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#801620000000
0!
0*
09
0>
0C
#801630000000
1!
1*
b1 6
19
1>
1C
b1 G
#801640000000
0!
0*
09
0>
0C
#801650000000
1!
1*
b10 6
19
1>
1C
b10 G
#801660000000
0!
0*
09
0>
0C
#801670000000
1!
1*
b11 6
19
1>
1C
b11 G
#801680000000
0!
0*
09
0>
0C
#801690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#801700000000
0!
0*
09
0>
0C
#801710000000
1!
1*
b101 6
19
1>
1C
b101 G
#801720000000
0!
0*
09
0>
0C
#801730000000
1!
1*
b110 6
19
1>
1C
b110 G
#801740000000
0!
0*
09
0>
0C
#801750000000
1!
1*
b111 6
19
1>
1C
b111 G
#801760000000
0!
1"
0*
1+
09
1:
0>
0C
#801770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#801780000000
0!
0*
09
0>
0C
#801790000000
1!
1*
b1 6
19
1>
1C
b1 G
#801800000000
0!
0*
09
0>
0C
#801810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#801820000000
0!
0*
09
0>
0C
#801830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#801840000000
0!
0*
09
0>
0C
#801850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#801860000000
0!
0*
09
0>
0C
#801870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#801880000000
0!
0#
0*
0,
09
0>
0?
0C
#801890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#801900000000
0!
0*
09
0>
0C
#801910000000
1!
1*
19
1>
1C
#801920000000
0!
0*
09
0>
0C
#801930000000
1!
1*
19
1>
1C
#801940000000
0!
0*
09
0>
0C
#801950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#801960000000
0!
0*
09
0>
0C
#801970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#801980000000
0!
0*
09
0>
0C
#801990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#802000000000
0!
0*
09
0>
0C
#802010000000
1!
1*
b10 6
19
1>
1C
b10 G
#802020000000
0!
0*
09
0>
0C
#802030000000
1!
1*
b11 6
19
1>
1C
b11 G
#802040000000
0!
0*
09
0>
0C
#802050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#802060000000
0!
0*
09
0>
0C
#802070000000
1!
1*
b101 6
19
1>
1C
b101 G
#802080000000
0!
0*
09
0>
0C
#802090000000
1!
1*
b110 6
19
1>
1C
b110 G
#802100000000
0!
0*
09
0>
0C
#802110000000
1!
1*
b111 6
19
1>
1C
b111 G
#802120000000
0!
0*
09
0>
0C
#802130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#802140000000
0!
0*
09
0>
0C
#802150000000
1!
1*
b1 6
19
1>
1C
b1 G
#802160000000
0!
0*
09
0>
0C
#802170000000
1!
1*
b10 6
19
1>
1C
b10 G
#802180000000
0!
0*
09
0>
0C
#802190000000
1!
1*
b11 6
19
1>
1C
b11 G
#802200000000
0!
0*
09
0>
0C
#802210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#802220000000
0!
0*
09
0>
0C
#802230000000
1!
1*
b101 6
19
1>
1C
b101 G
#802240000000
0!
0*
09
0>
0C
#802250000000
1!
1*
b110 6
19
1>
1C
b110 G
#802260000000
0!
0*
09
0>
0C
#802270000000
1!
1*
b111 6
19
1>
1C
b111 G
#802280000000
0!
0*
09
0>
0C
#802290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#802300000000
0!
0*
09
0>
0C
#802310000000
1!
1*
b1 6
19
1>
1C
b1 G
#802320000000
0!
0*
09
0>
0C
#802330000000
1!
1*
b10 6
19
1>
1C
b10 G
#802340000000
0!
0*
09
0>
0C
#802350000000
1!
1*
b11 6
19
1>
1C
b11 G
#802360000000
0!
0*
09
0>
0C
#802370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#802380000000
0!
0*
09
0>
0C
#802390000000
1!
1*
b101 6
19
1>
1C
b101 G
#802400000000
0!
0*
09
0>
0C
#802410000000
1!
1*
b110 6
19
1>
1C
b110 G
#802420000000
0!
0*
09
0>
0C
#802430000000
1!
1*
b111 6
19
1>
1C
b111 G
#802440000000
0!
1"
0*
1+
09
1:
0>
0C
#802450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#802460000000
0!
0*
09
0>
0C
#802470000000
1!
1*
b1 6
19
1>
1C
b1 G
#802480000000
0!
0*
09
0>
0C
#802490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#802500000000
0!
0*
09
0>
0C
#802510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#802520000000
0!
0*
09
0>
0C
#802530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#802540000000
0!
0*
09
0>
0C
#802550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#802560000000
0!
0#
0*
0,
09
0>
0?
0C
#802570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#802580000000
0!
0*
09
0>
0C
#802590000000
1!
1*
19
1>
1C
#802600000000
0!
0*
09
0>
0C
#802610000000
1!
1*
19
1>
1C
#802620000000
0!
0*
09
0>
0C
#802630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#802640000000
0!
0*
09
0>
0C
#802650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#802660000000
0!
0*
09
0>
0C
#802670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#802680000000
0!
0*
09
0>
0C
#802690000000
1!
1*
b10 6
19
1>
1C
b10 G
#802700000000
0!
0*
09
0>
0C
#802710000000
1!
1*
b11 6
19
1>
1C
b11 G
#802720000000
0!
0*
09
0>
0C
#802730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#802740000000
0!
0*
09
0>
0C
#802750000000
1!
1*
b101 6
19
1>
1C
b101 G
#802760000000
0!
0*
09
0>
0C
#802770000000
1!
1*
b110 6
19
1>
1C
b110 G
#802780000000
0!
0*
09
0>
0C
#802790000000
1!
1*
b111 6
19
1>
1C
b111 G
#802800000000
0!
0*
09
0>
0C
#802810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#802820000000
0!
0*
09
0>
0C
#802830000000
1!
1*
b1 6
19
1>
1C
b1 G
#802840000000
0!
0*
09
0>
0C
#802850000000
1!
1*
b10 6
19
1>
1C
b10 G
#802860000000
0!
0*
09
0>
0C
#802870000000
1!
1*
b11 6
19
1>
1C
b11 G
#802880000000
0!
0*
09
0>
0C
#802890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#802900000000
0!
0*
09
0>
0C
#802910000000
1!
1*
b101 6
19
1>
1C
b101 G
#802920000000
0!
0*
09
0>
0C
#802930000000
1!
1*
b110 6
19
1>
1C
b110 G
#802940000000
0!
0*
09
0>
0C
#802950000000
1!
1*
b111 6
19
1>
1C
b111 G
#802960000000
0!
0*
09
0>
0C
#802970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#802980000000
0!
0*
09
0>
0C
#802990000000
1!
1*
b1 6
19
1>
1C
b1 G
#803000000000
0!
0*
09
0>
0C
#803010000000
1!
1*
b10 6
19
1>
1C
b10 G
#803020000000
0!
0*
09
0>
0C
#803030000000
1!
1*
b11 6
19
1>
1C
b11 G
#803040000000
0!
0*
09
0>
0C
#803050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#803060000000
0!
0*
09
0>
0C
#803070000000
1!
1*
b101 6
19
1>
1C
b101 G
#803080000000
0!
0*
09
0>
0C
#803090000000
1!
1*
b110 6
19
1>
1C
b110 G
#803100000000
0!
0*
09
0>
0C
#803110000000
1!
1*
b111 6
19
1>
1C
b111 G
#803120000000
0!
1"
0*
1+
09
1:
0>
0C
#803130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#803140000000
0!
0*
09
0>
0C
#803150000000
1!
1*
b1 6
19
1>
1C
b1 G
#803160000000
0!
0*
09
0>
0C
#803170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#803180000000
0!
0*
09
0>
0C
#803190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#803200000000
0!
0*
09
0>
0C
#803210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#803220000000
0!
0*
09
0>
0C
#803230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#803240000000
0!
0#
0*
0,
09
0>
0?
0C
#803250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#803260000000
0!
0*
09
0>
0C
#803270000000
1!
1*
19
1>
1C
#803280000000
0!
0*
09
0>
0C
#803290000000
1!
1*
19
1>
1C
#803300000000
0!
0*
09
0>
0C
#803310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#803320000000
0!
0*
09
0>
0C
#803330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#803340000000
0!
0*
09
0>
0C
#803350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#803360000000
0!
0*
09
0>
0C
#803370000000
1!
1*
b10 6
19
1>
1C
b10 G
#803380000000
0!
0*
09
0>
0C
#803390000000
1!
1*
b11 6
19
1>
1C
b11 G
#803400000000
0!
0*
09
0>
0C
#803410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#803420000000
0!
0*
09
0>
0C
#803430000000
1!
1*
b101 6
19
1>
1C
b101 G
#803440000000
0!
0*
09
0>
0C
#803450000000
1!
1*
b110 6
19
1>
1C
b110 G
#803460000000
0!
0*
09
0>
0C
#803470000000
1!
1*
b111 6
19
1>
1C
b111 G
#803480000000
0!
0*
09
0>
0C
#803490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#803500000000
0!
0*
09
0>
0C
#803510000000
1!
1*
b1 6
19
1>
1C
b1 G
#803520000000
0!
0*
09
0>
0C
#803530000000
1!
1*
b10 6
19
1>
1C
b10 G
#803540000000
0!
0*
09
0>
0C
#803550000000
1!
1*
b11 6
19
1>
1C
b11 G
#803560000000
0!
0*
09
0>
0C
#803570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#803580000000
0!
0*
09
0>
0C
#803590000000
1!
1*
b101 6
19
1>
1C
b101 G
#803600000000
0!
0*
09
0>
0C
#803610000000
1!
1*
b110 6
19
1>
1C
b110 G
#803620000000
0!
0*
09
0>
0C
#803630000000
1!
1*
b111 6
19
1>
1C
b111 G
#803640000000
0!
0*
09
0>
0C
#803650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#803660000000
0!
0*
09
0>
0C
#803670000000
1!
1*
b1 6
19
1>
1C
b1 G
#803680000000
0!
0*
09
0>
0C
#803690000000
1!
1*
b10 6
19
1>
1C
b10 G
#803700000000
0!
0*
09
0>
0C
#803710000000
1!
1*
b11 6
19
1>
1C
b11 G
#803720000000
0!
0*
09
0>
0C
#803730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#803740000000
0!
0*
09
0>
0C
#803750000000
1!
1*
b101 6
19
1>
1C
b101 G
#803760000000
0!
0*
09
0>
0C
#803770000000
1!
1*
b110 6
19
1>
1C
b110 G
#803780000000
0!
0*
09
0>
0C
#803790000000
1!
1*
b111 6
19
1>
1C
b111 G
#803800000000
0!
1"
0*
1+
09
1:
0>
0C
#803810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#803820000000
0!
0*
09
0>
0C
#803830000000
1!
1*
b1 6
19
1>
1C
b1 G
#803840000000
0!
0*
09
0>
0C
#803850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#803860000000
0!
0*
09
0>
0C
#803870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#803880000000
0!
0*
09
0>
0C
#803890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#803900000000
0!
0*
09
0>
0C
#803910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#803920000000
0!
0#
0*
0,
09
0>
0?
0C
#803930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#803940000000
0!
0*
09
0>
0C
#803950000000
1!
1*
19
1>
1C
#803960000000
0!
0*
09
0>
0C
#803970000000
1!
1*
19
1>
1C
#803980000000
0!
0*
09
0>
0C
#803990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#804000000000
0!
0*
09
0>
0C
#804010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#804020000000
0!
0*
09
0>
0C
#804030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#804040000000
0!
0*
09
0>
0C
#804050000000
1!
1*
b10 6
19
1>
1C
b10 G
#804060000000
0!
0*
09
0>
0C
#804070000000
1!
1*
b11 6
19
1>
1C
b11 G
#804080000000
0!
0*
09
0>
0C
#804090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#804100000000
0!
0*
09
0>
0C
#804110000000
1!
1*
b101 6
19
1>
1C
b101 G
#804120000000
0!
0*
09
0>
0C
#804130000000
1!
1*
b110 6
19
1>
1C
b110 G
#804140000000
0!
0*
09
0>
0C
#804150000000
1!
1*
b111 6
19
1>
1C
b111 G
#804160000000
0!
0*
09
0>
0C
#804170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#804180000000
0!
0*
09
0>
0C
#804190000000
1!
1*
b1 6
19
1>
1C
b1 G
#804200000000
0!
0*
09
0>
0C
#804210000000
1!
1*
b10 6
19
1>
1C
b10 G
#804220000000
0!
0*
09
0>
0C
#804230000000
1!
1*
b11 6
19
1>
1C
b11 G
#804240000000
0!
0*
09
0>
0C
#804250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#804260000000
0!
0*
09
0>
0C
#804270000000
1!
1*
b101 6
19
1>
1C
b101 G
#804280000000
0!
0*
09
0>
0C
#804290000000
1!
1*
b110 6
19
1>
1C
b110 G
#804300000000
0!
0*
09
0>
0C
#804310000000
1!
1*
b111 6
19
1>
1C
b111 G
#804320000000
0!
0*
09
0>
0C
#804330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#804340000000
0!
0*
09
0>
0C
#804350000000
1!
1*
b1 6
19
1>
1C
b1 G
#804360000000
0!
0*
09
0>
0C
#804370000000
1!
1*
b10 6
19
1>
1C
b10 G
#804380000000
0!
0*
09
0>
0C
#804390000000
1!
1*
b11 6
19
1>
1C
b11 G
#804400000000
0!
0*
09
0>
0C
#804410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#804420000000
0!
0*
09
0>
0C
#804430000000
1!
1*
b101 6
19
1>
1C
b101 G
#804440000000
0!
0*
09
0>
0C
#804450000000
1!
1*
b110 6
19
1>
1C
b110 G
#804460000000
0!
0*
09
0>
0C
#804470000000
1!
1*
b111 6
19
1>
1C
b111 G
#804480000000
0!
1"
0*
1+
09
1:
0>
0C
#804490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#804500000000
0!
0*
09
0>
0C
#804510000000
1!
1*
b1 6
19
1>
1C
b1 G
#804520000000
0!
0*
09
0>
0C
#804530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#804540000000
0!
0*
09
0>
0C
#804550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#804560000000
0!
0*
09
0>
0C
#804570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#804580000000
0!
0*
09
0>
0C
#804590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#804600000000
0!
0#
0*
0,
09
0>
0?
0C
#804610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#804620000000
0!
0*
09
0>
0C
#804630000000
1!
1*
19
1>
1C
#804640000000
0!
0*
09
0>
0C
#804650000000
1!
1*
19
1>
1C
#804660000000
0!
0*
09
0>
0C
#804670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#804680000000
0!
0*
09
0>
0C
#804690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#804700000000
0!
0*
09
0>
0C
#804710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#804720000000
0!
0*
09
0>
0C
#804730000000
1!
1*
b10 6
19
1>
1C
b10 G
#804740000000
0!
0*
09
0>
0C
#804750000000
1!
1*
b11 6
19
1>
1C
b11 G
#804760000000
0!
0*
09
0>
0C
#804770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#804780000000
0!
0*
09
0>
0C
#804790000000
1!
1*
b101 6
19
1>
1C
b101 G
#804800000000
0!
0*
09
0>
0C
#804810000000
1!
1*
b110 6
19
1>
1C
b110 G
#804820000000
0!
0*
09
0>
0C
#804830000000
1!
1*
b111 6
19
1>
1C
b111 G
#804840000000
0!
0*
09
0>
0C
#804850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#804860000000
0!
0*
09
0>
0C
#804870000000
1!
1*
b1 6
19
1>
1C
b1 G
#804880000000
0!
0*
09
0>
0C
#804890000000
1!
1*
b10 6
19
1>
1C
b10 G
#804900000000
0!
0*
09
0>
0C
#804910000000
1!
1*
b11 6
19
1>
1C
b11 G
#804920000000
0!
0*
09
0>
0C
#804930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#804940000000
0!
0*
09
0>
0C
#804950000000
1!
1*
b101 6
19
1>
1C
b101 G
#804960000000
0!
0*
09
0>
0C
#804970000000
1!
1*
b110 6
19
1>
1C
b110 G
#804980000000
0!
0*
09
0>
0C
#804990000000
1!
1*
b111 6
19
1>
1C
b111 G
#805000000000
0!
0*
09
0>
0C
#805010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#805020000000
0!
0*
09
0>
0C
#805030000000
1!
1*
b1 6
19
1>
1C
b1 G
#805040000000
0!
0*
09
0>
0C
#805050000000
1!
1*
b10 6
19
1>
1C
b10 G
#805060000000
0!
0*
09
0>
0C
#805070000000
1!
1*
b11 6
19
1>
1C
b11 G
#805080000000
0!
0*
09
0>
0C
#805090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#805100000000
0!
0*
09
0>
0C
#805110000000
1!
1*
b101 6
19
1>
1C
b101 G
#805120000000
0!
0*
09
0>
0C
#805130000000
1!
1*
b110 6
19
1>
1C
b110 G
#805140000000
0!
0*
09
0>
0C
#805150000000
1!
1*
b111 6
19
1>
1C
b111 G
#805160000000
0!
1"
0*
1+
09
1:
0>
0C
#805170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#805180000000
0!
0*
09
0>
0C
#805190000000
1!
1*
b1 6
19
1>
1C
b1 G
#805200000000
0!
0*
09
0>
0C
#805210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#805220000000
0!
0*
09
0>
0C
#805230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#805240000000
0!
0*
09
0>
0C
#805250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#805260000000
0!
0*
09
0>
0C
#805270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#805280000000
0!
0#
0*
0,
09
0>
0?
0C
#805290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#805300000000
0!
0*
09
0>
0C
#805310000000
1!
1*
19
1>
1C
#805320000000
0!
0*
09
0>
0C
#805330000000
1!
1*
19
1>
1C
#805340000000
0!
0*
09
0>
0C
#805350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#805360000000
0!
0*
09
0>
0C
#805370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#805380000000
0!
0*
09
0>
0C
#805390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#805400000000
0!
0*
09
0>
0C
#805410000000
1!
1*
b10 6
19
1>
1C
b10 G
#805420000000
0!
0*
09
0>
0C
#805430000000
1!
1*
b11 6
19
1>
1C
b11 G
#805440000000
0!
0*
09
0>
0C
#805450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#805460000000
0!
0*
09
0>
0C
#805470000000
1!
1*
b101 6
19
1>
1C
b101 G
#805480000000
0!
0*
09
0>
0C
#805490000000
1!
1*
b110 6
19
1>
1C
b110 G
#805500000000
0!
0*
09
0>
0C
#805510000000
1!
1*
b111 6
19
1>
1C
b111 G
#805520000000
0!
0*
09
0>
0C
#805530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#805540000000
0!
0*
09
0>
0C
#805550000000
1!
1*
b1 6
19
1>
1C
b1 G
#805560000000
0!
0*
09
0>
0C
#805570000000
1!
1*
b10 6
19
1>
1C
b10 G
#805580000000
0!
0*
09
0>
0C
#805590000000
1!
1*
b11 6
19
1>
1C
b11 G
#805600000000
0!
0*
09
0>
0C
#805610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#805620000000
0!
0*
09
0>
0C
#805630000000
1!
1*
b101 6
19
1>
1C
b101 G
#805640000000
0!
0*
09
0>
0C
#805650000000
1!
1*
b110 6
19
1>
1C
b110 G
#805660000000
0!
0*
09
0>
0C
#805670000000
1!
1*
b111 6
19
1>
1C
b111 G
#805680000000
0!
0*
09
0>
0C
#805690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#805700000000
0!
0*
09
0>
0C
#805710000000
1!
1*
b1 6
19
1>
1C
b1 G
#805720000000
0!
0*
09
0>
0C
#805730000000
1!
1*
b10 6
19
1>
1C
b10 G
#805740000000
0!
0*
09
0>
0C
#805750000000
1!
1*
b11 6
19
1>
1C
b11 G
#805760000000
0!
0*
09
0>
0C
#805770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#805780000000
0!
0*
09
0>
0C
#805790000000
1!
1*
b101 6
19
1>
1C
b101 G
#805800000000
0!
0*
09
0>
0C
#805810000000
1!
1*
b110 6
19
1>
1C
b110 G
#805820000000
0!
0*
09
0>
0C
#805830000000
1!
1*
b111 6
19
1>
1C
b111 G
#805840000000
0!
1"
0*
1+
09
1:
0>
0C
#805850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#805860000000
0!
0*
09
0>
0C
#805870000000
1!
1*
b1 6
19
1>
1C
b1 G
#805880000000
0!
0*
09
0>
0C
#805890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#805900000000
0!
0*
09
0>
0C
#805910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#805920000000
0!
0*
09
0>
0C
#805930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#805940000000
0!
0*
09
0>
0C
#805950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#805960000000
0!
0#
0*
0,
09
0>
0?
0C
#805970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#805980000000
0!
0*
09
0>
0C
#805990000000
1!
1*
19
1>
1C
#806000000000
0!
0*
09
0>
0C
#806010000000
1!
1*
19
1>
1C
#806020000000
0!
0*
09
0>
0C
#806030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#806040000000
0!
0*
09
0>
0C
#806050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#806060000000
0!
0*
09
0>
0C
#806070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#806080000000
0!
0*
09
0>
0C
#806090000000
1!
1*
b10 6
19
1>
1C
b10 G
#806100000000
0!
0*
09
0>
0C
#806110000000
1!
1*
b11 6
19
1>
1C
b11 G
#806120000000
0!
0*
09
0>
0C
#806130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#806140000000
0!
0*
09
0>
0C
#806150000000
1!
1*
b101 6
19
1>
1C
b101 G
#806160000000
0!
0*
09
0>
0C
#806170000000
1!
1*
b110 6
19
1>
1C
b110 G
#806180000000
0!
0*
09
0>
0C
#806190000000
1!
1*
b111 6
19
1>
1C
b111 G
#806200000000
0!
0*
09
0>
0C
#806210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#806220000000
0!
0*
09
0>
0C
#806230000000
1!
1*
b1 6
19
1>
1C
b1 G
#806240000000
0!
0*
09
0>
0C
#806250000000
1!
1*
b10 6
19
1>
1C
b10 G
#806260000000
0!
0*
09
0>
0C
#806270000000
1!
1*
b11 6
19
1>
1C
b11 G
#806280000000
0!
0*
09
0>
0C
#806290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#806300000000
0!
0*
09
0>
0C
#806310000000
1!
1*
b101 6
19
1>
1C
b101 G
#806320000000
0!
0*
09
0>
0C
#806330000000
1!
1*
b110 6
19
1>
1C
b110 G
#806340000000
0!
0*
09
0>
0C
#806350000000
1!
1*
b111 6
19
1>
1C
b111 G
#806360000000
0!
0*
09
0>
0C
#806370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#806380000000
0!
0*
09
0>
0C
#806390000000
1!
1*
b1 6
19
1>
1C
b1 G
#806400000000
0!
0*
09
0>
0C
#806410000000
1!
1*
b10 6
19
1>
1C
b10 G
#806420000000
0!
0*
09
0>
0C
#806430000000
1!
1*
b11 6
19
1>
1C
b11 G
#806440000000
0!
0*
09
0>
0C
#806450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#806460000000
0!
0*
09
0>
0C
#806470000000
1!
1*
b101 6
19
1>
1C
b101 G
#806480000000
0!
0*
09
0>
0C
#806490000000
1!
1*
b110 6
19
1>
1C
b110 G
#806500000000
0!
0*
09
0>
0C
#806510000000
1!
1*
b111 6
19
1>
1C
b111 G
#806520000000
0!
1"
0*
1+
09
1:
0>
0C
#806530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#806540000000
0!
0*
09
0>
0C
#806550000000
1!
1*
b1 6
19
1>
1C
b1 G
#806560000000
0!
0*
09
0>
0C
#806570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#806580000000
0!
0*
09
0>
0C
#806590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#806600000000
0!
0*
09
0>
0C
#806610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#806620000000
0!
0*
09
0>
0C
#806630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#806640000000
0!
0#
0*
0,
09
0>
0?
0C
#806650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#806660000000
0!
0*
09
0>
0C
#806670000000
1!
1*
19
1>
1C
#806680000000
0!
0*
09
0>
0C
#806690000000
1!
1*
19
1>
1C
#806700000000
0!
0*
09
0>
0C
#806710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#806720000000
0!
0*
09
0>
0C
#806730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#806740000000
0!
0*
09
0>
0C
#806750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#806760000000
0!
0*
09
0>
0C
#806770000000
1!
1*
b10 6
19
1>
1C
b10 G
#806780000000
0!
0*
09
0>
0C
#806790000000
1!
1*
b11 6
19
1>
1C
b11 G
#806800000000
0!
0*
09
0>
0C
#806810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#806820000000
0!
0*
09
0>
0C
#806830000000
1!
1*
b101 6
19
1>
1C
b101 G
#806840000000
0!
0*
09
0>
0C
#806850000000
1!
1*
b110 6
19
1>
1C
b110 G
#806860000000
0!
0*
09
0>
0C
#806870000000
1!
1*
b111 6
19
1>
1C
b111 G
#806880000000
0!
0*
09
0>
0C
#806890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#806900000000
0!
0*
09
0>
0C
#806910000000
1!
1*
b1 6
19
1>
1C
b1 G
#806920000000
0!
0*
09
0>
0C
#806930000000
1!
1*
b10 6
19
1>
1C
b10 G
#806940000000
0!
0*
09
0>
0C
#806950000000
1!
1*
b11 6
19
1>
1C
b11 G
#806960000000
0!
0*
09
0>
0C
#806970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#806980000000
0!
0*
09
0>
0C
#806990000000
1!
1*
b101 6
19
1>
1C
b101 G
#807000000000
0!
0*
09
0>
0C
#807010000000
1!
1*
b110 6
19
1>
1C
b110 G
#807020000000
0!
0*
09
0>
0C
#807030000000
1!
1*
b111 6
19
1>
1C
b111 G
#807040000000
0!
0*
09
0>
0C
#807050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#807060000000
0!
0*
09
0>
0C
#807070000000
1!
1*
b1 6
19
1>
1C
b1 G
#807080000000
0!
0*
09
0>
0C
#807090000000
1!
1*
b10 6
19
1>
1C
b10 G
#807100000000
0!
0*
09
0>
0C
#807110000000
1!
1*
b11 6
19
1>
1C
b11 G
#807120000000
0!
0*
09
0>
0C
#807130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#807140000000
0!
0*
09
0>
0C
#807150000000
1!
1*
b101 6
19
1>
1C
b101 G
#807160000000
0!
0*
09
0>
0C
#807170000000
1!
1*
b110 6
19
1>
1C
b110 G
#807180000000
0!
0*
09
0>
0C
#807190000000
1!
1*
b111 6
19
1>
1C
b111 G
#807200000000
0!
1"
0*
1+
09
1:
0>
0C
#807210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#807220000000
0!
0*
09
0>
0C
#807230000000
1!
1*
b1 6
19
1>
1C
b1 G
#807240000000
0!
0*
09
0>
0C
#807250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#807260000000
0!
0*
09
0>
0C
#807270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#807280000000
0!
0*
09
0>
0C
#807290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#807300000000
0!
0*
09
0>
0C
#807310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#807320000000
0!
0#
0*
0,
09
0>
0?
0C
#807330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#807340000000
0!
0*
09
0>
0C
#807350000000
1!
1*
19
1>
1C
#807360000000
0!
0*
09
0>
0C
#807370000000
1!
1*
19
1>
1C
#807380000000
0!
0*
09
0>
0C
#807390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#807400000000
0!
0*
09
0>
0C
#807410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#807420000000
0!
0*
09
0>
0C
#807430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#807440000000
0!
0*
09
0>
0C
#807450000000
1!
1*
b10 6
19
1>
1C
b10 G
#807460000000
0!
0*
09
0>
0C
#807470000000
1!
1*
b11 6
19
1>
1C
b11 G
#807480000000
0!
0*
09
0>
0C
#807490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#807500000000
0!
0*
09
0>
0C
#807510000000
1!
1*
b101 6
19
1>
1C
b101 G
#807520000000
0!
0*
09
0>
0C
#807530000000
1!
1*
b110 6
19
1>
1C
b110 G
#807540000000
0!
0*
09
0>
0C
#807550000000
1!
1*
b111 6
19
1>
1C
b111 G
#807560000000
0!
0*
09
0>
0C
#807570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#807580000000
0!
0*
09
0>
0C
#807590000000
1!
1*
b1 6
19
1>
1C
b1 G
#807600000000
0!
0*
09
0>
0C
#807610000000
1!
1*
b10 6
19
1>
1C
b10 G
#807620000000
0!
0*
09
0>
0C
#807630000000
1!
1*
b11 6
19
1>
1C
b11 G
#807640000000
0!
0*
09
0>
0C
#807650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#807660000000
0!
0*
09
0>
0C
#807670000000
1!
1*
b101 6
19
1>
1C
b101 G
#807680000000
0!
0*
09
0>
0C
#807690000000
1!
1*
b110 6
19
1>
1C
b110 G
#807700000000
0!
0*
09
0>
0C
#807710000000
1!
1*
b111 6
19
1>
1C
b111 G
#807720000000
0!
0*
09
0>
0C
#807730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#807740000000
0!
0*
09
0>
0C
#807750000000
1!
1*
b1 6
19
1>
1C
b1 G
#807760000000
0!
0*
09
0>
0C
#807770000000
1!
1*
b10 6
19
1>
1C
b10 G
#807780000000
0!
0*
09
0>
0C
#807790000000
1!
1*
b11 6
19
1>
1C
b11 G
#807800000000
0!
0*
09
0>
0C
#807810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#807820000000
0!
0*
09
0>
0C
#807830000000
1!
1*
b101 6
19
1>
1C
b101 G
#807840000000
0!
0*
09
0>
0C
#807850000000
1!
1*
b110 6
19
1>
1C
b110 G
#807860000000
0!
0*
09
0>
0C
#807870000000
1!
1*
b111 6
19
1>
1C
b111 G
#807880000000
0!
1"
0*
1+
09
1:
0>
0C
#807890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#807900000000
0!
0*
09
0>
0C
#807910000000
1!
1*
b1 6
19
1>
1C
b1 G
#807920000000
0!
0*
09
0>
0C
#807930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#807940000000
0!
0*
09
0>
0C
#807950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#807960000000
0!
0*
09
0>
0C
#807970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#807980000000
0!
0*
09
0>
0C
#807990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#808000000000
0!
0#
0*
0,
09
0>
0?
0C
#808010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#808020000000
0!
0*
09
0>
0C
#808030000000
1!
1*
19
1>
1C
#808040000000
0!
0*
09
0>
0C
#808050000000
1!
1*
19
1>
1C
#808060000000
0!
0*
09
0>
0C
#808070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#808080000000
0!
0*
09
0>
0C
#808090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#808100000000
0!
0*
09
0>
0C
#808110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#808120000000
0!
0*
09
0>
0C
#808130000000
1!
1*
b10 6
19
1>
1C
b10 G
#808140000000
0!
0*
09
0>
0C
#808150000000
1!
1*
b11 6
19
1>
1C
b11 G
#808160000000
0!
0*
09
0>
0C
#808170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#808180000000
0!
0*
09
0>
0C
#808190000000
1!
1*
b101 6
19
1>
1C
b101 G
#808200000000
0!
0*
09
0>
0C
#808210000000
1!
1*
b110 6
19
1>
1C
b110 G
#808220000000
0!
0*
09
0>
0C
#808230000000
1!
1*
b111 6
19
1>
1C
b111 G
#808240000000
0!
0*
09
0>
0C
#808250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#808260000000
0!
0*
09
0>
0C
#808270000000
1!
1*
b1 6
19
1>
1C
b1 G
#808280000000
0!
0*
09
0>
0C
#808290000000
1!
1*
b10 6
19
1>
1C
b10 G
#808300000000
0!
0*
09
0>
0C
#808310000000
1!
1*
b11 6
19
1>
1C
b11 G
#808320000000
0!
0*
09
0>
0C
#808330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#808340000000
0!
0*
09
0>
0C
#808350000000
1!
1*
b101 6
19
1>
1C
b101 G
#808360000000
0!
0*
09
0>
0C
#808370000000
1!
1*
b110 6
19
1>
1C
b110 G
#808380000000
0!
0*
09
0>
0C
#808390000000
1!
1*
b111 6
19
1>
1C
b111 G
#808400000000
0!
0*
09
0>
0C
#808410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#808420000000
0!
0*
09
0>
0C
#808430000000
1!
1*
b1 6
19
1>
1C
b1 G
#808440000000
0!
0*
09
0>
0C
#808450000000
1!
1*
b10 6
19
1>
1C
b10 G
#808460000000
0!
0*
09
0>
0C
#808470000000
1!
1*
b11 6
19
1>
1C
b11 G
#808480000000
0!
0*
09
0>
0C
#808490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#808500000000
0!
0*
09
0>
0C
#808510000000
1!
1*
b101 6
19
1>
1C
b101 G
#808520000000
0!
0*
09
0>
0C
#808530000000
1!
1*
b110 6
19
1>
1C
b110 G
#808540000000
0!
0*
09
0>
0C
#808550000000
1!
1*
b111 6
19
1>
1C
b111 G
#808560000000
0!
1"
0*
1+
09
1:
0>
0C
#808570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#808580000000
0!
0*
09
0>
0C
#808590000000
1!
1*
b1 6
19
1>
1C
b1 G
#808600000000
0!
0*
09
0>
0C
#808610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#808620000000
0!
0*
09
0>
0C
#808630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#808640000000
0!
0*
09
0>
0C
#808650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#808660000000
0!
0*
09
0>
0C
#808670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#808680000000
0!
0#
0*
0,
09
0>
0?
0C
#808690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#808700000000
0!
0*
09
0>
0C
#808710000000
1!
1*
19
1>
1C
#808720000000
0!
0*
09
0>
0C
#808730000000
1!
1*
19
1>
1C
#808740000000
0!
0*
09
0>
0C
#808750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#808760000000
0!
0*
09
0>
0C
#808770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#808780000000
0!
0*
09
0>
0C
#808790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#808800000000
0!
0*
09
0>
0C
#808810000000
1!
1*
b10 6
19
1>
1C
b10 G
#808820000000
0!
0*
09
0>
0C
#808830000000
1!
1*
b11 6
19
1>
1C
b11 G
#808840000000
0!
0*
09
0>
0C
#808850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#808860000000
0!
0*
09
0>
0C
#808870000000
1!
1*
b101 6
19
1>
1C
b101 G
#808880000000
0!
0*
09
0>
0C
#808890000000
1!
1*
b110 6
19
1>
1C
b110 G
#808900000000
0!
0*
09
0>
0C
#808910000000
1!
1*
b111 6
19
1>
1C
b111 G
#808920000000
0!
0*
09
0>
0C
#808930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#808940000000
0!
0*
09
0>
0C
#808950000000
1!
1*
b1 6
19
1>
1C
b1 G
#808960000000
0!
0*
09
0>
0C
#808970000000
1!
1*
b10 6
19
1>
1C
b10 G
#808980000000
0!
0*
09
0>
0C
#808990000000
1!
1*
b11 6
19
1>
1C
b11 G
#809000000000
0!
0*
09
0>
0C
#809010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#809020000000
0!
0*
09
0>
0C
#809030000000
1!
1*
b101 6
19
1>
1C
b101 G
#809040000000
0!
0*
09
0>
0C
#809050000000
1!
1*
b110 6
19
1>
1C
b110 G
#809060000000
0!
0*
09
0>
0C
#809070000000
1!
1*
b111 6
19
1>
1C
b111 G
#809080000000
0!
0*
09
0>
0C
#809090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#809100000000
0!
0*
09
0>
0C
#809110000000
1!
1*
b1 6
19
1>
1C
b1 G
#809120000000
0!
0*
09
0>
0C
#809130000000
1!
1*
b10 6
19
1>
1C
b10 G
#809140000000
0!
0*
09
0>
0C
#809150000000
1!
1*
b11 6
19
1>
1C
b11 G
#809160000000
0!
0*
09
0>
0C
#809170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#809180000000
0!
0*
09
0>
0C
#809190000000
1!
1*
b101 6
19
1>
1C
b101 G
#809200000000
0!
0*
09
0>
0C
#809210000000
1!
1*
b110 6
19
1>
1C
b110 G
#809220000000
0!
0*
09
0>
0C
#809230000000
1!
1*
b111 6
19
1>
1C
b111 G
#809240000000
0!
1"
0*
1+
09
1:
0>
0C
#809250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#809260000000
0!
0*
09
0>
0C
#809270000000
1!
1*
b1 6
19
1>
1C
b1 G
#809280000000
0!
0*
09
0>
0C
#809290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#809300000000
0!
0*
09
0>
0C
#809310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#809320000000
0!
0*
09
0>
0C
#809330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#809340000000
0!
0*
09
0>
0C
#809350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#809360000000
0!
0#
0*
0,
09
0>
0?
0C
#809370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#809380000000
0!
0*
09
0>
0C
#809390000000
1!
1*
19
1>
1C
#809400000000
0!
0*
09
0>
0C
#809410000000
1!
1*
19
1>
1C
#809420000000
0!
0*
09
0>
0C
#809430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#809440000000
0!
0*
09
0>
0C
#809450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#809460000000
0!
0*
09
0>
0C
#809470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#809480000000
0!
0*
09
0>
0C
#809490000000
1!
1*
b10 6
19
1>
1C
b10 G
#809500000000
0!
0*
09
0>
0C
#809510000000
1!
1*
b11 6
19
1>
1C
b11 G
#809520000000
0!
0*
09
0>
0C
#809530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#809540000000
0!
0*
09
0>
0C
#809550000000
1!
1*
b101 6
19
1>
1C
b101 G
#809560000000
0!
0*
09
0>
0C
#809570000000
1!
1*
b110 6
19
1>
1C
b110 G
#809580000000
0!
0*
09
0>
0C
#809590000000
1!
1*
b111 6
19
1>
1C
b111 G
#809600000000
0!
0*
09
0>
0C
#809610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#809620000000
0!
0*
09
0>
0C
#809630000000
1!
1*
b1 6
19
1>
1C
b1 G
#809640000000
0!
0*
09
0>
0C
#809650000000
1!
1*
b10 6
19
1>
1C
b10 G
#809660000000
0!
0*
09
0>
0C
#809670000000
1!
1*
b11 6
19
1>
1C
b11 G
#809680000000
0!
0*
09
0>
0C
#809690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#809700000000
0!
0*
09
0>
0C
#809710000000
1!
1*
b101 6
19
1>
1C
b101 G
#809720000000
0!
0*
09
0>
0C
#809730000000
1!
1*
b110 6
19
1>
1C
b110 G
#809740000000
0!
0*
09
0>
0C
#809750000000
1!
1*
b111 6
19
1>
1C
b111 G
#809760000000
0!
0*
09
0>
0C
#809770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#809780000000
0!
0*
09
0>
0C
#809790000000
1!
1*
b1 6
19
1>
1C
b1 G
#809800000000
0!
0*
09
0>
0C
#809810000000
1!
1*
b10 6
19
1>
1C
b10 G
#809820000000
0!
0*
09
0>
0C
#809830000000
1!
1*
b11 6
19
1>
1C
b11 G
#809840000000
0!
0*
09
0>
0C
#809850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#809860000000
0!
0*
09
0>
0C
#809870000000
1!
1*
b101 6
19
1>
1C
b101 G
#809880000000
0!
0*
09
0>
0C
#809890000000
1!
1*
b110 6
19
1>
1C
b110 G
#809900000000
0!
0*
09
0>
0C
#809910000000
1!
1*
b111 6
19
1>
1C
b111 G
#809920000000
0!
1"
0*
1+
09
1:
0>
0C
#809930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#809940000000
0!
0*
09
0>
0C
#809950000000
1!
1*
b1 6
19
1>
1C
b1 G
#809960000000
0!
0*
09
0>
0C
#809970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#809980000000
0!
0*
09
0>
0C
#809990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#810000000000
0!
0*
09
0>
0C
#810010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#810020000000
0!
0*
09
0>
0C
#810030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#810040000000
0!
0#
0*
0,
09
0>
0?
0C
#810050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#810060000000
0!
0*
09
0>
0C
#810070000000
1!
1*
19
1>
1C
#810080000000
0!
0*
09
0>
0C
#810090000000
1!
1*
19
1>
1C
#810100000000
0!
0*
09
0>
0C
#810110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#810120000000
0!
0*
09
0>
0C
#810130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#810140000000
0!
0*
09
0>
0C
#810150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#810160000000
0!
0*
09
0>
0C
#810170000000
1!
1*
b10 6
19
1>
1C
b10 G
#810180000000
0!
0*
09
0>
0C
#810190000000
1!
1*
b11 6
19
1>
1C
b11 G
#810200000000
0!
0*
09
0>
0C
#810210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#810220000000
0!
0*
09
0>
0C
#810230000000
1!
1*
b101 6
19
1>
1C
b101 G
#810240000000
0!
0*
09
0>
0C
#810250000000
1!
1*
b110 6
19
1>
1C
b110 G
#810260000000
0!
0*
09
0>
0C
#810270000000
1!
1*
b111 6
19
1>
1C
b111 G
#810280000000
0!
0*
09
0>
0C
#810290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#810300000000
0!
0*
09
0>
0C
#810310000000
1!
1*
b1 6
19
1>
1C
b1 G
#810320000000
0!
0*
09
0>
0C
#810330000000
1!
1*
b10 6
19
1>
1C
b10 G
#810340000000
0!
0*
09
0>
0C
#810350000000
1!
1*
b11 6
19
1>
1C
b11 G
#810360000000
0!
0*
09
0>
0C
#810370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#810380000000
0!
0*
09
0>
0C
#810390000000
1!
1*
b101 6
19
1>
1C
b101 G
#810400000000
0!
0*
09
0>
0C
#810410000000
1!
1*
b110 6
19
1>
1C
b110 G
#810420000000
0!
0*
09
0>
0C
#810430000000
1!
1*
b111 6
19
1>
1C
b111 G
#810440000000
0!
0*
09
0>
0C
#810450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#810460000000
0!
0*
09
0>
0C
#810470000000
1!
1*
b1 6
19
1>
1C
b1 G
#810480000000
0!
0*
09
0>
0C
#810490000000
1!
1*
b10 6
19
1>
1C
b10 G
#810500000000
0!
0*
09
0>
0C
#810510000000
1!
1*
b11 6
19
1>
1C
b11 G
#810520000000
0!
0*
09
0>
0C
#810530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#810540000000
0!
0*
09
0>
0C
#810550000000
1!
1*
b101 6
19
1>
1C
b101 G
#810560000000
0!
0*
09
0>
0C
#810570000000
1!
1*
b110 6
19
1>
1C
b110 G
#810580000000
0!
0*
09
0>
0C
#810590000000
1!
1*
b111 6
19
1>
1C
b111 G
#810600000000
0!
1"
0*
1+
09
1:
0>
0C
#810610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#810620000000
0!
0*
09
0>
0C
#810630000000
1!
1*
b1 6
19
1>
1C
b1 G
#810640000000
0!
0*
09
0>
0C
#810650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#810660000000
0!
0*
09
0>
0C
#810670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#810680000000
0!
0*
09
0>
0C
#810690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#810700000000
0!
0*
09
0>
0C
#810710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#810720000000
0!
0#
0*
0,
09
0>
0?
0C
#810730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#810740000000
0!
0*
09
0>
0C
#810750000000
1!
1*
19
1>
1C
#810760000000
0!
0*
09
0>
0C
#810770000000
1!
1*
19
1>
1C
#810780000000
0!
0*
09
0>
0C
#810790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#810800000000
0!
0*
09
0>
0C
#810810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#810820000000
0!
0*
09
0>
0C
#810830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#810840000000
0!
0*
09
0>
0C
#810850000000
1!
1*
b10 6
19
1>
1C
b10 G
#810860000000
0!
0*
09
0>
0C
#810870000000
1!
1*
b11 6
19
1>
1C
b11 G
#810880000000
0!
0*
09
0>
0C
#810890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#810900000000
0!
0*
09
0>
0C
#810910000000
1!
1*
b101 6
19
1>
1C
b101 G
#810920000000
0!
0*
09
0>
0C
#810930000000
1!
1*
b110 6
19
1>
1C
b110 G
#810940000000
0!
0*
09
0>
0C
#810950000000
1!
1*
b111 6
19
1>
1C
b111 G
#810960000000
0!
0*
09
0>
0C
#810970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#810980000000
0!
0*
09
0>
0C
#810990000000
1!
1*
b1 6
19
1>
1C
b1 G
#811000000000
0!
0*
09
0>
0C
#811010000000
1!
1*
b10 6
19
1>
1C
b10 G
#811020000000
0!
0*
09
0>
0C
#811030000000
1!
1*
b11 6
19
1>
1C
b11 G
#811040000000
0!
0*
09
0>
0C
#811050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#811060000000
0!
0*
09
0>
0C
#811070000000
1!
1*
b101 6
19
1>
1C
b101 G
#811080000000
0!
0*
09
0>
0C
#811090000000
1!
1*
b110 6
19
1>
1C
b110 G
#811100000000
0!
0*
09
0>
0C
#811110000000
1!
1*
b111 6
19
1>
1C
b111 G
#811120000000
0!
0*
09
0>
0C
#811130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#811140000000
0!
0*
09
0>
0C
#811150000000
1!
1*
b1 6
19
1>
1C
b1 G
#811160000000
0!
0*
09
0>
0C
#811170000000
1!
1*
b10 6
19
1>
1C
b10 G
#811180000000
0!
0*
09
0>
0C
#811190000000
1!
1*
b11 6
19
1>
1C
b11 G
#811200000000
0!
0*
09
0>
0C
#811210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#811220000000
0!
0*
09
0>
0C
#811230000000
1!
1*
b101 6
19
1>
1C
b101 G
#811240000000
0!
0*
09
0>
0C
#811250000000
1!
1*
b110 6
19
1>
1C
b110 G
#811260000000
0!
0*
09
0>
0C
#811270000000
1!
1*
b111 6
19
1>
1C
b111 G
#811280000000
0!
1"
0*
1+
09
1:
0>
0C
#811290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#811300000000
0!
0*
09
0>
0C
#811310000000
1!
1*
b1 6
19
1>
1C
b1 G
#811320000000
0!
0*
09
0>
0C
#811330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#811340000000
0!
0*
09
0>
0C
#811350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#811360000000
0!
0*
09
0>
0C
#811370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#811380000000
0!
0*
09
0>
0C
#811390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#811400000000
0!
0#
0*
0,
09
0>
0?
0C
#811410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#811420000000
0!
0*
09
0>
0C
#811430000000
1!
1*
19
1>
1C
#811440000000
0!
0*
09
0>
0C
#811450000000
1!
1*
19
1>
1C
#811460000000
0!
0*
09
0>
0C
#811470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#811480000000
0!
0*
09
0>
0C
#811490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#811500000000
0!
0*
09
0>
0C
#811510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#811520000000
0!
0*
09
0>
0C
#811530000000
1!
1*
b10 6
19
1>
1C
b10 G
#811540000000
0!
0*
09
0>
0C
#811550000000
1!
1*
b11 6
19
1>
1C
b11 G
#811560000000
0!
0*
09
0>
0C
#811570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#811580000000
0!
0*
09
0>
0C
#811590000000
1!
1*
b101 6
19
1>
1C
b101 G
#811600000000
0!
0*
09
0>
0C
#811610000000
1!
1*
b110 6
19
1>
1C
b110 G
#811620000000
0!
0*
09
0>
0C
#811630000000
1!
1*
b111 6
19
1>
1C
b111 G
#811640000000
0!
0*
09
0>
0C
#811650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#811660000000
0!
0*
09
0>
0C
#811670000000
1!
1*
b1 6
19
1>
1C
b1 G
#811680000000
0!
0*
09
0>
0C
#811690000000
1!
1*
b10 6
19
1>
1C
b10 G
#811700000000
0!
0*
09
0>
0C
#811710000000
1!
1*
b11 6
19
1>
1C
b11 G
#811720000000
0!
0*
09
0>
0C
#811730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#811740000000
0!
0*
09
0>
0C
#811750000000
1!
1*
b101 6
19
1>
1C
b101 G
#811760000000
0!
0*
09
0>
0C
#811770000000
1!
1*
b110 6
19
1>
1C
b110 G
#811780000000
0!
0*
09
0>
0C
#811790000000
1!
1*
b111 6
19
1>
1C
b111 G
#811800000000
0!
0*
09
0>
0C
#811810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#811820000000
0!
0*
09
0>
0C
#811830000000
1!
1*
b1 6
19
1>
1C
b1 G
#811840000000
0!
0*
09
0>
0C
#811850000000
1!
1*
b10 6
19
1>
1C
b10 G
#811860000000
0!
0*
09
0>
0C
#811870000000
1!
1*
b11 6
19
1>
1C
b11 G
#811880000000
0!
0*
09
0>
0C
#811890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#811900000000
0!
0*
09
0>
0C
#811910000000
1!
1*
b101 6
19
1>
1C
b101 G
#811920000000
0!
0*
09
0>
0C
#811930000000
1!
1*
b110 6
19
1>
1C
b110 G
#811940000000
0!
0*
09
0>
0C
#811950000000
1!
1*
b111 6
19
1>
1C
b111 G
#811960000000
0!
1"
0*
1+
09
1:
0>
0C
#811970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#811980000000
0!
0*
09
0>
0C
#811990000000
1!
1*
b1 6
19
1>
1C
b1 G
#812000000000
0!
0*
09
0>
0C
#812010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#812020000000
0!
0*
09
0>
0C
#812030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#812040000000
0!
0*
09
0>
0C
#812050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#812060000000
0!
0*
09
0>
0C
#812070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#812080000000
0!
0#
0*
0,
09
0>
0?
0C
#812090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#812100000000
0!
0*
09
0>
0C
#812110000000
1!
1*
19
1>
1C
#812120000000
0!
0*
09
0>
0C
#812130000000
1!
1*
19
1>
1C
#812140000000
0!
0*
09
0>
0C
#812150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#812160000000
0!
0*
09
0>
0C
#812170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#812180000000
0!
0*
09
0>
0C
#812190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#812200000000
0!
0*
09
0>
0C
#812210000000
1!
1*
b10 6
19
1>
1C
b10 G
#812220000000
0!
0*
09
0>
0C
#812230000000
1!
1*
b11 6
19
1>
1C
b11 G
#812240000000
0!
0*
09
0>
0C
#812250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#812260000000
0!
0*
09
0>
0C
#812270000000
1!
1*
b101 6
19
1>
1C
b101 G
#812280000000
0!
0*
09
0>
0C
#812290000000
1!
1*
b110 6
19
1>
1C
b110 G
#812300000000
0!
0*
09
0>
0C
#812310000000
1!
1*
b111 6
19
1>
1C
b111 G
#812320000000
0!
0*
09
0>
0C
#812330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#812340000000
0!
0*
09
0>
0C
#812350000000
1!
1*
b1 6
19
1>
1C
b1 G
#812360000000
0!
0*
09
0>
0C
#812370000000
1!
1*
b10 6
19
1>
1C
b10 G
#812380000000
0!
0*
09
0>
0C
#812390000000
1!
1*
b11 6
19
1>
1C
b11 G
#812400000000
0!
0*
09
0>
0C
#812410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#812420000000
0!
0*
09
0>
0C
#812430000000
1!
1*
b101 6
19
1>
1C
b101 G
#812440000000
0!
0*
09
0>
0C
#812450000000
1!
1*
b110 6
19
1>
1C
b110 G
#812460000000
0!
0*
09
0>
0C
#812470000000
1!
1*
b111 6
19
1>
1C
b111 G
#812480000000
0!
0*
09
0>
0C
#812490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#812500000000
0!
0*
09
0>
0C
#812510000000
1!
1*
b1 6
19
1>
1C
b1 G
#812520000000
0!
0*
09
0>
0C
#812530000000
1!
1*
b10 6
19
1>
1C
b10 G
#812540000000
0!
0*
09
0>
0C
#812550000000
1!
1*
b11 6
19
1>
1C
b11 G
#812560000000
0!
0*
09
0>
0C
#812570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#812580000000
0!
0*
09
0>
0C
#812590000000
1!
1*
b101 6
19
1>
1C
b101 G
#812600000000
0!
0*
09
0>
0C
#812610000000
1!
1*
b110 6
19
1>
1C
b110 G
#812620000000
0!
0*
09
0>
0C
#812630000000
1!
1*
b111 6
19
1>
1C
b111 G
#812640000000
0!
1"
0*
1+
09
1:
0>
0C
#812650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#812660000000
0!
0*
09
0>
0C
#812670000000
1!
1*
b1 6
19
1>
1C
b1 G
#812680000000
0!
0*
09
0>
0C
#812690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#812700000000
0!
0*
09
0>
0C
#812710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#812720000000
0!
0*
09
0>
0C
#812730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#812740000000
0!
0*
09
0>
0C
#812750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#812760000000
0!
0#
0*
0,
09
0>
0?
0C
#812770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#812780000000
0!
0*
09
0>
0C
#812790000000
1!
1*
19
1>
1C
#812800000000
0!
0*
09
0>
0C
#812810000000
1!
1*
19
1>
1C
#812820000000
0!
0*
09
0>
0C
#812830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#812840000000
0!
0*
09
0>
0C
#812850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#812860000000
0!
0*
09
0>
0C
#812870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#812880000000
0!
0*
09
0>
0C
#812890000000
1!
1*
b10 6
19
1>
1C
b10 G
#812900000000
0!
0*
09
0>
0C
#812910000000
1!
1*
b11 6
19
1>
1C
b11 G
#812920000000
0!
0*
09
0>
0C
#812930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#812940000000
0!
0*
09
0>
0C
#812950000000
1!
1*
b101 6
19
1>
1C
b101 G
#812960000000
0!
0*
09
0>
0C
#812970000000
1!
1*
b110 6
19
1>
1C
b110 G
#812980000000
0!
0*
09
0>
0C
#812990000000
1!
1*
b111 6
19
1>
1C
b111 G
#813000000000
0!
0*
09
0>
0C
#813010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#813020000000
0!
0*
09
0>
0C
#813030000000
1!
1*
b1 6
19
1>
1C
b1 G
#813040000000
0!
0*
09
0>
0C
#813050000000
1!
1*
b10 6
19
1>
1C
b10 G
#813060000000
0!
0*
09
0>
0C
#813070000000
1!
1*
b11 6
19
1>
1C
b11 G
#813080000000
0!
0*
09
0>
0C
#813090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#813100000000
0!
0*
09
0>
0C
#813110000000
1!
1*
b101 6
19
1>
1C
b101 G
#813120000000
0!
0*
09
0>
0C
#813130000000
1!
1*
b110 6
19
1>
1C
b110 G
#813140000000
0!
0*
09
0>
0C
#813150000000
1!
1*
b111 6
19
1>
1C
b111 G
#813160000000
0!
0*
09
0>
0C
#813170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#813180000000
0!
0*
09
0>
0C
#813190000000
1!
1*
b1 6
19
1>
1C
b1 G
#813200000000
0!
0*
09
0>
0C
#813210000000
1!
1*
b10 6
19
1>
1C
b10 G
#813220000000
0!
0*
09
0>
0C
#813230000000
1!
1*
b11 6
19
1>
1C
b11 G
#813240000000
0!
0*
09
0>
0C
#813250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#813260000000
0!
0*
09
0>
0C
#813270000000
1!
1*
b101 6
19
1>
1C
b101 G
#813280000000
0!
0*
09
0>
0C
#813290000000
1!
1*
b110 6
19
1>
1C
b110 G
#813300000000
0!
0*
09
0>
0C
#813310000000
1!
1*
b111 6
19
1>
1C
b111 G
#813320000000
0!
1"
0*
1+
09
1:
0>
0C
#813330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#813340000000
0!
0*
09
0>
0C
#813350000000
1!
1*
b1 6
19
1>
1C
b1 G
#813360000000
0!
0*
09
0>
0C
#813370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#813380000000
0!
0*
09
0>
0C
#813390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#813400000000
0!
0*
09
0>
0C
#813410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#813420000000
0!
0*
09
0>
0C
#813430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#813440000000
0!
0#
0*
0,
09
0>
0?
0C
#813450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#813460000000
0!
0*
09
0>
0C
#813470000000
1!
1*
19
1>
1C
#813480000000
0!
0*
09
0>
0C
#813490000000
1!
1*
19
1>
1C
#813500000000
0!
0*
09
0>
0C
#813510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#813520000000
0!
0*
09
0>
0C
#813530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#813540000000
0!
0*
09
0>
0C
#813550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#813560000000
0!
0*
09
0>
0C
#813570000000
1!
1*
b10 6
19
1>
1C
b10 G
#813580000000
0!
0*
09
0>
0C
#813590000000
1!
1*
b11 6
19
1>
1C
b11 G
#813600000000
0!
0*
09
0>
0C
#813610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#813620000000
0!
0*
09
0>
0C
#813630000000
1!
1*
b101 6
19
1>
1C
b101 G
#813640000000
0!
0*
09
0>
0C
#813650000000
1!
1*
b110 6
19
1>
1C
b110 G
#813660000000
0!
0*
09
0>
0C
#813670000000
1!
1*
b111 6
19
1>
1C
b111 G
#813680000000
0!
0*
09
0>
0C
#813690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#813700000000
0!
0*
09
0>
0C
#813710000000
1!
1*
b1 6
19
1>
1C
b1 G
#813720000000
0!
0*
09
0>
0C
#813730000000
1!
1*
b10 6
19
1>
1C
b10 G
#813740000000
0!
0*
09
0>
0C
#813750000000
1!
1*
b11 6
19
1>
1C
b11 G
#813760000000
0!
0*
09
0>
0C
#813770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#813780000000
0!
0*
09
0>
0C
#813790000000
1!
1*
b101 6
19
1>
1C
b101 G
#813800000000
0!
0*
09
0>
0C
#813810000000
1!
1*
b110 6
19
1>
1C
b110 G
#813820000000
0!
0*
09
0>
0C
#813830000000
1!
1*
b111 6
19
1>
1C
b111 G
#813840000000
0!
0*
09
0>
0C
#813850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#813860000000
0!
0*
09
0>
0C
#813870000000
1!
1*
b1 6
19
1>
1C
b1 G
#813880000000
0!
0*
09
0>
0C
#813890000000
1!
1*
b10 6
19
1>
1C
b10 G
#813900000000
0!
0*
09
0>
0C
#813910000000
1!
1*
b11 6
19
1>
1C
b11 G
#813920000000
0!
0*
09
0>
0C
#813930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#813940000000
0!
0*
09
0>
0C
#813950000000
1!
1*
b101 6
19
1>
1C
b101 G
#813960000000
0!
0*
09
0>
0C
#813970000000
1!
1*
b110 6
19
1>
1C
b110 G
#813980000000
0!
0*
09
0>
0C
#813990000000
1!
1*
b111 6
19
1>
1C
b111 G
#814000000000
0!
1"
0*
1+
09
1:
0>
0C
#814010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#814020000000
0!
0*
09
0>
0C
#814030000000
1!
1*
b1 6
19
1>
1C
b1 G
#814040000000
0!
0*
09
0>
0C
#814050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#814060000000
0!
0*
09
0>
0C
#814070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#814080000000
0!
0*
09
0>
0C
#814090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#814100000000
0!
0*
09
0>
0C
#814110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#814120000000
0!
0#
0*
0,
09
0>
0?
0C
#814130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#814140000000
0!
0*
09
0>
0C
#814150000000
1!
1*
19
1>
1C
#814160000000
0!
0*
09
0>
0C
#814170000000
1!
1*
19
1>
1C
#814180000000
0!
0*
09
0>
0C
#814190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#814200000000
0!
0*
09
0>
0C
#814210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#814220000000
0!
0*
09
0>
0C
#814230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#814240000000
0!
0*
09
0>
0C
#814250000000
1!
1*
b10 6
19
1>
1C
b10 G
#814260000000
0!
0*
09
0>
0C
#814270000000
1!
1*
b11 6
19
1>
1C
b11 G
#814280000000
0!
0*
09
0>
0C
#814290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#814300000000
0!
0*
09
0>
0C
#814310000000
1!
1*
b101 6
19
1>
1C
b101 G
#814320000000
0!
0*
09
0>
0C
#814330000000
1!
1*
b110 6
19
1>
1C
b110 G
#814340000000
0!
0*
09
0>
0C
#814350000000
1!
1*
b111 6
19
1>
1C
b111 G
#814360000000
0!
0*
09
0>
0C
#814370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#814380000000
0!
0*
09
0>
0C
#814390000000
1!
1*
b1 6
19
1>
1C
b1 G
#814400000000
0!
0*
09
0>
0C
#814410000000
1!
1*
b10 6
19
1>
1C
b10 G
#814420000000
0!
0*
09
0>
0C
#814430000000
1!
1*
b11 6
19
1>
1C
b11 G
#814440000000
0!
0*
09
0>
0C
#814450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#814460000000
0!
0*
09
0>
0C
#814470000000
1!
1*
b101 6
19
1>
1C
b101 G
#814480000000
0!
0*
09
0>
0C
#814490000000
1!
1*
b110 6
19
1>
1C
b110 G
#814500000000
0!
0*
09
0>
0C
#814510000000
1!
1*
b111 6
19
1>
1C
b111 G
#814520000000
0!
0*
09
0>
0C
#814530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#814540000000
0!
0*
09
0>
0C
#814550000000
1!
1*
b1 6
19
1>
1C
b1 G
#814560000000
0!
0*
09
0>
0C
#814570000000
1!
1*
b10 6
19
1>
1C
b10 G
#814580000000
0!
0*
09
0>
0C
#814590000000
1!
1*
b11 6
19
1>
1C
b11 G
#814600000000
0!
0*
09
0>
0C
#814610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#814620000000
0!
0*
09
0>
0C
#814630000000
1!
1*
b101 6
19
1>
1C
b101 G
#814640000000
0!
0*
09
0>
0C
#814650000000
1!
1*
b110 6
19
1>
1C
b110 G
#814660000000
0!
0*
09
0>
0C
#814670000000
1!
1*
b111 6
19
1>
1C
b111 G
#814680000000
0!
1"
0*
1+
09
1:
0>
0C
#814690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#814700000000
0!
0*
09
0>
0C
#814710000000
1!
1*
b1 6
19
1>
1C
b1 G
#814720000000
0!
0*
09
0>
0C
#814730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#814740000000
0!
0*
09
0>
0C
#814750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#814760000000
0!
0*
09
0>
0C
#814770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#814780000000
0!
0*
09
0>
0C
#814790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#814800000000
0!
0#
0*
0,
09
0>
0?
0C
#814810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#814820000000
0!
0*
09
0>
0C
#814830000000
1!
1*
19
1>
1C
#814840000000
0!
0*
09
0>
0C
#814850000000
1!
1*
19
1>
1C
#814860000000
0!
0*
09
0>
0C
#814870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#814880000000
0!
0*
09
0>
0C
#814890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#814900000000
0!
0*
09
0>
0C
#814910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#814920000000
0!
0*
09
0>
0C
#814930000000
1!
1*
b10 6
19
1>
1C
b10 G
#814940000000
0!
0*
09
0>
0C
#814950000000
1!
1*
b11 6
19
1>
1C
b11 G
#814960000000
0!
0*
09
0>
0C
#814970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#814980000000
0!
0*
09
0>
0C
#814990000000
1!
1*
b101 6
19
1>
1C
b101 G
#815000000000
0!
0*
09
0>
0C
#815010000000
1!
1*
b110 6
19
1>
1C
b110 G
#815020000000
0!
0*
09
0>
0C
#815030000000
1!
1*
b111 6
19
1>
1C
b111 G
#815040000000
0!
0*
09
0>
0C
#815050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#815060000000
0!
0*
09
0>
0C
#815070000000
1!
1*
b1 6
19
1>
1C
b1 G
#815080000000
0!
0*
09
0>
0C
#815090000000
1!
1*
b10 6
19
1>
1C
b10 G
#815100000000
0!
0*
09
0>
0C
#815110000000
1!
1*
b11 6
19
1>
1C
b11 G
#815120000000
0!
0*
09
0>
0C
#815130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#815140000000
0!
0*
09
0>
0C
#815150000000
1!
1*
b101 6
19
1>
1C
b101 G
#815160000000
0!
0*
09
0>
0C
#815170000000
1!
1*
b110 6
19
1>
1C
b110 G
#815180000000
0!
0*
09
0>
0C
#815190000000
1!
1*
b111 6
19
1>
1C
b111 G
#815200000000
0!
0*
09
0>
0C
#815210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#815220000000
0!
0*
09
0>
0C
#815230000000
1!
1*
b1 6
19
1>
1C
b1 G
#815240000000
0!
0*
09
0>
0C
#815250000000
1!
1*
b10 6
19
1>
1C
b10 G
#815260000000
0!
0*
09
0>
0C
#815270000000
1!
1*
b11 6
19
1>
1C
b11 G
#815280000000
0!
0*
09
0>
0C
#815290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#815300000000
0!
0*
09
0>
0C
#815310000000
1!
1*
b101 6
19
1>
1C
b101 G
#815320000000
0!
0*
09
0>
0C
#815330000000
1!
1*
b110 6
19
1>
1C
b110 G
#815340000000
0!
0*
09
0>
0C
#815350000000
1!
1*
b111 6
19
1>
1C
b111 G
#815360000000
0!
1"
0*
1+
09
1:
0>
0C
#815370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#815380000000
0!
0*
09
0>
0C
#815390000000
1!
1*
b1 6
19
1>
1C
b1 G
#815400000000
0!
0*
09
0>
0C
#815410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#815420000000
0!
0*
09
0>
0C
#815430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#815440000000
0!
0*
09
0>
0C
#815450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#815460000000
0!
0*
09
0>
0C
#815470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#815480000000
0!
0#
0*
0,
09
0>
0?
0C
#815490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#815500000000
0!
0*
09
0>
0C
#815510000000
1!
1*
19
1>
1C
#815520000000
0!
0*
09
0>
0C
#815530000000
1!
1*
19
1>
1C
#815540000000
0!
0*
09
0>
0C
#815550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#815560000000
0!
0*
09
0>
0C
#815570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#815580000000
0!
0*
09
0>
0C
#815590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#815600000000
0!
0*
09
0>
0C
#815610000000
1!
1*
b10 6
19
1>
1C
b10 G
#815620000000
0!
0*
09
0>
0C
#815630000000
1!
1*
b11 6
19
1>
1C
b11 G
#815640000000
0!
0*
09
0>
0C
#815650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#815660000000
0!
0*
09
0>
0C
#815670000000
1!
1*
b101 6
19
1>
1C
b101 G
#815680000000
0!
0*
09
0>
0C
#815690000000
1!
1*
b110 6
19
1>
1C
b110 G
#815700000000
0!
0*
09
0>
0C
#815710000000
1!
1*
b111 6
19
1>
1C
b111 G
#815720000000
0!
0*
09
0>
0C
#815730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#815740000000
0!
0*
09
0>
0C
#815750000000
1!
1*
b1 6
19
1>
1C
b1 G
#815760000000
0!
0*
09
0>
0C
#815770000000
1!
1*
b10 6
19
1>
1C
b10 G
#815780000000
0!
0*
09
0>
0C
#815790000000
1!
1*
b11 6
19
1>
1C
b11 G
#815800000000
0!
0*
09
0>
0C
#815810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#815820000000
0!
0*
09
0>
0C
#815830000000
1!
1*
b101 6
19
1>
1C
b101 G
#815840000000
0!
0*
09
0>
0C
#815850000000
1!
1*
b110 6
19
1>
1C
b110 G
#815860000000
0!
0*
09
0>
0C
#815870000000
1!
1*
b111 6
19
1>
1C
b111 G
#815880000000
0!
0*
09
0>
0C
#815890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#815900000000
0!
0*
09
0>
0C
#815910000000
1!
1*
b1 6
19
1>
1C
b1 G
#815920000000
0!
0*
09
0>
0C
#815930000000
1!
1*
b10 6
19
1>
1C
b10 G
#815940000000
0!
0*
09
0>
0C
#815950000000
1!
1*
b11 6
19
1>
1C
b11 G
#815960000000
0!
0*
09
0>
0C
#815970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#815980000000
0!
0*
09
0>
0C
#815990000000
1!
1*
b101 6
19
1>
1C
b101 G
#816000000000
0!
0*
09
0>
0C
#816010000000
1!
1*
b110 6
19
1>
1C
b110 G
#816020000000
0!
0*
09
0>
0C
#816030000000
1!
1*
b111 6
19
1>
1C
b111 G
#816040000000
0!
1"
0*
1+
09
1:
0>
0C
#816050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#816060000000
0!
0*
09
0>
0C
#816070000000
1!
1*
b1 6
19
1>
1C
b1 G
#816080000000
0!
0*
09
0>
0C
#816090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#816100000000
0!
0*
09
0>
0C
#816110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#816120000000
0!
0*
09
0>
0C
#816130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#816140000000
0!
0*
09
0>
0C
#816150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#816160000000
0!
0#
0*
0,
09
0>
0?
0C
#816170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#816180000000
0!
0*
09
0>
0C
#816190000000
1!
1*
19
1>
1C
#816200000000
0!
0*
09
0>
0C
#816210000000
1!
1*
19
1>
1C
#816220000000
0!
0*
09
0>
0C
#816230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#816240000000
0!
0*
09
0>
0C
#816250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#816260000000
0!
0*
09
0>
0C
#816270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#816280000000
0!
0*
09
0>
0C
#816290000000
1!
1*
b10 6
19
1>
1C
b10 G
#816300000000
0!
0*
09
0>
0C
#816310000000
1!
1*
b11 6
19
1>
1C
b11 G
#816320000000
0!
0*
09
0>
0C
#816330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#816340000000
0!
0*
09
0>
0C
#816350000000
1!
1*
b101 6
19
1>
1C
b101 G
#816360000000
0!
0*
09
0>
0C
#816370000000
1!
1*
b110 6
19
1>
1C
b110 G
#816380000000
0!
0*
09
0>
0C
#816390000000
1!
1*
b111 6
19
1>
1C
b111 G
#816400000000
0!
0*
09
0>
0C
#816410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#816420000000
0!
0*
09
0>
0C
#816430000000
1!
1*
b1 6
19
1>
1C
b1 G
#816440000000
0!
0*
09
0>
0C
#816450000000
1!
1*
b10 6
19
1>
1C
b10 G
#816460000000
0!
0*
09
0>
0C
#816470000000
1!
1*
b11 6
19
1>
1C
b11 G
#816480000000
0!
0*
09
0>
0C
#816490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#816500000000
0!
0*
09
0>
0C
#816510000000
1!
1*
b101 6
19
1>
1C
b101 G
#816520000000
0!
0*
09
0>
0C
#816530000000
1!
1*
b110 6
19
1>
1C
b110 G
#816540000000
0!
0*
09
0>
0C
#816550000000
1!
1*
b111 6
19
1>
1C
b111 G
#816560000000
0!
0*
09
0>
0C
#816570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#816580000000
0!
0*
09
0>
0C
#816590000000
1!
1*
b1 6
19
1>
1C
b1 G
#816600000000
0!
0*
09
0>
0C
#816610000000
1!
1*
b10 6
19
1>
1C
b10 G
#816620000000
0!
0*
09
0>
0C
#816630000000
1!
1*
b11 6
19
1>
1C
b11 G
#816640000000
0!
0*
09
0>
0C
#816650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#816660000000
0!
0*
09
0>
0C
#816670000000
1!
1*
b101 6
19
1>
1C
b101 G
#816680000000
0!
0*
09
0>
0C
#816690000000
1!
1*
b110 6
19
1>
1C
b110 G
#816700000000
0!
0*
09
0>
0C
#816710000000
1!
1*
b111 6
19
1>
1C
b111 G
#816720000000
0!
1"
0*
1+
09
1:
0>
0C
#816730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#816740000000
0!
0*
09
0>
0C
#816750000000
1!
1*
b1 6
19
1>
1C
b1 G
#816760000000
0!
0*
09
0>
0C
#816770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#816780000000
0!
0*
09
0>
0C
#816790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#816800000000
0!
0*
09
0>
0C
#816810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#816820000000
0!
0*
09
0>
0C
#816830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#816840000000
0!
0#
0*
0,
09
0>
0?
0C
#816850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#816860000000
0!
0*
09
0>
0C
#816870000000
1!
1*
19
1>
1C
#816880000000
0!
0*
09
0>
0C
#816890000000
1!
1*
19
1>
1C
#816900000000
0!
0*
09
0>
0C
#816910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#816920000000
0!
0*
09
0>
0C
#816930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#816940000000
0!
0*
09
0>
0C
#816950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#816960000000
0!
0*
09
0>
0C
#816970000000
1!
1*
b10 6
19
1>
1C
b10 G
#816980000000
0!
0*
09
0>
0C
#816990000000
1!
1*
b11 6
19
1>
1C
b11 G
#817000000000
0!
0*
09
0>
0C
#817010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#817020000000
0!
0*
09
0>
0C
#817030000000
1!
1*
b101 6
19
1>
1C
b101 G
#817040000000
0!
0*
09
0>
0C
#817050000000
1!
1*
b110 6
19
1>
1C
b110 G
#817060000000
0!
0*
09
0>
0C
#817070000000
1!
1*
b111 6
19
1>
1C
b111 G
#817080000000
0!
0*
09
0>
0C
#817090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#817100000000
0!
0*
09
0>
0C
#817110000000
1!
1*
b1 6
19
1>
1C
b1 G
#817120000000
0!
0*
09
0>
0C
#817130000000
1!
1*
b10 6
19
1>
1C
b10 G
#817140000000
0!
0*
09
0>
0C
#817150000000
1!
1*
b11 6
19
1>
1C
b11 G
#817160000000
0!
0*
09
0>
0C
#817170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#817180000000
0!
0*
09
0>
0C
#817190000000
1!
1*
b101 6
19
1>
1C
b101 G
#817200000000
0!
0*
09
0>
0C
#817210000000
1!
1*
b110 6
19
1>
1C
b110 G
#817220000000
0!
0*
09
0>
0C
#817230000000
1!
1*
b111 6
19
1>
1C
b111 G
#817240000000
0!
0*
09
0>
0C
#817250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#817260000000
0!
0*
09
0>
0C
#817270000000
1!
1*
b1 6
19
1>
1C
b1 G
#817280000000
0!
0*
09
0>
0C
#817290000000
1!
1*
b10 6
19
1>
1C
b10 G
#817300000000
0!
0*
09
0>
0C
#817310000000
1!
1*
b11 6
19
1>
1C
b11 G
#817320000000
0!
0*
09
0>
0C
#817330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#817340000000
0!
0*
09
0>
0C
#817350000000
1!
1*
b101 6
19
1>
1C
b101 G
#817360000000
0!
0*
09
0>
0C
#817370000000
1!
1*
b110 6
19
1>
1C
b110 G
#817380000000
0!
0*
09
0>
0C
#817390000000
1!
1*
b111 6
19
1>
1C
b111 G
#817400000000
0!
1"
0*
1+
09
1:
0>
0C
#817410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#817420000000
0!
0*
09
0>
0C
#817430000000
1!
1*
b1 6
19
1>
1C
b1 G
#817440000000
0!
0*
09
0>
0C
#817450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#817460000000
0!
0*
09
0>
0C
#817470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#817480000000
0!
0*
09
0>
0C
#817490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#817500000000
0!
0*
09
0>
0C
#817510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#817520000000
0!
0#
0*
0,
09
0>
0?
0C
#817530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#817540000000
0!
0*
09
0>
0C
#817550000000
1!
1*
19
1>
1C
#817560000000
0!
0*
09
0>
0C
#817570000000
1!
1*
19
1>
1C
#817580000000
0!
0*
09
0>
0C
#817590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#817600000000
0!
0*
09
0>
0C
#817610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#817620000000
0!
0*
09
0>
0C
#817630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#817640000000
0!
0*
09
0>
0C
#817650000000
1!
1*
b10 6
19
1>
1C
b10 G
#817660000000
0!
0*
09
0>
0C
#817670000000
1!
1*
b11 6
19
1>
1C
b11 G
#817680000000
0!
0*
09
0>
0C
#817690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#817700000000
0!
0*
09
0>
0C
#817710000000
1!
1*
b101 6
19
1>
1C
b101 G
#817720000000
0!
0*
09
0>
0C
#817730000000
1!
1*
b110 6
19
1>
1C
b110 G
#817740000000
0!
0*
09
0>
0C
#817750000000
1!
1*
b111 6
19
1>
1C
b111 G
#817760000000
0!
0*
09
0>
0C
#817770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#817780000000
0!
0*
09
0>
0C
#817790000000
1!
1*
b1 6
19
1>
1C
b1 G
#817800000000
0!
0*
09
0>
0C
#817810000000
1!
1*
b10 6
19
1>
1C
b10 G
#817820000000
0!
0*
09
0>
0C
#817830000000
1!
1*
b11 6
19
1>
1C
b11 G
#817840000000
0!
0*
09
0>
0C
#817850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#817860000000
0!
0*
09
0>
0C
#817870000000
1!
1*
b101 6
19
1>
1C
b101 G
#817880000000
0!
0*
09
0>
0C
#817890000000
1!
1*
b110 6
19
1>
1C
b110 G
#817900000000
0!
0*
09
0>
0C
#817910000000
1!
1*
b111 6
19
1>
1C
b111 G
#817920000000
0!
0*
09
0>
0C
#817930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#817940000000
0!
0*
09
0>
0C
#817950000000
1!
1*
b1 6
19
1>
1C
b1 G
#817960000000
0!
0*
09
0>
0C
#817970000000
1!
1*
b10 6
19
1>
1C
b10 G
#817980000000
0!
0*
09
0>
0C
#817990000000
1!
1*
b11 6
19
1>
1C
b11 G
#818000000000
0!
0*
09
0>
0C
#818010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#818020000000
0!
0*
09
0>
0C
#818030000000
1!
1*
b101 6
19
1>
1C
b101 G
#818040000000
0!
0*
09
0>
0C
#818050000000
1!
1*
b110 6
19
1>
1C
b110 G
#818060000000
0!
0*
09
0>
0C
#818070000000
1!
1*
b111 6
19
1>
1C
b111 G
#818080000000
0!
1"
0*
1+
09
1:
0>
0C
#818090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#818100000000
0!
0*
09
0>
0C
#818110000000
1!
1*
b1 6
19
1>
1C
b1 G
#818120000000
0!
0*
09
0>
0C
#818130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#818140000000
0!
0*
09
0>
0C
#818150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#818160000000
0!
0*
09
0>
0C
#818170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#818180000000
0!
0*
09
0>
0C
#818190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#818200000000
0!
0#
0*
0,
09
0>
0?
0C
#818210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#818220000000
0!
0*
09
0>
0C
#818230000000
1!
1*
19
1>
1C
#818240000000
0!
0*
09
0>
0C
#818250000000
1!
1*
19
1>
1C
#818260000000
0!
0*
09
0>
0C
#818270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#818280000000
0!
0*
09
0>
0C
#818290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#818300000000
0!
0*
09
0>
0C
#818310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#818320000000
0!
0*
09
0>
0C
#818330000000
1!
1*
b10 6
19
1>
1C
b10 G
#818340000000
0!
0*
09
0>
0C
#818350000000
1!
1*
b11 6
19
1>
1C
b11 G
#818360000000
0!
0*
09
0>
0C
#818370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#818380000000
0!
0*
09
0>
0C
#818390000000
1!
1*
b101 6
19
1>
1C
b101 G
#818400000000
0!
0*
09
0>
0C
#818410000000
1!
1*
b110 6
19
1>
1C
b110 G
#818420000000
0!
0*
09
0>
0C
#818430000000
1!
1*
b111 6
19
1>
1C
b111 G
#818440000000
0!
0*
09
0>
0C
#818450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#818460000000
0!
0*
09
0>
0C
#818470000000
1!
1*
b1 6
19
1>
1C
b1 G
#818480000000
0!
0*
09
0>
0C
#818490000000
1!
1*
b10 6
19
1>
1C
b10 G
#818500000000
0!
0*
09
0>
0C
#818510000000
1!
1*
b11 6
19
1>
1C
b11 G
#818520000000
0!
0*
09
0>
0C
#818530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#818540000000
0!
0*
09
0>
0C
#818550000000
1!
1*
b101 6
19
1>
1C
b101 G
#818560000000
0!
0*
09
0>
0C
#818570000000
1!
1*
b110 6
19
1>
1C
b110 G
#818580000000
0!
0*
09
0>
0C
#818590000000
1!
1*
b111 6
19
1>
1C
b111 G
#818600000000
0!
0*
09
0>
0C
#818610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#818620000000
0!
0*
09
0>
0C
#818630000000
1!
1*
b1 6
19
1>
1C
b1 G
#818640000000
0!
0*
09
0>
0C
#818650000000
1!
1*
b10 6
19
1>
1C
b10 G
#818660000000
0!
0*
09
0>
0C
#818670000000
1!
1*
b11 6
19
1>
1C
b11 G
#818680000000
0!
0*
09
0>
0C
#818690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#818700000000
0!
0*
09
0>
0C
#818710000000
1!
1*
b101 6
19
1>
1C
b101 G
#818720000000
0!
0*
09
0>
0C
#818730000000
1!
1*
b110 6
19
1>
1C
b110 G
#818740000000
0!
0*
09
0>
0C
#818750000000
1!
1*
b111 6
19
1>
1C
b111 G
#818760000000
0!
1"
0*
1+
09
1:
0>
0C
#818770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#818780000000
0!
0*
09
0>
0C
#818790000000
1!
1*
b1 6
19
1>
1C
b1 G
#818800000000
0!
0*
09
0>
0C
#818810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#818820000000
0!
0*
09
0>
0C
#818830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#818840000000
0!
0*
09
0>
0C
#818850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#818860000000
0!
0*
09
0>
0C
#818870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#818880000000
0!
0#
0*
0,
09
0>
0?
0C
#818890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#818900000000
0!
0*
09
0>
0C
#818910000000
1!
1*
19
1>
1C
#818920000000
0!
0*
09
0>
0C
#818930000000
1!
1*
19
1>
1C
#818940000000
0!
0*
09
0>
0C
#818950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#818960000000
0!
0*
09
0>
0C
#818970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#818980000000
0!
0*
09
0>
0C
#818990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#819000000000
0!
0*
09
0>
0C
#819010000000
1!
1*
b10 6
19
1>
1C
b10 G
#819020000000
0!
0*
09
0>
0C
#819030000000
1!
1*
b11 6
19
1>
1C
b11 G
#819040000000
0!
0*
09
0>
0C
#819050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#819060000000
0!
0*
09
0>
0C
#819070000000
1!
1*
b101 6
19
1>
1C
b101 G
#819080000000
0!
0*
09
0>
0C
#819090000000
1!
1*
b110 6
19
1>
1C
b110 G
#819100000000
0!
0*
09
0>
0C
#819110000000
1!
1*
b111 6
19
1>
1C
b111 G
#819120000000
0!
0*
09
0>
0C
#819130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#819140000000
0!
0*
09
0>
0C
#819150000000
1!
1*
b1 6
19
1>
1C
b1 G
#819160000000
0!
0*
09
0>
0C
#819170000000
1!
1*
b10 6
19
1>
1C
b10 G
#819180000000
0!
0*
09
0>
0C
#819190000000
1!
1*
b11 6
19
1>
1C
b11 G
#819200000000
0!
0*
09
0>
0C
#819210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#819220000000
0!
0*
09
0>
0C
#819230000000
1!
1*
b101 6
19
1>
1C
b101 G
#819240000000
0!
0*
09
0>
0C
#819250000000
1!
1*
b110 6
19
1>
1C
b110 G
#819260000000
0!
0*
09
0>
0C
#819270000000
1!
1*
b111 6
19
1>
1C
b111 G
#819280000000
0!
0*
09
0>
0C
#819290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#819300000000
0!
0*
09
0>
0C
#819310000000
1!
1*
b1 6
19
1>
1C
b1 G
#819320000000
0!
0*
09
0>
0C
#819330000000
1!
1*
b10 6
19
1>
1C
b10 G
#819340000000
0!
0*
09
0>
0C
#819350000000
1!
1*
b11 6
19
1>
1C
b11 G
#819360000000
0!
0*
09
0>
0C
#819370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#819380000000
0!
0*
09
0>
0C
#819390000000
1!
1*
b101 6
19
1>
1C
b101 G
#819400000000
0!
0*
09
0>
0C
#819410000000
1!
1*
b110 6
19
1>
1C
b110 G
#819420000000
0!
0*
09
0>
0C
#819430000000
1!
1*
b111 6
19
1>
1C
b111 G
#819440000000
0!
1"
0*
1+
09
1:
0>
0C
#819450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#819460000000
0!
0*
09
0>
0C
#819470000000
1!
1*
b1 6
19
1>
1C
b1 G
#819480000000
0!
0*
09
0>
0C
#819490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#819500000000
0!
0*
09
0>
0C
#819510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#819520000000
0!
0*
09
0>
0C
#819530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#819540000000
0!
0*
09
0>
0C
#819550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#819560000000
0!
0#
0*
0,
09
0>
0?
0C
#819570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#819580000000
0!
0*
09
0>
0C
#819590000000
1!
1*
19
1>
1C
#819600000000
0!
0*
09
0>
0C
#819610000000
1!
1*
19
1>
1C
#819620000000
0!
0*
09
0>
0C
#819630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#819640000000
0!
0*
09
0>
0C
#819650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#819660000000
0!
0*
09
0>
0C
#819670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#819680000000
0!
0*
09
0>
0C
#819690000000
1!
1*
b10 6
19
1>
1C
b10 G
#819700000000
0!
0*
09
0>
0C
#819710000000
1!
1*
b11 6
19
1>
1C
b11 G
#819720000000
0!
0*
09
0>
0C
#819730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#819740000000
0!
0*
09
0>
0C
#819750000000
1!
1*
b101 6
19
1>
1C
b101 G
#819760000000
0!
0*
09
0>
0C
#819770000000
1!
1*
b110 6
19
1>
1C
b110 G
#819780000000
0!
0*
09
0>
0C
#819790000000
1!
1*
b111 6
19
1>
1C
b111 G
#819800000000
0!
0*
09
0>
0C
#819810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#819820000000
0!
0*
09
0>
0C
#819830000000
1!
1*
b1 6
19
1>
1C
b1 G
#819840000000
0!
0*
09
0>
0C
#819850000000
1!
1*
b10 6
19
1>
1C
b10 G
#819860000000
0!
0*
09
0>
0C
#819870000000
1!
1*
b11 6
19
1>
1C
b11 G
#819880000000
0!
0*
09
0>
0C
#819890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#819900000000
0!
0*
09
0>
0C
#819910000000
1!
1*
b101 6
19
1>
1C
b101 G
#819920000000
0!
0*
09
0>
0C
#819930000000
1!
1*
b110 6
19
1>
1C
b110 G
#819940000000
0!
0*
09
0>
0C
#819950000000
1!
1*
b111 6
19
1>
1C
b111 G
#819960000000
0!
0*
09
0>
0C
#819970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#819980000000
0!
0*
09
0>
0C
#819990000000
1!
1*
b1 6
19
1>
1C
b1 G
#820000000000
0!
0*
09
0>
0C
#820010000000
1!
1*
b10 6
19
1>
1C
b10 G
#820020000000
0!
0*
09
0>
0C
#820030000000
1!
1*
b11 6
19
1>
1C
b11 G
#820040000000
0!
0*
09
0>
0C
#820050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#820060000000
0!
0*
09
0>
0C
#820070000000
1!
1*
b101 6
19
1>
1C
b101 G
#820080000000
0!
0*
09
0>
0C
#820090000000
1!
1*
b110 6
19
1>
1C
b110 G
#820100000000
0!
0*
09
0>
0C
#820110000000
1!
1*
b111 6
19
1>
1C
b111 G
#820120000000
0!
1"
0*
1+
09
1:
0>
0C
#820130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#820140000000
0!
0*
09
0>
0C
#820150000000
1!
1*
b1 6
19
1>
1C
b1 G
#820160000000
0!
0*
09
0>
0C
#820170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#820180000000
0!
0*
09
0>
0C
#820190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#820200000000
0!
0*
09
0>
0C
#820210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#820220000000
0!
0*
09
0>
0C
#820230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#820240000000
0!
0#
0*
0,
09
0>
0?
0C
#820250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#820260000000
0!
0*
09
0>
0C
#820270000000
1!
1*
19
1>
1C
#820280000000
0!
0*
09
0>
0C
#820290000000
1!
1*
19
1>
1C
#820300000000
0!
0*
09
0>
0C
#820310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#820320000000
0!
0*
09
0>
0C
#820330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#820340000000
0!
0*
09
0>
0C
#820350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#820360000000
0!
0*
09
0>
0C
#820370000000
1!
1*
b10 6
19
1>
1C
b10 G
#820380000000
0!
0*
09
0>
0C
#820390000000
1!
1*
b11 6
19
1>
1C
b11 G
#820400000000
0!
0*
09
0>
0C
#820410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#820420000000
0!
0*
09
0>
0C
#820430000000
1!
1*
b101 6
19
1>
1C
b101 G
#820440000000
0!
0*
09
0>
0C
#820450000000
1!
1*
b110 6
19
1>
1C
b110 G
#820460000000
0!
0*
09
0>
0C
#820470000000
1!
1*
b111 6
19
1>
1C
b111 G
#820480000000
0!
0*
09
0>
0C
#820490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#820500000000
0!
0*
09
0>
0C
#820510000000
1!
1*
b1 6
19
1>
1C
b1 G
#820520000000
0!
0*
09
0>
0C
#820530000000
1!
1*
b10 6
19
1>
1C
b10 G
#820540000000
0!
0*
09
0>
0C
#820550000000
1!
1*
b11 6
19
1>
1C
b11 G
#820560000000
0!
0*
09
0>
0C
#820570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#820580000000
0!
0*
09
0>
0C
#820590000000
1!
1*
b101 6
19
1>
1C
b101 G
#820600000000
0!
0*
09
0>
0C
#820610000000
1!
1*
b110 6
19
1>
1C
b110 G
#820620000000
0!
0*
09
0>
0C
#820630000000
1!
1*
b111 6
19
1>
1C
b111 G
#820640000000
0!
0*
09
0>
0C
#820650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#820660000000
0!
0*
09
0>
0C
#820670000000
1!
1*
b1 6
19
1>
1C
b1 G
#820680000000
0!
0*
09
0>
0C
#820690000000
1!
1*
b10 6
19
1>
1C
b10 G
#820700000000
0!
0*
09
0>
0C
#820710000000
1!
1*
b11 6
19
1>
1C
b11 G
#820720000000
0!
0*
09
0>
0C
#820730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#820740000000
0!
0*
09
0>
0C
#820750000000
1!
1*
b101 6
19
1>
1C
b101 G
#820760000000
0!
0*
09
0>
0C
#820770000000
1!
1*
b110 6
19
1>
1C
b110 G
#820780000000
0!
0*
09
0>
0C
#820790000000
1!
1*
b111 6
19
1>
1C
b111 G
#820800000000
0!
1"
0*
1+
09
1:
0>
0C
#820810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#820820000000
0!
0*
09
0>
0C
#820830000000
1!
1*
b1 6
19
1>
1C
b1 G
#820840000000
0!
0*
09
0>
0C
#820850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#820860000000
0!
0*
09
0>
0C
#820870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#820880000000
0!
0*
09
0>
0C
#820890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#820900000000
0!
0*
09
0>
0C
#820910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#820920000000
0!
0#
0*
0,
09
0>
0?
0C
#820930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#820940000000
0!
0*
09
0>
0C
#820950000000
1!
1*
19
1>
1C
#820960000000
0!
0*
09
0>
0C
#820970000000
1!
1*
19
1>
1C
#820980000000
0!
0*
09
0>
0C
#820990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#821000000000
0!
0*
09
0>
0C
#821010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#821020000000
0!
0*
09
0>
0C
#821030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#821040000000
0!
0*
09
0>
0C
#821050000000
1!
1*
b10 6
19
1>
1C
b10 G
#821060000000
0!
0*
09
0>
0C
#821070000000
1!
1*
b11 6
19
1>
1C
b11 G
#821080000000
0!
0*
09
0>
0C
#821090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#821100000000
0!
0*
09
0>
0C
#821110000000
1!
1*
b101 6
19
1>
1C
b101 G
#821120000000
0!
0*
09
0>
0C
#821130000000
1!
1*
b110 6
19
1>
1C
b110 G
#821140000000
0!
0*
09
0>
0C
#821150000000
1!
1*
b111 6
19
1>
1C
b111 G
#821160000000
0!
0*
09
0>
0C
#821170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#821180000000
0!
0*
09
0>
0C
#821190000000
1!
1*
b1 6
19
1>
1C
b1 G
#821200000000
0!
0*
09
0>
0C
#821210000000
1!
1*
b10 6
19
1>
1C
b10 G
#821220000000
0!
0*
09
0>
0C
#821230000000
1!
1*
b11 6
19
1>
1C
b11 G
#821240000000
0!
0*
09
0>
0C
#821250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#821260000000
0!
0*
09
0>
0C
#821270000000
1!
1*
b101 6
19
1>
1C
b101 G
#821280000000
0!
0*
09
0>
0C
#821290000000
1!
1*
b110 6
19
1>
1C
b110 G
#821300000000
0!
0*
09
0>
0C
#821310000000
1!
1*
b111 6
19
1>
1C
b111 G
#821320000000
0!
0*
09
0>
0C
#821330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#821340000000
0!
0*
09
0>
0C
#821350000000
1!
1*
b1 6
19
1>
1C
b1 G
#821360000000
0!
0*
09
0>
0C
#821370000000
1!
1*
b10 6
19
1>
1C
b10 G
#821380000000
0!
0*
09
0>
0C
#821390000000
1!
1*
b11 6
19
1>
1C
b11 G
#821400000000
0!
0*
09
0>
0C
#821410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#821420000000
0!
0*
09
0>
0C
#821430000000
1!
1*
b101 6
19
1>
1C
b101 G
#821440000000
0!
0*
09
0>
0C
#821450000000
1!
1*
b110 6
19
1>
1C
b110 G
#821460000000
0!
0*
09
0>
0C
#821470000000
1!
1*
b111 6
19
1>
1C
b111 G
#821480000000
0!
1"
0*
1+
09
1:
0>
0C
#821490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#821500000000
0!
0*
09
0>
0C
#821510000000
1!
1*
b1 6
19
1>
1C
b1 G
#821520000000
0!
0*
09
0>
0C
#821530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#821540000000
0!
0*
09
0>
0C
#821550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#821560000000
0!
0*
09
0>
0C
#821570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#821580000000
0!
0*
09
0>
0C
#821590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#821600000000
0!
0#
0*
0,
09
0>
0?
0C
#821610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#821620000000
0!
0*
09
0>
0C
#821630000000
1!
1*
19
1>
1C
#821640000000
0!
0*
09
0>
0C
#821650000000
1!
1*
19
1>
1C
#821660000000
0!
0*
09
0>
0C
#821670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#821680000000
0!
0*
09
0>
0C
#821690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#821700000000
0!
0*
09
0>
0C
#821710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#821720000000
0!
0*
09
0>
0C
#821730000000
1!
1*
b10 6
19
1>
1C
b10 G
#821740000000
0!
0*
09
0>
0C
#821750000000
1!
1*
b11 6
19
1>
1C
b11 G
#821760000000
0!
0*
09
0>
0C
#821770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#821780000000
0!
0*
09
0>
0C
#821790000000
1!
1*
b101 6
19
1>
1C
b101 G
#821800000000
0!
0*
09
0>
0C
#821810000000
1!
1*
b110 6
19
1>
1C
b110 G
#821820000000
0!
0*
09
0>
0C
#821830000000
1!
1*
b111 6
19
1>
1C
b111 G
#821840000000
0!
0*
09
0>
0C
#821850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#821860000000
0!
0*
09
0>
0C
#821870000000
1!
1*
b1 6
19
1>
1C
b1 G
#821880000000
0!
0*
09
0>
0C
#821890000000
1!
1*
b10 6
19
1>
1C
b10 G
#821900000000
0!
0*
09
0>
0C
#821910000000
1!
1*
b11 6
19
1>
1C
b11 G
#821920000000
0!
0*
09
0>
0C
#821930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#821940000000
0!
0*
09
0>
0C
#821950000000
1!
1*
b101 6
19
1>
1C
b101 G
#821960000000
0!
0*
09
0>
0C
#821970000000
1!
1*
b110 6
19
1>
1C
b110 G
#821980000000
0!
0*
09
0>
0C
#821990000000
1!
1*
b111 6
19
1>
1C
b111 G
#822000000000
0!
0*
09
0>
0C
#822010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#822020000000
0!
0*
09
0>
0C
#822030000000
1!
1*
b1 6
19
1>
1C
b1 G
#822040000000
0!
0*
09
0>
0C
#822050000000
1!
1*
b10 6
19
1>
1C
b10 G
#822060000000
0!
0*
09
0>
0C
#822070000000
1!
1*
b11 6
19
1>
1C
b11 G
#822080000000
0!
0*
09
0>
0C
#822090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#822100000000
0!
0*
09
0>
0C
#822110000000
1!
1*
b101 6
19
1>
1C
b101 G
#822120000000
0!
0*
09
0>
0C
#822130000000
1!
1*
b110 6
19
1>
1C
b110 G
#822140000000
0!
0*
09
0>
0C
#822150000000
1!
1*
b111 6
19
1>
1C
b111 G
#822160000000
0!
1"
0*
1+
09
1:
0>
0C
#822170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#822180000000
0!
0*
09
0>
0C
#822190000000
1!
1*
b1 6
19
1>
1C
b1 G
#822200000000
0!
0*
09
0>
0C
#822210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#822220000000
0!
0*
09
0>
0C
#822230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#822240000000
0!
0*
09
0>
0C
#822250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#822260000000
0!
0*
09
0>
0C
#822270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#822280000000
0!
0#
0*
0,
09
0>
0?
0C
#822290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#822300000000
0!
0*
09
0>
0C
#822310000000
1!
1*
19
1>
1C
#822320000000
0!
0*
09
0>
0C
#822330000000
1!
1*
19
1>
1C
#822340000000
0!
0*
09
0>
0C
#822350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#822360000000
0!
0*
09
0>
0C
#822370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#822380000000
0!
0*
09
0>
0C
#822390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#822400000000
0!
0*
09
0>
0C
#822410000000
1!
1*
b10 6
19
1>
1C
b10 G
#822420000000
0!
0*
09
0>
0C
#822430000000
1!
1*
b11 6
19
1>
1C
b11 G
#822440000000
0!
0*
09
0>
0C
#822450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#822460000000
0!
0*
09
0>
0C
#822470000000
1!
1*
b101 6
19
1>
1C
b101 G
#822480000000
0!
0*
09
0>
0C
#822490000000
1!
1*
b110 6
19
1>
1C
b110 G
#822500000000
0!
0*
09
0>
0C
#822510000000
1!
1*
b111 6
19
1>
1C
b111 G
#822520000000
0!
0*
09
0>
0C
#822530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#822540000000
0!
0*
09
0>
0C
#822550000000
1!
1*
b1 6
19
1>
1C
b1 G
#822560000000
0!
0*
09
0>
0C
#822570000000
1!
1*
b10 6
19
1>
1C
b10 G
#822580000000
0!
0*
09
0>
0C
#822590000000
1!
1*
b11 6
19
1>
1C
b11 G
#822600000000
0!
0*
09
0>
0C
#822610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#822620000000
0!
0*
09
0>
0C
#822630000000
1!
1*
b101 6
19
1>
1C
b101 G
#822640000000
0!
0*
09
0>
0C
#822650000000
1!
1*
b110 6
19
1>
1C
b110 G
#822660000000
0!
0*
09
0>
0C
#822670000000
1!
1*
b111 6
19
1>
1C
b111 G
#822680000000
0!
0*
09
0>
0C
#822690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#822700000000
0!
0*
09
0>
0C
#822710000000
1!
1*
b1 6
19
1>
1C
b1 G
#822720000000
0!
0*
09
0>
0C
#822730000000
1!
1*
b10 6
19
1>
1C
b10 G
#822740000000
0!
0*
09
0>
0C
#822750000000
1!
1*
b11 6
19
1>
1C
b11 G
#822760000000
0!
0*
09
0>
0C
#822770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#822780000000
0!
0*
09
0>
0C
#822790000000
1!
1*
b101 6
19
1>
1C
b101 G
#822800000000
0!
0*
09
0>
0C
#822810000000
1!
1*
b110 6
19
1>
1C
b110 G
#822820000000
0!
0*
09
0>
0C
#822830000000
1!
1*
b111 6
19
1>
1C
b111 G
#822840000000
0!
1"
0*
1+
09
1:
0>
0C
#822850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#822860000000
0!
0*
09
0>
0C
#822870000000
1!
1*
b1 6
19
1>
1C
b1 G
#822880000000
0!
0*
09
0>
0C
#822890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#822900000000
0!
0*
09
0>
0C
#822910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#822920000000
0!
0*
09
0>
0C
#822930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#822940000000
0!
0*
09
0>
0C
#822950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#822960000000
0!
0#
0*
0,
09
0>
0?
0C
#822970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#822980000000
0!
0*
09
0>
0C
#822990000000
1!
1*
19
1>
1C
#823000000000
0!
0*
09
0>
0C
#823010000000
1!
1*
19
1>
1C
#823020000000
0!
0*
09
0>
0C
#823030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#823040000000
0!
0*
09
0>
0C
#823050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#823060000000
0!
0*
09
0>
0C
#823070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#823080000000
0!
0*
09
0>
0C
#823090000000
1!
1*
b10 6
19
1>
1C
b10 G
#823100000000
0!
0*
09
0>
0C
#823110000000
1!
1*
b11 6
19
1>
1C
b11 G
#823120000000
0!
0*
09
0>
0C
#823130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#823140000000
0!
0*
09
0>
0C
#823150000000
1!
1*
b101 6
19
1>
1C
b101 G
#823160000000
0!
0*
09
0>
0C
#823170000000
1!
1*
b110 6
19
1>
1C
b110 G
#823180000000
0!
0*
09
0>
0C
#823190000000
1!
1*
b111 6
19
1>
1C
b111 G
#823200000000
0!
0*
09
0>
0C
#823210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#823220000000
0!
0*
09
0>
0C
#823230000000
1!
1*
b1 6
19
1>
1C
b1 G
#823240000000
0!
0*
09
0>
0C
#823250000000
1!
1*
b10 6
19
1>
1C
b10 G
#823260000000
0!
0*
09
0>
0C
#823270000000
1!
1*
b11 6
19
1>
1C
b11 G
#823280000000
0!
0*
09
0>
0C
#823290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#823300000000
0!
0*
09
0>
0C
#823310000000
1!
1*
b101 6
19
1>
1C
b101 G
#823320000000
0!
0*
09
0>
0C
#823330000000
1!
1*
b110 6
19
1>
1C
b110 G
#823340000000
0!
0*
09
0>
0C
#823350000000
1!
1*
b111 6
19
1>
1C
b111 G
#823360000000
0!
0*
09
0>
0C
#823370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#823380000000
0!
0*
09
0>
0C
#823390000000
1!
1*
b1 6
19
1>
1C
b1 G
#823400000000
0!
0*
09
0>
0C
#823410000000
1!
1*
b10 6
19
1>
1C
b10 G
#823420000000
0!
0*
09
0>
0C
#823430000000
1!
1*
b11 6
19
1>
1C
b11 G
#823440000000
0!
0*
09
0>
0C
#823450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#823460000000
0!
0*
09
0>
0C
#823470000000
1!
1*
b101 6
19
1>
1C
b101 G
#823480000000
0!
0*
09
0>
0C
#823490000000
1!
1*
b110 6
19
1>
1C
b110 G
#823500000000
0!
0*
09
0>
0C
#823510000000
1!
1*
b111 6
19
1>
1C
b111 G
#823520000000
0!
1"
0*
1+
09
1:
0>
0C
#823530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#823540000000
0!
0*
09
0>
0C
#823550000000
1!
1*
b1 6
19
1>
1C
b1 G
#823560000000
0!
0*
09
0>
0C
#823570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#823580000000
0!
0*
09
0>
0C
#823590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#823600000000
0!
0*
09
0>
0C
#823610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#823620000000
0!
0*
09
0>
0C
#823630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#823640000000
0!
0#
0*
0,
09
0>
0?
0C
#823650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#823660000000
0!
0*
09
0>
0C
#823670000000
1!
1*
19
1>
1C
#823680000000
0!
0*
09
0>
0C
#823690000000
1!
1*
19
1>
1C
#823700000000
0!
0*
09
0>
0C
#823710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#823720000000
0!
0*
09
0>
0C
#823730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#823740000000
0!
0*
09
0>
0C
#823750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#823760000000
0!
0*
09
0>
0C
#823770000000
1!
1*
b10 6
19
1>
1C
b10 G
#823780000000
0!
0*
09
0>
0C
#823790000000
1!
1*
b11 6
19
1>
1C
b11 G
#823800000000
0!
0*
09
0>
0C
#823810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#823820000000
0!
0*
09
0>
0C
#823830000000
1!
1*
b101 6
19
1>
1C
b101 G
#823840000000
0!
0*
09
0>
0C
#823850000000
1!
1*
b110 6
19
1>
1C
b110 G
#823860000000
0!
0*
09
0>
0C
#823870000000
1!
1*
b111 6
19
1>
1C
b111 G
#823880000000
0!
0*
09
0>
0C
#823890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#823900000000
0!
0*
09
0>
0C
#823910000000
1!
1*
b1 6
19
1>
1C
b1 G
#823920000000
0!
0*
09
0>
0C
#823930000000
1!
1*
b10 6
19
1>
1C
b10 G
#823940000000
0!
0*
09
0>
0C
#823950000000
1!
1*
b11 6
19
1>
1C
b11 G
#823960000000
0!
0*
09
0>
0C
#823970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#823980000000
0!
0*
09
0>
0C
#823990000000
1!
1*
b101 6
19
1>
1C
b101 G
#824000000000
0!
0*
09
0>
0C
#824010000000
1!
1*
b110 6
19
1>
1C
b110 G
#824020000000
0!
0*
09
0>
0C
#824030000000
1!
1*
b111 6
19
1>
1C
b111 G
#824040000000
0!
0*
09
0>
0C
#824050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#824060000000
0!
0*
09
0>
0C
#824070000000
1!
1*
b1 6
19
1>
1C
b1 G
#824080000000
0!
0*
09
0>
0C
#824090000000
1!
1*
b10 6
19
1>
1C
b10 G
#824100000000
0!
0*
09
0>
0C
#824110000000
1!
1*
b11 6
19
1>
1C
b11 G
#824120000000
0!
0*
09
0>
0C
#824130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#824140000000
0!
0*
09
0>
0C
#824150000000
1!
1*
b101 6
19
1>
1C
b101 G
#824160000000
0!
0*
09
0>
0C
#824170000000
1!
1*
b110 6
19
1>
1C
b110 G
#824180000000
0!
0*
09
0>
0C
#824190000000
1!
1*
b111 6
19
1>
1C
b111 G
#824200000000
0!
1"
0*
1+
09
1:
0>
0C
#824210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#824220000000
0!
0*
09
0>
0C
#824230000000
1!
1*
b1 6
19
1>
1C
b1 G
#824240000000
0!
0*
09
0>
0C
#824250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#824260000000
0!
0*
09
0>
0C
#824270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#824280000000
0!
0*
09
0>
0C
#824290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#824300000000
0!
0*
09
0>
0C
#824310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#824320000000
0!
0#
0*
0,
09
0>
0?
0C
#824330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#824340000000
0!
0*
09
0>
0C
#824350000000
1!
1*
19
1>
1C
#824360000000
0!
0*
09
0>
0C
#824370000000
1!
1*
19
1>
1C
#824380000000
0!
0*
09
0>
0C
#824390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#824400000000
0!
0*
09
0>
0C
#824410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#824420000000
0!
0*
09
0>
0C
#824430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#824440000000
0!
0*
09
0>
0C
#824450000000
1!
1*
b10 6
19
1>
1C
b10 G
#824460000000
0!
0*
09
0>
0C
#824470000000
1!
1*
b11 6
19
1>
1C
b11 G
#824480000000
0!
0*
09
0>
0C
#824490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#824500000000
0!
0*
09
0>
0C
#824510000000
1!
1*
b101 6
19
1>
1C
b101 G
#824520000000
0!
0*
09
0>
0C
#824530000000
1!
1*
b110 6
19
1>
1C
b110 G
#824540000000
0!
0*
09
0>
0C
#824550000000
1!
1*
b111 6
19
1>
1C
b111 G
#824560000000
0!
0*
09
0>
0C
#824570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#824580000000
0!
0*
09
0>
0C
#824590000000
1!
1*
b1 6
19
1>
1C
b1 G
#824600000000
0!
0*
09
0>
0C
#824610000000
1!
1*
b10 6
19
1>
1C
b10 G
#824620000000
0!
0*
09
0>
0C
#824630000000
1!
1*
b11 6
19
1>
1C
b11 G
#824640000000
0!
0*
09
0>
0C
#824650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#824660000000
0!
0*
09
0>
0C
#824670000000
1!
1*
b101 6
19
1>
1C
b101 G
#824680000000
0!
0*
09
0>
0C
#824690000000
1!
1*
b110 6
19
1>
1C
b110 G
#824700000000
0!
0*
09
0>
0C
#824710000000
1!
1*
b111 6
19
1>
1C
b111 G
#824720000000
0!
0*
09
0>
0C
#824730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#824740000000
0!
0*
09
0>
0C
#824750000000
1!
1*
b1 6
19
1>
1C
b1 G
#824760000000
0!
0*
09
0>
0C
#824770000000
1!
1*
b10 6
19
1>
1C
b10 G
#824780000000
0!
0*
09
0>
0C
#824790000000
1!
1*
b11 6
19
1>
1C
b11 G
#824800000000
0!
0*
09
0>
0C
#824810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#824820000000
0!
0*
09
0>
0C
#824830000000
1!
1*
b101 6
19
1>
1C
b101 G
#824840000000
0!
0*
09
0>
0C
#824850000000
1!
1*
b110 6
19
1>
1C
b110 G
#824860000000
0!
0*
09
0>
0C
#824870000000
1!
1*
b111 6
19
1>
1C
b111 G
#824880000000
0!
1"
0*
1+
09
1:
0>
0C
#824890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#824900000000
0!
0*
09
0>
0C
#824910000000
1!
1*
b1 6
19
1>
1C
b1 G
#824920000000
0!
0*
09
0>
0C
#824930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#824940000000
0!
0*
09
0>
0C
#824950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#824960000000
0!
0*
09
0>
0C
#824970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#824980000000
0!
0*
09
0>
0C
#824990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#825000000000
0!
0#
0*
0,
09
0>
0?
0C
#825010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#825020000000
0!
0*
09
0>
0C
#825030000000
1!
1*
19
1>
1C
#825040000000
0!
0*
09
0>
0C
#825050000000
1!
1*
19
1>
1C
#825060000000
0!
0*
09
0>
0C
#825070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#825080000000
0!
0*
09
0>
0C
#825090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#825100000000
0!
0*
09
0>
0C
#825110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#825120000000
0!
0*
09
0>
0C
#825130000000
1!
1*
b10 6
19
1>
1C
b10 G
#825140000000
0!
0*
09
0>
0C
#825150000000
1!
1*
b11 6
19
1>
1C
b11 G
#825160000000
0!
0*
09
0>
0C
#825170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#825180000000
0!
0*
09
0>
0C
#825190000000
1!
1*
b101 6
19
1>
1C
b101 G
#825200000000
0!
0*
09
0>
0C
#825210000000
1!
1*
b110 6
19
1>
1C
b110 G
#825220000000
0!
0*
09
0>
0C
#825230000000
1!
1*
b111 6
19
1>
1C
b111 G
#825240000000
0!
0*
09
0>
0C
#825250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#825260000000
0!
0*
09
0>
0C
#825270000000
1!
1*
b1 6
19
1>
1C
b1 G
#825280000000
0!
0*
09
0>
0C
#825290000000
1!
1*
b10 6
19
1>
1C
b10 G
#825300000000
0!
0*
09
0>
0C
#825310000000
1!
1*
b11 6
19
1>
1C
b11 G
#825320000000
0!
0*
09
0>
0C
#825330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#825340000000
0!
0*
09
0>
0C
#825350000000
1!
1*
b101 6
19
1>
1C
b101 G
#825360000000
0!
0*
09
0>
0C
#825370000000
1!
1*
b110 6
19
1>
1C
b110 G
#825380000000
0!
0*
09
0>
0C
#825390000000
1!
1*
b111 6
19
1>
1C
b111 G
#825400000000
0!
0*
09
0>
0C
#825410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#825420000000
0!
0*
09
0>
0C
#825430000000
1!
1*
b1 6
19
1>
1C
b1 G
#825440000000
0!
0*
09
0>
0C
#825450000000
1!
1*
b10 6
19
1>
1C
b10 G
#825460000000
0!
0*
09
0>
0C
#825470000000
1!
1*
b11 6
19
1>
1C
b11 G
#825480000000
0!
0*
09
0>
0C
#825490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#825500000000
0!
0*
09
0>
0C
#825510000000
1!
1*
b101 6
19
1>
1C
b101 G
#825520000000
0!
0*
09
0>
0C
#825530000000
1!
1*
b110 6
19
1>
1C
b110 G
#825540000000
0!
0*
09
0>
0C
#825550000000
1!
1*
b111 6
19
1>
1C
b111 G
#825560000000
0!
1"
0*
1+
09
1:
0>
0C
#825570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#825580000000
0!
0*
09
0>
0C
#825590000000
1!
1*
b1 6
19
1>
1C
b1 G
#825600000000
0!
0*
09
0>
0C
#825610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#825620000000
0!
0*
09
0>
0C
#825630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#825640000000
0!
0*
09
0>
0C
#825650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#825660000000
0!
0*
09
0>
0C
#825670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#825680000000
0!
0#
0*
0,
09
0>
0?
0C
#825690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#825700000000
0!
0*
09
0>
0C
#825710000000
1!
1*
19
1>
1C
#825720000000
0!
0*
09
0>
0C
#825730000000
1!
1*
19
1>
1C
#825740000000
0!
0*
09
0>
0C
#825750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#825760000000
0!
0*
09
0>
0C
#825770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#825780000000
0!
0*
09
0>
0C
#825790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#825800000000
0!
0*
09
0>
0C
#825810000000
1!
1*
b10 6
19
1>
1C
b10 G
#825820000000
0!
0*
09
0>
0C
#825830000000
1!
1*
b11 6
19
1>
1C
b11 G
#825840000000
0!
0*
09
0>
0C
#825850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#825860000000
0!
0*
09
0>
0C
#825870000000
1!
1*
b101 6
19
1>
1C
b101 G
#825880000000
0!
0*
09
0>
0C
#825890000000
1!
1*
b110 6
19
1>
1C
b110 G
#825900000000
0!
0*
09
0>
0C
#825910000000
1!
1*
b111 6
19
1>
1C
b111 G
#825920000000
0!
0*
09
0>
0C
#825930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#825940000000
0!
0*
09
0>
0C
#825950000000
1!
1*
b1 6
19
1>
1C
b1 G
#825960000000
0!
0*
09
0>
0C
#825970000000
1!
1*
b10 6
19
1>
1C
b10 G
#825980000000
0!
0*
09
0>
0C
#825990000000
1!
1*
b11 6
19
1>
1C
b11 G
#826000000000
0!
0*
09
0>
0C
#826010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#826020000000
0!
0*
09
0>
0C
#826030000000
1!
1*
b101 6
19
1>
1C
b101 G
#826040000000
0!
0*
09
0>
0C
#826050000000
1!
1*
b110 6
19
1>
1C
b110 G
#826060000000
0!
0*
09
0>
0C
#826070000000
1!
1*
b111 6
19
1>
1C
b111 G
#826080000000
0!
0*
09
0>
0C
#826090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#826100000000
0!
0*
09
0>
0C
#826110000000
1!
1*
b1 6
19
1>
1C
b1 G
#826120000000
0!
0*
09
0>
0C
#826130000000
1!
1*
b10 6
19
1>
1C
b10 G
#826140000000
0!
0*
09
0>
0C
#826150000000
1!
1*
b11 6
19
1>
1C
b11 G
#826160000000
0!
0*
09
0>
0C
#826170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#826180000000
0!
0*
09
0>
0C
#826190000000
1!
1*
b101 6
19
1>
1C
b101 G
#826200000000
0!
0*
09
0>
0C
#826210000000
1!
1*
b110 6
19
1>
1C
b110 G
#826220000000
0!
0*
09
0>
0C
#826230000000
1!
1*
b111 6
19
1>
1C
b111 G
#826240000000
0!
1"
0*
1+
09
1:
0>
0C
#826250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#826260000000
0!
0*
09
0>
0C
#826270000000
1!
1*
b1 6
19
1>
1C
b1 G
#826280000000
0!
0*
09
0>
0C
#826290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#826300000000
0!
0*
09
0>
0C
#826310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#826320000000
0!
0*
09
0>
0C
#826330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#826340000000
0!
0*
09
0>
0C
#826350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#826360000000
0!
0#
0*
0,
09
0>
0?
0C
#826370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#826380000000
0!
0*
09
0>
0C
#826390000000
1!
1*
19
1>
1C
#826400000000
0!
0*
09
0>
0C
#826410000000
1!
1*
19
1>
1C
#826420000000
0!
0*
09
0>
0C
#826430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#826440000000
0!
0*
09
0>
0C
#826450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#826460000000
0!
0*
09
0>
0C
#826470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#826480000000
0!
0*
09
0>
0C
#826490000000
1!
1*
b10 6
19
1>
1C
b10 G
#826500000000
0!
0*
09
0>
0C
#826510000000
1!
1*
b11 6
19
1>
1C
b11 G
#826520000000
0!
0*
09
0>
0C
#826530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#826540000000
0!
0*
09
0>
0C
#826550000000
1!
1*
b101 6
19
1>
1C
b101 G
#826560000000
0!
0*
09
0>
0C
#826570000000
1!
1*
b110 6
19
1>
1C
b110 G
#826580000000
0!
0*
09
0>
0C
#826590000000
1!
1*
b111 6
19
1>
1C
b111 G
#826600000000
0!
0*
09
0>
0C
#826610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#826620000000
0!
0*
09
0>
0C
#826630000000
1!
1*
b1 6
19
1>
1C
b1 G
#826640000000
0!
0*
09
0>
0C
#826650000000
1!
1*
b10 6
19
1>
1C
b10 G
#826660000000
0!
0*
09
0>
0C
#826670000000
1!
1*
b11 6
19
1>
1C
b11 G
#826680000000
0!
0*
09
0>
0C
#826690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#826700000000
0!
0*
09
0>
0C
#826710000000
1!
1*
b101 6
19
1>
1C
b101 G
#826720000000
0!
0*
09
0>
0C
#826730000000
1!
1*
b110 6
19
1>
1C
b110 G
#826740000000
0!
0*
09
0>
0C
#826750000000
1!
1*
b111 6
19
1>
1C
b111 G
#826760000000
0!
0*
09
0>
0C
#826770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#826780000000
0!
0*
09
0>
0C
#826790000000
1!
1*
b1 6
19
1>
1C
b1 G
#826800000000
0!
0*
09
0>
0C
#826810000000
1!
1*
b10 6
19
1>
1C
b10 G
#826820000000
0!
0*
09
0>
0C
#826830000000
1!
1*
b11 6
19
1>
1C
b11 G
#826840000000
0!
0*
09
0>
0C
#826850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#826860000000
0!
0*
09
0>
0C
#826870000000
1!
1*
b101 6
19
1>
1C
b101 G
#826880000000
0!
0*
09
0>
0C
#826890000000
1!
1*
b110 6
19
1>
1C
b110 G
#826900000000
0!
0*
09
0>
0C
#826910000000
1!
1*
b111 6
19
1>
1C
b111 G
#826920000000
0!
1"
0*
1+
09
1:
0>
0C
#826930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#826940000000
0!
0*
09
0>
0C
#826950000000
1!
1*
b1 6
19
1>
1C
b1 G
#826960000000
0!
0*
09
0>
0C
#826970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#826980000000
0!
0*
09
0>
0C
#826990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#827000000000
0!
0*
09
0>
0C
#827010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#827020000000
0!
0*
09
0>
0C
#827030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#827040000000
0!
0#
0*
0,
09
0>
0?
0C
#827050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#827060000000
0!
0*
09
0>
0C
#827070000000
1!
1*
19
1>
1C
#827080000000
0!
0*
09
0>
0C
#827090000000
1!
1*
19
1>
1C
#827100000000
0!
0*
09
0>
0C
#827110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#827120000000
0!
0*
09
0>
0C
#827130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#827140000000
0!
0*
09
0>
0C
#827150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#827160000000
0!
0*
09
0>
0C
#827170000000
1!
1*
b10 6
19
1>
1C
b10 G
#827180000000
0!
0*
09
0>
0C
#827190000000
1!
1*
b11 6
19
1>
1C
b11 G
#827200000000
0!
0*
09
0>
0C
#827210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#827220000000
0!
0*
09
0>
0C
#827230000000
1!
1*
b101 6
19
1>
1C
b101 G
#827240000000
0!
0*
09
0>
0C
#827250000000
1!
1*
b110 6
19
1>
1C
b110 G
#827260000000
0!
0*
09
0>
0C
#827270000000
1!
1*
b111 6
19
1>
1C
b111 G
#827280000000
0!
0*
09
0>
0C
#827290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#827300000000
0!
0*
09
0>
0C
#827310000000
1!
1*
b1 6
19
1>
1C
b1 G
#827320000000
0!
0*
09
0>
0C
#827330000000
1!
1*
b10 6
19
1>
1C
b10 G
#827340000000
0!
0*
09
0>
0C
#827350000000
1!
1*
b11 6
19
1>
1C
b11 G
#827360000000
0!
0*
09
0>
0C
#827370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#827380000000
0!
0*
09
0>
0C
#827390000000
1!
1*
b101 6
19
1>
1C
b101 G
#827400000000
0!
0*
09
0>
0C
#827410000000
1!
1*
b110 6
19
1>
1C
b110 G
#827420000000
0!
0*
09
0>
0C
#827430000000
1!
1*
b111 6
19
1>
1C
b111 G
#827440000000
0!
0*
09
0>
0C
#827450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#827460000000
0!
0*
09
0>
0C
#827470000000
1!
1*
b1 6
19
1>
1C
b1 G
#827480000000
0!
0*
09
0>
0C
#827490000000
1!
1*
b10 6
19
1>
1C
b10 G
#827500000000
0!
0*
09
0>
0C
#827510000000
1!
1*
b11 6
19
1>
1C
b11 G
#827520000000
0!
0*
09
0>
0C
#827530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#827540000000
0!
0*
09
0>
0C
#827550000000
1!
1*
b101 6
19
1>
1C
b101 G
#827560000000
0!
0*
09
0>
0C
#827570000000
1!
1*
b110 6
19
1>
1C
b110 G
#827580000000
0!
0*
09
0>
0C
#827590000000
1!
1*
b111 6
19
1>
1C
b111 G
#827600000000
0!
1"
0*
1+
09
1:
0>
0C
#827610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#827620000000
0!
0*
09
0>
0C
#827630000000
1!
1*
b1 6
19
1>
1C
b1 G
#827640000000
0!
0*
09
0>
0C
#827650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#827660000000
0!
0*
09
0>
0C
#827670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#827680000000
0!
0*
09
0>
0C
#827690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#827700000000
0!
0*
09
0>
0C
#827710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#827720000000
0!
0#
0*
0,
09
0>
0?
0C
#827730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#827740000000
0!
0*
09
0>
0C
#827750000000
1!
1*
19
1>
1C
#827760000000
0!
0*
09
0>
0C
#827770000000
1!
1*
19
1>
1C
#827780000000
0!
0*
09
0>
0C
#827790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#827800000000
0!
0*
09
0>
0C
#827810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#827820000000
0!
0*
09
0>
0C
#827830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#827840000000
0!
0*
09
0>
0C
#827850000000
1!
1*
b10 6
19
1>
1C
b10 G
#827860000000
0!
0*
09
0>
0C
#827870000000
1!
1*
b11 6
19
1>
1C
b11 G
#827880000000
0!
0*
09
0>
0C
#827890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#827900000000
0!
0*
09
0>
0C
#827910000000
1!
1*
b101 6
19
1>
1C
b101 G
#827920000000
0!
0*
09
0>
0C
#827930000000
1!
1*
b110 6
19
1>
1C
b110 G
#827940000000
0!
0*
09
0>
0C
#827950000000
1!
1*
b111 6
19
1>
1C
b111 G
#827960000000
0!
0*
09
0>
0C
#827970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#827980000000
0!
0*
09
0>
0C
#827990000000
1!
1*
b1 6
19
1>
1C
b1 G
#828000000000
0!
0*
09
0>
0C
#828010000000
1!
1*
b10 6
19
1>
1C
b10 G
#828020000000
0!
0*
09
0>
0C
#828030000000
1!
1*
b11 6
19
1>
1C
b11 G
#828040000000
0!
0*
09
0>
0C
#828050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#828060000000
0!
0*
09
0>
0C
#828070000000
1!
1*
b101 6
19
1>
1C
b101 G
#828080000000
0!
0*
09
0>
0C
#828090000000
1!
1*
b110 6
19
1>
1C
b110 G
#828100000000
0!
0*
09
0>
0C
#828110000000
1!
1*
b111 6
19
1>
1C
b111 G
#828120000000
0!
0*
09
0>
0C
#828130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#828140000000
0!
0*
09
0>
0C
#828150000000
1!
1*
b1 6
19
1>
1C
b1 G
#828160000000
0!
0*
09
0>
0C
#828170000000
1!
1*
b10 6
19
1>
1C
b10 G
#828180000000
0!
0*
09
0>
0C
#828190000000
1!
1*
b11 6
19
1>
1C
b11 G
#828200000000
0!
0*
09
0>
0C
#828210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#828220000000
0!
0*
09
0>
0C
#828230000000
1!
1*
b101 6
19
1>
1C
b101 G
#828240000000
0!
0*
09
0>
0C
#828250000000
1!
1*
b110 6
19
1>
1C
b110 G
#828260000000
0!
0*
09
0>
0C
#828270000000
1!
1*
b111 6
19
1>
1C
b111 G
#828280000000
0!
1"
0*
1+
09
1:
0>
0C
#828290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#828300000000
0!
0*
09
0>
0C
#828310000000
1!
1*
b1 6
19
1>
1C
b1 G
#828320000000
0!
0*
09
0>
0C
#828330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#828340000000
0!
0*
09
0>
0C
#828350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#828360000000
0!
0*
09
0>
0C
#828370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#828380000000
0!
0*
09
0>
0C
#828390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#828400000000
0!
0#
0*
0,
09
0>
0?
0C
#828410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#828420000000
0!
0*
09
0>
0C
#828430000000
1!
1*
19
1>
1C
#828440000000
0!
0*
09
0>
0C
#828450000000
1!
1*
19
1>
1C
#828460000000
0!
0*
09
0>
0C
#828470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#828480000000
0!
0*
09
0>
0C
#828490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#828500000000
0!
0*
09
0>
0C
#828510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#828520000000
0!
0*
09
0>
0C
#828530000000
1!
1*
b10 6
19
1>
1C
b10 G
#828540000000
0!
0*
09
0>
0C
#828550000000
1!
1*
b11 6
19
1>
1C
b11 G
#828560000000
0!
0*
09
0>
0C
#828570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#828580000000
0!
0*
09
0>
0C
#828590000000
1!
1*
b101 6
19
1>
1C
b101 G
#828600000000
0!
0*
09
0>
0C
#828610000000
1!
1*
b110 6
19
1>
1C
b110 G
#828620000000
0!
0*
09
0>
0C
#828630000000
1!
1*
b111 6
19
1>
1C
b111 G
#828640000000
0!
0*
09
0>
0C
#828650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#828660000000
0!
0*
09
0>
0C
#828670000000
1!
1*
b1 6
19
1>
1C
b1 G
#828680000000
0!
0*
09
0>
0C
#828690000000
1!
1*
b10 6
19
1>
1C
b10 G
#828700000000
0!
0*
09
0>
0C
#828710000000
1!
1*
b11 6
19
1>
1C
b11 G
#828720000000
0!
0*
09
0>
0C
#828730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#828740000000
0!
0*
09
0>
0C
#828750000000
1!
1*
b101 6
19
1>
1C
b101 G
#828760000000
0!
0*
09
0>
0C
#828770000000
1!
1*
b110 6
19
1>
1C
b110 G
#828780000000
0!
0*
09
0>
0C
#828790000000
1!
1*
b111 6
19
1>
1C
b111 G
#828800000000
0!
0*
09
0>
0C
#828810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#828820000000
0!
0*
09
0>
0C
#828830000000
1!
1*
b1 6
19
1>
1C
b1 G
#828840000000
0!
0*
09
0>
0C
#828850000000
1!
1*
b10 6
19
1>
1C
b10 G
#828860000000
0!
0*
09
0>
0C
#828870000000
1!
1*
b11 6
19
1>
1C
b11 G
#828880000000
0!
0*
09
0>
0C
#828890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#828900000000
0!
0*
09
0>
0C
#828910000000
1!
1*
b101 6
19
1>
1C
b101 G
#828920000000
0!
0*
09
0>
0C
#828930000000
1!
1*
b110 6
19
1>
1C
b110 G
#828940000000
0!
0*
09
0>
0C
#828950000000
1!
1*
b111 6
19
1>
1C
b111 G
#828960000000
0!
1"
0*
1+
09
1:
0>
0C
#828970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#828980000000
0!
0*
09
0>
0C
#828990000000
1!
1*
b1 6
19
1>
1C
b1 G
#829000000000
0!
0*
09
0>
0C
#829010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#829020000000
0!
0*
09
0>
0C
#829030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#829040000000
0!
0*
09
0>
0C
#829050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#829060000000
0!
0*
09
0>
0C
#829070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#829080000000
0!
0#
0*
0,
09
0>
0?
0C
#829090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#829100000000
0!
0*
09
0>
0C
#829110000000
1!
1*
19
1>
1C
#829120000000
0!
0*
09
0>
0C
#829130000000
1!
1*
19
1>
1C
#829140000000
0!
0*
09
0>
0C
#829150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#829160000000
0!
0*
09
0>
0C
#829170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#829180000000
0!
0*
09
0>
0C
#829190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#829200000000
0!
0*
09
0>
0C
#829210000000
1!
1*
b10 6
19
1>
1C
b10 G
#829220000000
0!
0*
09
0>
0C
#829230000000
1!
1*
b11 6
19
1>
1C
b11 G
#829240000000
0!
0*
09
0>
0C
#829250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#829260000000
0!
0*
09
0>
0C
#829270000000
1!
1*
b101 6
19
1>
1C
b101 G
#829280000000
0!
0*
09
0>
0C
#829290000000
1!
1*
b110 6
19
1>
1C
b110 G
#829300000000
0!
0*
09
0>
0C
#829310000000
1!
1*
b111 6
19
1>
1C
b111 G
#829320000000
0!
0*
09
0>
0C
#829330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#829340000000
0!
0*
09
0>
0C
#829350000000
1!
1*
b1 6
19
1>
1C
b1 G
#829360000000
0!
0*
09
0>
0C
#829370000000
1!
1*
b10 6
19
1>
1C
b10 G
#829380000000
0!
0*
09
0>
0C
#829390000000
1!
1*
b11 6
19
1>
1C
b11 G
#829400000000
0!
0*
09
0>
0C
#829410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#829420000000
0!
0*
09
0>
0C
#829430000000
1!
1*
b101 6
19
1>
1C
b101 G
#829440000000
0!
0*
09
0>
0C
#829450000000
1!
1*
b110 6
19
1>
1C
b110 G
#829460000000
0!
0*
09
0>
0C
#829470000000
1!
1*
b111 6
19
1>
1C
b111 G
#829480000000
0!
0*
09
0>
0C
#829490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#829500000000
0!
0*
09
0>
0C
#829510000000
1!
1*
b1 6
19
1>
1C
b1 G
#829520000000
0!
0*
09
0>
0C
#829530000000
1!
1*
b10 6
19
1>
1C
b10 G
#829540000000
0!
0*
09
0>
0C
#829550000000
1!
1*
b11 6
19
1>
1C
b11 G
#829560000000
0!
0*
09
0>
0C
#829570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#829580000000
0!
0*
09
0>
0C
#829590000000
1!
1*
b101 6
19
1>
1C
b101 G
#829600000000
0!
0*
09
0>
0C
#829610000000
1!
1*
b110 6
19
1>
1C
b110 G
#829620000000
0!
0*
09
0>
0C
#829630000000
1!
1*
b111 6
19
1>
1C
b111 G
#829640000000
0!
1"
0*
1+
09
1:
0>
0C
#829650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#829660000000
0!
0*
09
0>
0C
#829670000000
1!
1*
b1 6
19
1>
1C
b1 G
#829680000000
0!
0*
09
0>
0C
#829690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#829700000000
0!
0*
09
0>
0C
#829710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#829720000000
0!
0*
09
0>
0C
#829730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#829740000000
0!
0*
09
0>
0C
#829750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#829760000000
0!
0#
0*
0,
09
0>
0?
0C
#829770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#829780000000
0!
0*
09
0>
0C
#829790000000
1!
1*
19
1>
1C
#829800000000
0!
0*
09
0>
0C
#829810000000
1!
1*
19
1>
1C
#829820000000
0!
0*
09
0>
0C
#829830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#829840000000
0!
0*
09
0>
0C
#829850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#829860000000
0!
0*
09
0>
0C
#829870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#829880000000
0!
0*
09
0>
0C
#829890000000
1!
1*
b10 6
19
1>
1C
b10 G
#829900000000
0!
0*
09
0>
0C
#829910000000
1!
1*
b11 6
19
1>
1C
b11 G
#829920000000
0!
0*
09
0>
0C
#829930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#829940000000
0!
0*
09
0>
0C
#829950000000
1!
1*
b101 6
19
1>
1C
b101 G
#829960000000
0!
0*
09
0>
0C
#829970000000
1!
1*
b110 6
19
1>
1C
b110 G
#829980000000
0!
0*
09
0>
0C
#829990000000
1!
1*
b111 6
19
1>
1C
b111 G
#830000000000
0!
0*
09
0>
0C
#830010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#830020000000
0!
0*
09
0>
0C
#830030000000
1!
1*
b1 6
19
1>
1C
b1 G
#830040000000
0!
0*
09
0>
0C
#830050000000
1!
1*
b10 6
19
1>
1C
b10 G
#830060000000
0!
0*
09
0>
0C
#830070000000
1!
1*
b11 6
19
1>
1C
b11 G
#830080000000
0!
0*
09
0>
0C
#830090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#830100000000
0!
0*
09
0>
0C
#830110000000
1!
1*
b101 6
19
1>
1C
b101 G
#830120000000
0!
0*
09
0>
0C
#830130000000
1!
1*
b110 6
19
1>
1C
b110 G
#830140000000
0!
0*
09
0>
0C
#830150000000
1!
1*
b111 6
19
1>
1C
b111 G
#830160000000
0!
0*
09
0>
0C
#830170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#830180000000
0!
0*
09
0>
0C
#830190000000
1!
1*
b1 6
19
1>
1C
b1 G
#830200000000
0!
0*
09
0>
0C
#830210000000
1!
1*
b10 6
19
1>
1C
b10 G
#830220000000
0!
0*
09
0>
0C
#830230000000
1!
1*
b11 6
19
1>
1C
b11 G
#830240000000
0!
0*
09
0>
0C
#830250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#830260000000
0!
0*
09
0>
0C
#830270000000
1!
1*
b101 6
19
1>
1C
b101 G
#830280000000
0!
0*
09
0>
0C
#830290000000
1!
1*
b110 6
19
1>
1C
b110 G
#830300000000
0!
0*
09
0>
0C
#830310000000
1!
1*
b111 6
19
1>
1C
b111 G
#830320000000
0!
1"
0*
1+
09
1:
0>
0C
#830330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#830340000000
0!
0*
09
0>
0C
#830350000000
1!
1*
b1 6
19
1>
1C
b1 G
#830360000000
0!
0*
09
0>
0C
#830370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#830380000000
0!
0*
09
0>
0C
#830390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#830400000000
0!
0*
09
0>
0C
#830410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#830420000000
0!
0*
09
0>
0C
#830430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#830440000000
0!
0#
0*
0,
09
0>
0?
0C
#830450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#830460000000
0!
0*
09
0>
0C
#830470000000
1!
1*
19
1>
1C
#830480000000
0!
0*
09
0>
0C
#830490000000
1!
1*
19
1>
1C
#830500000000
0!
0*
09
0>
0C
#830510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#830520000000
0!
0*
09
0>
0C
#830530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#830540000000
0!
0*
09
0>
0C
#830550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#830560000000
0!
0*
09
0>
0C
#830570000000
1!
1*
b10 6
19
1>
1C
b10 G
#830580000000
0!
0*
09
0>
0C
#830590000000
1!
1*
b11 6
19
1>
1C
b11 G
#830600000000
0!
0*
09
0>
0C
#830610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#830620000000
0!
0*
09
0>
0C
#830630000000
1!
1*
b101 6
19
1>
1C
b101 G
#830640000000
0!
0*
09
0>
0C
#830650000000
1!
1*
b110 6
19
1>
1C
b110 G
#830660000000
0!
0*
09
0>
0C
#830670000000
1!
1*
b111 6
19
1>
1C
b111 G
#830680000000
0!
0*
09
0>
0C
#830690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#830700000000
0!
0*
09
0>
0C
#830710000000
1!
1*
b1 6
19
1>
1C
b1 G
#830720000000
0!
0*
09
0>
0C
#830730000000
1!
1*
b10 6
19
1>
1C
b10 G
#830740000000
0!
0*
09
0>
0C
#830750000000
1!
1*
b11 6
19
1>
1C
b11 G
#830760000000
0!
0*
09
0>
0C
#830770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#830780000000
0!
0*
09
0>
0C
#830790000000
1!
1*
b101 6
19
1>
1C
b101 G
#830800000000
0!
0*
09
0>
0C
#830810000000
1!
1*
b110 6
19
1>
1C
b110 G
#830820000000
0!
0*
09
0>
0C
#830830000000
1!
1*
b111 6
19
1>
1C
b111 G
#830840000000
0!
0*
09
0>
0C
#830850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#830860000000
0!
0*
09
0>
0C
#830870000000
1!
1*
b1 6
19
1>
1C
b1 G
#830880000000
0!
0*
09
0>
0C
#830890000000
1!
1*
b10 6
19
1>
1C
b10 G
#830900000000
0!
0*
09
0>
0C
#830910000000
1!
1*
b11 6
19
1>
1C
b11 G
#830920000000
0!
0*
09
0>
0C
#830930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#830940000000
0!
0*
09
0>
0C
#830950000000
1!
1*
b101 6
19
1>
1C
b101 G
#830960000000
0!
0*
09
0>
0C
#830970000000
1!
1*
b110 6
19
1>
1C
b110 G
#830980000000
0!
0*
09
0>
0C
#830990000000
1!
1*
b111 6
19
1>
1C
b111 G
#831000000000
0!
1"
0*
1+
09
1:
0>
0C
#831010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#831020000000
0!
0*
09
0>
0C
#831030000000
1!
1*
b1 6
19
1>
1C
b1 G
#831040000000
0!
0*
09
0>
0C
#831050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#831060000000
0!
0*
09
0>
0C
#831070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#831080000000
0!
0*
09
0>
0C
#831090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#831100000000
0!
0*
09
0>
0C
#831110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#831120000000
0!
0#
0*
0,
09
0>
0?
0C
#831130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#831140000000
0!
0*
09
0>
0C
#831150000000
1!
1*
19
1>
1C
#831160000000
0!
0*
09
0>
0C
#831170000000
1!
1*
19
1>
1C
#831180000000
0!
0*
09
0>
0C
#831190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#831200000000
0!
0*
09
0>
0C
#831210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#831220000000
0!
0*
09
0>
0C
#831230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#831240000000
0!
0*
09
0>
0C
#831250000000
1!
1*
b10 6
19
1>
1C
b10 G
#831260000000
0!
0*
09
0>
0C
#831270000000
1!
1*
b11 6
19
1>
1C
b11 G
#831280000000
0!
0*
09
0>
0C
#831290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#831300000000
0!
0*
09
0>
0C
#831310000000
1!
1*
b101 6
19
1>
1C
b101 G
#831320000000
0!
0*
09
0>
0C
#831330000000
1!
1*
b110 6
19
1>
1C
b110 G
#831340000000
0!
0*
09
0>
0C
#831350000000
1!
1*
b111 6
19
1>
1C
b111 G
#831360000000
0!
0*
09
0>
0C
#831370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#831380000000
0!
0*
09
0>
0C
#831390000000
1!
1*
b1 6
19
1>
1C
b1 G
#831400000000
0!
0*
09
0>
0C
#831410000000
1!
1*
b10 6
19
1>
1C
b10 G
#831420000000
0!
0*
09
0>
0C
#831430000000
1!
1*
b11 6
19
1>
1C
b11 G
#831440000000
0!
0*
09
0>
0C
#831450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#831460000000
0!
0*
09
0>
0C
#831470000000
1!
1*
b101 6
19
1>
1C
b101 G
#831480000000
0!
0*
09
0>
0C
#831490000000
1!
1*
b110 6
19
1>
1C
b110 G
#831500000000
0!
0*
09
0>
0C
#831510000000
1!
1*
b111 6
19
1>
1C
b111 G
#831520000000
0!
0*
09
0>
0C
#831530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#831540000000
0!
0*
09
0>
0C
#831550000000
1!
1*
b1 6
19
1>
1C
b1 G
#831560000000
0!
0*
09
0>
0C
#831570000000
1!
1*
b10 6
19
1>
1C
b10 G
#831580000000
0!
0*
09
0>
0C
#831590000000
1!
1*
b11 6
19
1>
1C
b11 G
#831600000000
0!
0*
09
0>
0C
#831610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#831620000000
0!
0*
09
0>
0C
#831630000000
1!
1*
b101 6
19
1>
1C
b101 G
#831640000000
0!
0*
09
0>
0C
#831650000000
1!
1*
b110 6
19
1>
1C
b110 G
#831660000000
0!
0*
09
0>
0C
#831670000000
1!
1*
b111 6
19
1>
1C
b111 G
#831680000000
0!
1"
0*
1+
09
1:
0>
0C
#831690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#831700000000
0!
0*
09
0>
0C
#831710000000
1!
1*
b1 6
19
1>
1C
b1 G
#831720000000
0!
0*
09
0>
0C
#831730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#831740000000
0!
0*
09
0>
0C
#831750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#831760000000
0!
0*
09
0>
0C
#831770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#831780000000
0!
0*
09
0>
0C
#831790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#831800000000
0!
0#
0*
0,
09
0>
0?
0C
#831810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#831820000000
0!
0*
09
0>
0C
#831830000000
1!
1*
19
1>
1C
#831840000000
0!
0*
09
0>
0C
#831850000000
1!
1*
19
1>
1C
#831860000000
0!
0*
09
0>
0C
#831870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#831880000000
0!
0*
09
0>
0C
#831890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#831900000000
0!
0*
09
0>
0C
#831910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#831920000000
0!
0*
09
0>
0C
#831930000000
1!
1*
b10 6
19
1>
1C
b10 G
#831940000000
0!
0*
09
0>
0C
#831950000000
1!
1*
b11 6
19
1>
1C
b11 G
#831960000000
0!
0*
09
0>
0C
#831970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#831980000000
0!
0*
09
0>
0C
#831990000000
1!
1*
b101 6
19
1>
1C
b101 G
#832000000000
0!
0*
09
0>
0C
#832010000000
1!
1*
b110 6
19
1>
1C
b110 G
#832020000000
0!
0*
09
0>
0C
#832030000000
1!
1*
b111 6
19
1>
1C
b111 G
#832040000000
0!
0*
09
0>
0C
#832050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#832060000000
0!
0*
09
0>
0C
#832070000000
1!
1*
b1 6
19
1>
1C
b1 G
#832080000000
0!
0*
09
0>
0C
#832090000000
1!
1*
b10 6
19
1>
1C
b10 G
#832100000000
0!
0*
09
0>
0C
#832110000000
1!
1*
b11 6
19
1>
1C
b11 G
#832120000000
0!
0*
09
0>
0C
#832130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#832140000000
0!
0*
09
0>
0C
#832150000000
1!
1*
b101 6
19
1>
1C
b101 G
#832160000000
0!
0*
09
0>
0C
#832170000000
1!
1*
b110 6
19
1>
1C
b110 G
#832180000000
0!
0*
09
0>
0C
#832190000000
1!
1*
b111 6
19
1>
1C
b111 G
#832200000000
0!
0*
09
0>
0C
#832210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#832220000000
0!
0*
09
0>
0C
#832230000000
1!
1*
b1 6
19
1>
1C
b1 G
#832240000000
0!
0*
09
0>
0C
#832250000000
1!
1*
b10 6
19
1>
1C
b10 G
#832260000000
0!
0*
09
0>
0C
#832270000000
1!
1*
b11 6
19
1>
1C
b11 G
#832280000000
0!
0*
09
0>
0C
#832290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#832300000000
0!
0*
09
0>
0C
#832310000000
1!
1*
b101 6
19
1>
1C
b101 G
#832320000000
0!
0*
09
0>
0C
#832330000000
1!
1*
b110 6
19
1>
1C
b110 G
#832340000000
0!
0*
09
0>
0C
#832350000000
1!
1*
b111 6
19
1>
1C
b111 G
#832360000000
0!
1"
0*
1+
09
1:
0>
0C
#832370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#832380000000
0!
0*
09
0>
0C
#832390000000
1!
1*
b1 6
19
1>
1C
b1 G
#832400000000
0!
0*
09
0>
0C
#832410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#832420000000
0!
0*
09
0>
0C
#832430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#832440000000
0!
0*
09
0>
0C
#832450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#832460000000
0!
0*
09
0>
0C
#832470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#832480000000
0!
0#
0*
0,
09
0>
0?
0C
#832490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#832500000000
0!
0*
09
0>
0C
#832510000000
1!
1*
19
1>
1C
#832520000000
0!
0*
09
0>
0C
#832530000000
1!
1*
19
1>
1C
#832540000000
0!
0*
09
0>
0C
#832550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#832560000000
0!
0*
09
0>
0C
#832570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#832580000000
0!
0*
09
0>
0C
#832590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#832600000000
0!
0*
09
0>
0C
#832610000000
1!
1*
b10 6
19
1>
1C
b10 G
#832620000000
0!
0*
09
0>
0C
#832630000000
1!
1*
b11 6
19
1>
1C
b11 G
#832640000000
0!
0*
09
0>
0C
#832650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#832660000000
0!
0*
09
0>
0C
#832670000000
1!
1*
b101 6
19
1>
1C
b101 G
#832680000000
0!
0*
09
0>
0C
#832690000000
1!
1*
b110 6
19
1>
1C
b110 G
#832700000000
0!
0*
09
0>
0C
#832710000000
1!
1*
b111 6
19
1>
1C
b111 G
#832720000000
0!
0*
09
0>
0C
#832730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#832740000000
0!
0*
09
0>
0C
#832750000000
1!
1*
b1 6
19
1>
1C
b1 G
#832760000000
0!
0*
09
0>
0C
#832770000000
1!
1*
b10 6
19
1>
1C
b10 G
#832780000000
0!
0*
09
0>
0C
#832790000000
1!
1*
b11 6
19
1>
1C
b11 G
#832800000000
0!
0*
09
0>
0C
#832810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#832820000000
0!
0*
09
0>
0C
#832830000000
1!
1*
b101 6
19
1>
1C
b101 G
#832840000000
0!
0*
09
0>
0C
#832850000000
1!
1*
b110 6
19
1>
1C
b110 G
#832860000000
0!
0*
09
0>
0C
#832870000000
1!
1*
b111 6
19
1>
1C
b111 G
#832880000000
0!
0*
09
0>
0C
#832890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#832900000000
0!
0*
09
0>
0C
#832910000000
1!
1*
b1 6
19
1>
1C
b1 G
#832920000000
0!
0*
09
0>
0C
#832930000000
1!
1*
b10 6
19
1>
1C
b10 G
#832940000000
0!
0*
09
0>
0C
#832950000000
1!
1*
b11 6
19
1>
1C
b11 G
#832960000000
0!
0*
09
0>
0C
#832970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#832980000000
0!
0*
09
0>
0C
#832990000000
1!
1*
b101 6
19
1>
1C
b101 G
#833000000000
0!
0*
09
0>
0C
#833010000000
1!
1*
b110 6
19
1>
1C
b110 G
#833020000000
0!
0*
09
0>
0C
#833030000000
1!
1*
b111 6
19
1>
1C
b111 G
#833040000000
0!
1"
0*
1+
09
1:
0>
0C
#833050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#833060000000
0!
0*
09
0>
0C
#833070000000
1!
1*
b1 6
19
1>
1C
b1 G
#833080000000
0!
0*
09
0>
0C
#833090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#833100000000
0!
0*
09
0>
0C
#833110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#833120000000
0!
0*
09
0>
0C
#833130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#833140000000
0!
0*
09
0>
0C
#833150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#833160000000
0!
0#
0*
0,
09
0>
0?
0C
#833170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#833180000000
0!
0*
09
0>
0C
#833190000000
1!
1*
19
1>
1C
#833200000000
0!
0*
09
0>
0C
#833210000000
1!
1*
19
1>
1C
#833220000000
0!
0*
09
0>
0C
#833230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#833240000000
0!
0*
09
0>
0C
#833250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#833260000000
0!
0*
09
0>
0C
#833270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#833280000000
0!
0*
09
0>
0C
#833290000000
1!
1*
b10 6
19
1>
1C
b10 G
#833300000000
0!
0*
09
0>
0C
#833310000000
1!
1*
b11 6
19
1>
1C
b11 G
#833320000000
0!
0*
09
0>
0C
#833330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#833340000000
0!
0*
09
0>
0C
#833350000000
1!
1*
b101 6
19
1>
1C
b101 G
#833360000000
0!
0*
09
0>
0C
#833370000000
1!
1*
b110 6
19
1>
1C
b110 G
#833380000000
0!
0*
09
0>
0C
#833390000000
1!
1*
b111 6
19
1>
1C
b111 G
#833400000000
0!
0*
09
0>
0C
#833410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#833420000000
0!
0*
09
0>
0C
#833430000000
1!
1*
b1 6
19
1>
1C
b1 G
#833440000000
0!
0*
09
0>
0C
#833450000000
1!
1*
b10 6
19
1>
1C
b10 G
#833460000000
0!
0*
09
0>
0C
#833470000000
1!
1*
b11 6
19
1>
1C
b11 G
#833480000000
0!
0*
09
0>
0C
#833490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#833500000000
0!
0*
09
0>
0C
#833510000000
1!
1*
b101 6
19
1>
1C
b101 G
#833520000000
0!
0*
09
0>
0C
#833530000000
1!
1*
b110 6
19
1>
1C
b110 G
#833540000000
0!
0*
09
0>
0C
#833550000000
1!
1*
b111 6
19
1>
1C
b111 G
#833560000000
0!
0*
09
0>
0C
#833570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#833580000000
0!
0*
09
0>
0C
#833590000000
1!
1*
b1 6
19
1>
1C
b1 G
#833600000000
0!
0*
09
0>
0C
#833610000000
1!
1*
b10 6
19
1>
1C
b10 G
#833620000000
0!
0*
09
0>
0C
#833630000000
1!
1*
b11 6
19
1>
1C
b11 G
#833640000000
0!
0*
09
0>
0C
#833650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#833660000000
0!
0*
09
0>
0C
#833670000000
1!
1*
b101 6
19
1>
1C
b101 G
#833680000000
0!
0*
09
0>
0C
#833690000000
1!
1*
b110 6
19
1>
1C
b110 G
#833700000000
0!
0*
09
0>
0C
#833710000000
1!
1*
b111 6
19
1>
1C
b111 G
#833720000000
0!
1"
0*
1+
09
1:
0>
0C
#833730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#833740000000
0!
0*
09
0>
0C
#833750000000
1!
1*
b1 6
19
1>
1C
b1 G
#833760000000
0!
0*
09
0>
0C
#833770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#833780000000
0!
0*
09
0>
0C
#833790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#833800000000
0!
0*
09
0>
0C
#833810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#833820000000
0!
0*
09
0>
0C
#833830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#833840000000
0!
0#
0*
0,
09
0>
0?
0C
#833850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#833860000000
0!
0*
09
0>
0C
#833870000000
1!
1*
19
1>
1C
#833880000000
0!
0*
09
0>
0C
#833890000000
1!
1*
19
1>
1C
#833900000000
0!
0*
09
0>
0C
#833910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#833920000000
0!
0*
09
0>
0C
#833930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#833940000000
0!
0*
09
0>
0C
#833950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#833960000000
0!
0*
09
0>
0C
#833970000000
1!
1*
b10 6
19
1>
1C
b10 G
#833980000000
0!
0*
09
0>
0C
#833990000000
1!
1*
b11 6
19
1>
1C
b11 G
#834000000000
0!
0*
09
0>
0C
#834010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#834020000000
0!
0*
09
0>
0C
#834030000000
1!
1*
b101 6
19
1>
1C
b101 G
#834040000000
0!
0*
09
0>
0C
#834050000000
1!
1*
b110 6
19
1>
1C
b110 G
#834060000000
0!
0*
09
0>
0C
#834070000000
1!
1*
b111 6
19
1>
1C
b111 G
#834080000000
0!
0*
09
0>
0C
#834090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#834100000000
0!
0*
09
0>
0C
#834110000000
1!
1*
b1 6
19
1>
1C
b1 G
#834120000000
0!
0*
09
0>
0C
#834130000000
1!
1*
b10 6
19
1>
1C
b10 G
#834140000000
0!
0*
09
0>
0C
#834150000000
1!
1*
b11 6
19
1>
1C
b11 G
#834160000000
0!
0*
09
0>
0C
#834170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#834180000000
0!
0*
09
0>
0C
#834190000000
1!
1*
b101 6
19
1>
1C
b101 G
#834200000000
0!
0*
09
0>
0C
#834210000000
1!
1*
b110 6
19
1>
1C
b110 G
#834220000000
0!
0*
09
0>
0C
#834230000000
1!
1*
b111 6
19
1>
1C
b111 G
#834240000000
0!
0*
09
0>
0C
#834250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#834260000000
0!
0*
09
0>
0C
#834270000000
1!
1*
b1 6
19
1>
1C
b1 G
#834280000000
0!
0*
09
0>
0C
#834290000000
1!
1*
b10 6
19
1>
1C
b10 G
#834300000000
0!
0*
09
0>
0C
#834310000000
1!
1*
b11 6
19
1>
1C
b11 G
#834320000000
0!
0*
09
0>
0C
#834330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#834340000000
0!
0*
09
0>
0C
#834350000000
1!
1*
b101 6
19
1>
1C
b101 G
#834360000000
0!
0*
09
0>
0C
#834370000000
1!
1*
b110 6
19
1>
1C
b110 G
#834380000000
0!
0*
09
0>
0C
#834390000000
1!
1*
b111 6
19
1>
1C
b111 G
#834400000000
0!
1"
0*
1+
09
1:
0>
0C
#834410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#834420000000
0!
0*
09
0>
0C
#834430000000
1!
1*
b1 6
19
1>
1C
b1 G
#834440000000
0!
0*
09
0>
0C
#834450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#834460000000
0!
0*
09
0>
0C
#834470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#834480000000
0!
0*
09
0>
0C
#834490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#834500000000
0!
0*
09
0>
0C
#834510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#834520000000
0!
0#
0*
0,
09
0>
0?
0C
#834530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#834540000000
0!
0*
09
0>
0C
#834550000000
1!
1*
19
1>
1C
#834560000000
0!
0*
09
0>
0C
#834570000000
1!
1*
19
1>
1C
#834580000000
0!
0*
09
0>
0C
#834590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#834600000000
0!
0*
09
0>
0C
#834610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#834620000000
0!
0*
09
0>
0C
#834630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#834640000000
0!
0*
09
0>
0C
#834650000000
1!
1*
b10 6
19
1>
1C
b10 G
#834660000000
0!
0*
09
0>
0C
#834670000000
1!
1*
b11 6
19
1>
1C
b11 G
#834680000000
0!
0*
09
0>
0C
#834690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#834700000000
0!
0*
09
0>
0C
#834710000000
1!
1*
b101 6
19
1>
1C
b101 G
#834720000000
0!
0*
09
0>
0C
#834730000000
1!
1*
b110 6
19
1>
1C
b110 G
#834740000000
0!
0*
09
0>
0C
#834750000000
1!
1*
b111 6
19
1>
1C
b111 G
#834760000000
0!
0*
09
0>
0C
#834770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#834780000000
0!
0*
09
0>
0C
#834790000000
1!
1*
b1 6
19
1>
1C
b1 G
#834800000000
0!
0*
09
0>
0C
#834810000000
1!
1*
b10 6
19
1>
1C
b10 G
#834820000000
0!
0*
09
0>
0C
#834830000000
1!
1*
b11 6
19
1>
1C
b11 G
#834840000000
0!
0*
09
0>
0C
#834850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#834860000000
0!
0*
09
0>
0C
#834870000000
1!
1*
b101 6
19
1>
1C
b101 G
#834880000000
0!
0*
09
0>
0C
#834890000000
1!
1*
b110 6
19
1>
1C
b110 G
#834900000000
0!
0*
09
0>
0C
#834910000000
1!
1*
b111 6
19
1>
1C
b111 G
#834920000000
0!
0*
09
0>
0C
#834930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#834940000000
0!
0*
09
0>
0C
#834950000000
1!
1*
b1 6
19
1>
1C
b1 G
#834960000000
0!
0*
09
0>
0C
#834970000000
1!
1*
b10 6
19
1>
1C
b10 G
#834980000000
0!
0*
09
0>
0C
#834990000000
1!
1*
b11 6
19
1>
1C
b11 G
#835000000000
0!
0*
09
0>
0C
#835010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#835020000000
0!
0*
09
0>
0C
#835030000000
1!
1*
b101 6
19
1>
1C
b101 G
#835040000000
0!
0*
09
0>
0C
#835050000000
1!
1*
b110 6
19
1>
1C
b110 G
#835060000000
0!
0*
09
0>
0C
#835070000000
1!
1*
b111 6
19
1>
1C
b111 G
#835080000000
0!
1"
0*
1+
09
1:
0>
0C
#835090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#835100000000
0!
0*
09
0>
0C
#835110000000
1!
1*
b1 6
19
1>
1C
b1 G
#835120000000
0!
0*
09
0>
0C
#835130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#835140000000
0!
0*
09
0>
0C
#835150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#835160000000
0!
0*
09
0>
0C
#835170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#835180000000
0!
0*
09
0>
0C
#835190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#835200000000
0!
0#
0*
0,
09
0>
0?
0C
#835210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#835220000000
0!
0*
09
0>
0C
#835230000000
1!
1*
19
1>
1C
#835240000000
0!
0*
09
0>
0C
#835250000000
1!
1*
19
1>
1C
#835260000000
0!
0*
09
0>
0C
#835270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#835280000000
0!
0*
09
0>
0C
#835290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#835300000000
0!
0*
09
0>
0C
#835310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#835320000000
0!
0*
09
0>
0C
#835330000000
1!
1*
b10 6
19
1>
1C
b10 G
#835340000000
0!
0*
09
0>
0C
#835350000000
1!
1*
b11 6
19
1>
1C
b11 G
#835360000000
0!
0*
09
0>
0C
#835370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#835380000000
0!
0*
09
0>
0C
#835390000000
1!
1*
b101 6
19
1>
1C
b101 G
#835400000000
0!
0*
09
0>
0C
#835410000000
1!
1*
b110 6
19
1>
1C
b110 G
#835420000000
0!
0*
09
0>
0C
#835430000000
1!
1*
b111 6
19
1>
1C
b111 G
#835440000000
0!
0*
09
0>
0C
#835450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#835460000000
0!
0*
09
0>
0C
#835470000000
1!
1*
b1 6
19
1>
1C
b1 G
#835480000000
0!
0*
09
0>
0C
#835490000000
1!
1*
b10 6
19
1>
1C
b10 G
#835500000000
0!
0*
09
0>
0C
#835510000000
1!
1*
b11 6
19
1>
1C
b11 G
#835520000000
0!
0*
09
0>
0C
#835530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#835540000000
0!
0*
09
0>
0C
#835550000000
1!
1*
b101 6
19
1>
1C
b101 G
#835560000000
0!
0*
09
0>
0C
#835570000000
1!
1*
b110 6
19
1>
1C
b110 G
#835580000000
0!
0*
09
0>
0C
#835590000000
1!
1*
b111 6
19
1>
1C
b111 G
#835600000000
0!
0*
09
0>
0C
#835610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#835620000000
0!
0*
09
0>
0C
#835630000000
1!
1*
b1 6
19
1>
1C
b1 G
#835640000000
0!
0*
09
0>
0C
#835650000000
1!
1*
b10 6
19
1>
1C
b10 G
#835660000000
0!
0*
09
0>
0C
#835670000000
1!
1*
b11 6
19
1>
1C
b11 G
#835680000000
0!
0*
09
0>
0C
#835690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#835700000000
0!
0*
09
0>
0C
#835710000000
1!
1*
b101 6
19
1>
1C
b101 G
#835720000000
0!
0*
09
0>
0C
#835730000000
1!
1*
b110 6
19
1>
1C
b110 G
#835740000000
0!
0*
09
0>
0C
#835750000000
1!
1*
b111 6
19
1>
1C
b111 G
#835760000000
0!
1"
0*
1+
09
1:
0>
0C
#835770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#835780000000
0!
0*
09
0>
0C
#835790000000
1!
1*
b1 6
19
1>
1C
b1 G
#835800000000
0!
0*
09
0>
0C
#835810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#835820000000
0!
0*
09
0>
0C
#835830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#835840000000
0!
0*
09
0>
0C
#835850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#835860000000
0!
0*
09
0>
0C
#835870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#835880000000
0!
0#
0*
0,
09
0>
0?
0C
#835890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#835900000000
0!
0*
09
0>
0C
#835910000000
1!
1*
19
1>
1C
#835920000000
0!
0*
09
0>
0C
#835930000000
1!
1*
19
1>
1C
#835940000000
0!
0*
09
0>
0C
#835950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#835960000000
0!
0*
09
0>
0C
#835970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#835980000000
0!
0*
09
0>
0C
#835990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#836000000000
0!
0*
09
0>
0C
#836010000000
1!
1*
b10 6
19
1>
1C
b10 G
#836020000000
0!
0*
09
0>
0C
#836030000000
1!
1*
b11 6
19
1>
1C
b11 G
#836040000000
0!
0*
09
0>
0C
#836050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#836060000000
0!
0*
09
0>
0C
#836070000000
1!
1*
b101 6
19
1>
1C
b101 G
#836080000000
0!
0*
09
0>
0C
#836090000000
1!
1*
b110 6
19
1>
1C
b110 G
#836100000000
0!
0*
09
0>
0C
#836110000000
1!
1*
b111 6
19
1>
1C
b111 G
#836120000000
0!
0*
09
0>
0C
#836130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#836140000000
0!
0*
09
0>
0C
#836150000000
1!
1*
b1 6
19
1>
1C
b1 G
#836160000000
0!
0*
09
0>
0C
#836170000000
1!
1*
b10 6
19
1>
1C
b10 G
#836180000000
0!
0*
09
0>
0C
#836190000000
1!
1*
b11 6
19
1>
1C
b11 G
#836200000000
0!
0*
09
0>
0C
#836210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#836220000000
0!
0*
09
0>
0C
#836230000000
1!
1*
b101 6
19
1>
1C
b101 G
#836240000000
0!
0*
09
0>
0C
#836250000000
1!
1*
b110 6
19
1>
1C
b110 G
#836260000000
0!
0*
09
0>
0C
#836270000000
1!
1*
b111 6
19
1>
1C
b111 G
#836280000000
0!
0*
09
0>
0C
#836290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#836300000000
0!
0*
09
0>
0C
#836310000000
1!
1*
b1 6
19
1>
1C
b1 G
#836320000000
0!
0*
09
0>
0C
#836330000000
1!
1*
b10 6
19
1>
1C
b10 G
#836340000000
0!
0*
09
0>
0C
#836350000000
1!
1*
b11 6
19
1>
1C
b11 G
#836360000000
0!
0*
09
0>
0C
#836370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#836380000000
0!
0*
09
0>
0C
#836390000000
1!
1*
b101 6
19
1>
1C
b101 G
#836400000000
0!
0*
09
0>
0C
#836410000000
1!
1*
b110 6
19
1>
1C
b110 G
#836420000000
0!
0*
09
0>
0C
#836430000000
1!
1*
b111 6
19
1>
1C
b111 G
#836440000000
0!
1"
0*
1+
09
1:
0>
0C
#836450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#836460000000
0!
0*
09
0>
0C
#836470000000
1!
1*
b1 6
19
1>
1C
b1 G
#836480000000
0!
0*
09
0>
0C
#836490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#836500000000
0!
0*
09
0>
0C
#836510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#836520000000
0!
0*
09
0>
0C
#836530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#836540000000
0!
0*
09
0>
0C
#836550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#836560000000
0!
0#
0*
0,
09
0>
0?
0C
#836570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#836580000000
0!
0*
09
0>
0C
#836590000000
1!
1*
19
1>
1C
#836600000000
0!
0*
09
0>
0C
#836610000000
1!
1*
19
1>
1C
#836620000000
0!
0*
09
0>
0C
#836630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#836640000000
0!
0*
09
0>
0C
#836650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#836660000000
0!
0*
09
0>
0C
#836670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#836680000000
0!
0*
09
0>
0C
#836690000000
1!
1*
b10 6
19
1>
1C
b10 G
#836700000000
0!
0*
09
0>
0C
#836710000000
1!
1*
b11 6
19
1>
1C
b11 G
#836720000000
0!
0*
09
0>
0C
#836730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#836740000000
0!
0*
09
0>
0C
#836750000000
1!
1*
b101 6
19
1>
1C
b101 G
#836760000000
0!
0*
09
0>
0C
#836770000000
1!
1*
b110 6
19
1>
1C
b110 G
#836780000000
0!
0*
09
0>
0C
#836790000000
1!
1*
b111 6
19
1>
1C
b111 G
#836800000000
0!
0*
09
0>
0C
#836810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#836820000000
0!
0*
09
0>
0C
#836830000000
1!
1*
b1 6
19
1>
1C
b1 G
#836840000000
0!
0*
09
0>
0C
#836850000000
1!
1*
b10 6
19
1>
1C
b10 G
#836860000000
0!
0*
09
0>
0C
#836870000000
1!
1*
b11 6
19
1>
1C
b11 G
#836880000000
0!
0*
09
0>
0C
#836890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#836900000000
0!
0*
09
0>
0C
#836910000000
1!
1*
b101 6
19
1>
1C
b101 G
#836920000000
0!
0*
09
0>
0C
#836930000000
1!
1*
b110 6
19
1>
1C
b110 G
#836940000000
0!
0*
09
0>
0C
#836950000000
1!
1*
b111 6
19
1>
1C
b111 G
#836960000000
0!
0*
09
0>
0C
#836970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#836980000000
0!
0*
09
0>
0C
#836990000000
1!
1*
b1 6
19
1>
1C
b1 G
#837000000000
0!
0*
09
0>
0C
#837010000000
1!
1*
b10 6
19
1>
1C
b10 G
#837020000000
0!
0*
09
0>
0C
#837030000000
1!
1*
b11 6
19
1>
1C
b11 G
#837040000000
0!
0*
09
0>
0C
#837050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#837060000000
0!
0*
09
0>
0C
#837070000000
1!
1*
b101 6
19
1>
1C
b101 G
#837080000000
0!
0*
09
0>
0C
#837090000000
1!
1*
b110 6
19
1>
1C
b110 G
#837100000000
0!
0*
09
0>
0C
#837110000000
1!
1*
b111 6
19
1>
1C
b111 G
#837120000000
0!
1"
0*
1+
09
1:
0>
0C
#837130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#837140000000
0!
0*
09
0>
0C
#837150000000
1!
1*
b1 6
19
1>
1C
b1 G
#837160000000
0!
0*
09
0>
0C
#837170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#837180000000
0!
0*
09
0>
0C
#837190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#837200000000
0!
0*
09
0>
0C
#837210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#837220000000
0!
0*
09
0>
0C
#837230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#837240000000
0!
0#
0*
0,
09
0>
0?
0C
#837250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#837260000000
0!
0*
09
0>
0C
#837270000000
1!
1*
19
1>
1C
#837280000000
0!
0*
09
0>
0C
#837290000000
1!
1*
19
1>
1C
#837300000000
0!
0*
09
0>
0C
#837310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#837320000000
0!
0*
09
0>
0C
#837330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#837340000000
0!
0*
09
0>
0C
#837350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#837360000000
0!
0*
09
0>
0C
#837370000000
1!
1*
b10 6
19
1>
1C
b10 G
#837380000000
0!
0*
09
0>
0C
#837390000000
1!
1*
b11 6
19
1>
1C
b11 G
#837400000000
0!
0*
09
0>
0C
#837410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#837420000000
0!
0*
09
0>
0C
#837430000000
1!
1*
b101 6
19
1>
1C
b101 G
#837440000000
0!
0*
09
0>
0C
#837450000000
1!
1*
b110 6
19
1>
1C
b110 G
#837460000000
0!
0*
09
0>
0C
#837470000000
1!
1*
b111 6
19
1>
1C
b111 G
#837480000000
0!
0*
09
0>
0C
#837490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#837500000000
0!
0*
09
0>
0C
#837510000000
1!
1*
b1 6
19
1>
1C
b1 G
#837520000000
0!
0*
09
0>
0C
#837530000000
1!
1*
b10 6
19
1>
1C
b10 G
#837540000000
0!
0*
09
0>
0C
#837550000000
1!
1*
b11 6
19
1>
1C
b11 G
#837560000000
0!
0*
09
0>
0C
#837570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#837580000000
0!
0*
09
0>
0C
#837590000000
1!
1*
b101 6
19
1>
1C
b101 G
#837600000000
0!
0*
09
0>
0C
#837610000000
1!
1*
b110 6
19
1>
1C
b110 G
#837620000000
0!
0*
09
0>
0C
#837630000000
1!
1*
b111 6
19
1>
1C
b111 G
#837640000000
0!
0*
09
0>
0C
#837650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#837660000000
0!
0*
09
0>
0C
#837670000000
1!
1*
b1 6
19
1>
1C
b1 G
#837680000000
0!
0*
09
0>
0C
#837690000000
1!
1*
b10 6
19
1>
1C
b10 G
#837700000000
0!
0*
09
0>
0C
#837710000000
1!
1*
b11 6
19
1>
1C
b11 G
#837720000000
0!
0*
09
0>
0C
#837730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#837740000000
0!
0*
09
0>
0C
#837750000000
1!
1*
b101 6
19
1>
1C
b101 G
#837760000000
0!
0*
09
0>
0C
#837770000000
1!
1*
b110 6
19
1>
1C
b110 G
#837780000000
0!
0*
09
0>
0C
#837790000000
1!
1*
b111 6
19
1>
1C
b111 G
#837800000000
0!
1"
0*
1+
09
1:
0>
0C
#837810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#837820000000
0!
0*
09
0>
0C
#837830000000
1!
1*
b1 6
19
1>
1C
b1 G
#837840000000
0!
0*
09
0>
0C
#837850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#837860000000
0!
0*
09
0>
0C
#837870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#837880000000
0!
0*
09
0>
0C
#837890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#837900000000
0!
0*
09
0>
0C
#837910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#837920000000
0!
0#
0*
0,
09
0>
0?
0C
#837930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#837940000000
0!
0*
09
0>
0C
#837950000000
1!
1*
19
1>
1C
#837960000000
0!
0*
09
0>
0C
#837970000000
1!
1*
19
1>
1C
#837980000000
0!
0*
09
0>
0C
#837990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#838000000000
0!
0*
09
0>
0C
#838010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#838020000000
0!
0*
09
0>
0C
#838030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#838040000000
0!
0*
09
0>
0C
#838050000000
1!
1*
b10 6
19
1>
1C
b10 G
#838060000000
0!
0*
09
0>
0C
#838070000000
1!
1*
b11 6
19
1>
1C
b11 G
#838080000000
0!
0*
09
0>
0C
#838090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#838100000000
0!
0*
09
0>
0C
#838110000000
1!
1*
b101 6
19
1>
1C
b101 G
#838120000000
0!
0*
09
0>
0C
#838130000000
1!
1*
b110 6
19
1>
1C
b110 G
#838140000000
0!
0*
09
0>
0C
#838150000000
1!
1*
b111 6
19
1>
1C
b111 G
#838160000000
0!
0*
09
0>
0C
#838170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#838180000000
0!
0*
09
0>
0C
#838190000000
1!
1*
b1 6
19
1>
1C
b1 G
#838200000000
0!
0*
09
0>
0C
#838210000000
1!
1*
b10 6
19
1>
1C
b10 G
#838220000000
0!
0*
09
0>
0C
#838230000000
1!
1*
b11 6
19
1>
1C
b11 G
#838240000000
0!
0*
09
0>
0C
#838250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#838260000000
0!
0*
09
0>
0C
#838270000000
1!
1*
b101 6
19
1>
1C
b101 G
#838280000000
0!
0*
09
0>
0C
#838290000000
1!
1*
b110 6
19
1>
1C
b110 G
#838300000000
0!
0*
09
0>
0C
#838310000000
1!
1*
b111 6
19
1>
1C
b111 G
#838320000000
0!
0*
09
0>
0C
#838330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#838340000000
0!
0*
09
0>
0C
#838350000000
1!
1*
b1 6
19
1>
1C
b1 G
#838360000000
0!
0*
09
0>
0C
#838370000000
1!
1*
b10 6
19
1>
1C
b10 G
#838380000000
0!
0*
09
0>
0C
#838390000000
1!
1*
b11 6
19
1>
1C
b11 G
#838400000000
0!
0*
09
0>
0C
#838410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#838420000000
0!
0*
09
0>
0C
#838430000000
1!
1*
b101 6
19
1>
1C
b101 G
#838440000000
0!
0*
09
0>
0C
#838450000000
1!
1*
b110 6
19
1>
1C
b110 G
#838460000000
0!
0*
09
0>
0C
#838470000000
1!
1*
b111 6
19
1>
1C
b111 G
#838480000000
0!
1"
0*
1+
09
1:
0>
0C
#838490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#838500000000
0!
0*
09
0>
0C
#838510000000
1!
1*
b1 6
19
1>
1C
b1 G
#838520000000
0!
0*
09
0>
0C
#838530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#838540000000
0!
0*
09
0>
0C
#838550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#838560000000
0!
0*
09
0>
0C
#838570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#838580000000
0!
0*
09
0>
0C
#838590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#838600000000
0!
0#
0*
0,
09
0>
0?
0C
#838610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#838620000000
0!
0*
09
0>
0C
#838630000000
1!
1*
19
1>
1C
#838640000000
0!
0*
09
0>
0C
#838650000000
1!
1*
19
1>
1C
#838660000000
0!
0*
09
0>
0C
#838670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#838680000000
0!
0*
09
0>
0C
#838690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#838700000000
0!
0*
09
0>
0C
#838710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#838720000000
0!
0*
09
0>
0C
#838730000000
1!
1*
b10 6
19
1>
1C
b10 G
#838740000000
0!
0*
09
0>
0C
#838750000000
1!
1*
b11 6
19
1>
1C
b11 G
#838760000000
0!
0*
09
0>
0C
#838770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#838780000000
0!
0*
09
0>
0C
#838790000000
1!
1*
b101 6
19
1>
1C
b101 G
#838800000000
0!
0*
09
0>
0C
#838810000000
1!
1*
b110 6
19
1>
1C
b110 G
#838820000000
0!
0*
09
0>
0C
#838830000000
1!
1*
b111 6
19
1>
1C
b111 G
#838840000000
0!
0*
09
0>
0C
#838850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#838860000000
0!
0*
09
0>
0C
#838870000000
1!
1*
b1 6
19
1>
1C
b1 G
#838880000000
0!
0*
09
0>
0C
#838890000000
1!
1*
b10 6
19
1>
1C
b10 G
#838900000000
0!
0*
09
0>
0C
#838910000000
1!
1*
b11 6
19
1>
1C
b11 G
#838920000000
0!
0*
09
0>
0C
#838930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#838940000000
0!
0*
09
0>
0C
#838950000000
1!
1*
b101 6
19
1>
1C
b101 G
#838960000000
0!
0*
09
0>
0C
#838970000000
1!
1*
b110 6
19
1>
1C
b110 G
#838980000000
0!
0*
09
0>
0C
#838990000000
1!
1*
b111 6
19
1>
1C
b111 G
#839000000000
0!
0*
09
0>
0C
#839010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#839020000000
0!
0*
09
0>
0C
#839030000000
1!
1*
b1 6
19
1>
1C
b1 G
#839040000000
0!
0*
09
0>
0C
#839050000000
1!
1*
b10 6
19
1>
1C
b10 G
#839060000000
0!
0*
09
0>
0C
#839070000000
1!
1*
b11 6
19
1>
1C
b11 G
#839080000000
0!
0*
09
0>
0C
#839090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#839100000000
0!
0*
09
0>
0C
#839110000000
1!
1*
b101 6
19
1>
1C
b101 G
#839120000000
0!
0*
09
0>
0C
#839130000000
1!
1*
b110 6
19
1>
1C
b110 G
#839140000000
0!
0*
09
0>
0C
#839150000000
1!
1*
b111 6
19
1>
1C
b111 G
#839160000000
0!
1"
0*
1+
09
1:
0>
0C
#839170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#839180000000
0!
0*
09
0>
0C
#839190000000
1!
1*
b1 6
19
1>
1C
b1 G
#839200000000
0!
0*
09
0>
0C
#839210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#839220000000
0!
0*
09
0>
0C
#839230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#839240000000
0!
0*
09
0>
0C
#839250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#839260000000
0!
0*
09
0>
0C
#839270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#839280000000
0!
0#
0*
0,
09
0>
0?
0C
#839290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#839300000000
0!
0*
09
0>
0C
#839310000000
1!
1*
19
1>
1C
#839320000000
0!
0*
09
0>
0C
#839330000000
1!
1*
19
1>
1C
#839340000000
0!
0*
09
0>
0C
#839350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#839360000000
0!
0*
09
0>
0C
#839370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#839380000000
0!
0*
09
0>
0C
#839390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#839400000000
0!
0*
09
0>
0C
#839410000000
1!
1*
b10 6
19
1>
1C
b10 G
#839420000000
0!
0*
09
0>
0C
#839430000000
1!
1*
b11 6
19
1>
1C
b11 G
#839440000000
0!
0*
09
0>
0C
#839450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#839460000000
0!
0*
09
0>
0C
#839470000000
1!
1*
b101 6
19
1>
1C
b101 G
#839480000000
0!
0*
09
0>
0C
#839490000000
1!
1*
b110 6
19
1>
1C
b110 G
#839500000000
0!
0*
09
0>
0C
#839510000000
1!
1*
b111 6
19
1>
1C
b111 G
#839520000000
0!
0*
09
0>
0C
#839530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#839540000000
0!
0*
09
0>
0C
#839550000000
1!
1*
b1 6
19
1>
1C
b1 G
#839560000000
0!
0*
09
0>
0C
#839570000000
1!
1*
b10 6
19
1>
1C
b10 G
#839580000000
0!
0*
09
0>
0C
#839590000000
1!
1*
b11 6
19
1>
1C
b11 G
#839600000000
0!
0*
09
0>
0C
#839610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#839620000000
0!
0*
09
0>
0C
#839630000000
1!
1*
b101 6
19
1>
1C
b101 G
#839640000000
0!
0*
09
0>
0C
#839650000000
1!
1*
b110 6
19
1>
1C
b110 G
#839660000000
0!
0*
09
0>
0C
#839670000000
1!
1*
b111 6
19
1>
1C
b111 G
#839680000000
0!
0*
09
0>
0C
#839690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#839700000000
0!
0*
09
0>
0C
#839710000000
1!
1*
b1 6
19
1>
1C
b1 G
#839720000000
0!
0*
09
0>
0C
#839730000000
1!
1*
b10 6
19
1>
1C
b10 G
#839740000000
0!
0*
09
0>
0C
#839750000000
1!
1*
b11 6
19
1>
1C
b11 G
#839760000000
0!
0*
09
0>
0C
#839770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#839780000000
0!
0*
09
0>
0C
#839790000000
1!
1*
b101 6
19
1>
1C
b101 G
#839800000000
0!
0*
09
0>
0C
#839810000000
1!
1*
b110 6
19
1>
1C
b110 G
#839820000000
0!
0*
09
0>
0C
#839830000000
1!
1*
b111 6
19
1>
1C
b111 G
#839840000000
0!
1"
0*
1+
09
1:
0>
0C
#839850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#839860000000
0!
0*
09
0>
0C
#839870000000
1!
1*
b1 6
19
1>
1C
b1 G
#839880000000
0!
0*
09
0>
0C
#839890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#839900000000
0!
0*
09
0>
0C
#839910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#839920000000
0!
0*
09
0>
0C
#839930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#839940000000
0!
0*
09
0>
0C
#839950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#839960000000
0!
0#
0*
0,
09
0>
0?
0C
#839970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#839980000000
0!
0*
09
0>
0C
#839990000000
1!
1*
19
1>
1C
#840000000000
0!
0*
09
0>
0C
#840010000000
1!
1*
19
1>
1C
#840020000000
0!
0*
09
0>
0C
#840030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#840040000000
0!
0*
09
0>
0C
#840050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#840060000000
0!
0*
09
0>
0C
#840070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#840080000000
0!
0*
09
0>
0C
#840090000000
1!
1*
b10 6
19
1>
1C
b10 G
#840100000000
0!
0*
09
0>
0C
#840110000000
1!
1*
b11 6
19
1>
1C
b11 G
#840120000000
0!
0*
09
0>
0C
#840130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#840140000000
0!
0*
09
0>
0C
#840150000000
1!
1*
b101 6
19
1>
1C
b101 G
#840160000000
0!
0*
09
0>
0C
#840170000000
1!
1*
b110 6
19
1>
1C
b110 G
#840180000000
0!
0*
09
0>
0C
#840190000000
1!
1*
b111 6
19
1>
1C
b111 G
#840200000000
0!
0*
09
0>
0C
#840210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#840220000000
0!
0*
09
0>
0C
#840230000000
1!
1*
b1 6
19
1>
1C
b1 G
#840240000000
0!
0*
09
0>
0C
#840250000000
1!
1*
b10 6
19
1>
1C
b10 G
#840260000000
0!
0*
09
0>
0C
#840270000000
1!
1*
b11 6
19
1>
1C
b11 G
#840280000000
0!
0*
09
0>
0C
#840290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#840300000000
0!
0*
09
0>
0C
#840310000000
1!
1*
b101 6
19
1>
1C
b101 G
#840320000000
0!
0*
09
0>
0C
#840330000000
1!
1*
b110 6
19
1>
1C
b110 G
#840340000000
0!
0*
09
0>
0C
#840350000000
1!
1*
b111 6
19
1>
1C
b111 G
#840360000000
0!
0*
09
0>
0C
#840370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#840380000000
0!
0*
09
0>
0C
#840390000000
1!
1*
b1 6
19
1>
1C
b1 G
#840400000000
0!
0*
09
0>
0C
#840410000000
1!
1*
b10 6
19
1>
1C
b10 G
#840420000000
0!
0*
09
0>
0C
#840430000000
1!
1*
b11 6
19
1>
1C
b11 G
#840440000000
0!
0*
09
0>
0C
#840450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#840460000000
0!
0*
09
0>
0C
#840470000000
1!
1*
b101 6
19
1>
1C
b101 G
#840480000000
0!
0*
09
0>
0C
#840490000000
1!
1*
b110 6
19
1>
1C
b110 G
#840500000000
0!
0*
09
0>
0C
#840510000000
1!
1*
b111 6
19
1>
1C
b111 G
#840520000000
0!
1"
0*
1+
09
1:
0>
0C
#840530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#840540000000
0!
0*
09
0>
0C
#840550000000
1!
1*
b1 6
19
1>
1C
b1 G
#840560000000
0!
0*
09
0>
0C
#840570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#840580000000
0!
0*
09
0>
0C
#840590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#840600000000
0!
0*
09
0>
0C
#840610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#840620000000
0!
0*
09
0>
0C
#840630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#840640000000
0!
0#
0*
0,
09
0>
0?
0C
#840650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#840660000000
0!
0*
09
0>
0C
#840670000000
1!
1*
19
1>
1C
#840680000000
0!
0*
09
0>
0C
#840690000000
1!
1*
19
1>
1C
#840700000000
0!
0*
09
0>
0C
#840710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#840720000000
0!
0*
09
0>
0C
#840730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#840740000000
0!
0*
09
0>
0C
#840750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#840760000000
0!
0*
09
0>
0C
#840770000000
1!
1*
b10 6
19
1>
1C
b10 G
#840780000000
0!
0*
09
0>
0C
#840790000000
1!
1*
b11 6
19
1>
1C
b11 G
#840800000000
0!
0*
09
0>
0C
#840810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#840820000000
0!
0*
09
0>
0C
#840830000000
1!
1*
b101 6
19
1>
1C
b101 G
#840840000000
0!
0*
09
0>
0C
#840850000000
1!
1*
b110 6
19
1>
1C
b110 G
#840860000000
0!
0*
09
0>
0C
#840870000000
1!
1*
b111 6
19
1>
1C
b111 G
#840880000000
0!
0*
09
0>
0C
#840890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#840900000000
0!
0*
09
0>
0C
#840910000000
1!
1*
b1 6
19
1>
1C
b1 G
#840920000000
0!
0*
09
0>
0C
#840930000000
1!
1*
b10 6
19
1>
1C
b10 G
#840940000000
0!
0*
09
0>
0C
#840950000000
1!
1*
b11 6
19
1>
1C
b11 G
#840960000000
0!
0*
09
0>
0C
#840970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#840980000000
0!
0*
09
0>
0C
#840990000000
1!
1*
b101 6
19
1>
1C
b101 G
#841000000000
0!
0*
09
0>
0C
#841010000000
1!
1*
b110 6
19
1>
1C
b110 G
#841020000000
0!
0*
09
0>
0C
#841030000000
1!
1*
b111 6
19
1>
1C
b111 G
#841040000000
0!
0*
09
0>
0C
#841050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#841060000000
0!
0*
09
0>
0C
#841070000000
1!
1*
b1 6
19
1>
1C
b1 G
#841080000000
0!
0*
09
0>
0C
#841090000000
1!
1*
b10 6
19
1>
1C
b10 G
#841100000000
0!
0*
09
0>
0C
#841110000000
1!
1*
b11 6
19
1>
1C
b11 G
#841120000000
0!
0*
09
0>
0C
#841130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#841140000000
0!
0*
09
0>
0C
#841150000000
1!
1*
b101 6
19
1>
1C
b101 G
#841160000000
0!
0*
09
0>
0C
#841170000000
1!
1*
b110 6
19
1>
1C
b110 G
#841180000000
0!
0*
09
0>
0C
#841190000000
1!
1*
b111 6
19
1>
1C
b111 G
#841200000000
0!
1"
0*
1+
09
1:
0>
0C
#841210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#841220000000
0!
0*
09
0>
0C
#841230000000
1!
1*
b1 6
19
1>
1C
b1 G
#841240000000
0!
0*
09
0>
0C
#841250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#841260000000
0!
0*
09
0>
0C
#841270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#841280000000
0!
0*
09
0>
0C
#841290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#841300000000
0!
0*
09
0>
0C
#841310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#841320000000
0!
0#
0*
0,
09
0>
0?
0C
#841330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#841340000000
0!
0*
09
0>
0C
#841350000000
1!
1*
19
1>
1C
#841360000000
0!
0*
09
0>
0C
#841370000000
1!
1*
19
1>
1C
#841380000000
0!
0*
09
0>
0C
#841390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#841400000000
0!
0*
09
0>
0C
#841410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#841420000000
0!
0*
09
0>
0C
#841430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#841440000000
0!
0*
09
0>
0C
#841450000000
1!
1*
b10 6
19
1>
1C
b10 G
#841460000000
0!
0*
09
0>
0C
#841470000000
1!
1*
b11 6
19
1>
1C
b11 G
#841480000000
0!
0*
09
0>
0C
#841490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#841500000000
0!
0*
09
0>
0C
#841510000000
1!
1*
b101 6
19
1>
1C
b101 G
#841520000000
0!
0*
09
0>
0C
#841530000000
1!
1*
b110 6
19
1>
1C
b110 G
#841540000000
0!
0*
09
0>
0C
#841550000000
1!
1*
b111 6
19
1>
1C
b111 G
#841560000000
0!
0*
09
0>
0C
#841570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#841580000000
0!
0*
09
0>
0C
#841590000000
1!
1*
b1 6
19
1>
1C
b1 G
#841600000000
0!
0*
09
0>
0C
#841610000000
1!
1*
b10 6
19
1>
1C
b10 G
#841620000000
0!
0*
09
0>
0C
#841630000000
1!
1*
b11 6
19
1>
1C
b11 G
#841640000000
0!
0*
09
0>
0C
#841650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#841660000000
0!
0*
09
0>
0C
#841670000000
1!
1*
b101 6
19
1>
1C
b101 G
#841680000000
0!
0*
09
0>
0C
#841690000000
1!
1*
b110 6
19
1>
1C
b110 G
#841700000000
0!
0*
09
0>
0C
#841710000000
1!
1*
b111 6
19
1>
1C
b111 G
#841720000000
0!
0*
09
0>
0C
#841730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#841740000000
0!
0*
09
0>
0C
#841750000000
1!
1*
b1 6
19
1>
1C
b1 G
#841760000000
0!
0*
09
0>
0C
#841770000000
1!
1*
b10 6
19
1>
1C
b10 G
#841780000000
0!
0*
09
0>
0C
#841790000000
1!
1*
b11 6
19
1>
1C
b11 G
#841800000000
0!
0*
09
0>
0C
#841810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#841820000000
0!
0*
09
0>
0C
#841830000000
1!
1*
b101 6
19
1>
1C
b101 G
#841840000000
0!
0*
09
0>
0C
#841850000000
1!
1*
b110 6
19
1>
1C
b110 G
#841860000000
0!
0*
09
0>
0C
#841870000000
1!
1*
b111 6
19
1>
1C
b111 G
#841880000000
0!
1"
0*
1+
09
1:
0>
0C
#841890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#841900000000
0!
0*
09
0>
0C
#841910000000
1!
1*
b1 6
19
1>
1C
b1 G
#841920000000
0!
0*
09
0>
0C
#841930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#841940000000
0!
0*
09
0>
0C
#841950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#841960000000
0!
0*
09
0>
0C
#841970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#841980000000
0!
0*
09
0>
0C
#841990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#842000000000
0!
0#
0*
0,
09
0>
0?
0C
#842010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#842020000000
0!
0*
09
0>
0C
#842030000000
1!
1*
19
1>
1C
#842040000000
0!
0*
09
0>
0C
#842050000000
1!
1*
19
1>
1C
#842060000000
0!
0*
09
0>
0C
#842070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#842080000000
0!
0*
09
0>
0C
#842090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#842100000000
0!
0*
09
0>
0C
#842110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#842120000000
0!
0*
09
0>
0C
#842130000000
1!
1*
b10 6
19
1>
1C
b10 G
#842140000000
0!
0*
09
0>
0C
#842150000000
1!
1*
b11 6
19
1>
1C
b11 G
#842160000000
0!
0*
09
0>
0C
#842170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#842180000000
0!
0*
09
0>
0C
#842190000000
1!
1*
b101 6
19
1>
1C
b101 G
#842200000000
0!
0*
09
0>
0C
#842210000000
1!
1*
b110 6
19
1>
1C
b110 G
#842220000000
0!
0*
09
0>
0C
#842230000000
1!
1*
b111 6
19
1>
1C
b111 G
#842240000000
0!
0*
09
0>
0C
#842250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#842260000000
0!
0*
09
0>
0C
#842270000000
1!
1*
b1 6
19
1>
1C
b1 G
#842280000000
0!
0*
09
0>
0C
#842290000000
1!
1*
b10 6
19
1>
1C
b10 G
#842300000000
0!
0*
09
0>
0C
#842310000000
1!
1*
b11 6
19
1>
1C
b11 G
#842320000000
0!
0*
09
0>
0C
#842330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#842340000000
0!
0*
09
0>
0C
#842350000000
1!
1*
b101 6
19
1>
1C
b101 G
#842360000000
0!
0*
09
0>
0C
#842370000000
1!
1*
b110 6
19
1>
1C
b110 G
#842380000000
0!
0*
09
0>
0C
#842390000000
1!
1*
b111 6
19
1>
1C
b111 G
#842400000000
0!
0*
09
0>
0C
#842410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#842420000000
0!
0*
09
0>
0C
#842430000000
1!
1*
b1 6
19
1>
1C
b1 G
#842440000000
0!
0*
09
0>
0C
#842450000000
1!
1*
b10 6
19
1>
1C
b10 G
#842460000000
0!
0*
09
0>
0C
#842470000000
1!
1*
b11 6
19
1>
1C
b11 G
#842480000000
0!
0*
09
0>
0C
#842490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#842500000000
0!
0*
09
0>
0C
#842510000000
1!
1*
b101 6
19
1>
1C
b101 G
#842520000000
0!
0*
09
0>
0C
#842530000000
1!
1*
b110 6
19
1>
1C
b110 G
#842540000000
0!
0*
09
0>
0C
#842550000000
1!
1*
b111 6
19
1>
1C
b111 G
#842560000000
0!
1"
0*
1+
09
1:
0>
0C
#842570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#842580000000
0!
0*
09
0>
0C
#842590000000
1!
1*
b1 6
19
1>
1C
b1 G
#842600000000
0!
0*
09
0>
0C
#842610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#842620000000
0!
0*
09
0>
0C
#842630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#842640000000
0!
0*
09
0>
0C
#842650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#842660000000
0!
0*
09
0>
0C
#842670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#842680000000
0!
0#
0*
0,
09
0>
0?
0C
#842690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#842700000000
0!
0*
09
0>
0C
#842710000000
1!
1*
19
1>
1C
#842720000000
0!
0*
09
0>
0C
#842730000000
1!
1*
19
1>
1C
#842740000000
0!
0*
09
0>
0C
#842750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#842760000000
0!
0*
09
0>
0C
#842770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#842780000000
0!
0*
09
0>
0C
#842790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#842800000000
0!
0*
09
0>
0C
#842810000000
1!
1*
b10 6
19
1>
1C
b10 G
#842820000000
0!
0*
09
0>
0C
#842830000000
1!
1*
b11 6
19
1>
1C
b11 G
#842840000000
0!
0*
09
0>
0C
#842850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#842860000000
0!
0*
09
0>
0C
#842870000000
1!
1*
b101 6
19
1>
1C
b101 G
#842880000000
0!
0*
09
0>
0C
#842890000000
1!
1*
b110 6
19
1>
1C
b110 G
#842900000000
0!
0*
09
0>
0C
#842910000000
1!
1*
b111 6
19
1>
1C
b111 G
#842920000000
0!
0*
09
0>
0C
#842930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#842940000000
0!
0*
09
0>
0C
#842950000000
1!
1*
b1 6
19
1>
1C
b1 G
#842960000000
0!
0*
09
0>
0C
#842970000000
1!
1*
b10 6
19
1>
1C
b10 G
#842980000000
0!
0*
09
0>
0C
#842990000000
1!
1*
b11 6
19
1>
1C
b11 G
#843000000000
0!
0*
09
0>
0C
#843010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#843020000000
0!
0*
09
0>
0C
#843030000000
1!
1*
b101 6
19
1>
1C
b101 G
#843040000000
0!
0*
09
0>
0C
#843050000000
1!
1*
b110 6
19
1>
1C
b110 G
#843060000000
0!
0*
09
0>
0C
#843070000000
1!
1*
b111 6
19
1>
1C
b111 G
#843080000000
0!
0*
09
0>
0C
#843090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#843100000000
0!
0*
09
0>
0C
#843110000000
1!
1*
b1 6
19
1>
1C
b1 G
#843120000000
0!
0*
09
0>
0C
#843130000000
1!
1*
b10 6
19
1>
1C
b10 G
#843140000000
0!
0*
09
0>
0C
#843150000000
1!
1*
b11 6
19
1>
1C
b11 G
#843160000000
0!
0*
09
0>
0C
#843170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#843180000000
0!
0*
09
0>
0C
#843190000000
1!
1*
b101 6
19
1>
1C
b101 G
#843200000000
0!
0*
09
0>
0C
#843210000000
1!
1*
b110 6
19
1>
1C
b110 G
#843220000000
0!
0*
09
0>
0C
#843230000000
1!
1*
b111 6
19
1>
1C
b111 G
#843240000000
0!
1"
0*
1+
09
1:
0>
0C
#843250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#843260000000
0!
0*
09
0>
0C
#843270000000
1!
1*
b1 6
19
1>
1C
b1 G
#843280000000
0!
0*
09
0>
0C
#843290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#843300000000
0!
0*
09
0>
0C
#843310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#843320000000
0!
0*
09
0>
0C
#843330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#843340000000
0!
0*
09
0>
0C
#843350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#843360000000
0!
0#
0*
0,
09
0>
0?
0C
#843370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#843380000000
0!
0*
09
0>
0C
#843390000000
1!
1*
19
1>
1C
#843400000000
0!
0*
09
0>
0C
#843410000000
1!
1*
19
1>
1C
#843420000000
0!
0*
09
0>
0C
#843430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#843440000000
0!
0*
09
0>
0C
#843450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#843460000000
0!
0*
09
0>
0C
#843470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#843480000000
0!
0*
09
0>
0C
#843490000000
1!
1*
b10 6
19
1>
1C
b10 G
#843500000000
0!
0*
09
0>
0C
#843510000000
1!
1*
b11 6
19
1>
1C
b11 G
#843520000000
0!
0*
09
0>
0C
#843530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#843540000000
0!
0*
09
0>
0C
#843550000000
1!
1*
b101 6
19
1>
1C
b101 G
#843560000000
0!
0*
09
0>
0C
#843570000000
1!
1*
b110 6
19
1>
1C
b110 G
#843580000000
0!
0*
09
0>
0C
#843590000000
1!
1*
b111 6
19
1>
1C
b111 G
#843600000000
0!
0*
09
0>
0C
#843610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#843620000000
0!
0*
09
0>
0C
#843630000000
1!
1*
b1 6
19
1>
1C
b1 G
#843640000000
0!
0*
09
0>
0C
#843650000000
1!
1*
b10 6
19
1>
1C
b10 G
#843660000000
0!
0*
09
0>
0C
#843670000000
1!
1*
b11 6
19
1>
1C
b11 G
#843680000000
0!
0*
09
0>
0C
#843690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#843700000000
0!
0*
09
0>
0C
#843710000000
1!
1*
b101 6
19
1>
1C
b101 G
#843720000000
0!
0*
09
0>
0C
#843730000000
1!
1*
b110 6
19
1>
1C
b110 G
#843740000000
0!
0*
09
0>
0C
#843750000000
1!
1*
b111 6
19
1>
1C
b111 G
#843760000000
0!
0*
09
0>
0C
#843770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#843780000000
0!
0*
09
0>
0C
#843790000000
1!
1*
b1 6
19
1>
1C
b1 G
#843800000000
0!
0*
09
0>
0C
#843810000000
1!
1*
b10 6
19
1>
1C
b10 G
#843820000000
0!
0*
09
0>
0C
#843830000000
1!
1*
b11 6
19
1>
1C
b11 G
#843840000000
0!
0*
09
0>
0C
#843850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#843860000000
0!
0*
09
0>
0C
#843870000000
1!
1*
b101 6
19
1>
1C
b101 G
#843880000000
0!
0*
09
0>
0C
#843890000000
1!
1*
b110 6
19
1>
1C
b110 G
#843900000000
0!
0*
09
0>
0C
#843910000000
1!
1*
b111 6
19
1>
1C
b111 G
#843920000000
0!
1"
0*
1+
09
1:
0>
0C
#843930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#843940000000
0!
0*
09
0>
0C
#843950000000
1!
1*
b1 6
19
1>
1C
b1 G
#843960000000
0!
0*
09
0>
0C
#843970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#843980000000
0!
0*
09
0>
0C
#843990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#844000000000
0!
0*
09
0>
0C
#844010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#844020000000
0!
0*
09
0>
0C
#844030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#844040000000
0!
0#
0*
0,
09
0>
0?
0C
#844050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#844060000000
0!
0*
09
0>
0C
#844070000000
1!
1*
19
1>
1C
#844080000000
0!
0*
09
0>
0C
#844090000000
1!
1*
19
1>
1C
#844100000000
0!
0*
09
0>
0C
#844110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#844120000000
0!
0*
09
0>
0C
#844130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#844140000000
0!
0*
09
0>
0C
#844150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#844160000000
0!
0*
09
0>
0C
#844170000000
1!
1*
b10 6
19
1>
1C
b10 G
#844180000000
0!
0*
09
0>
0C
#844190000000
1!
1*
b11 6
19
1>
1C
b11 G
#844200000000
0!
0*
09
0>
0C
#844210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#844220000000
0!
0*
09
0>
0C
#844230000000
1!
1*
b101 6
19
1>
1C
b101 G
#844240000000
0!
0*
09
0>
0C
#844250000000
1!
1*
b110 6
19
1>
1C
b110 G
#844260000000
0!
0*
09
0>
0C
#844270000000
1!
1*
b111 6
19
1>
1C
b111 G
#844280000000
0!
0*
09
0>
0C
#844290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#844300000000
0!
0*
09
0>
0C
#844310000000
1!
1*
b1 6
19
1>
1C
b1 G
#844320000000
0!
0*
09
0>
0C
#844330000000
1!
1*
b10 6
19
1>
1C
b10 G
#844340000000
0!
0*
09
0>
0C
#844350000000
1!
1*
b11 6
19
1>
1C
b11 G
#844360000000
0!
0*
09
0>
0C
#844370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#844380000000
0!
0*
09
0>
0C
#844390000000
1!
1*
b101 6
19
1>
1C
b101 G
#844400000000
0!
0*
09
0>
0C
#844410000000
1!
1*
b110 6
19
1>
1C
b110 G
#844420000000
0!
0*
09
0>
0C
#844430000000
1!
1*
b111 6
19
1>
1C
b111 G
#844440000000
0!
0*
09
0>
0C
#844450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#844460000000
0!
0*
09
0>
0C
#844470000000
1!
1*
b1 6
19
1>
1C
b1 G
#844480000000
0!
0*
09
0>
0C
#844490000000
1!
1*
b10 6
19
1>
1C
b10 G
#844500000000
0!
0*
09
0>
0C
#844510000000
1!
1*
b11 6
19
1>
1C
b11 G
#844520000000
0!
0*
09
0>
0C
#844530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#844540000000
0!
0*
09
0>
0C
#844550000000
1!
1*
b101 6
19
1>
1C
b101 G
#844560000000
0!
0*
09
0>
0C
#844570000000
1!
1*
b110 6
19
1>
1C
b110 G
#844580000000
0!
0*
09
0>
0C
#844590000000
1!
1*
b111 6
19
1>
1C
b111 G
#844600000000
0!
1"
0*
1+
09
1:
0>
0C
#844610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#844620000000
0!
0*
09
0>
0C
#844630000000
1!
1*
b1 6
19
1>
1C
b1 G
#844640000000
0!
0*
09
0>
0C
#844650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#844660000000
0!
0*
09
0>
0C
#844670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#844680000000
0!
0*
09
0>
0C
#844690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#844700000000
0!
0*
09
0>
0C
#844710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#844720000000
0!
0#
0*
0,
09
0>
0?
0C
#844730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#844740000000
0!
0*
09
0>
0C
#844750000000
1!
1*
19
1>
1C
#844760000000
0!
0*
09
0>
0C
#844770000000
1!
1*
19
1>
1C
#844780000000
0!
0*
09
0>
0C
#844790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#844800000000
0!
0*
09
0>
0C
#844810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#844820000000
0!
0*
09
0>
0C
#844830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#844840000000
0!
0*
09
0>
0C
#844850000000
1!
1*
b10 6
19
1>
1C
b10 G
#844860000000
0!
0*
09
0>
0C
#844870000000
1!
1*
b11 6
19
1>
1C
b11 G
#844880000000
0!
0*
09
0>
0C
#844890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#844900000000
0!
0*
09
0>
0C
#844910000000
1!
1*
b101 6
19
1>
1C
b101 G
#844920000000
0!
0*
09
0>
0C
#844930000000
1!
1*
b110 6
19
1>
1C
b110 G
#844940000000
0!
0*
09
0>
0C
#844950000000
1!
1*
b111 6
19
1>
1C
b111 G
#844960000000
0!
0*
09
0>
0C
#844970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#844980000000
0!
0*
09
0>
0C
#844990000000
1!
1*
b1 6
19
1>
1C
b1 G
#845000000000
0!
0*
09
0>
0C
#845010000000
1!
1*
b10 6
19
1>
1C
b10 G
#845020000000
0!
0*
09
0>
0C
#845030000000
1!
1*
b11 6
19
1>
1C
b11 G
#845040000000
0!
0*
09
0>
0C
#845050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#845060000000
0!
0*
09
0>
0C
#845070000000
1!
1*
b101 6
19
1>
1C
b101 G
#845080000000
0!
0*
09
0>
0C
#845090000000
1!
1*
b110 6
19
1>
1C
b110 G
#845100000000
0!
0*
09
0>
0C
#845110000000
1!
1*
b111 6
19
1>
1C
b111 G
#845120000000
0!
0*
09
0>
0C
#845130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#845140000000
0!
0*
09
0>
0C
#845150000000
1!
1*
b1 6
19
1>
1C
b1 G
#845160000000
0!
0*
09
0>
0C
#845170000000
1!
1*
b10 6
19
1>
1C
b10 G
#845180000000
0!
0*
09
0>
0C
#845190000000
1!
1*
b11 6
19
1>
1C
b11 G
#845200000000
0!
0*
09
0>
0C
#845210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#845220000000
0!
0*
09
0>
0C
#845230000000
1!
1*
b101 6
19
1>
1C
b101 G
#845240000000
0!
0*
09
0>
0C
#845250000000
1!
1*
b110 6
19
1>
1C
b110 G
#845260000000
0!
0*
09
0>
0C
#845270000000
1!
1*
b111 6
19
1>
1C
b111 G
#845280000000
0!
1"
0*
1+
09
1:
0>
0C
#845290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#845300000000
0!
0*
09
0>
0C
#845310000000
1!
1*
b1 6
19
1>
1C
b1 G
#845320000000
0!
0*
09
0>
0C
#845330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#845340000000
0!
0*
09
0>
0C
#845350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#845360000000
0!
0*
09
0>
0C
#845370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#845380000000
0!
0*
09
0>
0C
#845390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#845400000000
0!
0#
0*
0,
09
0>
0?
0C
#845410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#845420000000
0!
0*
09
0>
0C
#845430000000
1!
1*
19
1>
1C
#845440000000
0!
0*
09
0>
0C
#845450000000
1!
1*
19
1>
1C
#845460000000
0!
0*
09
0>
0C
#845470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#845480000000
0!
0*
09
0>
0C
#845490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#845500000000
0!
0*
09
0>
0C
#845510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#845520000000
0!
0*
09
0>
0C
#845530000000
1!
1*
b10 6
19
1>
1C
b10 G
#845540000000
0!
0*
09
0>
0C
#845550000000
1!
1*
b11 6
19
1>
1C
b11 G
#845560000000
0!
0*
09
0>
0C
#845570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#845580000000
0!
0*
09
0>
0C
#845590000000
1!
1*
b101 6
19
1>
1C
b101 G
#845600000000
0!
0*
09
0>
0C
#845610000000
1!
1*
b110 6
19
1>
1C
b110 G
#845620000000
0!
0*
09
0>
0C
#845630000000
1!
1*
b111 6
19
1>
1C
b111 G
#845640000000
0!
0*
09
0>
0C
#845650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#845660000000
0!
0*
09
0>
0C
#845670000000
1!
1*
b1 6
19
1>
1C
b1 G
#845680000000
0!
0*
09
0>
0C
#845690000000
1!
1*
b10 6
19
1>
1C
b10 G
#845700000000
0!
0*
09
0>
0C
#845710000000
1!
1*
b11 6
19
1>
1C
b11 G
#845720000000
0!
0*
09
0>
0C
#845730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#845740000000
0!
0*
09
0>
0C
#845750000000
1!
1*
b101 6
19
1>
1C
b101 G
#845760000000
0!
0*
09
0>
0C
#845770000000
1!
1*
b110 6
19
1>
1C
b110 G
#845780000000
0!
0*
09
0>
0C
#845790000000
1!
1*
b111 6
19
1>
1C
b111 G
#845800000000
0!
0*
09
0>
0C
#845810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#845820000000
0!
0*
09
0>
0C
#845830000000
1!
1*
b1 6
19
1>
1C
b1 G
#845840000000
0!
0*
09
0>
0C
#845850000000
1!
1*
b10 6
19
1>
1C
b10 G
#845860000000
0!
0*
09
0>
0C
#845870000000
1!
1*
b11 6
19
1>
1C
b11 G
#845880000000
0!
0*
09
0>
0C
#845890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#845900000000
0!
0*
09
0>
0C
#845910000000
1!
1*
b101 6
19
1>
1C
b101 G
#845920000000
0!
0*
09
0>
0C
#845930000000
1!
1*
b110 6
19
1>
1C
b110 G
#845940000000
0!
0*
09
0>
0C
#845950000000
1!
1*
b111 6
19
1>
1C
b111 G
#845960000000
0!
1"
0*
1+
09
1:
0>
0C
#845970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#845980000000
0!
0*
09
0>
0C
#845990000000
1!
1*
b1 6
19
1>
1C
b1 G
#846000000000
0!
0*
09
0>
0C
#846010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#846020000000
0!
0*
09
0>
0C
#846030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#846040000000
0!
0*
09
0>
0C
#846050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#846060000000
0!
0*
09
0>
0C
#846070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#846080000000
0!
0#
0*
0,
09
0>
0?
0C
#846090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#846100000000
0!
0*
09
0>
0C
#846110000000
1!
1*
19
1>
1C
#846120000000
0!
0*
09
0>
0C
#846130000000
1!
1*
19
1>
1C
#846140000000
0!
0*
09
0>
0C
#846150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#846160000000
0!
0*
09
0>
0C
#846170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#846180000000
0!
0*
09
0>
0C
#846190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#846200000000
0!
0*
09
0>
0C
#846210000000
1!
1*
b10 6
19
1>
1C
b10 G
#846220000000
0!
0*
09
0>
0C
#846230000000
1!
1*
b11 6
19
1>
1C
b11 G
#846240000000
0!
0*
09
0>
0C
#846250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#846260000000
0!
0*
09
0>
0C
#846270000000
1!
1*
b101 6
19
1>
1C
b101 G
#846280000000
0!
0*
09
0>
0C
#846290000000
1!
1*
b110 6
19
1>
1C
b110 G
#846300000000
0!
0*
09
0>
0C
#846310000000
1!
1*
b111 6
19
1>
1C
b111 G
#846320000000
0!
0*
09
0>
0C
#846330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#846340000000
0!
0*
09
0>
0C
#846350000000
1!
1*
b1 6
19
1>
1C
b1 G
#846360000000
0!
0*
09
0>
0C
#846370000000
1!
1*
b10 6
19
1>
1C
b10 G
#846380000000
0!
0*
09
0>
0C
#846390000000
1!
1*
b11 6
19
1>
1C
b11 G
#846400000000
0!
0*
09
0>
0C
#846410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#846420000000
0!
0*
09
0>
0C
#846430000000
1!
1*
b101 6
19
1>
1C
b101 G
#846440000000
0!
0*
09
0>
0C
#846450000000
1!
1*
b110 6
19
1>
1C
b110 G
#846460000000
0!
0*
09
0>
0C
#846470000000
1!
1*
b111 6
19
1>
1C
b111 G
#846480000000
0!
0*
09
0>
0C
#846490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#846500000000
0!
0*
09
0>
0C
#846510000000
1!
1*
b1 6
19
1>
1C
b1 G
#846520000000
0!
0*
09
0>
0C
#846530000000
1!
1*
b10 6
19
1>
1C
b10 G
#846540000000
0!
0*
09
0>
0C
#846550000000
1!
1*
b11 6
19
1>
1C
b11 G
#846560000000
0!
0*
09
0>
0C
#846570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#846580000000
0!
0*
09
0>
0C
#846590000000
1!
1*
b101 6
19
1>
1C
b101 G
#846600000000
0!
0*
09
0>
0C
#846610000000
1!
1*
b110 6
19
1>
1C
b110 G
#846620000000
0!
0*
09
0>
0C
#846630000000
1!
1*
b111 6
19
1>
1C
b111 G
#846640000000
0!
1"
0*
1+
09
1:
0>
0C
#846650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#846660000000
0!
0*
09
0>
0C
#846670000000
1!
1*
b1 6
19
1>
1C
b1 G
#846680000000
0!
0*
09
0>
0C
#846690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#846700000000
0!
0*
09
0>
0C
#846710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#846720000000
0!
0*
09
0>
0C
#846730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#846740000000
0!
0*
09
0>
0C
#846750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#846760000000
0!
0#
0*
0,
09
0>
0?
0C
#846770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#846780000000
0!
0*
09
0>
0C
#846790000000
1!
1*
19
1>
1C
#846800000000
0!
0*
09
0>
0C
#846810000000
1!
1*
19
1>
1C
#846820000000
0!
0*
09
0>
0C
#846830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#846840000000
0!
0*
09
0>
0C
#846850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#846860000000
0!
0*
09
0>
0C
#846870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#846880000000
0!
0*
09
0>
0C
#846890000000
1!
1*
b10 6
19
1>
1C
b10 G
#846900000000
0!
0*
09
0>
0C
#846910000000
1!
1*
b11 6
19
1>
1C
b11 G
#846920000000
0!
0*
09
0>
0C
#846930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#846940000000
0!
0*
09
0>
0C
#846950000000
1!
1*
b101 6
19
1>
1C
b101 G
#846960000000
0!
0*
09
0>
0C
#846970000000
1!
1*
b110 6
19
1>
1C
b110 G
#846980000000
0!
0*
09
0>
0C
#846990000000
1!
1*
b111 6
19
1>
1C
b111 G
#847000000000
0!
0*
09
0>
0C
#847010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#847020000000
0!
0*
09
0>
0C
#847030000000
1!
1*
b1 6
19
1>
1C
b1 G
#847040000000
0!
0*
09
0>
0C
#847050000000
1!
1*
b10 6
19
1>
1C
b10 G
#847060000000
0!
0*
09
0>
0C
#847070000000
1!
1*
b11 6
19
1>
1C
b11 G
#847080000000
0!
0*
09
0>
0C
#847090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#847100000000
0!
0*
09
0>
0C
#847110000000
1!
1*
b101 6
19
1>
1C
b101 G
#847120000000
0!
0*
09
0>
0C
#847130000000
1!
1*
b110 6
19
1>
1C
b110 G
#847140000000
0!
0*
09
0>
0C
#847150000000
1!
1*
b111 6
19
1>
1C
b111 G
#847160000000
0!
0*
09
0>
0C
#847170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#847180000000
0!
0*
09
0>
0C
#847190000000
1!
1*
b1 6
19
1>
1C
b1 G
#847200000000
0!
0*
09
0>
0C
#847210000000
1!
1*
b10 6
19
1>
1C
b10 G
#847220000000
0!
0*
09
0>
0C
#847230000000
1!
1*
b11 6
19
1>
1C
b11 G
#847240000000
0!
0*
09
0>
0C
#847250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#847260000000
0!
0*
09
0>
0C
#847270000000
1!
1*
b101 6
19
1>
1C
b101 G
#847280000000
0!
0*
09
0>
0C
#847290000000
1!
1*
b110 6
19
1>
1C
b110 G
#847300000000
0!
0*
09
0>
0C
#847310000000
1!
1*
b111 6
19
1>
1C
b111 G
#847320000000
0!
1"
0*
1+
09
1:
0>
0C
#847330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#847340000000
0!
0*
09
0>
0C
#847350000000
1!
1*
b1 6
19
1>
1C
b1 G
#847360000000
0!
0*
09
0>
0C
#847370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#847380000000
0!
0*
09
0>
0C
#847390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#847400000000
0!
0*
09
0>
0C
#847410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#847420000000
0!
0*
09
0>
0C
#847430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#847440000000
0!
0#
0*
0,
09
0>
0?
0C
#847450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#847460000000
0!
0*
09
0>
0C
#847470000000
1!
1*
19
1>
1C
#847480000000
0!
0*
09
0>
0C
#847490000000
1!
1*
19
1>
1C
#847500000000
0!
0*
09
0>
0C
#847510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#847520000000
0!
0*
09
0>
0C
#847530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#847540000000
0!
0*
09
0>
0C
#847550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#847560000000
0!
0*
09
0>
0C
#847570000000
1!
1*
b10 6
19
1>
1C
b10 G
#847580000000
0!
0*
09
0>
0C
#847590000000
1!
1*
b11 6
19
1>
1C
b11 G
#847600000000
0!
0*
09
0>
0C
#847610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#847620000000
0!
0*
09
0>
0C
#847630000000
1!
1*
b101 6
19
1>
1C
b101 G
#847640000000
0!
0*
09
0>
0C
#847650000000
1!
1*
b110 6
19
1>
1C
b110 G
#847660000000
0!
0*
09
0>
0C
#847670000000
1!
1*
b111 6
19
1>
1C
b111 G
#847680000000
0!
0*
09
0>
0C
#847690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#847700000000
0!
0*
09
0>
0C
#847710000000
1!
1*
b1 6
19
1>
1C
b1 G
#847720000000
0!
0*
09
0>
0C
#847730000000
1!
1*
b10 6
19
1>
1C
b10 G
#847740000000
0!
0*
09
0>
0C
#847750000000
1!
1*
b11 6
19
1>
1C
b11 G
#847760000000
0!
0*
09
0>
0C
#847770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#847780000000
0!
0*
09
0>
0C
#847790000000
1!
1*
b101 6
19
1>
1C
b101 G
#847800000000
0!
0*
09
0>
0C
#847810000000
1!
1*
b110 6
19
1>
1C
b110 G
#847820000000
0!
0*
09
0>
0C
#847830000000
1!
1*
b111 6
19
1>
1C
b111 G
#847840000000
0!
0*
09
0>
0C
#847850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#847860000000
0!
0*
09
0>
0C
#847870000000
1!
1*
b1 6
19
1>
1C
b1 G
#847880000000
0!
0*
09
0>
0C
#847890000000
1!
1*
b10 6
19
1>
1C
b10 G
#847900000000
0!
0*
09
0>
0C
#847910000000
1!
1*
b11 6
19
1>
1C
b11 G
#847920000000
0!
0*
09
0>
0C
#847930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#847940000000
0!
0*
09
0>
0C
#847950000000
1!
1*
b101 6
19
1>
1C
b101 G
#847960000000
0!
0*
09
0>
0C
#847970000000
1!
1*
b110 6
19
1>
1C
b110 G
#847980000000
0!
0*
09
0>
0C
#847990000000
1!
1*
b111 6
19
1>
1C
b111 G
#848000000000
0!
1"
0*
1+
09
1:
0>
0C
#848010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#848020000000
0!
0*
09
0>
0C
#848030000000
1!
1*
b1 6
19
1>
1C
b1 G
#848040000000
0!
0*
09
0>
0C
#848050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#848060000000
0!
0*
09
0>
0C
#848070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#848080000000
0!
0*
09
0>
0C
#848090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#848100000000
0!
0*
09
0>
0C
#848110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#848120000000
0!
0#
0*
0,
09
0>
0?
0C
#848130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#848140000000
0!
0*
09
0>
0C
#848150000000
1!
1*
19
1>
1C
#848160000000
0!
0*
09
0>
0C
#848170000000
1!
1*
19
1>
1C
#848180000000
0!
0*
09
0>
0C
#848190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#848200000000
0!
0*
09
0>
0C
#848210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#848220000000
0!
0*
09
0>
0C
#848230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#848240000000
0!
0*
09
0>
0C
#848250000000
1!
1*
b10 6
19
1>
1C
b10 G
#848260000000
0!
0*
09
0>
0C
#848270000000
1!
1*
b11 6
19
1>
1C
b11 G
#848280000000
0!
0*
09
0>
0C
#848290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#848300000000
0!
0*
09
0>
0C
#848310000000
1!
1*
b101 6
19
1>
1C
b101 G
#848320000000
0!
0*
09
0>
0C
#848330000000
1!
1*
b110 6
19
1>
1C
b110 G
#848340000000
0!
0*
09
0>
0C
#848350000000
1!
1*
b111 6
19
1>
1C
b111 G
#848360000000
0!
0*
09
0>
0C
#848370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#848380000000
0!
0*
09
0>
0C
#848390000000
1!
1*
b1 6
19
1>
1C
b1 G
#848400000000
0!
0*
09
0>
0C
#848410000000
1!
1*
b10 6
19
1>
1C
b10 G
#848420000000
0!
0*
09
0>
0C
#848430000000
1!
1*
b11 6
19
1>
1C
b11 G
#848440000000
0!
0*
09
0>
0C
#848450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#848460000000
0!
0*
09
0>
0C
#848470000000
1!
1*
b101 6
19
1>
1C
b101 G
#848480000000
0!
0*
09
0>
0C
#848490000000
1!
1*
b110 6
19
1>
1C
b110 G
#848500000000
0!
0*
09
0>
0C
#848510000000
1!
1*
b111 6
19
1>
1C
b111 G
#848520000000
0!
0*
09
0>
0C
#848530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#848540000000
0!
0*
09
0>
0C
#848550000000
1!
1*
b1 6
19
1>
1C
b1 G
#848560000000
0!
0*
09
0>
0C
#848570000000
1!
1*
b10 6
19
1>
1C
b10 G
#848580000000
0!
0*
09
0>
0C
#848590000000
1!
1*
b11 6
19
1>
1C
b11 G
#848600000000
0!
0*
09
0>
0C
#848610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#848620000000
0!
0*
09
0>
0C
#848630000000
1!
1*
b101 6
19
1>
1C
b101 G
#848640000000
0!
0*
09
0>
0C
#848650000000
1!
1*
b110 6
19
1>
1C
b110 G
#848660000000
0!
0*
09
0>
0C
#848670000000
1!
1*
b111 6
19
1>
1C
b111 G
#848680000000
0!
1"
0*
1+
09
1:
0>
0C
#848690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#848700000000
0!
0*
09
0>
0C
#848710000000
1!
1*
b1 6
19
1>
1C
b1 G
#848720000000
0!
0*
09
0>
0C
#848730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#848740000000
0!
0*
09
0>
0C
#848750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#848760000000
0!
0*
09
0>
0C
#848770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#848780000000
0!
0*
09
0>
0C
#848790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#848800000000
0!
0#
0*
0,
09
0>
0?
0C
#848810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#848820000000
0!
0*
09
0>
0C
#848830000000
1!
1*
19
1>
1C
#848840000000
0!
0*
09
0>
0C
#848850000000
1!
1*
19
1>
1C
#848860000000
0!
0*
09
0>
0C
#848870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#848880000000
0!
0*
09
0>
0C
#848890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#848900000000
0!
0*
09
0>
0C
#848910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#848920000000
0!
0*
09
0>
0C
#848930000000
1!
1*
b10 6
19
1>
1C
b10 G
#848940000000
0!
0*
09
0>
0C
#848950000000
1!
1*
b11 6
19
1>
1C
b11 G
#848960000000
0!
0*
09
0>
0C
#848970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#848980000000
0!
0*
09
0>
0C
#848990000000
1!
1*
b101 6
19
1>
1C
b101 G
#849000000000
0!
0*
09
0>
0C
#849010000000
1!
1*
b110 6
19
1>
1C
b110 G
#849020000000
0!
0*
09
0>
0C
#849030000000
1!
1*
b111 6
19
1>
1C
b111 G
#849040000000
0!
0*
09
0>
0C
#849050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#849060000000
0!
0*
09
0>
0C
#849070000000
1!
1*
b1 6
19
1>
1C
b1 G
#849080000000
0!
0*
09
0>
0C
#849090000000
1!
1*
b10 6
19
1>
1C
b10 G
#849100000000
0!
0*
09
0>
0C
#849110000000
1!
1*
b11 6
19
1>
1C
b11 G
#849120000000
0!
0*
09
0>
0C
#849130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#849140000000
0!
0*
09
0>
0C
#849150000000
1!
1*
b101 6
19
1>
1C
b101 G
#849160000000
0!
0*
09
0>
0C
#849170000000
1!
1*
b110 6
19
1>
1C
b110 G
#849180000000
0!
0*
09
0>
0C
#849190000000
1!
1*
b111 6
19
1>
1C
b111 G
#849200000000
0!
0*
09
0>
0C
#849210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#849220000000
0!
0*
09
0>
0C
#849230000000
1!
1*
b1 6
19
1>
1C
b1 G
#849240000000
0!
0*
09
0>
0C
#849250000000
1!
1*
b10 6
19
1>
1C
b10 G
#849260000000
0!
0*
09
0>
0C
#849270000000
1!
1*
b11 6
19
1>
1C
b11 G
#849280000000
0!
0*
09
0>
0C
#849290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#849300000000
0!
0*
09
0>
0C
#849310000000
1!
1*
b101 6
19
1>
1C
b101 G
#849320000000
0!
0*
09
0>
0C
#849330000000
1!
1*
b110 6
19
1>
1C
b110 G
#849340000000
0!
0*
09
0>
0C
#849350000000
1!
1*
b111 6
19
1>
1C
b111 G
#849360000000
0!
1"
0*
1+
09
1:
0>
0C
#849370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#849380000000
0!
0*
09
0>
0C
#849390000000
1!
1*
b1 6
19
1>
1C
b1 G
#849400000000
0!
0*
09
0>
0C
#849410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#849420000000
0!
0*
09
0>
0C
#849430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#849440000000
0!
0*
09
0>
0C
#849450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#849460000000
0!
0*
09
0>
0C
#849470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#849480000000
0!
0#
0*
0,
09
0>
0?
0C
#849490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#849500000000
0!
0*
09
0>
0C
#849510000000
1!
1*
19
1>
1C
#849520000000
0!
0*
09
0>
0C
#849530000000
1!
1*
19
1>
1C
#849540000000
0!
0*
09
0>
0C
#849550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#849560000000
0!
0*
09
0>
0C
#849570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#849580000000
0!
0*
09
0>
0C
#849590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#849600000000
0!
0*
09
0>
0C
#849610000000
1!
1*
b10 6
19
1>
1C
b10 G
#849620000000
0!
0*
09
0>
0C
#849630000000
1!
1*
b11 6
19
1>
1C
b11 G
#849640000000
0!
0*
09
0>
0C
#849650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#849660000000
0!
0*
09
0>
0C
#849670000000
1!
1*
b101 6
19
1>
1C
b101 G
#849680000000
0!
0*
09
0>
0C
#849690000000
1!
1*
b110 6
19
1>
1C
b110 G
#849700000000
0!
0*
09
0>
0C
#849710000000
1!
1*
b111 6
19
1>
1C
b111 G
#849720000000
0!
0*
09
0>
0C
#849730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#849740000000
0!
0*
09
0>
0C
#849750000000
1!
1*
b1 6
19
1>
1C
b1 G
#849760000000
0!
0*
09
0>
0C
#849770000000
1!
1*
b10 6
19
1>
1C
b10 G
#849780000000
0!
0*
09
0>
0C
#849790000000
1!
1*
b11 6
19
1>
1C
b11 G
#849800000000
0!
0*
09
0>
0C
#849810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#849820000000
0!
0*
09
0>
0C
#849830000000
1!
1*
b101 6
19
1>
1C
b101 G
#849840000000
0!
0*
09
0>
0C
#849850000000
1!
1*
b110 6
19
1>
1C
b110 G
#849860000000
0!
0*
09
0>
0C
#849870000000
1!
1*
b111 6
19
1>
1C
b111 G
#849880000000
0!
0*
09
0>
0C
#849890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#849900000000
0!
0*
09
0>
0C
#849910000000
1!
1*
b1 6
19
1>
1C
b1 G
#849920000000
0!
0*
09
0>
0C
#849930000000
1!
1*
b10 6
19
1>
1C
b10 G
#849940000000
0!
0*
09
0>
0C
#849950000000
1!
1*
b11 6
19
1>
1C
b11 G
#849960000000
0!
0*
09
0>
0C
#849970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#849980000000
0!
0*
09
0>
0C
#849990000000
1!
1*
b101 6
19
1>
1C
b101 G
#850000000000
0!
0*
09
0>
0C
#850010000000
1!
1*
b110 6
19
1>
1C
b110 G
#850020000000
0!
0*
09
0>
0C
#850030000000
1!
1*
b111 6
19
1>
1C
b111 G
#850040000000
0!
1"
0*
1+
09
1:
0>
0C
#850050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#850060000000
0!
0*
09
0>
0C
#850070000000
1!
1*
b1 6
19
1>
1C
b1 G
#850080000000
0!
0*
09
0>
0C
#850090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#850100000000
0!
0*
09
0>
0C
#850110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#850120000000
0!
0*
09
0>
0C
#850130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#850140000000
0!
0*
09
0>
0C
#850150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#850160000000
0!
0#
0*
0,
09
0>
0?
0C
#850170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#850180000000
0!
0*
09
0>
0C
#850190000000
1!
1*
19
1>
1C
#850200000000
0!
0*
09
0>
0C
#850210000000
1!
1*
19
1>
1C
#850220000000
0!
0*
09
0>
0C
#850230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#850240000000
0!
0*
09
0>
0C
#850250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#850260000000
0!
0*
09
0>
0C
#850270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#850280000000
0!
0*
09
0>
0C
#850290000000
1!
1*
b10 6
19
1>
1C
b10 G
#850300000000
0!
0*
09
0>
0C
#850310000000
1!
1*
b11 6
19
1>
1C
b11 G
#850320000000
0!
0*
09
0>
0C
#850330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#850340000000
0!
0*
09
0>
0C
#850350000000
1!
1*
b101 6
19
1>
1C
b101 G
#850360000000
0!
0*
09
0>
0C
#850370000000
1!
1*
b110 6
19
1>
1C
b110 G
#850380000000
0!
0*
09
0>
0C
#850390000000
1!
1*
b111 6
19
1>
1C
b111 G
#850400000000
0!
0*
09
0>
0C
#850410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#850420000000
0!
0*
09
0>
0C
#850430000000
1!
1*
b1 6
19
1>
1C
b1 G
#850440000000
0!
0*
09
0>
0C
#850450000000
1!
1*
b10 6
19
1>
1C
b10 G
#850460000000
0!
0*
09
0>
0C
#850470000000
1!
1*
b11 6
19
1>
1C
b11 G
#850480000000
0!
0*
09
0>
0C
#850490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#850500000000
0!
0*
09
0>
0C
#850510000000
1!
1*
b101 6
19
1>
1C
b101 G
#850520000000
0!
0*
09
0>
0C
#850530000000
1!
1*
b110 6
19
1>
1C
b110 G
#850540000000
0!
0*
09
0>
0C
#850550000000
1!
1*
b111 6
19
1>
1C
b111 G
#850560000000
0!
0*
09
0>
0C
#850570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#850580000000
0!
0*
09
0>
0C
#850590000000
1!
1*
b1 6
19
1>
1C
b1 G
#850600000000
0!
0*
09
0>
0C
#850610000000
1!
1*
b10 6
19
1>
1C
b10 G
#850620000000
0!
0*
09
0>
0C
#850630000000
1!
1*
b11 6
19
1>
1C
b11 G
#850640000000
0!
0*
09
0>
0C
#850650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#850660000000
0!
0*
09
0>
0C
#850670000000
1!
1*
b101 6
19
1>
1C
b101 G
#850680000000
0!
0*
09
0>
0C
#850690000000
1!
1*
b110 6
19
1>
1C
b110 G
#850700000000
0!
0*
09
0>
0C
#850710000000
1!
1*
b111 6
19
1>
1C
b111 G
#850720000000
0!
1"
0*
1+
09
1:
0>
0C
#850730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#850740000000
0!
0*
09
0>
0C
#850750000000
1!
1*
b1 6
19
1>
1C
b1 G
#850760000000
0!
0*
09
0>
0C
#850770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#850780000000
0!
0*
09
0>
0C
#850790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#850800000000
0!
0*
09
0>
0C
#850810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#850820000000
0!
0*
09
0>
0C
#850830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#850840000000
0!
0#
0*
0,
09
0>
0?
0C
#850850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#850860000000
0!
0*
09
0>
0C
#850870000000
1!
1*
19
1>
1C
#850880000000
0!
0*
09
0>
0C
#850890000000
1!
1*
19
1>
1C
#850900000000
0!
0*
09
0>
0C
#850910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#850920000000
0!
0*
09
0>
0C
#850930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#850940000000
0!
0*
09
0>
0C
#850950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#850960000000
0!
0*
09
0>
0C
#850970000000
1!
1*
b10 6
19
1>
1C
b10 G
#850980000000
0!
0*
09
0>
0C
#850990000000
1!
1*
b11 6
19
1>
1C
b11 G
#851000000000
0!
0*
09
0>
0C
#851010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#851020000000
0!
0*
09
0>
0C
#851030000000
1!
1*
b101 6
19
1>
1C
b101 G
#851040000000
0!
0*
09
0>
0C
#851050000000
1!
1*
b110 6
19
1>
1C
b110 G
#851060000000
0!
0*
09
0>
0C
#851070000000
1!
1*
b111 6
19
1>
1C
b111 G
#851080000000
0!
0*
09
0>
0C
#851090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#851100000000
0!
0*
09
0>
0C
#851110000000
1!
1*
b1 6
19
1>
1C
b1 G
#851120000000
0!
0*
09
0>
0C
#851130000000
1!
1*
b10 6
19
1>
1C
b10 G
#851140000000
0!
0*
09
0>
0C
#851150000000
1!
1*
b11 6
19
1>
1C
b11 G
#851160000000
0!
0*
09
0>
0C
#851170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#851180000000
0!
0*
09
0>
0C
#851190000000
1!
1*
b101 6
19
1>
1C
b101 G
#851200000000
0!
0*
09
0>
0C
#851210000000
1!
1*
b110 6
19
1>
1C
b110 G
#851220000000
0!
0*
09
0>
0C
#851230000000
1!
1*
b111 6
19
1>
1C
b111 G
#851240000000
0!
0*
09
0>
0C
#851250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#851260000000
0!
0*
09
0>
0C
#851270000000
1!
1*
b1 6
19
1>
1C
b1 G
#851280000000
0!
0*
09
0>
0C
#851290000000
1!
1*
b10 6
19
1>
1C
b10 G
#851300000000
0!
0*
09
0>
0C
#851310000000
1!
1*
b11 6
19
1>
1C
b11 G
#851320000000
0!
0*
09
0>
0C
#851330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#851340000000
0!
0*
09
0>
0C
#851350000000
1!
1*
b101 6
19
1>
1C
b101 G
#851360000000
0!
0*
09
0>
0C
#851370000000
1!
1*
b110 6
19
1>
1C
b110 G
#851380000000
0!
0*
09
0>
0C
#851390000000
1!
1*
b111 6
19
1>
1C
b111 G
#851400000000
0!
1"
0*
1+
09
1:
0>
0C
#851410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#851420000000
0!
0*
09
0>
0C
#851430000000
1!
1*
b1 6
19
1>
1C
b1 G
#851440000000
0!
0*
09
0>
0C
#851450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#851460000000
0!
0*
09
0>
0C
#851470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#851480000000
0!
0*
09
0>
0C
#851490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#851500000000
0!
0*
09
0>
0C
#851510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#851520000000
0!
0#
0*
0,
09
0>
0?
0C
#851530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#851540000000
0!
0*
09
0>
0C
#851550000000
1!
1*
19
1>
1C
#851560000000
0!
0*
09
0>
0C
#851570000000
1!
1*
19
1>
1C
#851580000000
0!
0*
09
0>
0C
#851590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#851600000000
0!
0*
09
0>
0C
#851610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#851620000000
0!
0*
09
0>
0C
#851630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#851640000000
0!
0*
09
0>
0C
#851650000000
1!
1*
b10 6
19
1>
1C
b10 G
#851660000000
0!
0*
09
0>
0C
#851670000000
1!
1*
b11 6
19
1>
1C
b11 G
#851680000000
0!
0*
09
0>
0C
#851690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#851700000000
0!
0*
09
0>
0C
#851710000000
1!
1*
b101 6
19
1>
1C
b101 G
#851720000000
0!
0*
09
0>
0C
#851730000000
1!
1*
b110 6
19
1>
1C
b110 G
#851740000000
0!
0*
09
0>
0C
#851750000000
1!
1*
b111 6
19
1>
1C
b111 G
#851760000000
0!
0*
09
0>
0C
#851770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#851780000000
0!
0*
09
0>
0C
#851790000000
1!
1*
b1 6
19
1>
1C
b1 G
#851800000000
0!
0*
09
0>
0C
#851810000000
1!
1*
b10 6
19
1>
1C
b10 G
#851820000000
0!
0*
09
0>
0C
#851830000000
1!
1*
b11 6
19
1>
1C
b11 G
#851840000000
0!
0*
09
0>
0C
#851850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#851860000000
0!
0*
09
0>
0C
#851870000000
1!
1*
b101 6
19
1>
1C
b101 G
#851880000000
0!
0*
09
0>
0C
#851890000000
1!
1*
b110 6
19
1>
1C
b110 G
#851900000000
0!
0*
09
0>
0C
#851910000000
1!
1*
b111 6
19
1>
1C
b111 G
#851920000000
0!
0*
09
0>
0C
#851930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#851940000000
0!
0*
09
0>
0C
#851950000000
1!
1*
b1 6
19
1>
1C
b1 G
#851960000000
0!
0*
09
0>
0C
#851970000000
1!
1*
b10 6
19
1>
1C
b10 G
#851980000000
0!
0*
09
0>
0C
#851990000000
1!
1*
b11 6
19
1>
1C
b11 G
#852000000000
0!
0*
09
0>
0C
#852010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#852020000000
0!
0*
09
0>
0C
#852030000000
1!
1*
b101 6
19
1>
1C
b101 G
#852040000000
0!
0*
09
0>
0C
#852050000000
1!
1*
b110 6
19
1>
1C
b110 G
#852060000000
0!
0*
09
0>
0C
#852070000000
1!
1*
b111 6
19
1>
1C
b111 G
#852080000000
0!
1"
0*
1+
09
1:
0>
0C
#852090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#852100000000
0!
0*
09
0>
0C
#852110000000
1!
1*
b1 6
19
1>
1C
b1 G
#852120000000
0!
0*
09
0>
0C
#852130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#852140000000
0!
0*
09
0>
0C
#852150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#852160000000
0!
0*
09
0>
0C
#852170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#852180000000
0!
0*
09
0>
0C
#852190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#852200000000
0!
0#
0*
0,
09
0>
0?
0C
#852210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#852220000000
0!
0*
09
0>
0C
#852230000000
1!
1*
19
1>
1C
#852240000000
0!
0*
09
0>
0C
#852250000000
1!
1*
19
1>
1C
#852260000000
0!
0*
09
0>
0C
#852270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#852280000000
0!
0*
09
0>
0C
#852290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#852300000000
0!
0*
09
0>
0C
#852310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#852320000000
0!
0*
09
0>
0C
#852330000000
1!
1*
b10 6
19
1>
1C
b10 G
#852340000000
0!
0*
09
0>
0C
#852350000000
1!
1*
b11 6
19
1>
1C
b11 G
#852360000000
0!
0*
09
0>
0C
#852370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#852380000000
0!
0*
09
0>
0C
#852390000000
1!
1*
b101 6
19
1>
1C
b101 G
#852400000000
0!
0*
09
0>
0C
#852410000000
1!
1*
b110 6
19
1>
1C
b110 G
#852420000000
0!
0*
09
0>
0C
#852430000000
1!
1*
b111 6
19
1>
1C
b111 G
#852440000000
0!
0*
09
0>
0C
#852450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#852460000000
0!
0*
09
0>
0C
#852470000000
1!
1*
b1 6
19
1>
1C
b1 G
#852480000000
0!
0*
09
0>
0C
#852490000000
1!
1*
b10 6
19
1>
1C
b10 G
#852500000000
0!
0*
09
0>
0C
#852510000000
1!
1*
b11 6
19
1>
1C
b11 G
#852520000000
0!
0*
09
0>
0C
#852530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#852540000000
0!
0*
09
0>
0C
#852550000000
1!
1*
b101 6
19
1>
1C
b101 G
#852560000000
0!
0*
09
0>
0C
#852570000000
1!
1*
b110 6
19
1>
1C
b110 G
#852580000000
0!
0*
09
0>
0C
#852590000000
1!
1*
b111 6
19
1>
1C
b111 G
#852600000000
0!
0*
09
0>
0C
#852610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#852620000000
0!
0*
09
0>
0C
#852630000000
1!
1*
b1 6
19
1>
1C
b1 G
#852640000000
0!
0*
09
0>
0C
#852650000000
1!
1*
b10 6
19
1>
1C
b10 G
#852660000000
0!
0*
09
0>
0C
#852670000000
1!
1*
b11 6
19
1>
1C
b11 G
#852680000000
0!
0*
09
0>
0C
#852690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#852700000000
0!
0*
09
0>
0C
#852710000000
1!
1*
b101 6
19
1>
1C
b101 G
#852720000000
0!
0*
09
0>
0C
#852730000000
1!
1*
b110 6
19
1>
1C
b110 G
#852740000000
0!
0*
09
0>
0C
#852750000000
1!
1*
b111 6
19
1>
1C
b111 G
#852760000000
0!
1"
0*
1+
09
1:
0>
0C
#852770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#852780000000
0!
0*
09
0>
0C
#852790000000
1!
1*
b1 6
19
1>
1C
b1 G
#852800000000
0!
0*
09
0>
0C
#852810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#852820000000
0!
0*
09
0>
0C
#852830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#852840000000
0!
0*
09
0>
0C
#852850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#852860000000
0!
0*
09
0>
0C
#852870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#852880000000
0!
0#
0*
0,
09
0>
0?
0C
#852890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#852900000000
0!
0*
09
0>
0C
#852910000000
1!
1*
19
1>
1C
#852920000000
0!
0*
09
0>
0C
#852930000000
1!
1*
19
1>
1C
#852940000000
0!
0*
09
0>
0C
#852950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#852960000000
0!
0*
09
0>
0C
#852970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#852980000000
0!
0*
09
0>
0C
#852990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#853000000000
0!
0*
09
0>
0C
#853010000000
1!
1*
b10 6
19
1>
1C
b10 G
#853020000000
0!
0*
09
0>
0C
#853030000000
1!
1*
b11 6
19
1>
1C
b11 G
#853040000000
0!
0*
09
0>
0C
#853050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#853060000000
0!
0*
09
0>
0C
#853070000000
1!
1*
b101 6
19
1>
1C
b101 G
#853080000000
0!
0*
09
0>
0C
#853090000000
1!
1*
b110 6
19
1>
1C
b110 G
#853100000000
0!
0*
09
0>
0C
#853110000000
1!
1*
b111 6
19
1>
1C
b111 G
#853120000000
0!
0*
09
0>
0C
#853130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#853140000000
0!
0*
09
0>
0C
#853150000000
1!
1*
b1 6
19
1>
1C
b1 G
#853160000000
0!
0*
09
0>
0C
#853170000000
1!
1*
b10 6
19
1>
1C
b10 G
#853180000000
0!
0*
09
0>
0C
#853190000000
1!
1*
b11 6
19
1>
1C
b11 G
#853200000000
0!
0*
09
0>
0C
#853210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#853220000000
0!
0*
09
0>
0C
#853230000000
1!
1*
b101 6
19
1>
1C
b101 G
#853240000000
0!
0*
09
0>
0C
#853250000000
1!
1*
b110 6
19
1>
1C
b110 G
#853260000000
0!
0*
09
0>
0C
#853270000000
1!
1*
b111 6
19
1>
1C
b111 G
#853280000000
0!
0*
09
0>
0C
#853290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#853300000000
0!
0*
09
0>
0C
#853310000000
1!
1*
b1 6
19
1>
1C
b1 G
#853320000000
0!
0*
09
0>
0C
#853330000000
1!
1*
b10 6
19
1>
1C
b10 G
#853340000000
0!
0*
09
0>
0C
#853350000000
1!
1*
b11 6
19
1>
1C
b11 G
#853360000000
0!
0*
09
0>
0C
#853370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#853380000000
0!
0*
09
0>
0C
#853390000000
1!
1*
b101 6
19
1>
1C
b101 G
#853400000000
0!
0*
09
0>
0C
#853410000000
1!
1*
b110 6
19
1>
1C
b110 G
#853420000000
0!
0*
09
0>
0C
#853430000000
1!
1*
b111 6
19
1>
1C
b111 G
#853440000000
0!
1"
0*
1+
09
1:
0>
0C
#853450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#853460000000
0!
0*
09
0>
0C
#853470000000
1!
1*
b1 6
19
1>
1C
b1 G
#853480000000
0!
0*
09
0>
0C
#853490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#853500000000
0!
0*
09
0>
0C
#853510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#853520000000
0!
0*
09
0>
0C
#853530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#853540000000
0!
0*
09
0>
0C
#853550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#853560000000
0!
0#
0*
0,
09
0>
0?
0C
#853570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#853580000000
0!
0*
09
0>
0C
#853590000000
1!
1*
19
1>
1C
#853600000000
0!
0*
09
0>
0C
#853610000000
1!
1*
19
1>
1C
#853620000000
0!
0*
09
0>
0C
#853630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#853640000000
0!
0*
09
0>
0C
#853650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#853660000000
0!
0*
09
0>
0C
#853670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#853680000000
0!
0*
09
0>
0C
#853690000000
1!
1*
b10 6
19
1>
1C
b10 G
#853700000000
0!
0*
09
0>
0C
#853710000000
1!
1*
b11 6
19
1>
1C
b11 G
#853720000000
0!
0*
09
0>
0C
#853730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#853740000000
0!
0*
09
0>
0C
#853750000000
1!
1*
b101 6
19
1>
1C
b101 G
#853760000000
0!
0*
09
0>
0C
#853770000000
1!
1*
b110 6
19
1>
1C
b110 G
#853780000000
0!
0*
09
0>
0C
#853790000000
1!
1*
b111 6
19
1>
1C
b111 G
#853800000000
0!
0*
09
0>
0C
#853810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#853820000000
0!
0*
09
0>
0C
#853830000000
1!
1*
b1 6
19
1>
1C
b1 G
#853840000000
0!
0*
09
0>
0C
#853850000000
1!
1*
b10 6
19
1>
1C
b10 G
#853860000000
0!
0*
09
0>
0C
#853870000000
1!
1*
b11 6
19
1>
1C
b11 G
#853880000000
0!
0*
09
0>
0C
#853890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#853900000000
0!
0*
09
0>
0C
#853910000000
1!
1*
b101 6
19
1>
1C
b101 G
#853920000000
0!
0*
09
0>
0C
#853930000000
1!
1*
b110 6
19
1>
1C
b110 G
#853940000000
0!
0*
09
0>
0C
#853950000000
1!
1*
b111 6
19
1>
1C
b111 G
#853960000000
0!
0*
09
0>
0C
#853970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#853980000000
0!
0*
09
0>
0C
#853990000000
1!
1*
b1 6
19
1>
1C
b1 G
#854000000000
0!
0*
09
0>
0C
#854010000000
1!
1*
b10 6
19
1>
1C
b10 G
#854020000000
0!
0*
09
0>
0C
#854030000000
1!
1*
b11 6
19
1>
1C
b11 G
#854040000000
0!
0*
09
0>
0C
#854050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#854060000000
0!
0*
09
0>
0C
#854070000000
1!
1*
b101 6
19
1>
1C
b101 G
#854080000000
0!
0*
09
0>
0C
#854090000000
1!
1*
b110 6
19
1>
1C
b110 G
#854100000000
0!
0*
09
0>
0C
#854110000000
1!
1*
b111 6
19
1>
1C
b111 G
#854120000000
0!
1"
0*
1+
09
1:
0>
0C
#854130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#854140000000
0!
0*
09
0>
0C
#854150000000
1!
1*
b1 6
19
1>
1C
b1 G
#854160000000
0!
0*
09
0>
0C
#854170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#854180000000
0!
0*
09
0>
0C
#854190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#854200000000
0!
0*
09
0>
0C
#854210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#854220000000
0!
0*
09
0>
0C
#854230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#854240000000
0!
0#
0*
0,
09
0>
0?
0C
#854250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#854260000000
0!
0*
09
0>
0C
#854270000000
1!
1*
19
1>
1C
#854280000000
0!
0*
09
0>
0C
#854290000000
1!
1*
19
1>
1C
#854300000000
0!
0*
09
0>
0C
#854310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#854320000000
0!
0*
09
0>
0C
#854330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#854340000000
0!
0*
09
0>
0C
#854350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#854360000000
0!
0*
09
0>
0C
#854370000000
1!
1*
b10 6
19
1>
1C
b10 G
#854380000000
0!
0*
09
0>
0C
#854390000000
1!
1*
b11 6
19
1>
1C
b11 G
#854400000000
0!
0*
09
0>
0C
#854410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#854420000000
0!
0*
09
0>
0C
#854430000000
1!
1*
b101 6
19
1>
1C
b101 G
#854440000000
0!
0*
09
0>
0C
#854450000000
1!
1*
b110 6
19
1>
1C
b110 G
#854460000000
0!
0*
09
0>
0C
#854470000000
1!
1*
b111 6
19
1>
1C
b111 G
#854480000000
0!
0*
09
0>
0C
#854490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#854500000000
0!
0*
09
0>
0C
#854510000000
1!
1*
b1 6
19
1>
1C
b1 G
#854520000000
0!
0*
09
0>
0C
#854530000000
1!
1*
b10 6
19
1>
1C
b10 G
#854540000000
0!
0*
09
0>
0C
#854550000000
1!
1*
b11 6
19
1>
1C
b11 G
#854560000000
0!
0*
09
0>
0C
#854570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#854580000000
0!
0*
09
0>
0C
#854590000000
1!
1*
b101 6
19
1>
1C
b101 G
#854600000000
0!
0*
09
0>
0C
#854610000000
1!
1*
b110 6
19
1>
1C
b110 G
#854620000000
0!
0*
09
0>
0C
#854630000000
1!
1*
b111 6
19
1>
1C
b111 G
#854640000000
0!
0*
09
0>
0C
#854650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#854660000000
0!
0*
09
0>
0C
#854670000000
1!
1*
b1 6
19
1>
1C
b1 G
#854680000000
0!
0*
09
0>
0C
#854690000000
1!
1*
b10 6
19
1>
1C
b10 G
#854700000000
0!
0*
09
0>
0C
#854710000000
1!
1*
b11 6
19
1>
1C
b11 G
#854720000000
0!
0*
09
0>
0C
#854730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#854740000000
0!
0*
09
0>
0C
#854750000000
1!
1*
b101 6
19
1>
1C
b101 G
#854760000000
0!
0*
09
0>
0C
#854770000000
1!
1*
b110 6
19
1>
1C
b110 G
#854780000000
0!
0*
09
0>
0C
#854790000000
1!
1*
b111 6
19
1>
1C
b111 G
#854800000000
0!
1"
0*
1+
09
1:
0>
0C
#854810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#854820000000
0!
0*
09
0>
0C
#854830000000
1!
1*
b1 6
19
1>
1C
b1 G
#854840000000
0!
0*
09
0>
0C
#854850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#854860000000
0!
0*
09
0>
0C
#854870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#854880000000
0!
0*
09
0>
0C
#854890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#854900000000
0!
0*
09
0>
0C
#854910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#854920000000
0!
0#
0*
0,
09
0>
0?
0C
#854930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#854940000000
0!
0*
09
0>
0C
#854950000000
1!
1*
19
1>
1C
#854960000000
0!
0*
09
0>
0C
#854970000000
1!
1*
19
1>
1C
#854980000000
0!
0*
09
0>
0C
#854990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#855000000000
0!
0*
09
0>
0C
#855010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#855020000000
0!
0*
09
0>
0C
#855030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#855040000000
0!
0*
09
0>
0C
#855050000000
1!
1*
b10 6
19
1>
1C
b10 G
#855060000000
0!
0*
09
0>
0C
#855070000000
1!
1*
b11 6
19
1>
1C
b11 G
#855080000000
0!
0*
09
0>
0C
#855090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#855100000000
0!
0*
09
0>
0C
#855110000000
1!
1*
b101 6
19
1>
1C
b101 G
#855120000000
0!
0*
09
0>
0C
#855130000000
1!
1*
b110 6
19
1>
1C
b110 G
#855140000000
0!
0*
09
0>
0C
#855150000000
1!
1*
b111 6
19
1>
1C
b111 G
#855160000000
0!
0*
09
0>
0C
#855170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#855180000000
0!
0*
09
0>
0C
#855190000000
1!
1*
b1 6
19
1>
1C
b1 G
#855200000000
0!
0*
09
0>
0C
#855210000000
1!
1*
b10 6
19
1>
1C
b10 G
#855220000000
0!
0*
09
0>
0C
#855230000000
1!
1*
b11 6
19
1>
1C
b11 G
#855240000000
0!
0*
09
0>
0C
#855250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#855260000000
0!
0*
09
0>
0C
#855270000000
1!
1*
b101 6
19
1>
1C
b101 G
#855280000000
0!
0*
09
0>
0C
#855290000000
1!
1*
b110 6
19
1>
1C
b110 G
#855300000000
0!
0*
09
0>
0C
#855310000000
1!
1*
b111 6
19
1>
1C
b111 G
#855320000000
0!
0*
09
0>
0C
#855330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#855340000000
0!
0*
09
0>
0C
#855350000000
1!
1*
b1 6
19
1>
1C
b1 G
#855360000000
0!
0*
09
0>
0C
#855370000000
1!
1*
b10 6
19
1>
1C
b10 G
#855380000000
0!
0*
09
0>
0C
#855390000000
1!
1*
b11 6
19
1>
1C
b11 G
#855400000000
0!
0*
09
0>
0C
#855410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#855420000000
0!
0*
09
0>
0C
#855430000000
1!
1*
b101 6
19
1>
1C
b101 G
#855440000000
0!
0*
09
0>
0C
#855450000000
1!
1*
b110 6
19
1>
1C
b110 G
#855460000000
0!
0*
09
0>
0C
#855470000000
1!
1*
b111 6
19
1>
1C
b111 G
#855480000000
0!
1"
0*
1+
09
1:
0>
0C
#855490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#855500000000
0!
0*
09
0>
0C
#855510000000
1!
1*
b1 6
19
1>
1C
b1 G
#855520000000
0!
0*
09
0>
0C
#855530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#855540000000
0!
0*
09
0>
0C
#855550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#855560000000
0!
0*
09
0>
0C
#855570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#855580000000
0!
0*
09
0>
0C
#855590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#855600000000
0!
0#
0*
0,
09
0>
0?
0C
#855610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#855620000000
0!
0*
09
0>
0C
#855630000000
1!
1*
19
1>
1C
#855640000000
0!
0*
09
0>
0C
#855650000000
1!
1*
19
1>
1C
#855660000000
0!
0*
09
0>
0C
#855670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#855680000000
0!
0*
09
0>
0C
#855690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#855700000000
0!
0*
09
0>
0C
#855710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#855720000000
0!
0*
09
0>
0C
#855730000000
1!
1*
b10 6
19
1>
1C
b10 G
#855740000000
0!
0*
09
0>
0C
#855750000000
1!
1*
b11 6
19
1>
1C
b11 G
#855760000000
0!
0*
09
0>
0C
#855770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#855780000000
0!
0*
09
0>
0C
#855790000000
1!
1*
b101 6
19
1>
1C
b101 G
#855800000000
0!
0*
09
0>
0C
#855810000000
1!
1*
b110 6
19
1>
1C
b110 G
#855820000000
0!
0*
09
0>
0C
#855830000000
1!
1*
b111 6
19
1>
1C
b111 G
#855840000000
0!
0*
09
0>
0C
#855850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#855860000000
0!
0*
09
0>
0C
#855870000000
1!
1*
b1 6
19
1>
1C
b1 G
#855880000000
0!
0*
09
0>
0C
#855890000000
1!
1*
b10 6
19
1>
1C
b10 G
#855900000000
0!
0*
09
0>
0C
#855910000000
1!
1*
b11 6
19
1>
1C
b11 G
#855920000000
0!
0*
09
0>
0C
#855930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#855940000000
0!
0*
09
0>
0C
#855950000000
1!
1*
b101 6
19
1>
1C
b101 G
#855960000000
0!
0*
09
0>
0C
#855970000000
1!
1*
b110 6
19
1>
1C
b110 G
#855980000000
0!
0*
09
0>
0C
#855990000000
1!
1*
b111 6
19
1>
1C
b111 G
#856000000000
0!
0*
09
0>
0C
#856010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#856020000000
0!
0*
09
0>
0C
#856030000000
1!
1*
b1 6
19
1>
1C
b1 G
#856040000000
0!
0*
09
0>
0C
#856050000000
1!
1*
b10 6
19
1>
1C
b10 G
#856060000000
0!
0*
09
0>
0C
#856070000000
1!
1*
b11 6
19
1>
1C
b11 G
#856080000000
0!
0*
09
0>
0C
#856090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#856100000000
0!
0*
09
0>
0C
#856110000000
1!
1*
b101 6
19
1>
1C
b101 G
#856120000000
0!
0*
09
0>
0C
#856130000000
1!
1*
b110 6
19
1>
1C
b110 G
#856140000000
0!
0*
09
0>
0C
#856150000000
1!
1*
b111 6
19
1>
1C
b111 G
#856160000000
0!
1"
0*
1+
09
1:
0>
0C
#856170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#856180000000
0!
0*
09
0>
0C
#856190000000
1!
1*
b1 6
19
1>
1C
b1 G
#856200000000
0!
0*
09
0>
0C
#856210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#856220000000
0!
0*
09
0>
0C
#856230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#856240000000
0!
0*
09
0>
0C
#856250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#856260000000
0!
0*
09
0>
0C
#856270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#856280000000
0!
0#
0*
0,
09
0>
0?
0C
#856290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#856300000000
0!
0*
09
0>
0C
#856310000000
1!
1*
19
1>
1C
#856320000000
0!
0*
09
0>
0C
#856330000000
1!
1*
19
1>
1C
#856340000000
0!
0*
09
0>
0C
#856350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#856360000000
0!
0*
09
0>
0C
#856370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#856380000000
0!
0*
09
0>
0C
#856390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#856400000000
0!
0*
09
0>
0C
#856410000000
1!
1*
b10 6
19
1>
1C
b10 G
#856420000000
0!
0*
09
0>
0C
#856430000000
1!
1*
b11 6
19
1>
1C
b11 G
#856440000000
0!
0*
09
0>
0C
#856450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#856460000000
0!
0*
09
0>
0C
#856470000000
1!
1*
b101 6
19
1>
1C
b101 G
#856480000000
0!
0*
09
0>
0C
#856490000000
1!
1*
b110 6
19
1>
1C
b110 G
#856500000000
0!
0*
09
0>
0C
#856510000000
1!
1*
b111 6
19
1>
1C
b111 G
#856520000000
0!
0*
09
0>
0C
#856530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#856540000000
0!
0*
09
0>
0C
#856550000000
1!
1*
b1 6
19
1>
1C
b1 G
#856560000000
0!
0*
09
0>
0C
#856570000000
1!
1*
b10 6
19
1>
1C
b10 G
#856580000000
0!
0*
09
0>
0C
#856590000000
1!
1*
b11 6
19
1>
1C
b11 G
#856600000000
0!
0*
09
0>
0C
#856610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#856620000000
0!
0*
09
0>
0C
#856630000000
1!
1*
b101 6
19
1>
1C
b101 G
#856640000000
0!
0*
09
0>
0C
#856650000000
1!
1*
b110 6
19
1>
1C
b110 G
#856660000000
0!
0*
09
0>
0C
#856670000000
1!
1*
b111 6
19
1>
1C
b111 G
#856680000000
0!
0*
09
0>
0C
#856690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#856700000000
0!
0*
09
0>
0C
#856710000000
1!
1*
b1 6
19
1>
1C
b1 G
#856720000000
0!
0*
09
0>
0C
#856730000000
1!
1*
b10 6
19
1>
1C
b10 G
#856740000000
0!
0*
09
0>
0C
#856750000000
1!
1*
b11 6
19
1>
1C
b11 G
#856760000000
0!
0*
09
0>
0C
#856770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#856780000000
0!
0*
09
0>
0C
#856790000000
1!
1*
b101 6
19
1>
1C
b101 G
#856800000000
0!
0*
09
0>
0C
#856810000000
1!
1*
b110 6
19
1>
1C
b110 G
#856820000000
0!
0*
09
0>
0C
#856830000000
1!
1*
b111 6
19
1>
1C
b111 G
#856840000000
0!
1"
0*
1+
09
1:
0>
0C
#856850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#856860000000
0!
0*
09
0>
0C
#856870000000
1!
1*
b1 6
19
1>
1C
b1 G
#856880000000
0!
0*
09
0>
0C
#856890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#856900000000
0!
0*
09
0>
0C
#856910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#856920000000
0!
0*
09
0>
0C
#856930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#856940000000
0!
0*
09
0>
0C
#856950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#856960000000
0!
0#
0*
0,
09
0>
0?
0C
#856970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#856980000000
0!
0*
09
0>
0C
#856990000000
1!
1*
19
1>
1C
#857000000000
0!
0*
09
0>
0C
#857010000000
1!
1*
19
1>
1C
#857020000000
0!
0*
09
0>
0C
#857030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#857040000000
0!
0*
09
0>
0C
#857050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#857060000000
0!
0*
09
0>
0C
#857070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#857080000000
0!
0*
09
0>
0C
#857090000000
1!
1*
b10 6
19
1>
1C
b10 G
#857100000000
0!
0*
09
0>
0C
#857110000000
1!
1*
b11 6
19
1>
1C
b11 G
#857120000000
0!
0*
09
0>
0C
#857130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#857140000000
0!
0*
09
0>
0C
#857150000000
1!
1*
b101 6
19
1>
1C
b101 G
#857160000000
0!
0*
09
0>
0C
#857170000000
1!
1*
b110 6
19
1>
1C
b110 G
#857180000000
0!
0*
09
0>
0C
#857190000000
1!
1*
b111 6
19
1>
1C
b111 G
#857200000000
0!
0*
09
0>
0C
#857210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#857220000000
0!
0*
09
0>
0C
#857230000000
1!
1*
b1 6
19
1>
1C
b1 G
#857240000000
0!
0*
09
0>
0C
#857250000000
1!
1*
b10 6
19
1>
1C
b10 G
#857260000000
0!
0*
09
0>
0C
#857270000000
1!
1*
b11 6
19
1>
1C
b11 G
#857280000000
0!
0*
09
0>
0C
#857290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#857300000000
0!
0*
09
0>
0C
#857310000000
1!
1*
b101 6
19
1>
1C
b101 G
#857320000000
0!
0*
09
0>
0C
#857330000000
1!
1*
b110 6
19
1>
1C
b110 G
#857340000000
0!
0*
09
0>
0C
#857350000000
1!
1*
b111 6
19
1>
1C
b111 G
#857360000000
0!
0*
09
0>
0C
#857370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#857380000000
0!
0*
09
0>
0C
#857390000000
1!
1*
b1 6
19
1>
1C
b1 G
#857400000000
0!
0*
09
0>
0C
#857410000000
1!
1*
b10 6
19
1>
1C
b10 G
#857420000000
0!
0*
09
0>
0C
#857430000000
1!
1*
b11 6
19
1>
1C
b11 G
#857440000000
0!
0*
09
0>
0C
#857450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#857460000000
0!
0*
09
0>
0C
#857470000000
1!
1*
b101 6
19
1>
1C
b101 G
#857480000000
0!
0*
09
0>
0C
#857490000000
1!
1*
b110 6
19
1>
1C
b110 G
#857500000000
0!
0*
09
0>
0C
#857510000000
1!
1*
b111 6
19
1>
1C
b111 G
#857520000000
0!
1"
0*
1+
09
1:
0>
0C
#857530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#857540000000
0!
0*
09
0>
0C
#857550000000
1!
1*
b1 6
19
1>
1C
b1 G
#857560000000
0!
0*
09
0>
0C
#857570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#857580000000
0!
0*
09
0>
0C
#857590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#857600000000
0!
0*
09
0>
0C
#857610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#857620000000
0!
0*
09
0>
0C
#857630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#857640000000
0!
0#
0*
0,
09
0>
0?
0C
#857650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#857660000000
0!
0*
09
0>
0C
#857670000000
1!
1*
19
1>
1C
#857680000000
0!
0*
09
0>
0C
#857690000000
1!
1*
19
1>
1C
#857700000000
0!
0*
09
0>
0C
#857710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#857720000000
0!
0*
09
0>
0C
#857730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#857740000000
0!
0*
09
0>
0C
#857750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#857760000000
0!
0*
09
0>
0C
#857770000000
1!
1*
b10 6
19
1>
1C
b10 G
#857780000000
0!
0*
09
0>
0C
#857790000000
1!
1*
b11 6
19
1>
1C
b11 G
#857800000000
0!
0*
09
0>
0C
#857810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#857820000000
0!
0*
09
0>
0C
#857830000000
1!
1*
b101 6
19
1>
1C
b101 G
#857840000000
0!
0*
09
0>
0C
#857850000000
1!
1*
b110 6
19
1>
1C
b110 G
#857860000000
0!
0*
09
0>
0C
#857870000000
1!
1*
b111 6
19
1>
1C
b111 G
#857880000000
0!
0*
09
0>
0C
#857890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#857900000000
0!
0*
09
0>
0C
#857910000000
1!
1*
b1 6
19
1>
1C
b1 G
#857920000000
0!
0*
09
0>
0C
#857930000000
1!
1*
b10 6
19
1>
1C
b10 G
#857940000000
0!
0*
09
0>
0C
#857950000000
1!
1*
b11 6
19
1>
1C
b11 G
#857960000000
0!
0*
09
0>
0C
#857970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#857980000000
0!
0*
09
0>
0C
#857990000000
1!
1*
b101 6
19
1>
1C
b101 G
#858000000000
0!
0*
09
0>
0C
#858010000000
1!
1*
b110 6
19
1>
1C
b110 G
#858020000000
0!
0*
09
0>
0C
#858030000000
1!
1*
b111 6
19
1>
1C
b111 G
#858040000000
0!
0*
09
0>
0C
#858050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#858060000000
0!
0*
09
0>
0C
#858070000000
1!
1*
b1 6
19
1>
1C
b1 G
#858080000000
0!
0*
09
0>
0C
#858090000000
1!
1*
b10 6
19
1>
1C
b10 G
#858100000000
0!
0*
09
0>
0C
#858110000000
1!
1*
b11 6
19
1>
1C
b11 G
#858120000000
0!
0*
09
0>
0C
#858130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#858140000000
0!
0*
09
0>
0C
#858150000000
1!
1*
b101 6
19
1>
1C
b101 G
#858160000000
0!
0*
09
0>
0C
#858170000000
1!
1*
b110 6
19
1>
1C
b110 G
#858180000000
0!
0*
09
0>
0C
#858190000000
1!
1*
b111 6
19
1>
1C
b111 G
#858200000000
0!
1"
0*
1+
09
1:
0>
0C
#858210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#858220000000
0!
0*
09
0>
0C
#858230000000
1!
1*
b1 6
19
1>
1C
b1 G
#858240000000
0!
0*
09
0>
0C
#858250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#858260000000
0!
0*
09
0>
0C
#858270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#858280000000
0!
0*
09
0>
0C
#858290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#858300000000
0!
0*
09
0>
0C
#858310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#858320000000
0!
0#
0*
0,
09
0>
0?
0C
#858330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#858340000000
0!
0*
09
0>
0C
#858350000000
1!
1*
19
1>
1C
#858360000000
0!
0*
09
0>
0C
#858370000000
1!
1*
19
1>
1C
#858380000000
0!
0*
09
0>
0C
#858390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#858400000000
0!
0*
09
0>
0C
#858410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#858420000000
0!
0*
09
0>
0C
#858430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#858440000000
0!
0*
09
0>
0C
#858450000000
1!
1*
b10 6
19
1>
1C
b10 G
#858460000000
0!
0*
09
0>
0C
#858470000000
1!
1*
b11 6
19
1>
1C
b11 G
#858480000000
0!
0*
09
0>
0C
#858490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#858500000000
0!
0*
09
0>
0C
#858510000000
1!
1*
b101 6
19
1>
1C
b101 G
#858520000000
0!
0*
09
0>
0C
#858530000000
1!
1*
b110 6
19
1>
1C
b110 G
#858540000000
0!
0*
09
0>
0C
#858550000000
1!
1*
b111 6
19
1>
1C
b111 G
#858560000000
0!
0*
09
0>
0C
#858570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#858580000000
0!
0*
09
0>
0C
#858590000000
1!
1*
b1 6
19
1>
1C
b1 G
#858600000000
0!
0*
09
0>
0C
#858610000000
1!
1*
b10 6
19
1>
1C
b10 G
#858620000000
0!
0*
09
0>
0C
#858630000000
1!
1*
b11 6
19
1>
1C
b11 G
#858640000000
0!
0*
09
0>
0C
#858650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#858660000000
0!
0*
09
0>
0C
#858670000000
1!
1*
b101 6
19
1>
1C
b101 G
#858680000000
0!
0*
09
0>
0C
#858690000000
1!
1*
b110 6
19
1>
1C
b110 G
#858700000000
0!
0*
09
0>
0C
#858710000000
1!
1*
b111 6
19
1>
1C
b111 G
#858720000000
0!
0*
09
0>
0C
#858730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#858740000000
0!
0*
09
0>
0C
#858750000000
1!
1*
b1 6
19
1>
1C
b1 G
#858760000000
0!
0*
09
0>
0C
#858770000000
1!
1*
b10 6
19
1>
1C
b10 G
#858780000000
0!
0*
09
0>
0C
#858790000000
1!
1*
b11 6
19
1>
1C
b11 G
#858800000000
0!
0*
09
0>
0C
#858810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#858820000000
0!
0*
09
0>
0C
#858830000000
1!
1*
b101 6
19
1>
1C
b101 G
#858840000000
0!
0*
09
0>
0C
#858850000000
1!
1*
b110 6
19
1>
1C
b110 G
#858860000000
0!
0*
09
0>
0C
#858870000000
1!
1*
b111 6
19
1>
1C
b111 G
#858880000000
0!
1"
0*
1+
09
1:
0>
0C
#858890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#858900000000
0!
0*
09
0>
0C
#858910000000
1!
1*
b1 6
19
1>
1C
b1 G
#858920000000
0!
0*
09
0>
0C
#858930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#858940000000
0!
0*
09
0>
0C
#858950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#858960000000
0!
0*
09
0>
0C
#858970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#858980000000
0!
0*
09
0>
0C
#858990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#859000000000
0!
0#
0*
0,
09
0>
0?
0C
#859010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#859020000000
0!
0*
09
0>
0C
#859030000000
1!
1*
19
1>
1C
#859040000000
0!
0*
09
0>
0C
#859050000000
1!
1*
19
1>
1C
#859060000000
0!
0*
09
0>
0C
#859070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#859080000000
0!
0*
09
0>
0C
#859090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#859100000000
0!
0*
09
0>
0C
#859110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#859120000000
0!
0*
09
0>
0C
#859130000000
1!
1*
b10 6
19
1>
1C
b10 G
#859140000000
0!
0*
09
0>
0C
#859150000000
1!
1*
b11 6
19
1>
1C
b11 G
#859160000000
0!
0*
09
0>
0C
#859170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#859180000000
0!
0*
09
0>
0C
#859190000000
1!
1*
b101 6
19
1>
1C
b101 G
#859200000000
0!
0*
09
0>
0C
#859210000000
1!
1*
b110 6
19
1>
1C
b110 G
#859220000000
0!
0*
09
0>
0C
#859230000000
1!
1*
b111 6
19
1>
1C
b111 G
#859240000000
0!
0*
09
0>
0C
#859250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#859260000000
0!
0*
09
0>
0C
#859270000000
1!
1*
b1 6
19
1>
1C
b1 G
#859280000000
0!
0*
09
0>
0C
#859290000000
1!
1*
b10 6
19
1>
1C
b10 G
#859300000000
0!
0*
09
0>
0C
#859310000000
1!
1*
b11 6
19
1>
1C
b11 G
#859320000000
0!
0*
09
0>
0C
#859330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#859340000000
0!
0*
09
0>
0C
#859350000000
1!
1*
b101 6
19
1>
1C
b101 G
#859360000000
0!
0*
09
0>
0C
#859370000000
1!
1*
b110 6
19
1>
1C
b110 G
#859380000000
0!
0*
09
0>
0C
#859390000000
1!
1*
b111 6
19
1>
1C
b111 G
#859400000000
0!
0*
09
0>
0C
#859410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#859420000000
0!
0*
09
0>
0C
#859430000000
1!
1*
b1 6
19
1>
1C
b1 G
#859440000000
0!
0*
09
0>
0C
#859450000000
1!
1*
b10 6
19
1>
1C
b10 G
#859460000000
0!
0*
09
0>
0C
#859470000000
1!
1*
b11 6
19
1>
1C
b11 G
#859480000000
0!
0*
09
0>
0C
#859490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#859500000000
0!
0*
09
0>
0C
#859510000000
1!
1*
b101 6
19
1>
1C
b101 G
#859520000000
0!
0*
09
0>
0C
#859530000000
1!
1*
b110 6
19
1>
1C
b110 G
#859540000000
0!
0*
09
0>
0C
#859550000000
1!
1*
b111 6
19
1>
1C
b111 G
#859560000000
0!
1"
0*
1+
09
1:
0>
0C
#859570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#859580000000
0!
0*
09
0>
0C
#859590000000
1!
1*
b1 6
19
1>
1C
b1 G
#859600000000
0!
0*
09
0>
0C
#859610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#859620000000
0!
0*
09
0>
0C
#859630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#859640000000
0!
0*
09
0>
0C
#859650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#859660000000
0!
0*
09
0>
0C
#859670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#859680000000
0!
0#
0*
0,
09
0>
0?
0C
#859690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#859700000000
0!
0*
09
0>
0C
#859710000000
1!
1*
19
1>
1C
#859720000000
0!
0*
09
0>
0C
#859730000000
1!
1*
19
1>
1C
#859740000000
0!
0*
09
0>
0C
#859750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#859760000000
0!
0*
09
0>
0C
#859770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#859780000000
0!
0*
09
0>
0C
#859790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#859800000000
0!
0*
09
0>
0C
#859810000000
1!
1*
b10 6
19
1>
1C
b10 G
#859820000000
0!
0*
09
0>
0C
#859830000000
1!
1*
b11 6
19
1>
1C
b11 G
#859840000000
0!
0*
09
0>
0C
#859850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#859860000000
0!
0*
09
0>
0C
#859870000000
1!
1*
b101 6
19
1>
1C
b101 G
#859880000000
0!
0*
09
0>
0C
#859890000000
1!
1*
b110 6
19
1>
1C
b110 G
#859900000000
0!
0*
09
0>
0C
#859910000000
1!
1*
b111 6
19
1>
1C
b111 G
#859920000000
0!
0*
09
0>
0C
#859930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#859940000000
0!
0*
09
0>
0C
#859950000000
1!
1*
b1 6
19
1>
1C
b1 G
#859960000000
0!
0*
09
0>
0C
#859970000000
1!
1*
b10 6
19
1>
1C
b10 G
#859980000000
0!
0*
09
0>
0C
#859990000000
1!
1*
b11 6
19
1>
1C
b11 G
#860000000000
0!
0*
09
0>
0C
#860010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#860020000000
0!
0*
09
0>
0C
#860030000000
1!
1*
b101 6
19
1>
1C
b101 G
#860040000000
0!
0*
09
0>
0C
#860050000000
1!
1*
b110 6
19
1>
1C
b110 G
#860060000000
0!
0*
09
0>
0C
#860070000000
1!
1*
b111 6
19
1>
1C
b111 G
#860080000000
0!
0*
09
0>
0C
#860090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#860100000000
0!
0*
09
0>
0C
#860110000000
1!
1*
b1 6
19
1>
1C
b1 G
#860120000000
0!
0*
09
0>
0C
#860130000000
1!
1*
b10 6
19
1>
1C
b10 G
#860140000000
0!
0*
09
0>
0C
#860150000000
1!
1*
b11 6
19
1>
1C
b11 G
#860160000000
0!
0*
09
0>
0C
#860170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#860180000000
0!
0*
09
0>
0C
#860190000000
1!
1*
b101 6
19
1>
1C
b101 G
#860200000000
0!
0*
09
0>
0C
#860210000000
1!
1*
b110 6
19
1>
1C
b110 G
#860220000000
0!
0*
09
0>
0C
#860230000000
1!
1*
b111 6
19
1>
1C
b111 G
#860240000000
0!
1"
0*
1+
09
1:
0>
0C
#860250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#860260000000
0!
0*
09
0>
0C
#860270000000
1!
1*
b1 6
19
1>
1C
b1 G
#860280000000
0!
0*
09
0>
0C
#860290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#860300000000
0!
0*
09
0>
0C
#860310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#860320000000
0!
0*
09
0>
0C
#860330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#860340000000
0!
0*
09
0>
0C
#860350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#860360000000
0!
0#
0*
0,
09
0>
0?
0C
#860370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#860380000000
0!
0*
09
0>
0C
#860390000000
1!
1*
19
1>
1C
#860400000000
0!
0*
09
0>
0C
#860410000000
1!
1*
19
1>
1C
#860420000000
0!
0*
09
0>
0C
#860430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#860440000000
0!
0*
09
0>
0C
#860450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#860460000000
0!
0*
09
0>
0C
#860470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#860480000000
0!
0*
09
0>
0C
#860490000000
1!
1*
b10 6
19
1>
1C
b10 G
#860500000000
0!
0*
09
0>
0C
#860510000000
1!
1*
b11 6
19
1>
1C
b11 G
#860520000000
0!
0*
09
0>
0C
#860530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#860540000000
0!
0*
09
0>
0C
#860550000000
1!
1*
b101 6
19
1>
1C
b101 G
#860560000000
0!
0*
09
0>
0C
#860570000000
1!
1*
b110 6
19
1>
1C
b110 G
#860580000000
0!
0*
09
0>
0C
#860590000000
1!
1*
b111 6
19
1>
1C
b111 G
#860600000000
0!
0*
09
0>
0C
#860610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#860620000000
0!
0*
09
0>
0C
#860630000000
1!
1*
b1 6
19
1>
1C
b1 G
#860640000000
0!
0*
09
0>
0C
#860650000000
1!
1*
b10 6
19
1>
1C
b10 G
#860660000000
0!
0*
09
0>
0C
#860670000000
1!
1*
b11 6
19
1>
1C
b11 G
#860680000000
0!
0*
09
0>
0C
#860690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#860700000000
0!
0*
09
0>
0C
#860710000000
1!
1*
b101 6
19
1>
1C
b101 G
#860720000000
0!
0*
09
0>
0C
#860730000000
1!
1*
b110 6
19
1>
1C
b110 G
#860740000000
0!
0*
09
0>
0C
#860750000000
1!
1*
b111 6
19
1>
1C
b111 G
#860760000000
0!
0*
09
0>
0C
#860770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#860780000000
0!
0*
09
0>
0C
#860790000000
1!
1*
b1 6
19
1>
1C
b1 G
#860800000000
0!
0*
09
0>
0C
#860810000000
1!
1*
b10 6
19
1>
1C
b10 G
#860820000000
0!
0*
09
0>
0C
#860830000000
1!
1*
b11 6
19
1>
1C
b11 G
#860840000000
0!
0*
09
0>
0C
#860850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#860860000000
0!
0*
09
0>
0C
#860870000000
1!
1*
b101 6
19
1>
1C
b101 G
#860880000000
0!
0*
09
0>
0C
#860890000000
1!
1*
b110 6
19
1>
1C
b110 G
#860900000000
0!
0*
09
0>
0C
#860910000000
1!
1*
b111 6
19
1>
1C
b111 G
#860920000000
0!
1"
0*
1+
09
1:
0>
0C
#860930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#860940000000
0!
0*
09
0>
0C
#860950000000
1!
1*
b1 6
19
1>
1C
b1 G
#860960000000
0!
0*
09
0>
0C
#860970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#860980000000
0!
0*
09
0>
0C
#860990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#861000000000
0!
0*
09
0>
0C
#861010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#861020000000
0!
0*
09
0>
0C
#861030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#861040000000
0!
0#
0*
0,
09
0>
0?
0C
#861050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#861060000000
0!
0*
09
0>
0C
#861070000000
1!
1*
19
1>
1C
#861080000000
0!
0*
09
0>
0C
#861090000000
1!
1*
19
1>
1C
#861100000000
0!
0*
09
0>
0C
#861110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#861120000000
0!
0*
09
0>
0C
#861130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#861140000000
0!
0*
09
0>
0C
#861150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#861160000000
0!
0*
09
0>
0C
#861170000000
1!
1*
b10 6
19
1>
1C
b10 G
#861180000000
0!
0*
09
0>
0C
#861190000000
1!
1*
b11 6
19
1>
1C
b11 G
#861200000000
0!
0*
09
0>
0C
#861210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#861220000000
0!
0*
09
0>
0C
#861230000000
1!
1*
b101 6
19
1>
1C
b101 G
#861240000000
0!
0*
09
0>
0C
#861250000000
1!
1*
b110 6
19
1>
1C
b110 G
#861260000000
0!
0*
09
0>
0C
#861270000000
1!
1*
b111 6
19
1>
1C
b111 G
#861280000000
0!
0*
09
0>
0C
#861290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#861300000000
0!
0*
09
0>
0C
#861310000000
1!
1*
b1 6
19
1>
1C
b1 G
#861320000000
0!
0*
09
0>
0C
#861330000000
1!
1*
b10 6
19
1>
1C
b10 G
#861340000000
0!
0*
09
0>
0C
#861350000000
1!
1*
b11 6
19
1>
1C
b11 G
#861360000000
0!
0*
09
0>
0C
#861370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#861380000000
0!
0*
09
0>
0C
#861390000000
1!
1*
b101 6
19
1>
1C
b101 G
#861400000000
0!
0*
09
0>
0C
#861410000000
1!
1*
b110 6
19
1>
1C
b110 G
#861420000000
0!
0*
09
0>
0C
#861430000000
1!
1*
b111 6
19
1>
1C
b111 G
#861440000000
0!
0*
09
0>
0C
#861450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#861460000000
0!
0*
09
0>
0C
#861470000000
1!
1*
b1 6
19
1>
1C
b1 G
#861480000000
0!
0*
09
0>
0C
#861490000000
1!
1*
b10 6
19
1>
1C
b10 G
#861500000000
0!
0*
09
0>
0C
#861510000000
1!
1*
b11 6
19
1>
1C
b11 G
#861520000000
0!
0*
09
0>
0C
#861530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#861540000000
0!
0*
09
0>
0C
#861550000000
1!
1*
b101 6
19
1>
1C
b101 G
#861560000000
0!
0*
09
0>
0C
#861570000000
1!
1*
b110 6
19
1>
1C
b110 G
#861580000000
0!
0*
09
0>
0C
#861590000000
1!
1*
b111 6
19
1>
1C
b111 G
#861600000000
0!
1"
0*
1+
09
1:
0>
0C
#861610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#861620000000
0!
0*
09
0>
0C
#861630000000
1!
1*
b1 6
19
1>
1C
b1 G
#861640000000
0!
0*
09
0>
0C
#861650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#861660000000
0!
0*
09
0>
0C
#861670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#861680000000
0!
0*
09
0>
0C
#861690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#861700000000
0!
0*
09
0>
0C
#861710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#861720000000
0!
0#
0*
0,
09
0>
0?
0C
#861730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#861740000000
0!
0*
09
0>
0C
#861750000000
1!
1*
19
1>
1C
#861760000000
0!
0*
09
0>
0C
#861770000000
1!
1*
19
1>
1C
#861780000000
0!
0*
09
0>
0C
#861790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#861800000000
0!
0*
09
0>
0C
#861810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#861820000000
0!
0*
09
0>
0C
#861830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#861840000000
0!
0*
09
0>
0C
#861850000000
1!
1*
b10 6
19
1>
1C
b10 G
#861860000000
0!
0*
09
0>
0C
#861870000000
1!
1*
b11 6
19
1>
1C
b11 G
#861880000000
0!
0*
09
0>
0C
#861890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#861900000000
0!
0*
09
0>
0C
#861910000000
1!
1*
b101 6
19
1>
1C
b101 G
#861920000000
0!
0*
09
0>
0C
#861930000000
1!
1*
b110 6
19
1>
1C
b110 G
#861940000000
0!
0*
09
0>
0C
#861950000000
1!
1*
b111 6
19
1>
1C
b111 G
#861960000000
0!
0*
09
0>
0C
#861970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#861980000000
0!
0*
09
0>
0C
#861990000000
1!
1*
b1 6
19
1>
1C
b1 G
#862000000000
0!
0*
09
0>
0C
#862010000000
1!
1*
b10 6
19
1>
1C
b10 G
#862020000000
0!
0*
09
0>
0C
#862030000000
1!
1*
b11 6
19
1>
1C
b11 G
#862040000000
0!
0*
09
0>
0C
#862050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#862060000000
0!
0*
09
0>
0C
#862070000000
1!
1*
b101 6
19
1>
1C
b101 G
#862080000000
0!
0*
09
0>
0C
#862090000000
1!
1*
b110 6
19
1>
1C
b110 G
#862100000000
0!
0*
09
0>
0C
#862110000000
1!
1*
b111 6
19
1>
1C
b111 G
#862120000000
0!
0*
09
0>
0C
#862130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#862140000000
0!
0*
09
0>
0C
#862150000000
1!
1*
b1 6
19
1>
1C
b1 G
#862160000000
0!
0*
09
0>
0C
#862170000000
1!
1*
b10 6
19
1>
1C
b10 G
#862180000000
0!
0*
09
0>
0C
#862190000000
1!
1*
b11 6
19
1>
1C
b11 G
#862200000000
0!
0*
09
0>
0C
#862210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#862220000000
0!
0*
09
0>
0C
#862230000000
1!
1*
b101 6
19
1>
1C
b101 G
#862240000000
0!
0*
09
0>
0C
#862250000000
1!
1*
b110 6
19
1>
1C
b110 G
#862260000000
0!
0*
09
0>
0C
#862270000000
1!
1*
b111 6
19
1>
1C
b111 G
#862280000000
0!
1"
0*
1+
09
1:
0>
0C
#862290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#862300000000
0!
0*
09
0>
0C
#862310000000
1!
1*
b1 6
19
1>
1C
b1 G
#862320000000
0!
0*
09
0>
0C
#862330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#862340000000
0!
0*
09
0>
0C
#862350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#862360000000
0!
0*
09
0>
0C
#862370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#862380000000
0!
0*
09
0>
0C
#862390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#862400000000
0!
0#
0*
0,
09
0>
0?
0C
#862410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#862420000000
0!
0*
09
0>
0C
#862430000000
1!
1*
19
1>
1C
#862440000000
0!
0*
09
0>
0C
#862450000000
1!
1*
19
1>
1C
#862460000000
0!
0*
09
0>
0C
#862470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#862480000000
0!
0*
09
0>
0C
#862490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#862500000000
0!
0*
09
0>
0C
#862510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#862520000000
0!
0*
09
0>
0C
#862530000000
1!
1*
b10 6
19
1>
1C
b10 G
#862540000000
0!
0*
09
0>
0C
#862550000000
1!
1*
b11 6
19
1>
1C
b11 G
#862560000000
0!
0*
09
0>
0C
#862570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#862580000000
0!
0*
09
0>
0C
#862590000000
1!
1*
b101 6
19
1>
1C
b101 G
#862600000000
0!
0*
09
0>
0C
#862610000000
1!
1*
b110 6
19
1>
1C
b110 G
#862620000000
0!
0*
09
0>
0C
#862630000000
1!
1*
b111 6
19
1>
1C
b111 G
#862640000000
0!
0*
09
0>
0C
#862650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#862660000000
0!
0*
09
0>
0C
#862670000000
1!
1*
b1 6
19
1>
1C
b1 G
#862680000000
0!
0*
09
0>
0C
#862690000000
1!
1*
b10 6
19
1>
1C
b10 G
#862700000000
0!
0*
09
0>
0C
#862710000000
1!
1*
b11 6
19
1>
1C
b11 G
#862720000000
0!
0*
09
0>
0C
#862730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#862740000000
0!
0*
09
0>
0C
#862750000000
1!
1*
b101 6
19
1>
1C
b101 G
#862760000000
0!
0*
09
0>
0C
#862770000000
1!
1*
b110 6
19
1>
1C
b110 G
#862780000000
0!
0*
09
0>
0C
#862790000000
1!
1*
b111 6
19
1>
1C
b111 G
#862800000000
0!
0*
09
0>
0C
#862810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#862820000000
0!
0*
09
0>
0C
#862830000000
1!
1*
b1 6
19
1>
1C
b1 G
#862840000000
0!
0*
09
0>
0C
#862850000000
1!
1*
b10 6
19
1>
1C
b10 G
#862860000000
0!
0*
09
0>
0C
#862870000000
1!
1*
b11 6
19
1>
1C
b11 G
#862880000000
0!
0*
09
0>
0C
#862890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#862900000000
0!
0*
09
0>
0C
#862910000000
1!
1*
b101 6
19
1>
1C
b101 G
#862920000000
0!
0*
09
0>
0C
#862930000000
1!
1*
b110 6
19
1>
1C
b110 G
#862940000000
0!
0*
09
0>
0C
#862950000000
1!
1*
b111 6
19
1>
1C
b111 G
#862960000000
0!
1"
0*
1+
09
1:
0>
0C
#862970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#862980000000
0!
0*
09
0>
0C
#862990000000
1!
1*
b1 6
19
1>
1C
b1 G
#863000000000
0!
0*
09
0>
0C
#863010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#863020000000
0!
0*
09
0>
0C
#863030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#863040000000
0!
0*
09
0>
0C
#863050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#863060000000
0!
0*
09
0>
0C
#863070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#863080000000
0!
0#
0*
0,
09
0>
0?
0C
#863090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#863100000000
0!
0*
09
0>
0C
#863110000000
1!
1*
19
1>
1C
#863120000000
0!
0*
09
0>
0C
#863130000000
1!
1*
19
1>
1C
#863140000000
0!
0*
09
0>
0C
#863150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#863160000000
0!
0*
09
0>
0C
#863170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#863180000000
0!
0*
09
0>
0C
#863190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#863200000000
0!
0*
09
0>
0C
#863210000000
1!
1*
b10 6
19
1>
1C
b10 G
#863220000000
0!
0*
09
0>
0C
#863230000000
1!
1*
b11 6
19
1>
1C
b11 G
#863240000000
0!
0*
09
0>
0C
#863250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#863260000000
0!
0*
09
0>
0C
#863270000000
1!
1*
b101 6
19
1>
1C
b101 G
#863280000000
0!
0*
09
0>
0C
#863290000000
1!
1*
b110 6
19
1>
1C
b110 G
#863300000000
0!
0*
09
0>
0C
#863310000000
1!
1*
b111 6
19
1>
1C
b111 G
#863320000000
0!
0*
09
0>
0C
#863330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#863340000000
0!
0*
09
0>
0C
#863350000000
1!
1*
b1 6
19
1>
1C
b1 G
#863360000000
0!
0*
09
0>
0C
#863370000000
1!
1*
b10 6
19
1>
1C
b10 G
#863380000000
0!
0*
09
0>
0C
#863390000000
1!
1*
b11 6
19
1>
1C
b11 G
#863400000000
0!
0*
09
0>
0C
#863410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#863420000000
0!
0*
09
0>
0C
#863430000000
1!
1*
b101 6
19
1>
1C
b101 G
#863440000000
0!
0*
09
0>
0C
#863450000000
1!
1*
b110 6
19
1>
1C
b110 G
#863460000000
0!
0*
09
0>
0C
#863470000000
1!
1*
b111 6
19
1>
1C
b111 G
#863480000000
0!
0*
09
0>
0C
#863490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#863500000000
0!
0*
09
0>
0C
#863510000000
1!
1*
b1 6
19
1>
1C
b1 G
#863520000000
0!
0*
09
0>
0C
#863530000000
1!
1*
b10 6
19
1>
1C
b10 G
#863540000000
0!
0*
09
0>
0C
#863550000000
1!
1*
b11 6
19
1>
1C
b11 G
#863560000000
0!
0*
09
0>
0C
#863570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#863580000000
0!
0*
09
0>
0C
#863590000000
1!
1*
b101 6
19
1>
1C
b101 G
#863600000000
0!
0*
09
0>
0C
#863610000000
1!
1*
b110 6
19
1>
1C
b110 G
#863620000000
0!
0*
09
0>
0C
#863630000000
1!
1*
b111 6
19
1>
1C
b111 G
#863640000000
0!
1"
0*
1+
09
1:
0>
0C
#863650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#863660000000
0!
0*
09
0>
0C
#863670000000
1!
1*
b1 6
19
1>
1C
b1 G
#863680000000
0!
0*
09
0>
0C
#863690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#863700000000
0!
0*
09
0>
0C
#863710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#863720000000
0!
0*
09
0>
0C
#863730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#863740000000
0!
0*
09
0>
0C
#863750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#863760000000
0!
0#
0*
0,
09
0>
0?
0C
#863770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#863780000000
0!
0*
09
0>
0C
#863790000000
1!
1*
19
1>
1C
#863800000000
0!
0*
09
0>
0C
#863810000000
1!
1*
19
1>
1C
#863820000000
0!
0*
09
0>
0C
#863830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#863840000000
0!
0*
09
0>
0C
#863850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#863860000000
0!
0*
09
0>
0C
#863870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#863880000000
0!
0*
09
0>
0C
#863890000000
1!
1*
b10 6
19
1>
1C
b10 G
#863900000000
0!
0*
09
0>
0C
#863910000000
1!
1*
b11 6
19
1>
1C
b11 G
#863920000000
0!
0*
09
0>
0C
#863930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#863940000000
0!
0*
09
0>
0C
#863950000000
1!
1*
b101 6
19
1>
1C
b101 G
#863960000000
0!
0*
09
0>
0C
#863970000000
1!
1*
b110 6
19
1>
1C
b110 G
#863980000000
0!
0*
09
0>
0C
#863990000000
1!
1*
b111 6
19
1>
1C
b111 G
#864000000000
0!
0*
09
0>
0C
#864010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#864020000000
0!
0*
09
0>
0C
#864030000000
1!
1*
b1 6
19
1>
1C
b1 G
#864040000000
0!
0*
09
0>
0C
#864050000000
1!
1*
b10 6
19
1>
1C
b10 G
#864060000000
0!
0*
09
0>
0C
#864070000000
1!
1*
b11 6
19
1>
1C
b11 G
#864080000000
0!
0*
09
0>
0C
#864090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#864100000000
0!
0*
09
0>
0C
#864110000000
1!
1*
b101 6
19
1>
1C
b101 G
#864120000000
0!
0*
09
0>
0C
#864130000000
1!
1*
b110 6
19
1>
1C
b110 G
#864140000000
0!
0*
09
0>
0C
#864150000000
1!
1*
b111 6
19
1>
1C
b111 G
#864160000000
0!
0*
09
0>
0C
#864170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#864180000000
0!
0*
09
0>
0C
#864190000000
1!
1*
b1 6
19
1>
1C
b1 G
#864200000000
0!
0*
09
0>
0C
#864210000000
1!
1*
b10 6
19
1>
1C
b10 G
#864220000000
0!
0*
09
0>
0C
#864230000000
1!
1*
b11 6
19
1>
1C
b11 G
#864240000000
0!
0*
09
0>
0C
#864250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#864260000000
0!
0*
09
0>
0C
#864270000000
1!
1*
b101 6
19
1>
1C
b101 G
#864280000000
0!
0*
09
0>
0C
#864290000000
1!
1*
b110 6
19
1>
1C
b110 G
#864300000000
0!
0*
09
0>
0C
#864310000000
1!
1*
b111 6
19
1>
1C
b111 G
#864320000000
0!
1"
0*
1+
09
1:
0>
0C
#864330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#864340000000
0!
0*
09
0>
0C
#864350000000
1!
1*
b1 6
19
1>
1C
b1 G
#864360000000
0!
0*
09
0>
0C
#864370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#864380000000
0!
0*
09
0>
0C
#864390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#864400000000
0!
0*
09
0>
0C
#864410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#864420000000
0!
0*
09
0>
0C
#864430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#864440000000
0!
0#
0*
0,
09
0>
0?
0C
#864450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#864460000000
0!
0*
09
0>
0C
#864470000000
1!
1*
19
1>
1C
#864480000000
0!
0*
09
0>
0C
#864490000000
1!
1*
19
1>
1C
#864500000000
0!
0*
09
0>
0C
#864510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#864520000000
0!
0*
09
0>
0C
#864530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#864540000000
0!
0*
09
0>
0C
#864550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#864560000000
0!
0*
09
0>
0C
#864570000000
1!
1*
b10 6
19
1>
1C
b10 G
#864580000000
0!
0*
09
0>
0C
#864590000000
1!
1*
b11 6
19
1>
1C
b11 G
#864600000000
0!
0*
09
0>
0C
#864610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#864620000000
0!
0*
09
0>
0C
#864630000000
1!
1*
b101 6
19
1>
1C
b101 G
#864640000000
0!
0*
09
0>
0C
#864650000000
1!
1*
b110 6
19
1>
1C
b110 G
#864660000000
0!
0*
09
0>
0C
#864670000000
1!
1*
b111 6
19
1>
1C
b111 G
#864680000000
0!
0*
09
0>
0C
#864690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#864700000000
0!
0*
09
0>
0C
#864710000000
1!
1*
b1 6
19
1>
1C
b1 G
#864720000000
0!
0*
09
0>
0C
#864730000000
1!
1*
b10 6
19
1>
1C
b10 G
#864740000000
0!
0*
09
0>
0C
#864750000000
1!
1*
b11 6
19
1>
1C
b11 G
#864760000000
0!
0*
09
0>
0C
#864770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#864780000000
0!
0*
09
0>
0C
#864790000000
1!
1*
b101 6
19
1>
1C
b101 G
#864800000000
0!
0*
09
0>
0C
#864810000000
1!
1*
b110 6
19
1>
1C
b110 G
#864820000000
0!
0*
09
0>
0C
#864830000000
1!
1*
b111 6
19
1>
1C
b111 G
#864840000000
0!
0*
09
0>
0C
#864850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#864860000000
0!
0*
09
0>
0C
#864870000000
1!
1*
b1 6
19
1>
1C
b1 G
#864880000000
0!
0*
09
0>
0C
#864890000000
1!
1*
b10 6
19
1>
1C
b10 G
#864900000000
0!
0*
09
0>
0C
#864910000000
1!
1*
b11 6
19
1>
1C
b11 G
#864920000000
0!
0*
09
0>
0C
#864930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#864940000000
0!
0*
09
0>
0C
#864950000000
1!
1*
b101 6
19
1>
1C
b101 G
#864960000000
0!
0*
09
0>
0C
#864970000000
1!
1*
b110 6
19
1>
1C
b110 G
#864980000000
0!
0*
09
0>
0C
#864990000000
1!
1*
b111 6
19
1>
1C
b111 G
#865000000000
0!
1"
0*
1+
09
1:
0>
0C
#865010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#865020000000
0!
0*
09
0>
0C
#865030000000
1!
1*
b1 6
19
1>
1C
b1 G
#865040000000
0!
0*
09
0>
0C
#865050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#865060000000
0!
0*
09
0>
0C
#865070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#865080000000
0!
0*
09
0>
0C
#865090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#865100000000
0!
0*
09
0>
0C
#865110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#865120000000
0!
0#
0*
0,
09
0>
0?
0C
#865130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#865140000000
0!
0*
09
0>
0C
#865150000000
1!
1*
19
1>
1C
#865160000000
0!
0*
09
0>
0C
#865170000000
1!
1*
19
1>
1C
#865180000000
0!
0*
09
0>
0C
#865190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#865200000000
0!
0*
09
0>
0C
#865210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#865220000000
0!
0*
09
0>
0C
#865230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#865240000000
0!
0*
09
0>
0C
#865250000000
1!
1*
b10 6
19
1>
1C
b10 G
#865260000000
0!
0*
09
0>
0C
#865270000000
1!
1*
b11 6
19
1>
1C
b11 G
#865280000000
0!
0*
09
0>
0C
#865290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#865300000000
0!
0*
09
0>
0C
#865310000000
1!
1*
b101 6
19
1>
1C
b101 G
#865320000000
0!
0*
09
0>
0C
#865330000000
1!
1*
b110 6
19
1>
1C
b110 G
#865340000000
0!
0*
09
0>
0C
#865350000000
1!
1*
b111 6
19
1>
1C
b111 G
#865360000000
0!
0*
09
0>
0C
#865370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#865380000000
0!
0*
09
0>
0C
#865390000000
1!
1*
b1 6
19
1>
1C
b1 G
#865400000000
0!
0*
09
0>
0C
#865410000000
1!
1*
b10 6
19
1>
1C
b10 G
#865420000000
0!
0*
09
0>
0C
#865430000000
1!
1*
b11 6
19
1>
1C
b11 G
#865440000000
0!
0*
09
0>
0C
#865450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#865460000000
0!
0*
09
0>
0C
#865470000000
1!
1*
b101 6
19
1>
1C
b101 G
#865480000000
0!
0*
09
0>
0C
#865490000000
1!
1*
b110 6
19
1>
1C
b110 G
#865500000000
0!
0*
09
0>
0C
#865510000000
1!
1*
b111 6
19
1>
1C
b111 G
#865520000000
0!
0*
09
0>
0C
#865530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#865540000000
0!
0*
09
0>
0C
#865550000000
1!
1*
b1 6
19
1>
1C
b1 G
#865560000000
0!
0*
09
0>
0C
#865570000000
1!
1*
b10 6
19
1>
1C
b10 G
#865580000000
0!
0*
09
0>
0C
#865590000000
1!
1*
b11 6
19
1>
1C
b11 G
#865600000000
0!
0*
09
0>
0C
#865610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#865620000000
0!
0*
09
0>
0C
#865630000000
1!
1*
b101 6
19
1>
1C
b101 G
#865640000000
0!
0*
09
0>
0C
#865650000000
1!
1*
b110 6
19
1>
1C
b110 G
#865660000000
0!
0*
09
0>
0C
#865670000000
1!
1*
b111 6
19
1>
1C
b111 G
#865680000000
0!
1"
0*
1+
09
1:
0>
0C
#865690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#865700000000
0!
0*
09
0>
0C
#865710000000
1!
1*
b1 6
19
1>
1C
b1 G
#865720000000
0!
0*
09
0>
0C
#865730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#865740000000
0!
0*
09
0>
0C
#865750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#865760000000
0!
0*
09
0>
0C
#865770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#865780000000
0!
0*
09
0>
0C
#865790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#865800000000
0!
0#
0*
0,
09
0>
0?
0C
#865810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#865820000000
0!
0*
09
0>
0C
#865830000000
1!
1*
19
1>
1C
#865840000000
0!
0*
09
0>
0C
#865850000000
1!
1*
19
1>
1C
#865860000000
0!
0*
09
0>
0C
#865870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#865880000000
0!
0*
09
0>
0C
#865890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#865900000000
0!
0*
09
0>
0C
#865910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#865920000000
0!
0*
09
0>
0C
#865930000000
1!
1*
b10 6
19
1>
1C
b10 G
#865940000000
0!
0*
09
0>
0C
#865950000000
1!
1*
b11 6
19
1>
1C
b11 G
#865960000000
0!
0*
09
0>
0C
#865970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#865980000000
0!
0*
09
0>
0C
#865990000000
1!
1*
b101 6
19
1>
1C
b101 G
#866000000000
0!
0*
09
0>
0C
#866010000000
1!
1*
b110 6
19
1>
1C
b110 G
#866020000000
0!
0*
09
0>
0C
#866030000000
1!
1*
b111 6
19
1>
1C
b111 G
#866040000000
0!
0*
09
0>
0C
#866050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#866060000000
0!
0*
09
0>
0C
#866070000000
1!
1*
b1 6
19
1>
1C
b1 G
#866080000000
0!
0*
09
0>
0C
#866090000000
1!
1*
b10 6
19
1>
1C
b10 G
#866100000000
0!
0*
09
0>
0C
#866110000000
1!
1*
b11 6
19
1>
1C
b11 G
#866120000000
0!
0*
09
0>
0C
#866130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#866140000000
0!
0*
09
0>
0C
#866150000000
1!
1*
b101 6
19
1>
1C
b101 G
#866160000000
0!
0*
09
0>
0C
#866170000000
1!
1*
b110 6
19
1>
1C
b110 G
#866180000000
0!
0*
09
0>
0C
#866190000000
1!
1*
b111 6
19
1>
1C
b111 G
#866200000000
0!
0*
09
0>
0C
#866210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#866220000000
0!
0*
09
0>
0C
#866230000000
1!
1*
b1 6
19
1>
1C
b1 G
#866240000000
0!
0*
09
0>
0C
#866250000000
1!
1*
b10 6
19
1>
1C
b10 G
#866260000000
0!
0*
09
0>
0C
#866270000000
1!
1*
b11 6
19
1>
1C
b11 G
#866280000000
0!
0*
09
0>
0C
#866290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#866300000000
0!
0*
09
0>
0C
#866310000000
1!
1*
b101 6
19
1>
1C
b101 G
#866320000000
0!
0*
09
0>
0C
#866330000000
1!
1*
b110 6
19
1>
1C
b110 G
#866340000000
0!
0*
09
0>
0C
#866350000000
1!
1*
b111 6
19
1>
1C
b111 G
#866360000000
0!
1"
0*
1+
09
1:
0>
0C
#866370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#866380000000
0!
0*
09
0>
0C
#866390000000
1!
1*
b1 6
19
1>
1C
b1 G
#866400000000
0!
0*
09
0>
0C
#866410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#866420000000
0!
0*
09
0>
0C
#866430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#866440000000
0!
0*
09
0>
0C
#866450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#866460000000
0!
0*
09
0>
0C
#866470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#866480000000
0!
0#
0*
0,
09
0>
0?
0C
#866490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#866500000000
0!
0*
09
0>
0C
#866510000000
1!
1*
19
1>
1C
#866520000000
0!
0*
09
0>
0C
#866530000000
1!
1*
19
1>
1C
#866540000000
0!
0*
09
0>
0C
#866550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#866560000000
0!
0*
09
0>
0C
#866570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#866580000000
0!
0*
09
0>
0C
#866590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#866600000000
0!
0*
09
0>
0C
#866610000000
1!
1*
b10 6
19
1>
1C
b10 G
#866620000000
0!
0*
09
0>
0C
#866630000000
1!
1*
b11 6
19
1>
1C
b11 G
#866640000000
0!
0*
09
0>
0C
#866650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#866660000000
0!
0*
09
0>
0C
#866670000000
1!
1*
b101 6
19
1>
1C
b101 G
#866680000000
0!
0*
09
0>
0C
#866690000000
1!
1*
b110 6
19
1>
1C
b110 G
#866700000000
0!
0*
09
0>
0C
#866710000000
1!
1*
b111 6
19
1>
1C
b111 G
#866720000000
0!
0*
09
0>
0C
#866730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#866740000000
0!
0*
09
0>
0C
#866750000000
1!
1*
b1 6
19
1>
1C
b1 G
#866760000000
0!
0*
09
0>
0C
#866770000000
1!
1*
b10 6
19
1>
1C
b10 G
#866780000000
0!
0*
09
0>
0C
#866790000000
1!
1*
b11 6
19
1>
1C
b11 G
#866800000000
0!
0*
09
0>
0C
#866810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#866820000000
0!
0*
09
0>
0C
#866830000000
1!
1*
b101 6
19
1>
1C
b101 G
#866840000000
0!
0*
09
0>
0C
#866850000000
1!
1*
b110 6
19
1>
1C
b110 G
#866860000000
0!
0*
09
0>
0C
#866870000000
1!
1*
b111 6
19
1>
1C
b111 G
#866880000000
0!
0*
09
0>
0C
#866890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#866900000000
0!
0*
09
0>
0C
#866910000000
1!
1*
b1 6
19
1>
1C
b1 G
#866920000000
0!
0*
09
0>
0C
#866930000000
1!
1*
b10 6
19
1>
1C
b10 G
#866940000000
0!
0*
09
0>
0C
#866950000000
1!
1*
b11 6
19
1>
1C
b11 G
#866960000000
0!
0*
09
0>
0C
#866970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#866980000000
0!
0*
09
0>
0C
#866990000000
1!
1*
b101 6
19
1>
1C
b101 G
#867000000000
0!
0*
09
0>
0C
#867010000000
1!
1*
b110 6
19
1>
1C
b110 G
#867020000000
0!
0*
09
0>
0C
#867030000000
1!
1*
b111 6
19
1>
1C
b111 G
#867040000000
0!
1"
0*
1+
09
1:
0>
0C
#867050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#867060000000
0!
0*
09
0>
0C
#867070000000
1!
1*
b1 6
19
1>
1C
b1 G
#867080000000
0!
0*
09
0>
0C
#867090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#867100000000
0!
0*
09
0>
0C
#867110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#867120000000
0!
0*
09
0>
0C
#867130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#867140000000
0!
0*
09
0>
0C
#867150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#867160000000
0!
0#
0*
0,
09
0>
0?
0C
#867170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#867180000000
0!
0*
09
0>
0C
#867190000000
1!
1*
19
1>
1C
#867200000000
0!
0*
09
0>
0C
#867210000000
1!
1*
19
1>
1C
#867220000000
0!
0*
09
0>
0C
#867230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#867240000000
0!
0*
09
0>
0C
#867250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#867260000000
0!
0*
09
0>
0C
#867270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#867280000000
0!
0*
09
0>
0C
#867290000000
1!
1*
b10 6
19
1>
1C
b10 G
#867300000000
0!
0*
09
0>
0C
#867310000000
1!
1*
b11 6
19
1>
1C
b11 G
#867320000000
0!
0*
09
0>
0C
#867330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#867340000000
0!
0*
09
0>
0C
#867350000000
1!
1*
b101 6
19
1>
1C
b101 G
#867360000000
0!
0*
09
0>
0C
#867370000000
1!
1*
b110 6
19
1>
1C
b110 G
#867380000000
0!
0*
09
0>
0C
#867390000000
1!
1*
b111 6
19
1>
1C
b111 G
#867400000000
0!
0*
09
0>
0C
#867410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#867420000000
0!
0*
09
0>
0C
#867430000000
1!
1*
b1 6
19
1>
1C
b1 G
#867440000000
0!
0*
09
0>
0C
#867450000000
1!
1*
b10 6
19
1>
1C
b10 G
#867460000000
0!
0*
09
0>
0C
#867470000000
1!
1*
b11 6
19
1>
1C
b11 G
#867480000000
0!
0*
09
0>
0C
#867490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#867500000000
0!
0*
09
0>
0C
#867510000000
1!
1*
b101 6
19
1>
1C
b101 G
#867520000000
0!
0*
09
0>
0C
#867530000000
1!
1*
b110 6
19
1>
1C
b110 G
#867540000000
0!
0*
09
0>
0C
#867550000000
1!
1*
b111 6
19
1>
1C
b111 G
#867560000000
0!
0*
09
0>
0C
#867570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#867580000000
0!
0*
09
0>
0C
#867590000000
1!
1*
b1 6
19
1>
1C
b1 G
#867600000000
0!
0*
09
0>
0C
#867610000000
1!
1*
b10 6
19
1>
1C
b10 G
#867620000000
0!
0*
09
0>
0C
#867630000000
1!
1*
b11 6
19
1>
1C
b11 G
#867640000000
0!
0*
09
0>
0C
#867650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#867660000000
0!
0*
09
0>
0C
#867670000000
1!
1*
b101 6
19
1>
1C
b101 G
#867680000000
0!
0*
09
0>
0C
#867690000000
1!
1*
b110 6
19
1>
1C
b110 G
#867700000000
0!
0*
09
0>
0C
#867710000000
1!
1*
b111 6
19
1>
1C
b111 G
#867720000000
0!
1"
0*
1+
09
1:
0>
0C
#867730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#867740000000
0!
0*
09
0>
0C
#867750000000
1!
1*
b1 6
19
1>
1C
b1 G
#867760000000
0!
0*
09
0>
0C
#867770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#867780000000
0!
0*
09
0>
0C
#867790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#867800000000
0!
0*
09
0>
0C
#867810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#867820000000
0!
0*
09
0>
0C
#867830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#867840000000
0!
0#
0*
0,
09
0>
0?
0C
#867850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#867860000000
0!
0*
09
0>
0C
#867870000000
1!
1*
19
1>
1C
#867880000000
0!
0*
09
0>
0C
#867890000000
1!
1*
19
1>
1C
#867900000000
0!
0*
09
0>
0C
#867910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#867920000000
0!
0*
09
0>
0C
#867930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#867940000000
0!
0*
09
0>
0C
#867950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#867960000000
0!
0*
09
0>
0C
#867970000000
1!
1*
b10 6
19
1>
1C
b10 G
#867980000000
0!
0*
09
0>
0C
#867990000000
1!
1*
b11 6
19
1>
1C
b11 G
#868000000000
0!
0*
09
0>
0C
#868010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#868020000000
0!
0*
09
0>
0C
#868030000000
1!
1*
b101 6
19
1>
1C
b101 G
#868040000000
0!
0*
09
0>
0C
#868050000000
1!
1*
b110 6
19
1>
1C
b110 G
#868060000000
0!
0*
09
0>
0C
#868070000000
1!
1*
b111 6
19
1>
1C
b111 G
#868080000000
0!
0*
09
0>
0C
#868090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#868100000000
0!
0*
09
0>
0C
#868110000000
1!
1*
b1 6
19
1>
1C
b1 G
#868120000000
0!
0*
09
0>
0C
#868130000000
1!
1*
b10 6
19
1>
1C
b10 G
#868140000000
0!
0*
09
0>
0C
#868150000000
1!
1*
b11 6
19
1>
1C
b11 G
#868160000000
0!
0*
09
0>
0C
#868170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#868180000000
0!
0*
09
0>
0C
#868190000000
1!
1*
b101 6
19
1>
1C
b101 G
#868200000000
0!
0*
09
0>
0C
#868210000000
1!
1*
b110 6
19
1>
1C
b110 G
#868220000000
0!
0*
09
0>
0C
#868230000000
1!
1*
b111 6
19
1>
1C
b111 G
#868240000000
0!
0*
09
0>
0C
#868250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#868260000000
0!
0*
09
0>
0C
#868270000000
1!
1*
b1 6
19
1>
1C
b1 G
#868280000000
0!
0*
09
0>
0C
#868290000000
1!
1*
b10 6
19
1>
1C
b10 G
#868300000000
0!
0*
09
0>
0C
#868310000000
1!
1*
b11 6
19
1>
1C
b11 G
#868320000000
0!
0*
09
0>
0C
#868330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#868340000000
0!
0*
09
0>
0C
#868350000000
1!
1*
b101 6
19
1>
1C
b101 G
#868360000000
0!
0*
09
0>
0C
#868370000000
1!
1*
b110 6
19
1>
1C
b110 G
#868380000000
0!
0*
09
0>
0C
#868390000000
1!
1*
b111 6
19
1>
1C
b111 G
#868400000000
0!
1"
0*
1+
09
1:
0>
0C
#868410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#868420000000
0!
0*
09
0>
0C
#868430000000
1!
1*
b1 6
19
1>
1C
b1 G
#868440000000
0!
0*
09
0>
0C
#868450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#868460000000
0!
0*
09
0>
0C
#868470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#868480000000
0!
0*
09
0>
0C
#868490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#868500000000
0!
0*
09
0>
0C
#868510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#868520000000
0!
0#
0*
0,
09
0>
0?
0C
#868530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#868540000000
0!
0*
09
0>
0C
#868550000000
1!
1*
19
1>
1C
#868560000000
0!
0*
09
0>
0C
#868570000000
1!
1*
19
1>
1C
#868580000000
0!
0*
09
0>
0C
#868590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#868600000000
0!
0*
09
0>
0C
#868610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#868620000000
0!
0*
09
0>
0C
#868630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#868640000000
0!
0*
09
0>
0C
#868650000000
1!
1*
b10 6
19
1>
1C
b10 G
#868660000000
0!
0*
09
0>
0C
#868670000000
1!
1*
b11 6
19
1>
1C
b11 G
#868680000000
0!
0*
09
0>
0C
#868690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#868700000000
0!
0*
09
0>
0C
#868710000000
1!
1*
b101 6
19
1>
1C
b101 G
#868720000000
0!
0*
09
0>
0C
#868730000000
1!
1*
b110 6
19
1>
1C
b110 G
#868740000000
0!
0*
09
0>
0C
#868750000000
1!
1*
b111 6
19
1>
1C
b111 G
#868760000000
0!
0*
09
0>
0C
#868770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#868780000000
0!
0*
09
0>
0C
#868790000000
1!
1*
b1 6
19
1>
1C
b1 G
#868800000000
0!
0*
09
0>
0C
#868810000000
1!
1*
b10 6
19
1>
1C
b10 G
#868820000000
0!
0*
09
0>
0C
#868830000000
1!
1*
b11 6
19
1>
1C
b11 G
#868840000000
0!
0*
09
0>
0C
#868850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#868860000000
0!
0*
09
0>
0C
#868870000000
1!
1*
b101 6
19
1>
1C
b101 G
#868880000000
0!
0*
09
0>
0C
#868890000000
1!
1*
b110 6
19
1>
1C
b110 G
#868900000000
0!
0*
09
0>
0C
#868910000000
1!
1*
b111 6
19
1>
1C
b111 G
#868920000000
0!
0*
09
0>
0C
#868930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#868940000000
0!
0*
09
0>
0C
#868950000000
1!
1*
b1 6
19
1>
1C
b1 G
#868960000000
0!
0*
09
0>
0C
#868970000000
1!
1*
b10 6
19
1>
1C
b10 G
#868980000000
0!
0*
09
0>
0C
#868990000000
1!
1*
b11 6
19
1>
1C
b11 G
#869000000000
0!
0*
09
0>
0C
#869010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#869020000000
0!
0*
09
0>
0C
#869030000000
1!
1*
b101 6
19
1>
1C
b101 G
#869040000000
0!
0*
09
0>
0C
#869050000000
1!
1*
b110 6
19
1>
1C
b110 G
#869060000000
0!
0*
09
0>
0C
#869070000000
1!
1*
b111 6
19
1>
1C
b111 G
#869080000000
0!
1"
0*
1+
09
1:
0>
0C
#869090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#869100000000
0!
0*
09
0>
0C
#869110000000
1!
1*
b1 6
19
1>
1C
b1 G
#869120000000
0!
0*
09
0>
0C
#869130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#869140000000
0!
0*
09
0>
0C
#869150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#869160000000
0!
0*
09
0>
0C
#869170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#869180000000
0!
0*
09
0>
0C
#869190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#869200000000
0!
0#
0*
0,
09
0>
0?
0C
#869210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#869220000000
0!
0*
09
0>
0C
#869230000000
1!
1*
19
1>
1C
#869240000000
0!
0*
09
0>
0C
#869250000000
1!
1*
19
1>
1C
#869260000000
0!
0*
09
0>
0C
#869270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#869280000000
0!
0*
09
0>
0C
#869290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#869300000000
0!
0*
09
0>
0C
#869310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#869320000000
0!
0*
09
0>
0C
#869330000000
1!
1*
b10 6
19
1>
1C
b10 G
#869340000000
0!
0*
09
0>
0C
#869350000000
1!
1*
b11 6
19
1>
1C
b11 G
#869360000000
0!
0*
09
0>
0C
#869370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#869380000000
0!
0*
09
0>
0C
#869390000000
1!
1*
b101 6
19
1>
1C
b101 G
#869400000000
0!
0*
09
0>
0C
#869410000000
1!
1*
b110 6
19
1>
1C
b110 G
#869420000000
0!
0*
09
0>
0C
#869430000000
1!
1*
b111 6
19
1>
1C
b111 G
#869440000000
0!
0*
09
0>
0C
#869450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#869460000000
0!
0*
09
0>
0C
#869470000000
1!
1*
b1 6
19
1>
1C
b1 G
#869480000000
0!
0*
09
0>
0C
#869490000000
1!
1*
b10 6
19
1>
1C
b10 G
#869500000000
0!
0*
09
0>
0C
#869510000000
1!
1*
b11 6
19
1>
1C
b11 G
#869520000000
0!
0*
09
0>
0C
#869530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#869540000000
0!
0*
09
0>
0C
#869550000000
1!
1*
b101 6
19
1>
1C
b101 G
#869560000000
0!
0*
09
0>
0C
#869570000000
1!
1*
b110 6
19
1>
1C
b110 G
#869580000000
0!
0*
09
0>
0C
#869590000000
1!
1*
b111 6
19
1>
1C
b111 G
#869600000000
0!
0*
09
0>
0C
#869610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#869620000000
0!
0*
09
0>
0C
#869630000000
1!
1*
b1 6
19
1>
1C
b1 G
#869640000000
0!
0*
09
0>
0C
#869650000000
1!
1*
b10 6
19
1>
1C
b10 G
#869660000000
0!
0*
09
0>
0C
#869670000000
1!
1*
b11 6
19
1>
1C
b11 G
#869680000000
0!
0*
09
0>
0C
#869690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#869700000000
0!
0*
09
0>
0C
#869710000000
1!
1*
b101 6
19
1>
1C
b101 G
#869720000000
0!
0*
09
0>
0C
#869730000000
1!
1*
b110 6
19
1>
1C
b110 G
#869740000000
0!
0*
09
0>
0C
#869750000000
1!
1*
b111 6
19
1>
1C
b111 G
#869760000000
0!
1"
0*
1+
09
1:
0>
0C
#869770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#869780000000
0!
0*
09
0>
0C
#869790000000
1!
1*
b1 6
19
1>
1C
b1 G
#869800000000
0!
0*
09
0>
0C
#869810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#869820000000
0!
0*
09
0>
0C
#869830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#869840000000
0!
0*
09
0>
0C
#869850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#869860000000
0!
0*
09
0>
0C
#869870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#869880000000
0!
0#
0*
0,
09
0>
0?
0C
#869890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#869900000000
0!
0*
09
0>
0C
#869910000000
1!
1*
19
1>
1C
#869920000000
0!
0*
09
0>
0C
#869930000000
1!
1*
19
1>
1C
#869940000000
0!
0*
09
0>
0C
#869950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#869960000000
0!
0*
09
0>
0C
#869970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#869980000000
0!
0*
09
0>
0C
#869990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#870000000000
0!
0*
09
0>
0C
#870010000000
1!
1*
b10 6
19
1>
1C
b10 G
#870020000000
0!
0*
09
0>
0C
#870030000000
1!
1*
b11 6
19
1>
1C
b11 G
#870040000000
0!
0*
09
0>
0C
#870050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#870060000000
0!
0*
09
0>
0C
#870070000000
1!
1*
b101 6
19
1>
1C
b101 G
#870080000000
0!
0*
09
0>
0C
#870090000000
1!
1*
b110 6
19
1>
1C
b110 G
#870100000000
0!
0*
09
0>
0C
#870110000000
1!
1*
b111 6
19
1>
1C
b111 G
#870120000000
0!
0*
09
0>
0C
#870130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#870140000000
0!
0*
09
0>
0C
#870150000000
1!
1*
b1 6
19
1>
1C
b1 G
#870160000000
0!
0*
09
0>
0C
#870170000000
1!
1*
b10 6
19
1>
1C
b10 G
#870180000000
0!
0*
09
0>
0C
#870190000000
1!
1*
b11 6
19
1>
1C
b11 G
#870200000000
0!
0*
09
0>
0C
#870210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#870220000000
0!
0*
09
0>
0C
#870230000000
1!
1*
b101 6
19
1>
1C
b101 G
#870240000000
0!
0*
09
0>
0C
#870250000000
1!
1*
b110 6
19
1>
1C
b110 G
#870260000000
0!
0*
09
0>
0C
#870270000000
1!
1*
b111 6
19
1>
1C
b111 G
#870280000000
0!
0*
09
0>
0C
#870290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#870300000000
0!
0*
09
0>
0C
#870310000000
1!
1*
b1 6
19
1>
1C
b1 G
#870320000000
0!
0*
09
0>
0C
#870330000000
1!
1*
b10 6
19
1>
1C
b10 G
#870340000000
0!
0*
09
0>
0C
#870350000000
1!
1*
b11 6
19
1>
1C
b11 G
#870360000000
0!
0*
09
0>
0C
#870370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#870380000000
0!
0*
09
0>
0C
#870390000000
1!
1*
b101 6
19
1>
1C
b101 G
#870400000000
0!
0*
09
0>
0C
#870410000000
1!
1*
b110 6
19
1>
1C
b110 G
#870420000000
0!
0*
09
0>
0C
#870430000000
1!
1*
b111 6
19
1>
1C
b111 G
#870440000000
0!
1"
0*
1+
09
1:
0>
0C
#870450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#870460000000
0!
0*
09
0>
0C
#870470000000
1!
1*
b1 6
19
1>
1C
b1 G
#870480000000
0!
0*
09
0>
0C
#870490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#870500000000
0!
0*
09
0>
0C
#870510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#870520000000
0!
0*
09
0>
0C
#870530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#870540000000
0!
0*
09
0>
0C
#870550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#870560000000
0!
0#
0*
0,
09
0>
0?
0C
#870570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#870580000000
0!
0*
09
0>
0C
#870590000000
1!
1*
19
1>
1C
#870600000000
0!
0*
09
0>
0C
#870610000000
1!
1*
19
1>
1C
#870620000000
0!
0*
09
0>
0C
#870630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#870640000000
0!
0*
09
0>
0C
#870650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#870660000000
0!
0*
09
0>
0C
#870670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#870680000000
0!
0*
09
0>
0C
#870690000000
1!
1*
b10 6
19
1>
1C
b10 G
#870700000000
0!
0*
09
0>
0C
#870710000000
1!
1*
b11 6
19
1>
1C
b11 G
#870720000000
0!
0*
09
0>
0C
#870730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#870740000000
0!
0*
09
0>
0C
#870750000000
1!
1*
b101 6
19
1>
1C
b101 G
#870760000000
0!
0*
09
0>
0C
#870770000000
1!
1*
b110 6
19
1>
1C
b110 G
#870780000000
0!
0*
09
0>
0C
#870790000000
1!
1*
b111 6
19
1>
1C
b111 G
#870800000000
0!
0*
09
0>
0C
#870810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#870820000000
0!
0*
09
0>
0C
#870830000000
1!
1*
b1 6
19
1>
1C
b1 G
#870840000000
0!
0*
09
0>
0C
#870850000000
1!
1*
b10 6
19
1>
1C
b10 G
#870860000000
0!
0*
09
0>
0C
#870870000000
1!
1*
b11 6
19
1>
1C
b11 G
#870880000000
0!
0*
09
0>
0C
#870890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#870900000000
0!
0*
09
0>
0C
#870910000000
1!
1*
b101 6
19
1>
1C
b101 G
#870920000000
0!
0*
09
0>
0C
#870930000000
1!
1*
b110 6
19
1>
1C
b110 G
#870940000000
0!
0*
09
0>
0C
#870950000000
1!
1*
b111 6
19
1>
1C
b111 G
#870960000000
0!
0*
09
0>
0C
#870970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#870980000000
0!
0*
09
0>
0C
#870990000000
1!
1*
b1 6
19
1>
1C
b1 G
#871000000000
0!
0*
09
0>
0C
#871010000000
1!
1*
b10 6
19
1>
1C
b10 G
#871020000000
0!
0*
09
0>
0C
#871030000000
1!
1*
b11 6
19
1>
1C
b11 G
#871040000000
0!
0*
09
0>
0C
#871050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#871060000000
0!
0*
09
0>
0C
#871070000000
1!
1*
b101 6
19
1>
1C
b101 G
#871080000000
0!
0*
09
0>
0C
#871090000000
1!
1*
b110 6
19
1>
1C
b110 G
#871100000000
0!
0*
09
0>
0C
#871110000000
1!
1*
b111 6
19
1>
1C
b111 G
#871120000000
0!
1"
0*
1+
09
1:
0>
0C
#871130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#871140000000
0!
0*
09
0>
0C
#871150000000
1!
1*
b1 6
19
1>
1C
b1 G
#871160000000
0!
0*
09
0>
0C
#871170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#871180000000
0!
0*
09
0>
0C
#871190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#871200000000
0!
0*
09
0>
0C
#871210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#871220000000
0!
0*
09
0>
0C
#871230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#871240000000
0!
0#
0*
0,
09
0>
0?
0C
#871250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#871260000000
0!
0*
09
0>
0C
#871270000000
1!
1*
19
1>
1C
#871280000000
0!
0*
09
0>
0C
#871290000000
1!
1*
19
1>
1C
#871300000000
0!
0*
09
0>
0C
#871310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#871320000000
0!
0*
09
0>
0C
#871330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#871340000000
0!
0*
09
0>
0C
#871350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#871360000000
0!
0*
09
0>
0C
#871370000000
1!
1*
b10 6
19
1>
1C
b10 G
#871380000000
0!
0*
09
0>
0C
#871390000000
1!
1*
b11 6
19
1>
1C
b11 G
#871400000000
0!
0*
09
0>
0C
#871410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#871420000000
0!
0*
09
0>
0C
#871430000000
1!
1*
b101 6
19
1>
1C
b101 G
#871440000000
0!
0*
09
0>
0C
#871450000000
1!
1*
b110 6
19
1>
1C
b110 G
#871460000000
0!
0*
09
0>
0C
#871470000000
1!
1*
b111 6
19
1>
1C
b111 G
#871480000000
0!
0*
09
0>
0C
#871490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#871500000000
0!
0*
09
0>
0C
#871510000000
1!
1*
b1 6
19
1>
1C
b1 G
#871520000000
0!
0*
09
0>
0C
#871530000000
1!
1*
b10 6
19
1>
1C
b10 G
#871540000000
0!
0*
09
0>
0C
#871550000000
1!
1*
b11 6
19
1>
1C
b11 G
#871560000000
0!
0*
09
0>
0C
#871570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#871580000000
0!
0*
09
0>
0C
#871590000000
1!
1*
b101 6
19
1>
1C
b101 G
#871600000000
0!
0*
09
0>
0C
#871610000000
1!
1*
b110 6
19
1>
1C
b110 G
#871620000000
0!
0*
09
0>
0C
#871630000000
1!
1*
b111 6
19
1>
1C
b111 G
#871640000000
0!
0*
09
0>
0C
#871650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#871660000000
0!
0*
09
0>
0C
#871670000000
1!
1*
b1 6
19
1>
1C
b1 G
#871680000000
0!
0*
09
0>
0C
#871690000000
1!
1*
b10 6
19
1>
1C
b10 G
#871700000000
0!
0*
09
0>
0C
#871710000000
1!
1*
b11 6
19
1>
1C
b11 G
#871720000000
0!
0*
09
0>
0C
#871730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#871740000000
0!
0*
09
0>
0C
#871750000000
1!
1*
b101 6
19
1>
1C
b101 G
#871760000000
0!
0*
09
0>
0C
#871770000000
1!
1*
b110 6
19
1>
1C
b110 G
#871780000000
0!
0*
09
0>
0C
#871790000000
1!
1*
b111 6
19
1>
1C
b111 G
#871800000000
0!
1"
0*
1+
09
1:
0>
0C
#871810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#871820000000
0!
0*
09
0>
0C
#871830000000
1!
1*
b1 6
19
1>
1C
b1 G
#871840000000
0!
0*
09
0>
0C
#871850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#871860000000
0!
0*
09
0>
0C
#871870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#871880000000
0!
0*
09
0>
0C
#871890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#871900000000
0!
0*
09
0>
0C
#871910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#871920000000
0!
0#
0*
0,
09
0>
0?
0C
#871930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#871940000000
0!
0*
09
0>
0C
#871950000000
1!
1*
19
1>
1C
#871960000000
0!
0*
09
0>
0C
#871970000000
1!
1*
19
1>
1C
#871980000000
0!
0*
09
0>
0C
#871990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#872000000000
0!
0*
09
0>
0C
#872010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#872020000000
0!
0*
09
0>
0C
#872030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#872040000000
0!
0*
09
0>
0C
#872050000000
1!
1*
b10 6
19
1>
1C
b10 G
#872060000000
0!
0*
09
0>
0C
#872070000000
1!
1*
b11 6
19
1>
1C
b11 G
#872080000000
0!
0*
09
0>
0C
#872090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#872100000000
0!
0*
09
0>
0C
#872110000000
1!
1*
b101 6
19
1>
1C
b101 G
#872120000000
0!
0*
09
0>
0C
#872130000000
1!
1*
b110 6
19
1>
1C
b110 G
#872140000000
0!
0*
09
0>
0C
#872150000000
1!
1*
b111 6
19
1>
1C
b111 G
#872160000000
0!
0*
09
0>
0C
#872170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#872180000000
0!
0*
09
0>
0C
#872190000000
1!
1*
b1 6
19
1>
1C
b1 G
#872200000000
0!
0*
09
0>
0C
#872210000000
1!
1*
b10 6
19
1>
1C
b10 G
#872220000000
0!
0*
09
0>
0C
#872230000000
1!
1*
b11 6
19
1>
1C
b11 G
#872240000000
0!
0*
09
0>
0C
#872250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#872260000000
0!
0*
09
0>
0C
#872270000000
1!
1*
b101 6
19
1>
1C
b101 G
#872280000000
0!
0*
09
0>
0C
#872290000000
1!
1*
b110 6
19
1>
1C
b110 G
#872300000000
0!
0*
09
0>
0C
#872310000000
1!
1*
b111 6
19
1>
1C
b111 G
#872320000000
0!
0*
09
0>
0C
#872330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#872340000000
0!
0*
09
0>
0C
#872350000000
1!
1*
b1 6
19
1>
1C
b1 G
#872360000000
0!
0*
09
0>
0C
#872370000000
1!
1*
b10 6
19
1>
1C
b10 G
#872380000000
0!
0*
09
0>
0C
#872390000000
1!
1*
b11 6
19
1>
1C
b11 G
#872400000000
0!
0*
09
0>
0C
#872410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#872420000000
0!
0*
09
0>
0C
#872430000000
1!
1*
b101 6
19
1>
1C
b101 G
#872440000000
0!
0*
09
0>
0C
#872450000000
1!
1*
b110 6
19
1>
1C
b110 G
#872460000000
0!
0*
09
0>
0C
#872470000000
1!
1*
b111 6
19
1>
1C
b111 G
#872480000000
0!
1"
0*
1+
09
1:
0>
0C
#872490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#872500000000
0!
0*
09
0>
0C
#872510000000
1!
1*
b1 6
19
1>
1C
b1 G
#872520000000
0!
0*
09
0>
0C
#872530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#872540000000
0!
0*
09
0>
0C
#872550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#872560000000
0!
0*
09
0>
0C
#872570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#872580000000
0!
0*
09
0>
0C
#872590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#872600000000
0!
0#
0*
0,
09
0>
0?
0C
#872610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#872620000000
0!
0*
09
0>
0C
#872630000000
1!
1*
19
1>
1C
#872640000000
0!
0*
09
0>
0C
#872650000000
1!
1*
19
1>
1C
#872660000000
0!
0*
09
0>
0C
#872670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#872680000000
0!
0*
09
0>
0C
#872690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#872700000000
0!
0*
09
0>
0C
#872710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#872720000000
0!
0*
09
0>
0C
#872730000000
1!
1*
b10 6
19
1>
1C
b10 G
#872740000000
0!
0*
09
0>
0C
#872750000000
1!
1*
b11 6
19
1>
1C
b11 G
#872760000000
0!
0*
09
0>
0C
#872770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#872780000000
0!
0*
09
0>
0C
#872790000000
1!
1*
b101 6
19
1>
1C
b101 G
#872800000000
0!
0*
09
0>
0C
#872810000000
1!
1*
b110 6
19
1>
1C
b110 G
#872820000000
0!
0*
09
0>
0C
#872830000000
1!
1*
b111 6
19
1>
1C
b111 G
#872840000000
0!
0*
09
0>
0C
#872850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#872860000000
0!
0*
09
0>
0C
#872870000000
1!
1*
b1 6
19
1>
1C
b1 G
#872880000000
0!
0*
09
0>
0C
#872890000000
1!
1*
b10 6
19
1>
1C
b10 G
#872900000000
0!
0*
09
0>
0C
#872910000000
1!
1*
b11 6
19
1>
1C
b11 G
#872920000000
0!
0*
09
0>
0C
#872930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#872940000000
0!
0*
09
0>
0C
#872950000000
1!
1*
b101 6
19
1>
1C
b101 G
#872960000000
0!
0*
09
0>
0C
#872970000000
1!
1*
b110 6
19
1>
1C
b110 G
#872980000000
0!
0*
09
0>
0C
#872990000000
1!
1*
b111 6
19
1>
1C
b111 G
#873000000000
0!
0*
09
0>
0C
#873010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#873020000000
0!
0*
09
0>
0C
#873030000000
1!
1*
b1 6
19
1>
1C
b1 G
#873040000000
0!
0*
09
0>
0C
#873050000000
1!
1*
b10 6
19
1>
1C
b10 G
#873060000000
0!
0*
09
0>
0C
#873070000000
1!
1*
b11 6
19
1>
1C
b11 G
#873080000000
0!
0*
09
0>
0C
#873090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#873100000000
0!
0*
09
0>
0C
#873110000000
1!
1*
b101 6
19
1>
1C
b101 G
#873120000000
0!
0*
09
0>
0C
#873130000000
1!
1*
b110 6
19
1>
1C
b110 G
#873140000000
0!
0*
09
0>
0C
#873150000000
1!
1*
b111 6
19
1>
1C
b111 G
#873160000000
0!
1"
0*
1+
09
1:
0>
0C
#873170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#873180000000
0!
0*
09
0>
0C
#873190000000
1!
1*
b1 6
19
1>
1C
b1 G
#873200000000
0!
0*
09
0>
0C
#873210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#873220000000
0!
0*
09
0>
0C
#873230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#873240000000
0!
0*
09
0>
0C
#873250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#873260000000
0!
0*
09
0>
0C
#873270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#873280000000
0!
0#
0*
0,
09
0>
0?
0C
#873290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#873300000000
0!
0*
09
0>
0C
#873310000000
1!
1*
19
1>
1C
#873320000000
0!
0*
09
0>
0C
#873330000000
1!
1*
19
1>
1C
#873340000000
0!
0*
09
0>
0C
#873350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#873360000000
0!
0*
09
0>
0C
#873370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#873380000000
0!
0*
09
0>
0C
#873390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#873400000000
0!
0*
09
0>
0C
#873410000000
1!
1*
b10 6
19
1>
1C
b10 G
#873420000000
0!
0*
09
0>
0C
#873430000000
1!
1*
b11 6
19
1>
1C
b11 G
#873440000000
0!
0*
09
0>
0C
#873450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#873460000000
0!
0*
09
0>
0C
#873470000000
1!
1*
b101 6
19
1>
1C
b101 G
#873480000000
0!
0*
09
0>
0C
#873490000000
1!
1*
b110 6
19
1>
1C
b110 G
#873500000000
0!
0*
09
0>
0C
#873510000000
1!
1*
b111 6
19
1>
1C
b111 G
#873520000000
0!
0*
09
0>
0C
#873530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#873540000000
0!
0*
09
0>
0C
#873550000000
1!
1*
b1 6
19
1>
1C
b1 G
#873560000000
0!
0*
09
0>
0C
#873570000000
1!
1*
b10 6
19
1>
1C
b10 G
#873580000000
0!
0*
09
0>
0C
#873590000000
1!
1*
b11 6
19
1>
1C
b11 G
#873600000000
0!
0*
09
0>
0C
#873610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#873620000000
0!
0*
09
0>
0C
#873630000000
1!
1*
b101 6
19
1>
1C
b101 G
#873640000000
0!
0*
09
0>
0C
#873650000000
1!
1*
b110 6
19
1>
1C
b110 G
#873660000000
0!
0*
09
0>
0C
#873670000000
1!
1*
b111 6
19
1>
1C
b111 G
#873680000000
0!
0*
09
0>
0C
#873690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#873700000000
0!
0*
09
0>
0C
#873710000000
1!
1*
b1 6
19
1>
1C
b1 G
#873720000000
0!
0*
09
0>
0C
#873730000000
1!
1*
b10 6
19
1>
1C
b10 G
#873740000000
0!
0*
09
0>
0C
#873750000000
1!
1*
b11 6
19
1>
1C
b11 G
#873760000000
0!
0*
09
0>
0C
#873770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#873780000000
0!
0*
09
0>
0C
#873790000000
1!
1*
b101 6
19
1>
1C
b101 G
#873800000000
0!
0*
09
0>
0C
#873810000000
1!
1*
b110 6
19
1>
1C
b110 G
#873820000000
0!
0*
09
0>
0C
#873830000000
1!
1*
b111 6
19
1>
1C
b111 G
#873840000000
0!
1"
0*
1+
09
1:
0>
0C
#873850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#873860000000
0!
0*
09
0>
0C
#873870000000
1!
1*
b1 6
19
1>
1C
b1 G
#873880000000
0!
0*
09
0>
0C
#873890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#873900000000
0!
0*
09
0>
0C
#873910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#873920000000
0!
0*
09
0>
0C
#873930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#873940000000
0!
0*
09
0>
0C
#873950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#873960000000
0!
0#
0*
0,
09
0>
0?
0C
#873970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#873980000000
0!
0*
09
0>
0C
#873990000000
1!
1*
19
1>
1C
#874000000000
0!
0*
09
0>
0C
#874010000000
1!
1*
19
1>
1C
#874020000000
0!
0*
09
0>
0C
#874030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#874040000000
0!
0*
09
0>
0C
#874050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#874060000000
0!
0*
09
0>
0C
#874070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#874080000000
0!
0*
09
0>
0C
#874090000000
1!
1*
b10 6
19
1>
1C
b10 G
#874100000000
0!
0*
09
0>
0C
#874110000000
1!
1*
b11 6
19
1>
1C
b11 G
#874120000000
0!
0*
09
0>
0C
#874130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#874140000000
0!
0*
09
0>
0C
#874150000000
1!
1*
b101 6
19
1>
1C
b101 G
#874160000000
0!
0*
09
0>
0C
#874170000000
1!
1*
b110 6
19
1>
1C
b110 G
#874180000000
0!
0*
09
0>
0C
#874190000000
1!
1*
b111 6
19
1>
1C
b111 G
#874200000000
0!
0*
09
0>
0C
#874210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#874220000000
0!
0*
09
0>
0C
#874230000000
1!
1*
b1 6
19
1>
1C
b1 G
#874240000000
0!
0*
09
0>
0C
#874250000000
1!
1*
b10 6
19
1>
1C
b10 G
#874260000000
0!
0*
09
0>
0C
#874270000000
1!
1*
b11 6
19
1>
1C
b11 G
#874280000000
0!
0*
09
0>
0C
#874290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#874300000000
0!
0*
09
0>
0C
#874310000000
1!
1*
b101 6
19
1>
1C
b101 G
#874320000000
0!
0*
09
0>
0C
#874330000000
1!
1*
b110 6
19
1>
1C
b110 G
#874340000000
0!
0*
09
0>
0C
#874350000000
1!
1*
b111 6
19
1>
1C
b111 G
#874360000000
0!
0*
09
0>
0C
#874370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#874380000000
0!
0*
09
0>
0C
#874390000000
1!
1*
b1 6
19
1>
1C
b1 G
#874400000000
0!
0*
09
0>
0C
#874410000000
1!
1*
b10 6
19
1>
1C
b10 G
#874420000000
0!
0*
09
0>
0C
#874430000000
1!
1*
b11 6
19
1>
1C
b11 G
#874440000000
0!
0*
09
0>
0C
#874450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#874460000000
0!
0*
09
0>
0C
#874470000000
1!
1*
b101 6
19
1>
1C
b101 G
#874480000000
0!
0*
09
0>
0C
#874490000000
1!
1*
b110 6
19
1>
1C
b110 G
#874500000000
0!
0*
09
0>
0C
#874510000000
1!
1*
b111 6
19
1>
1C
b111 G
#874520000000
0!
1"
0*
1+
09
1:
0>
0C
#874530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#874540000000
0!
0*
09
0>
0C
#874550000000
1!
1*
b1 6
19
1>
1C
b1 G
#874560000000
0!
0*
09
0>
0C
#874570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#874580000000
0!
0*
09
0>
0C
#874590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#874600000000
0!
0*
09
0>
0C
#874610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#874620000000
0!
0*
09
0>
0C
#874630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#874640000000
0!
0#
0*
0,
09
0>
0?
0C
#874650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#874660000000
0!
0*
09
0>
0C
#874670000000
1!
1*
19
1>
1C
#874680000000
0!
0*
09
0>
0C
#874690000000
1!
1*
19
1>
1C
#874700000000
0!
0*
09
0>
0C
#874710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#874720000000
0!
0*
09
0>
0C
#874730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#874740000000
0!
0*
09
0>
0C
#874750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#874760000000
0!
0*
09
0>
0C
#874770000000
1!
1*
b10 6
19
1>
1C
b10 G
#874780000000
0!
0*
09
0>
0C
#874790000000
1!
1*
b11 6
19
1>
1C
b11 G
#874800000000
0!
0*
09
0>
0C
#874810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#874820000000
0!
0*
09
0>
0C
#874830000000
1!
1*
b101 6
19
1>
1C
b101 G
#874840000000
0!
0*
09
0>
0C
#874850000000
1!
1*
b110 6
19
1>
1C
b110 G
#874860000000
0!
0*
09
0>
0C
#874870000000
1!
1*
b111 6
19
1>
1C
b111 G
#874880000000
0!
0*
09
0>
0C
#874890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#874900000000
0!
0*
09
0>
0C
#874910000000
1!
1*
b1 6
19
1>
1C
b1 G
#874920000000
0!
0*
09
0>
0C
#874930000000
1!
1*
b10 6
19
1>
1C
b10 G
#874940000000
0!
0*
09
0>
0C
#874950000000
1!
1*
b11 6
19
1>
1C
b11 G
#874960000000
0!
0*
09
0>
0C
#874970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#874980000000
0!
0*
09
0>
0C
#874990000000
1!
1*
b101 6
19
1>
1C
b101 G
#875000000000
0!
0*
09
0>
0C
#875010000000
1!
1*
b110 6
19
1>
1C
b110 G
#875020000000
0!
0*
09
0>
0C
#875030000000
1!
1*
b111 6
19
1>
1C
b111 G
#875040000000
0!
0*
09
0>
0C
#875050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#875060000000
0!
0*
09
0>
0C
#875070000000
1!
1*
b1 6
19
1>
1C
b1 G
#875080000000
0!
0*
09
0>
0C
#875090000000
1!
1*
b10 6
19
1>
1C
b10 G
#875100000000
0!
0*
09
0>
0C
#875110000000
1!
1*
b11 6
19
1>
1C
b11 G
#875120000000
0!
0*
09
0>
0C
#875130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#875140000000
0!
0*
09
0>
0C
#875150000000
1!
1*
b101 6
19
1>
1C
b101 G
#875160000000
0!
0*
09
0>
0C
#875170000000
1!
1*
b110 6
19
1>
1C
b110 G
#875180000000
0!
0*
09
0>
0C
#875190000000
1!
1*
b111 6
19
1>
1C
b111 G
#875200000000
0!
1"
0*
1+
09
1:
0>
0C
#875210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#875220000000
0!
0*
09
0>
0C
#875230000000
1!
1*
b1 6
19
1>
1C
b1 G
#875240000000
0!
0*
09
0>
0C
#875250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#875260000000
0!
0*
09
0>
0C
#875270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#875280000000
0!
0*
09
0>
0C
#875290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#875300000000
0!
0*
09
0>
0C
#875310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#875320000000
0!
0#
0*
0,
09
0>
0?
0C
#875330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#875340000000
0!
0*
09
0>
0C
#875350000000
1!
1*
19
1>
1C
#875360000000
0!
0*
09
0>
0C
#875370000000
1!
1*
19
1>
1C
#875380000000
0!
0*
09
0>
0C
#875390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#875400000000
0!
0*
09
0>
0C
#875410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#875420000000
0!
0*
09
0>
0C
#875430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#875440000000
0!
0*
09
0>
0C
#875450000000
1!
1*
b10 6
19
1>
1C
b10 G
#875460000000
0!
0*
09
0>
0C
#875470000000
1!
1*
b11 6
19
1>
1C
b11 G
#875480000000
0!
0*
09
0>
0C
#875490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#875500000000
0!
0*
09
0>
0C
#875510000000
1!
1*
b101 6
19
1>
1C
b101 G
#875520000000
0!
0*
09
0>
0C
#875530000000
1!
1*
b110 6
19
1>
1C
b110 G
#875540000000
0!
0*
09
0>
0C
#875550000000
1!
1*
b111 6
19
1>
1C
b111 G
#875560000000
0!
0*
09
0>
0C
#875570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#875580000000
0!
0*
09
0>
0C
#875590000000
1!
1*
b1 6
19
1>
1C
b1 G
#875600000000
0!
0*
09
0>
0C
#875610000000
1!
1*
b10 6
19
1>
1C
b10 G
#875620000000
0!
0*
09
0>
0C
#875630000000
1!
1*
b11 6
19
1>
1C
b11 G
#875640000000
0!
0*
09
0>
0C
#875650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#875660000000
0!
0*
09
0>
0C
#875670000000
1!
1*
b101 6
19
1>
1C
b101 G
#875680000000
0!
0*
09
0>
0C
#875690000000
1!
1*
b110 6
19
1>
1C
b110 G
#875700000000
0!
0*
09
0>
0C
#875710000000
1!
1*
b111 6
19
1>
1C
b111 G
#875720000000
0!
0*
09
0>
0C
#875730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#875740000000
0!
0*
09
0>
0C
#875750000000
1!
1*
b1 6
19
1>
1C
b1 G
#875760000000
0!
0*
09
0>
0C
#875770000000
1!
1*
b10 6
19
1>
1C
b10 G
#875780000000
0!
0*
09
0>
0C
#875790000000
1!
1*
b11 6
19
1>
1C
b11 G
#875800000000
0!
0*
09
0>
0C
#875810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#875820000000
0!
0*
09
0>
0C
#875830000000
1!
1*
b101 6
19
1>
1C
b101 G
#875840000000
0!
0*
09
0>
0C
#875850000000
1!
1*
b110 6
19
1>
1C
b110 G
#875860000000
0!
0*
09
0>
0C
#875870000000
1!
1*
b111 6
19
1>
1C
b111 G
#875880000000
0!
1"
0*
1+
09
1:
0>
0C
#875890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#875900000000
0!
0*
09
0>
0C
#875910000000
1!
1*
b1 6
19
1>
1C
b1 G
#875920000000
0!
0*
09
0>
0C
#875930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#875940000000
0!
0*
09
0>
0C
#875950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#875960000000
0!
0*
09
0>
0C
#875970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#875980000000
0!
0*
09
0>
0C
#875990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#876000000000
0!
0#
0*
0,
09
0>
0?
0C
#876010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#876020000000
0!
0*
09
0>
0C
#876030000000
1!
1*
19
1>
1C
#876040000000
0!
0*
09
0>
0C
#876050000000
1!
1*
19
1>
1C
#876060000000
0!
0*
09
0>
0C
#876070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#876080000000
0!
0*
09
0>
0C
#876090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#876100000000
0!
0*
09
0>
0C
#876110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#876120000000
0!
0*
09
0>
0C
#876130000000
1!
1*
b10 6
19
1>
1C
b10 G
#876140000000
0!
0*
09
0>
0C
#876150000000
1!
1*
b11 6
19
1>
1C
b11 G
#876160000000
0!
0*
09
0>
0C
#876170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#876180000000
0!
0*
09
0>
0C
#876190000000
1!
1*
b101 6
19
1>
1C
b101 G
#876200000000
0!
0*
09
0>
0C
#876210000000
1!
1*
b110 6
19
1>
1C
b110 G
#876220000000
0!
0*
09
0>
0C
#876230000000
1!
1*
b111 6
19
1>
1C
b111 G
#876240000000
0!
0*
09
0>
0C
#876250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#876260000000
0!
0*
09
0>
0C
#876270000000
1!
1*
b1 6
19
1>
1C
b1 G
#876280000000
0!
0*
09
0>
0C
#876290000000
1!
1*
b10 6
19
1>
1C
b10 G
#876300000000
0!
0*
09
0>
0C
#876310000000
1!
1*
b11 6
19
1>
1C
b11 G
#876320000000
0!
0*
09
0>
0C
#876330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#876340000000
0!
0*
09
0>
0C
#876350000000
1!
1*
b101 6
19
1>
1C
b101 G
#876360000000
0!
0*
09
0>
0C
#876370000000
1!
1*
b110 6
19
1>
1C
b110 G
#876380000000
0!
0*
09
0>
0C
#876390000000
1!
1*
b111 6
19
1>
1C
b111 G
#876400000000
0!
0*
09
0>
0C
#876410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#876420000000
0!
0*
09
0>
0C
#876430000000
1!
1*
b1 6
19
1>
1C
b1 G
#876440000000
0!
0*
09
0>
0C
#876450000000
1!
1*
b10 6
19
1>
1C
b10 G
#876460000000
0!
0*
09
0>
0C
#876470000000
1!
1*
b11 6
19
1>
1C
b11 G
#876480000000
0!
0*
09
0>
0C
#876490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#876500000000
0!
0*
09
0>
0C
#876510000000
1!
1*
b101 6
19
1>
1C
b101 G
#876520000000
0!
0*
09
0>
0C
#876530000000
1!
1*
b110 6
19
1>
1C
b110 G
#876540000000
0!
0*
09
0>
0C
#876550000000
1!
1*
b111 6
19
1>
1C
b111 G
#876560000000
0!
1"
0*
1+
09
1:
0>
0C
#876570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#876580000000
0!
0*
09
0>
0C
#876590000000
1!
1*
b1 6
19
1>
1C
b1 G
#876600000000
0!
0*
09
0>
0C
#876610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#876620000000
0!
0*
09
0>
0C
#876630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#876640000000
0!
0*
09
0>
0C
#876650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#876660000000
0!
0*
09
0>
0C
#876670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#876680000000
0!
0#
0*
0,
09
0>
0?
0C
#876690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#876700000000
0!
0*
09
0>
0C
#876710000000
1!
1*
19
1>
1C
#876720000000
0!
0*
09
0>
0C
#876730000000
1!
1*
19
1>
1C
#876740000000
0!
0*
09
0>
0C
#876750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#876760000000
0!
0*
09
0>
0C
#876770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#876780000000
0!
0*
09
0>
0C
#876790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#876800000000
0!
0*
09
0>
0C
#876810000000
1!
1*
b10 6
19
1>
1C
b10 G
#876820000000
0!
0*
09
0>
0C
#876830000000
1!
1*
b11 6
19
1>
1C
b11 G
#876840000000
0!
0*
09
0>
0C
#876850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#876860000000
0!
0*
09
0>
0C
#876870000000
1!
1*
b101 6
19
1>
1C
b101 G
#876880000000
0!
0*
09
0>
0C
#876890000000
1!
1*
b110 6
19
1>
1C
b110 G
#876900000000
0!
0*
09
0>
0C
#876910000000
1!
1*
b111 6
19
1>
1C
b111 G
#876920000000
0!
0*
09
0>
0C
#876930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#876940000000
0!
0*
09
0>
0C
#876950000000
1!
1*
b1 6
19
1>
1C
b1 G
#876960000000
0!
0*
09
0>
0C
#876970000000
1!
1*
b10 6
19
1>
1C
b10 G
#876980000000
0!
0*
09
0>
0C
#876990000000
1!
1*
b11 6
19
1>
1C
b11 G
#877000000000
0!
0*
09
0>
0C
#877010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#877020000000
0!
0*
09
0>
0C
#877030000000
1!
1*
b101 6
19
1>
1C
b101 G
#877040000000
0!
0*
09
0>
0C
#877050000000
1!
1*
b110 6
19
1>
1C
b110 G
#877060000000
0!
0*
09
0>
0C
#877070000000
1!
1*
b111 6
19
1>
1C
b111 G
#877080000000
0!
0*
09
0>
0C
#877090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#877100000000
0!
0*
09
0>
0C
#877110000000
1!
1*
b1 6
19
1>
1C
b1 G
#877120000000
0!
0*
09
0>
0C
#877130000000
1!
1*
b10 6
19
1>
1C
b10 G
#877140000000
0!
0*
09
0>
0C
#877150000000
1!
1*
b11 6
19
1>
1C
b11 G
#877160000000
0!
0*
09
0>
0C
#877170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#877180000000
0!
0*
09
0>
0C
#877190000000
1!
1*
b101 6
19
1>
1C
b101 G
#877200000000
0!
0*
09
0>
0C
#877210000000
1!
1*
b110 6
19
1>
1C
b110 G
#877220000000
0!
0*
09
0>
0C
#877230000000
1!
1*
b111 6
19
1>
1C
b111 G
#877240000000
0!
1"
0*
1+
09
1:
0>
0C
#877250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#877260000000
0!
0*
09
0>
0C
#877270000000
1!
1*
b1 6
19
1>
1C
b1 G
#877280000000
0!
0*
09
0>
0C
#877290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#877300000000
0!
0*
09
0>
0C
#877310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#877320000000
0!
0*
09
0>
0C
#877330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#877340000000
0!
0*
09
0>
0C
#877350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#877360000000
0!
0#
0*
0,
09
0>
0?
0C
#877370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#877380000000
0!
0*
09
0>
0C
#877390000000
1!
1*
19
1>
1C
#877400000000
0!
0*
09
0>
0C
#877410000000
1!
1*
19
1>
1C
#877420000000
0!
0*
09
0>
0C
#877430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#877440000000
0!
0*
09
0>
0C
#877450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#877460000000
0!
0*
09
0>
0C
#877470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#877480000000
0!
0*
09
0>
0C
#877490000000
1!
1*
b10 6
19
1>
1C
b10 G
#877500000000
0!
0*
09
0>
0C
#877510000000
1!
1*
b11 6
19
1>
1C
b11 G
#877520000000
0!
0*
09
0>
0C
#877530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#877540000000
0!
0*
09
0>
0C
#877550000000
1!
1*
b101 6
19
1>
1C
b101 G
#877560000000
0!
0*
09
0>
0C
#877570000000
1!
1*
b110 6
19
1>
1C
b110 G
#877580000000
0!
0*
09
0>
0C
#877590000000
1!
1*
b111 6
19
1>
1C
b111 G
#877600000000
0!
0*
09
0>
0C
#877610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#877620000000
0!
0*
09
0>
0C
#877630000000
1!
1*
b1 6
19
1>
1C
b1 G
#877640000000
0!
0*
09
0>
0C
#877650000000
1!
1*
b10 6
19
1>
1C
b10 G
#877660000000
0!
0*
09
0>
0C
#877670000000
1!
1*
b11 6
19
1>
1C
b11 G
#877680000000
0!
0*
09
0>
0C
#877690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#877700000000
0!
0*
09
0>
0C
#877710000000
1!
1*
b101 6
19
1>
1C
b101 G
#877720000000
0!
0*
09
0>
0C
#877730000000
1!
1*
b110 6
19
1>
1C
b110 G
#877740000000
0!
0*
09
0>
0C
#877750000000
1!
1*
b111 6
19
1>
1C
b111 G
#877760000000
0!
0*
09
0>
0C
#877770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#877780000000
0!
0*
09
0>
0C
#877790000000
1!
1*
b1 6
19
1>
1C
b1 G
#877800000000
0!
0*
09
0>
0C
#877810000000
1!
1*
b10 6
19
1>
1C
b10 G
#877820000000
0!
0*
09
0>
0C
#877830000000
1!
1*
b11 6
19
1>
1C
b11 G
#877840000000
0!
0*
09
0>
0C
#877850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#877860000000
0!
0*
09
0>
0C
#877870000000
1!
1*
b101 6
19
1>
1C
b101 G
#877880000000
0!
0*
09
0>
0C
#877890000000
1!
1*
b110 6
19
1>
1C
b110 G
#877900000000
0!
0*
09
0>
0C
#877910000000
1!
1*
b111 6
19
1>
1C
b111 G
#877920000000
0!
1"
0*
1+
09
1:
0>
0C
#877930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#877940000000
0!
0*
09
0>
0C
#877950000000
1!
1*
b1 6
19
1>
1C
b1 G
#877960000000
0!
0*
09
0>
0C
#877970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#877980000000
0!
0*
09
0>
0C
#877990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#878000000000
0!
0*
09
0>
0C
#878010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#878020000000
0!
0*
09
0>
0C
#878030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#878040000000
0!
0#
0*
0,
09
0>
0?
0C
#878050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#878060000000
0!
0*
09
0>
0C
#878070000000
1!
1*
19
1>
1C
#878080000000
0!
0*
09
0>
0C
#878090000000
1!
1*
19
1>
1C
#878100000000
0!
0*
09
0>
0C
#878110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#878120000000
0!
0*
09
0>
0C
#878130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#878140000000
0!
0*
09
0>
0C
#878150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#878160000000
0!
0*
09
0>
0C
#878170000000
1!
1*
b10 6
19
1>
1C
b10 G
#878180000000
0!
0*
09
0>
0C
#878190000000
1!
1*
b11 6
19
1>
1C
b11 G
#878200000000
0!
0*
09
0>
0C
#878210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#878220000000
0!
0*
09
0>
0C
#878230000000
1!
1*
b101 6
19
1>
1C
b101 G
#878240000000
0!
0*
09
0>
0C
#878250000000
1!
1*
b110 6
19
1>
1C
b110 G
#878260000000
0!
0*
09
0>
0C
#878270000000
1!
1*
b111 6
19
1>
1C
b111 G
#878280000000
0!
0*
09
0>
0C
#878290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#878300000000
0!
0*
09
0>
0C
#878310000000
1!
1*
b1 6
19
1>
1C
b1 G
#878320000000
0!
0*
09
0>
0C
#878330000000
1!
1*
b10 6
19
1>
1C
b10 G
#878340000000
0!
0*
09
0>
0C
#878350000000
1!
1*
b11 6
19
1>
1C
b11 G
#878360000000
0!
0*
09
0>
0C
#878370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#878380000000
0!
0*
09
0>
0C
#878390000000
1!
1*
b101 6
19
1>
1C
b101 G
#878400000000
0!
0*
09
0>
0C
#878410000000
1!
1*
b110 6
19
1>
1C
b110 G
#878420000000
0!
0*
09
0>
0C
#878430000000
1!
1*
b111 6
19
1>
1C
b111 G
#878440000000
0!
0*
09
0>
0C
#878450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#878460000000
0!
0*
09
0>
0C
#878470000000
1!
1*
b1 6
19
1>
1C
b1 G
#878480000000
0!
0*
09
0>
0C
#878490000000
1!
1*
b10 6
19
1>
1C
b10 G
#878500000000
0!
0*
09
0>
0C
#878510000000
1!
1*
b11 6
19
1>
1C
b11 G
#878520000000
0!
0*
09
0>
0C
#878530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#878540000000
0!
0*
09
0>
0C
#878550000000
1!
1*
b101 6
19
1>
1C
b101 G
#878560000000
0!
0*
09
0>
0C
#878570000000
1!
1*
b110 6
19
1>
1C
b110 G
#878580000000
0!
0*
09
0>
0C
#878590000000
1!
1*
b111 6
19
1>
1C
b111 G
#878600000000
0!
1"
0*
1+
09
1:
0>
0C
#878610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#878620000000
0!
0*
09
0>
0C
#878630000000
1!
1*
b1 6
19
1>
1C
b1 G
#878640000000
0!
0*
09
0>
0C
#878650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#878660000000
0!
0*
09
0>
0C
#878670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#878680000000
0!
0*
09
0>
0C
#878690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#878700000000
0!
0*
09
0>
0C
#878710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#878720000000
0!
0#
0*
0,
09
0>
0?
0C
#878730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#878740000000
0!
0*
09
0>
0C
#878750000000
1!
1*
19
1>
1C
#878760000000
0!
0*
09
0>
0C
#878770000000
1!
1*
19
1>
1C
#878780000000
0!
0*
09
0>
0C
#878790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#878800000000
0!
0*
09
0>
0C
#878810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#878820000000
0!
0*
09
0>
0C
#878830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#878840000000
0!
0*
09
0>
0C
#878850000000
1!
1*
b10 6
19
1>
1C
b10 G
#878860000000
0!
0*
09
0>
0C
#878870000000
1!
1*
b11 6
19
1>
1C
b11 G
#878880000000
0!
0*
09
0>
0C
#878890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#878900000000
0!
0*
09
0>
0C
#878910000000
1!
1*
b101 6
19
1>
1C
b101 G
#878920000000
0!
0*
09
0>
0C
#878930000000
1!
1*
b110 6
19
1>
1C
b110 G
#878940000000
0!
0*
09
0>
0C
#878950000000
1!
1*
b111 6
19
1>
1C
b111 G
#878960000000
0!
0*
09
0>
0C
#878970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#878980000000
0!
0*
09
0>
0C
#878990000000
1!
1*
b1 6
19
1>
1C
b1 G
#879000000000
0!
0*
09
0>
0C
#879010000000
1!
1*
b10 6
19
1>
1C
b10 G
#879020000000
0!
0*
09
0>
0C
#879030000000
1!
1*
b11 6
19
1>
1C
b11 G
#879040000000
0!
0*
09
0>
0C
#879050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#879060000000
0!
0*
09
0>
0C
#879070000000
1!
1*
b101 6
19
1>
1C
b101 G
#879080000000
0!
0*
09
0>
0C
#879090000000
1!
1*
b110 6
19
1>
1C
b110 G
#879100000000
0!
0*
09
0>
0C
#879110000000
1!
1*
b111 6
19
1>
1C
b111 G
#879120000000
0!
0*
09
0>
0C
#879130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#879140000000
0!
0*
09
0>
0C
#879150000000
1!
1*
b1 6
19
1>
1C
b1 G
#879160000000
0!
0*
09
0>
0C
#879170000000
1!
1*
b10 6
19
1>
1C
b10 G
#879180000000
0!
0*
09
0>
0C
#879190000000
1!
1*
b11 6
19
1>
1C
b11 G
#879200000000
0!
0*
09
0>
0C
#879210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#879220000000
0!
0*
09
0>
0C
#879230000000
1!
1*
b101 6
19
1>
1C
b101 G
#879240000000
0!
0*
09
0>
0C
#879250000000
1!
1*
b110 6
19
1>
1C
b110 G
#879260000000
0!
0*
09
0>
0C
#879270000000
1!
1*
b111 6
19
1>
1C
b111 G
#879280000000
0!
1"
0*
1+
09
1:
0>
0C
#879290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#879300000000
0!
0*
09
0>
0C
#879310000000
1!
1*
b1 6
19
1>
1C
b1 G
#879320000000
0!
0*
09
0>
0C
#879330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#879340000000
0!
0*
09
0>
0C
#879350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#879360000000
0!
0*
09
0>
0C
#879370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#879380000000
0!
0*
09
0>
0C
#879390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#879400000000
0!
0#
0*
0,
09
0>
0?
0C
#879410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#879420000000
0!
0*
09
0>
0C
#879430000000
1!
1*
19
1>
1C
#879440000000
0!
0*
09
0>
0C
#879450000000
1!
1*
19
1>
1C
#879460000000
0!
0*
09
0>
0C
#879470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#879480000000
0!
0*
09
0>
0C
#879490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#879500000000
0!
0*
09
0>
0C
#879510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#879520000000
0!
0*
09
0>
0C
#879530000000
1!
1*
b10 6
19
1>
1C
b10 G
#879540000000
0!
0*
09
0>
0C
#879550000000
1!
1*
b11 6
19
1>
1C
b11 G
#879560000000
0!
0*
09
0>
0C
#879570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#879580000000
0!
0*
09
0>
0C
#879590000000
1!
1*
b101 6
19
1>
1C
b101 G
#879600000000
0!
0*
09
0>
0C
#879610000000
1!
1*
b110 6
19
1>
1C
b110 G
#879620000000
0!
0*
09
0>
0C
#879630000000
1!
1*
b111 6
19
1>
1C
b111 G
#879640000000
0!
0*
09
0>
0C
#879650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#879660000000
0!
0*
09
0>
0C
#879670000000
1!
1*
b1 6
19
1>
1C
b1 G
#879680000000
0!
0*
09
0>
0C
#879690000000
1!
1*
b10 6
19
1>
1C
b10 G
#879700000000
0!
0*
09
0>
0C
#879710000000
1!
1*
b11 6
19
1>
1C
b11 G
#879720000000
0!
0*
09
0>
0C
#879730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#879740000000
0!
0*
09
0>
0C
#879750000000
1!
1*
b101 6
19
1>
1C
b101 G
#879760000000
0!
0*
09
0>
0C
#879770000000
1!
1*
b110 6
19
1>
1C
b110 G
#879780000000
0!
0*
09
0>
0C
#879790000000
1!
1*
b111 6
19
1>
1C
b111 G
#879800000000
0!
0*
09
0>
0C
#879810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#879820000000
0!
0*
09
0>
0C
#879830000000
1!
1*
b1 6
19
1>
1C
b1 G
#879840000000
0!
0*
09
0>
0C
#879850000000
1!
1*
b10 6
19
1>
1C
b10 G
#879860000000
0!
0*
09
0>
0C
#879870000000
1!
1*
b11 6
19
1>
1C
b11 G
#879880000000
0!
0*
09
0>
0C
#879890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#879900000000
0!
0*
09
0>
0C
#879910000000
1!
1*
b101 6
19
1>
1C
b101 G
#879920000000
0!
0*
09
0>
0C
#879930000000
1!
1*
b110 6
19
1>
1C
b110 G
#879940000000
0!
0*
09
0>
0C
#879950000000
1!
1*
b111 6
19
1>
1C
b111 G
#879960000000
0!
1"
0*
1+
09
1:
0>
0C
#879970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#879980000000
0!
0*
09
0>
0C
#879990000000
1!
1*
b1 6
19
1>
1C
b1 G
#880000000000
0!
0*
09
0>
0C
#880010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#880020000000
0!
0*
09
0>
0C
#880030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#880040000000
0!
0*
09
0>
0C
#880050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#880060000000
0!
0*
09
0>
0C
#880070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#880080000000
0!
0#
0*
0,
09
0>
0?
0C
#880090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#880100000000
0!
0*
09
0>
0C
#880110000000
1!
1*
19
1>
1C
#880120000000
0!
0*
09
0>
0C
#880130000000
1!
1*
19
1>
1C
#880140000000
0!
0*
09
0>
0C
#880150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#880160000000
0!
0*
09
0>
0C
#880170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#880180000000
0!
0*
09
0>
0C
#880190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#880200000000
0!
0*
09
0>
0C
#880210000000
1!
1*
b10 6
19
1>
1C
b10 G
#880220000000
0!
0*
09
0>
0C
#880230000000
1!
1*
b11 6
19
1>
1C
b11 G
#880240000000
0!
0*
09
0>
0C
#880250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#880260000000
0!
0*
09
0>
0C
#880270000000
1!
1*
b101 6
19
1>
1C
b101 G
#880280000000
0!
0*
09
0>
0C
#880290000000
1!
1*
b110 6
19
1>
1C
b110 G
#880300000000
0!
0*
09
0>
0C
#880310000000
1!
1*
b111 6
19
1>
1C
b111 G
#880320000000
0!
0*
09
0>
0C
#880330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#880340000000
0!
0*
09
0>
0C
#880350000000
1!
1*
b1 6
19
1>
1C
b1 G
#880360000000
0!
0*
09
0>
0C
#880370000000
1!
1*
b10 6
19
1>
1C
b10 G
#880380000000
0!
0*
09
0>
0C
#880390000000
1!
1*
b11 6
19
1>
1C
b11 G
#880400000000
0!
0*
09
0>
0C
#880410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#880420000000
0!
0*
09
0>
0C
#880430000000
1!
1*
b101 6
19
1>
1C
b101 G
#880440000000
0!
0*
09
0>
0C
#880450000000
1!
1*
b110 6
19
1>
1C
b110 G
#880460000000
0!
0*
09
0>
0C
#880470000000
1!
1*
b111 6
19
1>
1C
b111 G
#880480000000
0!
0*
09
0>
0C
#880490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#880500000000
0!
0*
09
0>
0C
#880510000000
1!
1*
b1 6
19
1>
1C
b1 G
#880520000000
0!
0*
09
0>
0C
#880530000000
1!
1*
b10 6
19
1>
1C
b10 G
#880540000000
0!
0*
09
0>
0C
#880550000000
1!
1*
b11 6
19
1>
1C
b11 G
#880560000000
0!
0*
09
0>
0C
#880570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#880580000000
0!
0*
09
0>
0C
#880590000000
1!
1*
b101 6
19
1>
1C
b101 G
#880600000000
0!
0*
09
0>
0C
#880610000000
1!
1*
b110 6
19
1>
1C
b110 G
#880620000000
0!
0*
09
0>
0C
#880630000000
1!
1*
b111 6
19
1>
1C
b111 G
#880640000000
0!
1"
0*
1+
09
1:
0>
0C
#880650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#880660000000
0!
0*
09
0>
0C
#880670000000
1!
1*
b1 6
19
1>
1C
b1 G
#880680000000
0!
0*
09
0>
0C
#880690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#880700000000
0!
0*
09
0>
0C
#880710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#880720000000
0!
0*
09
0>
0C
#880730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#880740000000
0!
0*
09
0>
0C
#880750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#880760000000
0!
0#
0*
0,
09
0>
0?
0C
#880770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#880780000000
0!
0*
09
0>
0C
#880790000000
1!
1*
19
1>
1C
#880800000000
0!
0*
09
0>
0C
#880810000000
1!
1*
19
1>
1C
#880820000000
0!
0*
09
0>
0C
#880830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#880840000000
0!
0*
09
0>
0C
#880850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#880860000000
0!
0*
09
0>
0C
#880870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#880880000000
0!
0*
09
0>
0C
#880890000000
1!
1*
b10 6
19
1>
1C
b10 G
#880900000000
0!
0*
09
0>
0C
#880910000000
1!
1*
b11 6
19
1>
1C
b11 G
#880920000000
0!
0*
09
0>
0C
#880930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#880940000000
0!
0*
09
0>
0C
#880950000000
1!
1*
b101 6
19
1>
1C
b101 G
#880960000000
0!
0*
09
0>
0C
#880970000000
1!
1*
b110 6
19
1>
1C
b110 G
#880980000000
0!
0*
09
0>
0C
#880990000000
1!
1*
b111 6
19
1>
1C
b111 G
#881000000000
0!
0*
09
0>
0C
#881010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#881020000000
0!
0*
09
0>
0C
#881030000000
1!
1*
b1 6
19
1>
1C
b1 G
#881040000000
0!
0*
09
0>
0C
#881050000000
1!
1*
b10 6
19
1>
1C
b10 G
#881060000000
0!
0*
09
0>
0C
#881070000000
1!
1*
b11 6
19
1>
1C
b11 G
#881080000000
0!
0*
09
0>
0C
#881090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#881100000000
0!
0*
09
0>
0C
#881110000000
1!
1*
b101 6
19
1>
1C
b101 G
#881120000000
0!
0*
09
0>
0C
#881130000000
1!
1*
b110 6
19
1>
1C
b110 G
#881140000000
0!
0*
09
0>
0C
#881150000000
1!
1*
b111 6
19
1>
1C
b111 G
#881160000000
0!
0*
09
0>
0C
#881170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#881180000000
0!
0*
09
0>
0C
#881190000000
1!
1*
b1 6
19
1>
1C
b1 G
#881200000000
0!
0*
09
0>
0C
#881210000000
1!
1*
b10 6
19
1>
1C
b10 G
#881220000000
0!
0*
09
0>
0C
#881230000000
1!
1*
b11 6
19
1>
1C
b11 G
#881240000000
0!
0*
09
0>
0C
#881250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#881260000000
0!
0*
09
0>
0C
#881270000000
1!
1*
b101 6
19
1>
1C
b101 G
#881280000000
0!
0*
09
0>
0C
#881290000000
1!
1*
b110 6
19
1>
1C
b110 G
#881300000000
0!
0*
09
0>
0C
#881310000000
1!
1*
b111 6
19
1>
1C
b111 G
#881320000000
0!
1"
0*
1+
09
1:
0>
0C
#881330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#881340000000
0!
0*
09
0>
0C
#881350000000
1!
1*
b1 6
19
1>
1C
b1 G
#881360000000
0!
0*
09
0>
0C
#881370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#881380000000
0!
0*
09
0>
0C
#881390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#881400000000
0!
0*
09
0>
0C
#881410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#881420000000
0!
0*
09
0>
0C
#881430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#881440000000
0!
0#
0*
0,
09
0>
0?
0C
#881450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#881460000000
0!
0*
09
0>
0C
#881470000000
1!
1*
19
1>
1C
#881480000000
0!
0*
09
0>
0C
#881490000000
1!
1*
19
1>
1C
#881500000000
0!
0*
09
0>
0C
#881510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#881520000000
0!
0*
09
0>
0C
#881530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#881540000000
0!
0*
09
0>
0C
#881550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#881560000000
0!
0*
09
0>
0C
#881570000000
1!
1*
b10 6
19
1>
1C
b10 G
#881580000000
0!
0*
09
0>
0C
#881590000000
1!
1*
b11 6
19
1>
1C
b11 G
#881600000000
0!
0*
09
0>
0C
#881610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#881620000000
0!
0*
09
0>
0C
#881630000000
1!
1*
b101 6
19
1>
1C
b101 G
#881640000000
0!
0*
09
0>
0C
#881650000000
1!
1*
b110 6
19
1>
1C
b110 G
#881660000000
0!
0*
09
0>
0C
#881670000000
1!
1*
b111 6
19
1>
1C
b111 G
#881680000000
0!
0*
09
0>
0C
#881690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#881700000000
0!
0*
09
0>
0C
#881710000000
1!
1*
b1 6
19
1>
1C
b1 G
#881720000000
0!
0*
09
0>
0C
#881730000000
1!
1*
b10 6
19
1>
1C
b10 G
#881740000000
0!
0*
09
0>
0C
#881750000000
1!
1*
b11 6
19
1>
1C
b11 G
#881760000000
0!
0*
09
0>
0C
#881770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#881780000000
0!
0*
09
0>
0C
#881790000000
1!
1*
b101 6
19
1>
1C
b101 G
#881800000000
0!
0*
09
0>
0C
#881810000000
1!
1*
b110 6
19
1>
1C
b110 G
#881820000000
0!
0*
09
0>
0C
#881830000000
1!
1*
b111 6
19
1>
1C
b111 G
#881840000000
0!
0*
09
0>
0C
#881850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#881860000000
0!
0*
09
0>
0C
#881870000000
1!
1*
b1 6
19
1>
1C
b1 G
#881880000000
0!
0*
09
0>
0C
#881890000000
1!
1*
b10 6
19
1>
1C
b10 G
#881900000000
0!
0*
09
0>
0C
#881910000000
1!
1*
b11 6
19
1>
1C
b11 G
#881920000000
0!
0*
09
0>
0C
#881930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#881940000000
0!
0*
09
0>
0C
#881950000000
1!
1*
b101 6
19
1>
1C
b101 G
#881960000000
0!
0*
09
0>
0C
#881970000000
1!
1*
b110 6
19
1>
1C
b110 G
#881980000000
0!
0*
09
0>
0C
#881990000000
1!
1*
b111 6
19
1>
1C
b111 G
#882000000000
0!
1"
0*
1+
09
1:
0>
0C
#882010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#882020000000
0!
0*
09
0>
0C
#882030000000
1!
1*
b1 6
19
1>
1C
b1 G
#882040000000
0!
0*
09
0>
0C
#882050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#882060000000
0!
0*
09
0>
0C
#882070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#882080000000
0!
0*
09
0>
0C
#882090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#882100000000
0!
0*
09
0>
0C
#882110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#882120000000
0!
0#
0*
0,
09
0>
0?
0C
#882130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#882140000000
0!
0*
09
0>
0C
#882150000000
1!
1*
19
1>
1C
#882160000000
0!
0*
09
0>
0C
#882170000000
1!
1*
19
1>
1C
#882180000000
0!
0*
09
0>
0C
#882190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#882200000000
0!
0*
09
0>
0C
#882210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#882220000000
0!
0*
09
0>
0C
#882230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#882240000000
0!
0*
09
0>
0C
#882250000000
1!
1*
b10 6
19
1>
1C
b10 G
#882260000000
0!
0*
09
0>
0C
#882270000000
1!
1*
b11 6
19
1>
1C
b11 G
#882280000000
0!
0*
09
0>
0C
#882290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#882300000000
0!
0*
09
0>
0C
#882310000000
1!
1*
b101 6
19
1>
1C
b101 G
#882320000000
0!
0*
09
0>
0C
#882330000000
1!
1*
b110 6
19
1>
1C
b110 G
#882340000000
0!
0*
09
0>
0C
#882350000000
1!
1*
b111 6
19
1>
1C
b111 G
#882360000000
0!
0*
09
0>
0C
#882370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#882380000000
0!
0*
09
0>
0C
#882390000000
1!
1*
b1 6
19
1>
1C
b1 G
#882400000000
0!
0*
09
0>
0C
#882410000000
1!
1*
b10 6
19
1>
1C
b10 G
#882420000000
0!
0*
09
0>
0C
#882430000000
1!
1*
b11 6
19
1>
1C
b11 G
#882440000000
0!
0*
09
0>
0C
#882450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#882460000000
0!
0*
09
0>
0C
#882470000000
1!
1*
b101 6
19
1>
1C
b101 G
#882480000000
0!
0*
09
0>
0C
#882490000000
1!
1*
b110 6
19
1>
1C
b110 G
#882500000000
0!
0*
09
0>
0C
#882510000000
1!
1*
b111 6
19
1>
1C
b111 G
#882520000000
0!
0*
09
0>
0C
#882530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#882540000000
0!
0*
09
0>
0C
#882550000000
1!
1*
b1 6
19
1>
1C
b1 G
#882560000000
0!
0*
09
0>
0C
#882570000000
1!
1*
b10 6
19
1>
1C
b10 G
#882580000000
0!
0*
09
0>
0C
#882590000000
1!
1*
b11 6
19
1>
1C
b11 G
#882600000000
0!
0*
09
0>
0C
#882610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#882620000000
0!
0*
09
0>
0C
#882630000000
1!
1*
b101 6
19
1>
1C
b101 G
#882640000000
0!
0*
09
0>
0C
#882650000000
1!
1*
b110 6
19
1>
1C
b110 G
#882660000000
0!
0*
09
0>
0C
#882670000000
1!
1*
b111 6
19
1>
1C
b111 G
#882680000000
0!
1"
0*
1+
09
1:
0>
0C
#882690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#882700000000
0!
0*
09
0>
0C
#882710000000
1!
1*
b1 6
19
1>
1C
b1 G
#882720000000
0!
0*
09
0>
0C
#882730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#882740000000
0!
0*
09
0>
0C
#882750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#882760000000
0!
0*
09
0>
0C
#882770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#882780000000
0!
0*
09
0>
0C
#882790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#882800000000
0!
0#
0*
0,
09
0>
0?
0C
#882810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#882820000000
0!
0*
09
0>
0C
#882830000000
1!
1*
19
1>
1C
#882840000000
0!
0*
09
0>
0C
#882850000000
1!
1*
19
1>
1C
#882860000000
0!
0*
09
0>
0C
#882870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#882880000000
0!
0*
09
0>
0C
#882890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#882900000000
0!
0*
09
0>
0C
#882910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#882920000000
0!
0*
09
0>
0C
#882930000000
1!
1*
b10 6
19
1>
1C
b10 G
#882940000000
0!
0*
09
0>
0C
#882950000000
1!
1*
b11 6
19
1>
1C
b11 G
#882960000000
0!
0*
09
0>
0C
#882970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#882980000000
0!
0*
09
0>
0C
#882990000000
1!
1*
b101 6
19
1>
1C
b101 G
#883000000000
0!
0*
09
0>
0C
#883010000000
1!
1*
b110 6
19
1>
1C
b110 G
#883020000000
0!
0*
09
0>
0C
#883030000000
1!
1*
b111 6
19
1>
1C
b111 G
#883040000000
0!
0*
09
0>
0C
#883050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#883060000000
0!
0*
09
0>
0C
#883070000000
1!
1*
b1 6
19
1>
1C
b1 G
#883080000000
0!
0*
09
0>
0C
#883090000000
1!
1*
b10 6
19
1>
1C
b10 G
#883100000000
0!
0*
09
0>
0C
#883110000000
1!
1*
b11 6
19
1>
1C
b11 G
#883120000000
0!
0*
09
0>
0C
#883130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#883140000000
0!
0*
09
0>
0C
#883150000000
1!
1*
b101 6
19
1>
1C
b101 G
#883160000000
0!
0*
09
0>
0C
#883170000000
1!
1*
b110 6
19
1>
1C
b110 G
#883180000000
0!
0*
09
0>
0C
#883190000000
1!
1*
b111 6
19
1>
1C
b111 G
#883200000000
0!
0*
09
0>
0C
#883210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#883220000000
0!
0*
09
0>
0C
#883230000000
1!
1*
b1 6
19
1>
1C
b1 G
#883240000000
0!
0*
09
0>
0C
#883250000000
1!
1*
b10 6
19
1>
1C
b10 G
#883260000000
0!
0*
09
0>
0C
#883270000000
1!
1*
b11 6
19
1>
1C
b11 G
#883280000000
0!
0*
09
0>
0C
#883290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#883300000000
0!
0*
09
0>
0C
#883310000000
1!
1*
b101 6
19
1>
1C
b101 G
#883320000000
0!
0*
09
0>
0C
#883330000000
1!
1*
b110 6
19
1>
1C
b110 G
#883340000000
0!
0*
09
0>
0C
#883350000000
1!
1*
b111 6
19
1>
1C
b111 G
#883360000000
0!
1"
0*
1+
09
1:
0>
0C
#883370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#883380000000
0!
0*
09
0>
0C
#883390000000
1!
1*
b1 6
19
1>
1C
b1 G
#883400000000
0!
0*
09
0>
0C
#883410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#883420000000
0!
0*
09
0>
0C
#883430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#883440000000
0!
0*
09
0>
0C
#883450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#883460000000
0!
0*
09
0>
0C
#883470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#883480000000
0!
0#
0*
0,
09
0>
0?
0C
#883490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#883500000000
0!
0*
09
0>
0C
#883510000000
1!
1*
19
1>
1C
#883520000000
0!
0*
09
0>
0C
#883530000000
1!
1*
19
1>
1C
#883540000000
0!
0*
09
0>
0C
#883550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#883560000000
0!
0*
09
0>
0C
#883570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#883580000000
0!
0*
09
0>
0C
#883590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#883600000000
0!
0*
09
0>
0C
#883610000000
1!
1*
b10 6
19
1>
1C
b10 G
#883620000000
0!
0*
09
0>
0C
#883630000000
1!
1*
b11 6
19
1>
1C
b11 G
#883640000000
0!
0*
09
0>
0C
#883650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#883660000000
0!
0*
09
0>
0C
#883670000000
1!
1*
b101 6
19
1>
1C
b101 G
#883680000000
0!
0*
09
0>
0C
#883690000000
1!
1*
b110 6
19
1>
1C
b110 G
#883700000000
0!
0*
09
0>
0C
#883710000000
1!
1*
b111 6
19
1>
1C
b111 G
#883720000000
0!
0*
09
0>
0C
#883730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#883740000000
0!
0*
09
0>
0C
#883750000000
1!
1*
b1 6
19
1>
1C
b1 G
#883760000000
0!
0*
09
0>
0C
#883770000000
1!
1*
b10 6
19
1>
1C
b10 G
#883780000000
0!
0*
09
0>
0C
#883790000000
1!
1*
b11 6
19
1>
1C
b11 G
#883800000000
0!
0*
09
0>
0C
#883810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#883820000000
0!
0*
09
0>
0C
#883830000000
1!
1*
b101 6
19
1>
1C
b101 G
#883840000000
0!
0*
09
0>
0C
#883850000000
1!
1*
b110 6
19
1>
1C
b110 G
#883860000000
0!
0*
09
0>
0C
#883870000000
1!
1*
b111 6
19
1>
1C
b111 G
#883880000000
0!
0*
09
0>
0C
#883890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#883900000000
0!
0*
09
0>
0C
#883910000000
1!
1*
b1 6
19
1>
1C
b1 G
#883920000000
0!
0*
09
0>
0C
#883930000000
1!
1*
b10 6
19
1>
1C
b10 G
#883940000000
0!
0*
09
0>
0C
#883950000000
1!
1*
b11 6
19
1>
1C
b11 G
#883960000000
0!
0*
09
0>
0C
#883970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#883980000000
0!
0*
09
0>
0C
#883990000000
1!
1*
b101 6
19
1>
1C
b101 G
#884000000000
0!
0*
09
0>
0C
#884010000000
1!
1*
b110 6
19
1>
1C
b110 G
#884020000000
0!
0*
09
0>
0C
#884030000000
1!
1*
b111 6
19
1>
1C
b111 G
#884040000000
0!
1"
0*
1+
09
1:
0>
0C
#884050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#884060000000
0!
0*
09
0>
0C
#884070000000
1!
1*
b1 6
19
1>
1C
b1 G
#884080000000
0!
0*
09
0>
0C
#884090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#884100000000
0!
0*
09
0>
0C
#884110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#884120000000
0!
0*
09
0>
0C
#884130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#884140000000
0!
0*
09
0>
0C
#884150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#884160000000
0!
0#
0*
0,
09
0>
0?
0C
#884170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#884180000000
0!
0*
09
0>
0C
#884190000000
1!
1*
19
1>
1C
#884200000000
0!
0*
09
0>
0C
#884210000000
1!
1*
19
1>
1C
#884220000000
0!
0*
09
0>
0C
#884230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#884240000000
0!
0*
09
0>
0C
#884250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#884260000000
0!
0*
09
0>
0C
#884270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#884280000000
0!
0*
09
0>
0C
#884290000000
1!
1*
b10 6
19
1>
1C
b10 G
#884300000000
0!
0*
09
0>
0C
#884310000000
1!
1*
b11 6
19
1>
1C
b11 G
#884320000000
0!
0*
09
0>
0C
#884330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#884340000000
0!
0*
09
0>
0C
#884350000000
1!
1*
b101 6
19
1>
1C
b101 G
#884360000000
0!
0*
09
0>
0C
#884370000000
1!
1*
b110 6
19
1>
1C
b110 G
#884380000000
0!
0*
09
0>
0C
#884390000000
1!
1*
b111 6
19
1>
1C
b111 G
#884400000000
0!
0*
09
0>
0C
#884410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#884420000000
0!
0*
09
0>
0C
#884430000000
1!
1*
b1 6
19
1>
1C
b1 G
#884440000000
0!
0*
09
0>
0C
#884450000000
1!
1*
b10 6
19
1>
1C
b10 G
#884460000000
0!
0*
09
0>
0C
#884470000000
1!
1*
b11 6
19
1>
1C
b11 G
#884480000000
0!
0*
09
0>
0C
#884490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#884500000000
0!
0*
09
0>
0C
#884510000000
1!
1*
b101 6
19
1>
1C
b101 G
#884520000000
0!
0*
09
0>
0C
#884530000000
1!
1*
b110 6
19
1>
1C
b110 G
#884540000000
0!
0*
09
0>
0C
#884550000000
1!
1*
b111 6
19
1>
1C
b111 G
#884560000000
0!
0*
09
0>
0C
#884570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#884580000000
0!
0*
09
0>
0C
#884590000000
1!
1*
b1 6
19
1>
1C
b1 G
#884600000000
0!
0*
09
0>
0C
#884610000000
1!
1*
b10 6
19
1>
1C
b10 G
#884620000000
0!
0*
09
0>
0C
#884630000000
1!
1*
b11 6
19
1>
1C
b11 G
#884640000000
0!
0*
09
0>
0C
#884650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#884660000000
0!
0*
09
0>
0C
#884670000000
1!
1*
b101 6
19
1>
1C
b101 G
#884680000000
0!
0*
09
0>
0C
#884690000000
1!
1*
b110 6
19
1>
1C
b110 G
#884700000000
0!
0*
09
0>
0C
#884710000000
1!
1*
b111 6
19
1>
1C
b111 G
#884720000000
0!
1"
0*
1+
09
1:
0>
0C
#884730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#884740000000
0!
0*
09
0>
0C
#884750000000
1!
1*
b1 6
19
1>
1C
b1 G
#884760000000
0!
0*
09
0>
0C
#884770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#884780000000
0!
0*
09
0>
0C
#884790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#884800000000
0!
0*
09
0>
0C
#884810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#884820000000
0!
0*
09
0>
0C
#884830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#884840000000
0!
0#
0*
0,
09
0>
0?
0C
#884850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#884860000000
0!
0*
09
0>
0C
#884870000000
1!
1*
19
1>
1C
#884880000000
0!
0*
09
0>
0C
#884890000000
1!
1*
19
1>
1C
#884900000000
0!
0*
09
0>
0C
#884910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#884920000000
0!
0*
09
0>
0C
#884930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#884940000000
0!
0*
09
0>
0C
#884950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#884960000000
0!
0*
09
0>
0C
#884970000000
1!
1*
b10 6
19
1>
1C
b10 G
#884980000000
0!
0*
09
0>
0C
#884990000000
1!
1*
b11 6
19
1>
1C
b11 G
#885000000000
0!
0*
09
0>
0C
#885010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#885020000000
0!
0*
09
0>
0C
#885030000000
1!
1*
b101 6
19
1>
1C
b101 G
#885040000000
0!
0*
09
0>
0C
#885050000000
1!
1*
b110 6
19
1>
1C
b110 G
#885060000000
0!
0*
09
0>
0C
#885070000000
1!
1*
b111 6
19
1>
1C
b111 G
#885080000000
0!
0*
09
0>
0C
#885090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#885100000000
0!
0*
09
0>
0C
#885110000000
1!
1*
b1 6
19
1>
1C
b1 G
#885120000000
0!
0*
09
0>
0C
#885130000000
1!
1*
b10 6
19
1>
1C
b10 G
#885140000000
0!
0*
09
0>
0C
#885150000000
1!
1*
b11 6
19
1>
1C
b11 G
#885160000000
0!
0*
09
0>
0C
#885170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#885180000000
0!
0*
09
0>
0C
#885190000000
1!
1*
b101 6
19
1>
1C
b101 G
#885200000000
0!
0*
09
0>
0C
#885210000000
1!
1*
b110 6
19
1>
1C
b110 G
#885220000000
0!
0*
09
0>
0C
#885230000000
1!
1*
b111 6
19
1>
1C
b111 G
#885240000000
0!
0*
09
0>
0C
#885250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#885260000000
0!
0*
09
0>
0C
#885270000000
1!
1*
b1 6
19
1>
1C
b1 G
#885280000000
0!
0*
09
0>
0C
#885290000000
1!
1*
b10 6
19
1>
1C
b10 G
#885300000000
0!
0*
09
0>
0C
#885310000000
1!
1*
b11 6
19
1>
1C
b11 G
#885320000000
0!
0*
09
0>
0C
#885330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#885340000000
0!
0*
09
0>
0C
#885350000000
1!
1*
b101 6
19
1>
1C
b101 G
#885360000000
0!
0*
09
0>
0C
#885370000000
1!
1*
b110 6
19
1>
1C
b110 G
#885380000000
0!
0*
09
0>
0C
#885390000000
1!
1*
b111 6
19
1>
1C
b111 G
#885400000000
0!
1"
0*
1+
09
1:
0>
0C
#885410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#885420000000
0!
0*
09
0>
0C
#885430000000
1!
1*
b1 6
19
1>
1C
b1 G
#885440000000
0!
0*
09
0>
0C
#885450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#885460000000
0!
0*
09
0>
0C
#885470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#885480000000
0!
0*
09
0>
0C
#885490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#885500000000
0!
0*
09
0>
0C
#885510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#885520000000
0!
0#
0*
0,
09
0>
0?
0C
#885530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#885540000000
0!
0*
09
0>
0C
#885550000000
1!
1*
19
1>
1C
#885560000000
0!
0*
09
0>
0C
#885570000000
1!
1*
19
1>
1C
#885580000000
0!
0*
09
0>
0C
#885590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#885600000000
0!
0*
09
0>
0C
#885610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#885620000000
0!
0*
09
0>
0C
#885630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#885640000000
0!
0*
09
0>
0C
#885650000000
1!
1*
b10 6
19
1>
1C
b10 G
#885660000000
0!
0*
09
0>
0C
#885670000000
1!
1*
b11 6
19
1>
1C
b11 G
#885680000000
0!
0*
09
0>
0C
#885690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#885700000000
0!
0*
09
0>
0C
#885710000000
1!
1*
b101 6
19
1>
1C
b101 G
#885720000000
0!
0*
09
0>
0C
#885730000000
1!
1*
b110 6
19
1>
1C
b110 G
#885740000000
0!
0*
09
0>
0C
#885750000000
1!
1*
b111 6
19
1>
1C
b111 G
#885760000000
0!
0*
09
0>
0C
#885770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#885780000000
0!
0*
09
0>
0C
#885790000000
1!
1*
b1 6
19
1>
1C
b1 G
#885800000000
0!
0*
09
0>
0C
#885810000000
1!
1*
b10 6
19
1>
1C
b10 G
#885820000000
0!
0*
09
0>
0C
#885830000000
1!
1*
b11 6
19
1>
1C
b11 G
#885840000000
0!
0*
09
0>
0C
#885850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#885860000000
0!
0*
09
0>
0C
#885870000000
1!
1*
b101 6
19
1>
1C
b101 G
#885880000000
0!
0*
09
0>
0C
#885890000000
1!
1*
b110 6
19
1>
1C
b110 G
#885900000000
0!
0*
09
0>
0C
#885910000000
1!
1*
b111 6
19
1>
1C
b111 G
#885920000000
0!
0*
09
0>
0C
#885930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#885940000000
0!
0*
09
0>
0C
#885950000000
1!
1*
b1 6
19
1>
1C
b1 G
#885960000000
0!
0*
09
0>
0C
#885970000000
1!
1*
b10 6
19
1>
1C
b10 G
#885980000000
0!
0*
09
0>
0C
#885990000000
1!
1*
b11 6
19
1>
1C
b11 G
#886000000000
0!
0*
09
0>
0C
#886010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#886020000000
0!
0*
09
0>
0C
#886030000000
1!
1*
b101 6
19
1>
1C
b101 G
#886040000000
0!
0*
09
0>
0C
#886050000000
1!
1*
b110 6
19
1>
1C
b110 G
#886060000000
0!
0*
09
0>
0C
#886070000000
1!
1*
b111 6
19
1>
1C
b111 G
#886080000000
0!
1"
0*
1+
09
1:
0>
0C
#886090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#886100000000
0!
0*
09
0>
0C
#886110000000
1!
1*
b1 6
19
1>
1C
b1 G
#886120000000
0!
0*
09
0>
0C
#886130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#886140000000
0!
0*
09
0>
0C
#886150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#886160000000
0!
0*
09
0>
0C
#886170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#886180000000
0!
0*
09
0>
0C
#886190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#886200000000
0!
0#
0*
0,
09
0>
0?
0C
#886210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#886220000000
0!
0*
09
0>
0C
#886230000000
1!
1*
19
1>
1C
#886240000000
0!
0*
09
0>
0C
#886250000000
1!
1*
19
1>
1C
#886260000000
0!
0*
09
0>
0C
#886270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#886280000000
0!
0*
09
0>
0C
#886290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#886300000000
0!
0*
09
0>
0C
#886310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#886320000000
0!
0*
09
0>
0C
#886330000000
1!
1*
b10 6
19
1>
1C
b10 G
#886340000000
0!
0*
09
0>
0C
#886350000000
1!
1*
b11 6
19
1>
1C
b11 G
#886360000000
0!
0*
09
0>
0C
#886370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#886380000000
0!
0*
09
0>
0C
#886390000000
1!
1*
b101 6
19
1>
1C
b101 G
#886400000000
0!
0*
09
0>
0C
#886410000000
1!
1*
b110 6
19
1>
1C
b110 G
#886420000000
0!
0*
09
0>
0C
#886430000000
1!
1*
b111 6
19
1>
1C
b111 G
#886440000000
0!
0*
09
0>
0C
#886450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#886460000000
0!
0*
09
0>
0C
#886470000000
1!
1*
b1 6
19
1>
1C
b1 G
#886480000000
0!
0*
09
0>
0C
#886490000000
1!
1*
b10 6
19
1>
1C
b10 G
#886500000000
0!
0*
09
0>
0C
#886510000000
1!
1*
b11 6
19
1>
1C
b11 G
#886520000000
0!
0*
09
0>
0C
#886530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#886540000000
0!
0*
09
0>
0C
#886550000000
1!
1*
b101 6
19
1>
1C
b101 G
#886560000000
0!
0*
09
0>
0C
#886570000000
1!
1*
b110 6
19
1>
1C
b110 G
#886580000000
0!
0*
09
0>
0C
#886590000000
1!
1*
b111 6
19
1>
1C
b111 G
#886600000000
0!
0*
09
0>
0C
#886610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#886620000000
0!
0*
09
0>
0C
#886630000000
1!
1*
b1 6
19
1>
1C
b1 G
#886640000000
0!
0*
09
0>
0C
#886650000000
1!
1*
b10 6
19
1>
1C
b10 G
#886660000000
0!
0*
09
0>
0C
#886670000000
1!
1*
b11 6
19
1>
1C
b11 G
#886680000000
0!
0*
09
0>
0C
#886690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#886700000000
0!
0*
09
0>
0C
#886710000000
1!
1*
b101 6
19
1>
1C
b101 G
#886720000000
0!
0*
09
0>
0C
#886730000000
1!
1*
b110 6
19
1>
1C
b110 G
#886740000000
0!
0*
09
0>
0C
#886750000000
1!
1*
b111 6
19
1>
1C
b111 G
#886760000000
0!
1"
0*
1+
09
1:
0>
0C
#886770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#886780000000
0!
0*
09
0>
0C
#886790000000
1!
1*
b1 6
19
1>
1C
b1 G
#886800000000
0!
0*
09
0>
0C
#886810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#886820000000
0!
0*
09
0>
0C
#886830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#886840000000
0!
0*
09
0>
0C
#886850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#886860000000
0!
0*
09
0>
0C
#886870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#886880000000
0!
0#
0*
0,
09
0>
0?
0C
#886890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#886900000000
0!
0*
09
0>
0C
#886910000000
1!
1*
19
1>
1C
#886920000000
0!
0*
09
0>
0C
#886930000000
1!
1*
19
1>
1C
#886940000000
0!
0*
09
0>
0C
#886950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#886960000000
0!
0*
09
0>
0C
#886970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#886980000000
0!
0*
09
0>
0C
#886990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#887000000000
0!
0*
09
0>
0C
#887010000000
1!
1*
b10 6
19
1>
1C
b10 G
#887020000000
0!
0*
09
0>
0C
#887030000000
1!
1*
b11 6
19
1>
1C
b11 G
#887040000000
0!
0*
09
0>
0C
#887050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#887060000000
0!
0*
09
0>
0C
#887070000000
1!
1*
b101 6
19
1>
1C
b101 G
#887080000000
0!
0*
09
0>
0C
#887090000000
1!
1*
b110 6
19
1>
1C
b110 G
#887100000000
0!
0*
09
0>
0C
#887110000000
1!
1*
b111 6
19
1>
1C
b111 G
#887120000000
0!
0*
09
0>
0C
#887130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#887140000000
0!
0*
09
0>
0C
#887150000000
1!
1*
b1 6
19
1>
1C
b1 G
#887160000000
0!
0*
09
0>
0C
#887170000000
1!
1*
b10 6
19
1>
1C
b10 G
#887180000000
0!
0*
09
0>
0C
#887190000000
1!
1*
b11 6
19
1>
1C
b11 G
#887200000000
0!
0*
09
0>
0C
#887210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#887220000000
0!
0*
09
0>
0C
#887230000000
1!
1*
b101 6
19
1>
1C
b101 G
#887240000000
0!
0*
09
0>
0C
#887250000000
1!
1*
b110 6
19
1>
1C
b110 G
#887260000000
0!
0*
09
0>
0C
#887270000000
1!
1*
b111 6
19
1>
1C
b111 G
#887280000000
0!
0*
09
0>
0C
#887290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#887300000000
0!
0*
09
0>
0C
#887310000000
1!
1*
b1 6
19
1>
1C
b1 G
#887320000000
0!
0*
09
0>
0C
#887330000000
1!
1*
b10 6
19
1>
1C
b10 G
#887340000000
0!
0*
09
0>
0C
#887350000000
1!
1*
b11 6
19
1>
1C
b11 G
#887360000000
0!
0*
09
0>
0C
#887370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#887380000000
0!
0*
09
0>
0C
#887390000000
1!
1*
b101 6
19
1>
1C
b101 G
#887400000000
0!
0*
09
0>
0C
#887410000000
1!
1*
b110 6
19
1>
1C
b110 G
#887420000000
0!
0*
09
0>
0C
#887430000000
1!
1*
b111 6
19
1>
1C
b111 G
#887440000000
0!
1"
0*
1+
09
1:
0>
0C
#887450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#887460000000
0!
0*
09
0>
0C
#887470000000
1!
1*
b1 6
19
1>
1C
b1 G
#887480000000
0!
0*
09
0>
0C
#887490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#887500000000
0!
0*
09
0>
0C
#887510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#887520000000
0!
0*
09
0>
0C
#887530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#887540000000
0!
0*
09
0>
0C
#887550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#887560000000
0!
0#
0*
0,
09
0>
0?
0C
#887570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#887580000000
0!
0*
09
0>
0C
#887590000000
1!
1*
19
1>
1C
#887600000000
0!
0*
09
0>
0C
#887610000000
1!
1*
19
1>
1C
#887620000000
0!
0*
09
0>
0C
#887630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#887640000000
0!
0*
09
0>
0C
#887650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#887660000000
0!
0*
09
0>
0C
#887670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#887680000000
0!
0*
09
0>
0C
#887690000000
1!
1*
b10 6
19
1>
1C
b10 G
#887700000000
0!
0*
09
0>
0C
#887710000000
1!
1*
b11 6
19
1>
1C
b11 G
#887720000000
0!
0*
09
0>
0C
#887730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#887740000000
0!
0*
09
0>
0C
#887750000000
1!
1*
b101 6
19
1>
1C
b101 G
#887760000000
0!
0*
09
0>
0C
#887770000000
1!
1*
b110 6
19
1>
1C
b110 G
#887780000000
0!
0*
09
0>
0C
#887790000000
1!
1*
b111 6
19
1>
1C
b111 G
#887800000000
0!
0*
09
0>
0C
#887810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#887820000000
0!
0*
09
0>
0C
#887830000000
1!
1*
b1 6
19
1>
1C
b1 G
#887840000000
0!
0*
09
0>
0C
#887850000000
1!
1*
b10 6
19
1>
1C
b10 G
#887860000000
0!
0*
09
0>
0C
#887870000000
1!
1*
b11 6
19
1>
1C
b11 G
#887880000000
0!
0*
09
0>
0C
#887890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#887900000000
0!
0*
09
0>
0C
#887910000000
1!
1*
b101 6
19
1>
1C
b101 G
#887920000000
0!
0*
09
0>
0C
#887930000000
1!
1*
b110 6
19
1>
1C
b110 G
#887940000000
0!
0*
09
0>
0C
#887950000000
1!
1*
b111 6
19
1>
1C
b111 G
#887960000000
0!
0*
09
0>
0C
#887970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#887980000000
0!
0*
09
0>
0C
#887990000000
1!
1*
b1 6
19
1>
1C
b1 G
#888000000000
0!
0*
09
0>
0C
#888010000000
1!
1*
b10 6
19
1>
1C
b10 G
#888020000000
0!
0*
09
0>
0C
#888030000000
1!
1*
b11 6
19
1>
1C
b11 G
#888040000000
0!
0*
09
0>
0C
#888050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#888060000000
0!
0*
09
0>
0C
#888070000000
1!
1*
b101 6
19
1>
1C
b101 G
#888080000000
0!
0*
09
0>
0C
#888090000000
1!
1*
b110 6
19
1>
1C
b110 G
#888100000000
0!
0*
09
0>
0C
#888110000000
1!
1*
b111 6
19
1>
1C
b111 G
#888120000000
0!
1"
0*
1+
09
1:
0>
0C
#888130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#888140000000
0!
0*
09
0>
0C
#888150000000
1!
1*
b1 6
19
1>
1C
b1 G
#888160000000
0!
0*
09
0>
0C
#888170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#888180000000
0!
0*
09
0>
0C
#888190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#888200000000
0!
0*
09
0>
0C
#888210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#888220000000
0!
0*
09
0>
0C
#888230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#888240000000
0!
0#
0*
0,
09
0>
0?
0C
#888250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#888260000000
0!
0*
09
0>
0C
#888270000000
1!
1*
19
1>
1C
#888280000000
0!
0*
09
0>
0C
#888290000000
1!
1*
19
1>
1C
#888300000000
0!
0*
09
0>
0C
#888310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#888320000000
0!
0*
09
0>
0C
#888330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#888340000000
0!
0*
09
0>
0C
#888350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#888360000000
0!
0*
09
0>
0C
#888370000000
1!
1*
b10 6
19
1>
1C
b10 G
#888380000000
0!
0*
09
0>
0C
#888390000000
1!
1*
b11 6
19
1>
1C
b11 G
#888400000000
0!
0*
09
0>
0C
#888410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#888420000000
0!
0*
09
0>
0C
#888430000000
1!
1*
b101 6
19
1>
1C
b101 G
#888440000000
0!
0*
09
0>
0C
#888450000000
1!
1*
b110 6
19
1>
1C
b110 G
#888460000000
0!
0*
09
0>
0C
#888470000000
1!
1*
b111 6
19
1>
1C
b111 G
#888480000000
0!
0*
09
0>
0C
#888490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#888500000000
0!
0*
09
0>
0C
#888510000000
1!
1*
b1 6
19
1>
1C
b1 G
#888520000000
0!
0*
09
0>
0C
#888530000000
1!
1*
b10 6
19
1>
1C
b10 G
#888540000000
0!
0*
09
0>
0C
#888550000000
1!
1*
b11 6
19
1>
1C
b11 G
#888560000000
0!
0*
09
0>
0C
#888570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#888580000000
0!
0*
09
0>
0C
#888590000000
1!
1*
b101 6
19
1>
1C
b101 G
#888600000000
0!
0*
09
0>
0C
#888610000000
1!
1*
b110 6
19
1>
1C
b110 G
#888620000000
0!
0*
09
0>
0C
#888630000000
1!
1*
b111 6
19
1>
1C
b111 G
#888640000000
0!
0*
09
0>
0C
#888650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#888660000000
0!
0*
09
0>
0C
#888670000000
1!
1*
b1 6
19
1>
1C
b1 G
#888680000000
0!
0*
09
0>
0C
#888690000000
1!
1*
b10 6
19
1>
1C
b10 G
#888700000000
0!
0*
09
0>
0C
#888710000000
1!
1*
b11 6
19
1>
1C
b11 G
#888720000000
0!
0*
09
0>
0C
#888730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#888740000000
0!
0*
09
0>
0C
#888750000000
1!
1*
b101 6
19
1>
1C
b101 G
#888760000000
0!
0*
09
0>
0C
#888770000000
1!
1*
b110 6
19
1>
1C
b110 G
#888780000000
0!
0*
09
0>
0C
#888790000000
1!
1*
b111 6
19
1>
1C
b111 G
#888800000000
0!
1"
0*
1+
09
1:
0>
0C
#888810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#888820000000
0!
0*
09
0>
0C
#888830000000
1!
1*
b1 6
19
1>
1C
b1 G
#888840000000
0!
0*
09
0>
0C
#888850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#888860000000
0!
0*
09
0>
0C
#888870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#888880000000
0!
0*
09
0>
0C
#888890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#888900000000
0!
0*
09
0>
0C
#888910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#888920000000
0!
0#
0*
0,
09
0>
0?
0C
#888930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#888940000000
0!
0*
09
0>
0C
#888950000000
1!
1*
19
1>
1C
#888960000000
0!
0*
09
0>
0C
#888970000000
1!
1*
19
1>
1C
#888980000000
0!
0*
09
0>
0C
#888990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#889000000000
0!
0*
09
0>
0C
#889010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#889020000000
0!
0*
09
0>
0C
#889030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#889040000000
0!
0*
09
0>
0C
#889050000000
1!
1*
b10 6
19
1>
1C
b10 G
#889060000000
0!
0*
09
0>
0C
#889070000000
1!
1*
b11 6
19
1>
1C
b11 G
#889080000000
0!
0*
09
0>
0C
#889090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#889100000000
0!
0*
09
0>
0C
#889110000000
1!
1*
b101 6
19
1>
1C
b101 G
#889120000000
0!
0*
09
0>
0C
#889130000000
1!
1*
b110 6
19
1>
1C
b110 G
#889140000000
0!
0*
09
0>
0C
#889150000000
1!
1*
b111 6
19
1>
1C
b111 G
#889160000000
0!
0*
09
0>
0C
#889170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#889180000000
0!
0*
09
0>
0C
#889190000000
1!
1*
b1 6
19
1>
1C
b1 G
#889200000000
0!
0*
09
0>
0C
#889210000000
1!
1*
b10 6
19
1>
1C
b10 G
#889220000000
0!
0*
09
0>
0C
#889230000000
1!
1*
b11 6
19
1>
1C
b11 G
#889240000000
0!
0*
09
0>
0C
#889250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#889260000000
0!
0*
09
0>
0C
#889270000000
1!
1*
b101 6
19
1>
1C
b101 G
#889280000000
0!
0*
09
0>
0C
#889290000000
1!
1*
b110 6
19
1>
1C
b110 G
#889300000000
0!
0*
09
0>
0C
#889310000000
1!
1*
b111 6
19
1>
1C
b111 G
#889320000000
0!
0*
09
0>
0C
#889330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#889340000000
0!
0*
09
0>
0C
#889350000000
1!
1*
b1 6
19
1>
1C
b1 G
#889360000000
0!
0*
09
0>
0C
#889370000000
1!
1*
b10 6
19
1>
1C
b10 G
#889380000000
0!
0*
09
0>
0C
#889390000000
1!
1*
b11 6
19
1>
1C
b11 G
#889400000000
0!
0*
09
0>
0C
#889410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#889420000000
0!
0*
09
0>
0C
#889430000000
1!
1*
b101 6
19
1>
1C
b101 G
#889440000000
0!
0*
09
0>
0C
#889450000000
1!
1*
b110 6
19
1>
1C
b110 G
#889460000000
0!
0*
09
0>
0C
#889470000000
1!
1*
b111 6
19
1>
1C
b111 G
#889480000000
0!
1"
0*
1+
09
1:
0>
0C
#889490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#889500000000
0!
0*
09
0>
0C
#889510000000
1!
1*
b1 6
19
1>
1C
b1 G
#889520000000
0!
0*
09
0>
0C
#889530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#889540000000
0!
0*
09
0>
0C
#889550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#889560000000
0!
0*
09
0>
0C
#889570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#889580000000
0!
0*
09
0>
0C
#889590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#889600000000
0!
0#
0*
0,
09
0>
0?
0C
#889610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#889620000000
0!
0*
09
0>
0C
#889630000000
1!
1*
19
1>
1C
#889640000000
0!
0*
09
0>
0C
#889650000000
1!
1*
19
1>
1C
#889660000000
0!
0*
09
0>
0C
#889670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#889680000000
0!
0*
09
0>
0C
#889690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#889700000000
0!
0*
09
0>
0C
#889710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#889720000000
0!
0*
09
0>
0C
#889730000000
1!
1*
b10 6
19
1>
1C
b10 G
#889740000000
0!
0*
09
0>
0C
#889750000000
1!
1*
b11 6
19
1>
1C
b11 G
#889760000000
0!
0*
09
0>
0C
#889770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#889780000000
0!
0*
09
0>
0C
#889790000000
1!
1*
b101 6
19
1>
1C
b101 G
#889800000000
0!
0*
09
0>
0C
#889810000000
1!
1*
b110 6
19
1>
1C
b110 G
#889820000000
0!
0*
09
0>
0C
#889830000000
1!
1*
b111 6
19
1>
1C
b111 G
#889840000000
0!
0*
09
0>
0C
#889850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#889860000000
0!
0*
09
0>
0C
#889870000000
1!
1*
b1 6
19
1>
1C
b1 G
#889880000000
0!
0*
09
0>
0C
#889890000000
1!
1*
b10 6
19
1>
1C
b10 G
#889900000000
0!
0*
09
0>
0C
#889910000000
1!
1*
b11 6
19
1>
1C
b11 G
#889920000000
0!
0*
09
0>
0C
#889930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#889940000000
0!
0*
09
0>
0C
#889950000000
1!
1*
b101 6
19
1>
1C
b101 G
#889960000000
0!
0*
09
0>
0C
#889970000000
1!
1*
b110 6
19
1>
1C
b110 G
#889980000000
0!
0*
09
0>
0C
#889990000000
1!
1*
b111 6
19
1>
1C
b111 G
#890000000000
0!
0*
09
0>
0C
#890010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#890020000000
0!
0*
09
0>
0C
#890030000000
1!
1*
b1 6
19
1>
1C
b1 G
#890040000000
0!
0*
09
0>
0C
#890050000000
1!
1*
b10 6
19
1>
1C
b10 G
#890060000000
0!
0*
09
0>
0C
#890070000000
1!
1*
b11 6
19
1>
1C
b11 G
#890080000000
0!
0*
09
0>
0C
#890090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#890100000000
0!
0*
09
0>
0C
#890110000000
1!
1*
b101 6
19
1>
1C
b101 G
#890120000000
0!
0*
09
0>
0C
#890130000000
1!
1*
b110 6
19
1>
1C
b110 G
#890140000000
0!
0*
09
0>
0C
#890150000000
1!
1*
b111 6
19
1>
1C
b111 G
#890160000000
0!
1"
0*
1+
09
1:
0>
0C
#890170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#890180000000
0!
0*
09
0>
0C
#890190000000
1!
1*
b1 6
19
1>
1C
b1 G
#890200000000
0!
0*
09
0>
0C
#890210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#890220000000
0!
0*
09
0>
0C
#890230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#890240000000
0!
0*
09
0>
0C
#890250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#890260000000
0!
0*
09
0>
0C
#890270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#890280000000
0!
0#
0*
0,
09
0>
0?
0C
#890290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#890300000000
0!
0*
09
0>
0C
#890310000000
1!
1*
19
1>
1C
#890320000000
0!
0*
09
0>
0C
#890330000000
1!
1*
19
1>
1C
#890340000000
0!
0*
09
0>
0C
#890350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#890360000000
0!
0*
09
0>
0C
#890370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#890380000000
0!
0*
09
0>
0C
#890390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#890400000000
0!
0*
09
0>
0C
#890410000000
1!
1*
b10 6
19
1>
1C
b10 G
#890420000000
0!
0*
09
0>
0C
#890430000000
1!
1*
b11 6
19
1>
1C
b11 G
#890440000000
0!
0*
09
0>
0C
#890450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#890460000000
0!
0*
09
0>
0C
#890470000000
1!
1*
b101 6
19
1>
1C
b101 G
#890480000000
0!
0*
09
0>
0C
#890490000000
1!
1*
b110 6
19
1>
1C
b110 G
#890500000000
0!
0*
09
0>
0C
#890510000000
1!
1*
b111 6
19
1>
1C
b111 G
#890520000000
0!
0*
09
0>
0C
#890530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#890540000000
0!
0*
09
0>
0C
#890550000000
1!
1*
b1 6
19
1>
1C
b1 G
#890560000000
0!
0*
09
0>
0C
#890570000000
1!
1*
b10 6
19
1>
1C
b10 G
#890580000000
0!
0*
09
0>
0C
#890590000000
1!
1*
b11 6
19
1>
1C
b11 G
#890600000000
0!
0*
09
0>
0C
#890610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#890620000000
0!
0*
09
0>
0C
#890630000000
1!
1*
b101 6
19
1>
1C
b101 G
#890640000000
0!
0*
09
0>
0C
#890650000000
1!
1*
b110 6
19
1>
1C
b110 G
#890660000000
0!
0*
09
0>
0C
#890670000000
1!
1*
b111 6
19
1>
1C
b111 G
#890680000000
0!
0*
09
0>
0C
#890690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#890700000000
0!
0*
09
0>
0C
#890710000000
1!
1*
b1 6
19
1>
1C
b1 G
#890720000000
0!
0*
09
0>
0C
#890730000000
1!
1*
b10 6
19
1>
1C
b10 G
#890740000000
0!
0*
09
0>
0C
#890750000000
1!
1*
b11 6
19
1>
1C
b11 G
#890760000000
0!
0*
09
0>
0C
#890770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#890780000000
0!
0*
09
0>
0C
#890790000000
1!
1*
b101 6
19
1>
1C
b101 G
#890800000000
0!
0*
09
0>
0C
#890810000000
1!
1*
b110 6
19
1>
1C
b110 G
#890820000000
0!
0*
09
0>
0C
#890830000000
1!
1*
b111 6
19
1>
1C
b111 G
#890840000000
0!
1"
0*
1+
09
1:
0>
0C
#890850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#890860000000
0!
0*
09
0>
0C
#890870000000
1!
1*
b1 6
19
1>
1C
b1 G
#890880000000
0!
0*
09
0>
0C
#890890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#890900000000
0!
0*
09
0>
0C
#890910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#890920000000
0!
0*
09
0>
0C
#890930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#890940000000
0!
0*
09
0>
0C
#890950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#890960000000
0!
0#
0*
0,
09
0>
0?
0C
#890970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#890980000000
0!
0*
09
0>
0C
#890990000000
1!
1*
19
1>
1C
#891000000000
0!
0*
09
0>
0C
#891010000000
1!
1*
19
1>
1C
#891020000000
0!
0*
09
0>
0C
#891030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#891040000000
0!
0*
09
0>
0C
#891050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#891060000000
0!
0*
09
0>
0C
#891070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#891080000000
0!
0*
09
0>
0C
#891090000000
1!
1*
b10 6
19
1>
1C
b10 G
#891100000000
0!
0*
09
0>
0C
#891110000000
1!
1*
b11 6
19
1>
1C
b11 G
#891120000000
0!
0*
09
0>
0C
#891130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#891140000000
0!
0*
09
0>
0C
#891150000000
1!
1*
b101 6
19
1>
1C
b101 G
#891160000000
0!
0*
09
0>
0C
#891170000000
1!
1*
b110 6
19
1>
1C
b110 G
#891180000000
0!
0*
09
0>
0C
#891190000000
1!
1*
b111 6
19
1>
1C
b111 G
#891200000000
0!
0*
09
0>
0C
#891210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#891220000000
0!
0*
09
0>
0C
#891230000000
1!
1*
b1 6
19
1>
1C
b1 G
#891240000000
0!
0*
09
0>
0C
#891250000000
1!
1*
b10 6
19
1>
1C
b10 G
#891260000000
0!
0*
09
0>
0C
#891270000000
1!
1*
b11 6
19
1>
1C
b11 G
#891280000000
0!
0*
09
0>
0C
#891290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#891300000000
0!
0*
09
0>
0C
#891310000000
1!
1*
b101 6
19
1>
1C
b101 G
#891320000000
0!
0*
09
0>
0C
#891330000000
1!
1*
b110 6
19
1>
1C
b110 G
#891340000000
0!
0*
09
0>
0C
#891350000000
1!
1*
b111 6
19
1>
1C
b111 G
#891360000000
0!
0*
09
0>
0C
#891370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#891380000000
0!
0*
09
0>
0C
#891390000000
1!
1*
b1 6
19
1>
1C
b1 G
#891400000000
0!
0*
09
0>
0C
#891410000000
1!
1*
b10 6
19
1>
1C
b10 G
#891420000000
0!
0*
09
0>
0C
#891430000000
1!
1*
b11 6
19
1>
1C
b11 G
#891440000000
0!
0*
09
0>
0C
#891450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#891460000000
0!
0*
09
0>
0C
#891470000000
1!
1*
b101 6
19
1>
1C
b101 G
#891480000000
0!
0*
09
0>
0C
#891490000000
1!
1*
b110 6
19
1>
1C
b110 G
#891500000000
0!
0*
09
0>
0C
#891510000000
1!
1*
b111 6
19
1>
1C
b111 G
#891520000000
0!
1"
0*
1+
09
1:
0>
0C
#891530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#891540000000
0!
0*
09
0>
0C
#891550000000
1!
1*
b1 6
19
1>
1C
b1 G
#891560000000
0!
0*
09
0>
0C
#891570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#891580000000
0!
0*
09
0>
0C
#891590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#891600000000
0!
0*
09
0>
0C
#891610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#891620000000
0!
0*
09
0>
0C
#891630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#891640000000
0!
0#
0*
0,
09
0>
0?
0C
#891650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#891660000000
0!
0*
09
0>
0C
#891670000000
1!
1*
19
1>
1C
#891680000000
0!
0*
09
0>
0C
#891690000000
1!
1*
19
1>
1C
#891700000000
0!
0*
09
0>
0C
#891710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#891720000000
0!
0*
09
0>
0C
#891730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#891740000000
0!
0*
09
0>
0C
#891750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#891760000000
0!
0*
09
0>
0C
#891770000000
1!
1*
b10 6
19
1>
1C
b10 G
#891780000000
0!
0*
09
0>
0C
#891790000000
1!
1*
b11 6
19
1>
1C
b11 G
#891800000000
0!
0*
09
0>
0C
#891810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#891820000000
0!
0*
09
0>
0C
#891830000000
1!
1*
b101 6
19
1>
1C
b101 G
#891840000000
0!
0*
09
0>
0C
#891850000000
1!
1*
b110 6
19
1>
1C
b110 G
#891860000000
0!
0*
09
0>
0C
#891870000000
1!
1*
b111 6
19
1>
1C
b111 G
#891880000000
0!
0*
09
0>
0C
#891890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#891900000000
0!
0*
09
0>
0C
#891910000000
1!
1*
b1 6
19
1>
1C
b1 G
#891920000000
0!
0*
09
0>
0C
#891930000000
1!
1*
b10 6
19
1>
1C
b10 G
#891940000000
0!
0*
09
0>
0C
#891950000000
1!
1*
b11 6
19
1>
1C
b11 G
#891960000000
0!
0*
09
0>
0C
#891970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#891980000000
0!
0*
09
0>
0C
#891990000000
1!
1*
b101 6
19
1>
1C
b101 G
#892000000000
0!
0*
09
0>
0C
#892010000000
1!
1*
b110 6
19
1>
1C
b110 G
#892020000000
0!
0*
09
0>
0C
#892030000000
1!
1*
b111 6
19
1>
1C
b111 G
#892040000000
0!
0*
09
0>
0C
#892050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#892060000000
0!
0*
09
0>
0C
#892070000000
1!
1*
b1 6
19
1>
1C
b1 G
#892080000000
0!
0*
09
0>
0C
#892090000000
1!
1*
b10 6
19
1>
1C
b10 G
#892100000000
0!
0*
09
0>
0C
#892110000000
1!
1*
b11 6
19
1>
1C
b11 G
#892120000000
0!
0*
09
0>
0C
#892130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#892140000000
0!
0*
09
0>
0C
#892150000000
1!
1*
b101 6
19
1>
1C
b101 G
#892160000000
0!
0*
09
0>
0C
#892170000000
1!
1*
b110 6
19
1>
1C
b110 G
#892180000000
0!
0*
09
0>
0C
#892190000000
1!
1*
b111 6
19
1>
1C
b111 G
#892200000000
0!
1"
0*
1+
09
1:
0>
0C
#892210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#892220000000
0!
0*
09
0>
0C
#892230000000
1!
1*
b1 6
19
1>
1C
b1 G
#892240000000
0!
0*
09
0>
0C
#892250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#892260000000
0!
0*
09
0>
0C
#892270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#892280000000
0!
0*
09
0>
0C
#892290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#892300000000
0!
0*
09
0>
0C
#892310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#892320000000
0!
0#
0*
0,
09
0>
0?
0C
#892330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#892340000000
0!
0*
09
0>
0C
#892350000000
1!
1*
19
1>
1C
#892360000000
0!
0*
09
0>
0C
#892370000000
1!
1*
19
1>
1C
#892380000000
0!
0*
09
0>
0C
#892390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#892400000000
0!
0*
09
0>
0C
#892410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#892420000000
0!
0*
09
0>
0C
#892430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#892440000000
0!
0*
09
0>
0C
#892450000000
1!
1*
b10 6
19
1>
1C
b10 G
#892460000000
0!
0*
09
0>
0C
#892470000000
1!
1*
b11 6
19
1>
1C
b11 G
#892480000000
0!
0*
09
0>
0C
#892490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#892500000000
0!
0*
09
0>
0C
#892510000000
1!
1*
b101 6
19
1>
1C
b101 G
#892520000000
0!
0*
09
0>
0C
#892530000000
1!
1*
b110 6
19
1>
1C
b110 G
#892540000000
0!
0*
09
0>
0C
#892550000000
1!
1*
b111 6
19
1>
1C
b111 G
#892560000000
0!
0*
09
0>
0C
#892570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#892580000000
0!
0*
09
0>
0C
#892590000000
1!
1*
b1 6
19
1>
1C
b1 G
#892600000000
0!
0*
09
0>
0C
#892610000000
1!
1*
b10 6
19
1>
1C
b10 G
#892620000000
0!
0*
09
0>
0C
#892630000000
1!
1*
b11 6
19
1>
1C
b11 G
#892640000000
0!
0*
09
0>
0C
#892650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#892660000000
0!
0*
09
0>
0C
#892670000000
1!
1*
b101 6
19
1>
1C
b101 G
#892680000000
0!
0*
09
0>
0C
#892690000000
1!
1*
b110 6
19
1>
1C
b110 G
#892700000000
0!
0*
09
0>
0C
#892710000000
1!
1*
b111 6
19
1>
1C
b111 G
#892720000000
0!
0*
09
0>
0C
#892730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#892740000000
0!
0*
09
0>
0C
#892750000000
1!
1*
b1 6
19
1>
1C
b1 G
#892760000000
0!
0*
09
0>
0C
#892770000000
1!
1*
b10 6
19
1>
1C
b10 G
#892780000000
0!
0*
09
0>
0C
#892790000000
1!
1*
b11 6
19
1>
1C
b11 G
#892800000000
0!
0*
09
0>
0C
#892810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#892820000000
0!
0*
09
0>
0C
#892830000000
1!
1*
b101 6
19
1>
1C
b101 G
#892840000000
0!
0*
09
0>
0C
#892850000000
1!
1*
b110 6
19
1>
1C
b110 G
#892860000000
0!
0*
09
0>
0C
#892870000000
1!
1*
b111 6
19
1>
1C
b111 G
#892880000000
0!
1"
0*
1+
09
1:
0>
0C
#892890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#892900000000
0!
0*
09
0>
0C
#892910000000
1!
1*
b1 6
19
1>
1C
b1 G
#892920000000
0!
0*
09
0>
0C
#892930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#892940000000
0!
0*
09
0>
0C
#892950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#892960000000
0!
0*
09
0>
0C
#892970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#892980000000
0!
0*
09
0>
0C
#892990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#893000000000
0!
0#
0*
0,
09
0>
0?
0C
#893010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#893020000000
0!
0*
09
0>
0C
#893030000000
1!
1*
19
1>
1C
#893040000000
0!
0*
09
0>
0C
#893050000000
1!
1*
19
1>
1C
#893060000000
0!
0*
09
0>
0C
#893070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#893080000000
0!
0*
09
0>
0C
#893090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#893100000000
0!
0*
09
0>
0C
#893110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#893120000000
0!
0*
09
0>
0C
#893130000000
1!
1*
b10 6
19
1>
1C
b10 G
#893140000000
0!
0*
09
0>
0C
#893150000000
1!
1*
b11 6
19
1>
1C
b11 G
#893160000000
0!
0*
09
0>
0C
#893170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#893180000000
0!
0*
09
0>
0C
#893190000000
1!
1*
b101 6
19
1>
1C
b101 G
#893200000000
0!
0*
09
0>
0C
#893210000000
1!
1*
b110 6
19
1>
1C
b110 G
#893220000000
0!
0*
09
0>
0C
#893230000000
1!
1*
b111 6
19
1>
1C
b111 G
#893240000000
0!
0*
09
0>
0C
#893250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#893260000000
0!
0*
09
0>
0C
#893270000000
1!
1*
b1 6
19
1>
1C
b1 G
#893280000000
0!
0*
09
0>
0C
#893290000000
1!
1*
b10 6
19
1>
1C
b10 G
#893300000000
0!
0*
09
0>
0C
#893310000000
1!
1*
b11 6
19
1>
1C
b11 G
#893320000000
0!
0*
09
0>
0C
#893330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#893340000000
0!
0*
09
0>
0C
#893350000000
1!
1*
b101 6
19
1>
1C
b101 G
#893360000000
0!
0*
09
0>
0C
#893370000000
1!
1*
b110 6
19
1>
1C
b110 G
#893380000000
0!
0*
09
0>
0C
#893390000000
1!
1*
b111 6
19
1>
1C
b111 G
#893400000000
0!
0*
09
0>
0C
#893410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#893420000000
0!
0*
09
0>
0C
#893430000000
1!
1*
b1 6
19
1>
1C
b1 G
#893440000000
0!
0*
09
0>
0C
#893450000000
1!
1*
b10 6
19
1>
1C
b10 G
#893460000000
0!
0*
09
0>
0C
#893470000000
1!
1*
b11 6
19
1>
1C
b11 G
#893480000000
0!
0*
09
0>
0C
#893490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#893500000000
0!
0*
09
0>
0C
#893510000000
1!
1*
b101 6
19
1>
1C
b101 G
#893520000000
0!
0*
09
0>
0C
#893530000000
1!
1*
b110 6
19
1>
1C
b110 G
#893540000000
0!
0*
09
0>
0C
#893550000000
1!
1*
b111 6
19
1>
1C
b111 G
#893560000000
0!
1"
0*
1+
09
1:
0>
0C
#893570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#893580000000
0!
0*
09
0>
0C
#893590000000
1!
1*
b1 6
19
1>
1C
b1 G
#893600000000
0!
0*
09
0>
0C
#893610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#893620000000
0!
0*
09
0>
0C
#893630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#893640000000
0!
0*
09
0>
0C
#893650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#893660000000
0!
0*
09
0>
0C
#893670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#893680000000
0!
0#
0*
0,
09
0>
0?
0C
#893690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#893700000000
0!
0*
09
0>
0C
#893710000000
1!
1*
19
1>
1C
#893720000000
0!
0*
09
0>
0C
#893730000000
1!
1*
19
1>
1C
#893740000000
0!
0*
09
0>
0C
#893750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#893760000000
0!
0*
09
0>
0C
#893770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#893780000000
0!
0*
09
0>
0C
#893790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#893800000000
0!
0*
09
0>
0C
#893810000000
1!
1*
b10 6
19
1>
1C
b10 G
#893820000000
0!
0*
09
0>
0C
#893830000000
1!
1*
b11 6
19
1>
1C
b11 G
#893840000000
0!
0*
09
0>
0C
#893850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#893860000000
0!
0*
09
0>
0C
#893870000000
1!
1*
b101 6
19
1>
1C
b101 G
#893880000000
0!
0*
09
0>
0C
#893890000000
1!
1*
b110 6
19
1>
1C
b110 G
#893900000000
0!
0*
09
0>
0C
#893910000000
1!
1*
b111 6
19
1>
1C
b111 G
#893920000000
0!
0*
09
0>
0C
#893930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#893940000000
0!
0*
09
0>
0C
#893950000000
1!
1*
b1 6
19
1>
1C
b1 G
#893960000000
0!
0*
09
0>
0C
#893970000000
1!
1*
b10 6
19
1>
1C
b10 G
#893980000000
0!
0*
09
0>
0C
#893990000000
1!
1*
b11 6
19
1>
1C
b11 G
#894000000000
0!
0*
09
0>
0C
#894010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#894020000000
0!
0*
09
0>
0C
#894030000000
1!
1*
b101 6
19
1>
1C
b101 G
#894040000000
0!
0*
09
0>
0C
#894050000000
1!
1*
b110 6
19
1>
1C
b110 G
#894060000000
0!
0*
09
0>
0C
#894070000000
1!
1*
b111 6
19
1>
1C
b111 G
#894080000000
0!
0*
09
0>
0C
#894090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#894100000000
0!
0*
09
0>
0C
#894110000000
1!
1*
b1 6
19
1>
1C
b1 G
#894120000000
0!
0*
09
0>
0C
#894130000000
1!
1*
b10 6
19
1>
1C
b10 G
#894140000000
0!
0*
09
0>
0C
#894150000000
1!
1*
b11 6
19
1>
1C
b11 G
#894160000000
0!
0*
09
0>
0C
#894170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#894180000000
0!
0*
09
0>
0C
#894190000000
1!
1*
b101 6
19
1>
1C
b101 G
#894200000000
0!
0*
09
0>
0C
#894210000000
1!
1*
b110 6
19
1>
1C
b110 G
#894220000000
0!
0*
09
0>
0C
#894230000000
1!
1*
b111 6
19
1>
1C
b111 G
#894240000000
0!
1"
0*
1+
09
1:
0>
0C
#894250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#894260000000
0!
0*
09
0>
0C
#894270000000
1!
1*
b1 6
19
1>
1C
b1 G
#894280000000
0!
0*
09
0>
0C
#894290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#894300000000
0!
0*
09
0>
0C
#894310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#894320000000
0!
0*
09
0>
0C
#894330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#894340000000
0!
0*
09
0>
0C
#894350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#894360000000
0!
0#
0*
0,
09
0>
0?
0C
#894370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#894380000000
0!
0*
09
0>
0C
#894390000000
1!
1*
19
1>
1C
#894400000000
0!
0*
09
0>
0C
#894410000000
1!
1*
19
1>
1C
#894420000000
0!
0*
09
0>
0C
#894430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#894440000000
0!
0*
09
0>
0C
#894450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#894460000000
0!
0*
09
0>
0C
#894470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#894480000000
0!
0*
09
0>
0C
#894490000000
1!
1*
b10 6
19
1>
1C
b10 G
#894500000000
0!
0*
09
0>
0C
#894510000000
1!
1*
b11 6
19
1>
1C
b11 G
#894520000000
0!
0*
09
0>
0C
#894530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#894540000000
0!
0*
09
0>
0C
#894550000000
1!
1*
b101 6
19
1>
1C
b101 G
#894560000000
0!
0*
09
0>
0C
#894570000000
1!
1*
b110 6
19
1>
1C
b110 G
#894580000000
0!
0*
09
0>
0C
#894590000000
1!
1*
b111 6
19
1>
1C
b111 G
#894600000000
0!
0*
09
0>
0C
#894610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#894620000000
0!
0*
09
0>
0C
#894630000000
1!
1*
b1 6
19
1>
1C
b1 G
#894640000000
0!
0*
09
0>
0C
#894650000000
1!
1*
b10 6
19
1>
1C
b10 G
#894660000000
0!
0*
09
0>
0C
#894670000000
1!
1*
b11 6
19
1>
1C
b11 G
#894680000000
0!
0*
09
0>
0C
#894690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#894700000000
0!
0*
09
0>
0C
#894710000000
1!
1*
b101 6
19
1>
1C
b101 G
#894720000000
0!
0*
09
0>
0C
#894730000000
1!
1*
b110 6
19
1>
1C
b110 G
#894740000000
0!
0*
09
0>
0C
#894750000000
1!
1*
b111 6
19
1>
1C
b111 G
#894760000000
0!
0*
09
0>
0C
#894770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#894780000000
0!
0*
09
0>
0C
#894790000000
1!
1*
b1 6
19
1>
1C
b1 G
#894800000000
0!
0*
09
0>
0C
#894810000000
1!
1*
b10 6
19
1>
1C
b10 G
#894820000000
0!
0*
09
0>
0C
#894830000000
1!
1*
b11 6
19
1>
1C
b11 G
#894840000000
0!
0*
09
0>
0C
#894850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#894860000000
0!
0*
09
0>
0C
#894870000000
1!
1*
b101 6
19
1>
1C
b101 G
#894880000000
0!
0*
09
0>
0C
#894890000000
1!
1*
b110 6
19
1>
1C
b110 G
#894900000000
0!
0*
09
0>
0C
#894910000000
1!
1*
b111 6
19
1>
1C
b111 G
#894920000000
0!
1"
0*
1+
09
1:
0>
0C
#894930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#894940000000
0!
0*
09
0>
0C
#894950000000
1!
1*
b1 6
19
1>
1C
b1 G
#894960000000
0!
0*
09
0>
0C
#894970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#894980000000
0!
0*
09
0>
0C
#894990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#895000000000
0!
0*
09
0>
0C
#895010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#895020000000
0!
0*
09
0>
0C
#895030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#895040000000
0!
0#
0*
0,
09
0>
0?
0C
#895050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#895060000000
0!
0*
09
0>
0C
#895070000000
1!
1*
19
1>
1C
#895080000000
0!
0*
09
0>
0C
#895090000000
1!
1*
19
1>
1C
#895100000000
0!
0*
09
0>
0C
#895110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#895120000000
0!
0*
09
0>
0C
#895130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#895140000000
0!
0*
09
0>
0C
#895150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#895160000000
0!
0*
09
0>
0C
#895170000000
1!
1*
b10 6
19
1>
1C
b10 G
#895180000000
0!
0*
09
0>
0C
#895190000000
1!
1*
b11 6
19
1>
1C
b11 G
#895200000000
0!
0*
09
0>
0C
#895210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#895220000000
0!
0*
09
0>
0C
#895230000000
1!
1*
b101 6
19
1>
1C
b101 G
#895240000000
0!
0*
09
0>
0C
#895250000000
1!
1*
b110 6
19
1>
1C
b110 G
#895260000000
0!
0*
09
0>
0C
#895270000000
1!
1*
b111 6
19
1>
1C
b111 G
#895280000000
0!
0*
09
0>
0C
#895290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#895300000000
0!
0*
09
0>
0C
#895310000000
1!
1*
b1 6
19
1>
1C
b1 G
#895320000000
0!
0*
09
0>
0C
#895330000000
1!
1*
b10 6
19
1>
1C
b10 G
#895340000000
0!
0*
09
0>
0C
#895350000000
1!
1*
b11 6
19
1>
1C
b11 G
#895360000000
0!
0*
09
0>
0C
#895370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#895380000000
0!
0*
09
0>
0C
#895390000000
1!
1*
b101 6
19
1>
1C
b101 G
#895400000000
0!
0*
09
0>
0C
#895410000000
1!
1*
b110 6
19
1>
1C
b110 G
#895420000000
0!
0*
09
0>
0C
#895430000000
1!
1*
b111 6
19
1>
1C
b111 G
#895440000000
0!
0*
09
0>
0C
#895450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#895460000000
0!
0*
09
0>
0C
#895470000000
1!
1*
b1 6
19
1>
1C
b1 G
#895480000000
0!
0*
09
0>
0C
#895490000000
1!
1*
b10 6
19
1>
1C
b10 G
#895500000000
0!
0*
09
0>
0C
#895510000000
1!
1*
b11 6
19
1>
1C
b11 G
#895520000000
0!
0*
09
0>
0C
#895530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#895540000000
0!
0*
09
0>
0C
#895550000000
1!
1*
b101 6
19
1>
1C
b101 G
#895560000000
0!
0*
09
0>
0C
#895570000000
1!
1*
b110 6
19
1>
1C
b110 G
#895580000000
0!
0*
09
0>
0C
#895590000000
1!
1*
b111 6
19
1>
1C
b111 G
#895600000000
0!
1"
0*
1+
09
1:
0>
0C
#895610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#895620000000
0!
0*
09
0>
0C
#895630000000
1!
1*
b1 6
19
1>
1C
b1 G
#895640000000
0!
0*
09
0>
0C
#895650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#895660000000
0!
0*
09
0>
0C
#895670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#895680000000
0!
0*
09
0>
0C
#895690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#895700000000
0!
0*
09
0>
0C
#895710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#895720000000
0!
0#
0*
0,
09
0>
0?
0C
#895730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#895740000000
0!
0*
09
0>
0C
#895750000000
1!
1*
19
1>
1C
#895760000000
0!
0*
09
0>
0C
#895770000000
1!
1*
19
1>
1C
#895780000000
0!
0*
09
0>
0C
#895790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#895800000000
0!
0*
09
0>
0C
#895810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#895820000000
0!
0*
09
0>
0C
#895830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#895840000000
0!
0*
09
0>
0C
#895850000000
1!
1*
b10 6
19
1>
1C
b10 G
#895860000000
0!
0*
09
0>
0C
#895870000000
1!
1*
b11 6
19
1>
1C
b11 G
#895880000000
0!
0*
09
0>
0C
#895890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#895900000000
0!
0*
09
0>
0C
#895910000000
1!
1*
b101 6
19
1>
1C
b101 G
#895920000000
0!
0*
09
0>
0C
#895930000000
1!
1*
b110 6
19
1>
1C
b110 G
#895940000000
0!
0*
09
0>
0C
#895950000000
1!
1*
b111 6
19
1>
1C
b111 G
#895960000000
0!
0*
09
0>
0C
#895970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#895980000000
0!
0*
09
0>
0C
#895990000000
1!
1*
b1 6
19
1>
1C
b1 G
#896000000000
0!
0*
09
0>
0C
#896010000000
1!
1*
b10 6
19
1>
1C
b10 G
#896020000000
0!
0*
09
0>
0C
#896030000000
1!
1*
b11 6
19
1>
1C
b11 G
#896040000000
0!
0*
09
0>
0C
#896050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#896060000000
0!
0*
09
0>
0C
#896070000000
1!
1*
b101 6
19
1>
1C
b101 G
#896080000000
0!
0*
09
0>
0C
#896090000000
1!
1*
b110 6
19
1>
1C
b110 G
#896100000000
0!
0*
09
0>
0C
#896110000000
1!
1*
b111 6
19
1>
1C
b111 G
#896120000000
0!
0*
09
0>
0C
#896130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#896140000000
0!
0*
09
0>
0C
#896150000000
1!
1*
b1 6
19
1>
1C
b1 G
#896160000000
0!
0*
09
0>
0C
#896170000000
1!
1*
b10 6
19
1>
1C
b10 G
#896180000000
0!
0*
09
0>
0C
#896190000000
1!
1*
b11 6
19
1>
1C
b11 G
#896200000000
0!
0*
09
0>
0C
#896210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#896220000000
0!
0*
09
0>
0C
#896230000000
1!
1*
b101 6
19
1>
1C
b101 G
#896240000000
0!
0*
09
0>
0C
#896250000000
1!
1*
b110 6
19
1>
1C
b110 G
#896260000000
0!
0*
09
0>
0C
#896270000000
1!
1*
b111 6
19
1>
1C
b111 G
#896280000000
0!
1"
0*
1+
09
1:
0>
0C
#896290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#896300000000
0!
0*
09
0>
0C
#896310000000
1!
1*
b1 6
19
1>
1C
b1 G
#896320000000
0!
0*
09
0>
0C
#896330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#896340000000
0!
0*
09
0>
0C
#896350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#896360000000
0!
0*
09
0>
0C
#896370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#896380000000
0!
0*
09
0>
0C
#896390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#896400000000
0!
0#
0*
0,
09
0>
0?
0C
#896410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#896420000000
0!
0*
09
0>
0C
#896430000000
1!
1*
19
1>
1C
#896440000000
0!
0*
09
0>
0C
#896450000000
1!
1*
19
1>
1C
#896460000000
0!
0*
09
0>
0C
#896470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#896480000000
0!
0*
09
0>
0C
#896490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#896500000000
0!
0*
09
0>
0C
#896510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#896520000000
0!
0*
09
0>
0C
#896530000000
1!
1*
b10 6
19
1>
1C
b10 G
#896540000000
0!
0*
09
0>
0C
#896550000000
1!
1*
b11 6
19
1>
1C
b11 G
#896560000000
0!
0*
09
0>
0C
#896570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#896580000000
0!
0*
09
0>
0C
#896590000000
1!
1*
b101 6
19
1>
1C
b101 G
#896600000000
0!
0*
09
0>
0C
#896610000000
1!
1*
b110 6
19
1>
1C
b110 G
#896620000000
0!
0*
09
0>
0C
#896630000000
1!
1*
b111 6
19
1>
1C
b111 G
#896640000000
0!
0*
09
0>
0C
#896650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#896660000000
0!
0*
09
0>
0C
#896670000000
1!
1*
b1 6
19
1>
1C
b1 G
#896680000000
0!
0*
09
0>
0C
#896690000000
1!
1*
b10 6
19
1>
1C
b10 G
#896700000000
0!
0*
09
0>
0C
#896710000000
1!
1*
b11 6
19
1>
1C
b11 G
#896720000000
0!
0*
09
0>
0C
#896730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#896740000000
0!
0*
09
0>
0C
#896750000000
1!
1*
b101 6
19
1>
1C
b101 G
#896760000000
0!
0*
09
0>
0C
#896770000000
1!
1*
b110 6
19
1>
1C
b110 G
#896780000000
0!
0*
09
0>
0C
#896790000000
1!
1*
b111 6
19
1>
1C
b111 G
#896800000000
0!
0*
09
0>
0C
#896810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#896820000000
0!
0*
09
0>
0C
#896830000000
1!
1*
b1 6
19
1>
1C
b1 G
#896840000000
0!
0*
09
0>
0C
#896850000000
1!
1*
b10 6
19
1>
1C
b10 G
#896860000000
0!
0*
09
0>
0C
#896870000000
1!
1*
b11 6
19
1>
1C
b11 G
#896880000000
0!
0*
09
0>
0C
#896890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#896900000000
0!
0*
09
0>
0C
#896910000000
1!
1*
b101 6
19
1>
1C
b101 G
#896920000000
0!
0*
09
0>
0C
#896930000000
1!
1*
b110 6
19
1>
1C
b110 G
#896940000000
0!
0*
09
0>
0C
#896950000000
1!
1*
b111 6
19
1>
1C
b111 G
#896960000000
0!
1"
0*
1+
09
1:
0>
0C
#896970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#896980000000
0!
0*
09
0>
0C
#896990000000
1!
1*
b1 6
19
1>
1C
b1 G
#897000000000
0!
0*
09
0>
0C
#897010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#897020000000
0!
0*
09
0>
0C
#897030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#897040000000
0!
0*
09
0>
0C
#897050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#897060000000
0!
0*
09
0>
0C
#897070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#897080000000
0!
0#
0*
0,
09
0>
0?
0C
#897090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#897100000000
0!
0*
09
0>
0C
#897110000000
1!
1*
19
1>
1C
#897120000000
0!
0*
09
0>
0C
#897130000000
1!
1*
19
1>
1C
#897140000000
0!
0*
09
0>
0C
#897150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#897160000000
0!
0*
09
0>
0C
#897170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#897180000000
0!
0*
09
0>
0C
#897190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#897200000000
0!
0*
09
0>
0C
#897210000000
1!
1*
b10 6
19
1>
1C
b10 G
#897220000000
0!
0*
09
0>
0C
#897230000000
1!
1*
b11 6
19
1>
1C
b11 G
#897240000000
0!
0*
09
0>
0C
#897250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#897260000000
0!
0*
09
0>
0C
#897270000000
1!
1*
b101 6
19
1>
1C
b101 G
#897280000000
0!
0*
09
0>
0C
#897290000000
1!
1*
b110 6
19
1>
1C
b110 G
#897300000000
0!
0*
09
0>
0C
#897310000000
1!
1*
b111 6
19
1>
1C
b111 G
#897320000000
0!
0*
09
0>
0C
#897330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#897340000000
0!
0*
09
0>
0C
#897350000000
1!
1*
b1 6
19
1>
1C
b1 G
#897360000000
0!
0*
09
0>
0C
#897370000000
1!
1*
b10 6
19
1>
1C
b10 G
#897380000000
0!
0*
09
0>
0C
#897390000000
1!
1*
b11 6
19
1>
1C
b11 G
#897400000000
0!
0*
09
0>
0C
#897410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#897420000000
0!
0*
09
0>
0C
#897430000000
1!
1*
b101 6
19
1>
1C
b101 G
#897440000000
0!
0*
09
0>
0C
#897450000000
1!
1*
b110 6
19
1>
1C
b110 G
#897460000000
0!
0*
09
0>
0C
#897470000000
1!
1*
b111 6
19
1>
1C
b111 G
#897480000000
0!
0*
09
0>
0C
#897490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#897500000000
0!
0*
09
0>
0C
#897510000000
1!
1*
b1 6
19
1>
1C
b1 G
#897520000000
0!
0*
09
0>
0C
#897530000000
1!
1*
b10 6
19
1>
1C
b10 G
#897540000000
0!
0*
09
0>
0C
#897550000000
1!
1*
b11 6
19
1>
1C
b11 G
#897560000000
0!
0*
09
0>
0C
#897570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#897580000000
0!
0*
09
0>
0C
#897590000000
1!
1*
b101 6
19
1>
1C
b101 G
#897600000000
0!
0*
09
0>
0C
#897610000000
1!
1*
b110 6
19
1>
1C
b110 G
#897620000000
0!
0*
09
0>
0C
#897630000000
1!
1*
b111 6
19
1>
1C
b111 G
#897640000000
0!
1"
0*
1+
09
1:
0>
0C
#897650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#897660000000
0!
0*
09
0>
0C
#897670000000
1!
1*
b1 6
19
1>
1C
b1 G
#897680000000
0!
0*
09
0>
0C
#897690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#897700000000
0!
0*
09
0>
0C
#897710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#897720000000
0!
0*
09
0>
0C
#897730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#897740000000
0!
0*
09
0>
0C
#897750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#897760000000
0!
0#
0*
0,
09
0>
0?
0C
#897770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#897780000000
0!
0*
09
0>
0C
#897790000000
1!
1*
19
1>
1C
#897800000000
0!
0*
09
0>
0C
#897810000000
1!
1*
19
1>
1C
#897820000000
0!
0*
09
0>
0C
#897830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#897840000000
0!
0*
09
0>
0C
#897850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#897860000000
0!
0*
09
0>
0C
#897870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#897880000000
0!
0*
09
0>
0C
#897890000000
1!
1*
b10 6
19
1>
1C
b10 G
#897900000000
0!
0*
09
0>
0C
#897910000000
1!
1*
b11 6
19
1>
1C
b11 G
#897920000000
0!
0*
09
0>
0C
#897930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#897940000000
0!
0*
09
0>
0C
#897950000000
1!
1*
b101 6
19
1>
1C
b101 G
#897960000000
0!
0*
09
0>
0C
#897970000000
1!
1*
b110 6
19
1>
1C
b110 G
#897980000000
0!
0*
09
0>
0C
#897990000000
1!
1*
b111 6
19
1>
1C
b111 G
#898000000000
0!
0*
09
0>
0C
#898010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#898020000000
0!
0*
09
0>
0C
#898030000000
1!
1*
b1 6
19
1>
1C
b1 G
#898040000000
0!
0*
09
0>
0C
#898050000000
1!
1*
b10 6
19
1>
1C
b10 G
#898060000000
0!
0*
09
0>
0C
#898070000000
1!
1*
b11 6
19
1>
1C
b11 G
#898080000000
0!
0*
09
0>
0C
#898090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#898100000000
0!
0*
09
0>
0C
#898110000000
1!
1*
b101 6
19
1>
1C
b101 G
#898120000000
0!
0*
09
0>
0C
#898130000000
1!
1*
b110 6
19
1>
1C
b110 G
#898140000000
0!
0*
09
0>
0C
#898150000000
1!
1*
b111 6
19
1>
1C
b111 G
#898160000000
0!
0*
09
0>
0C
#898170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#898180000000
0!
0*
09
0>
0C
#898190000000
1!
1*
b1 6
19
1>
1C
b1 G
#898200000000
0!
0*
09
0>
0C
#898210000000
1!
1*
b10 6
19
1>
1C
b10 G
#898220000000
0!
0*
09
0>
0C
#898230000000
1!
1*
b11 6
19
1>
1C
b11 G
#898240000000
0!
0*
09
0>
0C
#898250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#898260000000
0!
0*
09
0>
0C
#898270000000
1!
1*
b101 6
19
1>
1C
b101 G
#898280000000
0!
0*
09
0>
0C
#898290000000
1!
1*
b110 6
19
1>
1C
b110 G
#898300000000
0!
0*
09
0>
0C
#898310000000
1!
1*
b111 6
19
1>
1C
b111 G
#898320000000
0!
1"
0*
1+
09
1:
0>
0C
#898330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#898340000000
0!
0*
09
0>
0C
#898350000000
1!
1*
b1 6
19
1>
1C
b1 G
#898360000000
0!
0*
09
0>
0C
#898370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#898380000000
0!
0*
09
0>
0C
#898390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#898400000000
0!
0*
09
0>
0C
#898410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#898420000000
0!
0*
09
0>
0C
#898430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#898440000000
0!
0#
0*
0,
09
0>
0?
0C
#898450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#898460000000
0!
0*
09
0>
0C
#898470000000
1!
1*
19
1>
1C
#898480000000
0!
0*
09
0>
0C
#898490000000
1!
1*
19
1>
1C
#898500000000
0!
0*
09
0>
0C
#898510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#898520000000
0!
0*
09
0>
0C
#898530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#898540000000
0!
0*
09
0>
0C
#898550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#898560000000
0!
0*
09
0>
0C
#898570000000
1!
1*
b10 6
19
1>
1C
b10 G
#898580000000
0!
0*
09
0>
0C
#898590000000
1!
1*
b11 6
19
1>
1C
b11 G
#898600000000
0!
0*
09
0>
0C
#898610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#898620000000
0!
0*
09
0>
0C
#898630000000
1!
1*
b101 6
19
1>
1C
b101 G
#898640000000
0!
0*
09
0>
0C
#898650000000
1!
1*
b110 6
19
1>
1C
b110 G
#898660000000
0!
0*
09
0>
0C
#898670000000
1!
1*
b111 6
19
1>
1C
b111 G
#898680000000
0!
0*
09
0>
0C
#898690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#898700000000
0!
0*
09
0>
0C
#898710000000
1!
1*
b1 6
19
1>
1C
b1 G
#898720000000
0!
0*
09
0>
0C
#898730000000
1!
1*
b10 6
19
1>
1C
b10 G
#898740000000
0!
0*
09
0>
0C
#898750000000
1!
1*
b11 6
19
1>
1C
b11 G
#898760000000
0!
0*
09
0>
0C
#898770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#898780000000
0!
0*
09
0>
0C
#898790000000
1!
1*
b101 6
19
1>
1C
b101 G
#898800000000
0!
0*
09
0>
0C
#898810000000
1!
1*
b110 6
19
1>
1C
b110 G
#898820000000
0!
0*
09
0>
0C
#898830000000
1!
1*
b111 6
19
1>
1C
b111 G
#898840000000
0!
0*
09
0>
0C
#898850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#898860000000
0!
0*
09
0>
0C
#898870000000
1!
1*
b1 6
19
1>
1C
b1 G
#898880000000
0!
0*
09
0>
0C
#898890000000
1!
1*
b10 6
19
1>
1C
b10 G
#898900000000
0!
0*
09
0>
0C
#898910000000
1!
1*
b11 6
19
1>
1C
b11 G
#898920000000
0!
0*
09
0>
0C
#898930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#898940000000
0!
0*
09
0>
0C
#898950000000
1!
1*
b101 6
19
1>
1C
b101 G
#898960000000
0!
0*
09
0>
0C
#898970000000
1!
1*
b110 6
19
1>
1C
b110 G
#898980000000
0!
0*
09
0>
0C
#898990000000
1!
1*
b111 6
19
1>
1C
b111 G
#899000000000
0!
1"
0*
1+
09
1:
0>
0C
#899010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#899020000000
0!
0*
09
0>
0C
#899030000000
1!
1*
b1 6
19
1>
1C
b1 G
#899040000000
0!
0*
09
0>
0C
#899050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#899060000000
0!
0*
09
0>
0C
#899070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#899080000000
0!
0*
09
0>
0C
#899090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#899100000000
0!
0*
09
0>
0C
#899110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#899120000000
0!
0#
0*
0,
09
0>
0?
0C
#899130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#899140000000
0!
0*
09
0>
0C
#899150000000
1!
1*
19
1>
1C
#899160000000
0!
0*
09
0>
0C
#899170000000
1!
1*
19
1>
1C
#899180000000
0!
0*
09
0>
0C
#899190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#899200000000
0!
0*
09
0>
0C
#899210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#899220000000
0!
0*
09
0>
0C
#899230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#899240000000
0!
0*
09
0>
0C
#899250000000
1!
1*
b10 6
19
1>
1C
b10 G
#899260000000
0!
0*
09
0>
0C
#899270000000
1!
1*
b11 6
19
1>
1C
b11 G
#899280000000
0!
0*
09
0>
0C
#899290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#899300000000
0!
0*
09
0>
0C
#899310000000
1!
1*
b101 6
19
1>
1C
b101 G
#899320000000
0!
0*
09
0>
0C
#899330000000
1!
1*
b110 6
19
1>
1C
b110 G
#899340000000
0!
0*
09
0>
0C
#899350000000
1!
1*
b111 6
19
1>
1C
b111 G
#899360000000
0!
0*
09
0>
0C
#899370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#899380000000
0!
0*
09
0>
0C
#899390000000
1!
1*
b1 6
19
1>
1C
b1 G
#899400000000
0!
0*
09
0>
0C
#899410000000
1!
1*
b10 6
19
1>
1C
b10 G
#899420000000
0!
0*
09
0>
0C
#899430000000
1!
1*
b11 6
19
1>
1C
b11 G
#899440000000
0!
0*
09
0>
0C
#899450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#899460000000
0!
0*
09
0>
0C
#899470000000
1!
1*
b101 6
19
1>
1C
b101 G
#899480000000
0!
0*
09
0>
0C
#899490000000
1!
1*
b110 6
19
1>
1C
b110 G
#899500000000
0!
0*
09
0>
0C
#899510000000
1!
1*
b111 6
19
1>
1C
b111 G
#899520000000
0!
0*
09
0>
0C
#899530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#899540000000
0!
0*
09
0>
0C
#899550000000
1!
1*
b1 6
19
1>
1C
b1 G
#899560000000
0!
0*
09
0>
0C
#899570000000
1!
1*
b10 6
19
1>
1C
b10 G
#899580000000
0!
0*
09
0>
0C
#899590000000
1!
1*
b11 6
19
1>
1C
b11 G
#899600000000
0!
0*
09
0>
0C
#899610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#899620000000
0!
0*
09
0>
0C
#899630000000
1!
1*
b101 6
19
1>
1C
b101 G
#899640000000
0!
0*
09
0>
0C
#899650000000
1!
1*
b110 6
19
1>
1C
b110 G
#899660000000
0!
0*
09
0>
0C
#899670000000
1!
1*
b111 6
19
1>
1C
b111 G
#899680000000
0!
1"
0*
1+
09
1:
0>
0C
#899690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#899700000000
0!
0*
09
0>
0C
#899710000000
1!
1*
b1 6
19
1>
1C
b1 G
#899720000000
0!
0*
09
0>
0C
#899730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#899740000000
0!
0*
09
0>
0C
#899750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#899760000000
0!
0*
09
0>
0C
#899770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#899780000000
0!
0*
09
0>
0C
#899790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#899800000000
0!
0#
0*
0,
09
0>
0?
0C
#899810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#899820000000
0!
0*
09
0>
0C
#899830000000
1!
1*
19
1>
1C
#899840000000
0!
0*
09
0>
0C
#899850000000
1!
1*
19
1>
1C
#899860000000
0!
0*
09
0>
0C
#899870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#899880000000
0!
0*
09
0>
0C
#899890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#899900000000
0!
0*
09
0>
0C
#899910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#899920000000
0!
0*
09
0>
0C
#899930000000
1!
1*
b10 6
19
1>
1C
b10 G
#899940000000
0!
0*
09
0>
0C
#899950000000
1!
1*
b11 6
19
1>
1C
b11 G
#899960000000
0!
0*
09
0>
0C
#899970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#899980000000
0!
0*
09
0>
0C
#899990000000
1!
1*
b101 6
19
1>
1C
b101 G
#900000000000
0!
0*
09
0>
0C
#900010000000
1!
1*
b110 6
19
1>
1C
b110 G
#900020000000
0!
0*
09
0>
0C
#900030000000
1!
1*
b111 6
19
1>
1C
b111 G
#900040000000
0!
0*
09
0>
0C
#900050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#900060000000
0!
0*
09
0>
0C
#900070000000
1!
1*
b1 6
19
1>
1C
b1 G
#900080000000
0!
0*
09
0>
0C
#900090000000
1!
1*
b10 6
19
1>
1C
b10 G
#900100000000
0!
0*
09
0>
0C
#900110000000
1!
1*
b11 6
19
1>
1C
b11 G
#900120000000
0!
0*
09
0>
0C
#900130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#900140000000
0!
0*
09
0>
0C
#900150000000
1!
1*
b101 6
19
1>
1C
b101 G
#900160000000
0!
0*
09
0>
0C
#900170000000
1!
1*
b110 6
19
1>
1C
b110 G
#900180000000
0!
0*
09
0>
0C
#900190000000
1!
1*
b111 6
19
1>
1C
b111 G
#900200000000
0!
0*
09
0>
0C
#900210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#900220000000
0!
0*
09
0>
0C
#900230000000
1!
1*
b1 6
19
1>
1C
b1 G
#900240000000
0!
0*
09
0>
0C
#900250000000
1!
1*
b10 6
19
1>
1C
b10 G
#900260000000
0!
0*
09
0>
0C
#900270000000
1!
1*
b11 6
19
1>
1C
b11 G
#900280000000
0!
0*
09
0>
0C
#900290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#900300000000
0!
0*
09
0>
0C
#900310000000
1!
1*
b101 6
19
1>
1C
b101 G
#900320000000
0!
0*
09
0>
0C
#900330000000
1!
1*
b110 6
19
1>
1C
b110 G
#900340000000
0!
0*
09
0>
0C
#900350000000
1!
1*
b111 6
19
1>
1C
b111 G
#900360000000
0!
1"
0*
1+
09
1:
0>
0C
#900370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#900380000000
0!
0*
09
0>
0C
#900390000000
1!
1*
b1 6
19
1>
1C
b1 G
#900400000000
0!
0*
09
0>
0C
#900410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#900420000000
0!
0*
09
0>
0C
#900430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#900440000000
0!
0*
09
0>
0C
#900450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#900460000000
0!
0*
09
0>
0C
#900470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#900480000000
0!
0#
0*
0,
09
0>
0?
0C
#900490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#900500000000
0!
0*
09
0>
0C
#900510000000
1!
1*
19
1>
1C
#900520000000
0!
0*
09
0>
0C
#900530000000
1!
1*
19
1>
1C
#900540000000
0!
0*
09
0>
0C
#900550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#900560000000
0!
0*
09
0>
0C
#900570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#900580000000
0!
0*
09
0>
0C
#900590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#900600000000
0!
0*
09
0>
0C
#900610000000
1!
1*
b10 6
19
1>
1C
b10 G
#900620000000
0!
0*
09
0>
0C
#900630000000
1!
1*
b11 6
19
1>
1C
b11 G
#900640000000
0!
0*
09
0>
0C
#900650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#900660000000
0!
0*
09
0>
0C
#900670000000
1!
1*
b101 6
19
1>
1C
b101 G
#900680000000
0!
0*
09
0>
0C
#900690000000
1!
1*
b110 6
19
1>
1C
b110 G
#900700000000
0!
0*
09
0>
0C
#900710000000
1!
1*
b111 6
19
1>
1C
b111 G
#900720000000
0!
0*
09
0>
0C
#900730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#900740000000
0!
0*
09
0>
0C
#900750000000
1!
1*
b1 6
19
1>
1C
b1 G
#900760000000
0!
0*
09
0>
0C
#900770000000
1!
1*
b10 6
19
1>
1C
b10 G
#900780000000
0!
0*
09
0>
0C
#900790000000
1!
1*
b11 6
19
1>
1C
b11 G
#900800000000
0!
0*
09
0>
0C
#900810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#900820000000
0!
0*
09
0>
0C
#900830000000
1!
1*
b101 6
19
1>
1C
b101 G
#900840000000
0!
0*
09
0>
0C
#900850000000
1!
1*
b110 6
19
1>
1C
b110 G
#900860000000
0!
0*
09
0>
0C
#900870000000
1!
1*
b111 6
19
1>
1C
b111 G
#900880000000
0!
0*
09
0>
0C
#900890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#900900000000
0!
0*
09
0>
0C
#900910000000
1!
1*
b1 6
19
1>
1C
b1 G
#900920000000
0!
0*
09
0>
0C
#900930000000
1!
1*
b10 6
19
1>
1C
b10 G
#900940000000
0!
0*
09
0>
0C
#900950000000
1!
1*
b11 6
19
1>
1C
b11 G
#900960000000
0!
0*
09
0>
0C
#900970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#900980000000
0!
0*
09
0>
0C
#900990000000
1!
1*
b101 6
19
1>
1C
b101 G
#901000000000
0!
0*
09
0>
0C
#901010000000
1!
1*
b110 6
19
1>
1C
b110 G
#901020000000
0!
0*
09
0>
0C
#901030000000
1!
1*
b111 6
19
1>
1C
b111 G
#901040000000
0!
1"
0*
1+
09
1:
0>
0C
#901050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#901060000000
0!
0*
09
0>
0C
#901070000000
1!
1*
b1 6
19
1>
1C
b1 G
#901080000000
0!
0*
09
0>
0C
#901090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#901100000000
0!
0*
09
0>
0C
#901110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#901120000000
0!
0*
09
0>
0C
#901130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#901140000000
0!
0*
09
0>
0C
#901150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#901160000000
0!
0#
0*
0,
09
0>
0?
0C
#901170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#901180000000
0!
0*
09
0>
0C
#901190000000
1!
1*
19
1>
1C
#901200000000
0!
0*
09
0>
0C
#901210000000
1!
1*
19
1>
1C
#901220000000
0!
0*
09
0>
0C
#901230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#901240000000
0!
0*
09
0>
0C
#901250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#901260000000
0!
0*
09
0>
0C
#901270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#901280000000
0!
0*
09
0>
0C
#901290000000
1!
1*
b10 6
19
1>
1C
b10 G
#901300000000
0!
0*
09
0>
0C
#901310000000
1!
1*
b11 6
19
1>
1C
b11 G
#901320000000
0!
0*
09
0>
0C
#901330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#901340000000
0!
0*
09
0>
0C
#901350000000
1!
1*
b101 6
19
1>
1C
b101 G
#901360000000
0!
0*
09
0>
0C
#901370000000
1!
1*
b110 6
19
1>
1C
b110 G
#901380000000
0!
0*
09
0>
0C
#901390000000
1!
1*
b111 6
19
1>
1C
b111 G
#901400000000
0!
0*
09
0>
0C
#901410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#901420000000
0!
0*
09
0>
0C
#901430000000
1!
1*
b1 6
19
1>
1C
b1 G
#901440000000
0!
0*
09
0>
0C
#901450000000
1!
1*
b10 6
19
1>
1C
b10 G
#901460000000
0!
0*
09
0>
0C
#901470000000
1!
1*
b11 6
19
1>
1C
b11 G
#901480000000
0!
0*
09
0>
0C
#901490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#901500000000
0!
0*
09
0>
0C
#901510000000
1!
1*
b101 6
19
1>
1C
b101 G
#901520000000
0!
0*
09
0>
0C
#901530000000
1!
1*
b110 6
19
1>
1C
b110 G
#901540000000
0!
0*
09
0>
0C
#901550000000
1!
1*
b111 6
19
1>
1C
b111 G
#901560000000
0!
0*
09
0>
0C
#901570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#901580000000
0!
0*
09
0>
0C
#901590000000
1!
1*
b1 6
19
1>
1C
b1 G
#901600000000
0!
0*
09
0>
0C
#901610000000
1!
1*
b10 6
19
1>
1C
b10 G
#901620000000
0!
0*
09
0>
0C
#901630000000
1!
1*
b11 6
19
1>
1C
b11 G
#901640000000
0!
0*
09
0>
0C
#901650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#901660000000
0!
0*
09
0>
0C
#901670000000
1!
1*
b101 6
19
1>
1C
b101 G
#901680000000
0!
0*
09
0>
0C
#901690000000
1!
1*
b110 6
19
1>
1C
b110 G
#901700000000
0!
0*
09
0>
0C
#901710000000
1!
1*
b111 6
19
1>
1C
b111 G
#901720000000
0!
1"
0*
1+
09
1:
0>
0C
#901730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#901740000000
0!
0*
09
0>
0C
#901750000000
1!
1*
b1 6
19
1>
1C
b1 G
#901760000000
0!
0*
09
0>
0C
#901770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#901780000000
0!
0*
09
0>
0C
#901790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#901800000000
0!
0*
09
0>
0C
#901810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#901820000000
0!
0*
09
0>
0C
#901830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#901840000000
0!
0#
0*
0,
09
0>
0?
0C
#901850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#901860000000
0!
0*
09
0>
0C
#901870000000
1!
1*
19
1>
1C
#901880000000
0!
0*
09
0>
0C
#901890000000
1!
1*
19
1>
1C
#901900000000
0!
0*
09
0>
0C
#901910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#901920000000
0!
0*
09
0>
0C
#901930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#901940000000
0!
0*
09
0>
0C
#901950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#901960000000
0!
0*
09
0>
0C
#901970000000
1!
1*
b10 6
19
1>
1C
b10 G
#901980000000
0!
0*
09
0>
0C
#901990000000
1!
1*
b11 6
19
1>
1C
b11 G
#902000000000
0!
0*
09
0>
0C
#902010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#902020000000
0!
0*
09
0>
0C
#902030000000
1!
1*
b101 6
19
1>
1C
b101 G
#902040000000
0!
0*
09
0>
0C
#902050000000
1!
1*
b110 6
19
1>
1C
b110 G
#902060000000
0!
0*
09
0>
0C
#902070000000
1!
1*
b111 6
19
1>
1C
b111 G
#902080000000
0!
0*
09
0>
0C
#902090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#902100000000
0!
0*
09
0>
0C
#902110000000
1!
1*
b1 6
19
1>
1C
b1 G
#902120000000
0!
0*
09
0>
0C
#902130000000
1!
1*
b10 6
19
1>
1C
b10 G
#902140000000
0!
0*
09
0>
0C
#902150000000
1!
1*
b11 6
19
1>
1C
b11 G
#902160000000
0!
0*
09
0>
0C
#902170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#902180000000
0!
0*
09
0>
0C
#902190000000
1!
1*
b101 6
19
1>
1C
b101 G
#902200000000
0!
0*
09
0>
0C
#902210000000
1!
1*
b110 6
19
1>
1C
b110 G
#902220000000
0!
0*
09
0>
0C
#902230000000
1!
1*
b111 6
19
1>
1C
b111 G
#902240000000
0!
0*
09
0>
0C
#902250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#902260000000
0!
0*
09
0>
0C
#902270000000
1!
1*
b1 6
19
1>
1C
b1 G
#902280000000
0!
0*
09
0>
0C
#902290000000
1!
1*
b10 6
19
1>
1C
b10 G
#902300000000
0!
0*
09
0>
0C
#902310000000
1!
1*
b11 6
19
1>
1C
b11 G
#902320000000
0!
0*
09
0>
0C
#902330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#902340000000
0!
0*
09
0>
0C
#902350000000
1!
1*
b101 6
19
1>
1C
b101 G
#902360000000
0!
0*
09
0>
0C
#902370000000
1!
1*
b110 6
19
1>
1C
b110 G
#902380000000
0!
0*
09
0>
0C
#902390000000
1!
1*
b111 6
19
1>
1C
b111 G
#902400000000
0!
1"
0*
1+
09
1:
0>
0C
#902410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#902420000000
0!
0*
09
0>
0C
#902430000000
1!
1*
b1 6
19
1>
1C
b1 G
#902440000000
0!
0*
09
0>
0C
#902450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#902460000000
0!
0*
09
0>
0C
#902470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#902480000000
0!
0*
09
0>
0C
#902490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#902500000000
0!
0*
09
0>
0C
#902510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#902520000000
0!
0#
0*
0,
09
0>
0?
0C
#902530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#902540000000
0!
0*
09
0>
0C
#902550000000
1!
1*
19
1>
1C
#902560000000
0!
0*
09
0>
0C
#902570000000
1!
1*
19
1>
1C
#902580000000
0!
0*
09
0>
0C
#902590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#902600000000
0!
0*
09
0>
0C
#902610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#902620000000
0!
0*
09
0>
0C
#902630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#902640000000
0!
0*
09
0>
0C
#902650000000
1!
1*
b10 6
19
1>
1C
b10 G
#902660000000
0!
0*
09
0>
0C
#902670000000
1!
1*
b11 6
19
1>
1C
b11 G
#902680000000
0!
0*
09
0>
0C
#902690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#902700000000
0!
0*
09
0>
0C
#902710000000
1!
1*
b101 6
19
1>
1C
b101 G
#902720000000
0!
0*
09
0>
0C
#902730000000
1!
1*
b110 6
19
1>
1C
b110 G
#902740000000
0!
0*
09
0>
0C
#902750000000
1!
1*
b111 6
19
1>
1C
b111 G
#902760000000
0!
0*
09
0>
0C
#902770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#902780000000
0!
0*
09
0>
0C
#902790000000
1!
1*
b1 6
19
1>
1C
b1 G
#902800000000
0!
0*
09
0>
0C
#902810000000
1!
1*
b10 6
19
1>
1C
b10 G
#902820000000
0!
0*
09
0>
0C
#902830000000
1!
1*
b11 6
19
1>
1C
b11 G
#902840000000
0!
0*
09
0>
0C
#902850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#902860000000
0!
0*
09
0>
0C
#902870000000
1!
1*
b101 6
19
1>
1C
b101 G
#902880000000
0!
0*
09
0>
0C
#902890000000
1!
1*
b110 6
19
1>
1C
b110 G
#902900000000
0!
0*
09
0>
0C
#902910000000
1!
1*
b111 6
19
1>
1C
b111 G
#902920000000
0!
0*
09
0>
0C
#902930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#902940000000
0!
0*
09
0>
0C
#902950000000
1!
1*
b1 6
19
1>
1C
b1 G
#902960000000
0!
0*
09
0>
0C
#902970000000
1!
1*
b10 6
19
1>
1C
b10 G
#902980000000
0!
0*
09
0>
0C
#902990000000
1!
1*
b11 6
19
1>
1C
b11 G
#903000000000
0!
0*
09
0>
0C
#903010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#903020000000
0!
0*
09
0>
0C
#903030000000
1!
1*
b101 6
19
1>
1C
b101 G
#903040000000
0!
0*
09
0>
0C
#903050000000
1!
1*
b110 6
19
1>
1C
b110 G
#903060000000
0!
0*
09
0>
0C
#903070000000
1!
1*
b111 6
19
1>
1C
b111 G
#903080000000
0!
1"
0*
1+
09
1:
0>
0C
#903090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#903100000000
0!
0*
09
0>
0C
#903110000000
1!
1*
b1 6
19
1>
1C
b1 G
#903120000000
0!
0*
09
0>
0C
#903130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#903140000000
0!
0*
09
0>
0C
#903150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#903160000000
0!
0*
09
0>
0C
#903170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#903180000000
0!
0*
09
0>
0C
#903190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#903200000000
0!
0#
0*
0,
09
0>
0?
0C
#903210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#903220000000
0!
0*
09
0>
0C
#903230000000
1!
1*
19
1>
1C
#903240000000
0!
0*
09
0>
0C
#903250000000
1!
1*
19
1>
1C
#903260000000
0!
0*
09
0>
0C
#903270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#903280000000
0!
0*
09
0>
0C
#903290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#903300000000
0!
0*
09
0>
0C
#903310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#903320000000
0!
0*
09
0>
0C
#903330000000
1!
1*
b10 6
19
1>
1C
b10 G
#903340000000
0!
0*
09
0>
0C
#903350000000
1!
1*
b11 6
19
1>
1C
b11 G
#903360000000
0!
0*
09
0>
0C
#903370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#903380000000
0!
0*
09
0>
0C
#903390000000
1!
1*
b101 6
19
1>
1C
b101 G
#903400000000
0!
0*
09
0>
0C
#903410000000
1!
1*
b110 6
19
1>
1C
b110 G
#903420000000
0!
0*
09
0>
0C
#903430000000
1!
1*
b111 6
19
1>
1C
b111 G
#903440000000
0!
0*
09
0>
0C
#903450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#903460000000
0!
0*
09
0>
0C
#903470000000
1!
1*
b1 6
19
1>
1C
b1 G
#903480000000
0!
0*
09
0>
0C
#903490000000
1!
1*
b10 6
19
1>
1C
b10 G
#903500000000
0!
0*
09
0>
0C
#903510000000
1!
1*
b11 6
19
1>
1C
b11 G
#903520000000
0!
0*
09
0>
0C
#903530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#903540000000
0!
0*
09
0>
0C
#903550000000
1!
1*
b101 6
19
1>
1C
b101 G
#903560000000
0!
0*
09
0>
0C
#903570000000
1!
1*
b110 6
19
1>
1C
b110 G
#903580000000
0!
0*
09
0>
0C
#903590000000
1!
1*
b111 6
19
1>
1C
b111 G
#903600000000
0!
0*
09
0>
0C
#903610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#903620000000
0!
0*
09
0>
0C
#903630000000
1!
1*
b1 6
19
1>
1C
b1 G
#903640000000
0!
0*
09
0>
0C
#903650000000
1!
1*
b10 6
19
1>
1C
b10 G
#903660000000
0!
0*
09
0>
0C
#903670000000
1!
1*
b11 6
19
1>
1C
b11 G
#903680000000
0!
0*
09
0>
0C
#903690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#903700000000
0!
0*
09
0>
0C
#903710000000
1!
1*
b101 6
19
1>
1C
b101 G
#903720000000
0!
0*
09
0>
0C
#903730000000
1!
1*
b110 6
19
1>
1C
b110 G
#903740000000
0!
0*
09
0>
0C
#903750000000
1!
1*
b111 6
19
1>
1C
b111 G
#903760000000
0!
1"
0*
1+
09
1:
0>
0C
#903770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#903780000000
0!
0*
09
0>
0C
#903790000000
1!
1*
b1 6
19
1>
1C
b1 G
#903800000000
0!
0*
09
0>
0C
#903810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#903820000000
0!
0*
09
0>
0C
#903830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#903840000000
0!
0*
09
0>
0C
#903850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#903860000000
0!
0*
09
0>
0C
#903870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#903880000000
0!
0#
0*
0,
09
0>
0?
0C
#903890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#903900000000
0!
0*
09
0>
0C
#903910000000
1!
1*
19
1>
1C
#903920000000
0!
0*
09
0>
0C
#903930000000
1!
1*
19
1>
1C
#903940000000
0!
0*
09
0>
0C
#903950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#903960000000
0!
0*
09
0>
0C
#903970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#903980000000
0!
0*
09
0>
0C
#903990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#904000000000
0!
0*
09
0>
0C
#904010000000
1!
1*
b10 6
19
1>
1C
b10 G
#904020000000
0!
0*
09
0>
0C
#904030000000
1!
1*
b11 6
19
1>
1C
b11 G
#904040000000
0!
0*
09
0>
0C
#904050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#904060000000
0!
0*
09
0>
0C
#904070000000
1!
1*
b101 6
19
1>
1C
b101 G
#904080000000
0!
0*
09
0>
0C
#904090000000
1!
1*
b110 6
19
1>
1C
b110 G
#904100000000
0!
0*
09
0>
0C
#904110000000
1!
1*
b111 6
19
1>
1C
b111 G
#904120000000
0!
0*
09
0>
0C
#904130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#904140000000
0!
0*
09
0>
0C
#904150000000
1!
1*
b1 6
19
1>
1C
b1 G
#904160000000
0!
0*
09
0>
0C
#904170000000
1!
1*
b10 6
19
1>
1C
b10 G
#904180000000
0!
0*
09
0>
0C
#904190000000
1!
1*
b11 6
19
1>
1C
b11 G
#904200000000
0!
0*
09
0>
0C
#904210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#904220000000
0!
0*
09
0>
0C
#904230000000
1!
1*
b101 6
19
1>
1C
b101 G
#904240000000
0!
0*
09
0>
0C
#904250000000
1!
1*
b110 6
19
1>
1C
b110 G
#904260000000
0!
0*
09
0>
0C
#904270000000
1!
1*
b111 6
19
1>
1C
b111 G
#904280000000
0!
0*
09
0>
0C
#904290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#904300000000
0!
0*
09
0>
0C
#904310000000
1!
1*
b1 6
19
1>
1C
b1 G
#904320000000
0!
0*
09
0>
0C
#904330000000
1!
1*
b10 6
19
1>
1C
b10 G
#904340000000
0!
0*
09
0>
0C
#904350000000
1!
1*
b11 6
19
1>
1C
b11 G
#904360000000
0!
0*
09
0>
0C
#904370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#904380000000
0!
0*
09
0>
0C
#904390000000
1!
1*
b101 6
19
1>
1C
b101 G
#904400000000
0!
0*
09
0>
0C
#904410000000
1!
1*
b110 6
19
1>
1C
b110 G
#904420000000
0!
0*
09
0>
0C
#904430000000
1!
1*
b111 6
19
1>
1C
b111 G
#904440000000
0!
1"
0*
1+
09
1:
0>
0C
#904450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#904460000000
0!
0*
09
0>
0C
#904470000000
1!
1*
b1 6
19
1>
1C
b1 G
#904480000000
0!
0*
09
0>
0C
#904490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#904500000000
0!
0*
09
0>
0C
#904510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#904520000000
0!
0*
09
0>
0C
#904530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#904540000000
0!
0*
09
0>
0C
#904550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#904560000000
0!
0#
0*
0,
09
0>
0?
0C
#904570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#904580000000
0!
0*
09
0>
0C
#904590000000
1!
1*
19
1>
1C
#904600000000
0!
0*
09
0>
0C
#904610000000
1!
1*
19
1>
1C
#904620000000
0!
0*
09
0>
0C
#904630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#904640000000
0!
0*
09
0>
0C
#904650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#904660000000
0!
0*
09
0>
0C
#904670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#904680000000
0!
0*
09
0>
0C
#904690000000
1!
1*
b10 6
19
1>
1C
b10 G
#904700000000
0!
0*
09
0>
0C
#904710000000
1!
1*
b11 6
19
1>
1C
b11 G
#904720000000
0!
0*
09
0>
0C
#904730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#904740000000
0!
0*
09
0>
0C
#904750000000
1!
1*
b101 6
19
1>
1C
b101 G
#904760000000
0!
0*
09
0>
0C
#904770000000
1!
1*
b110 6
19
1>
1C
b110 G
#904780000000
0!
0*
09
0>
0C
#904790000000
1!
1*
b111 6
19
1>
1C
b111 G
#904800000000
0!
0*
09
0>
0C
#904810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#904820000000
0!
0*
09
0>
0C
#904830000000
1!
1*
b1 6
19
1>
1C
b1 G
#904840000000
0!
0*
09
0>
0C
#904850000000
1!
1*
b10 6
19
1>
1C
b10 G
#904860000000
0!
0*
09
0>
0C
#904870000000
1!
1*
b11 6
19
1>
1C
b11 G
#904880000000
0!
0*
09
0>
0C
#904890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#904900000000
0!
0*
09
0>
0C
#904910000000
1!
1*
b101 6
19
1>
1C
b101 G
#904920000000
0!
0*
09
0>
0C
#904930000000
1!
1*
b110 6
19
1>
1C
b110 G
#904940000000
0!
0*
09
0>
0C
#904950000000
1!
1*
b111 6
19
1>
1C
b111 G
#904960000000
0!
0*
09
0>
0C
#904970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#904980000000
0!
0*
09
0>
0C
#904990000000
1!
1*
b1 6
19
1>
1C
b1 G
#905000000000
0!
0*
09
0>
0C
#905010000000
1!
1*
b10 6
19
1>
1C
b10 G
#905020000000
0!
0*
09
0>
0C
#905030000000
1!
1*
b11 6
19
1>
1C
b11 G
#905040000000
0!
0*
09
0>
0C
#905050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#905060000000
0!
0*
09
0>
0C
#905070000000
1!
1*
b101 6
19
1>
1C
b101 G
#905080000000
0!
0*
09
0>
0C
#905090000000
1!
1*
b110 6
19
1>
1C
b110 G
#905100000000
0!
0*
09
0>
0C
#905110000000
1!
1*
b111 6
19
1>
1C
b111 G
#905120000000
0!
1"
0*
1+
09
1:
0>
0C
#905130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#905140000000
0!
0*
09
0>
0C
#905150000000
1!
1*
b1 6
19
1>
1C
b1 G
#905160000000
0!
0*
09
0>
0C
#905170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#905180000000
0!
0*
09
0>
0C
#905190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#905200000000
0!
0*
09
0>
0C
#905210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#905220000000
0!
0*
09
0>
0C
#905230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#905240000000
0!
0#
0*
0,
09
0>
0?
0C
#905250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#905260000000
0!
0*
09
0>
0C
#905270000000
1!
1*
19
1>
1C
#905280000000
0!
0*
09
0>
0C
#905290000000
1!
1*
19
1>
1C
#905300000000
0!
0*
09
0>
0C
#905310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#905320000000
0!
0*
09
0>
0C
#905330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#905340000000
0!
0*
09
0>
0C
#905350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#905360000000
0!
0*
09
0>
0C
#905370000000
1!
1*
b10 6
19
1>
1C
b10 G
#905380000000
0!
0*
09
0>
0C
#905390000000
1!
1*
b11 6
19
1>
1C
b11 G
#905400000000
0!
0*
09
0>
0C
#905410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#905420000000
0!
0*
09
0>
0C
#905430000000
1!
1*
b101 6
19
1>
1C
b101 G
#905440000000
0!
0*
09
0>
0C
#905450000000
1!
1*
b110 6
19
1>
1C
b110 G
#905460000000
0!
0*
09
0>
0C
#905470000000
1!
1*
b111 6
19
1>
1C
b111 G
#905480000000
0!
0*
09
0>
0C
#905490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#905500000000
0!
0*
09
0>
0C
#905510000000
1!
1*
b1 6
19
1>
1C
b1 G
#905520000000
0!
0*
09
0>
0C
#905530000000
1!
1*
b10 6
19
1>
1C
b10 G
#905540000000
0!
0*
09
0>
0C
#905550000000
1!
1*
b11 6
19
1>
1C
b11 G
#905560000000
0!
0*
09
0>
0C
#905570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#905580000000
0!
0*
09
0>
0C
#905590000000
1!
1*
b101 6
19
1>
1C
b101 G
#905600000000
0!
0*
09
0>
0C
#905610000000
1!
1*
b110 6
19
1>
1C
b110 G
#905620000000
0!
0*
09
0>
0C
#905630000000
1!
1*
b111 6
19
1>
1C
b111 G
#905640000000
0!
0*
09
0>
0C
#905650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#905660000000
0!
0*
09
0>
0C
#905670000000
1!
1*
b1 6
19
1>
1C
b1 G
#905680000000
0!
0*
09
0>
0C
#905690000000
1!
1*
b10 6
19
1>
1C
b10 G
#905700000000
0!
0*
09
0>
0C
#905710000000
1!
1*
b11 6
19
1>
1C
b11 G
#905720000000
0!
0*
09
0>
0C
#905730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#905740000000
0!
0*
09
0>
0C
#905750000000
1!
1*
b101 6
19
1>
1C
b101 G
#905760000000
0!
0*
09
0>
0C
#905770000000
1!
1*
b110 6
19
1>
1C
b110 G
#905780000000
0!
0*
09
0>
0C
#905790000000
1!
1*
b111 6
19
1>
1C
b111 G
#905800000000
0!
1"
0*
1+
09
1:
0>
0C
#905810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#905820000000
0!
0*
09
0>
0C
#905830000000
1!
1*
b1 6
19
1>
1C
b1 G
#905840000000
0!
0*
09
0>
0C
#905850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#905860000000
0!
0*
09
0>
0C
#905870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#905880000000
0!
0*
09
0>
0C
#905890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#905900000000
0!
0*
09
0>
0C
#905910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#905920000000
0!
0#
0*
0,
09
0>
0?
0C
#905930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#905940000000
0!
0*
09
0>
0C
#905950000000
1!
1*
19
1>
1C
#905960000000
0!
0*
09
0>
0C
#905970000000
1!
1*
19
1>
1C
#905980000000
0!
0*
09
0>
0C
#905990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#906000000000
0!
0*
09
0>
0C
#906010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#906020000000
0!
0*
09
0>
0C
#906030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#906040000000
0!
0*
09
0>
0C
#906050000000
1!
1*
b10 6
19
1>
1C
b10 G
#906060000000
0!
0*
09
0>
0C
#906070000000
1!
1*
b11 6
19
1>
1C
b11 G
#906080000000
0!
0*
09
0>
0C
#906090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#906100000000
0!
0*
09
0>
0C
#906110000000
1!
1*
b101 6
19
1>
1C
b101 G
#906120000000
0!
0*
09
0>
0C
#906130000000
1!
1*
b110 6
19
1>
1C
b110 G
#906140000000
0!
0*
09
0>
0C
#906150000000
1!
1*
b111 6
19
1>
1C
b111 G
#906160000000
0!
0*
09
0>
0C
#906170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#906180000000
0!
0*
09
0>
0C
#906190000000
1!
1*
b1 6
19
1>
1C
b1 G
#906200000000
0!
0*
09
0>
0C
#906210000000
1!
1*
b10 6
19
1>
1C
b10 G
#906220000000
0!
0*
09
0>
0C
#906230000000
1!
1*
b11 6
19
1>
1C
b11 G
#906240000000
0!
0*
09
0>
0C
#906250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#906260000000
0!
0*
09
0>
0C
#906270000000
1!
1*
b101 6
19
1>
1C
b101 G
#906280000000
0!
0*
09
0>
0C
#906290000000
1!
1*
b110 6
19
1>
1C
b110 G
#906300000000
0!
0*
09
0>
0C
#906310000000
1!
1*
b111 6
19
1>
1C
b111 G
#906320000000
0!
0*
09
0>
0C
#906330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#906340000000
0!
0*
09
0>
0C
#906350000000
1!
1*
b1 6
19
1>
1C
b1 G
#906360000000
0!
0*
09
0>
0C
#906370000000
1!
1*
b10 6
19
1>
1C
b10 G
#906380000000
0!
0*
09
0>
0C
#906390000000
1!
1*
b11 6
19
1>
1C
b11 G
#906400000000
0!
0*
09
0>
0C
#906410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#906420000000
0!
0*
09
0>
0C
#906430000000
1!
1*
b101 6
19
1>
1C
b101 G
#906440000000
0!
0*
09
0>
0C
#906450000000
1!
1*
b110 6
19
1>
1C
b110 G
#906460000000
0!
0*
09
0>
0C
#906470000000
1!
1*
b111 6
19
1>
1C
b111 G
#906480000000
0!
1"
0*
1+
09
1:
0>
0C
#906490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#906500000000
0!
0*
09
0>
0C
#906510000000
1!
1*
b1 6
19
1>
1C
b1 G
#906520000000
0!
0*
09
0>
0C
#906530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#906540000000
0!
0*
09
0>
0C
#906550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#906560000000
0!
0*
09
0>
0C
#906570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#906580000000
0!
0*
09
0>
0C
#906590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#906600000000
0!
0#
0*
0,
09
0>
0?
0C
#906610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#906620000000
0!
0*
09
0>
0C
#906630000000
1!
1*
19
1>
1C
#906640000000
0!
0*
09
0>
0C
#906650000000
1!
1*
19
1>
1C
#906660000000
0!
0*
09
0>
0C
#906670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#906680000000
0!
0*
09
0>
0C
#906690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#906700000000
0!
0*
09
0>
0C
#906710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#906720000000
0!
0*
09
0>
0C
#906730000000
1!
1*
b10 6
19
1>
1C
b10 G
#906740000000
0!
0*
09
0>
0C
#906750000000
1!
1*
b11 6
19
1>
1C
b11 G
#906760000000
0!
0*
09
0>
0C
#906770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#906780000000
0!
0*
09
0>
0C
#906790000000
1!
1*
b101 6
19
1>
1C
b101 G
#906800000000
0!
0*
09
0>
0C
#906810000000
1!
1*
b110 6
19
1>
1C
b110 G
#906820000000
0!
0*
09
0>
0C
#906830000000
1!
1*
b111 6
19
1>
1C
b111 G
#906840000000
0!
0*
09
0>
0C
#906850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#906860000000
0!
0*
09
0>
0C
#906870000000
1!
1*
b1 6
19
1>
1C
b1 G
#906880000000
0!
0*
09
0>
0C
#906890000000
1!
1*
b10 6
19
1>
1C
b10 G
#906900000000
0!
0*
09
0>
0C
#906910000000
1!
1*
b11 6
19
1>
1C
b11 G
#906920000000
0!
0*
09
0>
0C
#906930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#906940000000
0!
0*
09
0>
0C
#906950000000
1!
1*
b101 6
19
1>
1C
b101 G
#906960000000
0!
0*
09
0>
0C
#906970000000
1!
1*
b110 6
19
1>
1C
b110 G
#906980000000
0!
0*
09
0>
0C
#906990000000
1!
1*
b111 6
19
1>
1C
b111 G
#907000000000
0!
0*
09
0>
0C
#907010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#907020000000
0!
0*
09
0>
0C
#907030000000
1!
1*
b1 6
19
1>
1C
b1 G
#907040000000
0!
0*
09
0>
0C
#907050000000
1!
1*
b10 6
19
1>
1C
b10 G
#907060000000
0!
0*
09
0>
0C
#907070000000
1!
1*
b11 6
19
1>
1C
b11 G
#907080000000
0!
0*
09
0>
0C
#907090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#907100000000
0!
0*
09
0>
0C
#907110000000
1!
1*
b101 6
19
1>
1C
b101 G
#907120000000
0!
0*
09
0>
0C
#907130000000
1!
1*
b110 6
19
1>
1C
b110 G
#907140000000
0!
0*
09
0>
0C
#907150000000
1!
1*
b111 6
19
1>
1C
b111 G
#907160000000
0!
1"
0*
1+
09
1:
0>
0C
#907170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#907180000000
0!
0*
09
0>
0C
#907190000000
1!
1*
b1 6
19
1>
1C
b1 G
#907200000000
0!
0*
09
0>
0C
#907210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#907220000000
0!
0*
09
0>
0C
#907230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#907240000000
0!
0*
09
0>
0C
#907250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#907260000000
0!
0*
09
0>
0C
#907270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#907280000000
0!
0#
0*
0,
09
0>
0?
0C
#907290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#907300000000
0!
0*
09
0>
0C
#907310000000
1!
1*
19
1>
1C
#907320000000
0!
0*
09
0>
0C
#907330000000
1!
1*
19
1>
1C
#907340000000
0!
0*
09
0>
0C
#907350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#907360000000
0!
0*
09
0>
0C
#907370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#907380000000
0!
0*
09
0>
0C
#907390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#907400000000
0!
0*
09
0>
0C
#907410000000
1!
1*
b10 6
19
1>
1C
b10 G
#907420000000
0!
0*
09
0>
0C
#907430000000
1!
1*
b11 6
19
1>
1C
b11 G
#907440000000
0!
0*
09
0>
0C
#907450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#907460000000
0!
0*
09
0>
0C
#907470000000
1!
1*
b101 6
19
1>
1C
b101 G
#907480000000
0!
0*
09
0>
0C
#907490000000
1!
1*
b110 6
19
1>
1C
b110 G
#907500000000
0!
0*
09
0>
0C
#907510000000
1!
1*
b111 6
19
1>
1C
b111 G
#907520000000
0!
0*
09
0>
0C
#907530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#907540000000
0!
0*
09
0>
0C
#907550000000
1!
1*
b1 6
19
1>
1C
b1 G
#907560000000
0!
0*
09
0>
0C
#907570000000
1!
1*
b10 6
19
1>
1C
b10 G
#907580000000
0!
0*
09
0>
0C
#907590000000
1!
1*
b11 6
19
1>
1C
b11 G
#907600000000
0!
0*
09
0>
0C
#907610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#907620000000
0!
0*
09
0>
0C
#907630000000
1!
1*
b101 6
19
1>
1C
b101 G
#907640000000
0!
0*
09
0>
0C
#907650000000
1!
1*
b110 6
19
1>
1C
b110 G
#907660000000
0!
0*
09
0>
0C
#907670000000
1!
1*
b111 6
19
1>
1C
b111 G
#907680000000
0!
0*
09
0>
0C
#907690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#907700000000
0!
0*
09
0>
0C
#907710000000
1!
1*
b1 6
19
1>
1C
b1 G
#907720000000
0!
0*
09
0>
0C
#907730000000
1!
1*
b10 6
19
1>
1C
b10 G
#907740000000
0!
0*
09
0>
0C
#907750000000
1!
1*
b11 6
19
1>
1C
b11 G
#907760000000
0!
0*
09
0>
0C
#907770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#907780000000
0!
0*
09
0>
0C
#907790000000
1!
1*
b101 6
19
1>
1C
b101 G
#907800000000
0!
0*
09
0>
0C
#907810000000
1!
1*
b110 6
19
1>
1C
b110 G
#907820000000
0!
0*
09
0>
0C
#907830000000
1!
1*
b111 6
19
1>
1C
b111 G
#907840000000
0!
1"
0*
1+
09
1:
0>
0C
#907850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#907860000000
0!
0*
09
0>
0C
#907870000000
1!
1*
b1 6
19
1>
1C
b1 G
#907880000000
0!
0*
09
0>
0C
#907890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#907900000000
0!
0*
09
0>
0C
#907910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#907920000000
0!
0*
09
0>
0C
#907930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#907940000000
0!
0*
09
0>
0C
#907950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#907960000000
0!
0#
0*
0,
09
0>
0?
0C
#907970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#907980000000
0!
0*
09
0>
0C
#907990000000
1!
1*
19
1>
1C
#908000000000
0!
0*
09
0>
0C
#908010000000
1!
1*
19
1>
1C
#908020000000
0!
0*
09
0>
0C
#908030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#908040000000
0!
0*
09
0>
0C
#908050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#908060000000
0!
0*
09
0>
0C
#908070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#908080000000
0!
0*
09
0>
0C
#908090000000
1!
1*
b10 6
19
1>
1C
b10 G
#908100000000
0!
0*
09
0>
0C
#908110000000
1!
1*
b11 6
19
1>
1C
b11 G
#908120000000
0!
0*
09
0>
0C
#908130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#908140000000
0!
0*
09
0>
0C
#908150000000
1!
1*
b101 6
19
1>
1C
b101 G
#908160000000
0!
0*
09
0>
0C
#908170000000
1!
1*
b110 6
19
1>
1C
b110 G
#908180000000
0!
0*
09
0>
0C
#908190000000
1!
1*
b111 6
19
1>
1C
b111 G
#908200000000
0!
0*
09
0>
0C
#908210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#908220000000
0!
0*
09
0>
0C
#908230000000
1!
1*
b1 6
19
1>
1C
b1 G
#908240000000
0!
0*
09
0>
0C
#908250000000
1!
1*
b10 6
19
1>
1C
b10 G
#908260000000
0!
0*
09
0>
0C
#908270000000
1!
1*
b11 6
19
1>
1C
b11 G
#908280000000
0!
0*
09
0>
0C
#908290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#908300000000
0!
0*
09
0>
0C
#908310000000
1!
1*
b101 6
19
1>
1C
b101 G
#908320000000
0!
0*
09
0>
0C
#908330000000
1!
1*
b110 6
19
1>
1C
b110 G
#908340000000
0!
0*
09
0>
0C
#908350000000
1!
1*
b111 6
19
1>
1C
b111 G
#908360000000
0!
0*
09
0>
0C
#908370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#908380000000
0!
0*
09
0>
0C
#908390000000
1!
1*
b1 6
19
1>
1C
b1 G
#908400000000
0!
0*
09
0>
0C
#908410000000
1!
1*
b10 6
19
1>
1C
b10 G
#908420000000
0!
0*
09
0>
0C
#908430000000
1!
1*
b11 6
19
1>
1C
b11 G
#908440000000
0!
0*
09
0>
0C
#908450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#908460000000
0!
0*
09
0>
0C
#908470000000
1!
1*
b101 6
19
1>
1C
b101 G
#908480000000
0!
0*
09
0>
0C
#908490000000
1!
1*
b110 6
19
1>
1C
b110 G
#908500000000
0!
0*
09
0>
0C
#908510000000
1!
1*
b111 6
19
1>
1C
b111 G
#908520000000
0!
1"
0*
1+
09
1:
0>
0C
#908530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#908540000000
0!
0*
09
0>
0C
#908550000000
1!
1*
b1 6
19
1>
1C
b1 G
#908560000000
0!
0*
09
0>
0C
#908570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#908580000000
0!
0*
09
0>
0C
#908590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#908600000000
0!
0*
09
0>
0C
#908610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#908620000000
0!
0*
09
0>
0C
#908630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#908640000000
0!
0#
0*
0,
09
0>
0?
0C
#908650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#908660000000
0!
0*
09
0>
0C
#908670000000
1!
1*
19
1>
1C
#908680000000
0!
0*
09
0>
0C
#908690000000
1!
1*
19
1>
1C
#908700000000
0!
0*
09
0>
0C
#908710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#908720000000
0!
0*
09
0>
0C
#908730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#908740000000
0!
0*
09
0>
0C
#908750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#908760000000
0!
0*
09
0>
0C
#908770000000
1!
1*
b10 6
19
1>
1C
b10 G
#908780000000
0!
0*
09
0>
0C
#908790000000
1!
1*
b11 6
19
1>
1C
b11 G
#908800000000
0!
0*
09
0>
0C
#908810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#908820000000
0!
0*
09
0>
0C
#908830000000
1!
1*
b101 6
19
1>
1C
b101 G
#908840000000
0!
0*
09
0>
0C
#908850000000
1!
1*
b110 6
19
1>
1C
b110 G
#908860000000
0!
0*
09
0>
0C
#908870000000
1!
1*
b111 6
19
1>
1C
b111 G
#908880000000
0!
0*
09
0>
0C
#908890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#908900000000
0!
0*
09
0>
0C
#908910000000
1!
1*
b1 6
19
1>
1C
b1 G
#908920000000
0!
0*
09
0>
0C
#908930000000
1!
1*
b10 6
19
1>
1C
b10 G
#908940000000
0!
0*
09
0>
0C
#908950000000
1!
1*
b11 6
19
1>
1C
b11 G
#908960000000
0!
0*
09
0>
0C
#908970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#908980000000
0!
0*
09
0>
0C
#908990000000
1!
1*
b101 6
19
1>
1C
b101 G
#909000000000
0!
0*
09
0>
0C
#909010000000
1!
1*
b110 6
19
1>
1C
b110 G
#909020000000
0!
0*
09
0>
0C
#909030000000
1!
1*
b111 6
19
1>
1C
b111 G
#909040000000
0!
0*
09
0>
0C
#909050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#909060000000
0!
0*
09
0>
0C
#909070000000
1!
1*
b1 6
19
1>
1C
b1 G
#909080000000
0!
0*
09
0>
0C
#909090000000
1!
1*
b10 6
19
1>
1C
b10 G
#909100000000
0!
0*
09
0>
0C
#909110000000
1!
1*
b11 6
19
1>
1C
b11 G
#909120000000
0!
0*
09
0>
0C
#909130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#909140000000
0!
0*
09
0>
0C
#909150000000
1!
1*
b101 6
19
1>
1C
b101 G
#909160000000
0!
0*
09
0>
0C
#909170000000
1!
1*
b110 6
19
1>
1C
b110 G
#909180000000
0!
0*
09
0>
0C
#909190000000
1!
1*
b111 6
19
1>
1C
b111 G
#909200000000
0!
1"
0*
1+
09
1:
0>
0C
#909210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#909220000000
0!
0*
09
0>
0C
#909230000000
1!
1*
b1 6
19
1>
1C
b1 G
#909240000000
0!
0*
09
0>
0C
#909250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#909260000000
0!
0*
09
0>
0C
#909270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#909280000000
0!
0*
09
0>
0C
#909290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#909300000000
0!
0*
09
0>
0C
#909310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#909320000000
0!
0#
0*
0,
09
0>
0?
0C
#909330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#909340000000
0!
0*
09
0>
0C
#909350000000
1!
1*
19
1>
1C
#909360000000
0!
0*
09
0>
0C
#909370000000
1!
1*
19
1>
1C
#909380000000
0!
0*
09
0>
0C
#909390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#909400000000
0!
0*
09
0>
0C
#909410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#909420000000
0!
0*
09
0>
0C
#909430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#909440000000
0!
0*
09
0>
0C
#909450000000
1!
1*
b10 6
19
1>
1C
b10 G
#909460000000
0!
0*
09
0>
0C
#909470000000
1!
1*
b11 6
19
1>
1C
b11 G
#909480000000
0!
0*
09
0>
0C
#909490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#909500000000
0!
0*
09
0>
0C
#909510000000
1!
1*
b101 6
19
1>
1C
b101 G
#909520000000
0!
0*
09
0>
0C
#909530000000
1!
1*
b110 6
19
1>
1C
b110 G
#909540000000
0!
0*
09
0>
0C
#909550000000
1!
1*
b111 6
19
1>
1C
b111 G
#909560000000
0!
0*
09
0>
0C
#909570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#909580000000
0!
0*
09
0>
0C
#909590000000
1!
1*
b1 6
19
1>
1C
b1 G
#909600000000
0!
0*
09
0>
0C
#909610000000
1!
1*
b10 6
19
1>
1C
b10 G
#909620000000
0!
0*
09
0>
0C
#909630000000
1!
1*
b11 6
19
1>
1C
b11 G
#909640000000
0!
0*
09
0>
0C
#909650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#909660000000
0!
0*
09
0>
0C
#909670000000
1!
1*
b101 6
19
1>
1C
b101 G
#909680000000
0!
0*
09
0>
0C
#909690000000
1!
1*
b110 6
19
1>
1C
b110 G
#909700000000
0!
0*
09
0>
0C
#909710000000
1!
1*
b111 6
19
1>
1C
b111 G
#909720000000
0!
0*
09
0>
0C
#909730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#909740000000
0!
0*
09
0>
0C
#909750000000
1!
1*
b1 6
19
1>
1C
b1 G
#909760000000
0!
0*
09
0>
0C
#909770000000
1!
1*
b10 6
19
1>
1C
b10 G
#909780000000
0!
0*
09
0>
0C
#909790000000
1!
1*
b11 6
19
1>
1C
b11 G
#909800000000
0!
0*
09
0>
0C
#909810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#909820000000
0!
0*
09
0>
0C
#909830000000
1!
1*
b101 6
19
1>
1C
b101 G
#909840000000
0!
0*
09
0>
0C
#909850000000
1!
1*
b110 6
19
1>
1C
b110 G
#909860000000
0!
0*
09
0>
0C
#909870000000
1!
1*
b111 6
19
1>
1C
b111 G
#909880000000
0!
1"
0*
1+
09
1:
0>
0C
#909890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#909900000000
0!
0*
09
0>
0C
#909910000000
1!
1*
b1 6
19
1>
1C
b1 G
#909920000000
0!
0*
09
0>
0C
#909930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#909940000000
0!
0*
09
0>
0C
#909950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#909960000000
0!
0*
09
0>
0C
#909970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#909980000000
0!
0*
09
0>
0C
#909990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#910000000000
0!
0#
0*
0,
09
0>
0?
0C
#910010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#910020000000
0!
0*
09
0>
0C
#910030000000
1!
1*
19
1>
1C
#910040000000
0!
0*
09
0>
0C
#910050000000
1!
1*
19
1>
1C
#910060000000
0!
0*
09
0>
0C
#910070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#910080000000
0!
0*
09
0>
0C
#910090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#910100000000
0!
0*
09
0>
0C
#910110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#910120000000
0!
0*
09
0>
0C
#910130000000
1!
1*
b10 6
19
1>
1C
b10 G
#910140000000
0!
0*
09
0>
0C
#910150000000
1!
1*
b11 6
19
1>
1C
b11 G
#910160000000
0!
0*
09
0>
0C
#910170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#910180000000
0!
0*
09
0>
0C
#910190000000
1!
1*
b101 6
19
1>
1C
b101 G
#910200000000
0!
0*
09
0>
0C
#910210000000
1!
1*
b110 6
19
1>
1C
b110 G
#910220000000
0!
0*
09
0>
0C
#910230000000
1!
1*
b111 6
19
1>
1C
b111 G
#910240000000
0!
0*
09
0>
0C
#910250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#910260000000
0!
0*
09
0>
0C
#910270000000
1!
1*
b1 6
19
1>
1C
b1 G
#910280000000
0!
0*
09
0>
0C
#910290000000
1!
1*
b10 6
19
1>
1C
b10 G
#910300000000
0!
0*
09
0>
0C
#910310000000
1!
1*
b11 6
19
1>
1C
b11 G
#910320000000
0!
0*
09
0>
0C
#910330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#910340000000
0!
0*
09
0>
0C
#910350000000
1!
1*
b101 6
19
1>
1C
b101 G
#910360000000
0!
0*
09
0>
0C
#910370000000
1!
1*
b110 6
19
1>
1C
b110 G
#910380000000
0!
0*
09
0>
0C
#910390000000
1!
1*
b111 6
19
1>
1C
b111 G
#910400000000
0!
0*
09
0>
0C
#910410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#910420000000
0!
0*
09
0>
0C
#910430000000
1!
1*
b1 6
19
1>
1C
b1 G
#910440000000
0!
0*
09
0>
0C
#910450000000
1!
1*
b10 6
19
1>
1C
b10 G
#910460000000
0!
0*
09
0>
0C
#910470000000
1!
1*
b11 6
19
1>
1C
b11 G
#910480000000
0!
0*
09
0>
0C
#910490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#910500000000
0!
0*
09
0>
0C
#910510000000
1!
1*
b101 6
19
1>
1C
b101 G
#910520000000
0!
0*
09
0>
0C
#910530000000
1!
1*
b110 6
19
1>
1C
b110 G
#910540000000
0!
0*
09
0>
0C
#910550000000
1!
1*
b111 6
19
1>
1C
b111 G
#910560000000
0!
1"
0*
1+
09
1:
0>
0C
#910570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#910580000000
0!
0*
09
0>
0C
#910590000000
1!
1*
b1 6
19
1>
1C
b1 G
#910600000000
0!
0*
09
0>
0C
#910610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#910620000000
0!
0*
09
0>
0C
#910630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#910640000000
0!
0*
09
0>
0C
#910650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#910660000000
0!
0*
09
0>
0C
#910670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#910680000000
0!
0#
0*
0,
09
0>
0?
0C
#910690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#910700000000
0!
0*
09
0>
0C
#910710000000
1!
1*
19
1>
1C
#910720000000
0!
0*
09
0>
0C
#910730000000
1!
1*
19
1>
1C
#910740000000
0!
0*
09
0>
0C
#910750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#910760000000
0!
0*
09
0>
0C
#910770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#910780000000
0!
0*
09
0>
0C
#910790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#910800000000
0!
0*
09
0>
0C
#910810000000
1!
1*
b10 6
19
1>
1C
b10 G
#910820000000
0!
0*
09
0>
0C
#910830000000
1!
1*
b11 6
19
1>
1C
b11 G
#910840000000
0!
0*
09
0>
0C
#910850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#910860000000
0!
0*
09
0>
0C
#910870000000
1!
1*
b101 6
19
1>
1C
b101 G
#910880000000
0!
0*
09
0>
0C
#910890000000
1!
1*
b110 6
19
1>
1C
b110 G
#910900000000
0!
0*
09
0>
0C
#910910000000
1!
1*
b111 6
19
1>
1C
b111 G
#910920000000
0!
0*
09
0>
0C
#910930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#910940000000
0!
0*
09
0>
0C
#910950000000
1!
1*
b1 6
19
1>
1C
b1 G
#910960000000
0!
0*
09
0>
0C
#910970000000
1!
1*
b10 6
19
1>
1C
b10 G
#910980000000
0!
0*
09
0>
0C
#910990000000
1!
1*
b11 6
19
1>
1C
b11 G
#911000000000
0!
0*
09
0>
0C
#911010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#911020000000
0!
0*
09
0>
0C
#911030000000
1!
1*
b101 6
19
1>
1C
b101 G
#911040000000
0!
0*
09
0>
0C
#911050000000
1!
1*
b110 6
19
1>
1C
b110 G
#911060000000
0!
0*
09
0>
0C
#911070000000
1!
1*
b111 6
19
1>
1C
b111 G
#911080000000
0!
0*
09
0>
0C
#911090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#911100000000
0!
0*
09
0>
0C
#911110000000
1!
1*
b1 6
19
1>
1C
b1 G
#911120000000
0!
0*
09
0>
0C
#911130000000
1!
1*
b10 6
19
1>
1C
b10 G
#911140000000
0!
0*
09
0>
0C
#911150000000
1!
1*
b11 6
19
1>
1C
b11 G
#911160000000
0!
0*
09
0>
0C
#911170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#911180000000
0!
0*
09
0>
0C
#911190000000
1!
1*
b101 6
19
1>
1C
b101 G
#911200000000
0!
0*
09
0>
0C
#911210000000
1!
1*
b110 6
19
1>
1C
b110 G
#911220000000
0!
0*
09
0>
0C
#911230000000
1!
1*
b111 6
19
1>
1C
b111 G
#911240000000
0!
1"
0*
1+
09
1:
0>
0C
#911250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#911260000000
0!
0*
09
0>
0C
#911270000000
1!
1*
b1 6
19
1>
1C
b1 G
#911280000000
0!
0*
09
0>
0C
#911290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#911300000000
0!
0*
09
0>
0C
#911310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#911320000000
0!
0*
09
0>
0C
#911330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#911340000000
0!
0*
09
0>
0C
#911350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#911360000000
0!
0#
0*
0,
09
0>
0?
0C
#911370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#911380000000
0!
0*
09
0>
0C
#911390000000
1!
1*
19
1>
1C
#911400000000
0!
0*
09
0>
0C
#911410000000
1!
1*
19
1>
1C
#911420000000
0!
0*
09
0>
0C
#911430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#911440000000
0!
0*
09
0>
0C
#911450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#911460000000
0!
0*
09
0>
0C
#911470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#911480000000
0!
0*
09
0>
0C
#911490000000
1!
1*
b10 6
19
1>
1C
b10 G
#911500000000
0!
0*
09
0>
0C
#911510000000
1!
1*
b11 6
19
1>
1C
b11 G
#911520000000
0!
0*
09
0>
0C
#911530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#911540000000
0!
0*
09
0>
0C
#911550000000
1!
1*
b101 6
19
1>
1C
b101 G
#911560000000
0!
0*
09
0>
0C
#911570000000
1!
1*
b110 6
19
1>
1C
b110 G
#911580000000
0!
0*
09
0>
0C
#911590000000
1!
1*
b111 6
19
1>
1C
b111 G
#911600000000
0!
0*
09
0>
0C
#911610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#911620000000
0!
0*
09
0>
0C
#911630000000
1!
1*
b1 6
19
1>
1C
b1 G
#911640000000
0!
0*
09
0>
0C
#911650000000
1!
1*
b10 6
19
1>
1C
b10 G
#911660000000
0!
0*
09
0>
0C
#911670000000
1!
1*
b11 6
19
1>
1C
b11 G
#911680000000
0!
0*
09
0>
0C
#911690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#911700000000
0!
0*
09
0>
0C
#911710000000
1!
1*
b101 6
19
1>
1C
b101 G
#911720000000
0!
0*
09
0>
0C
#911730000000
1!
1*
b110 6
19
1>
1C
b110 G
#911740000000
0!
0*
09
0>
0C
#911750000000
1!
1*
b111 6
19
1>
1C
b111 G
#911760000000
0!
0*
09
0>
0C
#911770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#911780000000
0!
0*
09
0>
0C
#911790000000
1!
1*
b1 6
19
1>
1C
b1 G
#911800000000
0!
0*
09
0>
0C
#911810000000
1!
1*
b10 6
19
1>
1C
b10 G
#911820000000
0!
0*
09
0>
0C
#911830000000
1!
1*
b11 6
19
1>
1C
b11 G
#911840000000
0!
0*
09
0>
0C
#911850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#911860000000
0!
0*
09
0>
0C
#911870000000
1!
1*
b101 6
19
1>
1C
b101 G
#911880000000
0!
0*
09
0>
0C
#911890000000
1!
1*
b110 6
19
1>
1C
b110 G
#911900000000
0!
0*
09
0>
0C
#911910000000
1!
1*
b111 6
19
1>
1C
b111 G
#911920000000
0!
1"
0*
1+
09
1:
0>
0C
#911930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#911940000000
0!
0*
09
0>
0C
#911950000000
1!
1*
b1 6
19
1>
1C
b1 G
#911960000000
0!
0*
09
0>
0C
#911970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#911980000000
0!
0*
09
0>
0C
#911990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#912000000000
0!
0*
09
0>
0C
#912010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#912020000000
0!
0*
09
0>
0C
#912030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#912040000000
0!
0#
0*
0,
09
0>
0?
0C
#912050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#912060000000
0!
0*
09
0>
0C
#912070000000
1!
1*
19
1>
1C
#912080000000
0!
0*
09
0>
0C
#912090000000
1!
1*
19
1>
1C
#912100000000
0!
0*
09
0>
0C
#912110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#912120000000
0!
0*
09
0>
0C
#912130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#912140000000
0!
0*
09
0>
0C
#912150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#912160000000
0!
0*
09
0>
0C
#912170000000
1!
1*
b10 6
19
1>
1C
b10 G
#912180000000
0!
0*
09
0>
0C
#912190000000
1!
1*
b11 6
19
1>
1C
b11 G
#912200000000
0!
0*
09
0>
0C
#912210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#912220000000
0!
0*
09
0>
0C
#912230000000
1!
1*
b101 6
19
1>
1C
b101 G
#912240000000
0!
0*
09
0>
0C
#912250000000
1!
1*
b110 6
19
1>
1C
b110 G
#912260000000
0!
0*
09
0>
0C
#912270000000
1!
1*
b111 6
19
1>
1C
b111 G
#912280000000
0!
0*
09
0>
0C
#912290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#912300000000
0!
0*
09
0>
0C
#912310000000
1!
1*
b1 6
19
1>
1C
b1 G
#912320000000
0!
0*
09
0>
0C
#912330000000
1!
1*
b10 6
19
1>
1C
b10 G
#912340000000
0!
0*
09
0>
0C
#912350000000
1!
1*
b11 6
19
1>
1C
b11 G
#912360000000
0!
0*
09
0>
0C
#912370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#912380000000
0!
0*
09
0>
0C
#912390000000
1!
1*
b101 6
19
1>
1C
b101 G
#912400000000
0!
0*
09
0>
0C
#912410000000
1!
1*
b110 6
19
1>
1C
b110 G
#912420000000
0!
0*
09
0>
0C
#912430000000
1!
1*
b111 6
19
1>
1C
b111 G
#912440000000
0!
0*
09
0>
0C
#912450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#912460000000
0!
0*
09
0>
0C
#912470000000
1!
1*
b1 6
19
1>
1C
b1 G
#912480000000
0!
0*
09
0>
0C
#912490000000
1!
1*
b10 6
19
1>
1C
b10 G
#912500000000
0!
0*
09
0>
0C
#912510000000
1!
1*
b11 6
19
1>
1C
b11 G
#912520000000
0!
0*
09
0>
0C
#912530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#912540000000
0!
0*
09
0>
0C
#912550000000
1!
1*
b101 6
19
1>
1C
b101 G
#912560000000
0!
0*
09
0>
0C
#912570000000
1!
1*
b110 6
19
1>
1C
b110 G
#912580000000
0!
0*
09
0>
0C
#912590000000
1!
1*
b111 6
19
1>
1C
b111 G
#912600000000
0!
1"
0*
1+
09
1:
0>
0C
#912610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#912620000000
0!
0*
09
0>
0C
#912630000000
1!
1*
b1 6
19
1>
1C
b1 G
#912640000000
0!
0*
09
0>
0C
#912650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#912660000000
0!
0*
09
0>
0C
#912670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#912680000000
0!
0*
09
0>
0C
#912690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#912700000000
0!
0*
09
0>
0C
#912710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#912720000000
0!
0#
0*
0,
09
0>
0?
0C
#912730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#912740000000
0!
0*
09
0>
0C
#912750000000
1!
1*
19
1>
1C
#912760000000
0!
0*
09
0>
0C
#912770000000
1!
1*
19
1>
1C
#912780000000
0!
0*
09
0>
0C
#912790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#912800000000
0!
0*
09
0>
0C
#912810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#912820000000
0!
0*
09
0>
0C
#912830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#912840000000
0!
0*
09
0>
0C
#912850000000
1!
1*
b10 6
19
1>
1C
b10 G
#912860000000
0!
0*
09
0>
0C
#912870000000
1!
1*
b11 6
19
1>
1C
b11 G
#912880000000
0!
0*
09
0>
0C
#912890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#912900000000
0!
0*
09
0>
0C
#912910000000
1!
1*
b101 6
19
1>
1C
b101 G
#912920000000
0!
0*
09
0>
0C
#912930000000
1!
1*
b110 6
19
1>
1C
b110 G
#912940000000
0!
0*
09
0>
0C
#912950000000
1!
1*
b111 6
19
1>
1C
b111 G
#912960000000
0!
0*
09
0>
0C
#912970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#912980000000
0!
0*
09
0>
0C
#912990000000
1!
1*
b1 6
19
1>
1C
b1 G
#913000000000
0!
0*
09
0>
0C
#913010000000
1!
1*
b10 6
19
1>
1C
b10 G
#913020000000
0!
0*
09
0>
0C
#913030000000
1!
1*
b11 6
19
1>
1C
b11 G
#913040000000
0!
0*
09
0>
0C
#913050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#913060000000
0!
0*
09
0>
0C
#913070000000
1!
1*
b101 6
19
1>
1C
b101 G
#913080000000
0!
0*
09
0>
0C
#913090000000
1!
1*
b110 6
19
1>
1C
b110 G
#913100000000
0!
0*
09
0>
0C
#913110000000
1!
1*
b111 6
19
1>
1C
b111 G
#913120000000
0!
0*
09
0>
0C
#913130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#913140000000
0!
0*
09
0>
0C
#913150000000
1!
1*
b1 6
19
1>
1C
b1 G
#913160000000
0!
0*
09
0>
0C
#913170000000
1!
1*
b10 6
19
1>
1C
b10 G
#913180000000
0!
0*
09
0>
0C
#913190000000
1!
1*
b11 6
19
1>
1C
b11 G
#913200000000
0!
0*
09
0>
0C
#913210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#913220000000
0!
0*
09
0>
0C
#913230000000
1!
1*
b101 6
19
1>
1C
b101 G
#913240000000
0!
0*
09
0>
0C
#913250000000
1!
1*
b110 6
19
1>
1C
b110 G
#913260000000
0!
0*
09
0>
0C
#913270000000
1!
1*
b111 6
19
1>
1C
b111 G
#913280000000
0!
1"
0*
1+
09
1:
0>
0C
#913290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#913300000000
0!
0*
09
0>
0C
#913310000000
1!
1*
b1 6
19
1>
1C
b1 G
#913320000000
0!
0*
09
0>
0C
#913330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#913340000000
0!
0*
09
0>
0C
#913350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#913360000000
0!
0*
09
0>
0C
#913370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#913380000000
0!
0*
09
0>
0C
#913390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#913400000000
0!
0#
0*
0,
09
0>
0?
0C
#913410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#913420000000
0!
0*
09
0>
0C
#913430000000
1!
1*
19
1>
1C
#913440000000
0!
0*
09
0>
0C
#913450000000
1!
1*
19
1>
1C
#913460000000
0!
0*
09
0>
0C
#913470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#913480000000
0!
0*
09
0>
0C
#913490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#913500000000
0!
0*
09
0>
0C
#913510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#913520000000
0!
0*
09
0>
0C
#913530000000
1!
1*
b10 6
19
1>
1C
b10 G
#913540000000
0!
0*
09
0>
0C
#913550000000
1!
1*
b11 6
19
1>
1C
b11 G
#913560000000
0!
0*
09
0>
0C
#913570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#913580000000
0!
0*
09
0>
0C
#913590000000
1!
1*
b101 6
19
1>
1C
b101 G
#913600000000
0!
0*
09
0>
0C
#913610000000
1!
1*
b110 6
19
1>
1C
b110 G
#913620000000
0!
0*
09
0>
0C
#913630000000
1!
1*
b111 6
19
1>
1C
b111 G
#913640000000
0!
0*
09
0>
0C
#913650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#913660000000
0!
0*
09
0>
0C
#913670000000
1!
1*
b1 6
19
1>
1C
b1 G
#913680000000
0!
0*
09
0>
0C
#913690000000
1!
1*
b10 6
19
1>
1C
b10 G
#913700000000
0!
0*
09
0>
0C
#913710000000
1!
1*
b11 6
19
1>
1C
b11 G
#913720000000
0!
0*
09
0>
0C
#913730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#913740000000
0!
0*
09
0>
0C
#913750000000
1!
1*
b101 6
19
1>
1C
b101 G
#913760000000
0!
0*
09
0>
0C
#913770000000
1!
1*
b110 6
19
1>
1C
b110 G
#913780000000
0!
0*
09
0>
0C
#913790000000
1!
1*
b111 6
19
1>
1C
b111 G
#913800000000
0!
0*
09
0>
0C
#913810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#913820000000
0!
0*
09
0>
0C
#913830000000
1!
1*
b1 6
19
1>
1C
b1 G
#913840000000
0!
0*
09
0>
0C
#913850000000
1!
1*
b10 6
19
1>
1C
b10 G
#913860000000
0!
0*
09
0>
0C
#913870000000
1!
1*
b11 6
19
1>
1C
b11 G
#913880000000
0!
0*
09
0>
0C
#913890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#913900000000
0!
0*
09
0>
0C
#913910000000
1!
1*
b101 6
19
1>
1C
b101 G
#913920000000
0!
0*
09
0>
0C
#913930000000
1!
1*
b110 6
19
1>
1C
b110 G
#913940000000
0!
0*
09
0>
0C
#913950000000
1!
1*
b111 6
19
1>
1C
b111 G
#913960000000
0!
1"
0*
1+
09
1:
0>
0C
#913970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#913980000000
0!
0*
09
0>
0C
#913990000000
1!
1*
b1 6
19
1>
1C
b1 G
#914000000000
0!
0*
09
0>
0C
#914010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#914020000000
0!
0*
09
0>
0C
#914030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#914040000000
0!
0*
09
0>
0C
#914050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#914060000000
0!
0*
09
0>
0C
#914070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#914080000000
0!
0#
0*
0,
09
0>
0?
0C
#914090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#914100000000
0!
0*
09
0>
0C
#914110000000
1!
1*
19
1>
1C
#914120000000
0!
0*
09
0>
0C
#914130000000
1!
1*
19
1>
1C
#914140000000
0!
0*
09
0>
0C
#914150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#914160000000
0!
0*
09
0>
0C
#914170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#914180000000
0!
0*
09
0>
0C
#914190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#914200000000
0!
0*
09
0>
0C
#914210000000
1!
1*
b10 6
19
1>
1C
b10 G
#914220000000
0!
0*
09
0>
0C
#914230000000
1!
1*
b11 6
19
1>
1C
b11 G
#914240000000
0!
0*
09
0>
0C
#914250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#914260000000
0!
0*
09
0>
0C
#914270000000
1!
1*
b101 6
19
1>
1C
b101 G
#914280000000
0!
0*
09
0>
0C
#914290000000
1!
1*
b110 6
19
1>
1C
b110 G
#914300000000
0!
0*
09
0>
0C
#914310000000
1!
1*
b111 6
19
1>
1C
b111 G
#914320000000
0!
0*
09
0>
0C
#914330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#914340000000
0!
0*
09
0>
0C
#914350000000
1!
1*
b1 6
19
1>
1C
b1 G
#914360000000
0!
0*
09
0>
0C
#914370000000
1!
1*
b10 6
19
1>
1C
b10 G
#914380000000
0!
0*
09
0>
0C
#914390000000
1!
1*
b11 6
19
1>
1C
b11 G
#914400000000
0!
0*
09
0>
0C
#914410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#914420000000
0!
0*
09
0>
0C
#914430000000
1!
1*
b101 6
19
1>
1C
b101 G
#914440000000
0!
0*
09
0>
0C
#914450000000
1!
1*
b110 6
19
1>
1C
b110 G
#914460000000
0!
0*
09
0>
0C
#914470000000
1!
1*
b111 6
19
1>
1C
b111 G
#914480000000
0!
0*
09
0>
0C
#914490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#914500000000
0!
0*
09
0>
0C
#914510000000
1!
1*
b1 6
19
1>
1C
b1 G
#914520000000
0!
0*
09
0>
0C
#914530000000
1!
1*
b10 6
19
1>
1C
b10 G
#914540000000
0!
0*
09
0>
0C
#914550000000
1!
1*
b11 6
19
1>
1C
b11 G
#914560000000
0!
0*
09
0>
0C
#914570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#914580000000
0!
0*
09
0>
0C
#914590000000
1!
1*
b101 6
19
1>
1C
b101 G
#914600000000
0!
0*
09
0>
0C
#914610000000
1!
1*
b110 6
19
1>
1C
b110 G
#914620000000
0!
0*
09
0>
0C
#914630000000
1!
1*
b111 6
19
1>
1C
b111 G
#914640000000
0!
1"
0*
1+
09
1:
0>
0C
#914650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#914660000000
0!
0*
09
0>
0C
#914670000000
1!
1*
b1 6
19
1>
1C
b1 G
#914680000000
0!
0*
09
0>
0C
#914690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#914700000000
0!
0*
09
0>
0C
#914710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#914720000000
0!
0*
09
0>
0C
#914730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#914740000000
0!
0*
09
0>
0C
#914750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#914760000000
0!
0#
0*
0,
09
0>
0?
0C
#914770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#914780000000
0!
0*
09
0>
0C
#914790000000
1!
1*
19
1>
1C
#914800000000
0!
0*
09
0>
0C
#914810000000
1!
1*
19
1>
1C
#914820000000
0!
0*
09
0>
0C
#914830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#914840000000
0!
0*
09
0>
0C
#914850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#914860000000
0!
0*
09
0>
0C
#914870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#914880000000
0!
0*
09
0>
0C
#914890000000
1!
1*
b10 6
19
1>
1C
b10 G
#914900000000
0!
0*
09
0>
0C
#914910000000
1!
1*
b11 6
19
1>
1C
b11 G
#914920000000
0!
0*
09
0>
0C
#914930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#914940000000
0!
0*
09
0>
0C
#914950000000
1!
1*
b101 6
19
1>
1C
b101 G
#914960000000
0!
0*
09
0>
0C
#914970000000
1!
1*
b110 6
19
1>
1C
b110 G
#914980000000
0!
0*
09
0>
0C
#914990000000
1!
1*
b111 6
19
1>
1C
b111 G
#915000000000
0!
0*
09
0>
0C
#915010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#915020000000
0!
0*
09
0>
0C
#915030000000
1!
1*
b1 6
19
1>
1C
b1 G
#915040000000
0!
0*
09
0>
0C
#915050000000
1!
1*
b10 6
19
1>
1C
b10 G
#915060000000
0!
0*
09
0>
0C
#915070000000
1!
1*
b11 6
19
1>
1C
b11 G
#915080000000
0!
0*
09
0>
0C
#915090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#915100000000
0!
0*
09
0>
0C
#915110000000
1!
1*
b101 6
19
1>
1C
b101 G
#915120000000
0!
0*
09
0>
0C
#915130000000
1!
1*
b110 6
19
1>
1C
b110 G
#915140000000
0!
0*
09
0>
0C
#915150000000
1!
1*
b111 6
19
1>
1C
b111 G
#915160000000
0!
0*
09
0>
0C
#915170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#915180000000
0!
0*
09
0>
0C
#915190000000
1!
1*
b1 6
19
1>
1C
b1 G
#915200000000
0!
0*
09
0>
0C
#915210000000
1!
1*
b10 6
19
1>
1C
b10 G
#915220000000
0!
0*
09
0>
0C
#915230000000
1!
1*
b11 6
19
1>
1C
b11 G
#915240000000
0!
0*
09
0>
0C
#915250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#915260000000
0!
0*
09
0>
0C
#915270000000
1!
1*
b101 6
19
1>
1C
b101 G
#915280000000
0!
0*
09
0>
0C
#915290000000
1!
1*
b110 6
19
1>
1C
b110 G
#915300000000
0!
0*
09
0>
0C
#915310000000
1!
1*
b111 6
19
1>
1C
b111 G
#915320000000
0!
1"
0*
1+
09
1:
0>
0C
#915330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#915340000000
0!
0*
09
0>
0C
#915350000000
1!
1*
b1 6
19
1>
1C
b1 G
#915360000000
0!
0*
09
0>
0C
#915370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#915380000000
0!
0*
09
0>
0C
#915390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#915400000000
0!
0*
09
0>
0C
#915410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#915420000000
0!
0*
09
0>
0C
#915430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#915440000000
0!
0#
0*
0,
09
0>
0?
0C
#915450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#915460000000
0!
0*
09
0>
0C
#915470000000
1!
1*
19
1>
1C
#915480000000
0!
0*
09
0>
0C
#915490000000
1!
1*
19
1>
1C
#915500000000
0!
0*
09
0>
0C
#915510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#915520000000
0!
0*
09
0>
0C
#915530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#915540000000
0!
0*
09
0>
0C
#915550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#915560000000
0!
0*
09
0>
0C
#915570000000
1!
1*
b10 6
19
1>
1C
b10 G
#915580000000
0!
0*
09
0>
0C
#915590000000
1!
1*
b11 6
19
1>
1C
b11 G
#915600000000
0!
0*
09
0>
0C
#915610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#915620000000
0!
0*
09
0>
0C
#915630000000
1!
1*
b101 6
19
1>
1C
b101 G
#915640000000
0!
0*
09
0>
0C
#915650000000
1!
1*
b110 6
19
1>
1C
b110 G
#915660000000
0!
0*
09
0>
0C
#915670000000
1!
1*
b111 6
19
1>
1C
b111 G
#915680000000
0!
0*
09
0>
0C
#915690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#915700000000
0!
0*
09
0>
0C
#915710000000
1!
1*
b1 6
19
1>
1C
b1 G
#915720000000
0!
0*
09
0>
0C
#915730000000
1!
1*
b10 6
19
1>
1C
b10 G
#915740000000
0!
0*
09
0>
0C
#915750000000
1!
1*
b11 6
19
1>
1C
b11 G
#915760000000
0!
0*
09
0>
0C
#915770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#915780000000
0!
0*
09
0>
0C
#915790000000
1!
1*
b101 6
19
1>
1C
b101 G
#915800000000
0!
0*
09
0>
0C
#915810000000
1!
1*
b110 6
19
1>
1C
b110 G
#915820000000
0!
0*
09
0>
0C
#915830000000
1!
1*
b111 6
19
1>
1C
b111 G
#915840000000
0!
0*
09
0>
0C
#915850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#915860000000
0!
0*
09
0>
0C
#915870000000
1!
1*
b1 6
19
1>
1C
b1 G
#915880000000
0!
0*
09
0>
0C
#915890000000
1!
1*
b10 6
19
1>
1C
b10 G
#915900000000
0!
0*
09
0>
0C
#915910000000
1!
1*
b11 6
19
1>
1C
b11 G
#915920000000
0!
0*
09
0>
0C
#915930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#915940000000
0!
0*
09
0>
0C
#915950000000
1!
1*
b101 6
19
1>
1C
b101 G
#915960000000
0!
0*
09
0>
0C
#915970000000
1!
1*
b110 6
19
1>
1C
b110 G
#915980000000
0!
0*
09
0>
0C
#915990000000
1!
1*
b111 6
19
1>
1C
b111 G
#916000000000
0!
1"
0*
1+
09
1:
0>
0C
#916010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#916020000000
0!
0*
09
0>
0C
#916030000000
1!
1*
b1 6
19
1>
1C
b1 G
#916040000000
0!
0*
09
0>
0C
#916050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#916060000000
0!
0*
09
0>
0C
#916070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#916080000000
0!
0*
09
0>
0C
#916090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#916100000000
0!
0*
09
0>
0C
#916110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#916120000000
0!
0#
0*
0,
09
0>
0?
0C
#916130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#916140000000
0!
0*
09
0>
0C
#916150000000
1!
1*
19
1>
1C
#916160000000
0!
0*
09
0>
0C
#916170000000
1!
1*
19
1>
1C
#916180000000
0!
0*
09
0>
0C
#916190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#916200000000
0!
0*
09
0>
0C
#916210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#916220000000
0!
0*
09
0>
0C
#916230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#916240000000
0!
0*
09
0>
0C
#916250000000
1!
1*
b10 6
19
1>
1C
b10 G
#916260000000
0!
0*
09
0>
0C
#916270000000
1!
1*
b11 6
19
1>
1C
b11 G
#916280000000
0!
0*
09
0>
0C
#916290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#916300000000
0!
0*
09
0>
0C
#916310000000
1!
1*
b101 6
19
1>
1C
b101 G
#916320000000
0!
0*
09
0>
0C
#916330000000
1!
1*
b110 6
19
1>
1C
b110 G
#916340000000
0!
0*
09
0>
0C
#916350000000
1!
1*
b111 6
19
1>
1C
b111 G
#916360000000
0!
0*
09
0>
0C
#916370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#916380000000
0!
0*
09
0>
0C
#916390000000
1!
1*
b1 6
19
1>
1C
b1 G
#916400000000
0!
0*
09
0>
0C
#916410000000
1!
1*
b10 6
19
1>
1C
b10 G
#916420000000
0!
0*
09
0>
0C
#916430000000
1!
1*
b11 6
19
1>
1C
b11 G
#916440000000
0!
0*
09
0>
0C
#916450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#916460000000
0!
0*
09
0>
0C
#916470000000
1!
1*
b101 6
19
1>
1C
b101 G
#916480000000
0!
0*
09
0>
0C
#916490000000
1!
1*
b110 6
19
1>
1C
b110 G
#916500000000
0!
0*
09
0>
0C
#916510000000
1!
1*
b111 6
19
1>
1C
b111 G
#916520000000
0!
0*
09
0>
0C
#916530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#916540000000
0!
0*
09
0>
0C
#916550000000
1!
1*
b1 6
19
1>
1C
b1 G
#916560000000
0!
0*
09
0>
0C
#916570000000
1!
1*
b10 6
19
1>
1C
b10 G
#916580000000
0!
0*
09
0>
0C
#916590000000
1!
1*
b11 6
19
1>
1C
b11 G
#916600000000
0!
0*
09
0>
0C
#916610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#916620000000
0!
0*
09
0>
0C
#916630000000
1!
1*
b101 6
19
1>
1C
b101 G
#916640000000
0!
0*
09
0>
0C
#916650000000
1!
1*
b110 6
19
1>
1C
b110 G
#916660000000
0!
0*
09
0>
0C
#916670000000
1!
1*
b111 6
19
1>
1C
b111 G
#916680000000
0!
1"
0*
1+
09
1:
0>
0C
#916690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#916700000000
0!
0*
09
0>
0C
#916710000000
1!
1*
b1 6
19
1>
1C
b1 G
#916720000000
0!
0*
09
0>
0C
#916730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#916740000000
0!
0*
09
0>
0C
#916750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#916760000000
0!
0*
09
0>
0C
#916770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#916780000000
0!
0*
09
0>
0C
#916790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#916800000000
0!
0#
0*
0,
09
0>
0?
0C
#916810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#916820000000
0!
0*
09
0>
0C
#916830000000
1!
1*
19
1>
1C
#916840000000
0!
0*
09
0>
0C
#916850000000
1!
1*
19
1>
1C
#916860000000
0!
0*
09
0>
0C
#916870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#916880000000
0!
0*
09
0>
0C
#916890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#916900000000
0!
0*
09
0>
0C
#916910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#916920000000
0!
0*
09
0>
0C
#916930000000
1!
1*
b10 6
19
1>
1C
b10 G
#916940000000
0!
0*
09
0>
0C
#916950000000
1!
1*
b11 6
19
1>
1C
b11 G
#916960000000
0!
0*
09
0>
0C
#916970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#916980000000
0!
0*
09
0>
0C
#916990000000
1!
1*
b101 6
19
1>
1C
b101 G
#917000000000
0!
0*
09
0>
0C
#917010000000
1!
1*
b110 6
19
1>
1C
b110 G
#917020000000
0!
0*
09
0>
0C
#917030000000
1!
1*
b111 6
19
1>
1C
b111 G
#917040000000
0!
0*
09
0>
0C
#917050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#917060000000
0!
0*
09
0>
0C
#917070000000
1!
1*
b1 6
19
1>
1C
b1 G
#917080000000
0!
0*
09
0>
0C
#917090000000
1!
1*
b10 6
19
1>
1C
b10 G
#917100000000
0!
0*
09
0>
0C
#917110000000
1!
1*
b11 6
19
1>
1C
b11 G
#917120000000
0!
0*
09
0>
0C
#917130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#917140000000
0!
0*
09
0>
0C
#917150000000
1!
1*
b101 6
19
1>
1C
b101 G
#917160000000
0!
0*
09
0>
0C
#917170000000
1!
1*
b110 6
19
1>
1C
b110 G
#917180000000
0!
0*
09
0>
0C
#917190000000
1!
1*
b111 6
19
1>
1C
b111 G
#917200000000
0!
0*
09
0>
0C
#917210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#917220000000
0!
0*
09
0>
0C
#917230000000
1!
1*
b1 6
19
1>
1C
b1 G
#917240000000
0!
0*
09
0>
0C
#917250000000
1!
1*
b10 6
19
1>
1C
b10 G
#917260000000
0!
0*
09
0>
0C
#917270000000
1!
1*
b11 6
19
1>
1C
b11 G
#917280000000
0!
0*
09
0>
0C
#917290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#917300000000
0!
0*
09
0>
0C
#917310000000
1!
1*
b101 6
19
1>
1C
b101 G
#917320000000
0!
0*
09
0>
0C
#917330000000
1!
1*
b110 6
19
1>
1C
b110 G
#917340000000
0!
0*
09
0>
0C
#917350000000
1!
1*
b111 6
19
1>
1C
b111 G
#917360000000
0!
1"
0*
1+
09
1:
0>
0C
#917370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#917380000000
0!
0*
09
0>
0C
#917390000000
1!
1*
b1 6
19
1>
1C
b1 G
#917400000000
0!
0*
09
0>
0C
#917410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#917420000000
0!
0*
09
0>
0C
#917430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#917440000000
0!
0*
09
0>
0C
#917450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#917460000000
0!
0*
09
0>
0C
#917470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#917480000000
0!
0#
0*
0,
09
0>
0?
0C
#917490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#917500000000
0!
0*
09
0>
0C
#917510000000
1!
1*
19
1>
1C
#917520000000
0!
0*
09
0>
0C
#917530000000
1!
1*
19
1>
1C
#917540000000
0!
0*
09
0>
0C
#917550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#917560000000
0!
0*
09
0>
0C
#917570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#917580000000
0!
0*
09
0>
0C
#917590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#917600000000
0!
0*
09
0>
0C
#917610000000
1!
1*
b10 6
19
1>
1C
b10 G
#917620000000
0!
0*
09
0>
0C
#917630000000
1!
1*
b11 6
19
1>
1C
b11 G
#917640000000
0!
0*
09
0>
0C
#917650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#917660000000
0!
0*
09
0>
0C
#917670000000
1!
1*
b101 6
19
1>
1C
b101 G
#917680000000
0!
0*
09
0>
0C
#917690000000
1!
1*
b110 6
19
1>
1C
b110 G
#917700000000
0!
0*
09
0>
0C
#917710000000
1!
1*
b111 6
19
1>
1C
b111 G
#917720000000
0!
0*
09
0>
0C
#917730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#917740000000
0!
0*
09
0>
0C
#917750000000
1!
1*
b1 6
19
1>
1C
b1 G
#917760000000
0!
0*
09
0>
0C
#917770000000
1!
1*
b10 6
19
1>
1C
b10 G
#917780000000
0!
0*
09
0>
0C
#917790000000
1!
1*
b11 6
19
1>
1C
b11 G
#917800000000
0!
0*
09
0>
0C
#917810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#917820000000
0!
0*
09
0>
0C
#917830000000
1!
1*
b101 6
19
1>
1C
b101 G
#917840000000
0!
0*
09
0>
0C
#917850000000
1!
1*
b110 6
19
1>
1C
b110 G
#917860000000
0!
0*
09
0>
0C
#917870000000
1!
1*
b111 6
19
1>
1C
b111 G
#917880000000
0!
0*
09
0>
0C
#917890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#917900000000
0!
0*
09
0>
0C
#917910000000
1!
1*
b1 6
19
1>
1C
b1 G
#917920000000
0!
0*
09
0>
0C
#917930000000
1!
1*
b10 6
19
1>
1C
b10 G
#917940000000
0!
0*
09
0>
0C
#917950000000
1!
1*
b11 6
19
1>
1C
b11 G
#917960000000
0!
0*
09
0>
0C
#917970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#917980000000
0!
0*
09
0>
0C
#917990000000
1!
1*
b101 6
19
1>
1C
b101 G
#918000000000
0!
0*
09
0>
0C
#918010000000
1!
1*
b110 6
19
1>
1C
b110 G
#918020000000
0!
0*
09
0>
0C
#918030000000
1!
1*
b111 6
19
1>
1C
b111 G
#918040000000
0!
1"
0*
1+
09
1:
0>
0C
#918050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#918060000000
0!
0*
09
0>
0C
#918070000000
1!
1*
b1 6
19
1>
1C
b1 G
#918080000000
0!
0*
09
0>
0C
#918090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#918100000000
0!
0*
09
0>
0C
#918110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#918120000000
0!
0*
09
0>
0C
#918130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#918140000000
0!
0*
09
0>
0C
#918150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#918160000000
0!
0#
0*
0,
09
0>
0?
0C
#918170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#918180000000
0!
0*
09
0>
0C
#918190000000
1!
1*
19
1>
1C
#918200000000
0!
0*
09
0>
0C
#918210000000
1!
1*
19
1>
1C
#918220000000
0!
0*
09
0>
0C
#918230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#918240000000
0!
0*
09
0>
0C
#918250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#918260000000
0!
0*
09
0>
0C
#918270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#918280000000
0!
0*
09
0>
0C
#918290000000
1!
1*
b10 6
19
1>
1C
b10 G
#918300000000
0!
0*
09
0>
0C
#918310000000
1!
1*
b11 6
19
1>
1C
b11 G
#918320000000
0!
0*
09
0>
0C
#918330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#918340000000
0!
0*
09
0>
0C
#918350000000
1!
1*
b101 6
19
1>
1C
b101 G
#918360000000
0!
0*
09
0>
0C
#918370000000
1!
1*
b110 6
19
1>
1C
b110 G
#918380000000
0!
0*
09
0>
0C
#918390000000
1!
1*
b111 6
19
1>
1C
b111 G
#918400000000
0!
0*
09
0>
0C
#918410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#918420000000
0!
0*
09
0>
0C
#918430000000
1!
1*
b1 6
19
1>
1C
b1 G
#918440000000
0!
0*
09
0>
0C
#918450000000
1!
1*
b10 6
19
1>
1C
b10 G
#918460000000
0!
0*
09
0>
0C
#918470000000
1!
1*
b11 6
19
1>
1C
b11 G
#918480000000
0!
0*
09
0>
0C
#918490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#918500000000
0!
0*
09
0>
0C
#918510000000
1!
1*
b101 6
19
1>
1C
b101 G
#918520000000
0!
0*
09
0>
0C
#918530000000
1!
1*
b110 6
19
1>
1C
b110 G
#918540000000
0!
0*
09
0>
0C
#918550000000
1!
1*
b111 6
19
1>
1C
b111 G
#918560000000
0!
0*
09
0>
0C
#918570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#918580000000
0!
0*
09
0>
0C
#918590000000
1!
1*
b1 6
19
1>
1C
b1 G
#918600000000
0!
0*
09
0>
0C
#918610000000
1!
1*
b10 6
19
1>
1C
b10 G
#918620000000
0!
0*
09
0>
0C
#918630000000
1!
1*
b11 6
19
1>
1C
b11 G
#918640000000
0!
0*
09
0>
0C
#918650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#918660000000
0!
0*
09
0>
0C
#918670000000
1!
1*
b101 6
19
1>
1C
b101 G
#918680000000
0!
0*
09
0>
0C
#918690000000
1!
1*
b110 6
19
1>
1C
b110 G
#918700000000
0!
0*
09
0>
0C
#918710000000
1!
1*
b111 6
19
1>
1C
b111 G
#918720000000
0!
1"
0*
1+
09
1:
0>
0C
#918730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#918740000000
0!
0*
09
0>
0C
#918750000000
1!
1*
b1 6
19
1>
1C
b1 G
#918760000000
0!
0*
09
0>
0C
#918770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#918780000000
0!
0*
09
0>
0C
#918790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#918800000000
0!
0*
09
0>
0C
#918810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#918820000000
0!
0*
09
0>
0C
#918830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#918840000000
0!
0#
0*
0,
09
0>
0?
0C
#918850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#918860000000
0!
0*
09
0>
0C
#918870000000
1!
1*
19
1>
1C
#918880000000
0!
0*
09
0>
0C
#918890000000
1!
1*
19
1>
1C
#918900000000
0!
0*
09
0>
0C
#918910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#918920000000
0!
0*
09
0>
0C
#918930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#918940000000
0!
0*
09
0>
0C
#918950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#918960000000
0!
0*
09
0>
0C
#918970000000
1!
1*
b10 6
19
1>
1C
b10 G
#918980000000
0!
0*
09
0>
0C
#918990000000
1!
1*
b11 6
19
1>
1C
b11 G
#919000000000
0!
0*
09
0>
0C
#919010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#919020000000
0!
0*
09
0>
0C
#919030000000
1!
1*
b101 6
19
1>
1C
b101 G
#919040000000
0!
0*
09
0>
0C
#919050000000
1!
1*
b110 6
19
1>
1C
b110 G
#919060000000
0!
0*
09
0>
0C
#919070000000
1!
1*
b111 6
19
1>
1C
b111 G
#919080000000
0!
0*
09
0>
0C
#919090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#919100000000
0!
0*
09
0>
0C
#919110000000
1!
1*
b1 6
19
1>
1C
b1 G
#919120000000
0!
0*
09
0>
0C
#919130000000
1!
1*
b10 6
19
1>
1C
b10 G
#919140000000
0!
0*
09
0>
0C
#919150000000
1!
1*
b11 6
19
1>
1C
b11 G
#919160000000
0!
0*
09
0>
0C
#919170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#919180000000
0!
0*
09
0>
0C
#919190000000
1!
1*
b101 6
19
1>
1C
b101 G
#919200000000
0!
0*
09
0>
0C
#919210000000
1!
1*
b110 6
19
1>
1C
b110 G
#919220000000
0!
0*
09
0>
0C
#919230000000
1!
1*
b111 6
19
1>
1C
b111 G
#919240000000
0!
0*
09
0>
0C
#919250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#919260000000
0!
0*
09
0>
0C
#919270000000
1!
1*
b1 6
19
1>
1C
b1 G
#919280000000
0!
0*
09
0>
0C
#919290000000
1!
1*
b10 6
19
1>
1C
b10 G
#919300000000
0!
0*
09
0>
0C
#919310000000
1!
1*
b11 6
19
1>
1C
b11 G
#919320000000
0!
0*
09
0>
0C
#919330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#919340000000
0!
0*
09
0>
0C
#919350000000
1!
1*
b101 6
19
1>
1C
b101 G
#919360000000
0!
0*
09
0>
0C
#919370000000
1!
1*
b110 6
19
1>
1C
b110 G
#919380000000
0!
0*
09
0>
0C
#919390000000
1!
1*
b111 6
19
1>
1C
b111 G
#919400000000
0!
1"
0*
1+
09
1:
0>
0C
#919410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#919420000000
0!
0*
09
0>
0C
#919430000000
1!
1*
b1 6
19
1>
1C
b1 G
#919440000000
0!
0*
09
0>
0C
#919450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#919460000000
0!
0*
09
0>
0C
#919470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#919480000000
0!
0*
09
0>
0C
#919490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#919500000000
0!
0*
09
0>
0C
#919510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#919520000000
0!
0#
0*
0,
09
0>
0?
0C
#919530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#919540000000
0!
0*
09
0>
0C
#919550000000
1!
1*
19
1>
1C
#919560000000
0!
0*
09
0>
0C
#919570000000
1!
1*
19
1>
1C
#919580000000
0!
0*
09
0>
0C
#919590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#919600000000
0!
0*
09
0>
0C
#919610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#919620000000
0!
0*
09
0>
0C
#919630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#919640000000
0!
0*
09
0>
0C
#919650000000
1!
1*
b10 6
19
1>
1C
b10 G
#919660000000
0!
0*
09
0>
0C
#919670000000
1!
1*
b11 6
19
1>
1C
b11 G
#919680000000
0!
0*
09
0>
0C
#919690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#919700000000
0!
0*
09
0>
0C
#919710000000
1!
1*
b101 6
19
1>
1C
b101 G
#919720000000
0!
0*
09
0>
0C
#919730000000
1!
1*
b110 6
19
1>
1C
b110 G
#919740000000
0!
0*
09
0>
0C
#919750000000
1!
1*
b111 6
19
1>
1C
b111 G
#919760000000
0!
0*
09
0>
0C
#919770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#919780000000
0!
0*
09
0>
0C
#919790000000
1!
1*
b1 6
19
1>
1C
b1 G
#919800000000
0!
0*
09
0>
0C
#919810000000
1!
1*
b10 6
19
1>
1C
b10 G
#919820000000
0!
0*
09
0>
0C
#919830000000
1!
1*
b11 6
19
1>
1C
b11 G
#919840000000
0!
0*
09
0>
0C
#919850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#919860000000
0!
0*
09
0>
0C
#919870000000
1!
1*
b101 6
19
1>
1C
b101 G
#919880000000
0!
0*
09
0>
0C
#919890000000
1!
1*
b110 6
19
1>
1C
b110 G
#919900000000
0!
0*
09
0>
0C
#919910000000
1!
1*
b111 6
19
1>
1C
b111 G
#919920000000
0!
0*
09
0>
0C
#919930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#919940000000
0!
0*
09
0>
0C
#919950000000
1!
1*
b1 6
19
1>
1C
b1 G
#919960000000
0!
0*
09
0>
0C
#919970000000
1!
1*
b10 6
19
1>
1C
b10 G
#919980000000
0!
0*
09
0>
0C
#919990000000
1!
1*
b11 6
19
1>
1C
b11 G
#920000000000
0!
0*
09
0>
0C
#920010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#920020000000
0!
0*
09
0>
0C
#920030000000
1!
1*
b101 6
19
1>
1C
b101 G
#920040000000
0!
0*
09
0>
0C
#920050000000
1!
1*
b110 6
19
1>
1C
b110 G
#920060000000
0!
0*
09
0>
0C
#920070000000
1!
1*
b111 6
19
1>
1C
b111 G
#920080000000
0!
1"
0*
1+
09
1:
0>
0C
#920090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#920100000000
0!
0*
09
0>
0C
#920110000000
1!
1*
b1 6
19
1>
1C
b1 G
#920120000000
0!
0*
09
0>
0C
#920130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#920140000000
0!
0*
09
0>
0C
#920150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#920160000000
0!
0*
09
0>
0C
#920170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#920180000000
0!
0*
09
0>
0C
#920190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#920200000000
0!
0#
0*
0,
09
0>
0?
0C
#920210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#920220000000
0!
0*
09
0>
0C
#920230000000
1!
1*
19
1>
1C
#920240000000
0!
0*
09
0>
0C
#920250000000
1!
1*
19
1>
1C
#920260000000
0!
0*
09
0>
0C
#920270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#920280000000
0!
0*
09
0>
0C
#920290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#920300000000
0!
0*
09
0>
0C
#920310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#920320000000
0!
0*
09
0>
0C
#920330000000
1!
1*
b10 6
19
1>
1C
b10 G
#920340000000
0!
0*
09
0>
0C
#920350000000
1!
1*
b11 6
19
1>
1C
b11 G
#920360000000
0!
0*
09
0>
0C
#920370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#920380000000
0!
0*
09
0>
0C
#920390000000
1!
1*
b101 6
19
1>
1C
b101 G
#920400000000
0!
0*
09
0>
0C
#920410000000
1!
1*
b110 6
19
1>
1C
b110 G
#920420000000
0!
0*
09
0>
0C
#920430000000
1!
1*
b111 6
19
1>
1C
b111 G
#920440000000
0!
0*
09
0>
0C
#920450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#920460000000
0!
0*
09
0>
0C
#920470000000
1!
1*
b1 6
19
1>
1C
b1 G
#920480000000
0!
0*
09
0>
0C
#920490000000
1!
1*
b10 6
19
1>
1C
b10 G
#920500000000
0!
0*
09
0>
0C
#920510000000
1!
1*
b11 6
19
1>
1C
b11 G
#920520000000
0!
0*
09
0>
0C
#920530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#920540000000
0!
0*
09
0>
0C
#920550000000
1!
1*
b101 6
19
1>
1C
b101 G
#920560000000
0!
0*
09
0>
0C
#920570000000
1!
1*
b110 6
19
1>
1C
b110 G
#920580000000
0!
0*
09
0>
0C
#920590000000
1!
1*
b111 6
19
1>
1C
b111 G
#920600000000
0!
0*
09
0>
0C
#920610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#920620000000
0!
0*
09
0>
0C
#920630000000
1!
1*
b1 6
19
1>
1C
b1 G
#920640000000
0!
0*
09
0>
0C
#920650000000
1!
1*
b10 6
19
1>
1C
b10 G
#920660000000
0!
0*
09
0>
0C
#920670000000
1!
1*
b11 6
19
1>
1C
b11 G
#920680000000
0!
0*
09
0>
0C
#920690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#920700000000
0!
0*
09
0>
0C
#920710000000
1!
1*
b101 6
19
1>
1C
b101 G
#920720000000
0!
0*
09
0>
0C
#920730000000
1!
1*
b110 6
19
1>
1C
b110 G
#920740000000
0!
0*
09
0>
0C
#920750000000
1!
1*
b111 6
19
1>
1C
b111 G
#920760000000
0!
1"
0*
1+
09
1:
0>
0C
#920770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#920780000000
0!
0*
09
0>
0C
#920790000000
1!
1*
b1 6
19
1>
1C
b1 G
#920800000000
0!
0*
09
0>
0C
#920810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#920820000000
0!
0*
09
0>
0C
#920830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#920840000000
0!
0*
09
0>
0C
#920850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#920860000000
0!
0*
09
0>
0C
#920870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#920880000000
0!
0#
0*
0,
09
0>
0?
0C
#920890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#920900000000
0!
0*
09
0>
0C
#920910000000
1!
1*
19
1>
1C
#920920000000
0!
0*
09
0>
0C
#920930000000
1!
1*
19
1>
1C
#920940000000
0!
0*
09
0>
0C
#920950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#920960000000
0!
0*
09
0>
0C
#920970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#920980000000
0!
0*
09
0>
0C
#920990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#921000000000
0!
0*
09
0>
0C
#921010000000
1!
1*
b10 6
19
1>
1C
b10 G
#921020000000
0!
0*
09
0>
0C
#921030000000
1!
1*
b11 6
19
1>
1C
b11 G
#921040000000
0!
0*
09
0>
0C
#921050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#921060000000
0!
0*
09
0>
0C
#921070000000
1!
1*
b101 6
19
1>
1C
b101 G
#921080000000
0!
0*
09
0>
0C
#921090000000
1!
1*
b110 6
19
1>
1C
b110 G
#921100000000
0!
0*
09
0>
0C
#921110000000
1!
1*
b111 6
19
1>
1C
b111 G
#921120000000
0!
0*
09
0>
0C
#921130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#921140000000
0!
0*
09
0>
0C
#921150000000
1!
1*
b1 6
19
1>
1C
b1 G
#921160000000
0!
0*
09
0>
0C
#921170000000
1!
1*
b10 6
19
1>
1C
b10 G
#921180000000
0!
0*
09
0>
0C
#921190000000
1!
1*
b11 6
19
1>
1C
b11 G
#921200000000
0!
0*
09
0>
0C
#921210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#921220000000
0!
0*
09
0>
0C
#921230000000
1!
1*
b101 6
19
1>
1C
b101 G
#921240000000
0!
0*
09
0>
0C
#921250000000
1!
1*
b110 6
19
1>
1C
b110 G
#921260000000
0!
0*
09
0>
0C
#921270000000
1!
1*
b111 6
19
1>
1C
b111 G
#921280000000
0!
0*
09
0>
0C
#921290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#921300000000
0!
0*
09
0>
0C
#921310000000
1!
1*
b1 6
19
1>
1C
b1 G
#921320000000
0!
0*
09
0>
0C
#921330000000
1!
1*
b10 6
19
1>
1C
b10 G
#921340000000
0!
0*
09
0>
0C
#921350000000
1!
1*
b11 6
19
1>
1C
b11 G
#921360000000
0!
0*
09
0>
0C
#921370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#921380000000
0!
0*
09
0>
0C
#921390000000
1!
1*
b101 6
19
1>
1C
b101 G
#921400000000
0!
0*
09
0>
0C
#921410000000
1!
1*
b110 6
19
1>
1C
b110 G
#921420000000
0!
0*
09
0>
0C
#921430000000
1!
1*
b111 6
19
1>
1C
b111 G
#921440000000
0!
1"
0*
1+
09
1:
0>
0C
#921450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#921460000000
0!
0*
09
0>
0C
#921470000000
1!
1*
b1 6
19
1>
1C
b1 G
#921480000000
0!
0*
09
0>
0C
#921490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#921500000000
0!
0*
09
0>
0C
#921510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#921520000000
0!
0*
09
0>
0C
#921530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#921540000000
0!
0*
09
0>
0C
#921550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#921560000000
0!
0#
0*
0,
09
0>
0?
0C
#921570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#921580000000
0!
0*
09
0>
0C
#921590000000
1!
1*
19
1>
1C
#921600000000
0!
0*
09
0>
0C
#921610000000
1!
1*
19
1>
1C
#921620000000
0!
0*
09
0>
0C
#921630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#921640000000
0!
0*
09
0>
0C
#921650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#921660000000
0!
0*
09
0>
0C
#921670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#921680000000
0!
0*
09
0>
0C
#921690000000
1!
1*
b10 6
19
1>
1C
b10 G
#921700000000
0!
0*
09
0>
0C
#921710000000
1!
1*
b11 6
19
1>
1C
b11 G
#921720000000
0!
0*
09
0>
0C
#921730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#921740000000
0!
0*
09
0>
0C
#921750000000
1!
1*
b101 6
19
1>
1C
b101 G
#921760000000
0!
0*
09
0>
0C
#921770000000
1!
1*
b110 6
19
1>
1C
b110 G
#921780000000
0!
0*
09
0>
0C
#921790000000
1!
1*
b111 6
19
1>
1C
b111 G
#921800000000
0!
0*
09
0>
0C
#921810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#921820000000
0!
0*
09
0>
0C
#921830000000
1!
1*
b1 6
19
1>
1C
b1 G
#921840000000
0!
0*
09
0>
0C
#921850000000
1!
1*
b10 6
19
1>
1C
b10 G
#921860000000
0!
0*
09
0>
0C
#921870000000
1!
1*
b11 6
19
1>
1C
b11 G
#921880000000
0!
0*
09
0>
0C
#921890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#921900000000
0!
0*
09
0>
0C
#921910000000
1!
1*
b101 6
19
1>
1C
b101 G
#921920000000
0!
0*
09
0>
0C
#921930000000
1!
1*
b110 6
19
1>
1C
b110 G
#921940000000
0!
0*
09
0>
0C
#921950000000
1!
1*
b111 6
19
1>
1C
b111 G
#921960000000
0!
0*
09
0>
0C
#921970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#921980000000
0!
0*
09
0>
0C
#921990000000
1!
1*
b1 6
19
1>
1C
b1 G
#922000000000
0!
0*
09
0>
0C
#922010000000
1!
1*
b10 6
19
1>
1C
b10 G
#922020000000
0!
0*
09
0>
0C
#922030000000
1!
1*
b11 6
19
1>
1C
b11 G
#922040000000
0!
0*
09
0>
0C
#922050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#922060000000
0!
0*
09
0>
0C
#922070000000
1!
1*
b101 6
19
1>
1C
b101 G
#922080000000
0!
0*
09
0>
0C
#922090000000
1!
1*
b110 6
19
1>
1C
b110 G
#922100000000
0!
0*
09
0>
0C
#922110000000
1!
1*
b111 6
19
1>
1C
b111 G
#922120000000
0!
1"
0*
1+
09
1:
0>
0C
#922130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#922140000000
0!
0*
09
0>
0C
#922150000000
1!
1*
b1 6
19
1>
1C
b1 G
#922160000000
0!
0*
09
0>
0C
#922170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#922180000000
0!
0*
09
0>
0C
#922190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#922200000000
0!
0*
09
0>
0C
#922210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#922220000000
0!
0*
09
0>
0C
#922230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#922240000000
0!
0#
0*
0,
09
0>
0?
0C
#922250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#922260000000
0!
0*
09
0>
0C
#922270000000
1!
1*
19
1>
1C
#922280000000
0!
0*
09
0>
0C
#922290000000
1!
1*
19
1>
1C
#922300000000
0!
0*
09
0>
0C
#922310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#922320000000
0!
0*
09
0>
0C
#922330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#922340000000
0!
0*
09
0>
0C
#922350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#922360000000
0!
0*
09
0>
0C
#922370000000
1!
1*
b10 6
19
1>
1C
b10 G
#922380000000
0!
0*
09
0>
0C
#922390000000
1!
1*
b11 6
19
1>
1C
b11 G
#922400000000
0!
0*
09
0>
0C
#922410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#922420000000
0!
0*
09
0>
0C
#922430000000
1!
1*
b101 6
19
1>
1C
b101 G
#922440000000
0!
0*
09
0>
0C
#922450000000
1!
1*
b110 6
19
1>
1C
b110 G
#922460000000
0!
0*
09
0>
0C
#922470000000
1!
1*
b111 6
19
1>
1C
b111 G
#922480000000
0!
0*
09
0>
0C
#922490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#922500000000
0!
0*
09
0>
0C
#922510000000
1!
1*
b1 6
19
1>
1C
b1 G
#922520000000
0!
0*
09
0>
0C
#922530000000
1!
1*
b10 6
19
1>
1C
b10 G
#922540000000
0!
0*
09
0>
0C
#922550000000
1!
1*
b11 6
19
1>
1C
b11 G
#922560000000
0!
0*
09
0>
0C
#922570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#922580000000
0!
0*
09
0>
0C
#922590000000
1!
1*
b101 6
19
1>
1C
b101 G
#922600000000
0!
0*
09
0>
0C
#922610000000
1!
1*
b110 6
19
1>
1C
b110 G
#922620000000
0!
0*
09
0>
0C
#922630000000
1!
1*
b111 6
19
1>
1C
b111 G
#922640000000
0!
0*
09
0>
0C
#922650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#922660000000
0!
0*
09
0>
0C
#922670000000
1!
1*
b1 6
19
1>
1C
b1 G
#922680000000
0!
0*
09
0>
0C
#922690000000
1!
1*
b10 6
19
1>
1C
b10 G
#922700000000
0!
0*
09
0>
0C
#922710000000
1!
1*
b11 6
19
1>
1C
b11 G
#922720000000
0!
0*
09
0>
0C
#922730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#922740000000
0!
0*
09
0>
0C
#922750000000
1!
1*
b101 6
19
1>
1C
b101 G
#922760000000
0!
0*
09
0>
0C
#922770000000
1!
1*
b110 6
19
1>
1C
b110 G
#922780000000
0!
0*
09
0>
0C
#922790000000
1!
1*
b111 6
19
1>
1C
b111 G
#922800000000
0!
1"
0*
1+
09
1:
0>
0C
#922810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#922820000000
0!
0*
09
0>
0C
#922830000000
1!
1*
b1 6
19
1>
1C
b1 G
#922840000000
0!
0*
09
0>
0C
#922850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#922860000000
0!
0*
09
0>
0C
#922870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#922880000000
0!
0*
09
0>
0C
#922890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#922900000000
0!
0*
09
0>
0C
#922910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#922920000000
0!
0#
0*
0,
09
0>
0?
0C
#922930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#922940000000
0!
0*
09
0>
0C
#922950000000
1!
1*
19
1>
1C
#922960000000
0!
0*
09
0>
0C
#922970000000
1!
1*
19
1>
1C
#922980000000
0!
0*
09
0>
0C
#922990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#923000000000
0!
0*
09
0>
0C
#923010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#923020000000
0!
0*
09
0>
0C
#923030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#923040000000
0!
0*
09
0>
0C
#923050000000
1!
1*
b10 6
19
1>
1C
b10 G
#923060000000
0!
0*
09
0>
0C
#923070000000
1!
1*
b11 6
19
1>
1C
b11 G
#923080000000
0!
0*
09
0>
0C
#923090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#923100000000
0!
0*
09
0>
0C
#923110000000
1!
1*
b101 6
19
1>
1C
b101 G
#923120000000
0!
0*
09
0>
0C
#923130000000
1!
1*
b110 6
19
1>
1C
b110 G
#923140000000
0!
0*
09
0>
0C
#923150000000
1!
1*
b111 6
19
1>
1C
b111 G
#923160000000
0!
0*
09
0>
0C
#923170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#923180000000
0!
0*
09
0>
0C
#923190000000
1!
1*
b1 6
19
1>
1C
b1 G
#923200000000
0!
0*
09
0>
0C
#923210000000
1!
1*
b10 6
19
1>
1C
b10 G
#923220000000
0!
0*
09
0>
0C
#923230000000
1!
1*
b11 6
19
1>
1C
b11 G
#923240000000
0!
0*
09
0>
0C
#923250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#923260000000
0!
0*
09
0>
0C
#923270000000
1!
1*
b101 6
19
1>
1C
b101 G
#923280000000
0!
0*
09
0>
0C
#923290000000
1!
1*
b110 6
19
1>
1C
b110 G
#923300000000
0!
0*
09
0>
0C
#923310000000
1!
1*
b111 6
19
1>
1C
b111 G
#923320000000
0!
0*
09
0>
0C
#923330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#923340000000
0!
0*
09
0>
0C
#923350000000
1!
1*
b1 6
19
1>
1C
b1 G
#923360000000
0!
0*
09
0>
0C
#923370000000
1!
1*
b10 6
19
1>
1C
b10 G
#923380000000
0!
0*
09
0>
0C
#923390000000
1!
1*
b11 6
19
1>
1C
b11 G
#923400000000
0!
0*
09
0>
0C
#923410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#923420000000
0!
0*
09
0>
0C
#923430000000
1!
1*
b101 6
19
1>
1C
b101 G
#923440000000
0!
0*
09
0>
0C
#923450000000
1!
1*
b110 6
19
1>
1C
b110 G
#923460000000
0!
0*
09
0>
0C
#923470000000
1!
1*
b111 6
19
1>
1C
b111 G
#923480000000
0!
1"
0*
1+
09
1:
0>
0C
#923490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#923500000000
0!
0*
09
0>
0C
#923510000000
1!
1*
b1 6
19
1>
1C
b1 G
#923520000000
0!
0*
09
0>
0C
#923530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#923540000000
0!
0*
09
0>
0C
#923550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#923560000000
0!
0*
09
0>
0C
#923570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#923580000000
0!
0*
09
0>
0C
#923590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#923600000000
0!
0#
0*
0,
09
0>
0?
0C
#923610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#923620000000
0!
0*
09
0>
0C
#923630000000
1!
1*
19
1>
1C
#923640000000
0!
0*
09
0>
0C
#923650000000
1!
1*
19
1>
1C
#923660000000
0!
0*
09
0>
0C
#923670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#923680000000
0!
0*
09
0>
0C
#923690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#923700000000
0!
0*
09
0>
0C
#923710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#923720000000
0!
0*
09
0>
0C
#923730000000
1!
1*
b10 6
19
1>
1C
b10 G
#923740000000
0!
0*
09
0>
0C
#923750000000
1!
1*
b11 6
19
1>
1C
b11 G
#923760000000
0!
0*
09
0>
0C
#923770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#923780000000
0!
0*
09
0>
0C
#923790000000
1!
1*
b101 6
19
1>
1C
b101 G
#923800000000
0!
0*
09
0>
0C
#923810000000
1!
1*
b110 6
19
1>
1C
b110 G
#923820000000
0!
0*
09
0>
0C
#923830000000
1!
1*
b111 6
19
1>
1C
b111 G
#923840000000
0!
0*
09
0>
0C
#923850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#923860000000
0!
0*
09
0>
0C
#923870000000
1!
1*
b1 6
19
1>
1C
b1 G
#923880000000
0!
0*
09
0>
0C
#923890000000
1!
1*
b10 6
19
1>
1C
b10 G
#923900000000
0!
0*
09
0>
0C
#923910000000
1!
1*
b11 6
19
1>
1C
b11 G
#923920000000
0!
0*
09
0>
0C
#923930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#923940000000
0!
0*
09
0>
0C
#923950000000
1!
1*
b101 6
19
1>
1C
b101 G
#923960000000
0!
0*
09
0>
0C
#923970000000
1!
1*
b110 6
19
1>
1C
b110 G
#923980000000
0!
0*
09
0>
0C
#923990000000
1!
1*
b111 6
19
1>
1C
b111 G
#924000000000
0!
0*
09
0>
0C
#924010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#924020000000
0!
0*
09
0>
0C
#924030000000
1!
1*
b1 6
19
1>
1C
b1 G
#924040000000
0!
0*
09
0>
0C
#924050000000
1!
1*
b10 6
19
1>
1C
b10 G
#924060000000
0!
0*
09
0>
0C
#924070000000
1!
1*
b11 6
19
1>
1C
b11 G
#924080000000
0!
0*
09
0>
0C
#924090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#924100000000
0!
0*
09
0>
0C
#924110000000
1!
1*
b101 6
19
1>
1C
b101 G
#924120000000
0!
0*
09
0>
0C
#924130000000
1!
1*
b110 6
19
1>
1C
b110 G
#924140000000
0!
0*
09
0>
0C
#924150000000
1!
1*
b111 6
19
1>
1C
b111 G
#924160000000
0!
1"
0*
1+
09
1:
0>
0C
#924170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#924180000000
0!
0*
09
0>
0C
#924190000000
1!
1*
b1 6
19
1>
1C
b1 G
#924200000000
0!
0*
09
0>
0C
#924210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#924220000000
0!
0*
09
0>
0C
#924230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#924240000000
0!
0*
09
0>
0C
#924250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#924260000000
0!
0*
09
0>
0C
#924270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#924280000000
0!
0#
0*
0,
09
0>
0?
0C
#924290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#924300000000
0!
0*
09
0>
0C
#924310000000
1!
1*
19
1>
1C
#924320000000
0!
0*
09
0>
0C
#924330000000
1!
1*
19
1>
1C
#924340000000
0!
0*
09
0>
0C
#924350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#924360000000
0!
0*
09
0>
0C
#924370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#924380000000
0!
0*
09
0>
0C
#924390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#924400000000
0!
0*
09
0>
0C
#924410000000
1!
1*
b10 6
19
1>
1C
b10 G
#924420000000
0!
0*
09
0>
0C
#924430000000
1!
1*
b11 6
19
1>
1C
b11 G
#924440000000
0!
0*
09
0>
0C
#924450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#924460000000
0!
0*
09
0>
0C
#924470000000
1!
1*
b101 6
19
1>
1C
b101 G
#924480000000
0!
0*
09
0>
0C
#924490000000
1!
1*
b110 6
19
1>
1C
b110 G
#924500000000
0!
0*
09
0>
0C
#924510000000
1!
1*
b111 6
19
1>
1C
b111 G
#924520000000
0!
0*
09
0>
0C
#924530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#924540000000
0!
0*
09
0>
0C
#924550000000
1!
1*
b1 6
19
1>
1C
b1 G
#924560000000
0!
0*
09
0>
0C
#924570000000
1!
1*
b10 6
19
1>
1C
b10 G
#924580000000
0!
0*
09
0>
0C
#924590000000
1!
1*
b11 6
19
1>
1C
b11 G
#924600000000
0!
0*
09
0>
0C
#924610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#924620000000
0!
0*
09
0>
0C
#924630000000
1!
1*
b101 6
19
1>
1C
b101 G
#924640000000
0!
0*
09
0>
0C
#924650000000
1!
1*
b110 6
19
1>
1C
b110 G
#924660000000
0!
0*
09
0>
0C
#924670000000
1!
1*
b111 6
19
1>
1C
b111 G
#924680000000
0!
0*
09
0>
0C
#924690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#924700000000
0!
0*
09
0>
0C
#924710000000
1!
1*
b1 6
19
1>
1C
b1 G
#924720000000
0!
0*
09
0>
0C
#924730000000
1!
1*
b10 6
19
1>
1C
b10 G
#924740000000
0!
0*
09
0>
0C
#924750000000
1!
1*
b11 6
19
1>
1C
b11 G
#924760000000
0!
0*
09
0>
0C
#924770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#924780000000
0!
0*
09
0>
0C
#924790000000
1!
1*
b101 6
19
1>
1C
b101 G
#924800000000
0!
0*
09
0>
0C
#924810000000
1!
1*
b110 6
19
1>
1C
b110 G
#924820000000
0!
0*
09
0>
0C
#924830000000
1!
1*
b111 6
19
1>
1C
b111 G
#924840000000
0!
1"
0*
1+
09
1:
0>
0C
#924850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#924860000000
0!
0*
09
0>
0C
#924870000000
1!
1*
b1 6
19
1>
1C
b1 G
#924880000000
0!
0*
09
0>
0C
#924890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#924900000000
0!
0*
09
0>
0C
#924910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#924920000000
0!
0*
09
0>
0C
#924930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#924940000000
0!
0*
09
0>
0C
#924950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#924960000000
0!
0#
0*
0,
09
0>
0?
0C
#924970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#924980000000
0!
0*
09
0>
0C
#924990000000
1!
1*
19
1>
1C
#925000000000
0!
0*
09
0>
0C
#925010000000
1!
1*
19
1>
1C
#925020000000
0!
0*
09
0>
0C
#925030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#925040000000
0!
0*
09
0>
0C
#925050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#925060000000
0!
0*
09
0>
0C
#925070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#925080000000
0!
0*
09
0>
0C
#925090000000
1!
1*
b10 6
19
1>
1C
b10 G
#925100000000
0!
0*
09
0>
0C
#925110000000
1!
1*
b11 6
19
1>
1C
b11 G
#925120000000
0!
0*
09
0>
0C
#925130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#925140000000
0!
0*
09
0>
0C
#925150000000
1!
1*
b101 6
19
1>
1C
b101 G
#925160000000
0!
0*
09
0>
0C
#925170000000
1!
1*
b110 6
19
1>
1C
b110 G
#925180000000
0!
0*
09
0>
0C
#925190000000
1!
1*
b111 6
19
1>
1C
b111 G
#925200000000
0!
0*
09
0>
0C
#925210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#925220000000
0!
0*
09
0>
0C
#925230000000
1!
1*
b1 6
19
1>
1C
b1 G
#925240000000
0!
0*
09
0>
0C
#925250000000
1!
1*
b10 6
19
1>
1C
b10 G
#925260000000
0!
0*
09
0>
0C
#925270000000
1!
1*
b11 6
19
1>
1C
b11 G
#925280000000
0!
0*
09
0>
0C
#925290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#925300000000
0!
0*
09
0>
0C
#925310000000
1!
1*
b101 6
19
1>
1C
b101 G
#925320000000
0!
0*
09
0>
0C
#925330000000
1!
1*
b110 6
19
1>
1C
b110 G
#925340000000
0!
0*
09
0>
0C
#925350000000
1!
1*
b111 6
19
1>
1C
b111 G
#925360000000
0!
0*
09
0>
0C
#925370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#925380000000
0!
0*
09
0>
0C
#925390000000
1!
1*
b1 6
19
1>
1C
b1 G
#925400000000
0!
0*
09
0>
0C
#925410000000
1!
1*
b10 6
19
1>
1C
b10 G
#925420000000
0!
0*
09
0>
0C
#925430000000
1!
1*
b11 6
19
1>
1C
b11 G
#925440000000
0!
0*
09
0>
0C
#925450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#925460000000
0!
0*
09
0>
0C
#925470000000
1!
1*
b101 6
19
1>
1C
b101 G
#925480000000
0!
0*
09
0>
0C
#925490000000
1!
1*
b110 6
19
1>
1C
b110 G
#925500000000
0!
0*
09
0>
0C
#925510000000
1!
1*
b111 6
19
1>
1C
b111 G
#925520000000
0!
1"
0*
1+
09
1:
0>
0C
#925530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#925540000000
0!
0*
09
0>
0C
#925550000000
1!
1*
b1 6
19
1>
1C
b1 G
#925560000000
0!
0*
09
0>
0C
#925570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#925580000000
0!
0*
09
0>
0C
#925590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#925600000000
0!
0*
09
0>
0C
#925610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#925620000000
0!
0*
09
0>
0C
#925630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#925640000000
0!
0#
0*
0,
09
0>
0?
0C
#925650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#925660000000
0!
0*
09
0>
0C
#925670000000
1!
1*
19
1>
1C
#925680000000
0!
0*
09
0>
0C
#925690000000
1!
1*
19
1>
1C
#925700000000
0!
0*
09
0>
0C
#925710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#925720000000
0!
0*
09
0>
0C
#925730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#925740000000
0!
0*
09
0>
0C
#925750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#925760000000
0!
0*
09
0>
0C
#925770000000
1!
1*
b10 6
19
1>
1C
b10 G
#925780000000
0!
0*
09
0>
0C
#925790000000
1!
1*
b11 6
19
1>
1C
b11 G
#925800000000
0!
0*
09
0>
0C
#925810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#925820000000
0!
0*
09
0>
0C
#925830000000
1!
1*
b101 6
19
1>
1C
b101 G
#925840000000
0!
0*
09
0>
0C
#925850000000
1!
1*
b110 6
19
1>
1C
b110 G
#925860000000
0!
0*
09
0>
0C
#925870000000
1!
1*
b111 6
19
1>
1C
b111 G
#925880000000
0!
0*
09
0>
0C
#925890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#925900000000
0!
0*
09
0>
0C
#925910000000
1!
1*
b1 6
19
1>
1C
b1 G
#925920000000
0!
0*
09
0>
0C
#925930000000
1!
1*
b10 6
19
1>
1C
b10 G
#925940000000
0!
0*
09
0>
0C
#925950000000
1!
1*
b11 6
19
1>
1C
b11 G
#925960000000
0!
0*
09
0>
0C
#925970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#925980000000
0!
0*
09
0>
0C
#925990000000
1!
1*
b101 6
19
1>
1C
b101 G
#926000000000
0!
0*
09
0>
0C
#926010000000
1!
1*
b110 6
19
1>
1C
b110 G
#926020000000
0!
0*
09
0>
0C
#926030000000
1!
1*
b111 6
19
1>
1C
b111 G
#926040000000
0!
0*
09
0>
0C
#926050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#926060000000
0!
0*
09
0>
0C
#926070000000
1!
1*
b1 6
19
1>
1C
b1 G
#926080000000
0!
0*
09
0>
0C
#926090000000
1!
1*
b10 6
19
1>
1C
b10 G
#926100000000
0!
0*
09
0>
0C
#926110000000
1!
1*
b11 6
19
1>
1C
b11 G
#926120000000
0!
0*
09
0>
0C
#926130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#926140000000
0!
0*
09
0>
0C
#926150000000
1!
1*
b101 6
19
1>
1C
b101 G
#926160000000
0!
0*
09
0>
0C
#926170000000
1!
1*
b110 6
19
1>
1C
b110 G
#926180000000
0!
0*
09
0>
0C
#926190000000
1!
1*
b111 6
19
1>
1C
b111 G
#926200000000
0!
1"
0*
1+
09
1:
0>
0C
#926210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#926220000000
0!
0*
09
0>
0C
#926230000000
1!
1*
b1 6
19
1>
1C
b1 G
#926240000000
0!
0*
09
0>
0C
#926250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#926260000000
0!
0*
09
0>
0C
#926270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#926280000000
0!
0*
09
0>
0C
#926290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#926300000000
0!
0*
09
0>
0C
#926310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#926320000000
0!
0#
0*
0,
09
0>
0?
0C
#926330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#926340000000
0!
0*
09
0>
0C
#926350000000
1!
1*
19
1>
1C
#926360000000
0!
0*
09
0>
0C
#926370000000
1!
1*
19
1>
1C
#926380000000
0!
0*
09
0>
0C
#926390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#926400000000
0!
0*
09
0>
0C
#926410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#926420000000
0!
0*
09
0>
0C
#926430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#926440000000
0!
0*
09
0>
0C
#926450000000
1!
1*
b10 6
19
1>
1C
b10 G
#926460000000
0!
0*
09
0>
0C
#926470000000
1!
1*
b11 6
19
1>
1C
b11 G
#926480000000
0!
0*
09
0>
0C
#926490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#926500000000
0!
0*
09
0>
0C
#926510000000
1!
1*
b101 6
19
1>
1C
b101 G
#926520000000
0!
0*
09
0>
0C
#926530000000
1!
1*
b110 6
19
1>
1C
b110 G
#926540000000
0!
0*
09
0>
0C
#926550000000
1!
1*
b111 6
19
1>
1C
b111 G
#926560000000
0!
0*
09
0>
0C
#926570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#926580000000
0!
0*
09
0>
0C
#926590000000
1!
1*
b1 6
19
1>
1C
b1 G
#926600000000
0!
0*
09
0>
0C
#926610000000
1!
1*
b10 6
19
1>
1C
b10 G
#926620000000
0!
0*
09
0>
0C
#926630000000
1!
1*
b11 6
19
1>
1C
b11 G
#926640000000
0!
0*
09
0>
0C
#926650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#926660000000
0!
0*
09
0>
0C
#926670000000
1!
1*
b101 6
19
1>
1C
b101 G
#926680000000
0!
0*
09
0>
0C
#926690000000
1!
1*
b110 6
19
1>
1C
b110 G
#926700000000
0!
0*
09
0>
0C
#926710000000
1!
1*
b111 6
19
1>
1C
b111 G
#926720000000
0!
0*
09
0>
0C
#926730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#926740000000
0!
0*
09
0>
0C
#926750000000
1!
1*
b1 6
19
1>
1C
b1 G
#926760000000
0!
0*
09
0>
0C
#926770000000
1!
1*
b10 6
19
1>
1C
b10 G
#926780000000
0!
0*
09
0>
0C
#926790000000
1!
1*
b11 6
19
1>
1C
b11 G
#926800000000
0!
0*
09
0>
0C
#926810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#926820000000
0!
0*
09
0>
0C
#926830000000
1!
1*
b101 6
19
1>
1C
b101 G
#926840000000
0!
0*
09
0>
0C
#926850000000
1!
1*
b110 6
19
1>
1C
b110 G
#926860000000
0!
0*
09
0>
0C
#926870000000
1!
1*
b111 6
19
1>
1C
b111 G
#926880000000
0!
1"
0*
1+
09
1:
0>
0C
#926890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#926900000000
0!
0*
09
0>
0C
#926910000000
1!
1*
b1 6
19
1>
1C
b1 G
#926920000000
0!
0*
09
0>
0C
#926930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#926940000000
0!
0*
09
0>
0C
#926950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#926960000000
0!
0*
09
0>
0C
#926970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#926980000000
0!
0*
09
0>
0C
#926990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#927000000000
0!
0#
0*
0,
09
0>
0?
0C
#927010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#927020000000
0!
0*
09
0>
0C
#927030000000
1!
1*
19
1>
1C
#927040000000
0!
0*
09
0>
0C
#927050000000
1!
1*
19
1>
1C
#927060000000
0!
0*
09
0>
0C
#927070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#927080000000
0!
0*
09
0>
0C
#927090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#927100000000
0!
0*
09
0>
0C
#927110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#927120000000
0!
0*
09
0>
0C
#927130000000
1!
1*
b10 6
19
1>
1C
b10 G
#927140000000
0!
0*
09
0>
0C
#927150000000
1!
1*
b11 6
19
1>
1C
b11 G
#927160000000
0!
0*
09
0>
0C
#927170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#927180000000
0!
0*
09
0>
0C
#927190000000
1!
1*
b101 6
19
1>
1C
b101 G
#927200000000
0!
0*
09
0>
0C
#927210000000
1!
1*
b110 6
19
1>
1C
b110 G
#927220000000
0!
0*
09
0>
0C
#927230000000
1!
1*
b111 6
19
1>
1C
b111 G
#927240000000
0!
0*
09
0>
0C
#927250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#927260000000
0!
0*
09
0>
0C
#927270000000
1!
1*
b1 6
19
1>
1C
b1 G
#927280000000
0!
0*
09
0>
0C
#927290000000
1!
1*
b10 6
19
1>
1C
b10 G
#927300000000
0!
0*
09
0>
0C
#927310000000
1!
1*
b11 6
19
1>
1C
b11 G
#927320000000
0!
0*
09
0>
0C
#927330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#927340000000
0!
0*
09
0>
0C
#927350000000
1!
1*
b101 6
19
1>
1C
b101 G
#927360000000
0!
0*
09
0>
0C
#927370000000
1!
1*
b110 6
19
1>
1C
b110 G
#927380000000
0!
0*
09
0>
0C
#927390000000
1!
1*
b111 6
19
1>
1C
b111 G
#927400000000
0!
0*
09
0>
0C
#927410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#927420000000
0!
0*
09
0>
0C
#927430000000
1!
1*
b1 6
19
1>
1C
b1 G
#927440000000
0!
0*
09
0>
0C
#927450000000
1!
1*
b10 6
19
1>
1C
b10 G
#927460000000
0!
0*
09
0>
0C
#927470000000
1!
1*
b11 6
19
1>
1C
b11 G
#927480000000
0!
0*
09
0>
0C
#927490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#927500000000
0!
0*
09
0>
0C
#927510000000
1!
1*
b101 6
19
1>
1C
b101 G
#927520000000
0!
0*
09
0>
0C
#927530000000
1!
1*
b110 6
19
1>
1C
b110 G
#927540000000
0!
0*
09
0>
0C
#927550000000
1!
1*
b111 6
19
1>
1C
b111 G
#927560000000
0!
1"
0*
1+
09
1:
0>
0C
#927570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#927580000000
0!
0*
09
0>
0C
#927590000000
1!
1*
b1 6
19
1>
1C
b1 G
#927600000000
0!
0*
09
0>
0C
#927610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#927620000000
0!
0*
09
0>
0C
#927630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#927640000000
0!
0*
09
0>
0C
#927650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#927660000000
0!
0*
09
0>
0C
#927670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#927680000000
0!
0#
0*
0,
09
0>
0?
0C
#927690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#927700000000
0!
0*
09
0>
0C
#927710000000
1!
1*
19
1>
1C
#927720000000
0!
0*
09
0>
0C
#927730000000
1!
1*
19
1>
1C
#927740000000
0!
0*
09
0>
0C
#927750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#927760000000
0!
0*
09
0>
0C
#927770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#927780000000
0!
0*
09
0>
0C
#927790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#927800000000
0!
0*
09
0>
0C
#927810000000
1!
1*
b10 6
19
1>
1C
b10 G
#927820000000
0!
0*
09
0>
0C
#927830000000
1!
1*
b11 6
19
1>
1C
b11 G
#927840000000
0!
0*
09
0>
0C
#927850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#927860000000
0!
0*
09
0>
0C
#927870000000
1!
1*
b101 6
19
1>
1C
b101 G
#927880000000
0!
0*
09
0>
0C
#927890000000
1!
1*
b110 6
19
1>
1C
b110 G
#927900000000
0!
0*
09
0>
0C
#927910000000
1!
1*
b111 6
19
1>
1C
b111 G
#927920000000
0!
0*
09
0>
0C
#927930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#927940000000
0!
0*
09
0>
0C
#927950000000
1!
1*
b1 6
19
1>
1C
b1 G
#927960000000
0!
0*
09
0>
0C
#927970000000
1!
1*
b10 6
19
1>
1C
b10 G
#927980000000
0!
0*
09
0>
0C
#927990000000
1!
1*
b11 6
19
1>
1C
b11 G
#928000000000
0!
0*
09
0>
0C
#928010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#928020000000
0!
0*
09
0>
0C
#928030000000
1!
1*
b101 6
19
1>
1C
b101 G
#928040000000
0!
0*
09
0>
0C
#928050000000
1!
1*
b110 6
19
1>
1C
b110 G
#928060000000
0!
0*
09
0>
0C
#928070000000
1!
1*
b111 6
19
1>
1C
b111 G
#928080000000
0!
0*
09
0>
0C
#928090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#928100000000
0!
0*
09
0>
0C
#928110000000
1!
1*
b1 6
19
1>
1C
b1 G
#928120000000
0!
0*
09
0>
0C
#928130000000
1!
1*
b10 6
19
1>
1C
b10 G
#928140000000
0!
0*
09
0>
0C
#928150000000
1!
1*
b11 6
19
1>
1C
b11 G
#928160000000
0!
0*
09
0>
0C
#928170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#928180000000
0!
0*
09
0>
0C
#928190000000
1!
1*
b101 6
19
1>
1C
b101 G
#928200000000
0!
0*
09
0>
0C
#928210000000
1!
1*
b110 6
19
1>
1C
b110 G
#928220000000
0!
0*
09
0>
0C
#928230000000
1!
1*
b111 6
19
1>
1C
b111 G
#928240000000
0!
1"
0*
1+
09
1:
0>
0C
#928250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#928260000000
0!
0*
09
0>
0C
#928270000000
1!
1*
b1 6
19
1>
1C
b1 G
#928280000000
0!
0*
09
0>
0C
#928290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#928300000000
0!
0*
09
0>
0C
#928310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#928320000000
0!
0*
09
0>
0C
#928330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#928340000000
0!
0*
09
0>
0C
#928350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#928360000000
0!
0#
0*
0,
09
0>
0?
0C
#928370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#928380000000
0!
0*
09
0>
0C
#928390000000
1!
1*
19
1>
1C
#928400000000
0!
0*
09
0>
0C
#928410000000
1!
1*
19
1>
1C
#928420000000
0!
0*
09
0>
0C
#928430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#928440000000
0!
0*
09
0>
0C
#928450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#928460000000
0!
0*
09
0>
0C
#928470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#928480000000
0!
0*
09
0>
0C
#928490000000
1!
1*
b10 6
19
1>
1C
b10 G
#928500000000
0!
0*
09
0>
0C
#928510000000
1!
1*
b11 6
19
1>
1C
b11 G
#928520000000
0!
0*
09
0>
0C
#928530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#928540000000
0!
0*
09
0>
0C
#928550000000
1!
1*
b101 6
19
1>
1C
b101 G
#928560000000
0!
0*
09
0>
0C
#928570000000
1!
1*
b110 6
19
1>
1C
b110 G
#928580000000
0!
0*
09
0>
0C
#928590000000
1!
1*
b111 6
19
1>
1C
b111 G
#928600000000
0!
0*
09
0>
0C
#928610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#928620000000
0!
0*
09
0>
0C
#928630000000
1!
1*
b1 6
19
1>
1C
b1 G
#928640000000
0!
0*
09
0>
0C
#928650000000
1!
1*
b10 6
19
1>
1C
b10 G
#928660000000
0!
0*
09
0>
0C
#928670000000
1!
1*
b11 6
19
1>
1C
b11 G
#928680000000
0!
0*
09
0>
0C
#928690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#928700000000
0!
0*
09
0>
0C
#928710000000
1!
1*
b101 6
19
1>
1C
b101 G
#928720000000
0!
0*
09
0>
0C
#928730000000
1!
1*
b110 6
19
1>
1C
b110 G
#928740000000
0!
0*
09
0>
0C
#928750000000
1!
1*
b111 6
19
1>
1C
b111 G
#928760000000
0!
0*
09
0>
0C
#928770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#928780000000
0!
0*
09
0>
0C
#928790000000
1!
1*
b1 6
19
1>
1C
b1 G
#928800000000
0!
0*
09
0>
0C
#928810000000
1!
1*
b10 6
19
1>
1C
b10 G
#928820000000
0!
0*
09
0>
0C
#928830000000
1!
1*
b11 6
19
1>
1C
b11 G
#928840000000
0!
0*
09
0>
0C
#928850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#928860000000
0!
0*
09
0>
0C
#928870000000
1!
1*
b101 6
19
1>
1C
b101 G
#928880000000
0!
0*
09
0>
0C
#928890000000
1!
1*
b110 6
19
1>
1C
b110 G
#928900000000
0!
0*
09
0>
0C
#928910000000
1!
1*
b111 6
19
1>
1C
b111 G
#928920000000
0!
1"
0*
1+
09
1:
0>
0C
#928930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#928940000000
0!
0*
09
0>
0C
#928950000000
1!
1*
b1 6
19
1>
1C
b1 G
#928960000000
0!
0*
09
0>
0C
#928970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#928980000000
0!
0*
09
0>
0C
#928990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#929000000000
0!
0*
09
0>
0C
#929010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#929020000000
0!
0*
09
0>
0C
#929030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#929040000000
0!
0#
0*
0,
09
0>
0?
0C
#929050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#929060000000
0!
0*
09
0>
0C
#929070000000
1!
1*
19
1>
1C
#929080000000
0!
0*
09
0>
0C
#929090000000
1!
1*
19
1>
1C
#929100000000
0!
0*
09
0>
0C
#929110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#929120000000
0!
0*
09
0>
0C
#929130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#929140000000
0!
0*
09
0>
0C
#929150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#929160000000
0!
0*
09
0>
0C
#929170000000
1!
1*
b10 6
19
1>
1C
b10 G
#929180000000
0!
0*
09
0>
0C
#929190000000
1!
1*
b11 6
19
1>
1C
b11 G
#929200000000
0!
0*
09
0>
0C
#929210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#929220000000
0!
0*
09
0>
0C
#929230000000
1!
1*
b101 6
19
1>
1C
b101 G
#929240000000
0!
0*
09
0>
0C
#929250000000
1!
1*
b110 6
19
1>
1C
b110 G
#929260000000
0!
0*
09
0>
0C
#929270000000
1!
1*
b111 6
19
1>
1C
b111 G
#929280000000
0!
0*
09
0>
0C
#929290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#929300000000
0!
0*
09
0>
0C
#929310000000
1!
1*
b1 6
19
1>
1C
b1 G
#929320000000
0!
0*
09
0>
0C
#929330000000
1!
1*
b10 6
19
1>
1C
b10 G
#929340000000
0!
0*
09
0>
0C
#929350000000
1!
1*
b11 6
19
1>
1C
b11 G
#929360000000
0!
0*
09
0>
0C
#929370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#929380000000
0!
0*
09
0>
0C
#929390000000
1!
1*
b101 6
19
1>
1C
b101 G
#929400000000
0!
0*
09
0>
0C
#929410000000
1!
1*
b110 6
19
1>
1C
b110 G
#929420000000
0!
0*
09
0>
0C
#929430000000
1!
1*
b111 6
19
1>
1C
b111 G
#929440000000
0!
0*
09
0>
0C
#929450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#929460000000
0!
0*
09
0>
0C
#929470000000
1!
1*
b1 6
19
1>
1C
b1 G
#929480000000
0!
0*
09
0>
0C
#929490000000
1!
1*
b10 6
19
1>
1C
b10 G
#929500000000
0!
0*
09
0>
0C
#929510000000
1!
1*
b11 6
19
1>
1C
b11 G
#929520000000
0!
0*
09
0>
0C
#929530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#929540000000
0!
0*
09
0>
0C
#929550000000
1!
1*
b101 6
19
1>
1C
b101 G
#929560000000
0!
0*
09
0>
0C
#929570000000
1!
1*
b110 6
19
1>
1C
b110 G
#929580000000
0!
0*
09
0>
0C
#929590000000
1!
1*
b111 6
19
1>
1C
b111 G
#929600000000
0!
1"
0*
1+
09
1:
0>
0C
#929610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#929620000000
0!
0*
09
0>
0C
#929630000000
1!
1*
b1 6
19
1>
1C
b1 G
#929640000000
0!
0*
09
0>
0C
#929650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#929660000000
0!
0*
09
0>
0C
#929670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#929680000000
0!
0*
09
0>
0C
#929690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#929700000000
0!
0*
09
0>
0C
#929710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#929720000000
0!
0#
0*
0,
09
0>
0?
0C
#929730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#929740000000
0!
0*
09
0>
0C
#929750000000
1!
1*
19
1>
1C
#929760000000
0!
0*
09
0>
0C
#929770000000
1!
1*
19
1>
1C
#929780000000
0!
0*
09
0>
0C
#929790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#929800000000
0!
0*
09
0>
0C
#929810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#929820000000
0!
0*
09
0>
0C
#929830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#929840000000
0!
0*
09
0>
0C
#929850000000
1!
1*
b10 6
19
1>
1C
b10 G
#929860000000
0!
0*
09
0>
0C
#929870000000
1!
1*
b11 6
19
1>
1C
b11 G
#929880000000
0!
0*
09
0>
0C
#929890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#929900000000
0!
0*
09
0>
0C
#929910000000
1!
1*
b101 6
19
1>
1C
b101 G
#929920000000
0!
0*
09
0>
0C
#929930000000
1!
1*
b110 6
19
1>
1C
b110 G
#929940000000
0!
0*
09
0>
0C
#929950000000
1!
1*
b111 6
19
1>
1C
b111 G
#929960000000
0!
0*
09
0>
0C
#929970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#929980000000
0!
0*
09
0>
0C
#929990000000
1!
1*
b1 6
19
1>
1C
b1 G
#930000000000
0!
0*
09
0>
0C
#930010000000
1!
1*
b10 6
19
1>
1C
b10 G
#930020000000
0!
0*
09
0>
0C
#930030000000
1!
1*
b11 6
19
1>
1C
b11 G
#930040000000
0!
0*
09
0>
0C
#930050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#930060000000
0!
0*
09
0>
0C
#930070000000
1!
1*
b101 6
19
1>
1C
b101 G
#930080000000
0!
0*
09
0>
0C
#930090000000
1!
1*
b110 6
19
1>
1C
b110 G
#930100000000
0!
0*
09
0>
0C
#930110000000
1!
1*
b111 6
19
1>
1C
b111 G
#930120000000
0!
0*
09
0>
0C
#930130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#930140000000
0!
0*
09
0>
0C
#930150000000
1!
1*
b1 6
19
1>
1C
b1 G
#930160000000
0!
0*
09
0>
0C
#930170000000
1!
1*
b10 6
19
1>
1C
b10 G
#930180000000
0!
0*
09
0>
0C
#930190000000
1!
1*
b11 6
19
1>
1C
b11 G
#930200000000
0!
0*
09
0>
0C
#930210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#930220000000
0!
0*
09
0>
0C
#930230000000
1!
1*
b101 6
19
1>
1C
b101 G
#930240000000
0!
0*
09
0>
0C
#930250000000
1!
1*
b110 6
19
1>
1C
b110 G
#930260000000
0!
0*
09
0>
0C
#930270000000
1!
1*
b111 6
19
1>
1C
b111 G
#930280000000
0!
1"
0*
1+
09
1:
0>
0C
#930290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#930300000000
0!
0*
09
0>
0C
#930310000000
1!
1*
b1 6
19
1>
1C
b1 G
#930320000000
0!
0*
09
0>
0C
#930330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#930340000000
0!
0*
09
0>
0C
#930350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#930360000000
0!
0*
09
0>
0C
#930370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#930380000000
0!
0*
09
0>
0C
#930390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#930400000000
0!
0#
0*
0,
09
0>
0?
0C
#930410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#930420000000
0!
0*
09
0>
0C
#930430000000
1!
1*
19
1>
1C
#930440000000
0!
0*
09
0>
0C
#930450000000
1!
1*
19
1>
1C
#930460000000
0!
0*
09
0>
0C
#930470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#930480000000
0!
0*
09
0>
0C
#930490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#930500000000
0!
0*
09
0>
0C
#930510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#930520000000
0!
0*
09
0>
0C
#930530000000
1!
1*
b10 6
19
1>
1C
b10 G
#930540000000
0!
0*
09
0>
0C
#930550000000
1!
1*
b11 6
19
1>
1C
b11 G
#930560000000
0!
0*
09
0>
0C
#930570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#930580000000
0!
0*
09
0>
0C
#930590000000
1!
1*
b101 6
19
1>
1C
b101 G
#930600000000
0!
0*
09
0>
0C
#930610000000
1!
1*
b110 6
19
1>
1C
b110 G
#930620000000
0!
0*
09
0>
0C
#930630000000
1!
1*
b111 6
19
1>
1C
b111 G
#930640000000
0!
0*
09
0>
0C
#930650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#930660000000
0!
0*
09
0>
0C
#930670000000
1!
1*
b1 6
19
1>
1C
b1 G
#930680000000
0!
0*
09
0>
0C
#930690000000
1!
1*
b10 6
19
1>
1C
b10 G
#930700000000
0!
0*
09
0>
0C
#930710000000
1!
1*
b11 6
19
1>
1C
b11 G
#930720000000
0!
0*
09
0>
0C
#930730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#930740000000
0!
0*
09
0>
0C
#930750000000
1!
1*
b101 6
19
1>
1C
b101 G
#930760000000
0!
0*
09
0>
0C
#930770000000
1!
1*
b110 6
19
1>
1C
b110 G
#930780000000
0!
0*
09
0>
0C
#930790000000
1!
1*
b111 6
19
1>
1C
b111 G
#930800000000
0!
0*
09
0>
0C
#930810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#930820000000
0!
0*
09
0>
0C
#930830000000
1!
1*
b1 6
19
1>
1C
b1 G
#930840000000
0!
0*
09
0>
0C
#930850000000
1!
1*
b10 6
19
1>
1C
b10 G
#930860000000
0!
0*
09
0>
0C
#930870000000
1!
1*
b11 6
19
1>
1C
b11 G
#930880000000
0!
0*
09
0>
0C
#930890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#930900000000
0!
0*
09
0>
0C
#930910000000
1!
1*
b101 6
19
1>
1C
b101 G
#930920000000
0!
0*
09
0>
0C
#930930000000
1!
1*
b110 6
19
1>
1C
b110 G
#930940000000
0!
0*
09
0>
0C
#930950000000
1!
1*
b111 6
19
1>
1C
b111 G
#930960000000
0!
1"
0*
1+
09
1:
0>
0C
#930970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#930980000000
0!
0*
09
0>
0C
#930990000000
1!
1*
b1 6
19
1>
1C
b1 G
#931000000000
0!
0*
09
0>
0C
#931010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#931020000000
0!
0*
09
0>
0C
#931030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#931040000000
0!
0*
09
0>
0C
#931050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#931060000000
0!
0*
09
0>
0C
#931070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#931080000000
0!
0#
0*
0,
09
0>
0?
0C
#931090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#931100000000
0!
0*
09
0>
0C
#931110000000
1!
1*
19
1>
1C
#931120000000
0!
0*
09
0>
0C
#931130000000
1!
1*
19
1>
1C
#931140000000
0!
0*
09
0>
0C
#931150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#931160000000
0!
0*
09
0>
0C
#931170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#931180000000
0!
0*
09
0>
0C
#931190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#931200000000
0!
0*
09
0>
0C
#931210000000
1!
1*
b10 6
19
1>
1C
b10 G
#931220000000
0!
0*
09
0>
0C
#931230000000
1!
1*
b11 6
19
1>
1C
b11 G
#931240000000
0!
0*
09
0>
0C
#931250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#931260000000
0!
0*
09
0>
0C
#931270000000
1!
1*
b101 6
19
1>
1C
b101 G
#931280000000
0!
0*
09
0>
0C
#931290000000
1!
1*
b110 6
19
1>
1C
b110 G
#931300000000
0!
0*
09
0>
0C
#931310000000
1!
1*
b111 6
19
1>
1C
b111 G
#931320000000
0!
0*
09
0>
0C
#931330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#931340000000
0!
0*
09
0>
0C
#931350000000
1!
1*
b1 6
19
1>
1C
b1 G
#931360000000
0!
0*
09
0>
0C
#931370000000
1!
1*
b10 6
19
1>
1C
b10 G
#931380000000
0!
0*
09
0>
0C
#931390000000
1!
1*
b11 6
19
1>
1C
b11 G
#931400000000
0!
0*
09
0>
0C
#931410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#931420000000
0!
0*
09
0>
0C
#931430000000
1!
1*
b101 6
19
1>
1C
b101 G
#931440000000
0!
0*
09
0>
0C
#931450000000
1!
1*
b110 6
19
1>
1C
b110 G
#931460000000
0!
0*
09
0>
0C
#931470000000
1!
1*
b111 6
19
1>
1C
b111 G
#931480000000
0!
0*
09
0>
0C
#931490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#931500000000
0!
0*
09
0>
0C
#931510000000
1!
1*
b1 6
19
1>
1C
b1 G
#931520000000
0!
0*
09
0>
0C
#931530000000
1!
1*
b10 6
19
1>
1C
b10 G
#931540000000
0!
0*
09
0>
0C
#931550000000
1!
1*
b11 6
19
1>
1C
b11 G
#931560000000
0!
0*
09
0>
0C
#931570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#931580000000
0!
0*
09
0>
0C
#931590000000
1!
1*
b101 6
19
1>
1C
b101 G
#931600000000
0!
0*
09
0>
0C
#931610000000
1!
1*
b110 6
19
1>
1C
b110 G
#931620000000
0!
0*
09
0>
0C
#931630000000
1!
1*
b111 6
19
1>
1C
b111 G
#931640000000
0!
1"
0*
1+
09
1:
0>
0C
#931650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#931660000000
0!
0*
09
0>
0C
#931670000000
1!
1*
b1 6
19
1>
1C
b1 G
#931680000000
0!
0*
09
0>
0C
#931690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#931700000000
0!
0*
09
0>
0C
#931710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#931720000000
0!
0*
09
0>
0C
#931730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#931740000000
0!
0*
09
0>
0C
#931750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#931760000000
0!
0#
0*
0,
09
0>
0?
0C
#931770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#931780000000
0!
0*
09
0>
0C
#931790000000
1!
1*
19
1>
1C
#931800000000
0!
0*
09
0>
0C
#931810000000
1!
1*
19
1>
1C
#931820000000
0!
0*
09
0>
0C
#931830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#931840000000
0!
0*
09
0>
0C
#931850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#931860000000
0!
0*
09
0>
0C
#931870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#931880000000
0!
0*
09
0>
0C
#931890000000
1!
1*
b10 6
19
1>
1C
b10 G
#931900000000
0!
0*
09
0>
0C
#931910000000
1!
1*
b11 6
19
1>
1C
b11 G
#931920000000
0!
0*
09
0>
0C
#931930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#931940000000
0!
0*
09
0>
0C
#931950000000
1!
1*
b101 6
19
1>
1C
b101 G
#931960000000
0!
0*
09
0>
0C
#931970000000
1!
1*
b110 6
19
1>
1C
b110 G
#931980000000
0!
0*
09
0>
0C
#931990000000
1!
1*
b111 6
19
1>
1C
b111 G
#932000000000
0!
0*
09
0>
0C
#932010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#932020000000
0!
0*
09
0>
0C
#932030000000
1!
1*
b1 6
19
1>
1C
b1 G
#932040000000
0!
0*
09
0>
0C
#932050000000
1!
1*
b10 6
19
1>
1C
b10 G
#932060000000
0!
0*
09
0>
0C
#932070000000
1!
1*
b11 6
19
1>
1C
b11 G
#932080000000
0!
0*
09
0>
0C
#932090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#932100000000
0!
0*
09
0>
0C
#932110000000
1!
1*
b101 6
19
1>
1C
b101 G
#932120000000
0!
0*
09
0>
0C
#932130000000
1!
1*
b110 6
19
1>
1C
b110 G
#932140000000
0!
0*
09
0>
0C
#932150000000
1!
1*
b111 6
19
1>
1C
b111 G
#932160000000
0!
0*
09
0>
0C
#932170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#932180000000
0!
0*
09
0>
0C
#932190000000
1!
1*
b1 6
19
1>
1C
b1 G
#932200000000
0!
0*
09
0>
0C
#932210000000
1!
1*
b10 6
19
1>
1C
b10 G
#932220000000
0!
0*
09
0>
0C
#932230000000
1!
1*
b11 6
19
1>
1C
b11 G
#932240000000
0!
0*
09
0>
0C
#932250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#932260000000
0!
0*
09
0>
0C
#932270000000
1!
1*
b101 6
19
1>
1C
b101 G
#932280000000
0!
0*
09
0>
0C
#932290000000
1!
1*
b110 6
19
1>
1C
b110 G
#932300000000
0!
0*
09
0>
0C
#932310000000
1!
1*
b111 6
19
1>
1C
b111 G
#932320000000
0!
1"
0*
1+
09
1:
0>
0C
#932330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#932340000000
0!
0*
09
0>
0C
#932350000000
1!
1*
b1 6
19
1>
1C
b1 G
#932360000000
0!
0*
09
0>
0C
#932370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#932380000000
0!
0*
09
0>
0C
#932390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#932400000000
0!
0*
09
0>
0C
#932410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#932420000000
0!
0*
09
0>
0C
#932430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#932440000000
0!
0#
0*
0,
09
0>
0?
0C
#932450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#932460000000
0!
0*
09
0>
0C
#932470000000
1!
1*
19
1>
1C
#932480000000
0!
0*
09
0>
0C
#932490000000
1!
1*
19
1>
1C
#932500000000
0!
0*
09
0>
0C
#932510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#932520000000
0!
0*
09
0>
0C
#932530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#932540000000
0!
0*
09
0>
0C
#932550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#932560000000
0!
0*
09
0>
0C
#932570000000
1!
1*
b10 6
19
1>
1C
b10 G
#932580000000
0!
0*
09
0>
0C
#932590000000
1!
1*
b11 6
19
1>
1C
b11 G
#932600000000
0!
0*
09
0>
0C
#932610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#932620000000
0!
0*
09
0>
0C
#932630000000
1!
1*
b101 6
19
1>
1C
b101 G
#932640000000
0!
0*
09
0>
0C
#932650000000
1!
1*
b110 6
19
1>
1C
b110 G
#932660000000
0!
0*
09
0>
0C
#932670000000
1!
1*
b111 6
19
1>
1C
b111 G
#932680000000
0!
0*
09
0>
0C
#932690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#932700000000
0!
0*
09
0>
0C
#932710000000
1!
1*
b1 6
19
1>
1C
b1 G
#932720000000
0!
0*
09
0>
0C
#932730000000
1!
1*
b10 6
19
1>
1C
b10 G
#932740000000
0!
0*
09
0>
0C
#932750000000
1!
1*
b11 6
19
1>
1C
b11 G
#932760000000
0!
0*
09
0>
0C
#932770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#932780000000
0!
0*
09
0>
0C
#932790000000
1!
1*
b101 6
19
1>
1C
b101 G
#932800000000
0!
0*
09
0>
0C
#932810000000
1!
1*
b110 6
19
1>
1C
b110 G
#932820000000
0!
0*
09
0>
0C
#932830000000
1!
1*
b111 6
19
1>
1C
b111 G
#932840000000
0!
0*
09
0>
0C
#932850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#932860000000
0!
0*
09
0>
0C
#932870000000
1!
1*
b1 6
19
1>
1C
b1 G
#932880000000
0!
0*
09
0>
0C
#932890000000
1!
1*
b10 6
19
1>
1C
b10 G
#932900000000
0!
0*
09
0>
0C
#932910000000
1!
1*
b11 6
19
1>
1C
b11 G
#932920000000
0!
0*
09
0>
0C
#932930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#932940000000
0!
0*
09
0>
0C
#932950000000
1!
1*
b101 6
19
1>
1C
b101 G
#932960000000
0!
0*
09
0>
0C
#932970000000
1!
1*
b110 6
19
1>
1C
b110 G
#932980000000
0!
0*
09
0>
0C
#932990000000
1!
1*
b111 6
19
1>
1C
b111 G
#933000000000
0!
1"
0*
1+
09
1:
0>
0C
#933010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#933020000000
0!
0*
09
0>
0C
#933030000000
1!
1*
b1 6
19
1>
1C
b1 G
#933040000000
0!
0*
09
0>
0C
#933050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#933060000000
0!
0*
09
0>
0C
#933070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#933080000000
0!
0*
09
0>
0C
#933090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#933100000000
0!
0*
09
0>
0C
#933110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#933120000000
0!
0#
0*
0,
09
0>
0?
0C
#933130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#933140000000
0!
0*
09
0>
0C
#933150000000
1!
1*
19
1>
1C
#933160000000
0!
0*
09
0>
0C
#933170000000
1!
1*
19
1>
1C
#933180000000
0!
0*
09
0>
0C
#933190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#933200000000
0!
0*
09
0>
0C
#933210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#933220000000
0!
0*
09
0>
0C
#933230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#933240000000
0!
0*
09
0>
0C
#933250000000
1!
1*
b10 6
19
1>
1C
b10 G
#933260000000
0!
0*
09
0>
0C
#933270000000
1!
1*
b11 6
19
1>
1C
b11 G
#933280000000
0!
0*
09
0>
0C
#933290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#933300000000
0!
0*
09
0>
0C
#933310000000
1!
1*
b101 6
19
1>
1C
b101 G
#933320000000
0!
0*
09
0>
0C
#933330000000
1!
1*
b110 6
19
1>
1C
b110 G
#933340000000
0!
0*
09
0>
0C
#933350000000
1!
1*
b111 6
19
1>
1C
b111 G
#933360000000
0!
0*
09
0>
0C
#933370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#933380000000
0!
0*
09
0>
0C
#933390000000
1!
1*
b1 6
19
1>
1C
b1 G
#933400000000
0!
0*
09
0>
0C
#933410000000
1!
1*
b10 6
19
1>
1C
b10 G
#933420000000
0!
0*
09
0>
0C
#933430000000
1!
1*
b11 6
19
1>
1C
b11 G
#933440000000
0!
0*
09
0>
0C
#933450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#933460000000
0!
0*
09
0>
0C
#933470000000
1!
1*
b101 6
19
1>
1C
b101 G
#933480000000
0!
0*
09
0>
0C
#933490000000
1!
1*
b110 6
19
1>
1C
b110 G
#933500000000
0!
0*
09
0>
0C
#933510000000
1!
1*
b111 6
19
1>
1C
b111 G
#933520000000
0!
0*
09
0>
0C
#933530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#933540000000
0!
0*
09
0>
0C
#933550000000
1!
1*
b1 6
19
1>
1C
b1 G
#933560000000
0!
0*
09
0>
0C
#933570000000
1!
1*
b10 6
19
1>
1C
b10 G
#933580000000
0!
0*
09
0>
0C
#933590000000
1!
1*
b11 6
19
1>
1C
b11 G
#933600000000
0!
0*
09
0>
0C
#933610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#933620000000
0!
0*
09
0>
0C
#933630000000
1!
1*
b101 6
19
1>
1C
b101 G
#933640000000
0!
0*
09
0>
0C
#933650000000
1!
1*
b110 6
19
1>
1C
b110 G
#933660000000
0!
0*
09
0>
0C
#933670000000
1!
1*
b111 6
19
1>
1C
b111 G
#933680000000
0!
1"
0*
1+
09
1:
0>
0C
#933690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#933700000000
0!
0*
09
0>
0C
#933710000000
1!
1*
b1 6
19
1>
1C
b1 G
#933720000000
0!
0*
09
0>
0C
#933730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#933740000000
0!
0*
09
0>
0C
#933750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#933760000000
0!
0*
09
0>
0C
#933770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#933780000000
0!
0*
09
0>
0C
#933790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#933800000000
0!
0#
0*
0,
09
0>
0?
0C
#933810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#933820000000
0!
0*
09
0>
0C
#933830000000
1!
1*
19
1>
1C
#933840000000
0!
0*
09
0>
0C
#933850000000
1!
1*
19
1>
1C
#933860000000
0!
0*
09
0>
0C
#933870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#933880000000
0!
0*
09
0>
0C
#933890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#933900000000
0!
0*
09
0>
0C
#933910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#933920000000
0!
0*
09
0>
0C
#933930000000
1!
1*
b10 6
19
1>
1C
b10 G
#933940000000
0!
0*
09
0>
0C
#933950000000
1!
1*
b11 6
19
1>
1C
b11 G
#933960000000
0!
0*
09
0>
0C
#933970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#933980000000
0!
0*
09
0>
0C
#933990000000
1!
1*
b101 6
19
1>
1C
b101 G
#934000000000
0!
0*
09
0>
0C
#934010000000
1!
1*
b110 6
19
1>
1C
b110 G
#934020000000
0!
0*
09
0>
0C
#934030000000
1!
1*
b111 6
19
1>
1C
b111 G
#934040000000
0!
0*
09
0>
0C
#934050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#934060000000
0!
0*
09
0>
0C
#934070000000
1!
1*
b1 6
19
1>
1C
b1 G
#934080000000
0!
0*
09
0>
0C
#934090000000
1!
1*
b10 6
19
1>
1C
b10 G
#934100000000
0!
0*
09
0>
0C
#934110000000
1!
1*
b11 6
19
1>
1C
b11 G
#934120000000
0!
0*
09
0>
0C
#934130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#934140000000
0!
0*
09
0>
0C
#934150000000
1!
1*
b101 6
19
1>
1C
b101 G
#934160000000
0!
0*
09
0>
0C
#934170000000
1!
1*
b110 6
19
1>
1C
b110 G
#934180000000
0!
0*
09
0>
0C
#934190000000
1!
1*
b111 6
19
1>
1C
b111 G
#934200000000
0!
0*
09
0>
0C
#934210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#934220000000
0!
0*
09
0>
0C
#934230000000
1!
1*
b1 6
19
1>
1C
b1 G
#934240000000
0!
0*
09
0>
0C
#934250000000
1!
1*
b10 6
19
1>
1C
b10 G
#934260000000
0!
0*
09
0>
0C
#934270000000
1!
1*
b11 6
19
1>
1C
b11 G
#934280000000
0!
0*
09
0>
0C
#934290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#934300000000
0!
0*
09
0>
0C
#934310000000
1!
1*
b101 6
19
1>
1C
b101 G
#934320000000
0!
0*
09
0>
0C
#934330000000
1!
1*
b110 6
19
1>
1C
b110 G
#934340000000
0!
0*
09
0>
0C
#934350000000
1!
1*
b111 6
19
1>
1C
b111 G
#934360000000
0!
1"
0*
1+
09
1:
0>
0C
#934370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#934380000000
0!
0*
09
0>
0C
#934390000000
1!
1*
b1 6
19
1>
1C
b1 G
#934400000000
0!
0*
09
0>
0C
#934410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#934420000000
0!
0*
09
0>
0C
#934430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#934440000000
0!
0*
09
0>
0C
#934450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#934460000000
0!
0*
09
0>
0C
#934470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#934480000000
0!
0#
0*
0,
09
0>
0?
0C
#934490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#934500000000
0!
0*
09
0>
0C
#934510000000
1!
1*
19
1>
1C
#934520000000
0!
0*
09
0>
0C
#934530000000
1!
1*
19
1>
1C
#934540000000
0!
0*
09
0>
0C
#934550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#934560000000
0!
0*
09
0>
0C
#934570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#934580000000
0!
0*
09
0>
0C
#934590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#934600000000
0!
0*
09
0>
0C
#934610000000
1!
1*
b10 6
19
1>
1C
b10 G
#934620000000
0!
0*
09
0>
0C
#934630000000
1!
1*
b11 6
19
1>
1C
b11 G
#934640000000
0!
0*
09
0>
0C
#934650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#934660000000
0!
0*
09
0>
0C
#934670000000
1!
1*
b101 6
19
1>
1C
b101 G
#934680000000
0!
0*
09
0>
0C
#934690000000
1!
1*
b110 6
19
1>
1C
b110 G
#934700000000
0!
0*
09
0>
0C
#934710000000
1!
1*
b111 6
19
1>
1C
b111 G
#934720000000
0!
0*
09
0>
0C
#934730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#934740000000
0!
0*
09
0>
0C
#934750000000
1!
1*
b1 6
19
1>
1C
b1 G
#934760000000
0!
0*
09
0>
0C
#934770000000
1!
1*
b10 6
19
1>
1C
b10 G
#934780000000
0!
0*
09
0>
0C
#934790000000
1!
1*
b11 6
19
1>
1C
b11 G
#934800000000
0!
0*
09
0>
0C
#934810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#934820000000
0!
0*
09
0>
0C
#934830000000
1!
1*
b101 6
19
1>
1C
b101 G
#934840000000
0!
0*
09
0>
0C
#934850000000
1!
1*
b110 6
19
1>
1C
b110 G
#934860000000
0!
0*
09
0>
0C
#934870000000
1!
1*
b111 6
19
1>
1C
b111 G
#934880000000
0!
0*
09
0>
0C
#934890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#934900000000
0!
0*
09
0>
0C
#934910000000
1!
1*
b1 6
19
1>
1C
b1 G
#934920000000
0!
0*
09
0>
0C
#934930000000
1!
1*
b10 6
19
1>
1C
b10 G
#934940000000
0!
0*
09
0>
0C
#934950000000
1!
1*
b11 6
19
1>
1C
b11 G
#934960000000
0!
0*
09
0>
0C
#934970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#934980000000
0!
0*
09
0>
0C
#934990000000
1!
1*
b101 6
19
1>
1C
b101 G
#935000000000
0!
0*
09
0>
0C
#935010000000
1!
1*
b110 6
19
1>
1C
b110 G
#935020000000
0!
0*
09
0>
0C
#935030000000
1!
1*
b111 6
19
1>
1C
b111 G
#935040000000
0!
1"
0*
1+
09
1:
0>
0C
#935050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#935060000000
0!
0*
09
0>
0C
#935070000000
1!
1*
b1 6
19
1>
1C
b1 G
#935080000000
0!
0*
09
0>
0C
#935090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#935100000000
0!
0*
09
0>
0C
#935110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#935120000000
0!
0*
09
0>
0C
#935130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#935140000000
0!
0*
09
0>
0C
#935150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#935160000000
0!
0#
0*
0,
09
0>
0?
0C
#935170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#935180000000
0!
0*
09
0>
0C
#935190000000
1!
1*
19
1>
1C
#935200000000
0!
0*
09
0>
0C
#935210000000
1!
1*
19
1>
1C
#935220000000
0!
0*
09
0>
0C
#935230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#935240000000
0!
0*
09
0>
0C
#935250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#935260000000
0!
0*
09
0>
0C
#935270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#935280000000
0!
0*
09
0>
0C
#935290000000
1!
1*
b10 6
19
1>
1C
b10 G
#935300000000
0!
0*
09
0>
0C
#935310000000
1!
1*
b11 6
19
1>
1C
b11 G
#935320000000
0!
0*
09
0>
0C
#935330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#935340000000
0!
0*
09
0>
0C
#935350000000
1!
1*
b101 6
19
1>
1C
b101 G
#935360000000
0!
0*
09
0>
0C
#935370000000
1!
1*
b110 6
19
1>
1C
b110 G
#935380000000
0!
0*
09
0>
0C
#935390000000
1!
1*
b111 6
19
1>
1C
b111 G
#935400000000
0!
0*
09
0>
0C
#935410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#935420000000
0!
0*
09
0>
0C
#935430000000
1!
1*
b1 6
19
1>
1C
b1 G
#935440000000
0!
0*
09
0>
0C
#935450000000
1!
1*
b10 6
19
1>
1C
b10 G
#935460000000
0!
0*
09
0>
0C
#935470000000
1!
1*
b11 6
19
1>
1C
b11 G
#935480000000
0!
0*
09
0>
0C
#935490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#935500000000
0!
0*
09
0>
0C
#935510000000
1!
1*
b101 6
19
1>
1C
b101 G
#935520000000
0!
0*
09
0>
0C
#935530000000
1!
1*
b110 6
19
1>
1C
b110 G
#935540000000
0!
0*
09
0>
0C
#935550000000
1!
1*
b111 6
19
1>
1C
b111 G
#935560000000
0!
0*
09
0>
0C
#935570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#935580000000
0!
0*
09
0>
0C
#935590000000
1!
1*
b1 6
19
1>
1C
b1 G
#935600000000
0!
0*
09
0>
0C
#935610000000
1!
1*
b10 6
19
1>
1C
b10 G
#935620000000
0!
0*
09
0>
0C
#935630000000
1!
1*
b11 6
19
1>
1C
b11 G
#935640000000
0!
0*
09
0>
0C
#935650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#935660000000
0!
0*
09
0>
0C
#935670000000
1!
1*
b101 6
19
1>
1C
b101 G
#935680000000
0!
0*
09
0>
0C
#935690000000
1!
1*
b110 6
19
1>
1C
b110 G
#935700000000
0!
0*
09
0>
0C
#935710000000
1!
1*
b111 6
19
1>
1C
b111 G
#935720000000
0!
1"
0*
1+
09
1:
0>
0C
#935730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#935740000000
0!
0*
09
0>
0C
#935750000000
1!
1*
b1 6
19
1>
1C
b1 G
#935760000000
0!
0*
09
0>
0C
#935770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#935780000000
0!
0*
09
0>
0C
#935790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#935800000000
0!
0*
09
0>
0C
#935810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#935820000000
0!
0*
09
0>
0C
#935830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#935840000000
0!
0#
0*
0,
09
0>
0?
0C
#935850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#935860000000
0!
0*
09
0>
0C
#935870000000
1!
1*
19
1>
1C
#935880000000
0!
0*
09
0>
0C
#935890000000
1!
1*
19
1>
1C
#935900000000
0!
0*
09
0>
0C
#935910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#935920000000
0!
0*
09
0>
0C
#935930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#935940000000
0!
0*
09
0>
0C
#935950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#935960000000
0!
0*
09
0>
0C
#935970000000
1!
1*
b10 6
19
1>
1C
b10 G
#935980000000
0!
0*
09
0>
0C
#935990000000
1!
1*
b11 6
19
1>
1C
b11 G
#936000000000
0!
0*
09
0>
0C
#936010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#936020000000
0!
0*
09
0>
0C
#936030000000
1!
1*
b101 6
19
1>
1C
b101 G
#936040000000
0!
0*
09
0>
0C
#936050000000
1!
1*
b110 6
19
1>
1C
b110 G
#936060000000
0!
0*
09
0>
0C
#936070000000
1!
1*
b111 6
19
1>
1C
b111 G
#936080000000
0!
0*
09
0>
0C
#936090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#936100000000
0!
0*
09
0>
0C
#936110000000
1!
1*
b1 6
19
1>
1C
b1 G
#936120000000
0!
0*
09
0>
0C
#936130000000
1!
1*
b10 6
19
1>
1C
b10 G
#936140000000
0!
0*
09
0>
0C
#936150000000
1!
1*
b11 6
19
1>
1C
b11 G
#936160000000
0!
0*
09
0>
0C
#936170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#936180000000
0!
0*
09
0>
0C
#936190000000
1!
1*
b101 6
19
1>
1C
b101 G
#936200000000
0!
0*
09
0>
0C
#936210000000
1!
1*
b110 6
19
1>
1C
b110 G
#936220000000
0!
0*
09
0>
0C
#936230000000
1!
1*
b111 6
19
1>
1C
b111 G
#936240000000
0!
0*
09
0>
0C
#936250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#936260000000
0!
0*
09
0>
0C
#936270000000
1!
1*
b1 6
19
1>
1C
b1 G
#936280000000
0!
0*
09
0>
0C
#936290000000
1!
1*
b10 6
19
1>
1C
b10 G
#936300000000
0!
0*
09
0>
0C
#936310000000
1!
1*
b11 6
19
1>
1C
b11 G
#936320000000
0!
0*
09
0>
0C
#936330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#936340000000
0!
0*
09
0>
0C
#936350000000
1!
1*
b101 6
19
1>
1C
b101 G
#936360000000
0!
0*
09
0>
0C
#936370000000
1!
1*
b110 6
19
1>
1C
b110 G
#936380000000
0!
0*
09
0>
0C
#936390000000
1!
1*
b111 6
19
1>
1C
b111 G
#936400000000
0!
1"
0*
1+
09
1:
0>
0C
#936410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#936420000000
0!
0*
09
0>
0C
#936430000000
1!
1*
b1 6
19
1>
1C
b1 G
#936440000000
0!
0*
09
0>
0C
#936450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#936460000000
0!
0*
09
0>
0C
#936470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#936480000000
0!
0*
09
0>
0C
#936490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#936500000000
0!
0*
09
0>
0C
#936510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#936520000000
0!
0#
0*
0,
09
0>
0?
0C
#936530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#936540000000
0!
0*
09
0>
0C
#936550000000
1!
1*
19
1>
1C
#936560000000
0!
0*
09
0>
0C
#936570000000
1!
1*
19
1>
1C
#936580000000
0!
0*
09
0>
0C
#936590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#936600000000
0!
0*
09
0>
0C
#936610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#936620000000
0!
0*
09
0>
0C
#936630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#936640000000
0!
0*
09
0>
0C
#936650000000
1!
1*
b10 6
19
1>
1C
b10 G
#936660000000
0!
0*
09
0>
0C
#936670000000
1!
1*
b11 6
19
1>
1C
b11 G
#936680000000
0!
0*
09
0>
0C
#936690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#936700000000
0!
0*
09
0>
0C
#936710000000
1!
1*
b101 6
19
1>
1C
b101 G
#936720000000
0!
0*
09
0>
0C
#936730000000
1!
1*
b110 6
19
1>
1C
b110 G
#936740000000
0!
0*
09
0>
0C
#936750000000
1!
1*
b111 6
19
1>
1C
b111 G
#936760000000
0!
0*
09
0>
0C
#936770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#936780000000
0!
0*
09
0>
0C
#936790000000
1!
1*
b1 6
19
1>
1C
b1 G
#936800000000
0!
0*
09
0>
0C
#936810000000
1!
1*
b10 6
19
1>
1C
b10 G
#936820000000
0!
0*
09
0>
0C
#936830000000
1!
1*
b11 6
19
1>
1C
b11 G
#936840000000
0!
0*
09
0>
0C
#936850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#936860000000
0!
0*
09
0>
0C
#936870000000
1!
1*
b101 6
19
1>
1C
b101 G
#936880000000
0!
0*
09
0>
0C
#936890000000
1!
1*
b110 6
19
1>
1C
b110 G
#936900000000
0!
0*
09
0>
0C
#936910000000
1!
1*
b111 6
19
1>
1C
b111 G
#936920000000
0!
0*
09
0>
0C
#936930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#936940000000
0!
0*
09
0>
0C
#936950000000
1!
1*
b1 6
19
1>
1C
b1 G
#936960000000
0!
0*
09
0>
0C
#936970000000
1!
1*
b10 6
19
1>
1C
b10 G
#936980000000
0!
0*
09
0>
0C
#936990000000
1!
1*
b11 6
19
1>
1C
b11 G
#937000000000
0!
0*
09
0>
0C
#937010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#937020000000
0!
0*
09
0>
0C
#937030000000
1!
1*
b101 6
19
1>
1C
b101 G
#937040000000
0!
0*
09
0>
0C
#937050000000
1!
1*
b110 6
19
1>
1C
b110 G
#937060000000
0!
0*
09
0>
0C
#937070000000
1!
1*
b111 6
19
1>
1C
b111 G
#937080000000
0!
1"
0*
1+
09
1:
0>
0C
#937090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#937100000000
0!
0*
09
0>
0C
#937110000000
1!
1*
b1 6
19
1>
1C
b1 G
#937120000000
0!
0*
09
0>
0C
#937130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#937140000000
0!
0*
09
0>
0C
#937150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#937160000000
0!
0*
09
0>
0C
#937170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#937180000000
0!
0*
09
0>
0C
#937190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#937200000000
0!
0#
0*
0,
09
0>
0?
0C
#937210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#937220000000
0!
0*
09
0>
0C
#937230000000
1!
1*
19
1>
1C
#937240000000
0!
0*
09
0>
0C
#937250000000
1!
1*
19
1>
1C
#937260000000
0!
0*
09
0>
0C
#937270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#937280000000
0!
0*
09
0>
0C
#937290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#937300000000
0!
0*
09
0>
0C
#937310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#937320000000
0!
0*
09
0>
0C
#937330000000
1!
1*
b10 6
19
1>
1C
b10 G
#937340000000
0!
0*
09
0>
0C
#937350000000
1!
1*
b11 6
19
1>
1C
b11 G
#937360000000
0!
0*
09
0>
0C
#937370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#937380000000
0!
0*
09
0>
0C
#937390000000
1!
1*
b101 6
19
1>
1C
b101 G
#937400000000
0!
0*
09
0>
0C
#937410000000
1!
1*
b110 6
19
1>
1C
b110 G
#937420000000
0!
0*
09
0>
0C
#937430000000
1!
1*
b111 6
19
1>
1C
b111 G
#937440000000
0!
0*
09
0>
0C
#937450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#937460000000
0!
0*
09
0>
0C
#937470000000
1!
1*
b1 6
19
1>
1C
b1 G
#937480000000
0!
0*
09
0>
0C
#937490000000
1!
1*
b10 6
19
1>
1C
b10 G
#937500000000
0!
0*
09
0>
0C
#937510000000
1!
1*
b11 6
19
1>
1C
b11 G
#937520000000
0!
0*
09
0>
0C
#937530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#937540000000
0!
0*
09
0>
0C
#937550000000
1!
1*
b101 6
19
1>
1C
b101 G
#937560000000
0!
0*
09
0>
0C
#937570000000
1!
1*
b110 6
19
1>
1C
b110 G
#937580000000
0!
0*
09
0>
0C
#937590000000
1!
1*
b111 6
19
1>
1C
b111 G
#937600000000
0!
0*
09
0>
0C
#937610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#937620000000
0!
0*
09
0>
0C
#937630000000
1!
1*
b1 6
19
1>
1C
b1 G
#937640000000
0!
0*
09
0>
0C
#937650000000
1!
1*
b10 6
19
1>
1C
b10 G
#937660000000
0!
0*
09
0>
0C
#937670000000
1!
1*
b11 6
19
1>
1C
b11 G
#937680000000
0!
0*
09
0>
0C
#937690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#937700000000
0!
0*
09
0>
0C
#937710000000
1!
1*
b101 6
19
1>
1C
b101 G
#937720000000
0!
0*
09
0>
0C
#937730000000
1!
1*
b110 6
19
1>
1C
b110 G
#937740000000
0!
0*
09
0>
0C
#937750000000
1!
1*
b111 6
19
1>
1C
b111 G
#937760000000
0!
1"
0*
1+
09
1:
0>
0C
#937770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#937780000000
0!
0*
09
0>
0C
#937790000000
1!
1*
b1 6
19
1>
1C
b1 G
#937800000000
0!
0*
09
0>
0C
#937810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#937820000000
0!
0*
09
0>
0C
#937830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#937840000000
0!
0*
09
0>
0C
#937850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#937860000000
0!
0*
09
0>
0C
#937870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#937880000000
0!
0#
0*
0,
09
0>
0?
0C
#937890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#937900000000
0!
0*
09
0>
0C
#937910000000
1!
1*
19
1>
1C
#937920000000
0!
0*
09
0>
0C
#937930000000
1!
1*
19
1>
1C
#937940000000
0!
0*
09
0>
0C
#937950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#937960000000
0!
0*
09
0>
0C
#937970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#937980000000
0!
0*
09
0>
0C
#937990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#938000000000
0!
0*
09
0>
0C
#938010000000
1!
1*
b10 6
19
1>
1C
b10 G
#938020000000
0!
0*
09
0>
0C
#938030000000
1!
1*
b11 6
19
1>
1C
b11 G
#938040000000
0!
0*
09
0>
0C
#938050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#938060000000
0!
0*
09
0>
0C
#938070000000
1!
1*
b101 6
19
1>
1C
b101 G
#938080000000
0!
0*
09
0>
0C
#938090000000
1!
1*
b110 6
19
1>
1C
b110 G
#938100000000
0!
0*
09
0>
0C
#938110000000
1!
1*
b111 6
19
1>
1C
b111 G
#938120000000
0!
0*
09
0>
0C
#938130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#938140000000
0!
0*
09
0>
0C
#938150000000
1!
1*
b1 6
19
1>
1C
b1 G
#938160000000
0!
0*
09
0>
0C
#938170000000
1!
1*
b10 6
19
1>
1C
b10 G
#938180000000
0!
0*
09
0>
0C
#938190000000
1!
1*
b11 6
19
1>
1C
b11 G
#938200000000
0!
0*
09
0>
0C
#938210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#938220000000
0!
0*
09
0>
0C
#938230000000
1!
1*
b101 6
19
1>
1C
b101 G
#938240000000
0!
0*
09
0>
0C
#938250000000
1!
1*
b110 6
19
1>
1C
b110 G
#938260000000
0!
0*
09
0>
0C
#938270000000
1!
1*
b111 6
19
1>
1C
b111 G
#938280000000
0!
0*
09
0>
0C
#938290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#938300000000
0!
0*
09
0>
0C
#938310000000
1!
1*
b1 6
19
1>
1C
b1 G
#938320000000
0!
0*
09
0>
0C
#938330000000
1!
1*
b10 6
19
1>
1C
b10 G
#938340000000
0!
0*
09
0>
0C
#938350000000
1!
1*
b11 6
19
1>
1C
b11 G
#938360000000
0!
0*
09
0>
0C
#938370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#938380000000
0!
0*
09
0>
0C
#938390000000
1!
1*
b101 6
19
1>
1C
b101 G
#938400000000
0!
0*
09
0>
0C
#938410000000
1!
1*
b110 6
19
1>
1C
b110 G
#938420000000
0!
0*
09
0>
0C
#938430000000
1!
1*
b111 6
19
1>
1C
b111 G
#938440000000
0!
1"
0*
1+
09
1:
0>
0C
#938450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#938460000000
0!
0*
09
0>
0C
#938470000000
1!
1*
b1 6
19
1>
1C
b1 G
#938480000000
0!
0*
09
0>
0C
#938490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#938500000000
0!
0*
09
0>
0C
#938510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#938520000000
0!
0*
09
0>
0C
#938530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#938540000000
0!
0*
09
0>
0C
#938550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#938560000000
0!
0#
0*
0,
09
0>
0?
0C
#938570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#938580000000
0!
0*
09
0>
0C
#938590000000
1!
1*
19
1>
1C
#938600000000
0!
0*
09
0>
0C
#938610000000
1!
1*
19
1>
1C
#938620000000
0!
0*
09
0>
0C
#938630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#938640000000
0!
0*
09
0>
0C
#938650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#938660000000
0!
0*
09
0>
0C
#938670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#938680000000
0!
0*
09
0>
0C
#938690000000
1!
1*
b10 6
19
1>
1C
b10 G
#938700000000
0!
0*
09
0>
0C
#938710000000
1!
1*
b11 6
19
1>
1C
b11 G
#938720000000
0!
0*
09
0>
0C
#938730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#938740000000
0!
0*
09
0>
0C
#938750000000
1!
1*
b101 6
19
1>
1C
b101 G
#938760000000
0!
0*
09
0>
0C
#938770000000
1!
1*
b110 6
19
1>
1C
b110 G
#938780000000
0!
0*
09
0>
0C
#938790000000
1!
1*
b111 6
19
1>
1C
b111 G
#938800000000
0!
0*
09
0>
0C
#938810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#938820000000
0!
0*
09
0>
0C
#938830000000
1!
1*
b1 6
19
1>
1C
b1 G
#938840000000
0!
0*
09
0>
0C
#938850000000
1!
1*
b10 6
19
1>
1C
b10 G
#938860000000
0!
0*
09
0>
0C
#938870000000
1!
1*
b11 6
19
1>
1C
b11 G
#938880000000
0!
0*
09
0>
0C
#938890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#938900000000
0!
0*
09
0>
0C
#938910000000
1!
1*
b101 6
19
1>
1C
b101 G
#938920000000
0!
0*
09
0>
0C
#938930000000
1!
1*
b110 6
19
1>
1C
b110 G
#938940000000
0!
0*
09
0>
0C
#938950000000
1!
1*
b111 6
19
1>
1C
b111 G
#938960000000
0!
0*
09
0>
0C
#938970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#938980000000
0!
0*
09
0>
0C
#938990000000
1!
1*
b1 6
19
1>
1C
b1 G
#939000000000
0!
0*
09
0>
0C
#939010000000
1!
1*
b10 6
19
1>
1C
b10 G
#939020000000
0!
0*
09
0>
0C
#939030000000
1!
1*
b11 6
19
1>
1C
b11 G
#939040000000
0!
0*
09
0>
0C
#939050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#939060000000
0!
0*
09
0>
0C
#939070000000
1!
1*
b101 6
19
1>
1C
b101 G
#939080000000
0!
0*
09
0>
0C
#939090000000
1!
1*
b110 6
19
1>
1C
b110 G
#939100000000
0!
0*
09
0>
0C
#939110000000
1!
1*
b111 6
19
1>
1C
b111 G
#939120000000
0!
1"
0*
1+
09
1:
0>
0C
#939130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#939140000000
0!
0*
09
0>
0C
#939150000000
1!
1*
b1 6
19
1>
1C
b1 G
#939160000000
0!
0*
09
0>
0C
#939170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#939180000000
0!
0*
09
0>
0C
#939190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#939200000000
0!
0*
09
0>
0C
#939210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#939220000000
0!
0*
09
0>
0C
#939230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#939240000000
0!
0#
0*
0,
09
0>
0?
0C
#939250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#939260000000
0!
0*
09
0>
0C
#939270000000
1!
1*
19
1>
1C
#939280000000
0!
0*
09
0>
0C
#939290000000
1!
1*
19
1>
1C
#939300000000
0!
0*
09
0>
0C
#939310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#939320000000
0!
0*
09
0>
0C
#939330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#939340000000
0!
0*
09
0>
0C
#939350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#939360000000
0!
0*
09
0>
0C
#939370000000
1!
1*
b10 6
19
1>
1C
b10 G
#939380000000
0!
0*
09
0>
0C
#939390000000
1!
1*
b11 6
19
1>
1C
b11 G
#939400000000
0!
0*
09
0>
0C
#939410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#939420000000
0!
0*
09
0>
0C
#939430000000
1!
1*
b101 6
19
1>
1C
b101 G
#939440000000
0!
0*
09
0>
0C
#939450000000
1!
1*
b110 6
19
1>
1C
b110 G
#939460000000
0!
0*
09
0>
0C
#939470000000
1!
1*
b111 6
19
1>
1C
b111 G
#939480000000
0!
0*
09
0>
0C
#939490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#939500000000
0!
0*
09
0>
0C
#939510000000
1!
1*
b1 6
19
1>
1C
b1 G
#939520000000
0!
0*
09
0>
0C
#939530000000
1!
1*
b10 6
19
1>
1C
b10 G
#939540000000
0!
0*
09
0>
0C
#939550000000
1!
1*
b11 6
19
1>
1C
b11 G
#939560000000
0!
0*
09
0>
0C
#939570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#939580000000
0!
0*
09
0>
0C
#939590000000
1!
1*
b101 6
19
1>
1C
b101 G
#939600000000
0!
0*
09
0>
0C
#939610000000
1!
1*
b110 6
19
1>
1C
b110 G
#939620000000
0!
0*
09
0>
0C
#939630000000
1!
1*
b111 6
19
1>
1C
b111 G
#939640000000
0!
0*
09
0>
0C
#939650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#939660000000
0!
0*
09
0>
0C
#939670000000
1!
1*
b1 6
19
1>
1C
b1 G
#939680000000
0!
0*
09
0>
0C
#939690000000
1!
1*
b10 6
19
1>
1C
b10 G
#939700000000
0!
0*
09
0>
0C
#939710000000
1!
1*
b11 6
19
1>
1C
b11 G
#939720000000
0!
0*
09
0>
0C
#939730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#939740000000
0!
0*
09
0>
0C
#939750000000
1!
1*
b101 6
19
1>
1C
b101 G
#939760000000
0!
0*
09
0>
0C
#939770000000
1!
1*
b110 6
19
1>
1C
b110 G
#939780000000
0!
0*
09
0>
0C
#939790000000
1!
1*
b111 6
19
1>
1C
b111 G
#939800000000
0!
1"
0*
1+
09
1:
0>
0C
#939810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#939820000000
0!
0*
09
0>
0C
#939830000000
1!
1*
b1 6
19
1>
1C
b1 G
#939840000000
0!
0*
09
0>
0C
#939850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#939860000000
0!
0*
09
0>
0C
#939870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#939880000000
0!
0*
09
0>
0C
#939890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#939900000000
0!
0*
09
0>
0C
#939910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#939920000000
0!
0#
0*
0,
09
0>
0?
0C
#939930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#939940000000
0!
0*
09
0>
0C
#939950000000
1!
1*
19
1>
1C
#939960000000
0!
0*
09
0>
0C
#939970000000
1!
1*
19
1>
1C
#939980000000
0!
0*
09
0>
0C
#939990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#940000000000
0!
0*
09
0>
0C
#940010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#940020000000
0!
0*
09
0>
0C
#940030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#940040000000
0!
0*
09
0>
0C
#940050000000
1!
1*
b10 6
19
1>
1C
b10 G
#940060000000
0!
0*
09
0>
0C
#940070000000
1!
1*
b11 6
19
1>
1C
b11 G
#940080000000
0!
0*
09
0>
0C
#940090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#940100000000
0!
0*
09
0>
0C
#940110000000
1!
1*
b101 6
19
1>
1C
b101 G
#940120000000
0!
0*
09
0>
0C
#940130000000
1!
1*
b110 6
19
1>
1C
b110 G
#940140000000
0!
0*
09
0>
0C
#940150000000
1!
1*
b111 6
19
1>
1C
b111 G
#940160000000
0!
0*
09
0>
0C
#940170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#940180000000
0!
0*
09
0>
0C
#940190000000
1!
1*
b1 6
19
1>
1C
b1 G
#940200000000
0!
0*
09
0>
0C
#940210000000
1!
1*
b10 6
19
1>
1C
b10 G
#940220000000
0!
0*
09
0>
0C
#940230000000
1!
1*
b11 6
19
1>
1C
b11 G
#940240000000
0!
0*
09
0>
0C
#940250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#940260000000
0!
0*
09
0>
0C
#940270000000
1!
1*
b101 6
19
1>
1C
b101 G
#940280000000
0!
0*
09
0>
0C
#940290000000
1!
1*
b110 6
19
1>
1C
b110 G
#940300000000
0!
0*
09
0>
0C
#940310000000
1!
1*
b111 6
19
1>
1C
b111 G
#940320000000
0!
0*
09
0>
0C
#940330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#940340000000
0!
0*
09
0>
0C
#940350000000
1!
1*
b1 6
19
1>
1C
b1 G
#940360000000
0!
0*
09
0>
0C
#940370000000
1!
1*
b10 6
19
1>
1C
b10 G
#940380000000
0!
0*
09
0>
0C
#940390000000
1!
1*
b11 6
19
1>
1C
b11 G
#940400000000
0!
0*
09
0>
0C
#940410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#940420000000
0!
0*
09
0>
0C
#940430000000
1!
1*
b101 6
19
1>
1C
b101 G
#940440000000
0!
0*
09
0>
0C
#940450000000
1!
1*
b110 6
19
1>
1C
b110 G
#940460000000
0!
0*
09
0>
0C
#940470000000
1!
1*
b111 6
19
1>
1C
b111 G
#940480000000
0!
1"
0*
1+
09
1:
0>
0C
#940490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#940500000000
0!
0*
09
0>
0C
#940510000000
1!
1*
b1 6
19
1>
1C
b1 G
#940520000000
0!
0*
09
0>
0C
#940530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#940540000000
0!
0*
09
0>
0C
#940550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#940560000000
0!
0*
09
0>
0C
#940570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#940580000000
0!
0*
09
0>
0C
#940590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#940600000000
0!
0#
0*
0,
09
0>
0?
0C
#940610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#940620000000
0!
0*
09
0>
0C
#940630000000
1!
1*
19
1>
1C
#940640000000
0!
0*
09
0>
0C
#940650000000
1!
1*
19
1>
1C
#940660000000
0!
0*
09
0>
0C
#940670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#940680000000
0!
0*
09
0>
0C
#940690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#940700000000
0!
0*
09
0>
0C
#940710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#940720000000
0!
0*
09
0>
0C
#940730000000
1!
1*
b10 6
19
1>
1C
b10 G
#940740000000
0!
0*
09
0>
0C
#940750000000
1!
1*
b11 6
19
1>
1C
b11 G
#940760000000
0!
0*
09
0>
0C
#940770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#940780000000
0!
0*
09
0>
0C
#940790000000
1!
1*
b101 6
19
1>
1C
b101 G
#940800000000
0!
0*
09
0>
0C
#940810000000
1!
1*
b110 6
19
1>
1C
b110 G
#940820000000
0!
0*
09
0>
0C
#940830000000
1!
1*
b111 6
19
1>
1C
b111 G
#940840000000
0!
0*
09
0>
0C
#940850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#940860000000
0!
0*
09
0>
0C
#940870000000
1!
1*
b1 6
19
1>
1C
b1 G
#940880000000
0!
0*
09
0>
0C
#940890000000
1!
1*
b10 6
19
1>
1C
b10 G
#940900000000
0!
0*
09
0>
0C
#940910000000
1!
1*
b11 6
19
1>
1C
b11 G
#940920000000
0!
0*
09
0>
0C
#940930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#940940000000
0!
0*
09
0>
0C
#940950000000
1!
1*
b101 6
19
1>
1C
b101 G
#940960000000
0!
0*
09
0>
0C
#940970000000
1!
1*
b110 6
19
1>
1C
b110 G
#940980000000
0!
0*
09
0>
0C
#940990000000
1!
1*
b111 6
19
1>
1C
b111 G
#941000000000
0!
0*
09
0>
0C
#941010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#941020000000
0!
0*
09
0>
0C
#941030000000
1!
1*
b1 6
19
1>
1C
b1 G
#941040000000
0!
0*
09
0>
0C
#941050000000
1!
1*
b10 6
19
1>
1C
b10 G
#941060000000
0!
0*
09
0>
0C
#941070000000
1!
1*
b11 6
19
1>
1C
b11 G
#941080000000
0!
0*
09
0>
0C
#941090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#941100000000
0!
0*
09
0>
0C
#941110000000
1!
1*
b101 6
19
1>
1C
b101 G
#941120000000
0!
0*
09
0>
0C
#941130000000
1!
1*
b110 6
19
1>
1C
b110 G
#941140000000
0!
0*
09
0>
0C
#941150000000
1!
1*
b111 6
19
1>
1C
b111 G
#941160000000
0!
1"
0*
1+
09
1:
0>
0C
#941170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#941180000000
0!
0*
09
0>
0C
#941190000000
1!
1*
b1 6
19
1>
1C
b1 G
#941200000000
0!
0*
09
0>
0C
#941210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#941220000000
0!
0*
09
0>
0C
#941230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#941240000000
0!
0*
09
0>
0C
#941250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#941260000000
0!
0*
09
0>
0C
#941270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#941280000000
0!
0#
0*
0,
09
0>
0?
0C
#941290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#941300000000
0!
0*
09
0>
0C
#941310000000
1!
1*
19
1>
1C
#941320000000
0!
0*
09
0>
0C
#941330000000
1!
1*
19
1>
1C
#941340000000
0!
0*
09
0>
0C
#941350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#941360000000
0!
0*
09
0>
0C
#941370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#941380000000
0!
0*
09
0>
0C
#941390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#941400000000
0!
0*
09
0>
0C
#941410000000
1!
1*
b10 6
19
1>
1C
b10 G
#941420000000
0!
0*
09
0>
0C
#941430000000
1!
1*
b11 6
19
1>
1C
b11 G
#941440000000
0!
0*
09
0>
0C
#941450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#941460000000
0!
0*
09
0>
0C
#941470000000
1!
1*
b101 6
19
1>
1C
b101 G
#941480000000
0!
0*
09
0>
0C
#941490000000
1!
1*
b110 6
19
1>
1C
b110 G
#941500000000
0!
0*
09
0>
0C
#941510000000
1!
1*
b111 6
19
1>
1C
b111 G
#941520000000
0!
0*
09
0>
0C
#941530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#941540000000
0!
0*
09
0>
0C
#941550000000
1!
1*
b1 6
19
1>
1C
b1 G
#941560000000
0!
0*
09
0>
0C
#941570000000
1!
1*
b10 6
19
1>
1C
b10 G
#941580000000
0!
0*
09
0>
0C
#941590000000
1!
1*
b11 6
19
1>
1C
b11 G
#941600000000
0!
0*
09
0>
0C
#941610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#941620000000
0!
0*
09
0>
0C
#941630000000
1!
1*
b101 6
19
1>
1C
b101 G
#941640000000
0!
0*
09
0>
0C
#941650000000
1!
1*
b110 6
19
1>
1C
b110 G
#941660000000
0!
0*
09
0>
0C
#941670000000
1!
1*
b111 6
19
1>
1C
b111 G
#941680000000
0!
0*
09
0>
0C
#941690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#941700000000
0!
0*
09
0>
0C
#941710000000
1!
1*
b1 6
19
1>
1C
b1 G
#941720000000
0!
0*
09
0>
0C
#941730000000
1!
1*
b10 6
19
1>
1C
b10 G
#941740000000
0!
0*
09
0>
0C
#941750000000
1!
1*
b11 6
19
1>
1C
b11 G
#941760000000
0!
0*
09
0>
0C
#941770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#941780000000
0!
0*
09
0>
0C
#941790000000
1!
1*
b101 6
19
1>
1C
b101 G
#941800000000
0!
0*
09
0>
0C
#941810000000
1!
1*
b110 6
19
1>
1C
b110 G
#941820000000
0!
0*
09
0>
0C
#941830000000
1!
1*
b111 6
19
1>
1C
b111 G
#941840000000
0!
1"
0*
1+
09
1:
0>
0C
#941850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#941860000000
0!
0*
09
0>
0C
#941870000000
1!
1*
b1 6
19
1>
1C
b1 G
#941880000000
0!
0*
09
0>
0C
#941890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#941900000000
0!
0*
09
0>
0C
#941910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#941920000000
0!
0*
09
0>
0C
#941930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#941940000000
0!
0*
09
0>
0C
#941950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#941960000000
0!
0#
0*
0,
09
0>
0?
0C
#941970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#941980000000
0!
0*
09
0>
0C
#941990000000
1!
1*
19
1>
1C
#942000000000
0!
0*
09
0>
0C
#942010000000
1!
1*
19
1>
1C
#942020000000
0!
0*
09
0>
0C
#942030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#942040000000
0!
0*
09
0>
0C
#942050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#942060000000
0!
0*
09
0>
0C
#942070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#942080000000
0!
0*
09
0>
0C
#942090000000
1!
1*
b10 6
19
1>
1C
b10 G
#942100000000
0!
0*
09
0>
0C
#942110000000
1!
1*
b11 6
19
1>
1C
b11 G
#942120000000
0!
0*
09
0>
0C
#942130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#942140000000
0!
0*
09
0>
0C
#942150000000
1!
1*
b101 6
19
1>
1C
b101 G
#942160000000
0!
0*
09
0>
0C
#942170000000
1!
1*
b110 6
19
1>
1C
b110 G
#942180000000
0!
0*
09
0>
0C
#942190000000
1!
1*
b111 6
19
1>
1C
b111 G
#942200000000
0!
0*
09
0>
0C
#942210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#942220000000
0!
0*
09
0>
0C
#942230000000
1!
1*
b1 6
19
1>
1C
b1 G
#942240000000
0!
0*
09
0>
0C
#942250000000
1!
1*
b10 6
19
1>
1C
b10 G
#942260000000
0!
0*
09
0>
0C
#942270000000
1!
1*
b11 6
19
1>
1C
b11 G
#942280000000
0!
0*
09
0>
0C
#942290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#942300000000
0!
0*
09
0>
0C
#942310000000
1!
1*
b101 6
19
1>
1C
b101 G
#942320000000
0!
0*
09
0>
0C
#942330000000
1!
1*
b110 6
19
1>
1C
b110 G
#942340000000
0!
0*
09
0>
0C
#942350000000
1!
1*
b111 6
19
1>
1C
b111 G
#942360000000
0!
0*
09
0>
0C
#942370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#942380000000
0!
0*
09
0>
0C
#942390000000
1!
1*
b1 6
19
1>
1C
b1 G
#942400000000
0!
0*
09
0>
0C
#942410000000
1!
1*
b10 6
19
1>
1C
b10 G
#942420000000
0!
0*
09
0>
0C
#942430000000
1!
1*
b11 6
19
1>
1C
b11 G
#942440000000
0!
0*
09
0>
0C
#942450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#942460000000
0!
0*
09
0>
0C
#942470000000
1!
1*
b101 6
19
1>
1C
b101 G
#942480000000
0!
0*
09
0>
0C
#942490000000
1!
1*
b110 6
19
1>
1C
b110 G
#942500000000
0!
0*
09
0>
0C
#942510000000
1!
1*
b111 6
19
1>
1C
b111 G
#942520000000
0!
1"
0*
1+
09
1:
0>
0C
#942530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#942540000000
0!
0*
09
0>
0C
#942550000000
1!
1*
b1 6
19
1>
1C
b1 G
#942560000000
0!
0*
09
0>
0C
#942570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#942580000000
0!
0*
09
0>
0C
#942590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#942600000000
0!
0*
09
0>
0C
#942610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#942620000000
0!
0*
09
0>
0C
#942630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#942640000000
0!
0#
0*
0,
09
0>
0?
0C
#942650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#942660000000
0!
0*
09
0>
0C
#942670000000
1!
1*
19
1>
1C
#942680000000
0!
0*
09
0>
0C
#942690000000
1!
1*
19
1>
1C
#942700000000
0!
0*
09
0>
0C
#942710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#942720000000
0!
0*
09
0>
0C
#942730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#942740000000
0!
0*
09
0>
0C
#942750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#942760000000
0!
0*
09
0>
0C
#942770000000
1!
1*
b10 6
19
1>
1C
b10 G
#942780000000
0!
0*
09
0>
0C
#942790000000
1!
1*
b11 6
19
1>
1C
b11 G
#942800000000
0!
0*
09
0>
0C
#942810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#942820000000
0!
0*
09
0>
0C
#942830000000
1!
1*
b101 6
19
1>
1C
b101 G
#942840000000
0!
0*
09
0>
0C
#942850000000
1!
1*
b110 6
19
1>
1C
b110 G
#942860000000
0!
0*
09
0>
0C
#942870000000
1!
1*
b111 6
19
1>
1C
b111 G
#942880000000
0!
0*
09
0>
0C
#942890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#942900000000
0!
0*
09
0>
0C
#942910000000
1!
1*
b1 6
19
1>
1C
b1 G
#942920000000
0!
0*
09
0>
0C
#942930000000
1!
1*
b10 6
19
1>
1C
b10 G
#942940000000
0!
0*
09
0>
0C
#942950000000
1!
1*
b11 6
19
1>
1C
b11 G
#942960000000
0!
0*
09
0>
0C
#942970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#942980000000
0!
0*
09
0>
0C
#942990000000
1!
1*
b101 6
19
1>
1C
b101 G
#943000000000
0!
0*
09
0>
0C
#943010000000
1!
1*
b110 6
19
1>
1C
b110 G
#943020000000
0!
0*
09
0>
0C
#943030000000
1!
1*
b111 6
19
1>
1C
b111 G
#943040000000
0!
0*
09
0>
0C
#943050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#943060000000
0!
0*
09
0>
0C
#943070000000
1!
1*
b1 6
19
1>
1C
b1 G
#943080000000
0!
0*
09
0>
0C
#943090000000
1!
1*
b10 6
19
1>
1C
b10 G
#943100000000
0!
0*
09
0>
0C
#943110000000
1!
1*
b11 6
19
1>
1C
b11 G
#943120000000
0!
0*
09
0>
0C
#943130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#943140000000
0!
0*
09
0>
0C
#943150000000
1!
1*
b101 6
19
1>
1C
b101 G
#943160000000
0!
0*
09
0>
0C
#943170000000
1!
1*
b110 6
19
1>
1C
b110 G
#943180000000
0!
0*
09
0>
0C
#943190000000
1!
1*
b111 6
19
1>
1C
b111 G
#943200000000
0!
1"
0*
1+
09
1:
0>
0C
#943210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#943220000000
0!
0*
09
0>
0C
#943230000000
1!
1*
b1 6
19
1>
1C
b1 G
#943240000000
0!
0*
09
0>
0C
#943250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#943260000000
0!
0*
09
0>
0C
#943270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#943280000000
0!
0*
09
0>
0C
#943290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#943300000000
0!
0*
09
0>
0C
#943310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#943320000000
0!
0#
0*
0,
09
0>
0?
0C
#943330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#943340000000
0!
0*
09
0>
0C
#943350000000
1!
1*
19
1>
1C
#943360000000
0!
0*
09
0>
0C
#943370000000
1!
1*
19
1>
1C
#943380000000
0!
0*
09
0>
0C
#943390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#943400000000
0!
0*
09
0>
0C
#943410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#943420000000
0!
0*
09
0>
0C
#943430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#943440000000
0!
0*
09
0>
0C
#943450000000
1!
1*
b10 6
19
1>
1C
b10 G
#943460000000
0!
0*
09
0>
0C
#943470000000
1!
1*
b11 6
19
1>
1C
b11 G
#943480000000
0!
0*
09
0>
0C
#943490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#943500000000
0!
0*
09
0>
0C
#943510000000
1!
1*
b101 6
19
1>
1C
b101 G
#943520000000
0!
0*
09
0>
0C
#943530000000
1!
1*
b110 6
19
1>
1C
b110 G
#943540000000
0!
0*
09
0>
0C
#943550000000
1!
1*
b111 6
19
1>
1C
b111 G
#943560000000
0!
0*
09
0>
0C
#943570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#943580000000
0!
0*
09
0>
0C
#943590000000
1!
1*
b1 6
19
1>
1C
b1 G
#943600000000
0!
0*
09
0>
0C
#943610000000
1!
1*
b10 6
19
1>
1C
b10 G
#943620000000
0!
0*
09
0>
0C
#943630000000
1!
1*
b11 6
19
1>
1C
b11 G
#943640000000
0!
0*
09
0>
0C
#943650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#943660000000
0!
0*
09
0>
0C
#943670000000
1!
1*
b101 6
19
1>
1C
b101 G
#943680000000
0!
0*
09
0>
0C
#943690000000
1!
1*
b110 6
19
1>
1C
b110 G
#943700000000
0!
0*
09
0>
0C
#943710000000
1!
1*
b111 6
19
1>
1C
b111 G
#943720000000
0!
0*
09
0>
0C
#943730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#943740000000
0!
0*
09
0>
0C
#943750000000
1!
1*
b1 6
19
1>
1C
b1 G
#943760000000
0!
0*
09
0>
0C
#943770000000
1!
1*
b10 6
19
1>
1C
b10 G
#943780000000
0!
0*
09
0>
0C
#943790000000
1!
1*
b11 6
19
1>
1C
b11 G
#943800000000
0!
0*
09
0>
0C
#943810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#943820000000
0!
0*
09
0>
0C
#943830000000
1!
1*
b101 6
19
1>
1C
b101 G
#943840000000
0!
0*
09
0>
0C
#943850000000
1!
1*
b110 6
19
1>
1C
b110 G
#943860000000
0!
0*
09
0>
0C
#943870000000
1!
1*
b111 6
19
1>
1C
b111 G
#943880000000
0!
1"
0*
1+
09
1:
0>
0C
#943890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#943900000000
0!
0*
09
0>
0C
#943910000000
1!
1*
b1 6
19
1>
1C
b1 G
#943920000000
0!
0*
09
0>
0C
#943930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#943940000000
0!
0*
09
0>
0C
#943950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#943960000000
0!
0*
09
0>
0C
#943970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#943980000000
0!
0*
09
0>
0C
#943990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#944000000000
0!
0#
0*
0,
09
0>
0?
0C
#944010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#944020000000
0!
0*
09
0>
0C
#944030000000
1!
1*
19
1>
1C
#944040000000
0!
0*
09
0>
0C
#944050000000
1!
1*
19
1>
1C
#944060000000
0!
0*
09
0>
0C
#944070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#944080000000
0!
0*
09
0>
0C
#944090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#944100000000
0!
0*
09
0>
0C
#944110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#944120000000
0!
0*
09
0>
0C
#944130000000
1!
1*
b10 6
19
1>
1C
b10 G
#944140000000
0!
0*
09
0>
0C
#944150000000
1!
1*
b11 6
19
1>
1C
b11 G
#944160000000
0!
0*
09
0>
0C
#944170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#944180000000
0!
0*
09
0>
0C
#944190000000
1!
1*
b101 6
19
1>
1C
b101 G
#944200000000
0!
0*
09
0>
0C
#944210000000
1!
1*
b110 6
19
1>
1C
b110 G
#944220000000
0!
0*
09
0>
0C
#944230000000
1!
1*
b111 6
19
1>
1C
b111 G
#944240000000
0!
0*
09
0>
0C
#944250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#944260000000
0!
0*
09
0>
0C
#944270000000
1!
1*
b1 6
19
1>
1C
b1 G
#944280000000
0!
0*
09
0>
0C
#944290000000
1!
1*
b10 6
19
1>
1C
b10 G
#944300000000
0!
0*
09
0>
0C
#944310000000
1!
1*
b11 6
19
1>
1C
b11 G
#944320000000
0!
0*
09
0>
0C
#944330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#944340000000
0!
0*
09
0>
0C
#944350000000
1!
1*
b101 6
19
1>
1C
b101 G
#944360000000
0!
0*
09
0>
0C
#944370000000
1!
1*
b110 6
19
1>
1C
b110 G
#944380000000
0!
0*
09
0>
0C
#944390000000
1!
1*
b111 6
19
1>
1C
b111 G
#944400000000
0!
0*
09
0>
0C
#944410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#944420000000
0!
0*
09
0>
0C
#944430000000
1!
1*
b1 6
19
1>
1C
b1 G
#944440000000
0!
0*
09
0>
0C
#944450000000
1!
1*
b10 6
19
1>
1C
b10 G
#944460000000
0!
0*
09
0>
0C
#944470000000
1!
1*
b11 6
19
1>
1C
b11 G
#944480000000
0!
0*
09
0>
0C
#944490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#944500000000
0!
0*
09
0>
0C
#944510000000
1!
1*
b101 6
19
1>
1C
b101 G
#944520000000
0!
0*
09
0>
0C
#944530000000
1!
1*
b110 6
19
1>
1C
b110 G
#944540000000
0!
0*
09
0>
0C
#944550000000
1!
1*
b111 6
19
1>
1C
b111 G
#944560000000
0!
1"
0*
1+
09
1:
0>
0C
#944570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#944580000000
0!
0*
09
0>
0C
#944590000000
1!
1*
b1 6
19
1>
1C
b1 G
#944600000000
0!
0*
09
0>
0C
#944610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#944620000000
0!
0*
09
0>
0C
#944630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#944640000000
0!
0*
09
0>
0C
#944650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#944660000000
0!
0*
09
0>
0C
#944670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#944680000000
0!
0#
0*
0,
09
0>
0?
0C
#944690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#944700000000
0!
0*
09
0>
0C
#944710000000
1!
1*
19
1>
1C
#944720000000
0!
0*
09
0>
0C
#944730000000
1!
1*
19
1>
1C
#944740000000
0!
0*
09
0>
0C
#944750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#944760000000
0!
0*
09
0>
0C
#944770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#944780000000
0!
0*
09
0>
0C
#944790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#944800000000
0!
0*
09
0>
0C
#944810000000
1!
1*
b10 6
19
1>
1C
b10 G
#944820000000
0!
0*
09
0>
0C
#944830000000
1!
1*
b11 6
19
1>
1C
b11 G
#944840000000
0!
0*
09
0>
0C
#944850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#944860000000
0!
0*
09
0>
0C
#944870000000
1!
1*
b101 6
19
1>
1C
b101 G
#944880000000
0!
0*
09
0>
0C
#944890000000
1!
1*
b110 6
19
1>
1C
b110 G
#944900000000
0!
0*
09
0>
0C
#944910000000
1!
1*
b111 6
19
1>
1C
b111 G
#944920000000
0!
0*
09
0>
0C
#944930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#944940000000
0!
0*
09
0>
0C
#944950000000
1!
1*
b1 6
19
1>
1C
b1 G
#944960000000
0!
0*
09
0>
0C
#944970000000
1!
1*
b10 6
19
1>
1C
b10 G
#944980000000
0!
0*
09
0>
0C
#944990000000
1!
1*
b11 6
19
1>
1C
b11 G
#945000000000
0!
0*
09
0>
0C
#945010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#945020000000
0!
0*
09
0>
0C
#945030000000
1!
1*
b101 6
19
1>
1C
b101 G
#945040000000
0!
0*
09
0>
0C
#945050000000
1!
1*
b110 6
19
1>
1C
b110 G
#945060000000
0!
0*
09
0>
0C
#945070000000
1!
1*
b111 6
19
1>
1C
b111 G
#945080000000
0!
0*
09
0>
0C
#945090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#945100000000
0!
0*
09
0>
0C
#945110000000
1!
1*
b1 6
19
1>
1C
b1 G
#945120000000
0!
0*
09
0>
0C
#945130000000
1!
1*
b10 6
19
1>
1C
b10 G
#945140000000
0!
0*
09
0>
0C
#945150000000
1!
1*
b11 6
19
1>
1C
b11 G
#945160000000
0!
0*
09
0>
0C
#945170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#945180000000
0!
0*
09
0>
0C
#945190000000
1!
1*
b101 6
19
1>
1C
b101 G
#945200000000
0!
0*
09
0>
0C
#945210000000
1!
1*
b110 6
19
1>
1C
b110 G
#945220000000
0!
0*
09
0>
0C
#945230000000
1!
1*
b111 6
19
1>
1C
b111 G
#945240000000
0!
1"
0*
1+
09
1:
0>
0C
#945250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#945260000000
0!
0*
09
0>
0C
#945270000000
1!
1*
b1 6
19
1>
1C
b1 G
#945280000000
0!
0*
09
0>
0C
#945290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#945300000000
0!
0*
09
0>
0C
#945310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#945320000000
0!
0*
09
0>
0C
#945330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#945340000000
0!
0*
09
0>
0C
#945350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#945360000000
0!
0#
0*
0,
09
0>
0?
0C
#945370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#945380000000
0!
0*
09
0>
0C
#945390000000
1!
1*
19
1>
1C
#945400000000
0!
0*
09
0>
0C
#945410000000
1!
1*
19
1>
1C
#945420000000
0!
0*
09
0>
0C
#945430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#945440000000
0!
0*
09
0>
0C
#945450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#945460000000
0!
0*
09
0>
0C
#945470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#945480000000
0!
0*
09
0>
0C
#945490000000
1!
1*
b10 6
19
1>
1C
b10 G
#945500000000
0!
0*
09
0>
0C
#945510000000
1!
1*
b11 6
19
1>
1C
b11 G
#945520000000
0!
0*
09
0>
0C
#945530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#945540000000
0!
0*
09
0>
0C
#945550000000
1!
1*
b101 6
19
1>
1C
b101 G
#945560000000
0!
0*
09
0>
0C
#945570000000
1!
1*
b110 6
19
1>
1C
b110 G
#945580000000
0!
0*
09
0>
0C
#945590000000
1!
1*
b111 6
19
1>
1C
b111 G
#945600000000
0!
0*
09
0>
0C
#945610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#945620000000
0!
0*
09
0>
0C
#945630000000
1!
1*
b1 6
19
1>
1C
b1 G
#945640000000
0!
0*
09
0>
0C
#945650000000
1!
1*
b10 6
19
1>
1C
b10 G
#945660000000
0!
0*
09
0>
0C
#945670000000
1!
1*
b11 6
19
1>
1C
b11 G
#945680000000
0!
0*
09
0>
0C
#945690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#945700000000
0!
0*
09
0>
0C
#945710000000
1!
1*
b101 6
19
1>
1C
b101 G
#945720000000
0!
0*
09
0>
0C
#945730000000
1!
1*
b110 6
19
1>
1C
b110 G
#945740000000
0!
0*
09
0>
0C
#945750000000
1!
1*
b111 6
19
1>
1C
b111 G
#945760000000
0!
0*
09
0>
0C
#945770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#945780000000
0!
0*
09
0>
0C
#945790000000
1!
1*
b1 6
19
1>
1C
b1 G
#945800000000
0!
0*
09
0>
0C
#945810000000
1!
1*
b10 6
19
1>
1C
b10 G
#945820000000
0!
0*
09
0>
0C
#945830000000
1!
1*
b11 6
19
1>
1C
b11 G
#945840000000
0!
0*
09
0>
0C
#945850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#945860000000
0!
0*
09
0>
0C
#945870000000
1!
1*
b101 6
19
1>
1C
b101 G
#945880000000
0!
0*
09
0>
0C
#945890000000
1!
1*
b110 6
19
1>
1C
b110 G
#945900000000
0!
0*
09
0>
0C
#945910000000
1!
1*
b111 6
19
1>
1C
b111 G
#945920000000
0!
1"
0*
1+
09
1:
0>
0C
#945930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#945940000000
0!
0*
09
0>
0C
#945950000000
1!
1*
b1 6
19
1>
1C
b1 G
#945960000000
0!
0*
09
0>
0C
#945970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#945980000000
0!
0*
09
0>
0C
#945990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#946000000000
0!
0*
09
0>
0C
#946010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#946020000000
0!
0*
09
0>
0C
#946030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#946040000000
0!
0#
0*
0,
09
0>
0?
0C
#946050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#946060000000
0!
0*
09
0>
0C
#946070000000
1!
1*
19
1>
1C
#946080000000
0!
0*
09
0>
0C
#946090000000
1!
1*
19
1>
1C
#946100000000
0!
0*
09
0>
0C
#946110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#946120000000
0!
0*
09
0>
0C
#946130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#946140000000
0!
0*
09
0>
0C
#946150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#946160000000
0!
0*
09
0>
0C
#946170000000
1!
1*
b10 6
19
1>
1C
b10 G
#946180000000
0!
0*
09
0>
0C
#946190000000
1!
1*
b11 6
19
1>
1C
b11 G
#946200000000
0!
0*
09
0>
0C
#946210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#946220000000
0!
0*
09
0>
0C
#946230000000
1!
1*
b101 6
19
1>
1C
b101 G
#946240000000
0!
0*
09
0>
0C
#946250000000
1!
1*
b110 6
19
1>
1C
b110 G
#946260000000
0!
0*
09
0>
0C
#946270000000
1!
1*
b111 6
19
1>
1C
b111 G
#946280000000
0!
0*
09
0>
0C
#946290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#946300000000
0!
0*
09
0>
0C
#946310000000
1!
1*
b1 6
19
1>
1C
b1 G
#946320000000
0!
0*
09
0>
0C
#946330000000
1!
1*
b10 6
19
1>
1C
b10 G
#946340000000
0!
0*
09
0>
0C
#946350000000
1!
1*
b11 6
19
1>
1C
b11 G
#946360000000
0!
0*
09
0>
0C
#946370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#946380000000
0!
0*
09
0>
0C
#946390000000
1!
1*
b101 6
19
1>
1C
b101 G
#946400000000
0!
0*
09
0>
0C
#946410000000
1!
1*
b110 6
19
1>
1C
b110 G
#946420000000
0!
0*
09
0>
0C
#946430000000
1!
1*
b111 6
19
1>
1C
b111 G
#946440000000
0!
0*
09
0>
0C
#946450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#946460000000
0!
0*
09
0>
0C
#946470000000
1!
1*
b1 6
19
1>
1C
b1 G
#946480000000
0!
0*
09
0>
0C
#946490000000
1!
1*
b10 6
19
1>
1C
b10 G
#946500000000
0!
0*
09
0>
0C
#946510000000
1!
1*
b11 6
19
1>
1C
b11 G
#946520000000
0!
0*
09
0>
0C
#946530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#946540000000
0!
0*
09
0>
0C
#946550000000
1!
1*
b101 6
19
1>
1C
b101 G
#946560000000
0!
0*
09
0>
0C
#946570000000
1!
1*
b110 6
19
1>
1C
b110 G
#946580000000
0!
0*
09
0>
0C
#946590000000
1!
1*
b111 6
19
1>
1C
b111 G
#946600000000
0!
1"
0*
1+
09
1:
0>
0C
#946610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#946620000000
0!
0*
09
0>
0C
#946630000000
1!
1*
b1 6
19
1>
1C
b1 G
#946640000000
0!
0*
09
0>
0C
#946650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#946660000000
0!
0*
09
0>
0C
#946670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#946680000000
0!
0*
09
0>
0C
#946690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#946700000000
0!
0*
09
0>
0C
#946710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#946720000000
0!
0#
0*
0,
09
0>
0?
0C
#946730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#946740000000
0!
0*
09
0>
0C
#946750000000
1!
1*
19
1>
1C
#946760000000
0!
0*
09
0>
0C
#946770000000
1!
1*
19
1>
1C
#946780000000
0!
0*
09
0>
0C
#946790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#946800000000
0!
0*
09
0>
0C
#946810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#946820000000
0!
0*
09
0>
0C
#946830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#946840000000
0!
0*
09
0>
0C
#946850000000
1!
1*
b10 6
19
1>
1C
b10 G
#946860000000
0!
0*
09
0>
0C
#946870000000
1!
1*
b11 6
19
1>
1C
b11 G
#946880000000
0!
0*
09
0>
0C
#946890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#946900000000
0!
0*
09
0>
0C
#946910000000
1!
1*
b101 6
19
1>
1C
b101 G
#946920000000
0!
0*
09
0>
0C
#946930000000
1!
1*
b110 6
19
1>
1C
b110 G
#946940000000
0!
0*
09
0>
0C
#946950000000
1!
1*
b111 6
19
1>
1C
b111 G
#946960000000
0!
0*
09
0>
0C
#946970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#946980000000
0!
0*
09
0>
0C
#946990000000
1!
1*
b1 6
19
1>
1C
b1 G
#947000000000
0!
0*
09
0>
0C
#947010000000
1!
1*
b10 6
19
1>
1C
b10 G
#947020000000
0!
0*
09
0>
0C
#947030000000
1!
1*
b11 6
19
1>
1C
b11 G
#947040000000
0!
0*
09
0>
0C
#947050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#947060000000
0!
0*
09
0>
0C
#947070000000
1!
1*
b101 6
19
1>
1C
b101 G
#947080000000
0!
0*
09
0>
0C
#947090000000
1!
1*
b110 6
19
1>
1C
b110 G
#947100000000
0!
0*
09
0>
0C
#947110000000
1!
1*
b111 6
19
1>
1C
b111 G
#947120000000
0!
0*
09
0>
0C
#947130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#947140000000
0!
0*
09
0>
0C
#947150000000
1!
1*
b1 6
19
1>
1C
b1 G
#947160000000
0!
0*
09
0>
0C
#947170000000
1!
1*
b10 6
19
1>
1C
b10 G
#947180000000
0!
0*
09
0>
0C
#947190000000
1!
1*
b11 6
19
1>
1C
b11 G
#947200000000
0!
0*
09
0>
0C
#947210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#947220000000
0!
0*
09
0>
0C
#947230000000
1!
1*
b101 6
19
1>
1C
b101 G
#947240000000
0!
0*
09
0>
0C
#947250000000
1!
1*
b110 6
19
1>
1C
b110 G
#947260000000
0!
0*
09
0>
0C
#947270000000
1!
1*
b111 6
19
1>
1C
b111 G
#947280000000
0!
1"
0*
1+
09
1:
0>
0C
#947290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#947300000000
0!
0*
09
0>
0C
#947310000000
1!
1*
b1 6
19
1>
1C
b1 G
#947320000000
0!
0*
09
0>
0C
#947330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#947340000000
0!
0*
09
0>
0C
#947350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#947360000000
0!
0*
09
0>
0C
#947370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#947380000000
0!
0*
09
0>
0C
#947390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#947400000000
0!
0#
0*
0,
09
0>
0?
0C
#947410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#947420000000
0!
0*
09
0>
0C
#947430000000
1!
1*
19
1>
1C
#947440000000
0!
0*
09
0>
0C
#947450000000
1!
1*
19
1>
1C
#947460000000
0!
0*
09
0>
0C
#947470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#947480000000
0!
0*
09
0>
0C
#947490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#947500000000
0!
0*
09
0>
0C
#947510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#947520000000
0!
0*
09
0>
0C
#947530000000
1!
1*
b10 6
19
1>
1C
b10 G
#947540000000
0!
0*
09
0>
0C
#947550000000
1!
1*
b11 6
19
1>
1C
b11 G
#947560000000
0!
0*
09
0>
0C
#947570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#947580000000
0!
0*
09
0>
0C
#947590000000
1!
1*
b101 6
19
1>
1C
b101 G
#947600000000
0!
0*
09
0>
0C
#947610000000
1!
1*
b110 6
19
1>
1C
b110 G
#947620000000
0!
0*
09
0>
0C
#947630000000
1!
1*
b111 6
19
1>
1C
b111 G
#947640000000
0!
0*
09
0>
0C
#947650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#947660000000
0!
0*
09
0>
0C
#947670000000
1!
1*
b1 6
19
1>
1C
b1 G
#947680000000
0!
0*
09
0>
0C
#947690000000
1!
1*
b10 6
19
1>
1C
b10 G
#947700000000
0!
0*
09
0>
0C
#947710000000
1!
1*
b11 6
19
1>
1C
b11 G
#947720000000
0!
0*
09
0>
0C
#947730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#947740000000
0!
0*
09
0>
0C
#947750000000
1!
1*
b101 6
19
1>
1C
b101 G
#947760000000
0!
0*
09
0>
0C
#947770000000
1!
1*
b110 6
19
1>
1C
b110 G
#947780000000
0!
0*
09
0>
0C
#947790000000
1!
1*
b111 6
19
1>
1C
b111 G
#947800000000
0!
0*
09
0>
0C
#947810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#947820000000
0!
0*
09
0>
0C
#947830000000
1!
1*
b1 6
19
1>
1C
b1 G
#947840000000
0!
0*
09
0>
0C
#947850000000
1!
1*
b10 6
19
1>
1C
b10 G
#947860000000
0!
0*
09
0>
0C
#947870000000
1!
1*
b11 6
19
1>
1C
b11 G
#947880000000
0!
0*
09
0>
0C
#947890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#947900000000
0!
0*
09
0>
0C
#947910000000
1!
1*
b101 6
19
1>
1C
b101 G
#947920000000
0!
0*
09
0>
0C
#947930000000
1!
1*
b110 6
19
1>
1C
b110 G
#947940000000
0!
0*
09
0>
0C
#947950000000
1!
1*
b111 6
19
1>
1C
b111 G
#947960000000
0!
1"
0*
1+
09
1:
0>
0C
#947970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#947980000000
0!
0*
09
0>
0C
#947990000000
1!
1*
b1 6
19
1>
1C
b1 G
#948000000000
0!
0*
09
0>
0C
#948010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#948020000000
0!
0*
09
0>
0C
#948030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#948040000000
0!
0*
09
0>
0C
#948050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#948060000000
0!
0*
09
0>
0C
#948070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#948080000000
0!
0#
0*
0,
09
0>
0?
0C
#948090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#948100000000
0!
0*
09
0>
0C
#948110000000
1!
1*
19
1>
1C
#948120000000
0!
0*
09
0>
0C
#948130000000
1!
1*
19
1>
1C
#948140000000
0!
0*
09
0>
0C
#948150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#948160000000
0!
0*
09
0>
0C
#948170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#948180000000
0!
0*
09
0>
0C
#948190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#948200000000
0!
0*
09
0>
0C
#948210000000
1!
1*
b10 6
19
1>
1C
b10 G
#948220000000
0!
0*
09
0>
0C
#948230000000
1!
1*
b11 6
19
1>
1C
b11 G
#948240000000
0!
0*
09
0>
0C
#948250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#948260000000
0!
0*
09
0>
0C
#948270000000
1!
1*
b101 6
19
1>
1C
b101 G
#948280000000
0!
0*
09
0>
0C
#948290000000
1!
1*
b110 6
19
1>
1C
b110 G
#948300000000
0!
0*
09
0>
0C
#948310000000
1!
1*
b111 6
19
1>
1C
b111 G
#948320000000
0!
0*
09
0>
0C
#948330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#948340000000
0!
0*
09
0>
0C
#948350000000
1!
1*
b1 6
19
1>
1C
b1 G
#948360000000
0!
0*
09
0>
0C
#948370000000
1!
1*
b10 6
19
1>
1C
b10 G
#948380000000
0!
0*
09
0>
0C
#948390000000
1!
1*
b11 6
19
1>
1C
b11 G
#948400000000
0!
0*
09
0>
0C
#948410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#948420000000
0!
0*
09
0>
0C
#948430000000
1!
1*
b101 6
19
1>
1C
b101 G
#948440000000
0!
0*
09
0>
0C
#948450000000
1!
1*
b110 6
19
1>
1C
b110 G
#948460000000
0!
0*
09
0>
0C
#948470000000
1!
1*
b111 6
19
1>
1C
b111 G
#948480000000
0!
0*
09
0>
0C
#948490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#948500000000
0!
0*
09
0>
0C
#948510000000
1!
1*
b1 6
19
1>
1C
b1 G
#948520000000
0!
0*
09
0>
0C
#948530000000
1!
1*
b10 6
19
1>
1C
b10 G
#948540000000
0!
0*
09
0>
0C
#948550000000
1!
1*
b11 6
19
1>
1C
b11 G
#948560000000
0!
0*
09
0>
0C
#948570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#948580000000
0!
0*
09
0>
0C
#948590000000
1!
1*
b101 6
19
1>
1C
b101 G
#948600000000
0!
0*
09
0>
0C
#948610000000
1!
1*
b110 6
19
1>
1C
b110 G
#948620000000
0!
0*
09
0>
0C
#948630000000
1!
1*
b111 6
19
1>
1C
b111 G
#948640000000
0!
1"
0*
1+
09
1:
0>
0C
#948650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#948660000000
0!
0*
09
0>
0C
#948670000000
1!
1*
b1 6
19
1>
1C
b1 G
#948680000000
0!
0*
09
0>
0C
#948690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#948700000000
0!
0*
09
0>
0C
#948710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#948720000000
0!
0*
09
0>
0C
#948730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#948740000000
0!
0*
09
0>
0C
#948750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#948760000000
0!
0#
0*
0,
09
0>
0?
0C
#948770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#948780000000
0!
0*
09
0>
0C
#948790000000
1!
1*
19
1>
1C
#948800000000
0!
0*
09
0>
0C
#948810000000
1!
1*
19
1>
1C
#948820000000
0!
0*
09
0>
0C
#948830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#948840000000
0!
0*
09
0>
0C
#948850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#948860000000
0!
0*
09
0>
0C
#948870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#948880000000
0!
0*
09
0>
0C
#948890000000
1!
1*
b10 6
19
1>
1C
b10 G
#948900000000
0!
0*
09
0>
0C
#948910000000
1!
1*
b11 6
19
1>
1C
b11 G
#948920000000
0!
0*
09
0>
0C
#948930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#948940000000
0!
0*
09
0>
0C
#948950000000
1!
1*
b101 6
19
1>
1C
b101 G
#948960000000
0!
0*
09
0>
0C
#948970000000
1!
1*
b110 6
19
1>
1C
b110 G
#948980000000
0!
0*
09
0>
0C
#948990000000
1!
1*
b111 6
19
1>
1C
b111 G
#949000000000
0!
0*
09
0>
0C
#949010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#949020000000
0!
0*
09
0>
0C
#949030000000
1!
1*
b1 6
19
1>
1C
b1 G
#949040000000
0!
0*
09
0>
0C
#949050000000
1!
1*
b10 6
19
1>
1C
b10 G
#949060000000
0!
0*
09
0>
0C
#949070000000
1!
1*
b11 6
19
1>
1C
b11 G
#949080000000
0!
0*
09
0>
0C
#949090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#949100000000
0!
0*
09
0>
0C
#949110000000
1!
1*
b101 6
19
1>
1C
b101 G
#949120000000
0!
0*
09
0>
0C
#949130000000
1!
1*
b110 6
19
1>
1C
b110 G
#949140000000
0!
0*
09
0>
0C
#949150000000
1!
1*
b111 6
19
1>
1C
b111 G
#949160000000
0!
0*
09
0>
0C
#949170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#949180000000
0!
0*
09
0>
0C
#949190000000
1!
1*
b1 6
19
1>
1C
b1 G
#949200000000
0!
0*
09
0>
0C
#949210000000
1!
1*
b10 6
19
1>
1C
b10 G
#949220000000
0!
0*
09
0>
0C
#949230000000
1!
1*
b11 6
19
1>
1C
b11 G
#949240000000
0!
0*
09
0>
0C
#949250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#949260000000
0!
0*
09
0>
0C
#949270000000
1!
1*
b101 6
19
1>
1C
b101 G
#949280000000
0!
0*
09
0>
0C
#949290000000
1!
1*
b110 6
19
1>
1C
b110 G
#949300000000
0!
0*
09
0>
0C
#949310000000
1!
1*
b111 6
19
1>
1C
b111 G
#949320000000
0!
1"
0*
1+
09
1:
0>
0C
#949330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#949340000000
0!
0*
09
0>
0C
#949350000000
1!
1*
b1 6
19
1>
1C
b1 G
#949360000000
0!
0*
09
0>
0C
#949370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#949380000000
0!
0*
09
0>
0C
#949390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#949400000000
0!
0*
09
0>
0C
#949410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#949420000000
0!
0*
09
0>
0C
#949430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#949440000000
0!
0#
0*
0,
09
0>
0?
0C
#949450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#949460000000
0!
0*
09
0>
0C
#949470000000
1!
1*
19
1>
1C
#949480000000
0!
0*
09
0>
0C
#949490000000
1!
1*
19
1>
1C
#949500000000
0!
0*
09
0>
0C
#949510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#949520000000
0!
0*
09
0>
0C
#949530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#949540000000
0!
0*
09
0>
0C
#949550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#949560000000
0!
0*
09
0>
0C
#949570000000
1!
1*
b10 6
19
1>
1C
b10 G
#949580000000
0!
0*
09
0>
0C
#949590000000
1!
1*
b11 6
19
1>
1C
b11 G
#949600000000
0!
0*
09
0>
0C
#949610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#949620000000
0!
0*
09
0>
0C
#949630000000
1!
1*
b101 6
19
1>
1C
b101 G
#949640000000
0!
0*
09
0>
0C
#949650000000
1!
1*
b110 6
19
1>
1C
b110 G
#949660000000
0!
0*
09
0>
0C
#949670000000
1!
1*
b111 6
19
1>
1C
b111 G
#949680000000
0!
0*
09
0>
0C
#949690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#949700000000
0!
0*
09
0>
0C
#949710000000
1!
1*
b1 6
19
1>
1C
b1 G
#949720000000
0!
0*
09
0>
0C
#949730000000
1!
1*
b10 6
19
1>
1C
b10 G
#949740000000
0!
0*
09
0>
0C
#949750000000
1!
1*
b11 6
19
1>
1C
b11 G
#949760000000
0!
0*
09
0>
0C
#949770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#949780000000
0!
0*
09
0>
0C
#949790000000
1!
1*
b101 6
19
1>
1C
b101 G
#949800000000
0!
0*
09
0>
0C
#949810000000
1!
1*
b110 6
19
1>
1C
b110 G
#949820000000
0!
0*
09
0>
0C
#949830000000
1!
1*
b111 6
19
1>
1C
b111 G
#949840000000
0!
0*
09
0>
0C
#949850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#949860000000
0!
0*
09
0>
0C
#949870000000
1!
1*
b1 6
19
1>
1C
b1 G
#949880000000
0!
0*
09
0>
0C
#949890000000
1!
1*
b10 6
19
1>
1C
b10 G
#949900000000
0!
0*
09
0>
0C
#949910000000
1!
1*
b11 6
19
1>
1C
b11 G
#949920000000
0!
0*
09
0>
0C
#949930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#949940000000
0!
0*
09
0>
0C
#949950000000
1!
1*
b101 6
19
1>
1C
b101 G
#949960000000
0!
0*
09
0>
0C
#949970000000
1!
1*
b110 6
19
1>
1C
b110 G
#949980000000
0!
0*
09
0>
0C
#949990000000
1!
1*
b111 6
19
1>
1C
b111 G
#950000000000
0!
1"
0*
1+
09
1:
0>
0C
#950010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#950020000000
0!
0*
09
0>
0C
#950030000000
1!
1*
b1 6
19
1>
1C
b1 G
#950040000000
0!
0*
09
0>
0C
#950050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#950060000000
0!
0*
09
0>
0C
#950070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#950080000000
0!
0*
09
0>
0C
#950090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#950100000000
0!
0*
09
0>
0C
#950110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#950120000000
0!
0#
0*
0,
09
0>
0?
0C
#950130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#950140000000
0!
0*
09
0>
0C
#950150000000
1!
1*
19
1>
1C
#950160000000
0!
0*
09
0>
0C
#950170000000
1!
1*
19
1>
1C
#950180000000
0!
0*
09
0>
0C
#950190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#950200000000
0!
0*
09
0>
0C
#950210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#950220000000
0!
0*
09
0>
0C
#950230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#950240000000
0!
0*
09
0>
0C
#950250000000
1!
1*
b10 6
19
1>
1C
b10 G
#950260000000
0!
0*
09
0>
0C
#950270000000
1!
1*
b11 6
19
1>
1C
b11 G
#950280000000
0!
0*
09
0>
0C
#950290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#950300000000
0!
0*
09
0>
0C
#950310000000
1!
1*
b101 6
19
1>
1C
b101 G
#950320000000
0!
0*
09
0>
0C
#950330000000
1!
1*
b110 6
19
1>
1C
b110 G
#950340000000
0!
0*
09
0>
0C
#950350000000
1!
1*
b111 6
19
1>
1C
b111 G
#950360000000
0!
0*
09
0>
0C
#950370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#950380000000
0!
0*
09
0>
0C
#950390000000
1!
1*
b1 6
19
1>
1C
b1 G
#950400000000
0!
0*
09
0>
0C
#950410000000
1!
1*
b10 6
19
1>
1C
b10 G
#950420000000
0!
0*
09
0>
0C
#950430000000
1!
1*
b11 6
19
1>
1C
b11 G
#950440000000
0!
0*
09
0>
0C
#950450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#950460000000
0!
0*
09
0>
0C
#950470000000
1!
1*
b101 6
19
1>
1C
b101 G
#950480000000
0!
0*
09
0>
0C
#950490000000
1!
1*
b110 6
19
1>
1C
b110 G
#950500000000
0!
0*
09
0>
0C
#950510000000
1!
1*
b111 6
19
1>
1C
b111 G
#950520000000
0!
0*
09
0>
0C
#950530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#950540000000
0!
0*
09
0>
0C
#950550000000
1!
1*
b1 6
19
1>
1C
b1 G
#950560000000
0!
0*
09
0>
0C
#950570000000
1!
1*
b10 6
19
1>
1C
b10 G
#950580000000
0!
0*
09
0>
0C
#950590000000
1!
1*
b11 6
19
1>
1C
b11 G
#950600000000
0!
0*
09
0>
0C
#950610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#950620000000
0!
0*
09
0>
0C
#950630000000
1!
1*
b101 6
19
1>
1C
b101 G
#950640000000
0!
0*
09
0>
0C
#950650000000
1!
1*
b110 6
19
1>
1C
b110 G
#950660000000
0!
0*
09
0>
0C
#950670000000
1!
1*
b111 6
19
1>
1C
b111 G
#950680000000
0!
1"
0*
1+
09
1:
0>
0C
#950690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#950700000000
0!
0*
09
0>
0C
#950710000000
1!
1*
b1 6
19
1>
1C
b1 G
#950720000000
0!
0*
09
0>
0C
#950730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#950740000000
0!
0*
09
0>
0C
#950750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#950760000000
0!
0*
09
0>
0C
#950770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#950780000000
0!
0*
09
0>
0C
#950790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#950800000000
0!
0#
0*
0,
09
0>
0?
0C
#950810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#950820000000
0!
0*
09
0>
0C
#950830000000
1!
1*
19
1>
1C
#950840000000
0!
0*
09
0>
0C
#950850000000
1!
1*
19
1>
1C
#950860000000
0!
0*
09
0>
0C
#950870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#950880000000
0!
0*
09
0>
0C
#950890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#950900000000
0!
0*
09
0>
0C
#950910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#950920000000
0!
0*
09
0>
0C
#950930000000
1!
1*
b10 6
19
1>
1C
b10 G
#950940000000
0!
0*
09
0>
0C
#950950000000
1!
1*
b11 6
19
1>
1C
b11 G
#950960000000
0!
0*
09
0>
0C
#950970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#950980000000
0!
0*
09
0>
0C
#950990000000
1!
1*
b101 6
19
1>
1C
b101 G
#951000000000
0!
0*
09
0>
0C
#951010000000
1!
1*
b110 6
19
1>
1C
b110 G
#951020000000
0!
0*
09
0>
0C
#951030000000
1!
1*
b111 6
19
1>
1C
b111 G
#951040000000
0!
0*
09
0>
0C
#951050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#951060000000
0!
0*
09
0>
0C
#951070000000
1!
1*
b1 6
19
1>
1C
b1 G
#951080000000
0!
0*
09
0>
0C
#951090000000
1!
1*
b10 6
19
1>
1C
b10 G
#951100000000
0!
0*
09
0>
0C
#951110000000
1!
1*
b11 6
19
1>
1C
b11 G
#951120000000
0!
0*
09
0>
0C
#951130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#951140000000
0!
0*
09
0>
0C
#951150000000
1!
1*
b101 6
19
1>
1C
b101 G
#951160000000
0!
0*
09
0>
0C
#951170000000
1!
1*
b110 6
19
1>
1C
b110 G
#951180000000
0!
0*
09
0>
0C
#951190000000
1!
1*
b111 6
19
1>
1C
b111 G
#951200000000
0!
0*
09
0>
0C
#951210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#951220000000
0!
0*
09
0>
0C
#951230000000
1!
1*
b1 6
19
1>
1C
b1 G
#951240000000
0!
0*
09
0>
0C
#951250000000
1!
1*
b10 6
19
1>
1C
b10 G
#951260000000
0!
0*
09
0>
0C
#951270000000
1!
1*
b11 6
19
1>
1C
b11 G
#951280000000
0!
0*
09
0>
0C
#951290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#951300000000
0!
0*
09
0>
0C
#951310000000
1!
1*
b101 6
19
1>
1C
b101 G
#951320000000
0!
0*
09
0>
0C
#951330000000
1!
1*
b110 6
19
1>
1C
b110 G
#951340000000
0!
0*
09
0>
0C
#951350000000
1!
1*
b111 6
19
1>
1C
b111 G
#951360000000
0!
1"
0*
1+
09
1:
0>
0C
#951370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#951380000000
0!
0*
09
0>
0C
#951390000000
1!
1*
b1 6
19
1>
1C
b1 G
#951400000000
0!
0*
09
0>
0C
#951410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#951420000000
0!
0*
09
0>
0C
#951430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#951440000000
0!
0*
09
0>
0C
#951450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#951460000000
0!
0*
09
0>
0C
#951470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#951480000000
0!
0#
0*
0,
09
0>
0?
0C
#951490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#951500000000
0!
0*
09
0>
0C
#951510000000
1!
1*
19
1>
1C
#951520000000
0!
0*
09
0>
0C
#951530000000
1!
1*
19
1>
1C
#951540000000
0!
0*
09
0>
0C
#951550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#951560000000
0!
0*
09
0>
0C
#951570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#951580000000
0!
0*
09
0>
0C
#951590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#951600000000
0!
0*
09
0>
0C
#951610000000
1!
1*
b10 6
19
1>
1C
b10 G
#951620000000
0!
0*
09
0>
0C
#951630000000
1!
1*
b11 6
19
1>
1C
b11 G
#951640000000
0!
0*
09
0>
0C
#951650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#951660000000
0!
0*
09
0>
0C
#951670000000
1!
1*
b101 6
19
1>
1C
b101 G
#951680000000
0!
0*
09
0>
0C
#951690000000
1!
1*
b110 6
19
1>
1C
b110 G
#951700000000
0!
0*
09
0>
0C
#951710000000
1!
1*
b111 6
19
1>
1C
b111 G
#951720000000
0!
0*
09
0>
0C
#951730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#951740000000
0!
0*
09
0>
0C
#951750000000
1!
1*
b1 6
19
1>
1C
b1 G
#951760000000
0!
0*
09
0>
0C
#951770000000
1!
1*
b10 6
19
1>
1C
b10 G
#951780000000
0!
0*
09
0>
0C
#951790000000
1!
1*
b11 6
19
1>
1C
b11 G
#951800000000
0!
0*
09
0>
0C
#951810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#951820000000
0!
0*
09
0>
0C
#951830000000
1!
1*
b101 6
19
1>
1C
b101 G
#951840000000
0!
0*
09
0>
0C
#951850000000
1!
1*
b110 6
19
1>
1C
b110 G
#951860000000
0!
0*
09
0>
0C
#951870000000
1!
1*
b111 6
19
1>
1C
b111 G
#951880000000
0!
0*
09
0>
0C
#951890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#951900000000
0!
0*
09
0>
0C
#951910000000
1!
1*
b1 6
19
1>
1C
b1 G
#951920000000
0!
0*
09
0>
0C
#951930000000
1!
1*
b10 6
19
1>
1C
b10 G
#951940000000
0!
0*
09
0>
0C
#951950000000
1!
1*
b11 6
19
1>
1C
b11 G
#951960000000
0!
0*
09
0>
0C
#951970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#951980000000
0!
0*
09
0>
0C
#951990000000
1!
1*
b101 6
19
1>
1C
b101 G
#952000000000
0!
0*
09
0>
0C
#952010000000
1!
1*
b110 6
19
1>
1C
b110 G
#952020000000
0!
0*
09
0>
0C
#952030000000
1!
1*
b111 6
19
1>
1C
b111 G
#952040000000
0!
1"
0*
1+
09
1:
0>
0C
#952050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#952060000000
0!
0*
09
0>
0C
#952070000000
1!
1*
b1 6
19
1>
1C
b1 G
#952080000000
0!
0*
09
0>
0C
#952090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#952100000000
0!
0*
09
0>
0C
#952110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#952120000000
0!
0*
09
0>
0C
#952130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#952140000000
0!
0*
09
0>
0C
#952150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#952160000000
0!
0#
0*
0,
09
0>
0?
0C
#952170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#952180000000
0!
0*
09
0>
0C
#952190000000
1!
1*
19
1>
1C
#952200000000
0!
0*
09
0>
0C
#952210000000
1!
1*
19
1>
1C
#952220000000
0!
0*
09
0>
0C
#952230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#952240000000
0!
0*
09
0>
0C
#952250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#952260000000
0!
0*
09
0>
0C
#952270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#952280000000
0!
0*
09
0>
0C
#952290000000
1!
1*
b10 6
19
1>
1C
b10 G
#952300000000
0!
0*
09
0>
0C
#952310000000
1!
1*
b11 6
19
1>
1C
b11 G
#952320000000
0!
0*
09
0>
0C
#952330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#952340000000
0!
0*
09
0>
0C
#952350000000
1!
1*
b101 6
19
1>
1C
b101 G
#952360000000
0!
0*
09
0>
0C
#952370000000
1!
1*
b110 6
19
1>
1C
b110 G
#952380000000
0!
0*
09
0>
0C
#952390000000
1!
1*
b111 6
19
1>
1C
b111 G
#952400000000
0!
0*
09
0>
0C
#952410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#952420000000
0!
0*
09
0>
0C
#952430000000
1!
1*
b1 6
19
1>
1C
b1 G
#952440000000
0!
0*
09
0>
0C
#952450000000
1!
1*
b10 6
19
1>
1C
b10 G
#952460000000
0!
0*
09
0>
0C
#952470000000
1!
1*
b11 6
19
1>
1C
b11 G
#952480000000
0!
0*
09
0>
0C
#952490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#952500000000
0!
0*
09
0>
0C
#952510000000
1!
1*
b101 6
19
1>
1C
b101 G
#952520000000
0!
0*
09
0>
0C
#952530000000
1!
1*
b110 6
19
1>
1C
b110 G
#952540000000
0!
0*
09
0>
0C
#952550000000
1!
1*
b111 6
19
1>
1C
b111 G
#952560000000
0!
0*
09
0>
0C
#952570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#952580000000
0!
0*
09
0>
0C
#952590000000
1!
1*
b1 6
19
1>
1C
b1 G
#952600000000
0!
0*
09
0>
0C
#952610000000
1!
1*
b10 6
19
1>
1C
b10 G
#952620000000
0!
0*
09
0>
0C
#952630000000
1!
1*
b11 6
19
1>
1C
b11 G
#952640000000
0!
0*
09
0>
0C
#952650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#952660000000
0!
0*
09
0>
0C
#952670000000
1!
1*
b101 6
19
1>
1C
b101 G
#952680000000
0!
0*
09
0>
0C
#952690000000
1!
1*
b110 6
19
1>
1C
b110 G
#952700000000
0!
0*
09
0>
0C
#952710000000
1!
1*
b111 6
19
1>
1C
b111 G
#952720000000
0!
1"
0*
1+
09
1:
0>
0C
#952730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#952740000000
0!
0*
09
0>
0C
#952750000000
1!
1*
b1 6
19
1>
1C
b1 G
#952760000000
0!
0*
09
0>
0C
#952770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#952780000000
0!
0*
09
0>
0C
#952790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#952800000000
0!
0*
09
0>
0C
#952810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#952820000000
0!
0*
09
0>
0C
#952830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#952840000000
0!
0#
0*
0,
09
0>
0?
0C
#952850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#952860000000
0!
0*
09
0>
0C
#952870000000
1!
1*
19
1>
1C
#952880000000
0!
0*
09
0>
0C
#952890000000
1!
1*
19
1>
1C
#952900000000
0!
0*
09
0>
0C
#952910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#952920000000
0!
0*
09
0>
0C
#952930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#952940000000
0!
0*
09
0>
0C
#952950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#952960000000
0!
0*
09
0>
0C
#952970000000
1!
1*
b10 6
19
1>
1C
b10 G
#952980000000
0!
0*
09
0>
0C
#952990000000
1!
1*
b11 6
19
1>
1C
b11 G
#953000000000
0!
0*
09
0>
0C
#953010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#953020000000
0!
0*
09
0>
0C
#953030000000
1!
1*
b101 6
19
1>
1C
b101 G
#953040000000
0!
0*
09
0>
0C
#953050000000
1!
1*
b110 6
19
1>
1C
b110 G
#953060000000
0!
0*
09
0>
0C
#953070000000
1!
1*
b111 6
19
1>
1C
b111 G
#953080000000
0!
0*
09
0>
0C
#953090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#953100000000
0!
0*
09
0>
0C
#953110000000
1!
1*
b1 6
19
1>
1C
b1 G
#953120000000
0!
0*
09
0>
0C
#953130000000
1!
1*
b10 6
19
1>
1C
b10 G
#953140000000
0!
0*
09
0>
0C
#953150000000
1!
1*
b11 6
19
1>
1C
b11 G
#953160000000
0!
0*
09
0>
0C
#953170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#953180000000
0!
0*
09
0>
0C
#953190000000
1!
1*
b101 6
19
1>
1C
b101 G
#953200000000
0!
0*
09
0>
0C
#953210000000
1!
1*
b110 6
19
1>
1C
b110 G
#953220000000
0!
0*
09
0>
0C
#953230000000
1!
1*
b111 6
19
1>
1C
b111 G
#953240000000
0!
0*
09
0>
0C
#953250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#953260000000
0!
0*
09
0>
0C
#953270000000
1!
1*
b1 6
19
1>
1C
b1 G
#953280000000
0!
0*
09
0>
0C
#953290000000
1!
1*
b10 6
19
1>
1C
b10 G
#953300000000
0!
0*
09
0>
0C
#953310000000
1!
1*
b11 6
19
1>
1C
b11 G
#953320000000
0!
0*
09
0>
0C
#953330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#953340000000
0!
0*
09
0>
0C
#953350000000
1!
1*
b101 6
19
1>
1C
b101 G
#953360000000
0!
0*
09
0>
0C
#953370000000
1!
1*
b110 6
19
1>
1C
b110 G
#953380000000
0!
0*
09
0>
0C
#953390000000
1!
1*
b111 6
19
1>
1C
b111 G
#953400000000
0!
1"
0*
1+
09
1:
0>
0C
#953410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#953420000000
0!
0*
09
0>
0C
#953430000000
1!
1*
b1 6
19
1>
1C
b1 G
#953440000000
0!
0*
09
0>
0C
#953450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#953460000000
0!
0*
09
0>
0C
#953470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#953480000000
0!
0*
09
0>
0C
#953490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#953500000000
0!
0*
09
0>
0C
#953510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#953520000000
0!
0#
0*
0,
09
0>
0?
0C
#953530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#953540000000
0!
0*
09
0>
0C
#953550000000
1!
1*
19
1>
1C
#953560000000
0!
0*
09
0>
0C
#953570000000
1!
1*
19
1>
1C
#953580000000
0!
0*
09
0>
0C
#953590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#953600000000
0!
0*
09
0>
0C
#953610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#953620000000
0!
0*
09
0>
0C
#953630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#953640000000
0!
0*
09
0>
0C
#953650000000
1!
1*
b10 6
19
1>
1C
b10 G
#953660000000
0!
0*
09
0>
0C
#953670000000
1!
1*
b11 6
19
1>
1C
b11 G
#953680000000
0!
0*
09
0>
0C
#953690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#953700000000
0!
0*
09
0>
0C
#953710000000
1!
1*
b101 6
19
1>
1C
b101 G
#953720000000
0!
0*
09
0>
0C
#953730000000
1!
1*
b110 6
19
1>
1C
b110 G
#953740000000
0!
0*
09
0>
0C
#953750000000
1!
1*
b111 6
19
1>
1C
b111 G
#953760000000
0!
0*
09
0>
0C
#953770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#953780000000
0!
0*
09
0>
0C
#953790000000
1!
1*
b1 6
19
1>
1C
b1 G
#953800000000
0!
0*
09
0>
0C
#953810000000
1!
1*
b10 6
19
1>
1C
b10 G
#953820000000
0!
0*
09
0>
0C
#953830000000
1!
1*
b11 6
19
1>
1C
b11 G
#953840000000
0!
0*
09
0>
0C
#953850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#953860000000
0!
0*
09
0>
0C
#953870000000
1!
1*
b101 6
19
1>
1C
b101 G
#953880000000
0!
0*
09
0>
0C
#953890000000
1!
1*
b110 6
19
1>
1C
b110 G
#953900000000
0!
0*
09
0>
0C
#953910000000
1!
1*
b111 6
19
1>
1C
b111 G
#953920000000
0!
0*
09
0>
0C
#953930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#953940000000
0!
0*
09
0>
0C
#953950000000
1!
1*
b1 6
19
1>
1C
b1 G
#953960000000
0!
0*
09
0>
0C
#953970000000
1!
1*
b10 6
19
1>
1C
b10 G
#953980000000
0!
0*
09
0>
0C
#953990000000
1!
1*
b11 6
19
1>
1C
b11 G
#954000000000
0!
0*
09
0>
0C
#954010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#954020000000
0!
0*
09
0>
0C
#954030000000
1!
1*
b101 6
19
1>
1C
b101 G
#954040000000
0!
0*
09
0>
0C
#954050000000
1!
1*
b110 6
19
1>
1C
b110 G
#954060000000
0!
0*
09
0>
0C
#954070000000
1!
1*
b111 6
19
1>
1C
b111 G
#954080000000
0!
1"
0*
1+
09
1:
0>
0C
#954090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#954100000000
0!
0*
09
0>
0C
#954110000000
1!
1*
b1 6
19
1>
1C
b1 G
#954120000000
0!
0*
09
0>
0C
#954130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#954140000000
0!
0*
09
0>
0C
#954150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#954160000000
0!
0*
09
0>
0C
#954170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#954180000000
0!
0*
09
0>
0C
#954190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#954200000000
0!
0#
0*
0,
09
0>
0?
0C
#954210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#954220000000
0!
0*
09
0>
0C
#954230000000
1!
1*
19
1>
1C
#954240000000
0!
0*
09
0>
0C
#954250000000
1!
1*
19
1>
1C
#954260000000
0!
0*
09
0>
0C
#954270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#954280000000
0!
0*
09
0>
0C
#954290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#954300000000
0!
0*
09
0>
0C
#954310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#954320000000
0!
0*
09
0>
0C
#954330000000
1!
1*
b10 6
19
1>
1C
b10 G
#954340000000
0!
0*
09
0>
0C
#954350000000
1!
1*
b11 6
19
1>
1C
b11 G
#954360000000
0!
0*
09
0>
0C
#954370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#954380000000
0!
0*
09
0>
0C
#954390000000
1!
1*
b101 6
19
1>
1C
b101 G
#954400000000
0!
0*
09
0>
0C
#954410000000
1!
1*
b110 6
19
1>
1C
b110 G
#954420000000
0!
0*
09
0>
0C
#954430000000
1!
1*
b111 6
19
1>
1C
b111 G
#954440000000
0!
0*
09
0>
0C
#954450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#954460000000
0!
0*
09
0>
0C
#954470000000
1!
1*
b1 6
19
1>
1C
b1 G
#954480000000
0!
0*
09
0>
0C
#954490000000
1!
1*
b10 6
19
1>
1C
b10 G
#954500000000
0!
0*
09
0>
0C
#954510000000
1!
1*
b11 6
19
1>
1C
b11 G
#954520000000
0!
0*
09
0>
0C
#954530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#954540000000
0!
0*
09
0>
0C
#954550000000
1!
1*
b101 6
19
1>
1C
b101 G
#954560000000
0!
0*
09
0>
0C
#954570000000
1!
1*
b110 6
19
1>
1C
b110 G
#954580000000
0!
0*
09
0>
0C
#954590000000
1!
1*
b111 6
19
1>
1C
b111 G
#954600000000
0!
0*
09
0>
0C
#954610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#954620000000
0!
0*
09
0>
0C
#954630000000
1!
1*
b1 6
19
1>
1C
b1 G
#954640000000
0!
0*
09
0>
0C
#954650000000
1!
1*
b10 6
19
1>
1C
b10 G
#954660000000
0!
0*
09
0>
0C
#954670000000
1!
1*
b11 6
19
1>
1C
b11 G
#954680000000
0!
0*
09
0>
0C
#954690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#954700000000
0!
0*
09
0>
0C
#954710000000
1!
1*
b101 6
19
1>
1C
b101 G
#954720000000
0!
0*
09
0>
0C
#954730000000
1!
1*
b110 6
19
1>
1C
b110 G
#954740000000
0!
0*
09
0>
0C
#954750000000
1!
1*
b111 6
19
1>
1C
b111 G
#954760000000
0!
1"
0*
1+
09
1:
0>
0C
#954770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#954780000000
0!
0*
09
0>
0C
#954790000000
1!
1*
b1 6
19
1>
1C
b1 G
#954800000000
0!
0*
09
0>
0C
#954810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#954820000000
0!
0*
09
0>
0C
#954830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#954840000000
0!
0*
09
0>
0C
#954850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#954860000000
0!
0*
09
0>
0C
#954870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#954880000000
0!
0#
0*
0,
09
0>
0?
0C
#954890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#954900000000
0!
0*
09
0>
0C
#954910000000
1!
1*
19
1>
1C
#954920000000
0!
0*
09
0>
0C
#954930000000
1!
1*
19
1>
1C
#954940000000
0!
0*
09
0>
0C
#954950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#954960000000
0!
0*
09
0>
0C
#954970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#954980000000
0!
0*
09
0>
0C
#954990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#955000000000
0!
0*
09
0>
0C
#955010000000
1!
1*
b10 6
19
1>
1C
b10 G
#955020000000
0!
0*
09
0>
0C
#955030000000
1!
1*
b11 6
19
1>
1C
b11 G
#955040000000
0!
0*
09
0>
0C
#955050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#955060000000
0!
0*
09
0>
0C
#955070000000
1!
1*
b101 6
19
1>
1C
b101 G
#955080000000
0!
0*
09
0>
0C
#955090000000
1!
1*
b110 6
19
1>
1C
b110 G
#955100000000
0!
0*
09
0>
0C
#955110000000
1!
1*
b111 6
19
1>
1C
b111 G
#955120000000
0!
0*
09
0>
0C
#955130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#955140000000
0!
0*
09
0>
0C
#955150000000
1!
1*
b1 6
19
1>
1C
b1 G
#955160000000
0!
0*
09
0>
0C
#955170000000
1!
1*
b10 6
19
1>
1C
b10 G
#955180000000
0!
0*
09
0>
0C
#955190000000
1!
1*
b11 6
19
1>
1C
b11 G
#955200000000
0!
0*
09
0>
0C
#955210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#955220000000
0!
0*
09
0>
0C
#955230000000
1!
1*
b101 6
19
1>
1C
b101 G
#955240000000
0!
0*
09
0>
0C
#955250000000
1!
1*
b110 6
19
1>
1C
b110 G
#955260000000
0!
0*
09
0>
0C
#955270000000
1!
1*
b111 6
19
1>
1C
b111 G
#955280000000
0!
0*
09
0>
0C
#955290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#955300000000
0!
0*
09
0>
0C
#955310000000
1!
1*
b1 6
19
1>
1C
b1 G
#955320000000
0!
0*
09
0>
0C
#955330000000
1!
1*
b10 6
19
1>
1C
b10 G
#955340000000
0!
0*
09
0>
0C
#955350000000
1!
1*
b11 6
19
1>
1C
b11 G
#955360000000
0!
0*
09
0>
0C
#955370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#955380000000
0!
0*
09
0>
0C
#955390000000
1!
1*
b101 6
19
1>
1C
b101 G
#955400000000
0!
0*
09
0>
0C
#955410000000
1!
1*
b110 6
19
1>
1C
b110 G
#955420000000
0!
0*
09
0>
0C
#955430000000
1!
1*
b111 6
19
1>
1C
b111 G
#955440000000
0!
1"
0*
1+
09
1:
0>
0C
#955450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#955460000000
0!
0*
09
0>
0C
#955470000000
1!
1*
b1 6
19
1>
1C
b1 G
#955480000000
0!
0*
09
0>
0C
#955490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#955500000000
0!
0*
09
0>
0C
#955510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#955520000000
0!
0*
09
0>
0C
#955530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#955540000000
0!
0*
09
0>
0C
#955550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#955560000000
0!
0#
0*
0,
09
0>
0?
0C
#955570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#955580000000
0!
0*
09
0>
0C
#955590000000
1!
1*
19
1>
1C
#955600000000
0!
0*
09
0>
0C
#955610000000
1!
1*
19
1>
1C
#955620000000
0!
0*
09
0>
0C
#955630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#955640000000
0!
0*
09
0>
0C
#955650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#955660000000
0!
0*
09
0>
0C
#955670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#955680000000
0!
0*
09
0>
0C
#955690000000
1!
1*
b10 6
19
1>
1C
b10 G
#955700000000
0!
0*
09
0>
0C
#955710000000
1!
1*
b11 6
19
1>
1C
b11 G
#955720000000
0!
0*
09
0>
0C
#955730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#955740000000
0!
0*
09
0>
0C
#955750000000
1!
1*
b101 6
19
1>
1C
b101 G
#955760000000
0!
0*
09
0>
0C
#955770000000
1!
1*
b110 6
19
1>
1C
b110 G
#955780000000
0!
0*
09
0>
0C
#955790000000
1!
1*
b111 6
19
1>
1C
b111 G
#955800000000
0!
0*
09
0>
0C
#955810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#955820000000
0!
0*
09
0>
0C
#955830000000
1!
1*
b1 6
19
1>
1C
b1 G
#955840000000
0!
0*
09
0>
0C
#955850000000
1!
1*
b10 6
19
1>
1C
b10 G
#955860000000
0!
0*
09
0>
0C
#955870000000
1!
1*
b11 6
19
1>
1C
b11 G
#955880000000
0!
0*
09
0>
0C
#955890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#955900000000
0!
0*
09
0>
0C
#955910000000
1!
1*
b101 6
19
1>
1C
b101 G
#955920000000
0!
0*
09
0>
0C
#955930000000
1!
1*
b110 6
19
1>
1C
b110 G
#955940000000
0!
0*
09
0>
0C
#955950000000
1!
1*
b111 6
19
1>
1C
b111 G
#955960000000
0!
0*
09
0>
0C
#955970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#955980000000
0!
0*
09
0>
0C
#955990000000
1!
1*
b1 6
19
1>
1C
b1 G
#956000000000
0!
0*
09
0>
0C
#956010000000
1!
1*
b10 6
19
1>
1C
b10 G
#956020000000
0!
0*
09
0>
0C
#956030000000
1!
1*
b11 6
19
1>
1C
b11 G
#956040000000
0!
0*
09
0>
0C
#956050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#956060000000
0!
0*
09
0>
0C
#956070000000
1!
1*
b101 6
19
1>
1C
b101 G
#956080000000
0!
0*
09
0>
0C
#956090000000
1!
1*
b110 6
19
1>
1C
b110 G
#956100000000
0!
0*
09
0>
0C
#956110000000
1!
1*
b111 6
19
1>
1C
b111 G
#956120000000
0!
1"
0*
1+
09
1:
0>
0C
#956130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#956140000000
0!
0*
09
0>
0C
#956150000000
1!
1*
b1 6
19
1>
1C
b1 G
#956160000000
0!
0*
09
0>
0C
#956170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#956180000000
0!
0*
09
0>
0C
#956190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#956200000000
0!
0*
09
0>
0C
#956210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#956220000000
0!
0*
09
0>
0C
#956230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#956240000000
0!
0#
0*
0,
09
0>
0?
0C
#956250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#956260000000
0!
0*
09
0>
0C
#956270000000
1!
1*
19
1>
1C
#956280000000
0!
0*
09
0>
0C
#956290000000
1!
1*
19
1>
1C
#956300000000
0!
0*
09
0>
0C
#956310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#956320000000
0!
0*
09
0>
0C
#956330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#956340000000
0!
0*
09
0>
0C
#956350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#956360000000
0!
0*
09
0>
0C
#956370000000
1!
1*
b10 6
19
1>
1C
b10 G
#956380000000
0!
0*
09
0>
0C
#956390000000
1!
1*
b11 6
19
1>
1C
b11 G
#956400000000
0!
0*
09
0>
0C
#956410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#956420000000
0!
0*
09
0>
0C
#956430000000
1!
1*
b101 6
19
1>
1C
b101 G
#956440000000
0!
0*
09
0>
0C
#956450000000
1!
1*
b110 6
19
1>
1C
b110 G
#956460000000
0!
0*
09
0>
0C
#956470000000
1!
1*
b111 6
19
1>
1C
b111 G
#956480000000
0!
0*
09
0>
0C
#956490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#956500000000
0!
0*
09
0>
0C
#956510000000
1!
1*
b1 6
19
1>
1C
b1 G
#956520000000
0!
0*
09
0>
0C
#956530000000
1!
1*
b10 6
19
1>
1C
b10 G
#956540000000
0!
0*
09
0>
0C
#956550000000
1!
1*
b11 6
19
1>
1C
b11 G
#956560000000
0!
0*
09
0>
0C
#956570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#956580000000
0!
0*
09
0>
0C
#956590000000
1!
1*
b101 6
19
1>
1C
b101 G
#956600000000
0!
0*
09
0>
0C
#956610000000
1!
1*
b110 6
19
1>
1C
b110 G
#956620000000
0!
0*
09
0>
0C
#956630000000
1!
1*
b111 6
19
1>
1C
b111 G
#956640000000
0!
0*
09
0>
0C
#956650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#956660000000
0!
0*
09
0>
0C
#956670000000
1!
1*
b1 6
19
1>
1C
b1 G
#956680000000
0!
0*
09
0>
0C
#956690000000
1!
1*
b10 6
19
1>
1C
b10 G
#956700000000
0!
0*
09
0>
0C
#956710000000
1!
1*
b11 6
19
1>
1C
b11 G
#956720000000
0!
0*
09
0>
0C
#956730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#956740000000
0!
0*
09
0>
0C
#956750000000
1!
1*
b101 6
19
1>
1C
b101 G
#956760000000
0!
0*
09
0>
0C
#956770000000
1!
1*
b110 6
19
1>
1C
b110 G
#956780000000
0!
0*
09
0>
0C
#956790000000
1!
1*
b111 6
19
1>
1C
b111 G
#956800000000
0!
1"
0*
1+
09
1:
0>
0C
#956810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#956820000000
0!
0*
09
0>
0C
#956830000000
1!
1*
b1 6
19
1>
1C
b1 G
#956840000000
0!
0*
09
0>
0C
#956850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#956860000000
0!
0*
09
0>
0C
#956870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#956880000000
0!
0*
09
0>
0C
#956890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#956900000000
0!
0*
09
0>
0C
#956910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#956920000000
0!
0#
0*
0,
09
0>
0?
0C
#956930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#956940000000
0!
0*
09
0>
0C
#956950000000
1!
1*
19
1>
1C
#956960000000
0!
0*
09
0>
0C
#956970000000
1!
1*
19
1>
1C
#956980000000
0!
0*
09
0>
0C
#956990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#957000000000
0!
0*
09
0>
0C
#957010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#957020000000
0!
0*
09
0>
0C
#957030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#957040000000
0!
0*
09
0>
0C
#957050000000
1!
1*
b10 6
19
1>
1C
b10 G
#957060000000
0!
0*
09
0>
0C
#957070000000
1!
1*
b11 6
19
1>
1C
b11 G
#957080000000
0!
0*
09
0>
0C
#957090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#957100000000
0!
0*
09
0>
0C
#957110000000
1!
1*
b101 6
19
1>
1C
b101 G
#957120000000
0!
0*
09
0>
0C
#957130000000
1!
1*
b110 6
19
1>
1C
b110 G
#957140000000
0!
0*
09
0>
0C
#957150000000
1!
1*
b111 6
19
1>
1C
b111 G
#957160000000
0!
0*
09
0>
0C
#957170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#957180000000
0!
0*
09
0>
0C
#957190000000
1!
1*
b1 6
19
1>
1C
b1 G
#957200000000
0!
0*
09
0>
0C
#957210000000
1!
1*
b10 6
19
1>
1C
b10 G
#957220000000
0!
0*
09
0>
0C
#957230000000
1!
1*
b11 6
19
1>
1C
b11 G
#957240000000
0!
0*
09
0>
0C
#957250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#957260000000
0!
0*
09
0>
0C
#957270000000
1!
1*
b101 6
19
1>
1C
b101 G
#957280000000
0!
0*
09
0>
0C
#957290000000
1!
1*
b110 6
19
1>
1C
b110 G
#957300000000
0!
0*
09
0>
0C
#957310000000
1!
1*
b111 6
19
1>
1C
b111 G
#957320000000
0!
0*
09
0>
0C
#957330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#957340000000
0!
0*
09
0>
0C
#957350000000
1!
1*
b1 6
19
1>
1C
b1 G
#957360000000
0!
0*
09
0>
0C
#957370000000
1!
1*
b10 6
19
1>
1C
b10 G
#957380000000
0!
0*
09
0>
0C
#957390000000
1!
1*
b11 6
19
1>
1C
b11 G
#957400000000
0!
0*
09
0>
0C
#957410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#957420000000
0!
0*
09
0>
0C
#957430000000
1!
1*
b101 6
19
1>
1C
b101 G
#957440000000
0!
0*
09
0>
0C
#957450000000
1!
1*
b110 6
19
1>
1C
b110 G
#957460000000
0!
0*
09
0>
0C
#957470000000
1!
1*
b111 6
19
1>
1C
b111 G
#957480000000
0!
1"
0*
1+
09
1:
0>
0C
#957490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#957500000000
0!
0*
09
0>
0C
#957510000000
1!
1*
b1 6
19
1>
1C
b1 G
#957520000000
0!
0*
09
0>
0C
#957530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#957540000000
0!
0*
09
0>
0C
#957550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#957560000000
0!
0*
09
0>
0C
#957570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#957580000000
0!
0*
09
0>
0C
#957590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#957600000000
0!
0#
0*
0,
09
0>
0?
0C
#957610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#957620000000
0!
0*
09
0>
0C
#957630000000
1!
1*
19
1>
1C
#957640000000
0!
0*
09
0>
0C
#957650000000
1!
1*
19
1>
1C
#957660000000
0!
0*
09
0>
0C
#957670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#957680000000
0!
0*
09
0>
0C
#957690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#957700000000
0!
0*
09
0>
0C
#957710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#957720000000
0!
0*
09
0>
0C
#957730000000
1!
1*
b10 6
19
1>
1C
b10 G
#957740000000
0!
0*
09
0>
0C
#957750000000
1!
1*
b11 6
19
1>
1C
b11 G
#957760000000
0!
0*
09
0>
0C
#957770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#957780000000
0!
0*
09
0>
0C
#957790000000
1!
1*
b101 6
19
1>
1C
b101 G
#957800000000
0!
0*
09
0>
0C
#957810000000
1!
1*
b110 6
19
1>
1C
b110 G
#957820000000
0!
0*
09
0>
0C
#957830000000
1!
1*
b111 6
19
1>
1C
b111 G
#957840000000
0!
0*
09
0>
0C
#957850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#957860000000
0!
0*
09
0>
0C
#957870000000
1!
1*
b1 6
19
1>
1C
b1 G
#957880000000
0!
0*
09
0>
0C
#957890000000
1!
1*
b10 6
19
1>
1C
b10 G
#957900000000
0!
0*
09
0>
0C
#957910000000
1!
1*
b11 6
19
1>
1C
b11 G
#957920000000
0!
0*
09
0>
0C
#957930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#957940000000
0!
0*
09
0>
0C
#957950000000
1!
1*
b101 6
19
1>
1C
b101 G
#957960000000
0!
0*
09
0>
0C
#957970000000
1!
1*
b110 6
19
1>
1C
b110 G
#957980000000
0!
0*
09
0>
0C
#957990000000
1!
1*
b111 6
19
1>
1C
b111 G
#958000000000
0!
0*
09
0>
0C
#958010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#958020000000
0!
0*
09
0>
0C
#958030000000
1!
1*
b1 6
19
1>
1C
b1 G
#958040000000
0!
0*
09
0>
0C
#958050000000
1!
1*
b10 6
19
1>
1C
b10 G
#958060000000
0!
0*
09
0>
0C
#958070000000
1!
1*
b11 6
19
1>
1C
b11 G
#958080000000
0!
0*
09
0>
0C
#958090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#958100000000
0!
0*
09
0>
0C
#958110000000
1!
1*
b101 6
19
1>
1C
b101 G
#958120000000
0!
0*
09
0>
0C
#958130000000
1!
1*
b110 6
19
1>
1C
b110 G
#958140000000
0!
0*
09
0>
0C
#958150000000
1!
1*
b111 6
19
1>
1C
b111 G
#958160000000
0!
1"
0*
1+
09
1:
0>
0C
#958170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#958180000000
0!
0*
09
0>
0C
#958190000000
1!
1*
b1 6
19
1>
1C
b1 G
#958200000000
0!
0*
09
0>
0C
#958210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#958220000000
0!
0*
09
0>
0C
#958230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#958240000000
0!
0*
09
0>
0C
#958250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#958260000000
0!
0*
09
0>
0C
#958270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#958280000000
0!
0#
0*
0,
09
0>
0?
0C
#958290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#958300000000
0!
0*
09
0>
0C
#958310000000
1!
1*
19
1>
1C
#958320000000
0!
0*
09
0>
0C
#958330000000
1!
1*
19
1>
1C
#958340000000
0!
0*
09
0>
0C
#958350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#958360000000
0!
0*
09
0>
0C
#958370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#958380000000
0!
0*
09
0>
0C
#958390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#958400000000
0!
0*
09
0>
0C
#958410000000
1!
1*
b10 6
19
1>
1C
b10 G
#958420000000
0!
0*
09
0>
0C
#958430000000
1!
1*
b11 6
19
1>
1C
b11 G
#958440000000
0!
0*
09
0>
0C
#958450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#958460000000
0!
0*
09
0>
0C
#958470000000
1!
1*
b101 6
19
1>
1C
b101 G
#958480000000
0!
0*
09
0>
0C
#958490000000
1!
1*
b110 6
19
1>
1C
b110 G
#958500000000
0!
0*
09
0>
0C
#958510000000
1!
1*
b111 6
19
1>
1C
b111 G
#958520000000
0!
0*
09
0>
0C
#958530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#958540000000
0!
0*
09
0>
0C
#958550000000
1!
1*
b1 6
19
1>
1C
b1 G
#958560000000
0!
0*
09
0>
0C
#958570000000
1!
1*
b10 6
19
1>
1C
b10 G
#958580000000
0!
0*
09
0>
0C
#958590000000
1!
1*
b11 6
19
1>
1C
b11 G
#958600000000
0!
0*
09
0>
0C
#958610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#958620000000
0!
0*
09
0>
0C
#958630000000
1!
1*
b101 6
19
1>
1C
b101 G
#958640000000
0!
0*
09
0>
0C
#958650000000
1!
1*
b110 6
19
1>
1C
b110 G
#958660000000
0!
0*
09
0>
0C
#958670000000
1!
1*
b111 6
19
1>
1C
b111 G
#958680000000
0!
0*
09
0>
0C
#958690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#958700000000
0!
0*
09
0>
0C
#958710000000
1!
1*
b1 6
19
1>
1C
b1 G
#958720000000
0!
0*
09
0>
0C
#958730000000
1!
1*
b10 6
19
1>
1C
b10 G
#958740000000
0!
0*
09
0>
0C
#958750000000
1!
1*
b11 6
19
1>
1C
b11 G
#958760000000
0!
0*
09
0>
0C
#958770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#958780000000
0!
0*
09
0>
0C
#958790000000
1!
1*
b101 6
19
1>
1C
b101 G
#958800000000
0!
0*
09
0>
0C
#958810000000
1!
1*
b110 6
19
1>
1C
b110 G
#958820000000
0!
0*
09
0>
0C
#958830000000
1!
1*
b111 6
19
1>
1C
b111 G
#958840000000
0!
1"
0*
1+
09
1:
0>
0C
#958850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#958860000000
0!
0*
09
0>
0C
#958870000000
1!
1*
b1 6
19
1>
1C
b1 G
#958880000000
0!
0*
09
0>
0C
#958890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#958900000000
0!
0*
09
0>
0C
#958910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#958920000000
0!
0*
09
0>
0C
#958930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#958940000000
0!
0*
09
0>
0C
#958950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#958960000000
0!
0#
0*
0,
09
0>
0?
0C
#958970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#958980000000
0!
0*
09
0>
0C
#958990000000
1!
1*
19
1>
1C
#959000000000
0!
0*
09
0>
0C
#959010000000
1!
1*
19
1>
1C
#959020000000
0!
0*
09
0>
0C
#959030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#959040000000
0!
0*
09
0>
0C
#959050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#959060000000
0!
0*
09
0>
0C
#959070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#959080000000
0!
0*
09
0>
0C
#959090000000
1!
1*
b10 6
19
1>
1C
b10 G
#959100000000
0!
0*
09
0>
0C
#959110000000
1!
1*
b11 6
19
1>
1C
b11 G
#959120000000
0!
0*
09
0>
0C
#959130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#959140000000
0!
0*
09
0>
0C
#959150000000
1!
1*
b101 6
19
1>
1C
b101 G
#959160000000
0!
0*
09
0>
0C
#959170000000
1!
1*
b110 6
19
1>
1C
b110 G
#959180000000
0!
0*
09
0>
0C
#959190000000
1!
1*
b111 6
19
1>
1C
b111 G
#959200000000
0!
0*
09
0>
0C
#959210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#959220000000
0!
0*
09
0>
0C
#959230000000
1!
1*
b1 6
19
1>
1C
b1 G
#959240000000
0!
0*
09
0>
0C
#959250000000
1!
1*
b10 6
19
1>
1C
b10 G
#959260000000
0!
0*
09
0>
0C
#959270000000
1!
1*
b11 6
19
1>
1C
b11 G
#959280000000
0!
0*
09
0>
0C
#959290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#959300000000
0!
0*
09
0>
0C
#959310000000
1!
1*
b101 6
19
1>
1C
b101 G
#959320000000
0!
0*
09
0>
0C
#959330000000
1!
1*
b110 6
19
1>
1C
b110 G
#959340000000
0!
0*
09
0>
0C
#959350000000
1!
1*
b111 6
19
1>
1C
b111 G
#959360000000
0!
0*
09
0>
0C
#959370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#959380000000
0!
0*
09
0>
0C
#959390000000
1!
1*
b1 6
19
1>
1C
b1 G
#959400000000
0!
0*
09
0>
0C
#959410000000
1!
1*
b10 6
19
1>
1C
b10 G
#959420000000
0!
0*
09
0>
0C
#959430000000
1!
1*
b11 6
19
1>
1C
b11 G
#959440000000
0!
0*
09
0>
0C
#959450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#959460000000
0!
0*
09
0>
0C
#959470000000
1!
1*
b101 6
19
1>
1C
b101 G
#959480000000
0!
0*
09
0>
0C
#959490000000
1!
1*
b110 6
19
1>
1C
b110 G
#959500000000
0!
0*
09
0>
0C
#959510000000
1!
1*
b111 6
19
1>
1C
b111 G
#959520000000
0!
1"
0*
1+
09
1:
0>
0C
#959530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#959540000000
0!
0*
09
0>
0C
#959550000000
1!
1*
b1 6
19
1>
1C
b1 G
#959560000000
0!
0*
09
0>
0C
#959570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#959580000000
0!
0*
09
0>
0C
#959590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#959600000000
0!
0*
09
0>
0C
#959610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#959620000000
0!
0*
09
0>
0C
#959630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#959640000000
0!
0#
0*
0,
09
0>
0?
0C
#959650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#959660000000
0!
0*
09
0>
0C
#959670000000
1!
1*
19
1>
1C
#959680000000
0!
0*
09
0>
0C
#959690000000
1!
1*
19
1>
1C
#959700000000
0!
0*
09
0>
0C
#959710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#959720000000
0!
0*
09
0>
0C
#959730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#959740000000
0!
0*
09
0>
0C
#959750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#959760000000
0!
0*
09
0>
0C
#959770000000
1!
1*
b10 6
19
1>
1C
b10 G
#959780000000
0!
0*
09
0>
0C
#959790000000
1!
1*
b11 6
19
1>
1C
b11 G
#959800000000
0!
0*
09
0>
0C
#959810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#959820000000
0!
0*
09
0>
0C
#959830000000
1!
1*
b101 6
19
1>
1C
b101 G
#959840000000
0!
0*
09
0>
0C
#959850000000
1!
1*
b110 6
19
1>
1C
b110 G
#959860000000
0!
0*
09
0>
0C
#959870000000
1!
1*
b111 6
19
1>
1C
b111 G
#959880000000
0!
0*
09
0>
0C
#959890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#959900000000
0!
0*
09
0>
0C
#959910000000
1!
1*
b1 6
19
1>
1C
b1 G
#959920000000
0!
0*
09
0>
0C
#959930000000
1!
1*
b10 6
19
1>
1C
b10 G
#959940000000
0!
0*
09
0>
0C
#959950000000
1!
1*
b11 6
19
1>
1C
b11 G
#959960000000
0!
0*
09
0>
0C
#959970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#959980000000
0!
0*
09
0>
0C
#959990000000
1!
1*
b101 6
19
1>
1C
b101 G
#960000000000
0!
0*
09
0>
0C
#960010000000
1!
1*
b110 6
19
1>
1C
b110 G
#960020000000
0!
0*
09
0>
0C
#960030000000
1!
1*
b111 6
19
1>
1C
b111 G
#960040000000
0!
0*
09
0>
0C
#960050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#960060000000
0!
0*
09
0>
0C
#960070000000
1!
1*
b1 6
19
1>
1C
b1 G
#960080000000
0!
0*
09
0>
0C
#960090000000
1!
1*
b10 6
19
1>
1C
b10 G
#960100000000
0!
0*
09
0>
0C
#960110000000
1!
1*
b11 6
19
1>
1C
b11 G
#960120000000
0!
0*
09
0>
0C
#960130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#960140000000
0!
0*
09
0>
0C
#960150000000
1!
1*
b101 6
19
1>
1C
b101 G
#960160000000
0!
0*
09
0>
0C
#960170000000
1!
1*
b110 6
19
1>
1C
b110 G
#960180000000
0!
0*
09
0>
0C
#960190000000
1!
1*
b111 6
19
1>
1C
b111 G
#960200000000
0!
1"
0*
1+
09
1:
0>
0C
#960210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#960220000000
0!
0*
09
0>
0C
#960230000000
1!
1*
b1 6
19
1>
1C
b1 G
#960240000000
0!
0*
09
0>
0C
#960250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#960260000000
0!
0*
09
0>
0C
#960270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#960280000000
0!
0*
09
0>
0C
#960290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#960300000000
0!
0*
09
0>
0C
#960310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#960320000000
0!
0#
0*
0,
09
0>
0?
0C
#960330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#960340000000
0!
0*
09
0>
0C
#960350000000
1!
1*
19
1>
1C
#960360000000
0!
0*
09
0>
0C
#960370000000
1!
1*
19
1>
1C
#960380000000
0!
0*
09
0>
0C
#960390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#960400000000
0!
0*
09
0>
0C
#960410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#960420000000
0!
0*
09
0>
0C
#960430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#960440000000
0!
0*
09
0>
0C
#960450000000
1!
1*
b10 6
19
1>
1C
b10 G
#960460000000
0!
0*
09
0>
0C
#960470000000
1!
1*
b11 6
19
1>
1C
b11 G
#960480000000
0!
0*
09
0>
0C
#960490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#960500000000
0!
0*
09
0>
0C
#960510000000
1!
1*
b101 6
19
1>
1C
b101 G
#960520000000
0!
0*
09
0>
0C
#960530000000
1!
1*
b110 6
19
1>
1C
b110 G
#960540000000
0!
0*
09
0>
0C
#960550000000
1!
1*
b111 6
19
1>
1C
b111 G
#960560000000
0!
0*
09
0>
0C
#960570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#960580000000
0!
0*
09
0>
0C
#960590000000
1!
1*
b1 6
19
1>
1C
b1 G
#960600000000
0!
0*
09
0>
0C
#960610000000
1!
1*
b10 6
19
1>
1C
b10 G
#960620000000
0!
0*
09
0>
0C
#960630000000
1!
1*
b11 6
19
1>
1C
b11 G
#960640000000
0!
0*
09
0>
0C
#960650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#960660000000
0!
0*
09
0>
0C
#960670000000
1!
1*
b101 6
19
1>
1C
b101 G
#960680000000
0!
0*
09
0>
0C
#960690000000
1!
1*
b110 6
19
1>
1C
b110 G
#960700000000
0!
0*
09
0>
0C
#960710000000
1!
1*
b111 6
19
1>
1C
b111 G
#960720000000
0!
0*
09
0>
0C
#960730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#960740000000
0!
0*
09
0>
0C
#960750000000
1!
1*
b1 6
19
1>
1C
b1 G
#960760000000
0!
0*
09
0>
0C
#960770000000
1!
1*
b10 6
19
1>
1C
b10 G
#960780000000
0!
0*
09
0>
0C
#960790000000
1!
1*
b11 6
19
1>
1C
b11 G
#960800000000
0!
0*
09
0>
0C
#960810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#960820000000
0!
0*
09
0>
0C
#960830000000
1!
1*
b101 6
19
1>
1C
b101 G
#960840000000
0!
0*
09
0>
0C
#960850000000
1!
1*
b110 6
19
1>
1C
b110 G
#960860000000
0!
0*
09
0>
0C
#960870000000
1!
1*
b111 6
19
1>
1C
b111 G
#960880000000
0!
1"
0*
1+
09
1:
0>
0C
#960890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#960900000000
0!
0*
09
0>
0C
#960910000000
1!
1*
b1 6
19
1>
1C
b1 G
#960920000000
0!
0*
09
0>
0C
#960930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#960940000000
0!
0*
09
0>
0C
#960950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#960960000000
0!
0*
09
0>
0C
#960970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#960980000000
0!
0*
09
0>
0C
#960990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#961000000000
0!
0#
0*
0,
09
0>
0?
0C
#961010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#961020000000
0!
0*
09
0>
0C
#961030000000
1!
1*
19
1>
1C
#961040000000
0!
0*
09
0>
0C
#961050000000
1!
1*
19
1>
1C
#961060000000
0!
0*
09
0>
0C
#961070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#961080000000
0!
0*
09
0>
0C
#961090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#961100000000
0!
0*
09
0>
0C
#961110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#961120000000
0!
0*
09
0>
0C
#961130000000
1!
1*
b10 6
19
1>
1C
b10 G
#961140000000
0!
0*
09
0>
0C
#961150000000
1!
1*
b11 6
19
1>
1C
b11 G
#961160000000
0!
0*
09
0>
0C
#961170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#961180000000
0!
0*
09
0>
0C
#961190000000
1!
1*
b101 6
19
1>
1C
b101 G
#961200000000
0!
0*
09
0>
0C
#961210000000
1!
1*
b110 6
19
1>
1C
b110 G
#961220000000
0!
0*
09
0>
0C
#961230000000
1!
1*
b111 6
19
1>
1C
b111 G
#961240000000
0!
0*
09
0>
0C
#961250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#961260000000
0!
0*
09
0>
0C
#961270000000
1!
1*
b1 6
19
1>
1C
b1 G
#961280000000
0!
0*
09
0>
0C
#961290000000
1!
1*
b10 6
19
1>
1C
b10 G
#961300000000
0!
0*
09
0>
0C
#961310000000
1!
1*
b11 6
19
1>
1C
b11 G
#961320000000
0!
0*
09
0>
0C
#961330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#961340000000
0!
0*
09
0>
0C
#961350000000
1!
1*
b101 6
19
1>
1C
b101 G
#961360000000
0!
0*
09
0>
0C
#961370000000
1!
1*
b110 6
19
1>
1C
b110 G
#961380000000
0!
0*
09
0>
0C
#961390000000
1!
1*
b111 6
19
1>
1C
b111 G
#961400000000
0!
0*
09
0>
0C
#961410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#961420000000
0!
0*
09
0>
0C
#961430000000
1!
1*
b1 6
19
1>
1C
b1 G
#961440000000
0!
0*
09
0>
0C
#961450000000
1!
1*
b10 6
19
1>
1C
b10 G
#961460000000
0!
0*
09
0>
0C
#961470000000
1!
1*
b11 6
19
1>
1C
b11 G
#961480000000
0!
0*
09
0>
0C
#961490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#961500000000
0!
0*
09
0>
0C
#961510000000
1!
1*
b101 6
19
1>
1C
b101 G
#961520000000
0!
0*
09
0>
0C
#961530000000
1!
1*
b110 6
19
1>
1C
b110 G
#961540000000
0!
0*
09
0>
0C
#961550000000
1!
1*
b111 6
19
1>
1C
b111 G
#961560000000
0!
1"
0*
1+
09
1:
0>
0C
#961570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#961580000000
0!
0*
09
0>
0C
#961590000000
1!
1*
b1 6
19
1>
1C
b1 G
#961600000000
0!
0*
09
0>
0C
#961610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#961620000000
0!
0*
09
0>
0C
#961630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#961640000000
0!
0*
09
0>
0C
#961650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#961660000000
0!
0*
09
0>
0C
#961670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#961680000000
0!
0#
0*
0,
09
0>
0?
0C
#961690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#961700000000
0!
0*
09
0>
0C
#961710000000
1!
1*
19
1>
1C
#961720000000
0!
0*
09
0>
0C
#961730000000
1!
1*
19
1>
1C
#961740000000
0!
0*
09
0>
0C
#961750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#961760000000
0!
0*
09
0>
0C
#961770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#961780000000
0!
0*
09
0>
0C
#961790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#961800000000
0!
0*
09
0>
0C
#961810000000
1!
1*
b10 6
19
1>
1C
b10 G
#961820000000
0!
0*
09
0>
0C
#961830000000
1!
1*
b11 6
19
1>
1C
b11 G
#961840000000
0!
0*
09
0>
0C
#961850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#961860000000
0!
0*
09
0>
0C
#961870000000
1!
1*
b101 6
19
1>
1C
b101 G
#961880000000
0!
0*
09
0>
0C
#961890000000
1!
1*
b110 6
19
1>
1C
b110 G
#961900000000
0!
0*
09
0>
0C
#961910000000
1!
1*
b111 6
19
1>
1C
b111 G
#961920000000
0!
0*
09
0>
0C
#961930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#961940000000
0!
0*
09
0>
0C
#961950000000
1!
1*
b1 6
19
1>
1C
b1 G
#961960000000
0!
0*
09
0>
0C
#961970000000
1!
1*
b10 6
19
1>
1C
b10 G
#961980000000
0!
0*
09
0>
0C
#961990000000
1!
1*
b11 6
19
1>
1C
b11 G
#962000000000
0!
0*
09
0>
0C
#962010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#962020000000
0!
0*
09
0>
0C
#962030000000
1!
1*
b101 6
19
1>
1C
b101 G
#962040000000
0!
0*
09
0>
0C
#962050000000
1!
1*
b110 6
19
1>
1C
b110 G
#962060000000
0!
0*
09
0>
0C
#962070000000
1!
1*
b111 6
19
1>
1C
b111 G
#962080000000
0!
0*
09
0>
0C
#962090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#962100000000
0!
0*
09
0>
0C
#962110000000
1!
1*
b1 6
19
1>
1C
b1 G
#962120000000
0!
0*
09
0>
0C
#962130000000
1!
1*
b10 6
19
1>
1C
b10 G
#962140000000
0!
0*
09
0>
0C
#962150000000
1!
1*
b11 6
19
1>
1C
b11 G
#962160000000
0!
0*
09
0>
0C
#962170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#962180000000
0!
0*
09
0>
0C
#962190000000
1!
1*
b101 6
19
1>
1C
b101 G
#962200000000
0!
0*
09
0>
0C
#962210000000
1!
1*
b110 6
19
1>
1C
b110 G
#962220000000
0!
0*
09
0>
0C
#962230000000
1!
1*
b111 6
19
1>
1C
b111 G
#962240000000
0!
1"
0*
1+
09
1:
0>
0C
#962250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#962260000000
0!
0*
09
0>
0C
#962270000000
1!
1*
b1 6
19
1>
1C
b1 G
#962280000000
0!
0*
09
0>
0C
#962290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#962300000000
0!
0*
09
0>
0C
#962310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#962320000000
0!
0*
09
0>
0C
#962330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#962340000000
0!
0*
09
0>
0C
#962350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#962360000000
0!
0#
0*
0,
09
0>
0?
0C
#962370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#962380000000
0!
0*
09
0>
0C
#962390000000
1!
1*
19
1>
1C
#962400000000
0!
0*
09
0>
0C
#962410000000
1!
1*
19
1>
1C
#962420000000
0!
0*
09
0>
0C
#962430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#962440000000
0!
0*
09
0>
0C
#962450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#962460000000
0!
0*
09
0>
0C
#962470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#962480000000
0!
0*
09
0>
0C
#962490000000
1!
1*
b10 6
19
1>
1C
b10 G
#962500000000
0!
0*
09
0>
0C
#962510000000
1!
1*
b11 6
19
1>
1C
b11 G
#962520000000
0!
0*
09
0>
0C
#962530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#962540000000
0!
0*
09
0>
0C
#962550000000
1!
1*
b101 6
19
1>
1C
b101 G
#962560000000
0!
0*
09
0>
0C
#962570000000
1!
1*
b110 6
19
1>
1C
b110 G
#962580000000
0!
0*
09
0>
0C
#962590000000
1!
1*
b111 6
19
1>
1C
b111 G
#962600000000
0!
0*
09
0>
0C
#962610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#962620000000
0!
0*
09
0>
0C
#962630000000
1!
1*
b1 6
19
1>
1C
b1 G
#962640000000
0!
0*
09
0>
0C
#962650000000
1!
1*
b10 6
19
1>
1C
b10 G
#962660000000
0!
0*
09
0>
0C
#962670000000
1!
1*
b11 6
19
1>
1C
b11 G
#962680000000
0!
0*
09
0>
0C
#962690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#962700000000
0!
0*
09
0>
0C
#962710000000
1!
1*
b101 6
19
1>
1C
b101 G
#962720000000
0!
0*
09
0>
0C
#962730000000
1!
1*
b110 6
19
1>
1C
b110 G
#962740000000
0!
0*
09
0>
0C
#962750000000
1!
1*
b111 6
19
1>
1C
b111 G
#962760000000
0!
0*
09
0>
0C
#962770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#962780000000
0!
0*
09
0>
0C
#962790000000
1!
1*
b1 6
19
1>
1C
b1 G
#962800000000
0!
0*
09
0>
0C
#962810000000
1!
1*
b10 6
19
1>
1C
b10 G
#962820000000
0!
0*
09
0>
0C
#962830000000
1!
1*
b11 6
19
1>
1C
b11 G
#962840000000
0!
0*
09
0>
0C
#962850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#962860000000
0!
0*
09
0>
0C
#962870000000
1!
1*
b101 6
19
1>
1C
b101 G
#962880000000
0!
0*
09
0>
0C
#962890000000
1!
1*
b110 6
19
1>
1C
b110 G
#962900000000
0!
0*
09
0>
0C
#962910000000
1!
1*
b111 6
19
1>
1C
b111 G
#962920000000
0!
1"
0*
1+
09
1:
0>
0C
#962930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#962940000000
0!
0*
09
0>
0C
#962950000000
1!
1*
b1 6
19
1>
1C
b1 G
#962960000000
0!
0*
09
0>
0C
#962970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#962980000000
0!
0*
09
0>
0C
#962990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#963000000000
0!
0*
09
0>
0C
#963010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#963020000000
0!
0*
09
0>
0C
#963030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#963040000000
0!
0#
0*
0,
09
0>
0?
0C
#963050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#963060000000
0!
0*
09
0>
0C
#963070000000
1!
1*
19
1>
1C
#963080000000
0!
0*
09
0>
0C
#963090000000
1!
1*
19
1>
1C
#963100000000
0!
0*
09
0>
0C
#963110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#963120000000
0!
0*
09
0>
0C
#963130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#963140000000
0!
0*
09
0>
0C
#963150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#963160000000
0!
0*
09
0>
0C
#963170000000
1!
1*
b10 6
19
1>
1C
b10 G
#963180000000
0!
0*
09
0>
0C
#963190000000
1!
1*
b11 6
19
1>
1C
b11 G
#963200000000
0!
0*
09
0>
0C
#963210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#963220000000
0!
0*
09
0>
0C
#963230000000
1!
1*
b101 6
19
1>
1C
b101 G
#963240000000
0!
0*
09
0>
0C
#963250000000
1!
1*
b110 6
19
1>
1C
b110 G
#963260000000
0!
0*
09
0>
0C
#963270000000
1!
1*
b111 6
19
1>
1C
b111 G
#963280000000
0!
0*
09
0>
0C
#963290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#963300000000
0!
0*
09
0>
0C
#963310000000
1!
1*
b1 6
19
1>
1C
b1 G
#963320000000
0!
0*
09
0>
0C
#963330000000
1!
1*
b10 6
19
1>
1C
b10 G
#963340000000
0!
0*
09
0>
0C
#963350000000
1!
1*
b11 6
19
1>
1C
b11 G
#963360000000
0!
0*
09
0>
0C
#963370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#963380000000
0!
0*
09
0>
0C
#963390000000
1!
1*
b101 6
19
1>
1C
b101 G
#963400000000
0!
0*
09
0>
0C
#963410000000
1!
1*
b110 6
19
1>
1C
b110 G
#963420000000
0!
0*
09
0>
0C
#963430000000
1!
1*
b111 6
19
1>
1C
b111 G
#963440000000
0!
0*
09
0>
0C
#963450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#963460000000
0!
0*
09
0>
0C
#963470000000
1!
1*
b1 6
19
1>
1C
b1 G
#963480000000
0!
0*
09
0>
0C
#963490000000
1!
1*
b10 6
19
1>
1C
b10 G
#963500000000
0!
0*
09
0>
0C
#963510000000
1!
1*
b11 6
19
1>
1C
b11 G
#963520000000
0!
0*
09
0>
0C
#963530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#963540000000
0!
0*
09
0>
0C
#963550000000
1!
1*
b101 6
19
1>
1C
b101 G
#963560000000
0!
0*
09
0>
0C
#963570000000
1!
1*
b110 6
19
1>
1C
b110 G
#963580000000
0!
0*
09
0>
0C
#963590000000
1!
1*
b111 6
19
1>
1C
b111 G
#963600000000
0!
1"
0*
1+
09
1:
0>
0C
#963610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#963620000000
0!
0*
09
0>
0C
#963630000000
1!
1*
b1 6
19
1>
1C
b1 G
#963640000000
0!
0*
09
0>
0C
#963650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#963660000000
0!
0*
09
0>
0C
#963670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#963680000000
0!
0*
09
0>
0C
#963690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#963700000000
0!
0*
09
0>
0C
#963710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#963720000000
0!
0#
0*
0,
09
0>
0?
0C
#963730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#963740000000
0!
0*
09
0>
0C
#963750000000
1!
1*
19
1>
1C
#963760000000
0!
0*
09
0>
0C
#963770000000
1!
1*
19
1>
1C
#963780000000
0!
0*
09
0>
0C
#963790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#963800000000
0!
0*
09
0>
0C
#963810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#963820000000
0!
0*
09
0>
0C
#963830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#963840000000
0!
0*
09
0>
0C
#963850000000
1!
1*
b10 6
19
1>
1C
b10 G
#963860000000
0!
0*
09
0>
0C
#963870000000
1!
1*
b11 6
19
1>
1C
b11 G
#963880000000
0!
0*
09
0>
0C
#963890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#963900000000
0!
0*
09
0>
0C
#963910000000
1!
1*
b101 6
19
1>
1C
b101 G
#963920000000
0!
0*
09
0>
0C
#963930000000
1!
1*
b110 6
19
1>
1C
b110 G
#963940000000
0!
0*
09
0>
0C
#963950000000
1!
1*
b111 6
19
1>
1C
b111 G
#963960000000
0!
0*
09
0>
0C
#963970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#963980000000
0!
0*
09
0>
0C
#963990000000
1!
1*
b1 6
19
1>
1C
b1 G
#964000000000
0!
0*
09
0>
0C
#964010000000
1!
1*
b10 6
19
1>
1C
b10 G
#964020000000
0!
0*
09
0>
0C
#964030000000
1!
1*
b11 6
19
1>
1C
b11 G
#964040000000
0!
0*
09
0>
0C
#964050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#964060000000
0!
0*
09
0>
0C
#964070000000
1!
1*
b101 6
19
1>
1C
b101 G
#964080000000
0!
0*
09
0>
0C
#964090000000
1!
1*
b110 6
19
1>
1C
b110 G
#964100000000
0!
0*
09
0>
0C
#964110000000
1!
1*
b111 6
19
1>
1C
b111 G
#964120000000
0!
0*
09
0>
0C
#964130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#964140000000
0!
0*
09
0>
0C
#964150000000
1!
1*
b1 6
19
1>
1C
b1 G
#964160000000
0!
0*
09
0>
0C
#964170000000
1!
1*
b10 6
19
1>
1C
b10 G
#964180000000
0!
0*
09
0>
0C
#964190000000
1!
1*
b11 6
19
1>
1C
b11 G
#964200000000
0!
0*
09
0>
0C
#964210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#964220000000
0!
0*
09
0>
0C
#964230000000
1!
1*
b101 6
19
1>
1C
b101 G
#964240000000
0!
0*
09
0>
0C
#964250000000
1!
1*
b110 6
19
1>
1C
b110 G
#964260000000
0!
0*
09
0>
0C
#964270000000
1!
1*
b111 6
19
1>
1C
b111 G
#964280000000
0!
1"
0*
1+
09
1:
0>
0C
#964290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#964300000000
0!
0*
09
0>
0C
#964310000000
1!
1*
b1 6
19
1>
1C
b1 G
#964320000000
0!
0*
09
0>
0C
#964330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#964340000000
0!
0*
09
0>
0C
#964350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#964360000000
0!
0*
09
0>
0C
#964370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#964380000000
0!
0*
09
0>
0C
#964390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#964400000000
0!
0#
0*
0,
09
0>
0?
0C
#964410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#964420000000
0!
0*
09
0>
0C
#964430000000
1!
1*
19
1>
1C
#964440000000
0!
0*
09
0>
0C
#964450000000
1!
1*
19
1>
1C
#964460000000
0!
0*
09
0>
0C
#964470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#964480000000
0!
0*
09
0>
0C
#964490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#964500000000
0!
0*
09
0>
0C
#964510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#964520000000
0!
0*
09
0>
0C
#964530000000
1!
1*
b10 6
19
1>
1C
b10 G
#964540000000
0!
0*
09
0>
0C
#964550000000
1!
1*
b11 6
19
1>
1C
b11 G
#964560000000
0!
0*
09
0>
0C
#964570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#964580000000
0!
0*
09
0>
0C
#964590000000
1!
1*
b101 6
19
1>
1C
b101 G
#964600000000
0!
0*
09
0>
0C
#964610000000
1!
1*
b110 6
19
1>
1C
b110 G
#964620000000
0!
0*
09
0>
0C
#964630000000
1!
1*
b111 6
19
1>
1C
b111 G
#964640000000
0!
0*
09
0>
0C
#964650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#964660000000
0!
0*
09
0>
0C
#964670000000
1!
1*
b1 6
19
1>
1C
b1 G
#964680000000
0!
0*
09
0>
0C
#964690000000
1!
1*
b10 6
19
1>
1C
b10 G
#964700000000
0!
0*
09
0>
0C
#964710000000
1!
1*
b11 6
19
1>
1C
b11 G
#964720000000
0!
0*
09
0>
0C
#964730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#964740000000
0!
0*
09
0>
0C
#964750000000
1!
1*
b101 6
19
1>
1C
b101 G
#964760000000
0!
0*
09
0>
0C
#964770000000
1!
1*
b110 6
19
1>
1C
b110 G
#964780000000
0!
0*
09
0>
0C
#964790000000
1!
1*
b111 6
19
1>
1C
b111 G
#964800000000
0!
0*
09
0>
0C
#964810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#964820000000
0!
0*
09
0>
0C
#964830000000
1!
1*
b1 6
19
1>
1C
b1 G
#964840000000
0!
0*
09
0>
0C
#964850000000
1!
1*
b10 6
19
1>
1C
b10 G
#964860000000
0!
0*
09
0>
0C
#964870000000
1!
1*
b11 6
19
1>
1C
b11 G
#964880000000
0!
0*
09
0>
0C
#964890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#964900000000
0!
0*
09
0>
0C
#964910000000
1!
1*
b101 6
19
1>
1C
b101 G
#964920000000
0!
0*
09
0>
0C
#964930000000
1!
1*
b110 6
19
1>
1C
b110 G
#964940000000
0!
0*
09
0>
0C
#964950000000
1!
1*
b111 6
19
1>
1C
b111 G
#964960000000
0!
1"
0*
1+
09
1:
0>
0C
#964970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#964980000000
0!
0*
09
0>
0C
#964990000000
1!
1*
b1 6
19
1>
1C
b1 G
#965000000000
0!
0*
09
0>
0C
#965010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#965020000000
0!
0*
09
0>
0C
#965030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#965040000000
0!
0*
09
0>
0C
#965050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#965060000000
0!
0*
09
0>
0C
#965070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#965080000000
0!
0#
0*
0,
09
0>
0?
0C
#965090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#965100000000
0!
0*
09
0>
0C
#965110000000
1!
1*
19
1>
1C
#965120000000
0!
0*
09
0>
0C
#965130000000
1!
1*
19
1>
1C
#965140000000
0!
0*
09
0>
0C
#965150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#965160000000
0!
0*
09
0>
0C
#965170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#965180000000
0!
0*
09
0>
0C
#965190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#965200000000
0!
0*
09
0>
0C
#965210000000
1!
1*
b10 6
19
1>
1C
b10 G
#965220000000
0!
0*
09
0>
0C
#965230000000
1!
1*
b11 6
19
1>
1C
b11 G
#965240000000
0!
0*
09
0>
0C
#965250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#965260000000
0!
0*
09
0>
0C
#965270000000
1!
1*
b101 6
19
1>
1C
b101 G
#965280000000
0!
0*
09
0>
0C
#965290000000
1!
1*
b110 6
19
1>
1C
b110 G
#965300000000
0!
0*
09
0>
0C
#965310000000
1!
1*
b111 6
19
1>
1C
b111 G
#965320000000
0!
0*
09
0>
0C
#965330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#965340000000
0!
0*
09
0>
0C
#965350000000
1!
1*
b1 6
19
1>
1C
b1 G
#965360000000
0!
0*
09
0>
0C
#965370000000
1!
1*
b10 6
19
1>
1C
b10 G
#965380000000
0!
0*
09
0>
0C
#965390000000
1!
1*
b11 6
19
1>
1C
b11 G
#965400000000
0!
0*
09
0>
0C
#965410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#965420000000
0!
0*
09
0>
0C
#965430000000
1!
1*
b101 6
19
1>
1C
b101 G
#965440000000
0!
0*
09
0>
0C
#965450000000
1!
1*
b110 6
19
1>
1C
b110 G
#965460000000
0!
0*
09
0>
0C
#965470000000
1!
1*
b111 6
19
1>
1C
b111 G
#965480000000
0!
0*
09
0>
0C
#965490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#965500000000
0!
0*
09
0>
0C
#965510000000
1!
1*
b1 6
19
1>
1C
b1 G
#965520000000
0!
0*
09
0>
0C
#965530000000
1!
1*
b10 6
19
1>
1C
b10 G
#965540000000
0!
0*
09
0>
0C
#965550000000
1!
1*
b11 6
19
1>
1C
b11 G
#965560000000
0!
0*
09
0>
0C
#965570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#965580000000
0!
0*
09
0>
0C
#965590000000
1!
1*
b101 6
19
1>
1C
b101 G
#965600000000
0!
0*
09
0>
0C
#965610000000
1!
1*
b110 6
19
1>
1C
b110 G
#965620000000
0!
0*
09
0>
0C
#965630000000
1!
1*
b111 6
19
1>
1C
b111 G
#965640000000
0!
1"
0*
1+
09
1:
0>
0C
#965650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#965660000000
0!
0*
09
0>
0C
#965670000000
1!
1*
b1 6
19
1>
1C
b1 G
#965680000000
0!
0*
09
0>
0C
#965690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#965700000000
0!
0*
09
0>
0C
#965710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#965720000000
0!
0*
09
0>
0C
#965730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#965740000000
0!
0*
09
0>
0C
#965750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#965760000000
0!
0#
0*
0,
09
0>
0?
0C
#965770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#965780000000
0!
0*
09
0>
0C
#965790000000
1!
1*
19
1>
1C
#965800000000
0!
0*
09
0>
0C
#965810000000
1!
1*
19
1>
1C
#965820000000
0!
0*
09
0>
0C
#965830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#965840000000
0!
0*
09
0>
0C
#965850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#965860000000
0!
0*
09
0>
0C
#965870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#965880000000
0!
0*
09
0>
0C
#965890000000
1!
1*
b10 6
19
1>
1C
b10 G
#965900000000
0!
0*
09
0>
0C
#965910000000
1!
1*
b11 6
19
1>
1C
b11 G
#965920000000
0!
0*
09
0>
0C
#965930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#965940000000
0!
0*
09
0>
0C
#965950000000
1!
1*
b101 6
19
1>
1C
b101 G
#965960000000
0!
0*
09
0>
0C
#965970000000
1!
1*
b110 6
19
1>
1C
b110 G
#965980000000
0!
0*
09
0>
0C
#965990000000
1!
1*
b111 6
19
1>
1C
b111 G
#966000000000
0!
0*
09
0>
0C
#966010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#966020000000
0!
0*
09
0>
0C
#966030000000
1!
1*
b1 6
19
1>
1C
b1 G
#966040000000
0!
0*
09
0>
0C
#966050000000
1!
1*
b10 6
19
1>
1C
b10 G
#966060000000
0!
0*
09
0>
0C
#966070000000
1!
1*
b11 6
19
1>
1C
b11 G
#966080000000
0!
0*
09
0>
0C
#966090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#966100000000
0!
0*
09
0>
0C
#966110000000
1!
1*
b101 6
19
1>
1C
b101 G
#966120000000
0!
0*
09
0>
0C
#966130000000
1!
1*
b110 6
19
1>
1C
b110 G
#966140000000
0!
0*
09
0>
0C
#966150000000
1!
1*
b111 6
19
1>
1C
b111 G
#966160000000
0!
0*
09
0>
0C
#966170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#966180000000
0!
0*
09
0>
0C
#966190000000
1!
1*
b1 6
19
1>
1C
b1 G
#966200000000
0!
0*
09
0>
0C
#966210000000
1!
1*
b10 6
19
1>
1C
b10 G
#966220000000
0!
0*
09
0>
0C
#966230000000
1!
1*
b11 6
19
1>
1C
b11 G
#966240000000
0!
0*
09
0>
0C
#966250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#966260000000
0!
0*
09
0>
0C
#966270000000
1!
1*
b101 6
19
1>
1C
b101 G
#966280000000
0!
0*
09
0>
0C
#966290000000
1!
1*
b110 6
19
1>
1C
b110 G
#966300000000
0!
0*
09
0>
0C
#966310000000
1!
1*
b111 6
19
1>
1C
b111 G
#966320000000
0!
1"
0*
1+
09
1:
0>
0C
#966330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#966340000000
0!
0*
09
0>
0C
#966350000000
1!
1*
b1 6
19
1>
1C
b1 G
#966360000000
0!
0*
09
0>
0C
#966370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#966380000000
0!
0*
09
0>
0C
#966390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#966400000000
0!
0*
09
0>
0C
#966410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#966420000000
0!
0*
09
0>
0C
#966430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#966440000000
0!
0#
0*
0,
09
0>
0?
0C
#966450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#966460000000
0!
0*
09
0>
0C
#966470000000
1!
1*
19
1>
1C
#966480000000
0!
0*
09
0>
0C
#966490000000
1!
1*
19
1>
1C
#966500000000
0!
0*
09
0>
0C
#966510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#966520000000
0!
0*
09
0>
0C
#966530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#966540000000
0!
0*
09
0>
0C
#966550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#966560000000
0!
0*
09
0>
0C
#966570000000
1!
1*
b10 6
19
1>
1C
b10 G
#966580000000
0!
0*
09
0>
0C
#966590000000
1!
1*
b11 6
19
1>
1C
b11 G
#966600000000
0!
0*
09
0>
0C
#966610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#966620000000
0!
0*
09
0>
0C
#966630000000
1!
1*
b101 6
19
1>
1C
b101 G
#966640000000
0!
0*
09
0>
0C
#966650000000
1!
1*
b110 6
19
1>
1C
b110 G
#966660000000
0!
0*
09
0>
0C
#966670000000
1!
1*
b111 6
19
1>
1C
b111 G
#966680000000
0!
0*
09
0>
0C
#966690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#966700000000
0!
0*
09
0>
0C
#966710000000
1!
1*
b1 6
19
1>
1C
b1 G
#966720000000
0!
0*
09
0>
0C
#966730000000
1!
1*
b10 6
19
1>
1C
b10 G
#966740000000
0!
0*
09
0>
0C
#966750000000
1!
1*
b11 6
19
1>
1C
b11 G
#966760000000
0!
0*
09
0>
0C
#966770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#966780000000
0!
0*
09
0>
0C
#966790000000
1!
1*
b101 6
19
1>
1C
b101 G
#966800000000
0!
0*
09
0>
0C
#966810000000
1!
1*
b110 6
19
1>
1C
b110 G
#966820000000
0!
0*
09
0>
0C
#966830000000
1!
1*
b111 6
19
1>
1C
b111 G
#966840000000
0!
0*
09
0>
0C
#966850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#966860000000
0!
0*
09
0>
0C
#966870000000
1!
1*
b1 6
19
1>
1C
b1 G
#966880000000
0!
0*
09
0>
0C
#966890000000
1!
1*
b10 6
19
1>
1C
b10 G
#966900000000
0!
0*
09
0>
0C
#966910000000
1!
1*
b11 6
19
1>
1C
b11 G
#966920000000
0!
0*
09
0>
0C
#966930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#966940000000
0!
0*
09
0>
0C
#966950000000
1!
1*
b101 6
19
1>
1C
b101 G
#966960000000
0!
0*
09
0>
0C
#966970000000
1!
1*
b110 6
19
1>
1C
b110 G
#966980000000
0!
0*
09
0>
0C
#966990000000
1!
1*
b111 6
19
1>
1C
b111 G
#967000000000
0!
1"
0*
1+
09
1:
0>
0C
#967010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#967020000000
0!
0*
09
0>
0C
#967030000000
1!
1*
b1 6
19
1>
1C
b1 G
#967040000000
0!
0*
09
0>
0C
#967050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#967060000000
0!
0*
09
0>
0C
#967070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#967080000000
0!
0*
09
0>
0C
#967090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#967100000000
0!
0*
09
0>
0C
#967110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#967120000000
0!
0#
0*
0,
09
0>
0?
0C
#967130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#967140000000
0!
0*
09
0>
0C
#967150000000
1!
1*
19
1>
1C
#967160000000
0!
0*
09
0>
0C
#967170000000
1!
1*
19
1>
1C
#967180000000
0!
0*
09
0>
0C
#967190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#967200000000
0!
0*
09
0>
0C
#967210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#967220000000
0!
0*
09
0>
0C
#967230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#967240000000
0!
0*
09
0>
0C
#967250000000
1!
1*
b10 6
19
1>
1C
b10 G
#967260000000
0!
0*
09
0>
0C
#967270000000
1!
1*
b11 6
19
1>
1C
b11 G
#967280000000
0!
0*
09
0>
0C
#967290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#967300000000
0!
0*
09
0>
0C
#967310000000
1!
1*
b101 6
19
1>
1C
b101 G
#967320000000
0!
0*
09
0>
0C
#967330000000
1!
1*
b110 6
19
1>
1C
b110 G
#967340000000
0!
0*
09
0>
0C
#967350000000
1!
1*
b111 6
19
1>
1C
b111 G
#967360000000
0!
0*
09
0>
0C
#967370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#967380000000
0!
0*
09
0>
0C
#967390000000
1!
1*
b1 6
19
1>
1C
b1 G
#967400000000
0!
0*
09
0>
0C
#967410000000
1!
1*
b10 6
19
1>
1C
b10 G
#967420000000
0!
0*
09
0>
0C
#967430000000
1!
1*
b11 6
19
1>
1C
b11 G
#967440000000
0!
0*
09
0>
0C
#967450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#967460000000
0!
0*
09
0>
0C
#967470000000
1!
1*
b101 6
19
1>
1C
b101 G
#967480000000
0!
0*
09
0>
0C
#967490000000
1!
1*
b110 6
19
1>
1C
b110 G
#967500000000
0!
0*
09
0>
0C
#967510000000
1!
1*
b111 6
19
1>
1C
b111 G
#967520000000
0!
0*
09
0>
0C
#967530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#967540000000
0!
0*
09
0>
0C
#967550000000
1!
1*
b1 6
19
1>
1C
b1 G
#967560000000
0!
0*
09
0>
0C
#967570000000
1!
1*
b10 6
19
1>
1C
b10 G
#967580000000
0!
0*
09
0>
0C
#967590000000
1!
1*
b11 6
19
1>
1C
b11 G
#967600000000
0!
0*
09
0>
0C
#967610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#967620000000
0!
0*
09
0>
0C
#967630000000
1!
1*
b101 6
19
1>
1C
b101 G
#967640000000
0!
0*
09
0>
0C
#967650000000
1!
1*
b110 6
19
1>
1C
b110 G
#967660000000
0!
0*
09
0>
0C
#967670000000
1!
1*
b111 6
19
1>
1C
b111 G
#967680000000
0!
1"
0*
1+
09
1:
0>
0C
#967690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#967700000000
0!
0*
09
0>
0C
#967710000000
1!
1*
b1 6
19
1>
1C
b1 G
#967720000000
0!
0*
09
0>
0C
#967730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#967740000000
0!
0*
09
0>
0C
#967750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#967760000000
0!
0*
09
0>
0C
#967770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#967780000000
0!
0*
09
0>
0C
#967790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#967800000000
0!
0#
0*
0,
09
0>
0?
0C
#967810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#967820000000
0!
0*
09
0>
0C
#967830000000
1!
1*
19
1>
1C
#967840000000
0!
0*
09
0>
0C
#967850000000
1!
1*
19
1>
1C
#967860000000
0!
0*
09
0>
0C
#967870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#967880000000
0!
0*
09
0>
0C
#967890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#967900000000
0!
0*
09
0>
0C
#967910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#967920000000
0!
0*
09
0>
0C
#967930000000
1!
1*
b10 6
19
1>
1C
b10 G
#967940000000
0!
0*
09
0>
0C
#967950000000
1!
1*
b11 6
19
1>
1C
b11 G
#967960000000
0!
0*
09
0>
0C
#967970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#967980000000
0!
0*
09
0>
0C
#967990000000
1!
1*
b101 6
19
1>
1C
b101 G
#968000000000
0!
0*
09
0>
0C
#968010000000
1!
1*
b110 6
19
1>
1C
b110 G
#968020000000
0!
0*
09
0>
0C
#968030000000
1!
1*
b111 6
19
1>
1C
b111 G
#968040000000
0!
0*
09
0>
0C
#968050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#968060000000
0!
0*
09
0>
0C
#968070000000
1!
1*
b1 6
19
1>
1C
b1 G
#968080000000
0!
0*
09
0>
0C
#968090000000
1!
1*
b10 6
19
1>
1C
b10 G
#968100000000
0!
0*
09
0>
0C
#968110000000
1!
1*
b11 6
19
1>
1C
b11 G
#968120000000
0!
0*
09
0>
0C
#968130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#968140000000
0!
0*
09
0>
0C
#968150000000
1!
1*
b101 6
19
1>
1C
b101 G
#968160000000
0!
0*
09
0>
0C
#968170000000
1!
1*
b110 6
19
1>
1C
b110 G
#968180000000
0!
0*
09
0>
0C
#968190000000
1!
1*
b111 6
19
1>
1C
b111 G
#968200000000
0!
0*
09
0>
0C
#968210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#968220000000
0!
0*
09
0>
0C
#968230000000
1!
1*
b1 6
19
1>
1C
b1 G
#968240000000
0!
0*
09
0>
0C
#968250000000
1!
1*
b10 6
19
1>
1C
b10 G
#968260000000
0!
0*
09
0>
0C
#968270000000
1!
1*
b11 6
19
1>
1C
b11 G
#968280000000
0!
0*
09
0>
0C
#968290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#968300000000
0!
0*
09
0>
0C
#968310000000
1!
1*
b101 6
19
1>
1C
b101 G
#968320000000
0!
0*
09
0>
0C
#968330000000
1!
1*
b110 6
19
1>
1C
b110 G
#968340000000
0!
0*
09
0>
0C
#968350000000
1!
1*
b111 6
19
1>
1C
b111 G
#968360000000
0!
1"
0*
1+
09
1:
0>
0C
#968370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#968380000000
0!
0*
09
0>
0C
#968390000000
1!
1*
b1 6
19
1>
1C
b1 G
#968400000000
0!
0*
09
0>
0C
#968410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#968420000000
0!
0*
09
0>
0C
#968430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#968440000000
0!
0*
09
0>
0C
#968450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#968460000000
0!
0*
09
0>
0C
#968470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#968480000000
0!
0#
0*
0,
09
0>
0?
0C
#968490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#968500000000
0!
0*
09
0>
0C
#968510000000
1!
1*
19
1>
1C
#968520000000
0!
0*
09
0>
0C
#968530000000
1!
1*
19
1>
1C
#968540000000
0!
0*
09
0>
0C
#968550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#968560000000
0!
0*
09
0>
0C
#968570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#968580000000
0!
0*
09
0>
0C
#968590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#968600000000
0!
0*
09
0>
0C
#968610000000
1!
1*
b10 6
19
1>
1C
b10 G
#968620000000
0!
0*
09
0>
0C
#968630000000
1!
1*
b11 6
19
1>
1C
b11 G
#968640000000
0!
0*
09
0>
0C
#968650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#968660000000
0!
0*
09
0>
0C
#968670000000
1!
1*
b101 6
19
1>
1C
b101 G
#968680000000
0!
0*
09
0>
0C
#968690000000
1!
1*
b110 6
19
1>
1C
b110 G
#968700000000
0!
0*
09
0>
0C
#968710000000
1!
1*
b111 6
19
1>
1C
b111 G
#968720000000
0!
0*
09
0>
0C
#968730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#968740000000
0!
0*
09
0>
0C
#968750000000
1!
1*
b1 6
19
1>
1C
b1 G
#968760000000
0!
0*
09
0>
0C
#968770000000
1!
1*
b10 6
19
1>
1C
b10 G
#968780000000
0!
0*
09
0>
0C
#968790000000
1!
1*
b11 6
19
1>
1C
b11 G
#968800000000
0!
0*
09
0>
0C
#968810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#968820000000
0!
0*
09
0>
0C
#968830000000
1!
1*
b101 6
19
1>
1C
b101 G
#968840000000
0!
0*
09
0>
0C
#968850000000
1!
1*
b110 6
19
1>
1C
b110 G
#968860000000
0!
0*
09
0>
0C
#968870000000
1!
1*
b111 6
19
1>
1C
b111 G
#968880000000
0!
0*
09
0>
0C
#968890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#968900000000
0!
0*
09
0>
0C
#968910000000
1!
1*
b1 6
19
1>
1C
b1 G
#968920000000
0!
0*
09
0>
0C
#968930000000
1!
1*
b10 6
19
1>
1C
b10 G
#968940000000
0!
0*
09
0>
0C
#968950000000
1!
1*
b11 6
19
1>
1C
b11 G
#968960000000
0!
0*
09
0>
0C
#968970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#968980000000
0!
0*
09
0>
0C
#968990000000
1!
1*
b101 6
19
1>
1C
b101 G
#969000000000
0!
0*
09
0>
0C
#969010000000
1!
1*
b110 6
19
1>
1C
b110 G
#969020000000
0!
0*
09
0>
0C
#969030000000
1!
1*
b111 6
19
1>
1C
b111 G
#969040000000
0!
1"
0*
1+
09
1:
0>
0C
#969050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#969060000000
0!
0*
09
0>
0C
#969070000000
1!
1*
b1 6
19
1>
1C
b1 G
#969080000000
0!
0*
09
0>
0C
#969090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#969100000000
0!
0*
09
0>
0C
#969110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#969120000000
0!
0*
09
0>
0C
#969130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#969140000000
0!
0*
09
0>
0C
#969150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#969160000000
0!
0#
0*
0,
09
0>
0?
0C
#969170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#969180000000
0!
0*
09
0>
0C
#969190000000
1!
1*
19
1>
1C
#969200000000
0!
0*
09
0>
0C
#969210000000
1!
1*
19
1>
1C
#969220000000
0!
0*
09
0>
0C
#969230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#969240000000
0!
0*
09
0>
0C
#969250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#969260000000
0!
0*
09
0>
0C
#969270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#969280000000
0!
0*
09
0>
0C
#969290000000
1!
1*
b10 6
19
1>
1C
b10 G
#969300000000
0!
0*
09
0>
0C
#969310000000
1!
1*
b11 6
19
1>
1C
b11 G
#969320000000
0!
0*
09
0>
0C
#969330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#969340000000
0!
0*
09
0>
0C
#969350000000
1!
1*
b101 6
19
1>
1C
b101 G
#969360000000
0!
0*
09
0>
0C
#969370000000
1!
1*
b110 6
19
1>
1C
b110 G
#969380000000
0!
0*
09
0>
0C
#969390000000
1!
1*
b111 6
19
1>
1C
b111 G
#969400000000
0!
0*
09
0>
0C
#969410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#969420000000
0!
0*
09
0>
0C
#969430000000
1!
1*
b1 6
19
1>
1C
b1 G
#969440000000
0!
0*
09
0>
0C
#969450000000
1!
1*
b10 6
19
1>
1C
b10 G
#969460000000
0!
0*
09
0>
0C
#969470000000
1!
1*
b11 6
19
1>
1C
b11 G
#969480000000
0!
0*
09
0>
0C
#969490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#969500000000
0!
0*
09
0>
0C
#969510000000
1!
1*
b101 6
19
1>
1C
b101 G
#969520000000
0!
0*
09
0>
0C
#969530000000
1!
1*
b110 6
19
1>
1C
b110 G
#969540000000
0!
0*
09
0>
0C
#969550000000
1!
1*
b111 6
19
1>
1C
b111 G
#969560000000
0!
0*
09
0>
0C
#969570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#969580000000
0!
0*
09
0>
0C
#969590000000
1!
1*
b1 6
19
1>
1C
b1 G
#969600000000
0!
0*
09
0>
0C
#969610000000
1!
1*
b10 6
19
1>
1C
b10 G
#969620000000
0!
0*
09
0>
0C
#969630000000
1!
1*
b11 6
19
1>
1C
b11 G
#969640000000
0!
0*
09
0>
0C
#969650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#969660000000
0!
0*
09
0>
0C
#969670000000
1!
1*
b101 6
19
1>
1C
b101 G
#969680000000
0!
0*
09
0>
0C
#969690000000
1!
1*
b110 6
19
1>
1C
b110 G
#969700000000
0!
0*
09
0>
0C
#969710000000
1!
1*
b111 6
19
1>
1C
b111 G
#969720000000
0!
1"
0*
1+
09
1:
0>
0C
#969730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#969740000000
0!
0*
09
0>
0C
#969750000000
1!
1*
b1 6
19
1>
1C
b1 G
#969760000000
0!
0*
09
0>
0C
#969770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#969780000000
0!
0*
09
0>
0C
#969790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#969800000000
0!
0*
09
0>
0C
#969810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#969820000000
0!
0*
09
0>
0C
#969830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#969840000000
0!
0#
0*
0,
09
0>
0?
0C
#969850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#969860000000
0!
0*
09
0>
0C
#969870000000
1!
1*
19
1>
1C
#969880000000
0!
0*
09
0>
0C
#969890000000
1!
1*
19
1>
1C
#969900000000
0!
0*
09
0>
0C
#969910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#969920000000
0!
0*
09
0>
0C
#969930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#969940000000
0!
0*
09
0>
0C
#969950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#969960000000
0!
0*
09
0>
0C
#969970000000
1!
1*
b10 6
19
1>
1C
b10 G
#969980000000
0!
0*
09
0>
0C
#969990000000
1!
1*
b11 6
19
1>
1C
b11 G
#970000000000
0!
0*
09
0>
0C
#970010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#970020000000
0!
0*
09
0>
0C
#970030000000
1!
1*
b101 6
19
1>
1C
b101 G
#970040000000
0!
0*
09
0>
0C
#970050000000
1!
1*
b110 6
19
1>
1C
b110 G
#970060000000
0!
0*
09
0>
0C
#970070000000
1!
1*
b111 6
19
1>
1C
b111 G
#970080000000
0!
0*
09
0>
0C
#970090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#970100000000
0!
0*
09
0>
0C
#970110000000
1!
1*
b1 6
19
1>
1C
b1 G
#970120000000
0!
0*
09
0>
0C
#970130000000
1!
1*
b10 6
19
1>
1C
b10 G
#970140000000
0!
0*
09
0>
0C
#970150000000
1!
1*
b11 6
19
1>
1C
b11 G
#970160000000
0!
0*
09
0>
0C
#970170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#970180000000
0!
0*
09
0>
0C
#970190000000
1!
1*
b101 6
19
1>
1C
b101 G
#970200000000
0!
0*
09
0>
0C
#970210000000
1!
1*
b110 6
19
1>
1C
b110 G
#970220000000
0!
0*
09
0>
0C
#970230000000
1!
1*
b111 6
19
1>
1C
b111 G
#970240000000
0!
0*
09
0>
0C
#970250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#970260000000
0!
0*
09
0>
0C
#970270000000
1!
1*
b1 6
19
1>
1C
b1 G
#970280000000
0!
0*
09
0>
0C
#970290000000
1!
1*
b10 6
19
1>
1C
b10 G
#970300000000
0!
0*
09
0>
0C
#970310000000
1!
1*
b11 6
19
1>
1C
b11 G
#970320000000
0!
0*
09
0>
0C
#970330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#970340000000
0!
0*
09
0>
0C
#970350000000
1!
1*
b101 6
19
1>
1C
b101 G
#970360000000
0!
0*
09
0>
0C
#970370000000
1!
1*
b110 6
19
1>
1C
b110 G
#970380000000
0!
0*
09
0>
0C
#970390000000
1!
1*
b111 6
19
1>
1C
b111 G
#970400000000
0!
1"
0*
1+
09
1:
0>
0C
#970410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#970420000000
0!
0*
09
0>
0C
#970430000000
1!
1*
b1 6
19
1>
1C
b1 G
#970440000000
0!
0*
09
0>
0C
#970450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#970460000000
0!
0*
09
0>
0C
#970470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#970480000000
0!
0*
09
0>
0C
#970490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#970500000000
0!
0*
09
0>
0C
#970510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#970520000000
0!
0#
0*
0,
09
0>
0?
0C
#970530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#970540000000
0!
0*
09
0>
0C
#970550000000
1!
1*
19
1>
1C
#970560000000
0!
0*
09
0>
0C
#970570000000
1!
1*
19
1>
1C
#970580000000
0!
0*
09
0>
0C
#970590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#970600000000
0!
0*
09
0>
0C
#970610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#970620000000
0!
0*
09
0>
0C
#970630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#970640000000
0!
0*
09
0>
0C
#970650000000
1!
1*
b10 6
19
1>
1C
b10 G
#970660000000
0!
0*
09
0>
0C
#970670000000
1!
1*
b11 6
19
1>
1C
b11 G
#970680000000
0!
0*
09
0>
0C
#970690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#970700000000
0!
0*
09
0>
0C
#970710000000
1!
1*
b101 6
19
1>
1C
b101 G
#970720000000
0!
0*
09
0>
0C
#970730000000
1!
1*
b110 6
19
1>
1C
b110 G
#970740000000
0!
0*
09
0>
0C
#970750000000
1!
1*
b111 6
19
1>
1C
b111 G
#970760000000
0!
0*
09
0>
0C
#970770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#970780000000
0!
0*
09
0>
0C
#970790000000
1!
1*
b1 6
19
1>
1C
b1 G
#970800000000
0!
0*
09
0>
0C
#970810000000
1!
1*
b10 6
19
1>
1C
b10 G
#970820000000
0!
0*
09
0>
0C
#970830000000
1!
1*
b11 6
19
1>
1C
b11 G
#970840000000
0!
0*
09
0>
0C
#970850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#970860000000
0!
0*
09
0>
0C
#970870000000
1!
1*
b101 6
19
1>
1C
b101 G
#970880000000
0!
0*
09
0>
0C
#970890000000
1!
1*
b110 6
19
1>
1C
b110 G
#970900000000
0!
0*
09
0>
0C
#970910000000
1!
1*
b111 6
19
1>
1C
b111 G
#970920000000
0!
0*
09
0>
0C
#970930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#970940000000
0!
0*
09
0>
0C
#970950000000
1!
1*
b1 6
19
1>
1C
b1 G
#970960000000
0!
0*
09
0>
0C
#970970000000
1!
1*
b10 6
19
1>
1C
b10 G
#970980000000
0!
0*
09
0>
0C
#970990000000
1!
1*
b11 6
19
1>
1C
b11 G
#971000000000
0!
0*
09
0>
0C
#971010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#971020000000
0!
0*
09
0>
0C
#971030000000
1!
1*
b101 6
19
1>
1C
b101 G
#971040000000
0!
0*
09
0>
0C
#971050000000
1!
1*
b110 6
19
1>
1C
b110 G
#971060000000
0!
0*
09
0>
0C
#971070000000
1!
1*
b111 6
19
1>
1C
b111 G
#971080000000
0!
1"
0*
1+
09
1:
0>
0C
#971090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#971100000000
0!
0*
09
0>
0C
#971110000000
1!
1*
b1 6
19
1>
1C
b1 G
#971120000000
0!
0*
09
0>
0C
#971130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#971140000000
0!
0*
09
0>
0C
#971150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#971160000000
0!
0*
09
0>
0C
#971170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#971180000000
0!
0*
09
0>
0C
#971190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#971200000000
0!
0#
0*
0,
09
0>
0?
0C
#971210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#971220000000
0!
0*
09
0>
0C
#971230000000
1!
1*
19
1>
1C
#971240000000
0!
0*
09
0>
0C
#971250000000
1!
1*
19
1>
1C
#971260000000
0!
0*
09
0>
0C
#971270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#971280000000
0!
0*
09
0>
0C
#971290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#971300000000
0!
0*
09
0>
0C
#971310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#971320000000
0!
0*
09
0>
0C
#971330000000
1!
1*
b10 6
19
1>
1C
b10 G
#971340000000
0!
0*
09
0>
0C
#971350000000
1!
1*
b11 6
19
1>
1C
b11 G
#971360000000
0!
0*
09
0>
0C
#971370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#971380000000
0!
0*
09
0>
0C
#971390000000
1!
1*
b101 6
19
1>
1C
b101 G
#971400000000
0!
0*
09
0>
0C
#971410000000
1!
1*
b110 6
19
1>
1C
b110 G
#971420000000
0!
0*
09
0>
0C
#971430000000
1!
1*
b111 6
19
1>
1C
b111 G
#971440000000
0!
0*
09
0>
0C
#971450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#971460000000
0!
0*
09
0>
0C
#971470000000
1!
1*
b1 6
19
1>
1C
b1 G
#971480000000
0!
0*
09
0>
0C
#971490000000
1!
1*
b10 6
19
1>
1C
b10 G
#971500000000
0!
0*
09
0>
0C
#971510000000
1!
1*
b11 6
19
1>
1C
b11 G
#971520000000
0!
0*
09
0>
0C
#971530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#971540000000
0!
0*
09
0>
0C
#971550000000
1!
1*
b101 6
19
1>
1C
b101 G
#971560000000
0!
0*
09
0>
0C
#971570000000
1!
1*
b110 6
19
1>
1C
b110 G
#971580000000
0!
0*
09
0>
0C
#971590000000
1!
1*
b111 6
19
1>
1C
b111 G
#971600000000
0!
0*
09
0>
0C
#971610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#971620000000
0!
0*
09
0>
0C
#971630000000
1!
1*
b1 6
19
1>
1C
b1 G
#971640000000
0!
0*
09
0>
0C
#971650000000
1!
1*
b10 6
19
1>
1C
b10 G
#971660000000
0!
0*
09
0>
0C
#971670000000
1!
1*
b11 6
19
1>
1C
b11 G
#971680000000
0!
0*
09
0>
0C
#971690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#971700000000
0!
0*
09
0>
0C
#971710000000
1!
1*
b101 6
19
1>
1C
b101 G
#971720000000
0!
0*
09
0>
0C
#971730000000
1!
1*
b110 6
19
1>
1C
b110 G
#971740000000
0!
0*
09
0>
0C
#971750000000
1!
1*
b111 6
19
1>
1C
b111 G
#971760000000
0!
1"
0*
1+
09
1:
0>
0C
#971770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#971780000000
0!
0*
09
0>
0C
#971790000000
1!
1*
b1 6
19
1>
1C
b1 G
#971800000000
0!
0*
09
0>
0C
#971810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#971820000000
0!
0*
09
0>
0C
#971830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#971840000000
0!
0*
09
0>
0C
#971850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#971860000000
0!
0*
09
0>
0C
#971870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#971880000000
0!
0#
0*
0,
09
0>
0?
0C
#971890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#971900000000
0!
0*
09
0>
0C
#971910000000
1!
1*
19
1>
1C
#971920000000
0!
0*
09
0>
0C
#971930000000
1!
1*
19
1>
1C
#971940000000
0!
0*
09
0>
0C
#971950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#971960000000
0!
0*
09
0>
0C
#971970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#971980000000
0!
0*
09
0>
0C
#971990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#972000000000
0!
0*
09
0>
0C
#972010000000
1!
1*
b10 6
19
1>
1C
b10 G
#972020000000
0!
0*
09
0>
0C
#972030000000
1!
1*
b11 6
19
1>
1C
b11 G
#972040000000
0!
0*
09
0>
0C
#972050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#972060000000
0!
0*
09
0>
0C
#972070000000
1!
1*
b101 6
19
1>
1C
b101 G
#972080000000
0!
0*
09
0>
0C
#972090000000
1!
1*
b110 6
19
1>
1C
b110 G
#972100000000
0!
0*
09
0>
0C
#972110000000
1!
1*
b111 6
19
1>
1C
b111 G
#972120000000
0!
0*
09
0>
0C
#972130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#972140000000
0!
0*
09
0>
0C
#972150000000
1!
1*
b1 6
19
1>
1C
b1 G
#972160000000
0!
0*
09
0>
0C
#972170000000
1!
1*
b10 6
19
1>
1C
b10 G
#972180000000
0!
0*
09
0>
0C
#972190000000
1!
1*
b11 6
19
1>
1C
b11 G
#972200000000
0!
0*
09
0>
0C
#972210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#972220000000
0!
0*
09
0>
0C
#972230000000
1!
1*
b101 6
19
1>
1C
b101 G
#972240000000
0!
0*
09
0>
0C
#972250000000
1!
1*
b110 6
19
1>
1C
b110 G
#972260000000
0!
0*
09
0>
0C
#972270000000
1!
1*
b111 6
19
1>
1C
b111 G
#972280000000
0!
0*
09
0>
0C
#972290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#972300000000
0!
0*
09
0>
0C
#972310000000
1!
1*
b1 6
19
1>
1C
b1 G
#972320000000
0!
0*
09
0>
0C
#972330000000
1!
1*
b10 6
19
1>
1C
b10 G
#972340000000
0!
0*
09
0>
0C
#972350000000
1!
1*
b11 6
19
1>
1C
b11 G
#972360000000
0!
0*
09
0>
0C
#972370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#972380000000
0!
0*
09
0>
0C
#972390000000
1!
1*
b101 6
19
1>
1C
b101 G
#972400000000
0!
0*
09
0>
0C
#972410000000
1!
1*
b110 6
19
1>
1C
b110 G
#972420000000
0!
0*
09
0>
0C
#972430000000
1!
1*
b111 6
19
1>
1C
b111 G
#972440000000
0!
1"
0*
1+
09
1:
0>
0C
#972450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#972460000000
0!
0*
09
0>
0C
#972470000000
1!
1*
b1 6
19
1>
1C
b1 G
#972480000000
0!
0*
09
0>
0C
#972490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#972500000000
0!
0*
09
0>
0C
#972510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#972520000000
0!
0*
09
0>
0C
#972530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#972540000000
0!
0*
09
0>
0C
#972550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#972560000000
0!
0#
0*
0,
09
0>
0?
0C
#972570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#972580000000
0!
0*
09
0>
0C
#972590000000
1!
1*
19
1>
1C
#972600000000
0!
0*
09
0>
0C
#972610000000
1!
1*
19
1>
1C
#972620000000
0!
0*
09
0>
0C
#972630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#972640000000
0!
0*
09
0>
0C
#972650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#972660000000
0!
0*
09
0>
0C
#972670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#972680000000
0!
0*
09
0>
0C
#972690000000
1!
1*
b10 6
19
1>
1C
b10 G
#972700000000
0!
0*
09
0>
0C
#972710000000
1!
1*
b11 6
19
1>
1C
b11 G
#972720000000
0!
0*
09
0>
0C
#972730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#972740000000
0!
0*
09
0>
0C
#972750000000
1!
1*
b101 6
19
1>
1C
b101 G
#972760000000
0!
0*
09
0>
0C
#972770000000
1!
1*
b110 6
19
1>
1C
b110 G
#972780000000
0!
0*
09
0>
0C
#972790000000
1!
1*
b111 6
19
1>
1C
b111 G
#972800000000
0!
0*
09
0>
0C
#972810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#972820000000
0!
0*
09
0>
0C
#972830000000
1!
1*
b1 6
19
1>
1C
b1 G
#972840000000
0!
0*
09
0>
0C
#972850000000
1!
1*
b10 6
19
1>
1C
b10 G
#972860000000
0!
0*
09
0>
0C
#972870000000
1!
1*
b11 6
19
1>
1C
b11 G
#972880000000
0!
0*
09
0>
0C
#972890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#972900000000
0!
0*
09
0>
0C
#972910000000
1!
1*
b101 6
19
1>
1C
b101 G
#972920000000
0!
0*
09
0>
0C
#972930000000
1!
1*
b110 6
19
1>
1C
b110 G
#972940000000
0!
0*
09
0>
0C
#972950000000
1!
1*
b111 6
19
1>
1C
b111 G
#972960000000
0!
0*
09
0>
0C
#972970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#972980000000
0!
0*
09
0>
0C
#972990000000
1!
1*
b1 6
19
1>
1C
b1 G
#973000000000
0!
0*
09
0>
0C
#973010000000
1!
1*
b10 6
19
1>
1C
b10 G
#973020000000
0!
0*
09
0>
0C
#973030000000
1!
1*
b11 6
19
1>
1C
b11 G
#973040000000
0!
0*
09
0>
0C
#973050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#973060000000
0!
0*
09
0>
0C
#973070000000
1!
1*
b101 6
19
1>
1C
b101 G
#973080000000
0!
0*
09
0>
0C
#973090000000
1!
1*
b110 6
19
1>
1C
b110 G
#973100000000
0!
0*
09
0>
0C
#973110000000
1!
1*
b111 6
19
1>
1C
b111 G
#973120000000
0!
1"
0*
1+
09
1:
0>
0C
#973130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#973140000000
0!
0*
09
0>
0C
#973150000000
1!
1*
b1 6
19
1>
1C
b1 G
#973160000000
0!
0*
09
0>
0C
#973170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#973180000000
0!
0*
09
0>
0C
#973190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#973200000000
0!
0*
09
0>
0C
#973210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#973220000000
0!
0*
09
0>
0C
#973230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#973240000000
0!
0#
0*
0,
09
0>
0?
0C
#973250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#973260000000
0!
0*
09
0>
0C
#973270000000
1!
1*
19
1>
1C
#973280000000
0!
0*
09
0>
0C
#973290000000
1!
1*
19
1>
1C
#973300000000
0!
0*
09
0>
0C
#973310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#973320000000
0!
0*
09
0>
0C
#973330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#973340000000
0!
0*
09
0>
0C
#973350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#973360000000
0!
0*
09
0>
0C
#973370000000
1!
1*
b10 6
19
1>
1C
b10 G
#973380000000
0!
0*
09
0>
0C
#973390000000
1!
1*
b11 6
19
1>
1C
b11 G
#973400000000
0!
0*
09
0>
0C
#973410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#973420000000
0!
0*
09
0>
0C
#973430000000
1!
1*
b101 6
19
1>
1C
b101 G
#973440000000
0!
0*
09
0>
0C
#973450000000
1!
1*
b110 6
19
1>
1C
b110 G
#973460000000
0!
0*
09
0>
0C
#973470000000
1!
1*
b111 6
19
1>
1C
b111 G
#973480000000
0!
0*
09
0>
0C
#973490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#973500000000
0!
0*
09
0>
0C
#973510000000
1!
1*
b1 6
19
1>
1C
b1 G
#973520000000
0!
0*
09
0>
0C
#973530000000
1!
1*
b10 6
19
1>
1C
b10 G
#973540000000
0!
0*
09
0>
0C
#973550000000
1!
1*
b11 6
19
1>
1C
b11 G
#973560000000
0!
0*
09
0>
0C
#973570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#973580000000
0!
0*
09
0>
0C
#973590000000
1!
1*
b101 6
19
1>
1C
b101 G
#973600000000
0!
0*
09
0>
0C
#973610000000
1!
1*
b110 6
19
1>
1C
b110 G
#973620000000
0!
0*
09
0>
0C
#973630000000
1!
1*
b111 6
19
1>
1C
b111 G
#973640000000
0!
0*
09
0>
0C
#973650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#973660000000
0!
0*
09
0>
0C
#973670000000
1!
1*
b1 6
19
1>
1C
b1 G
#973680000000
0!
0*
09
0>
0C
#973690000000
1!
1*
b10 6
19
1>
1C
b10 G
#973700000000
0!
0*
09
0>
0C
#973710000000
1!
1*
b11 6
19
1>
1C
b11 G
#973720000000
0!
0*
09
0>
0C
#973730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#973740000000
0!
0*
09
0>
0C
#973750000000
1!
1*
b101 6
19
1>
1C
b101 G
#973760000000
0!
0*
09
0>
0C
#973770000000
1!
1*
b110 6
19
1>
1C
b110 G
#973780000000
0!
0*
09
0>
0C
#973790000000
1!
1*
b111 6
19
1>
1C
b111 G
#973800000000
0!
1"
0*
1+
09
1:
0>
0C
#973810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#973820000000
0!
0*
09
0>
0C
#973830000000
1!
1*
b1 6
19
1>
1C
b1 G
#973840000000
0!
0*
09
0>
0C
#973850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#973860000000
0!
0*
09
0>
0C
#973870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#973880000000
0!
0*
09
0>
0C
#973890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#973900000000
0!
0*
09
0>
0C
#973910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#973920000000
0!
0#
0*
0,
09
0>
0?
0C
#973930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#973940000000
0!
0*
09
0>
0C
#973950000000
1!
1*
19
1>
1C
#973960000000
0!
0*
09
0>
0C
#973970000000
1!
1*
19
1>
1C
#973980000000
0!
0*
09
0>
0C
#973990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#974000000000
0!
0*
09
0>
0C
#974010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#974020000000
0!
0*
09
0>
0C
#974030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#974040000000
0!
0*
09
0>
0C
#974050000000
1!
1*
b10 6
19
1>
1C
b10 G
#974060000000
0!
0*
09
0>
0C
#974070000000
1!
1*
b11 6
19
1>
1C
b11 G
#974080000000
0!
0*
09
0>
0C
#974090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#974100000000
0!
0*
09
0>
0C
#974110000000
1!
1*
b101 6
19
1>
1C
b101 G
#974120000000
0!
0*
09
0>
0C
#974130000000
1!
1*
b110 6
19
1>
1C
b110 G
#974140000000
0!
0*
09
0>
0C
#974150000000
1!
1*
b111 6
19
1>
1C
b111 G
#974160000000
0!
0*
09
0>
0C
#974170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#974180000000
0!
0*
09
0>
0C
#974190000000
1!
1*
b1 6
19
1>
1C
b1 G
#974200000000
0!
0*
09
0>
0C
#974210000000
1!
1*
b10 6
19
1>
1C
b10 G
#974220000000
0!
0*
09
0>
0C
#974230000000
1!
1*
b11 6
19
1>
1C
b11 G
#974240000000
0!
0*
09
0>
0C
#974250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#974260000000
0!
0*
09
0>
0C
#974270000000
1!
1*
b101 6
19
1>
1C
b101 G
#974280000000
0!
0*
09
0>
0C
#974290000000
1!
1*
b110 6
19
1>
1C
b110 G
#974300000000
0!
0*
09
0>
0C
#974310000000
1!
1*
b111 6
19
1>
1C
b111 G
#974320000000
0!
0*
09
0>
0C
#974330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#974340000000
0!
0*
09
0>
0C
#974350000000
1!
1*
b1 6
19
1>
1C
b1 G
#974360000000
0!
0*
09
0>
0C
#974370000000
1!
1*
b10 6
19
1>
1C
b10 G
#974380000000
0!
0*
09
0>
0C
#974390000000
1!
1*
b11 6
19
1>
1C
b11 G
#974400000000
0!
0*
09
0>
0C
#974410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#974420000000
0!
0*
09
0>
0C
#974430000000
1!
1*
b101 6
19
1>
1C
b101 G
#974440000000
0!
0*
09
0>
0C
#974450000000
1!
1*
b110 6
19
1>
1C
b110 G
#974460000000
0!
0*
09
0>
0C
#974470000000
1!
1*
b111 6
19
1>
1C
b111 G
#974480000000
0!
1"
0*
1+
09
1:
0>
0C
#974490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#974500000000
0!
0*
09
0>
0C
#974510000000
1!
1*
b1 6
19
1>
1C
b1 G
#974520000000
0!
0*
09
0>
0C
#974530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#974540000000
0!
0*
09
0>
0C
#974550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#974560000000
0!
0*
09
0>
0C
#974570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#974580000000
0!
0*
09
0>
0C
#974590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#974600000000
0!
0#
0*
0,
09
0>
0?
0C
#974610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#974620000000
0!
0*
09
0>
0C
#974630000000
1!
1*
19
1>
1C
#974640000000
0!
0*
09
0>
0C
#974650000000
1!
1*
19
1>
1C
#974660000000
0!
0*
09
0>
0C
#974670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#974680000000
0!
0*
09
0>
0C
#974690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#974700000000
0!
0*
09
0>
0C
#974710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#974720000000
0!
0*
09
0>
0C
#974730000000
1!
1*
b10 6
19
1>
1C
b10 G
#974740000000
0!
0*
09
0>
0C
#974750000000
1!
1*
b11 6
19
1>
1C
b11 G
#974760000000
0!
0*
09
0>
0C
#974770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#974780000000
0!
0*
09
0>
0C
#974790000000
1!
1*
b101 6
19
1>
1C
b101 G
#974800000000
0!
0*
09
0>
0C
#974810000000
1!
1*
b110 6
19
1>
1C
b110 G
#974820000000
0!
0*
09
0>
0C
#974830000000
1!
1*
b111 6
19
1>
1C
b111 G
#974840000000
0!
0*
09
0>
0C
#974850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#974860000000
0!
0*
09
0>
0C
#974870000000
1!
1*
b1 6
19
1>
1C
b1 G
#974880000000
0!
0*
09
0>
0C
#974890000000
1!
1*
b10 6
19
1>
1C
b10 G
#974900000000
0!
0*
09
0>
0C
#974910000000
1!
1*
b11 6
19
1>
1C
b11 G
#974920000000
0!
0*
09
0>
0C
#974930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#974940000000
0!
0*
09
0>
0C
#974950000000
1!
1*
b101 6
19
1>
1C
b101 G
#974960000000
0!
0*
09
0>
0C
#974970000000
1!
1*
b110 6
19
1>
1C
b110 G
#974980000000
0!
0*
09
0>
0C
#974990000000
1!
1*
b111 6
19
1>
1C
b111 G
#975000000000
0!
0*
09
0>
0C
#975010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#975020000000
0!
0*
09
0>
0C
#975030000000
1!
1*
b1 6
19
1>
1C
b1 G
#975040000000
0!
0*
09
0>
0C
#975050000000
1!
1*
b10 6
19
1>
1C
b10 G
#975060000000
0!
0*
09
0>
0C
#975070000000
1!
1*
b11 6
19
1>
1C
b11 G
#975080000000
0!
0*
09
0>
0C
#975090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#975100000000
0!
0*
09
0>
0C
#975110000000
1!
1*
b101 6
19
1>
1C
b101 G
#975120000000
0!
0*
09
0>
0C
#975130000000
1!
1*
b110 6
19
1>
1C
b110 G
#975140000000
0!
0*
09
0>
0C
#975150000000
1!
1*
b111 6
19
1>
1C
b111 G
#975160000000
0!
1"
0*
1+
09
1:
0>
0C
#975170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#975180000000
0!
0*
09
0>
0C
#975190000000
1!
1*
b1 6
19
1>
1C
b1 G
#975200000000
0!
0*
09
0>
0C
#975210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#975220000000
0!
0*
09
0>
0C
#975230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#975240000000
0!
0*
09
0>
0C
#975250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#975260000000
0!
0*
09
0>
0C
#975270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#975280000000
0!
0#
0*
0,
09
0>
0?
0C
#975290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#975300000000
0!
0*
09
0>
0C
#975310000000
1!
1*
19
1>
1C
#975320000000
0!
0*
09
0>
0C
#975330000000
1!
1*
19
1>
1C
#975340000000
0!
0*
09
0>
0C
#975350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#975360000000
0!
0*
09
0>
0C
#975370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#975380000000
0!
0*
09
0>
0C
#975390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#975400000000
0!
0*
09
0>
0C
#975410000000
1!
1*
b10 6
19
1>
1C
b10 G
#975420000000
0!
0*
09
0>
0C
#975430000000
1!
1*
b11 6
19
1>
1C
b11 G
#975440000000
0!
0*
09
0>
0C
#975450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#975460000000
0!
0*
09
0>
0C
#975470000000
1!
1*
b101 6
19
1>
1C
b101 G
#975480000000
0!
0*
09
0>
0C
#975490000000
1!
1*
b110 6
19
1>
1C
b110 G
#975500000000
0!
0*
09
0>
0C
#975510000000
1!
1*
b111 6
19
1>
1C
b111 G
#975520000000
0!
0*
09
0>
0C
#975530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#975540000000
0!
0*
09
0>
0C
#975550000000
1!
1*
b1 6
19
1>
1C
b1 G
#975560000000
0!
0*
09
0>
0C
#975570000000
1!
1*
b10 6
19
1>
1C
b10 G
#975580000000
0!
0*
09
0>
0C
#975590000000
1!
1*
b11 6
19
1>
1C
b11 G
#975600000000
0!
0*
09
0>
0C
#975610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#975620000000
0!
0*
09
0>
0C
#975630000000
1!
1*
b101 6
19
1>
1C
b101 G
#975640000000
0!
0*
09
0>
0C
#975650000000
1!
1*
b110 6
19
1>
1C
b110 G
#975660000000
0!
0*
09
0>
0C
#975670000000
1!
1*
b111 6
19
1>
1C
b111 G
#975680000000
0!
0*
09
0>
0C
#975690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#975700000000
0!
0*
09
0>
0C
#975710000000
1!
1*
b1 6
19
1>
1C
b1 G
#975720000000
0!
0*
09
0>
0C
#975730000000
1!
1*
b10 6
19
1>
1C
b10 G
#975740000000
0!
0*
09
0>
0C
#975750000000
1!
1*
b11 6
19
1>
1C
b11 G
#975760000000
0!
0*
09
0>
0C
#975770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#975780000000
0!
0*
09
0>
0C
#975790000000
1!
1*
b101 6
19
1>
1C
b101 G
#975800000000
0!
0*
09
0>
0C
#975810000000
1!
1*
b110 6
19
1>
1C
b110 G
#975820000000
0!
0*
09
0>
0C
#975830000000
1!
1*
b111 6
19
1>
1C
b111 G
#975840000000
0!
1"
0*
1+
09
1:
0>
0C
#975850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#975860000000
0!
0*
09
0>
0C
#975870000000
1!
1*
b1 6
19
1>
1C
b1 G
#975880000000
0!
0*
09
0>
0C
#975890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#975900000000
0!
0*
09
0>
0C
#975910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#975920000000
0!
0*
09
0>
0C
#975930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#975940000000
0!
0*
09
0>
0C
#975950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#975960000000
0!
0#
0*
0,
09
0>
0?
0C
#975970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#975980000000
0!
0*
09
0>
0C
#975990000000
1!
1*
19
1>
1C
#976000000000
0!
0*
09
0>
0C
#976010000000
1!
1*
19
1>
1C
#976020000000
0!
0*
09
0>
0C
#976030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#976040000000
0!
0*
09
0>
0C
#976050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#976060000000
0!
0*
09
0>
0C
#976070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#976080000000
0!
0*
09
0>
0C
#976090000000
1!
1*
b10 6
19
1>
1C
b10 G
#976100000000
0!
0*
09
0>
0C
#976110000000
1!
1*
b11 6
19
1>
1C
b11 G
#976120000000
0!
0*
09
0>
0C
#976130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#976140000000
0!
0*
09
0>
0C
#976150000000
1!
1*
b101 6
19
1>
1C
b101 G
#976160000000
0!
0*
09
0>
0C
#976170000000
1!
1*
b110 6
19
1>
1C
b110 G
#976180000000
0!
0*
09
0>
0C
#976190000000
1!
1*
b111 6
19
1>
1C
b111 G
#976200000000
0!
0*
09
0>
0C
#976210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#976220000000
0!
0*
09
0>
0C
#976230000000
1!
1*
b1 6
19
1>
1C
b1 G
#976240000000
0!
0*
09
0>
0C
#976250000000
1!
1*
b10 6
19
1>
1C
b10 G
#976260000000
0!
0*
09
0>
0C
#976270000000
1!
1*
b11 6
19
1>
1C
b11 G
#976280000000
0!
0*
09
0>
0C
#976290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#976300000000
0!
0*
09
0>
0C
#976310000000
1!
1*
b101 6
19
1>
1C
b101 G
#976320000000
0!
0*
09
0>
0C
#976330000000
1!
1*
b110 6
19
1>
1C
b110 G
#976340000000
0!
0*
09
0>
0C
#976350000000
1!
1*
b111 6
19
1>
1C
b111 G
#976360000000
0!
0*
09
0>
0C
#976370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#976380000000
0!
0*
09
0>
0C
#976390000000
1!
1*
b1 6
19
1>
1C
b1 G
#976400000000
0!
0*
09
0>
0C
#976410000000
1!
1*
b10 6
19
1>
1C
b10 G
#976420000000
0!
0*
09
0>
0C
#976430000000
1!
1*
b11 6
19
1>
1C
b11 G
#976440000000
0!
0*
09
0>
0C
#976450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#976460000000
0!
0*
09
0>
0C
#976470000000
1!
1*
b101 6
19
1>
1C
b101 G
#976480000000
0!
0*
09
0>
0C
#976490000000
1!
1*
b110 6
19
1>
1C
b110 G
#976500000000
0!
0*
09
0>
0C
#976510000000
1!
1*
b111 6
19
1>
1C
b111 G
#976520000000
0!
1"
0*
1+
09
1:
0>
0C
#976530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#976540000000
0!
0*
09
0>
0C
#976550000000
1!
1*
b1 6
19
1>
1C
b1 G
#976560000000
0!
0*
09
0>
0C
#976570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#976580000000
0!
0*
09
0>
0C
#976590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#976600000000
0!
0*
09
0>
0C
#976610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#976620000000
0!
0*
09
0>
0C
#976630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#976640000000
0!
0#
0*
0,
09
0>
0?
0C
#976650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#976660000000
0!
0*
09
0>
0C
#976670000000
1!
1*
19
1>
1C
#976680000000
0!
0*
09
0>
0C
#976690000000
1!
1*
19
1>
1C
#976700000000
0!
0*
09
0>
0C
#976710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#976720000000
0!
0*
09
0>
0C
#976730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#976740000000
0!
0*
09
0>
0C
#976750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#976760000000
0!
0*
09
0>
0C
#976770000000
1!
1*
b10 6
19
1>
1C
b10 G
#976780000000
0!
0*
09
0>
0C
#976790000000
1!
1*
b11 6
19
1>
1C
b11 G
#976800000000
0!
0*
09
0>
0C
#976810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#976820000000
0!
0*
09
0>
0C
#976830000000
1!
1*
b101 6
19
1>
1C
b101 G
#976840000000
0!
0*
09
0>
0C
#976850000000
1!
1*
b110 6
19
1>
1C
b110 G
#976860000000
0!
0*
09
0>
0C
#976870000000
1!
1*
b111 6
19
1>
1C
b111 G
#976880000000
0!
0*
09
0>
0C
#976890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#976900000000
0!
0*
09
0>
0C
#976910000000
1!
1*
b1 6
19
1>
1C
b1 G
#976920000000
0!
0*
09
0>
0C
#976930000000
1!
1*
b10 6
19
1>
1C
b10 G
#976940000000
0!
0*
09
0>
0C
#976950000000
1!
1*
b11 6
19
1>
1C
b11 G
#976960000000
0!
0*
09
0>
0C
#976970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#976980000000
0!
0*
09
0>
0C
#976990000000
1!
1*
b101 6
19
1>
1C
b101 G
#977000000000
0!
0*
09
0>
0C
#977010000000
1!
1*
b110 6
19
1>
1C
b110 G
#977020000000
0!
0*
09
0>
0C
#977030000000
1!
1*
b111 6
19
1>
1C
b111 G
#977040000000
0!
0*
09
0>
0C
#977050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#977060000000
0!
0*
09
0>
0C
#977070000000
1!
1*
b1 6
19
1>
1C
b1 G
#977080000000
0!
0*
09
0>
0C
#977090000000
1!
1*
b10 6
19
1>
1C
b10 G
#977100000000
0!
0*
09
0>
0C
#977110000000
1!
1*
b11 6
19
1>
1C
b11 G
#977120000000
0!
0*
09
0>
0C
#977130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#977140000000
0!
0*
09
0>
0C
#977150000000
1!
1*
b101 6
19
1>
1C
b101 G
#977160000000
0!
0*
09
0>
0C
#977170000000
1!
1*
b110 6
19
1>
1C
b110 G
#977180000000
0!
0*
09
0>
0C
#977190000000
1!
1*
b111 6
19
1>
1C
b111 G
#977200000000
0!
1"
0*
1+
09
1:
0>
0C
#977210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#977220000000
0!
0*
09
0>
0C
#977230000000
1!
1*
b1 6
19
1>
1C
b1 G
#977240000000
0!
0*
09
0>
0C
#977250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#977260000000
0!
0*
09
0>
0C
#977270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#977280000000
0!
0*
09
0>
0C
#977290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#977300000000
0!
0*
09
0>
0C
#977310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#977320000000
0!
0#
0*
0,
09
0>
0?
0C
#977330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#977340000000
0!
0*
09
0>
0C
#977350000000
1!
1*
19
1>
1C
#977360000000
0!
0*
09
0>
0C
#977370000000
1!
1*
19
1>
1C
#977380000000
0!
0*
09
0>
0C
#977390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#977400000000
0!
0*
09
0>
0C
#977410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#977420000000
0!
0*
09
0>
0C
#977430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#977440000000
0!
0*
09
0>
0C
#977450000000
1!
1*
b10 6
19
1>
1C
b10 G
#977460000000
0!
0*
09
0>
0C
#977470000000
1!
1*
b11 6
19
1>
1C
b11 G
#977480000000
0!
0*
09
0>
0C
#977490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#977500000000
0!
0*
09
0>
0C
#977510000000
1!
1*
b101 6
19
1>
1C
b101 G
#977520000000
0!
0*
09
0>
0C
#977530000000
1!
1*
b110 6
19
1>
1C
b110 G
#977540000000
0!
0*
09
0>
0C
#977550000000
1!
1*
b111 6
19
1>
1C
b111 G
#977560000000
0!
0*
09
0>
0C
#977570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#977580000000
0!
0*
09
0>
0C
#977590000000
1!
1*
b1 6
19
1>
1C
b1 G
#977600000000
0!
0*
09
0>
0C
#977610000000
1!
1*
b10 6
19
1>
1C
b10 G
#977620000000
0!
0*
09
0>
0C
#977630000000
1!
1*
b11 6
19
1>
1C
b11 G
#977640000000
0!
0*
09
0>
0C
#977650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#977660000000
0!
0*
09
0>
0C
#977670000000
1!
1*
b101 6
19
1>
1C
b101 G
#977680000000
0!
0*
09
0>
0C
#977690000000
1!
1*
b110 6
19
1>
1C
b110 G
#977700000000
0!
0*
09
0>
0C
#977710000000
1!
1*
b111 6
19
1>
1C
b111 G
#977720000000
0!
0*
09
0>
0C
#977730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#977740000000
0!
0*
09
0>
0C
#977750000000
1!
1*
b1 6
19
1>
1C
b1 G
#977760000000
0!
0*
09
0>
0C
#977770000000
1!
1*
b10 6
19
1>
1C
b10 G
#977780000000
0!
0*
09
0>
0C
#977790000000
1!
1*
b11 6
19
1>
1C
b11 G
#977800000000
0!
0*
09
0>
0C
#977810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#977820000000
0!
0*
09
0>
0C
#977830000000
1!
1*
b101 6
19
1>
1C
b101 G
#977840000000
0!
0*
09
0>
0C
#977850000000
1!
1*
b110 6
19
1>
1C
b110 G
#977860000000
0!
0*
09
0>
0C
#977870000000
1!
1*
b111 6
19
1>
1C
b111 G
#977880000000
0!
1"
0*
1+
09
1:
0>
0C
#977890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#977900000000
0!
0*
09
0>
0C
#977910000000
1!
1*
b1 6
19
1>
1C
b1 G
#977920000000
0!
0*
09
0>
0C
#977930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#977940000000
0!
0*
09
0>
0C
#977950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#977960000000
0!
0*
09
0>
0C
#977970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#977980000000
0!
0*
09
0>
0C
#977990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#978000000000
0!
0#
0*
0,
09
0>
0?
0C
#978010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#978020000000
0!
0*
09
0>
0C
#978030000000
1!
1*
19
1>
1C
#978040000000
0!
0*
09
0>
0C
#978050000000
1!
1*
19
1>
1C
#978060000000
0!
0*
09
0>
0C
#978070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#978080000000
0!
0*
09
0>
0C
#978090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#978100000000
0!
0*
09
0>
0C
#978110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#978120000000
0!
0*
09
0>
0C
#978130000000
1!
1*
b10 6
19
1>
1C
b10 G
#978140000000
0!
0*
09
0>
0C
#978150000000
1!
1*
b11 6
19
1>
1C
b11 G
#978160000000
0!
0*
09
0>
0C
#978170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#978180000000
0!
0*
09
0>
0C
#978190000000
1!
1*
b101 6
19
1>
1C
b101 G
#978200000000
0!
0*
09
0>
0C
#978210000000
1!
1*
b110 6
19
1>
1C
b110 G
#978220000000
0!
0*
09
0>
0C
#978230000000
1!
1*
b111 6
19
1>
1C
b111 G
#978240000000
0!
0*
09
0>
0C
#978250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#978260000000
0!
0*
09
0>
0C
#978270000000
1!
1*
b1 6
19
1>
1C
b1 G
#978280000000
0!
0*
09
0>
0C
#978290000000
1!
1*
b10 6
19
1>
1C
b10 G
#978300000000
0!
0*
09
0>
0C
#978310000000
1!
1*
b11 6
19
1>
1C
b11 G
#978320000000
0!
0*
09
0>
0C
#978330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#978340000000
0!
0*
09
0>
0C
#978350000000
1!
1*
b101 6
19
1>
1C
b101 G
#978360000000
0!
0*
09
0>
0C
#978370000000
1!
1*
b110 6
19
1>
1C
b110 G
#978380000000
0!
0*
09
0>
0C
#978390000000
1!
1*
b111 6
19
1>
1C
b111 G
#978400000000
0!
0*
09
0>
0C
#978410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#978420000000
0!
0*
09
0>
0C
#978430000000
1!
1*
b1 6
19
1>
1C
b1 G
#978440000000
0!
0*
09
0>
0C
#978450000000
1!
1*
b10 6
19
1>
1C
b10 G
#978460000000
0!
0*
09
0>
0C
#978470000000
1!
1*
b11 6
19
1>
1C
b11 G
#978480000000
0!
0*
09
0>
0C
#978490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#978500000000
0!
0*
09
0>
0C
#978510000000
1!
1*
b101 6
19
1>
1C
b101 G
#978520000000
0!
0*
09
0>
0C
#978530000000
1!
1*
b110 6
19
1>
1C
b110 G
#978540000000
0!
0*
09
0>
0C
#978550000000
1!
1*
b111 6
19
1>
1C
b111 G
#978560000000
0!
1"
0*
1+
09
1:
0>
0C
#978570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#978580000000
0!
0*
09
0>
0C
#978590000000
1!
1*
b1 6
19
1>
1C
b1 G
#978600000000
0!
0*
09
0>
0C
#978610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#978620000000
0!
0*
09
0>
0C
#978630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#978640000000
0!
0*
09
0>
0C
#978650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#978660000000
0!
0*
09
0>
0C
#978670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#978680000000
0!
0#
0*
0,
09
0>
0?
0C
#978690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#978700000000
0!
0*
09
0>
0C
#978710000000
1!
1*
19
1>
1C
#978720000000
0!
0*
09
0>
0C
#978730000000
1!
1*
19
1>
1C
#978740000000
0!
0*
09
0>
0C
#978750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#978760000000
0!
0*
09
0>
0C
#978770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#978780000000
0!
0*
09
0>
0C
#978790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#978800000000
0!
0*
09
0>
0C
#978810000000
1!
1*
b10 6
19
1>
1C
b10 G
#978820000000
0!
0*
09
0>
0C
#978830000000
1!
1*
b11 6
19
1>
1C
b11 G
#978840000000
0!
0*
09
0>
0C
#978850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#978860000000
0!
0*
09
0>
0C
#978870000000
1!
1*
b101 6
19
1>
1C
b101 G
#978880000000
0!
0*
09
0>
0C
#978890000000
1!
1*
b110 6
19
1>
1C
b110 G
#978900000000
0!
0*
09
0>
0C
#978910000000
1!
1*
b111 6
19
1>
1C
b111 G
#978920000000
0!
0*
09
0>
0C
#978930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#978940000000
0!
0*
09
0>
0C
#978950000000
1!
1*
b1 6
19
1>
1C
b1 G
#978960000000
0!
0*
09
0>
0C
#978970000000
1!
1*
b10 6
19
1>
1C
b10 G
#978980000000
0!
0*
09
0>
0C
#978990000000
1!
1*
b11 6
19
1>
1C
b11 G
#979000000000
0!
0*
09
0>
0C
#979010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#979020000000
0!
0*
09
0>
0C
#979030000000
1!
1*
b101 6
19
1>
1C
b101 G
#979040000000
0!
0*
09
0>
0C
#979050000000
1!
1*
b110 6
19
1>
1C
b110 G
#979060000000
0!
0*
09
0>
0C
#979070000000
1!
1*
b111 6
19
1>
1C
b111 G
#979080000000
0!
0*
09
0>
0C
#979090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#979100000000
0!
0*
09
0>
0C
#979110000000
1!
1*
b1 6
19
1>
1C
b1 G
#979120000000
0!
0*
09
0>
0C
#979130000000
1!
1*
b10 6
19
1>
1C
b10 G
#979140000000
0!
0*
09
0>
0C
#979150000000
1!
1*
b11 6
19
1>
1C
b11 G
#979160000000
0!
0*
09
0>
0C
#979170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#979180000000
0!
0*
09
0>
0C
#979190000000
1!
1*
b101 6
19
1>
1C
b101 G
#979200000000
0!
0*
09
0>
0C
#979210000000
1!
1*
b110 6
19
1>
1C
b110 G
#979220000000
0!
0*
09
0>
0C
#979230000000
1!
1*
b111 6
19
1>
1C
b111 G
#979240000000
0!
1"
0*
1+
09
1:
0>
0C
#979250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#979260000000
0!
0*
09
0>
0C
#979270000000
1!
1*
b1 6
19
1>
1C
b1 G
#979280000000
0!
0*
09
0>
0C
#979290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#979300000000
0!
0*
09
0>
0C
#979310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#979320000000
0!
0*
09
0>
0C
#979330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#979340000000
0!
0*
09
0>
0C
#979350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#979360000000
0!
0#
0*
0,
09
0>
0?
0C
#979370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#979380000000
0!
0*
09
0>
0C
#979390000000
1!
1*
19
1>
1C
#979400000000
0!
0*
09
0>
0C
#979410000000
1!
1*
19
1>
1C
#979420000000
0!
0*
09
0>
0C
#979430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#979440000000
0!
0*
09
0>
0C
#979450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#979460000000
0!
0*
09
0>
0C
#979470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#979480000000
0!
0*
09
0>
0C
#979490000000
1!
1*
b10 6
19
1>
1C
b10 G
#979500000000
0!
0*
09
0>
0C
#979510000000
1!
1*
b11 6
19
1>
1C
b11 G
#979520000000
0!
0*
09
0>
0C
#979530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#979540000000
0!
0*
09
0>
0C
#979550000000
1!
1*
b101 6
19
1>
1C
b101 G
#979560000000
0!
0*
09
0>
0C
#979570000000
1!
1*
b110 6
19
1>
1C
b110 G
#979580000000
0!
0*
09
0>
0C
#979590000000
1!
1*
b111 6
19
1>
1C
b111 G
#979600000000
0!
0*
09
0>
0C
#979610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#979620000000
0!
0*
09
0>
0C
#979630000000
1!
1*
b1 6
19
1>
1C
b1 G
#979640000000
0!
0*
09
0>
0C
#979650000000
1!
1*
b10 6
19
1>
1C
b10 G
#979660000000
0!
0*
09
0>
0C
#979670000000
1!
1*
b11 6
19
1>
1C
b11 G
#979680000000
0!
0*
09
0>
0C
#979690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#979700000000
0!
0*
09
0>
0C
#979710000000
1!
1*
b101 6
19
1>
1C
b101 G
#979720000000
0!
0*
09
0>
0C
#979730000000
1!
1*
b110 6
19
1>
1C
b110 G
#979740000000
0!
0*
09
0>
0C
#979750000000
1!
1*
b111 6
19
1>
1C
b111 G
#979760000000
0!
0*
09
0>
0C
#979770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#979780000000
0!
0*
09
0>
0C
#979790000000
1!
1*
b1 6
19
1>
1C
b1 G
#979800000000
0!
0*
09
0>
0C
#979810000000
1!
1*
b10 6
19
1>
1C
b10 G
#979820000000
0!
0*
09
0>
0C
#979830000000
1!
1*
b11 6
19
1>
1C
b11 G
#979840000000
0!
0*
09
0>
0C
#979850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#979860000000
0!
0*
09
0>
0C
#979870000000
1!
1*
b101 6
19
1>
1C
b101 G
#979880000000
0!
0*
09
0>
0C
#979890000000
1!
1*
b110 6
19
1>
1C
b110 G
#979900000000
0!
0*
09
0>
0C
#979910000000
1!
1*
b111 6
19
1>
1C
b111 G
#979920000000
0!
1"
0*
1+
09
1:
0>
0C
#979930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#979940000000
0!
0*
09
0>
0C
#979950000000
1!
1*
b1 6
19
1>
1C
b1 G
#979960000000
0!
0*
09
0>
0C
#979970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#979980000000
0!
0*
09
0>
0C
#979990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#980000000000
0!
0*
09
0>
0C
#980010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#980020000000
0!
0*
09
0>
0C
#980030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#980040000000
0!
0#
0*
0,
09
0>
0?
0C
#980050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#980060000000
0!
0*
09
0>
0C
#980070000000
1!
1*
19
1>
1C
#980080000000
0!
0*
09
0>
0C
#980090000000
1!
1*
19
1>
1C
#980100000000
0!
0*
09
0>
0C
#980110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#980120000000
0!
0*
09
0>
0C
#980130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#980140000000
0!
0*
09
0>
0C
#980150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#980160000000
0!
0*
09
0>
0C
#980170000000
1!
1*
b10 6
19
1>
1C
b10 G
#980180000000
0!
0*
09
0>
0C
#980190000000
1!
1*
b11 6
19
1>
1C
b11 G
#980200000000
0!
0*
09
0>
0C
#980210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#980220000000
0!
0*
09
0>
0C
#980230000000
1!
1*
b101 6
19
1>
1C
b101 G
#980240000000
0!
0*
09
0>
0C
#980250000000
1!
1*
b110 6
19
1>
1C
b110 G
#980260000000
0!
0*
09
0>
0C
#980270000000
1!
1*
b111 6
19
1>
1C
b111 G
#980280000000
0!
0*
09
0>
0C
#980290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#980300000000
0!
0*
09
0>
0C
#980310000000
1!
1*
b1 6
19
1>
1C
b1 G
#980320000000
0!
0*
09
0>
0C
#980330000000
1!
1*
b10 6
19
1>
1C
b10 G
#980340000000
0!
0*
09
0>
0C
#980350000000
1!
1*
b11 6
19
1>
1C
b11 G
#980360000000
0!
0*
09
0>
0C
#980370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#980380000000
0!
0*
09
0>
0C
#980390000000
1!
1*
b101 6
19
1>
1C
b101 G
#980400000000
0!
0*
09
0>
0C
#980410000000
1!
1*
b110 6
19
1>
1C
b110 G
#980420000000
0!
0*
09
0>
0C
#980430000000
1!
1*
b111 6
19
1>
1C
b111 G
#980440000000
0!
0*
09
0>
0C
#980450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#980460000000
0!
0*
09
0>
0C
#980470000000
1!
1*
b1 6
19
1>
1C
b1 G
#980480000000
0!
0*
09
0>
0C
#980490000000
1!
1*
b10 6
19
1>
1C
b10 G
#980500000000
0!
0*
09
0>
0C
#980510000000
1!
1*
b11 6
19
1>
1C
b11 G
#980520000000
0!
0*
09
0>
0C
#980530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#980540000000
0!
0*
09
0>
0C
#980550000000
1!
1*
b101 6
19
1>
1C
b101 G
#980560000000
0!
0*
09
0>
0C
#980570000000
1!
1*
b110 6
19
1>
1C
b110 G
#980580000000
0!
0*
09
0>
0C
#980590000000
1!
1*
b111 6
19
1>
1C
b111 G
#980600000000
0!
1"
0*
1+
09
1:
0>
0C
#980610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#980620000000
0!
0*
09
0>
0C
#980630000000
1!
1*
b1 6
19
1>
1C
b1 G
#980640000000
0!
0*
09
0>
0C
#980650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#980660000000
0!
0*
09
0>
0C
#980670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#980680000000
0!
0*
09
0>
0C
#980690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#980700000000
0!
0*
09
0>
0C
#980710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#980720000000
0!
0#
0*
0,
09
0>
0?
0C
#980730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#980740000000
0!
0*
09
0>
0C
#980750000000
1!
1*
19
1>
1C
#980760000000
0!
0*
09
0>
0C
#980770000000
1!
1*
19
1>
1C
#980780000000
0!
0*
09
0>
0C
#980790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#980800000000
0!
0*
09
0>
0C
#980810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#980820000000
0!
0*
09
0>
0C
#980830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#980840000000
0!
0*
09
0>
0C
#980850000000
1!
1*
b10 6
19
1>
1C
b10 G
#980860000000
0!
0*
09
0>
0C
#980870000000
1!
1*
b11 6
19
1>
1C
b11 G
#980880000000
0!
0*
09
0>
0C
#980890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#980900000000
0!
0*
09
0>
0C
#980910000000
1!
1*
b101 6
19
1>
1C
b101 G
#980920000000
0!
0*
09
0>
0C
#980930000000
1!
1*
b110 6
19
1>
1C
b110 G
#980940000000
0!
0*
09
0>
0C
#980950000000
1!
1*
b111 6
19
1>
1C
b111 G
#980960000000
0!
0*
09
0>
0C
#980970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#980980000000
0!
0*
09
0>
0C
#980990000000
1!
1*
b1 6
19
1>
1C
b1 G
#981000000000
0!
0*
09
0>
0C
#981010000000
1!
1*
b10 6
19
1>
1C
b10 G
#981020000000
0!
0*
09
0>
0C
#981030000000
1!
1*
b11 6
19
1>
1C
b11 G
#981040000000
0!
0*
09
0>
0C
#981050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#981060000000
0!
0*
09
0>
0C
#981070000000
1!
1*
b101 6
19
1>
1C
b101 G
#981080000000
0!
0*
09
0>
0C
#981090000000
1!
1*
b110 6
19
1>
1C
b110 G
#981100000000
0!
0*
09
0>
0C
#981110000000
1!
1*
b111 6
19
1>
1C
b111 G
#981120000000
0!
0*
09
0>
0C
#981130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#981140000000
0!
0*
09
0>
0C
#981150000000
1!
1*
b1 6
19
1>
1C
b1 G
#981160000000
0!
0*
09
0>
0C
#981170000000
1!
1*
b10 6
19
1>
1C
b10 G
#981180000000
0!
0*
09
0>
0C
#981190000000
1!
1*
b11 6
19
1>
1C
b11 G
#981200000000
0!
0*
09
0>
0C
#981210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#981220000000
0!
0*
09
0>
0C
#981230000000
1!
1*
b101 6
19
1>
1C
b101 G
#981240000000
0!
0*
09
0>
0C
#981250000000
1!
1*
b110 6
19
1>
1C
b110 G
#981260000000
0!
0*
09
0>
0C
#981270000000
1!
1*
b111 6
19
1>
1C
b111 G
#981280000000
0!
1"
0*
1+
09
1:
0>
0C
#981290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#981300000000
0!
0*
09
0>
0C
#981310000000
1!
1*
b1 6
19
1>
1C
b1 G
#981320000000
0!
0*
09
0>
0C
#981330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#981340000000
0!
0*
09
0>
0C
#981350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#981360000000
0!
0*
09
0>
0C
#981370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#981380000000
0!
0*
09
0>
0C
#981390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#981400000000
0!
0#
0*
0,
09
0>
0?
0C
#981410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#981420000000
0!
0*
09
0>
0C
#981430000000
1!
1*
19
1>
1C
#981440000000
0!
0*
09
0>
0C
#981450000000
1!
1*
19
1>
1C
#981460000000
0!
0*
09
0>
0C
#981470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#981480000000
0!
0*
09
0>
0C
#981490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#981500000000
0!
0*
09
0>
0C
#981510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#981520000000
0!
0*
09
0>
0C
#981530000000
1!
1*
b10 6
19
1>
1C
b10 G
#981540000000
0!
0*
09
0>
0C
#981550000000
1!
1*
b11 6
19
1>
1C
b11 G
#981560000000
0!
0*
09
0>
0C
#981570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#981580000000
0!
0*
09
0>
0C
#981590000000
1!
1*
b101 6
19
1>
1C
b101 G
#981600000000
0!
0*
09
0>
0C
#981610000000
1!
1*
b110 6
19
1>
1C
b110 G
#981620000000
0!
0*
09
0>
0C
#981630000000
1!
1*
b111 6
19
1>
1C
b111 G
#981640000000
0!
0*
09
0>
0C
#981650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#981660000000
0!
0*
09
0>
0C
#981670000000
1!
1*
b1 6
19
1>
1C
b1 G
#981680000000
0!
0*
09
0>
0C
#981690000000
1!
1*
b10 6
19
1>
1C
b10 G
#981700000000
0!
0*
09
0>
0C
#981710000000
1!
1*
b11 6
19
1>
1C
b11 G
#981720000000
0!
0*
09
0>
0C
#981730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#981740000000
0!
0*
09
0>
0C
#981750000000
1!
1*
b101 6
19
1>
1C
b101 G
#981760000000
0!
0*
09
0>
0C
#981770000000
1!
1*
b110 6
19
1>
1C
b110 G
#981780000000
0!
0*
09
0>
0C
#981790000000
1!
1*
b111 6
19
1>
1C
b111 G
#981800000000
0!
0*
09
0>
0C
#981810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#981820000000
0!
0*
09
0>
0C
#981830000000
1!
1*
b1 6
19
1>
1C
b1 G
#981840000000
0!
0*
09
0>
0C
#981850000000
1!
1*
b10 6
19
1>
1C
b10 G
#981860000000
0!
0*
09
0>
0C
#981870000000
1!
1*
b11 6
19
1>
1C
b11 G
#981880000000
0!
0*
09
0>
0C
#981890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#981900000000
0!
0*
09
0>
0C
#981910000000
1!
1*
b101 6
19
1>
1C
b101 G
#981920000000
0!
0*
09
0>
0C
#981930000000
1!
1*
b110 6
19
1>
1C
b110 G
#981940000000
0!
0*
09
0>
0C
#981950000000
1!
1*
b111 6
19
1>
1C
b111 G
#981960000000
0!
1"
0*
1+
09
1:
0>
0C
#981970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#981980000000
0!
0*
09
0>
0C
#981990000000
1!
1*
b1 6
19
1>
1C
b1 G
#982000000000
0!
0*
09
0>
0C
#982010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#982020000000
0!
0*
09
0>
0C
#982030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#982040000000
0!
0*
09
0>
0C
#982050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#982060000000
0!
0*
09
0>
0C
#982070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#982080000000
0!
0#
0*
0,
09
0>
0?
0C
#982090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#982100000000
0!
0*
09
0>
0C
#982110000000
1!
1*
19
1>
1C
#982120000000
0!
0*
09
0>
0C
#982130000000
1!
1*
19
1>
1C
#982140000000
0!
0*
09
0>
0C
#982150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#982160000000
0!
0*
09
0>
0C
#982170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#982180000000
0!
0*
09
0>
0C
#982190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#982200000000
0!
0*
09
0>
0C
#982210000000
1!
1*
b10 6
19
1>
1C
b10 G
#982220000000
0!
0*
09
0>
0C
#982230000000
1!
1*
b11 6
19
1>
1C
b11 G
#982240000000
0!
0*
09
0>
0C
#982250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#982260000000
0!
0*
09
0>
0C
#982270000000
1!
1*
b101 6
19
1>
1C
b101 G
#982280000000
0!
0*
09
0>
0C
#982290000000
1!
1*
b110 6
19
1>
1C
b110 G
#982300000000
0!
0*
09
0>
0C
#982310000000
1!
1*
b111 6
19
1>
1C
b111 G
#982320000000
0!
0*
09
0>
0C
#982330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#982340000000
0!
0*
09
0>
0C
#982350000000
1!
1*
b1 6
19
1>
1C
b1 G
#982360000000
0!
0*
09
0>
0C
#982370000000
1!
1*
b10 6
19
1>
1C
b10 G
#982380000000
0!
0*
09
0>
0C
#982390000000
1!
1*
b11 6
19
1>
1C
b11 G
#982400000000
0!
0*
09
0>
0C
#982410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#982420000000
0!
0*
09
0>
0C
#982430000000
1!
1*
b101 6
19
1>
1C
b101 G
#982440000000
0!
0*
09
0>
0C
#982450000000
1!
1*
b110 6
19
1>
1C
b110 G
#982460000000
0!
0*
09
0>
0C
#982470000000
1!
1*
b111 6
19
1>
1C
b111 G
#982480000000
0!
0*
09
0>
0C
#982490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#982500000000
0!
0*
09
0>
0C
#982510000000
1!
1*
b1 6
19
1>
1C
b1 G
#982520000000
0!
0*
09
0>
0C
#982530000000
1!
1*
b10 6
19
1>
1C
b10 G
#982540000000
0!
0*
09
0>
0C
#982550000000
1!
1*
b11 6
19
1>
1C
b11 G
#982560000000
0!
0*
09
0>
0C
#982570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#982580000000
0!
0*
09
0>
0C
#982590000000
1!
1*
b101 6
19
1>
1C
b101 G
#982600000000
0!
0*
09
0>
0C
#982610000000
1!
1*
b110 6
19
1>
1C
b110 G
#982620000000
0!
0*
09
0>
0C
#982630000000
1!
1*
b111 6
19
1>
1C
b111 G
#982640000000
0!
1"
0*
1+
09
1:
0>
0C
#982650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#982660000000
0!
0*
09
0>
0C
#982670000000
1!
1*
b1 6
19
1>
1C
b1 G
#982680000000
0!
0*
09
0>
0C
#982690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#982700000000
0!
0*
09
0>
0C
#982710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#982720000000
0!
0*
09
0>
0C
#982730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#982740000000
0!
0*
09
0>
0C
#982750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#982760000000
0!
0#
0*
0,
09
0>
0?
0C
#982770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#982780000000
0!
0*
09
0>
0C
#982790000000
1!
1*
19
1>
1C
#982800000000
0!
0*
09
0>
0C
#982810000000
1!
1*
19
1>
1C
#982820000000
0!
0*
09
0>
0C
#982830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#982840000000
0!
0*
09
0>
0C
#982850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#982860000000
0!
0*
09
0>
0C
#982870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#982880000000
0!
0*
09
0>
0C
#982890000000
1!
1*
b10 6
19
1>
1C
b10 G
#982900000000
0!
0*
09
0>
0C
#982910000000
1!
1*
b11 6
19
1>
1C
b11 G
#982920000000
0!
0*
09
0>
0C
#982930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#982940000000
0!
0*
09
0>
0C
#982950000000
1!
1*
b101 6
19
1>
1C
b101 G
#982960000000
0!
0*
09
0>
0C
#982970000000
1!
1*
b110 6
19
1>
1C
b110 G
#982980000000
0!
0*
09
0>
0C
#982990000000
1!
1*
b111 6
19
1>
1C
b111 G
#983000000000
0!
0*
09
0>
0C
#983010000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#983020000000
0!
0*
09
0>
0C
#983030000000
1!
1*
b1 6
19
1>
1C
b1 G
#983040000000
0!
0*
09
0>
0C
#983050000000
1!
1*
b10 6
19
1>
1C
b10 G
#983060000000
0!
0*
09
0>
0C
#983070000000
1!
1*
b11 6
19
1>
1C
b11 G
#983080000000
0!
0*
09
0>
0C
#983090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#983100000000
0!
0*
09
0>
0C
#983110000000
1!
1*
b101 6
19
1>
1C
b101 G
#983120000000
0!
0*
09
0>
0C
#983130000000
1!
1*
b110 6
19
1>
1C
b110 G
#983140000000
0!
0*
09
0>
0C
#983150000000
1!
1*
b111 6
19
1>
1C
b111 G
#983160000000
0!
0*
09
0>
0C
#983170000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#983180000000
0!
0*
09
0>
0C
#983190000000
1!
1*
b1 6
19
1>
1C
b1 G
#983200000000
0!
0*
09
0>
0C
#983210000000
1!
1*
b10 6
19
1>
1C
b10 G
#983220000000
0!
0*
09
0>
0C
#983230000000
1!
1*
b11 6
19
1>
1C
b11 G
#983240000000
0!
0*
09
0>
0C
#983250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#983260000000
0!
0*
09
0>
0C
#983270000000
1!
1*
b101 6
19
1>
1C
b101 G
#983280000000
0!
0*
09
0>
0C
#983290000000
1!
1*
b110 6
19
1>
1C
b110 G
#983300000000
0!
0*
09
0>
0C
#983310000000
1!
1*
b111 6
19
1>
1C
b111 G
#983320000000
0!
1"
0*
1+
09
1:
0>
0C
#983330000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#983340000000
0!
0*
09
0>
0C
#983350000000
1!
1*
b1 6
19
1>
1C
b1 G
#983360000000
0!
0*
09
0>
0C
#983370000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#983380000000
0!
0*
09
0>
0C
#983390000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#983400000000
0!
0*
09
0>
0C
#983410000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#983420000000
0!
0*
09
0>
0C
#983430000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#983440000000
0!
0#
0*
0,
09
0>
0?
0C
#983450000000
1!
1*
02
19
1>
0@
0A
0B
1C
#983460000000
0!
0*
09
0>
0C
#983470000000
1!
1*
19
1>
1C
#983480000000
0!
0*
09
0>
0C
#983490000000
1!
1*
19
1>
1C
#983500000000
0!
0*
09
0>
0C
#983510000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#983520000000
0!
0*
09
0>
0C
#983530000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#983540000000
0!
0*
09
0>
0C
#983550000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#983560000000
0!
0*
09
0>
0C
#983570000000
1!
1*
b10 6
19
1>
1C
b10 G
#983580000000
0!
0*
09
0>
0C
#983590000000
1!
1*
b11 6
19
1>
1C
b11 G
#983600000000
0!
0*
09
0>
0C
#983610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#983620000000
0!
0*
09
0>
0C
#983630000000
1!
1*
b101 6
19
1>
1C
b101 G
#983640000000
0!
0*
09
0>
0C
#983650000000
1!
1*
b110 6
19
1>
1C
b110 G
#983660000000
0!
0*
09
0>
0C
#983670000000
1!
1*
b111 6
19
1>
1C
b111 G
#983680000000
0!
0*
09
0>
0C
#983690000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#983700000000
0!
0*
09
0>
0C
#983710000000
1!
1*
b1 6
19
1>
1C
b1 G
#983720000000
0!
0*
09
0>
0C
#983730000000
1!
1*
b10 6
19
1>
1C
b10 G
#983740000000
0!
0*
09
0>
0C
#983750000000
1!
1*
b11 6
19
1>
1C
b11 G
#983760000000
0!
0*
09
0>
0C
#983770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#983780000000
0!
0*
09
0>
0C
#983790000000
1!
1*
b101 6
19
1>
1C
b101 G
#983800000000
0!
0*
09
0>
0C
#983810000000
1!
1*
b110 6
19
1>
1C
b110 G
#983820000000
0!
0*
09
0>
0C
#983830000000
1!
1*
b111 6
19
1>
1C
b111 G
#983840000000
0!
0*
09
0>
0C
#983850000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#983860000000
0!
0*
09
0>
0C
#983870000000
1!
1*
b1 6
19
1>
1C
b1 G
#983880000000
0!
0*
09
0>
0C
#983890000000
1!
1*
b10 6
19
1>
1C
b10 G
#983900000000
0!
0*
09
0>
0C
#983910000000
1!
1*
b11 6
19
1>
1C
b11 G
#983920000000
0!
0*
09
0>
0C
#983930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#983940000000
0!
0*
09
0>
0C
#983950000000
1!
1*
b101 6
19
1>
1C
b101 G
#983960000000
0!
0*
09
0>
0C
#983970000000
1!
1*
b110 6
19
1>
1C
b110 G
#983980000000
0!
0*
09
0>
0C
#983990000000
1!
1*
b111 6
19
1>
1C
b111 G
#984000000000
0!
1"
0*
1+
09
1:
0>
0C
#984010000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#984020000000
0!
0*
09
0>
0C
#984030000000
1!
1*
b1 6
19
1>
1C
b1 G
#984040000000
0!
0*
09
0>
0C
#984050000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#984060000000
0!
0*
09
0>
0C
#984070000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#984080000000
0!
0*
09
0>
0C
#984090000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#984100000000
0!
0*
09
0>
0C
#984110000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#984120000000
0!
0#
0*
0,
09
0>
0?
0C
#984130000000
1!
1*
02
19
1>
0@
0A
0B
1C
#984140000000
0!
0*
09
0>
0C
#984150000000
1!
1*
19
1>
1C
#984160000000
0!
0*
09
0>
0C
#984170000000
1!
1*
19
1>
1C
#984180000000
0!
0*
09
0>
0C
#984190000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#984200000000
0!
0*
09
0>
0C
#984210000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#984220000000
0!
0*
09
0>
0C
#984230000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#984240000000
0!
0*
09
0>
0C
#984250000000
1!
1*
b10 6
19
1>
1C
b10 G
#984260000000
0!
0*
09
0>
0C
#984270000000
1!
1*
b11 6
19
1>
1C
b11 G
#984280000000
0!
0*
09
0>
0C
#984290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#984300000000
0!
0*
09
0>
0C
#984310000000
1!
1*
b101 6
19
1>
1C
b101 G
#984320000000
0!
0*
09
0>
0C
#984330000000
1!
1*
b110 6
19
1>
1C
b110 G
#984340000000
0!
0*
09
0>
0C
#984350000000
1!
1*
b111 6
19
1>
1C
b111 G
#984360000000
0!
0*
09
0>
0C
#984370000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#984380000000
0!
0*
09
0>
0C
#984390000000
1!
1*
b1 6
19
1>
1C
b1 G
#984400000000
0!
0*
09
0>
0C
#984410000000
1!
1*
b10 6
19
1>
1C
b10 G
#984420000000
0!
0*
09
0>
0C
#984430000000
1!
1*
b11 6
19
1>
1C
b11 G
#984440000000
0!
0*
09
0>
0C
#984450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#984460000000
0!
0*
09
0>
0C
#984470000000
1!
1*
b101 6
19
1>
1C
b101 G
#984480000000
0!
0*
09
0>
0C
#984490000000
1!
1*
b110 6
19
1>
1C
b110 G
#984500000000
0!
0*
09
0>
0C
#984510000000
1!
1*
b111 6
19
1>
1C
b111 G
#984520000000
0!
0*
09
0>
0C
#984530000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#984540000000
0!
0*
09
0>
0C
#984550000000
1!
1*
b1 6
19
1>
1C
b1 G
#984560000000
0!
0*
09
0>
0C
#984570000000
1!
1*
b10 6
19
1>
1C
b10 G
#984580000000
0!
0*
09
0>
0C
#984590000000
1!
1*
b11 6
19
1>
1C
b11 G
#984600000000
0!
0*
09
0>
0C
#984610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#984620000000
0!
0*
09
0>
0C
#984630000000
1!
1*
b101 6
19
1>
1C
b101 G
#984640000000
0!
0*
09
0>
0C
#984650000000
1!
1*
b110 6
19
1>
1C
b110 G
#984660000000
0!
0*
09
0>
0C
#984670000000
1!
1*
b111 6
19
1>
1C
b111 G
#984680000000
0!
1"
0*
1+
09
1:
0>
0C
#984690000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#984700000000
0!
0*
09
0>
0C
#984710000000
1!
1*
b1 6
19
1>
1C
b1 G
#984720000000
0!
0*
09
0>
0C
#984730000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#984740000000
0!
0*
09
0>
0C
#984750000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#984760000000
0!
0*
09
0>
0C
#984770000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#984780000000
0!
0*
09
0>
0C
#984790000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#984800000000
0!
0#
0*
0,
09
0>
0?
0C
#984810000000
1!
1*
02
19
1>
0@
0A
0B
1C
#984820000000
0!
0*
09
0>
0C
#984830000000
1!
1*
19
1>
1C
#984840000000
0!
0*
09
0>
0C
#984850000000
1!
1*
19
1>
1C
#984860000000
0!
0*
09
0>
0C
#984870000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#984880000000
0!
0*
09
0>
0C
#984890000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#984900000000
0!
0*
09
0>
0C
#984910000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#984920000000
0!
0*
09
0>
0C
#984930000000
1!
1*
b10 6
19
1>
1C
b10 G
#984940000000
0!
0*
09
0>
0C
#984950000000
1!
1*
b11 6
19
1>
1C
b11 G
#984960000000
0!
0*
09
0>
0C
#984970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#984980000000
0!
0*
09
0>
0C
#984990000000
1!
1*
b101 6
19
1>
1C
b101 G
#985000000000
0!
0*
09
0>
0C
#985010000000
1!
1*
b110 6
19
1>
1C
b110 G
#985020000000
0!
0*
09
0>
0C
#985030000000
1!
1*
b111 6
19
1>
1C
b111 G
#985040000000
0!
0*
09
0>
0C
#985050000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#985060000000
0!
0*
09
0>
0C
#985070000000
1!
1*
b1 6
19
1>
1C
b1 G
#985080000000
0!
0*
09
0>
0C
#985090000000
1!
1*
b10 6
19
1>
1C
b10 G
#985100000000
0!
0*
09
0>
0C
#985110000000
1!
1*
b11 6
19
1>
1C
b11 G
#985120000000
0!
0*
09
0>
0C
#985130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#985140000000
0!
0*
09
0>
0C
#985150000000
1!
1*
b101 6
19
1>
1C
b101 G
#985160000000
0!
0*
09
0>
0C
#985170000000
1!
1*
b110 6
19
1>
1C
b110 G
#985180000000
0!
0*
09
0>
0C
#985190000000
1!
1*
b111 6
19
1>
1C
b111 G
#985200000000
0!
0*
09
0>
0C
#985210000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#985220000000
0!
0*
09
0>
0C
#985230000000
1!
1*
b1 6
19
1>
1C
b1 G
#985240000000
0!
0*
09
0>
0C
#985250000000
1!
1*
b10 6
19
1>
1C
b10 G
#985260000000
0!
0*
09
0>
0C
#985270000000
1!
1*
b11 6
19
1>
1C
b11 G
#985280000000
0!
0*
09
0>
0C
#985290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#985300000000
0!
0*
09
0>
0C
#985310000000
1!
1*
b101 6
19
1>
1C
b101 G
#985320000000
0!
0*
09
0>
0C
#985330000000
1!
1*
b110 6
19
1>
1C
b110 G
#985340000000
0!
0*
09
0>
0C
#985350000000
1!
1*
b111 6
19
1>
1C
b111 G
#985360000000
0!
1"
0*
1+
09
1:
0>
0C
#985370000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#985380000000
0!
0*
09
0>
0C
#985390000000
1!
1*
b1 6
19
1>
1C
b1 G
#985400000000
0!
0*
09
0>
0C
#985410000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#985420000000
0!
0*
09
0>
0C
#985430000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#985440000000
0!
0*
09
0>
0C
#985450000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#985460000000
0!
0*
09
0>
0C
#985470000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#985480000000
0!
0#
0*
0,
09
0>
0?
0C
#985490000000
1!
1*
02
19
1>
0@
0A
0B
1C
#985500000000
0!
0*
09
0>
0C
#985510000000
1!
1*
19
1>
1C
#985520000000
0!
0*
09
0>
0C
#985530000000
1!
1*
19
1>
1C
#985540000000
0!
0*
09
0>
0C
#985550000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#985560000000
0!
0*
09
0>
0C
#985570000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#985580000000
0!
0*
09
0>
0C
#985590000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#985600000000
0!
0*
09
0>
0C
#985610000000
1!
1*
b10 6
19
1>
1C
b10 G
#985620000000
0!
0*
09
0>
0C
#985630000000
1!
1*
b11 6
19
1>
1C
b11 G
#985640000000
0!
0*
09
0>
0C
#985650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#985660000000
0!
0*
09
0>
0C
#985670000000
1!
1*
b101 6
19
1>
1C
b101 G
#985680000000
0!
0*
09
0>
0C
#985690000000
1!
1*
b110 6
19
1>
1C
b110 G
#985700000000
0!
0*
09
0>
0C
#985710000000
1!
1*
b111 6
19
1>
1C
b111 G
#985720000000
0!
0*
09
0>
0C
#985730000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#985740000000
0!
0*
09
0>
0C
#985750000000
1!
1*
b1 6
19
1>
1C
b1 G
#985760000000
0!
0*
09
0>
0C
#985770000000
1!
1*
b10 6
19
1>
1C
b10 G
#985780000000
0!
0*
09
0>
0C
#985790000000
1!
1*
b11 6
19
1>
1C
b11 G
#985800000000
0!
0*
09
0>
0C
#985810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#985820000000
0!
0*
09
0>
0C
#985830000000
1!
1*
b101 6
19
1>
1C
b101 G
#985840000000
0!
0*
09
0>
0C
#985850000000
1!
1*
b110 6
19
1>
1C
b110 G
#985860000000
0!
0*
09
0>
0C
#985870000000
1!
1*
b111 6
19
1>
1C
b111 G
#985880000000
0!
0*
09
0>
0C
#985890000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#985900000000
0!
0*
09
0>
0C
#985910000000
1!
1*
b1 6
19
1>
1C
b1 G
#985920000000
0!
0*
09
0>
0C
#985930000000
1!
1*
b10 6
19
1>
1C
b10 G
#985940000000
0!
0*
09
0>
0C
#985950000000
1!
1*
b11 6
19
1>
1C
b11 G
#985960000000
0!
0*
09
0>
0C
#985970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#985980000000
0!
0*
09
0>
0C
#985990000000
1!
1*
b101 6
19
1>
1C
b101 G
#986000000000
0!
0*
09
0>
0C
#986010000000
1!
1*
b110 6
19
1>
1C
b110 G
#986020000000
0!
0*
09
0>
0C
#986030000000
1!
1*
b111 6
19
1>
1C
b111 G
#986040000000
0!
1"
0*
1+
09
1:
0>
0C
#986050000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#986060000000
0!
0*
09
0>
0C
#986070000000
1!
1*
b1 6
19
1>
1C
b1 G
#986080000000
0!
0*
09
0>
0C
#986090000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#986100000000
0!
0*
09
0>
0C
#986110000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#986120000000
0!
0*
09
0>
0C
#986130000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#986140000000
0!
0*
09
0>
0C
#986150000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#986160000000
0!
0#
0*
0,
09
0>
0?
0C
#986170000000
1!
1*
02
19
1>
0@
0A
0B
1C
#986180000000
0!
0*
09
0>
0C
#986190000000
1!
1*
19
1>
1C
#986200000000
0!
0*
09
0>
0C
#986210000000
1!
1*
19
1>
1C
#986220000000
0!
0*
09
0>
0C
#986230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#986240000000
0!
0*
09
0>
0C
#986250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#986260000000
0!
0*
09
0>
0C
#986270000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#986280000000
0!
0*
09
0>
0C
#986290000000
1!
1*
b10 6
19
1>
1C
b10 G
#986300000000
0!
0*
09
0>
0C
#986310000000
1!
1*
b11 6
19
1>
1C
b11 G
#986320000000
0!
0*
09
0>
0C
#986330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#986340000000
0!
0*
09
0>
0C
#986350000000
1!
1*
b101 6
19
1>
1C
b101 G
#986360000000
0!
0*
09
0>
0C
#986370000000
1!
1*
b110 6
19
1>
1C
b110 G
#986380000000
0!
0*
09
0>
0C
#986390000000
1!
1*
b111 6
19
1>
1C
b111 G
#986400000000
0!
0*
09
0>
0C
#986410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#986420000000
0!
0*
09
0>
0C
#986430000000
1!
1*
b1 6
19
1>
1C
b1 G
#986440000000
0!
0*
09
0>
0C
#986450000000
1!
1*
b10 6
19
1>
1C
b10 G
#986460000000
0!
0*
09
0>
0C
#986470000000
1!
1*
b11 6
19
1>
1C
b11 G
#986480000000
0!
0*
09
0>
0C
#986490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#986500000000
0!
0*
09
0>
0C
#986510000000
1!
1*
b101 6
19
1>
1C
b101 G
#986520000000
0!
0*
09
0>
0C
#986530000000
1!
1*
b110 6
19
1>
1C
b110 G
#986540000000
0!
0*
09
0>
0C
#986550000000
1!
1*
b111 6
19
1>
1C
b111 G
#986560000000
0!
0*
09
0>
0C
#986570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#986580000000
0!
0*
09
0>
0C
#986590000000
1!
1*
b1 6
19
1>
1C
b1 G
#986600000000
0!
0*
09
0>
0C
#986610000000
1!
1*
b10 6
19
1>
1C
b10 G
#986620000000
0!
0*
09
0>
0C
#986630000000
1!
1*
b11 6
19
1>
1C
b11 G
#986640000000
0!
0*
09
0>
0C
#986650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#986660000000
0!
0*
09
0>
0C
#986670000000
1!
1*
b101 6
19
1>
1C
b101 G
#986680000000
0!
0*
09
0>
0C
#986690000000
1!
1*
b110 6
19
1>
1C
b110 G
#986700000000
0!
0*
09
0>
0C
#986710000000
1!
1*
b111 6
19
1>
1C
b111 G
#986720000000
0!
1"
0*
1+
09
1:
0>
0C
#986730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#986740000000
0!
0*
09
0>
0C
#986750000000
1!
1*
b1 6
19
1>
1C
b1 G
#986760000000
0!
0*
09
0>
0C
#986770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#986780000000
0!
0*
09
0>
0C
#986790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#986800000000
0!
0*
09
0>
0C
#986810000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#986820000000
0!
0*
09
0>
0C
#986830000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#986840000000
0!
0#
0*
0,
09
0>
0?
0C
#986850000000
1!
1*
02
19
1>
0@
0A
0B
1C
#986860000000
0!
0*
09
0>
0C
#986870000000
1!
1*
19
1>
1C
#986880000000
0!
0*
09
0>
0C
#986890000000
1!
1*
19
1>
1C
#986900000000
0!
0*
09
0>
0C
#986910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#986920000000
0!
0*
09
0>
0C
#986930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#986940000000
0!
0*
09
0>
0C
#986950000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#986960000000
0!
0*
09
0>
0C
#986970000000
1!
1*
b10 6
19
1>
1C
b10 G
#986980000000
0!
0*
09
0>
0C
#986990000000
1!
1*
b11 6
19
1>
1C
b11 G
#987000000000
0!
0*
09
0>
0C
#987010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#987020000000
0!
0*
09
0>
0C
#987030000000
1!
1*
b101 6
19
1>
1C
b101 G
#987040000000
0!
0*
09
0>
0C
#987050000000
1!
1*
b110 6
19
1>
1C
b110 G
#987060000000
0!
0*
09
0>
0C
#987070000000
1!
1*
b111 6
19
1>
1C
b111 G
#987080000000
0!
0*
09
0>
0C
#987090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#987100000000
0!
0*
09
0>
0C
#987110000000
1!
1*
b1 6
19
1>
1C
b1 G
#987120000000
0!
0*
09
0>
0C
#987130000000
1!
1*
b10 6
19
1>
1C
b10 G
#987140000000
0!
0*
09
0>
0C
#987150000000
1!
1*
b11 6
19
1>
1C
b11 G
#987160000000
0!
0*
09
0>
0C
#987170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#987180000000
0!
0*
09
0>
0C
#987190000000
1!
1*
b101 6
19
1>
1C
b101 G
#987200000000
0!
0*
09
0>
0C
#987210000000
1!
1*
b110 6
19
1>
1C
b110 G
#987220000000
0!
0*
09
0>
0C
#987230000000
1!
1*
b111 6
19
1>
1C
b111 G
#987240000000
0!
0*
09
0>
0C
#987250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#987260000000
0!
0*
09
0>
0C
#987270000000
1!
1*
b1 6
19
1>
1C
b1 G
#987280000000
0!
0*
09
0>
0C
#987290000000
1!
1*
b10 6
19
1>
1C
b10 G
#987300000000
0!
0*
09
0>
0C
#987310000000
1!
1*
b11 6
19
1>
1C
b11 G
#987320000000
0!
0*
09
0>
0C
#987330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#987340000000
0!
0*
09
0>
0C
#987350000000
1!
1*
b101 6
19
1>
1C
b101 G
#987360000000
0!
0*
09
0>
0C
#987370000000
1!
1*
b110 6
19
1>
1C
b110 G
#987380000000
0!
0*
09
0>
0C
#987390000000
1!
1*
b111 6
19
1>
1C
b111 G
#987400000000
0!
1"
0*
1+
09
1:
0>
0C
#987410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#987420000000
0!
0*
09
0>
0C
#987430000000
1!
1*
b1 6
19
1>
1C
b1 G
#987440000000
0!
0*
09
0>
0C
#987450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#987460000000
0!
0*
09
0>
0C
#987470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#987480000000
0!
0*
09
0>
0C
#987490000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#987500000000
0!
0*
09
0>
0C
#987510000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#987520000000
0!
0#
0*
0,
09
0>
0?
0C
#987530000000
1!
1*
02
19
1>
0@
0A
0B
1C
#987540000000
0!
0*
09
0>
0C
#987550000000
1!
1*
19
1>
1C
#987560000000
0!
0*
09
0>
0C
#987570000000
1!
1*
19
1>
1C
#987580000000
0!
0*
09
0>
0C
#987590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#987600000000
0!
0*
09
0>
0C
#987610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#987620000000
0!
0*
09
0>
0C
#987630000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#987640000000
0!
0*
09
0>
0C
#987650000000
1!
1*
b10 6
19
1>
1C
b10 G
#987660000000
0!
0*
09
0>
0C
#987670000000
1!
1*
b11 6
19
1>
1C
b11 G
#987680000000
0!
0*
09
0>
0C
#987690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#987700000000
0!
0*
09
0>
0C
#987710000000
1!
1*
b101 6
19
1>
1C
b101 G
#987720000000
0!
0*
09
0>
0C
#987730000000
1!
1*
b110 6
19
1>
1C
b110 G
#987740000000
0!
0*
09
0>
0C
#987750000000
1!
1*
b111 6
19
1>
1C
b111 G
#987760000000
0!
0*
09
0>
0C
#987770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#987780000000
0!
0*
09
0>
0C
#987790000000
1!
1*
b1 6
19
1>
1C
b1 G
#987800000000
0!
0*
09
0>
0C
#987810000000
1!
1*
b10 6
19
1>
1C
b10 G
#987820000000
0!
0*
09
0>
0C
#987830000000
1!
1*
b11 6
19
1>
1C
b11 G
#987840000000
0!
0*
09
0>
0C
#987850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#987860000000
0!
0*
09
0>
0C
#987870000000
1!
1*
b101 6
19
1>
1C
b101 G
#987880000000
0!
0*
09
0>
0C
#987890000000
1!
1*
b110 6
19
1>
1C
b110 G
#987900000000
0!
0*
09
0>
0C
#987910000000
1!
1*
b111 6
19
1>
1C
b111 G
#987920000000
0!
0*
09
0>
0C
#987930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#987940000000
0!
0*
09
0>
0C
#987950000000
1!
1*
b1 6
19
1>
1C
b1 G
#987960000000
0!
0*
09
0>
0C
#987970000000
1!
1*
b10 6
19
1>
1C
b10 G
#987980000000
0!
0*
09
0>
0C
#987990000000
1!
1*
b11 6
19
1>
1C
b11 G
#988000000000
0!
0*
09
0>
0C
#988010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#988020000000
0!
0*
09
0>
0C
#988030000000
1!
1*
b101 6
19
1>
1C
b101 G
#988040000000
0!
0*
09
0>
0C
#988050000000
1!
1*
b110 6
19
1>
1C
b110 G
#988060000000
0!
0*
09
0>
0C
#988070000000
1!
1*
b111 6
19
1>
1C
b111 G
#988080000000
0!
1"
0*
1+
09
1:
0>
0C
#988090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#988100000000
0!
0*
09
0>
0C
#988110000000
1!
1*
b1 6
19
1>
1C
b1 G
#988120000000
0!
0*
09
0>
0C
#988130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#988140000000
0!
0*
09
0>
0C
#988150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#988160000000
0!
0*
09
0>
0C
#988170000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#988180000000
0!
0*
09
0>
0C
#988190000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#988200000000
0!
0#
0*
0,
09
0>
0?
0C
#988210000000
1!
1*
02
19
1>
0@
0A
0B
1C
#988220000000
0!
0*
09
0>
0C
#988230000000
1!
1*
19
1>
1C
#988240000000
0!
0*
09
0>
0C
#988250000000
1!
1*
19
1>
1C
#988260000000
0!
0*
09
0>
0C
#988270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#988280000000
0!
0*
09
0>
0C
#988290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#988300000000
0!
0*
09
0>
0C
#988310000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#988320000000
0!
0*
09
0>
0C
#988330000000
1!
1*
b10 6
19
1>
1C
b10 G
#988340000000
0!
0*
09
0>
0C
#988350000000
1!
1*
b11 6
19
1>
1C
b11 G
#988360000000
0!
0*
09
0>
0C
#988370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#988380000000
0!
0*
09
0>
0C
#988390000000
1!
1*
b101 6
19
1>
1C
b101 G
#988400000000
0!
0*
09
0>
0C
#988410000000
1!
1*
b110 6
19
1>
1C
b110 G
#988420000000
0!
0*
09
0>
0C
#988430000000
1!
1*
b111 6
19
1>
1C
b111 G
#988440000000
0!
0*
09
0>
0C
#988450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#988460000000
0!
0*
09
0>
0C
#988470000000
1!
1*
b1 6
19
1>
1C
b1 G
#988480000000
0!
0*
09
0>
0C
#988490000000
1!
1*
b10 6
19
1>
1C
b10 G
#988500000000
0!
0*
09
0>
0C
#988510000000
1!
1*
b11 6
19
1>
1C
b11 G
#988520000000
0!
0*
09
0>
0C
#988530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#988540000000
0!
0*
09
0>
0C
#988550000000
1!
1*
b101 6
19
1>
1C
b101 G
#988560000000
0!
0*
09
0>
0C
#988570000000
1!
1*
b110 6
19
1>
1C
b110 G
#988580000000
0!
0*
09
0>
0C
#988590000000
1!
1*
b111 6
19
1>
1C
b111 G
#988600000000
0!
0*
09
0>
0C
#988610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#988620000000
0!
0*
09
0>
0C
#988630000000
1!
1*
b1 6
19
1>
1C
b1 G
#988640000000
0!
0*
09
0>
0C
#988650000000
1!
1*
b10 6
19
1>
1C
b10 G
#988660000000
0!
0*
09
0>
0C
#988670000000
1!
1*
b11 6
19
1>
1C
b11 G
#988680000000
0!
0*
09
0>
0C
#988690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#988700000000
0!
0*
09
0>
0C
#988710000000
1!
1*
b101 6
19
1>
1C
b101 G
#988720000000
0!
0*
09
0>
0C
#988730000000
1!
1*
b110 6
19
1>
1C
b110 G
#988740000000
0!
0*
09
0>
0C
#988750000000
1!
1*
b111 6
19
1>
1C
b111 G
#988760000000
0!
1"
0*
1+
09
1:
0>
0C
#988770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#988780000000
0!
0*
09
0>
0C
#988790000000
1!
1*
b1 6
19
1>
1C
b1 G
#988800000000
0!
0*
09
0>
0C
#988810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#988820000000
0!
0*
09
0>
0C
#988830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#988840000000
0!
0*
09
0>
0C
#988850000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#988860000000
0!
0*
09
0>
0C
#988870000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#988880000000
0!
0#
0*
0,
09
0>
0?
0C
#988890000000
1!
1*
02
19
1>
0@
0A
0B
1C
#988900000000
0!
0*
09
0>
0C
#988910000000
1!
1*
19
1>
1C
#988920000000
0!
0*
09
0>
0C
#988930000000
1!
1*
19
1>
1C
#988940000000
0!
0*
09
0>
0C
#988950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#988960000000
0!
0*
09
0>
0C
#988970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#988980000000
0!
0*
09
0>
0C
#988990000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#989000000000
0!
0*
09
0>
0C
#989010000000
1!
1*
b10 6
19
1>
1C
b10 G
#989020000000
0!
0*
09
0>
0C
#989030000000
1!
1*
b11 6
19
1>
1C
b11 G
#989040000000
0!
0*
09
0>
0C
#989050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#989060000000
0!
0*
09
0>
0C
#989070000000
1!
1*
b101 6
19
1>
1C
b101 G
#989080000000
0!
0*
09
0>
0C
#989090000000
1!
1*
b110 6
19
1>
1C
b110 G
#989100000000
0!
0*
09
0>
0C
#989110000000
1!
1*
b111 6
19
1>
1C
b111 G
#989120000000
0!
0*
09
0>
0C
#989130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#989140000000
0!
0*
09
0>
0C
#989150000000
1!
1*
b1 6
19
1>
1C
b1 G
#989160000000
0!
0*
09
0>
0C
#989170000000
1!
1*
b10 6
19
1>
1C
b10 G
#989180000000
0!
0*
09
0>
0C
#989190000000
1!
1*
b11 6
19
1>
1C
b11 G
#989200000000
0!
0*
09
0>
0C
#989210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#989220000000
0!
0*
09
0>
0C
#989230000000
1!
1*
b101 6
19
1>
1C
b101 G
#989240000000
0!
0*
09
0>
0C
#989250000000
1!
1*
b110 6
19
1>
1C
b110 G
#989260000000
0!
0*
09
0>
0C
#989270000000
1!
1*
b111 6
19
1>
1C
b111 G
#989280000000
0!
0*
09
0>
0C
#989290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#989300000000
0!
0*
09
0>
0C
#989310000000
1!
1*
b1 6
19
1>
1C
b1 G
#989320000000
0!
0*
09
0>
0C
#989330000000
1!
1*
b10 6
19
1>
1C
b10 G
#989340000000
0!
0*
09
0>
0C
#989350000000
1!
1*
b11 6
19
1>
1C
b11 G
#989360000000
0!
0*
09
0>
0C
#989370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#989380000000
0!
0*
09
0>
0C
#989390000000
1!
1*
b101 6
19
1>
1C
b101 G
#989400000000
0!
0*
09
0>
0C
#989410000000
1!
1*
b110 6
19
1>
1C
b110 G
#989420000000
0!
0*
09
0>
0C
#989430000000
1!
1*
b111 6
19
1>
1C
b111 G
#989440000000
0!
1"
0*
1+
09
1:
0>
0C
#989450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#989460000000
0!
0*
09
0>
0C
#989470000000
1!
1*
b1 6
19
1>
1C
b1 G
#989480000000
0!
0*
09
0>
0C
#989490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#989500000000
0!
0*
09
0>
0C
#989510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#989520000000
0!
0*
09
0>
0C
#989530000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#989540000000
0!
0*
09
0>
0C
#989550000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#989560000000
0!
0#
0*
0,
09
0>
0?
0C
#989570000000
1!
1*
02
19
1>
0@
0A
0B
1C
#989580000000
0!
0*
09
0>
0C
#989590000000
1!
1*
19
1>
1C
#989600000000
0!
0*
09
0>
0C
#989610000000
1!
1*
19
1>
1C
#989620000000
0!
0*
09
0>
0C
#989630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#989640000000
0!
0*
09
0>
0C
#989650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#989660000000
0!
0*
09
0>
0C
#989670000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#989680000000
0!
0*
09
0>
0C
#989690000000
1!
1*
b10 6
19
1>
1C
b10 G
#989700000000
0!
0*
09
0>
0C
#989710000000
1!
1*
b11 6
19
1>
1C
b11 G
#989720000000
0!
0*
09
0>
0C
#989730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#989740000000
0!
0*
09
0>
0C
#989750000000
1!
1*
b101 6
19
1>
1C
b101 G
#989760000000
0!
0*
09
0>
0C
#989770000000
1!
1*
b110 6
19
1>
1C
b110 G
#989780000000
0!
0*
09
0>
0C
#989790000000
1!
1*
b111 6
19
1>
1C
b111 G
#989800000000
0!
0*
09
0>
0C
#989810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#989820000000
0!
0*
09
0>
0C
#989830000000
1!
1*
b1 6
19
1>
1C
b1 G
#989840000000
0!
0*
09
0>
0C
#989850000000
1!
1*
b10 6
19
1>
1C
b10 G
#989860000000
0!
0*
09
0>
0C
#989870000000
1!
1*
b11 6
19
1>
1C
b11 G
#989880000000
0!
0*
09
0>
0C
#989890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#989900000000
0!
0*
09
0>
0C
#989910000000
1!
1*
b101 6
19
1>
1C
b101 G
#989920000000
0!
0*
09
0>
0C
#989930000000
1!
1*
b110 6
19
1>
1C
b110 G
#989940000000
0!
0*
09
0>
0C
#989950000000
1!
1*
b111 6
19
1>
1C
b111 G
#989960000000
0!
0*
09
0>
0C
#989970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#989980000000
0!
0*
09
0>
0C
#989990000000
1!
1*
b1 6
19
1>
1C
b1 G
#990000000000
0!
0*
09
0>
0C
#990010000000
1!
1*
b10 6
19
1>
1C
b10 G
#990020000000
0!
0*
09
0>
0C
#990030000000
1!
1*
b11 6
19
1>
1C
b11 G
#990040000000
0!
0*
09
0>
0C
#990050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#990060000000
0!
0*
09
0>
0C
#990070000000
1!
1*
b101 6
19
1>
1C
b101 G
#990080000000
0!
0*
09
0>
0C
#990090000000
1!
1*
b110 6
19
1>
1C
b110 G
#990100000000
0!
0*
09
0>
0C
#990110000000
1!
1*
b111 6
19
1>
1C
b111 G
#990120000000
0!
1"
0*
1+
09
1:
0>
0C
#990130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#990140000000
0!
0*
09
0>
0C
#990150000000
1!
1*
b1 6
19
1>
1C
b1 G
#990160000000
0!
0*
09
0>
0C
#990170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#990180000000
0!
0*
09
0>
0C
#990190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#990200000000
0!
0*
09
0>
0C
#990210000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#990220000000
0!
0*
09
0>
0C
#990230000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#990240000000
0!
0#
0*
0,
09
0>
0?
0C
#990250000000
1!
1*
02
19
1>
0@
0A
0B
1C
#990260000000
0!
0*
09
0>
0C
#990270000000
1!
1*
19
1>
1C
#990280000000
0!
0*
09
0>
0C
#990290000000
1!
1*
19
1>
1C
#990300000000
0!
0*
09
0>
0C
#990310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#990320000000
0!
0*
09
0>
0C
#990330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#990340000000
0!
0*
09
0>
0C
#990350000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#990360000000
0!
0*
09
0>
0C
#990370000000
1!
1*
b10 6
19
1>
1C
b10 G
#990380000000
0!
0*
09
0>
0C
#990390000000
1!
1*
b11 6
19
1>
1C
b11 G
#990400000000
0!
0*
09
0>
0C
#990410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#990420000000
0!
0*
09
0>
0C
#990430000000
1!
1*
b101 6
19
1>
1C
b101 G
#990440000000
0!
0*
09
0>
0C
#990450000000
1!
1*
b110 6
19
1>
1C
b110 G
#990460000000
0!
0*
09
0>
0C
#990470000000
1!
1*
b111 6
19
1>
1C
b111 G
#990480000000
0!
0*
09
0>
0C
#990490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#990500000000
0!
0*
09
0>
0C
#990510000000
1!
1*
b1 6
19
1>
1C
b1 G
#990520000000
0!
0*
09
0>
0C
#990530000000
1!
1*
b10 6
19
1>
1C
b10 G
#990540000000
0!
0*
09
0>
0C
#990550000000
1!
1*
b11 6
19
1>
1C
b11 G
#990560000000
0!
0*
09
0>
0C
#990570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#990580000000
0!
0*
09
0>
0C
#990590000000
1!
1*
b101 6
19
1>
1C
b101 G
#990600000000
0!
0*
09
0>
0C
#990610000000
1!
1*
b110 6
19
1>
1C
b110 G
#990620000000
0!
0*
09
0>
0C
#990630000000
1!
1*
b111 6
19
1>
1C
b111 G
#990640000000
0!
0*
09
0>
0C
#990650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#990660000000
0!
0*
09
0>
0C
#990670000000
1!
1*
b1 6
19
1>
1C
b1 G
#990680000000
0!
0*
09
0>
0C
#990690000000
1!
1*
b10 6
19
1>
1C
b10 G
#990700000000
0!
0*
09
0>
0C
#990710000000
1!
1*
b11 6
19
1>
1C
b11 G
#990720000000
0!
0*
09
0>
0C
#990730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#990740000000
0!
0*
09
0>
0C
#990750000000
1!
1*
b101 6
19
1>
1C
b101 G
#990760000000
0!
0*
09
0>
0C
#990770000000
1!
1*
b110 6
19
1>
1C
b110 G
#990780000000
0!
0*
09
0>
0C
#990790000000
1!
1*
b111 6
19
1>
1C
b111 G
#990800000000
0!
1"
0*
1+
09
1:
0>
0C
#990810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#990820000000
0!
0*
09
0>
0C
#990830000000
1!
1*
b1 6
19
1>
1C
b1 G
#990840000000
0!
0*
09
0>
0C
#990850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#990860000000
0!
0*
09
0>
0C
#990870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#990880000000
0!
0*
09
0>
0C
#990890000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#990900000000
0!
0*
09
0>
0C
#990910000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#990920000000
0!
0#
0*
0,
09
0>
0?
0C
#990930000000
1!
1*
02
19
1>
0@
0A
0B
1C
#990940000000
0!
0*
09
0>
0C
#990950000000
1!
1*
19
1>
1C
#990960000000
0!
0*
09
0>
0C
#990970000000
1!
1*
19
1>
1C
#990980000000
0!
0*
09
0>
0C
#990990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#991000000000
0!
0*
09
0>
0C
#991010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#991020000000
0!
0*
09
0>
0C
#991030000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#991040000000
0!
0*
09
0>
0C
#991050000000
1!
1*
b10 6
19
1>
1C
b10 G
#991060000000
0!
0*
09
0>
0C
#991070000000
1!
1*
b11 6
19
1>
1C
b11 G
#991080000000
0!
0*
09
0>
0C
#991090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#991100000000
0!
0*
09
0>
0C
#991110000000
1!
1*
b101 6
19
1>
1C
b101 G
#991120000000
0!
0*
09
0>
0C
#991130000000
1!
1*
b110 6
19
1>
1C
b110 G
#991140000000
0!
0*
09
0>
0C
#991150000000
1!
1*
b111 6
19
1>
1C
b111 G
#991160000000
0!
0*
09
0>
0C
#991170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#991180000000
0!
0*
09
0>
0C
#991190000000
1!
1*
b1 6
19
1>
1C
b1 G
#991200000000
0!
0*
09
0>
0C
#991210000000
1!
1*
b10 6
19
1>
1C
b10 G
#991220000000
0!
0*
09
0>
0C
#991230000000
1!
1*
b11 6
19
1>
1C
b11 G
#991240000000
0!
0*
09
0>
0C
#991250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#991260000000
0!
0*
09
0>
0C
#991270000000
1!
1*
b101 6
19
1>
1C
b101 G
#991280000000
0!
0*
09
0>
0C
#991290000000
1!
1*
b110 6
19
1>
1C
b110 G
#991300000000
0!
0*
09
0>
0C
#991310000000
1!
1*
b111 6
19
1>
1C
b111 G
#991320000000
0!
0*
09
0>
0C
#991330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#991340000000
0!
0*
09
0>
0C
#991350000000
1!
1*
b1 6
19
1>
1C
b1 G
#991360000000
0!
0*
09
0>
0C
#991370000000
1!
1*
b10 6
19
1>
1C
b10 G
#991380000000
0!
0*
09
0>
0C
#991390000000
1!
1*
b11 6
19
1>
1C
b11 G
#991400000000
0!
0*
09
0>
0C
#991410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#991420000000
0!
0*
09
0>
0C
#991430000000
1!
1*
b101 6
19
1>
1C
b101 G
#991440000000
0!
0*
09
0>
0C
#991450000000
1!
1*
b110 6
19
1>
1C
b110 G
#991460000000
0!
0*
09
0>
0C
#991470000000
1!
1*
b111 6
19
1>
1C
b111 G
#991480000000
0!
1"
0*
1+
09
1:
0>
0C
#991490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#991500000000
0!
0*
09
0>
0C
#991510000000
1!
1*
b1 6
19
1>
1C
b1 G
#991520000000
0!
0*
09
0>
0C
#991530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#991540000000
0!
0*
09
0>
0C
#991550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#991560000000
0!
0*
09
0>
0C
#991570000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#991580000000
0!
0*
09
0>
0C
#991590000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#991600000000
0!
0#
0*
0,
09
0>
0?
0C
#991610000000
1!
1*
02
19
1>
0@
0A
0B
1C
#991620000000
0!
0*
09
0>
0C
#991630000000
1!
1*
19
1>
1C
#991640000000
0!
0*
09
0>
0C
#991650000000
1!
1*
19
1>
1C
#991660000000
0!
0*
09
0>
0C
#991670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#991680000000
0!
0*
09
0>
0C
#991690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#991700000000
0!
0*
09
0>
0C
#991710000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#991720000000
0!
0*
09
0>
0C
#991730000000
1!
1*
b10 6
19
1>
1C
b10 G
#991740000000
0!
0*
09
0>
0C
#991750000000
1!
1*
b11 6
19
1>
1C
b11 G
#991760000000
0!
0*
09
0>
0C
#991770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#991780000000
0!
0*
09
0>
0C
#991790000000
1!
1*
b101 6
19
1>
1C
b101 G
#991800000000
0!
0*
09
0>
0C
#991810000000
1!
1*
b110 6
19
1>
1C
b110 G
#991820000000
0!
0*
09
0>
0C
#991830000000
1!
1*
b111 6
19
1>
1C
b111 G
#991840000000
0!
0*
09
0>
0C
#991850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#991860000000
0!
0*
09
0>
0C
#991870000000
1!
1*
b1 6
19
1>
1C
b1 G
#991880000000
0!
0*
09
0>
0C
#991890000000
1!
1*
b10 6
19
1>
1C
b10 G
#991900000000
0!
0*
09
0>
0C
#991910000000
1!
1*
b11 6
19
1>
1C
b11 G
#991920000000
0!
0*
09
0>
0C
#991930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#991940000000
0!
0*
09
0>
0C
#991950000000
1!
1*
b101 6
19
1>
1C
b101 G
#991960000000
0!
0*
09
0>
0C
#991970000000
1!
1*
b110 6
19
1>
1C
b110 G
#991980000000
0!
0*
09
0>
0C
#991990000000
1!
1*
b111 6
19
1>
1C
b111 G
#992000000000
0!
0*
09
0>
0C
#992010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#992020000000
0!
0*
09
0>
0C
#992030000000
1!
1*
b1 6
19
1>
1C
b1 G
#992040000000
0!
0*
09
0>
0C
#992050000000
1!
1*
b10 6
19
1>
1C
b10 G
#992060000000
0!
0*
09
0>
0C
#992070000000
1!
1*
b11 6
19
1>
1C
b11 G
#992080000000
0!
0*
09
0>
0C
#992090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#992100000000
0!
0*
09
0>
0C
#992110000000
1!
1*
b101 6
19
1>
1C
b101 G
#992120000000
0!
0*
09
0>
0C
#992130000000
1!
1*
b110 6
19
1>
1C
b110 G
#992140000000
0!
0*
09
0>
0C
#992150000000
1!
1*
b111 6
19
1>
1C
b111 G
#992160000000
0!
1"
0*
1+
09
1:
0>
0C
#992170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#992180000000
0!
0*
09
0>
0C
#992190000000
1!
1*
b1 6
19
1>
1C
b1 G
#992200000000
0!
0*
09
0>
0C
#992210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#992220000000
0!
0*
09
0>
0C
#992230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#992240000000
0!
0*
09
0>
0C
#992250000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#992260000000
0!
0*
09
0>
0C
#992270000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#992280000000
0!
0#
0*
0,
09
0>
0?
0C
#992290000000
1!
1*
02
19
1>
0@
0A
0B
1C
#992300000000
0!
0*
09
0>
0C
#992310000000
1!
1*
19
1>
1C
#992320000000
0!
0*
09
0>
0C
#992330000000
1!
1*
19
1>
1C
#992340000000
0!
0*
09
0>
0C
#992350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#992360000000
0!
0*
09
0>
0C
#992370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#992380000000
0!
0*
09
0>
0C
#992390000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#992400000000
0!
0*
09
0>
0C
#992410000000
1!
1*
b10 6
19
1>
1C
b10 G
#992420000000
0!
0*
09
0>
0C
#992430000000
1!
1*
b11 6
19
1>
1C
b11 G
#992440000000
0!
0*
09
0>
0C
#992450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#992460000000
0!
0*
09
0>
0C
#992470000000
1!
1*
b101 6
19
1>
1C
b101 G
#992480000000
0!
0*
09
0>
0C
#992490000000
1!
1*
b110 6
19
1>
1C
b110 G
#992500000000
0!
0*
09
0>
0C
#992510000000
1!
1*
b111 6
19
1>
1C
b111 G
#992520000000
0!
0*
09
0>
0C
#992530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#992540000000
0!
0*
09
0>
0C
#992550000000
1!
1*
b1 6
19
1>
1C
b1 G
#992560000000
0!
0*
09
0>
0C
#992570000000
1!
1*
b10 6
19
1>
1C
b10 G
#992580000000
0!
0*
09
0>
0C
#992590000000
1!
1*
b11 6
19
1>
1C
b11 G
#992600000000
0!
0*
09
0>
0C
#992610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#992620000000
0!
0*
09
0>
0C
#992630000000
1!
1*
b101 6
19
1>
1C
b101 G
#992640000000
0!
0*
09
0>
0C
#992650000000
1!
1*
b110 6
19
1>
1C
b110 G
#992660000000
0!
0*
09
0>
0C
#992670000000
1!
1*
b111 6
19
1>
1C
b111 G
#992680000000
0!
0*
09
0>
0C
#992690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#992700000000
0!
0*
09
0>
0C
#992710000000
1!
1*
b1 6
19
1>
1C
b1 G
#992720000000
0!
0*
09
0>
0C
#992730000000
1!
1*
b10 6
19
1>
1C
b10 G
#992740000000
0!
0*
09
0>
0C
#992750000000
1!
1*
b11 6
19
1>
1C
b11 G
#992760000000
0!
0*
09
0>
0C
#992770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#992780000000
0!
0*
09
0>
0C
#992790000000
1!
1*
b101 6
19
1>
1C
b101 G
#992800000000
0!
0*
09
0>
0C
#992810000000
1!
1*
b110 6
19
1>
1C
b110 G
#992820000000
0!
0*
09
0>
0C
#992830000000
1!
1*
b111 6
19
1>
1C
b111 G
#992840000000
0!
1"
0*
1+
09
1:
0>
0C
#992850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#992860000000
0!
0*
09
0>
0C
#992870000000
1!
1*
b1 6
19
1>
1C
b1 G
#992880000000
0!
0*
09
0>
0C
#992890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#992900000000
0!
0*
09
0>
0C
#992910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#992920000000
0!
0*
09
0>
0C
#992930000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#992940000000
0!
0*
09
0>
0C
#992950000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#992960000000
0!
0#
0*
0,
09
0>
0?
0C
#992970000000
1!
1*
02
19
1>
0@
0A
0B
1C
#992980000000
0!
0*
09
0>
0C
#992990000000
1!
1*
19
1>
1C
#993000000000
0!
0*
09
0>
0C
#993010000000
1!
1*
19
1>
1C
#993020000000
0!
0*
09
0>
0C
#993030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#993040000000
0!
0*
09
0>
0C
#993050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#993060000000
0!
0*
09
0>
0C
#993070000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#993080000000
0!
0*
09
0>
0C
#993090000000
1!
1*
b10 6
19
1>
1C
b10 G
#993100000000
0!
0*
09
0>
0C
#993110000000
1!
1*
b11 6
19
1>
1C
b11 G
#993120000000
0!
0*
09
0>
0C
#993130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#993140000000
0!
0*
09
0>
0C
#993150000000
1!
1*
b101 6
19
1>
1C
b101 G
#993160000000
0!
0*
09
0>
0C
#993170000000
1!
1*
b110 6
19
1>
1C
b110 G
#993180000000
0!
0*
09
0>
0C
#993190000000
1!
1*
b111 6
19
1>
1C
b111 G
#993200000000
0!
0*
09
0>
0C
#993210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#993220000000
0!
0*
09
0>
0C
#993230000000
1!
1*
b1 6
19
1>
1C
b1 G
#993240000000
0!
0*
09
0>
0C
#993250000000
1!
1*
b10 6
19
1>
1C
b10 G
#993260000000
0!
0*
09
0>
0C
#993270000000
1!
1*
b11 6
19
1>
1C
b11 G
#993280000000
0!
0*
09
0>
0C
#993290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#993300000000
0!
0*
09
0>
0C
#993310000000
1!
1*
b101 6
19
1>
1C
b101 G
#993320000000
0!
0*
09
0>
0C
#993330000000
1!
1*
b110 6
19
1>
1C
b110 G
#993340000000
0!
0*
09
0>
0C
#993350000000
1!
1*
b111 6
19
1>
1C
b111 G
#993360000000
0!
0*
09
0>
0C
#993370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#993380000000
0!
0*
09
0>
0C
#993390000000
1!
1*
b1 6
19
1>
1C
b1 G
#993400000000
0!
0*
09
0>
0C
#993410000000
1!
1*
b10 6
19
1>
1C
b10 G
#993420000000
0!
0*
09
0>
0C
#993430000000
1!
1*
b11 6
19
1>
1C
b11 G
#993440000000
0!
0*
09
0>
0C
#993450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#993460000000
0!
0*
09
0>
0C
#993470000000
1!
1*
b101 6
19
1>
1C
b101 G
#993480000000
0!
0*
09
0>
0C
#993490000000
1!
1*
b110 6
19
1>
1C
b110 G
#993500000000
0!
0*
09
0>
0C
#993510000000
1!
1*
b111 6
19
1>
1C
b111 G
#993520000000
0!
1"
0*
1+
09
1:
0>
0C
#993530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#993540000000
0!
0*
09
0>
0C
#993550000000
1!
1*
b1 6
19
1>
1C
b1 G
#993560000000
0!
0*
09
0>
0C
#993570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#993580000000
0!
0*
09
0>
0C
#993590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#993600000000
0!
0*
09
0>
0C
#993610000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#993620000000
0!
0*
09
0>
0C
#993630000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#993640000000
0!
0#
0*
0,
09
0>
0?
0C
#993650000000
1!
1*
02
19
1>
0@
0A
0B
1C
#993660000000
0!
0*
09
0>
0C
#993670000000
1!
1*
19
1>
1C
#993680000000
0!
0*
09
0>
0C
#993690000000
1!
1*
19
1>
1C
#993700000000
0!
0*
09
0>
0C
#993710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#993720000000
0!
0*
09
0>
0C
#993730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#993740000000
0!
0*
09
0>
0C
#993750000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#993760000000
0!
0*
09
0>
0C
#993770000000
1!
1*
b10 6
19
1>
1C
b10 G
#993780000000
0!
0*
09
0>
0C
#993790000000
1!
1*
b11 6
19
1>
1C
b11 G
#993800000000
0!
0*
09
0>
0C
#993810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#993820000000
0!
0*
09
0>
0C
#993830000000
1!
1*
b101 6
19
1>
1C
b101 G
#993840000000
0!
0*
09
0>
0C
#993850000000
1!
1*
b110 6
19
1>
1C
b110 G
#993860000000
0!
0*
09
0>
0C
#993870000000
1!
1*
b111 6
19
1>
1C
b111 G
#993880000000
0!
0*
09
0>
0C
#993890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#993900000000
0!
0*
09
0>
0C
#993910000000
1!
1*
b1 6
19
1>
1C
b1 G
#993920000000
0!
0*
09
0>
0C
#993930000000
1!
1*
b10 6
19
1>
1C
b10 G
#993940000000
0!
0*
09
0>
0C
#993950000000
1!
1*
b11 6
19
1>
1C
b11 G
#993960000000
0!
0*
09
0>
0C
#993970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#993980000000
0!
0*
09
0>
0C
#993990000000
1!
1*
b101 6
19
1>
1C
b101 G
#994000000000
0!
0*
09
0>
0C
#994010000000
1!
1*
b110 6
19
1>
1C
b110 G
#994020000000
0!
0*
09
0>
0C
#994030000000
1!
1*
b111 6
19
1>
1C
b111 G
#994040000000
0!
0*
09
0>
0C
#994050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#994060000000
0!
0*
09
0>
0C
#994070000000
1!
1*
b1 6
19
1>
1C
b1 G
#994080000000
0!
0*
09
0>
0C
#994090000000
1!
1*
b10 6
19
1>
1C
b10 G
#994100000000
0!
0*
09
0>
0C
#994110000000
1!
1*
b11 6
19
1>
1C
b11 G
#994120000000
0!
0*
09
0>
0C
#994130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#994140000000
0!
0*
09
0>
0C
#994150000000
1!
1*
b101 6
19
1>
1C
b101 G
#994160000000
0!
0*
09
0>
0C
#994170000000
1!
1*
b110 6
19
1>
1C
b110 G
#994180000000
0!
0*
09
0>
0C
#994190000000
1!
1*
b111 6
19
1>
1C
b111 G
#994200000000
0!
1"
0*
1+
09
1:
0>
0C
#994210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#994220000000
0!
0*
09
0>
0C
#994230000000
1!
1*
b1 6
19
1>
1C
b1 G
#994240000000
0!
0*
09
0>
0C
#994250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#994260000000
0!
0*
09
0>
0C
#994270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#994280000000
0!
0*
09
0>
0C
#994290000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#994300000000
0!
0*
09
0>
0C
#994310000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#994320000000
0!
0#
0*
0,
09
0>
0?
0C
#994330000000
1!
1*
02
19
1>
0@
0A
0B
1C
#994340000000
0!
0*
09
0>
0C
#994350000000
1!
1*
19
1>
1C
#994360000000
0!
0*
09
0>
0C
#994370000000
1!
1*
19
1>
1C
#994380000000
0!
0*
09
0>
0C
#994390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#994400000000
0!
0*
09
0>
0C
#994410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#994420000000
0!
0*
09
0>
0C
#994430000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#994440000000
0!
0*
09
0>
0C
#994450000000
1!
1*
b10 6
19
1>
1C
b10 G
#994460000000
0!
0*
09
0>
0C
#994470000000
1!
1*
b11 6
19
1>
1C
b11 G
#994480000000
0!
0*
09
0>
0C
#994490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#994500000000
0!
0*
09
0>
0C
#994510000000
1!
1*
b101 6
19
1>
1C
b101 G
#994520000000
0!
0*
09
0>
0C
#994530000000
1!
1*
b110 6
19
1>
1C
b110 G
#994540000000
0!
0*
09
0>
0C
#994550000000
1!
1*
b111 6
19
1>
1C
b111 G
#994560000000
0!
0*
09
0>
0C
#994570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#994580000000
0!
0*
09
0>
0C
#994590000000
1!
1*
b1 6
19
1>
1C
b1 G
#994600000000
0!
0*
09
0>
0C
#994610000000
1!
1*
b10 6
19
1>
1C
b10 G
#994620000000
0!
0*
09
0>
0C
#994630000000
1!
1*
b11 6
19
1>
1C
b11 G
#994640000000
0!
0*
09
0>
0C
#994650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#994660000000
0!
0*
09
0>
0C
#994670000000
1!
1*
b101 6
19
1>
1C
b101 G
#994680000000
0!
0*
09
0>
0C
#994690000000
1!
1*
b110 6
19
1>
1C
b110 G
#994700000000
0!
0*
09
0>
0C
#994710000000
1!
1*
b111 6
19
1>
1C
b111 G
#994720000000
0!
0*
09
0>
0C
#994730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#994740000000
0!
0*
09
0>
0C
#994750000000
1!
1*
b1 6
19
1>
1C
b1 G
#994760000000
0!
0*
09
0>
0C
#994770000000
1!
1*
b10 6
19
1>
1C
b10 G
#994780000000
0!
0*
09
0>
0C
#994790000000
1!
1*
b11 6
19
1>
1C
b11 G
#994800000000
0!
0*
09
0>
0C
#994810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#994820000000
0!
0*
09
0>
0C
#994830000000
1!
1*
b101 6
19
1>
1C
b101 G
#994840000000
0!
0*
09
0>
0C
#994850000000
1!
1*
b110 6
19
1>
1C
b110 G
#994860000000
0!
0*
09
0>
0C
#994870000000
1!
1*
b111 6
19
1>
1C
b111 G
#994880000000
0!
1"
0*
1+
09
1:
0>
0C
#994890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#994900000000
0!
0*
09
0>
0C
#994910000000
1!
1*
b1 6
19
1>
1C
b1 G
#994920000000
0!
0*
09
0>
0C
#994930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#994940000000
0!
0*
09
0>
0C
#994950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#994960000000
0!
0*
09
0>
0C
#994970000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#994980000000
0!
0*
09
0>
0C
#994990000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#995000000000
0!
0#
0*
0,
09
0>
0?
0C
#995010000000
1!
1*
02
19
1>
0@
0A
0B
1C
#995020000000
0!
0*
09
0>
0C
#995030000000
1!
1*
19
1>
1C
#995040000000
0!
0*
09
0>
0C
#995050000000
1!
1*
19
1>
1C
#995060000000
0!
0*
09
0>
0C
#995070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#995080000000
0!
0*
09
0>
0C
#995090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#995100000000
0!
0*
09
0>
0C
#995110000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#995120000000
0!
0*
09
0>
0C
#995130000000
1!
1*
b10 6
19
1>
1C
b10 G
#995140000000
0!
0*
09
0>
0C
#995150000000
1!
1*
b11 6
19
1>
1C
b11 G
#995160000000
0!
0*
09
0>
0C
#995170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#995180000000
0!
0*
09
0>
0C
#995190000000
1!
1*
b101 6
19
1>
1C
b101 G
#995200000000
0!
0*
09
0>
0C
#995210000000
1!
1*
b110 6
19
1>
1C
b110 G
#995220000000
0!
0*
09
0>
0C
#995230000000
1!
1*
b111 6
19
1>
1C
b111 G
#995240000000
0!
0*
09
0>
0C
#995250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#995260000000
0!
0*
09
0>
0C
#995270000000
1!
1*
b1 6
19
1>
1C
b1 G
#995280000000
0!
0*
09
0>
0C
#995290000000
1!
1*
b10 6
19
1>
1C
b10 G
#995300000000
0!
0*
09
0>
0C
#995310000000
1!
1*
b11 6
19
1>
1C
b11 G
#995320000000
0!
0*
09
0>
0C
#995330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#995340000000
0!
0*
09
0>
0C
#995350000000
1!
1*
b101 6
19
1>
1C
b101 G
#995360000000
0!
0*
09
0>
0C
#995370000000
1!
1*
b110 6
19
1>
1C
b110 G
#995380000000
0!
0*
09
0>
0C
#995390000000
1!
1*
b111 6
19
1>
1C
b111 G
#995400000000
0!
0*
09
0>
0C
#995410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#995420000000
0!
0*
09
0>
0C
#995430000000
1!
1*
b1 6
19
1>
1C
b1 G
#995440000000
0!
0*
09
0>
0C
#995450000000
1!
1*
b10 6
19
1>
1C
b10 G
#995460000000
0!
0*
09
0>
0C
#995470000000
1!
1*
b11 6
19
1>
1C
b11 G
#995480000000
0!
0*
09
0>
0C
#995490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#995500000000
0!
0*
09
0>
0C
#995510000000
1!
1*
b101 6
19
1>
1C
b101 G
#995520000000
0!
0*
09
0>
0C
#995530000000
1!
1*
b110 6
19
1>
1C
b110 G
#995540000000
0!
0*
09
0>
0C
#995550000000
1!
1*
b111 6
19
1>
1C
b111 G
#995560000000
0!
1"
0*
1+
09
1:
0>
0C
#995570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#995580000000
0!
0*
09
0>
0C
#995590000000
1!
1*
b1 6
19
1>
1C
b1 G
#995600000000
0!
0*
09
0>
0C
#995610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#995620000000
0!
0*
09
0>
0C
#995630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#995640000000
0!
0*
09
0>
0C
#995650000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#995660000000
0!
0*
09
0>
0C
#995670000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#995680000000
0!
0#
0*
0,
09
0>
0?
0C
#995690000000
1!
1*
02
19
1>
0@
0A
0B
1C
#995700000000
0!
0*
09
0>
0C
#995710000000
1!
1*
19
1>
1C
#995720000000
0!
0*
09
0>
0C
#995730000000
1!
1*
19
1>
1C
#995740000000
0!
0*
09
0>
0C
#995750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#995760000000
0!
0*
09
0>
0C
#995770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#995780000000
0!
0*
09
0>
0C
#995790000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#995800000000
0!
0*
09
0>
0C
#995810000000
1!
1*
b10 6
19
1>
1C
b10 G
#995820000000
0!
0*
09
0>
0C
#995830000000
1!
1*
b11 6
19
1>
1C
b11 G
#995840000000
0!
0*
09
0>
0C
#995850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#995860000000
0!
0*
09
0>
0C
#995870000000
1!
1*
b101 6
19
1>
1C
b101 G
#995880000000
0!
0*
09
0>
0C
#995890000000
1!
1*
b110 6
19
1>
1C
b110 G
#995900000000
0!
0*
09
0>
0C
#995910000000
1!
1*
b111 6
19
1>
1C
b111 G
#995920000000
0!
0*
09
0>
0C
#995930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#995940000000
0!
0*
09
0>
0C
#995950000000
1!
1*
b1 6
19
1>
1C
b1 G
#995960000000
0!
0*
09
0>
0C
#995970000000
1!
1*
b10 6
19
1>
1C
b10 G
#995980000000
0!
0*
09
0>
0C
#995990000000
1!
1*
b11 6
19
1>
1C
b11 G
#996000000000
0!
0*
09
0>
0C
#996010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#996020000000
0!
0*
09
0>
0C
#996030000000
1!
1*
b101 6
19
1>
1C
b101 G
#996040000000
0!
0*
09
0>
0C
#996050000000
1!
1*
b110 6
19
1>
1C
b110 G
#996060000000
0!
0*
09
0>
0C
#996070000000
1!
1*
b111 6
19
1>
1C
b111 G
#996080000000
0!
0*
09
0>
0C
#996090000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#996100000000
0!
0*
09
0>
0C
#996110000000
1!
1*
b1 6
19
1>
1C
b1 G
#996120000000
0!
0*
09
0>
0C
#996130000000
1!
1*
b10 6
19
1>
1C
b10 G
#996140000000
0!
0*
09
0>
0C
#996150000000
1!
1*
b11 6
19
1>
1C
b11 G
#996160000000
0!
0*
09
0>
0C
#996170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#996180000000
0!
0*
09
0>
0C
#996190000000
1!
1*
b101 6
19
1>
1C
b101 G
#996200000000
0!
0*
09
0>
0C
#996210000000
1!
1*
b110 6
19
1>
1C
b110 G
#996220000000
0!
0*
09
0>
0C
#996230000000
1!
1*
b111 6
19
1>
1C
b111 G
#996240000000
0!
1"
0*
1+
09
1:
0>
0C
#996250000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#996260000000
0!
0*
09
0>
0C
#996270000000
1!
1*
b1 6
19
1>
1C
b1 G
#996280000000
0!
0*
09
0>
0C
#996290000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#996300000000
0!
0*
09
0>
0C
#996310000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#996320000000
0!
0*
09
0>
0C
#996330000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#996340000000
0!
0*
09
0>
0C
#996350000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#996360000000
0!
0#
0*
0,
09
0>
0?
0C
#996370000000
1!
1*
02
19
1>
0@
0A
0B
1C
#996380000000
0!
0*
09
0>
0C
#996390000000
1!
1*
19
1>
1C
#996400000000
0!
0*
09
0>
0C
#996410000000
1!
1*
19
1>
1C
#996420000000
0!
0*
09
0>
0C
#996430000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#996440000000
0!
0*
09
0>
0C
#996450000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#996460000000
0!
0*
09
0>
0C
#996470000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#996480000000
0!
0*
09
0>
0C
#996490000000
1!
1*
b10 6
19
1>
1C
b10 G
#996500000000
0!
0*
09
0>
0C
#996510000000
1!
1*
b11 6
19
1>
1C
b11 G
#996520000000
0!
0*
09
0>
0C
#996530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#996540000000
0!
0*
09
0>
0C
#996550000000
1!
1*
b101 6
19
1>
1C
b101 G
#996560000000
0!
0*
09
0>
0C
#996570000000
1!
1*
b110 6
19
1>
1C
b110 G
#996580000000
0!
0*
09
0>
0C
#996590000000
1!
1*
b111 6
19
1>
1C
b111 G
#996600000000
0!
0*
09
0>
0C
#996610000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#996620000000
0!
0*
09
0>
0C
#996630000000
1!
1*
b1 6
19
1>
1C
b1 G
#996640000000
0!
0*
09
0>
0C
#996650000000
1!
1*
b10 6
19
1>
1C
b10 G
#996660000000
0!
0*
09
0>
0C
#996670000000
1!
1*
b11 6
19
1>
1C
b11 G
#996680000000
0!
0*
09
0>
0C
#996690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#996700000000
0!
0*
09
0>
0C
#996710000000
1!
1*
b101 6
19
1>
1C
b101 G
#996720000000
0!
0*
09
0>
0C
#996730000000
1!
1*
b110 6
19
1>
1C
b110 G
#996740000000
0!
0*
09
0>
0C
#996750000000
1!
1*
b111 6
19
1>
1C
b111 G
#996760000000
0!
0*
09
0>
0C
#996770000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#996780000000
0!
0*
09
0>
0C
#996790000000
1!
1*
b1 6
19
1>
1C
b1 G
#996800000000
0!
0*
09
0>
0C
#996810000000
1!
1*
b10 6
19
1>
1C
b10 G
#996820000000
0!
0*
09
0>
0C
#996830000000
1!
1*
b11 6
19
1>
1C
b11 G
#996840000000
0!
0*
09
0>
0C
#996850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#996860000000
0!
0*
09
0>
0C
#996870000000
1!
1*
b101 6
19
1>
1C
b101 G
#996880000000
0!
0*
09
0>
0C
#996890000000
1!
1*
b110 6
19
1>
1C
b110 G
#996900000000
0!
0*
09
0>
0C
#996910000000
1!
1*
b111 6
19
1>
1C
b111 G
#996920000000
0!
1"
0*
1+
09
1:
0>
0C
#996930000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#996940000000
0!
0*
09
0>
0C
#996950000000
1!
1*
b1 6
19
1>
1C
b1 G
#996960000000
0!
0*
09
0>
0C
#996970000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#996980000000
0!
0*
09
0>
0C
#996990000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#997000000000
0!
0*
09
0>
0C
#997010000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#997020000000
0!
0*
09
0>
0C
#997030000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#997040000000
0!
0#
0*
0,
09
0>
0?
0C
#997050000000
1!
1*
02
19
1>
0@
0A
0B
1C
#997060000000
0!
0*
09
0>
0C
#997070000000
1!
1*
19
1>
1C
#997080000000
0!
0*
09
0>
0C
#997090000000
1!
1*
19
1>
1C
#997100000000
0!
0*
09
0>
0C
#997110000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#997120000000
0!
0*
09
0>
0C
#997130000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#997140000000
0!
0*
09
0>
0C
#997150000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#997160000000
0!
0*
09
0>
0C
#997170000000
1!
1*
b10 6
19
1>
1C
b10 G
#997180000000
0!
0*
09
0>
0C
#997190000000
1!
1*
b11 6
19
1>
1C
b11 G
#997200000000
0!
0*
09
0>
0C
#997210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#997220000000
0!
0*
09
0>
0C
#997230000000
1!
1*
b101 6
19
1>
1C
b101 G
#997240000000
0!
0*
09
0>
0C
#997250000000
1!
1*
b110 6
19
1>
1C
b110 G
#997260000000
0!
0*
09
0>
0C
#997270000000
1!
1*
b111 6
19
1>
1C
b111 G
#997280000000
0!
0*
09
0>
0C
#997290000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#997300000000
0!
0*
09
0>
0C
#997310000000
1!
1*
b1 6
19
1>
1C
b1 G
#997320000000
0!
0*
09
0>
0C
#997330000000
1!
1*
b10 6
19
1>
1C
b10 G
#997340000000
0!
0*
09
0>
0C
#997350000000
1!
1*
b11 6
19
1>
1C
b11 G
#997360000000
0!
0*
09
0>
0C
#997370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#997380000000
0!
0*
09
0>
0C
#997390000000
1!
1*
b101 6
19
1>
1C
b101 G
#997400000000
0!
0*
09
0>
0C
#997410000000
1!
1*
b110 6
19
1>
1C
b110 G
#997420000000
0!
0*
09
0>
0C
#997430000000
1!
1*
b111 6
19
1>
1C
b111 G
#997440000000
0!
0*
09
0>
0C
#997450000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#997460000000
0!
0*
09
0>
0C
#997470000000
1!
1*
b1 6
19
1>
1C
b1 G
#997480000000
0!
0*
09
0>
0C
#997490000000
1!
1*
b10 6
19
1>
1C
b10 G
#997500000000
0!
0*
09
0>
0C
#997510000000
1!
1*
b11 6
19
1>
1C
b11 G
#997520000000
0!
0*
09
0>
0C
#997530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#997540000000
0!
0*
09
0>
0C
#997550000000
1!
1*
b101 6
19
1>
1C
b101 G
#997560000000
0!
0*
09
0>
0C
#997570000000
1!
1*
b110 6
19
1>
1C
b110 G
#997580000000
0!
0*
09
0>
0C
#997590000000
1!
1*
b111 6
19
1>
1C
b111 G
#997600000000
0!
1"
0*
1+
09
1:
0>
0C
#997610000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#997620000000
0!
0*
09
0>
0C
#997630000000
1!
1*
b1 6
19
1>
1C
b1 G
#997640000000
0!
0*
09
0>
0C
#997650000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#997660000000
0!
0*
09
0>
0C
#997670000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#997680000000
0!
0*
09
0>
0C
#997690000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#997700000000
0!
0*
09
0>
0C
#997710000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#997720000000
0!
0#
0*
0,
09
0>
0?
0C
#997730000000
1!
1*
02
19
1>
0@
0A
0B
1C
#997740000000
0!
0*
09
0>
0C
#997750000000
1!
1*
19
1>
1C
#997760000000
0!
0*
09
0>
0C
#997770000000
1!
1*
19
1>
1C
#997780000000
0!
0*
09
0>
0C
#997790000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#997800000000
0!
0*
09
0>
0C
#997810000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#997820000000
0!
0*
09
0>
0C
#997830000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#997840000000
0!
0*
09
0>
0C
#997850000000
1!
1*
b10 6
19
1>
1C
b10 G
#997860000000
0!
0*
09
0>
0C
#997870000000
1!
1*
b11 6
19
1>
1C
b11 G
#997880000000
0!
0*
09
0>
0C
#997890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#997900000000
0!
0*
09
0>
0C
#997910000000
1!
1*
b101 6
19
1>
1C
b101 G
#997920000000
0!
0*
09
0>
0C
#997930000000
1!
1*
b110 6
19
1>
1C
b110 G
#997940000000
0!
0*
09
0>
0C
#997950000000
1!
1*
b111 6
19
1>
1C
b111 G
#997960000000
0!
0*
09
0>
0C
#997970000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#997980000000
0!
0*
09
0>
0C
#997990000000
1!
1*
b1 6
19
1>
1C
b1 G
#998000000000
0!
0*
09
0>
0C
#998010000000
1!
1*
b10 6
19
1>
1C
b10 G
#998020000000
0!
0*
09
0>
0C
#998030000000
1!
1*
b11 6
19
1>
1C
b11 G
#998040000000
0!
0*
09
0>
0C
#998050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#998060000000
0!
0*
09
0>
0C
#998070000000
1!
1*
b101 6
19
1>
1C
b101 G
#998080000000
0!
0*
09
0>
0C
#998090000000
1!
1*
b110 6
19
1>
1C
b110 G
#998100000000
0!
0*
09
0>
0C
#998110000000
1!
1*
b111 6
19
1>
1C
b111 G
#998120000000
0!
0*
09
0>
0C
#998130000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#998140000000
0!
0*
09
0>
0C
#998150000000
1!
1*
b1 6
19
1>
1C
b1 G
#998160000000
0!
0*
09
0>
0C
#998170000000
1!
1*
b10 6
19
1>
1C
b10 G
#998180000000
0!
0*
09
0>
0C
#998190000000
1!
1*
b11 6
19
1>
1C
b11 G
#998200000000
0!
0*
09
0>
0C
#998210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#998220000000
0!
0*
09
0>
0C
#998230000000
1!
1*
b101 6
19
1>
1C
b101 G
#998240000000
0!
0*
09
0>
0C
#998250000000
1!
1*
b110 6
19
1>
1C
b110 G
#998260000000
0!
0*
09
0>
0C
#998270000000
1!
1*
b111 6
19
1>
1C
b111 G
#998280000000
0!
1"
0*
1+
09
1:
0>
0C
#998290000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#998300000000
0!
0*
09
0>
0C
#998310000000
1!
1*
b1 6
19
1>
1C
b1 G
#998320000000
0!
0*
09
0>
0C
#998330000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#998340000000
0!
0*
09
0>
0C
#998350000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#998360000000
0!
0*
09
0>
0C
#998370000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#998380000000
0!
0*
09
0>
0C
#998390000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#998400000000
0!
0#
0*
0,
09
0>
0?
0C
#998410000000
1!
1*
02
19
1>
0@
0A
0B
1C
#998420000000
0!
0*
09
0>
0C
#998430000000
1!
1*
19
1>
1C
#998440000000
0!
0*
09
0>
0C
#998450000000
1!
1*
19
1>
1C
#998460000000
0!
0*
09
0>
0C
#998470000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#998480000000
0!
0*
09
0>
0C
#998490000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#998500000000
0!
0*
09
0>
0C
#998510000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#998520000000
0!
0*
09
0>
0C
#998530000000
1!
1*
b10 6
19
1>
1C
b10 G
#998540000000
0!
0*
09
0>
0C
#998550000000
1!
1*
b11 6
19
1>
1C
b11 G
#998560000000
0!
0*
09
0>
0C
#998570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#998580000000
0!
0*
09
0>
0C
#998590000000
1!
1*
b101 6
19
1>
1C
b101 G
#998600000000
0!
0*
09
0>
0C
#998610000000
1!
1*
b110 6
19
1>
1C
b110 G
#998620000000
0!
0*
09
0>
0C
#998630000000
1!
1*
b111 6
19
1>
1C
b111 G
#998640000000
0!
0*
09
0>
0C
#998650000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#998660000000
0!
0*
09
0>
0C
#998670000000
1!
1*
b1 6
19
1>
1C
b1 G
#998680000000
0!
0*
09
0>
0C
#998690000000
1!
1*
b10 6
19
1>
1C
b10 G
#998700000000
0!
0*
09
0>
0C
#998710000000
1!
1*
b11 6
19
1>
1C
b11 G
#998720000000
0!
0*
09
0>
0C
#998730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#998740000000
0!
0*
09
0>
0C
#998750000000
1!
1*
b101 6
19
1>
1C
b101 G
#998760000000
0!
0*
09
0>
0C
#998770000000
1!
1*
b110 6
19
1>
1C
b110 G
#998780000000
0!
0*
09
0>
0C
#998790000000
1!
1*
b111 6
19
1>
1C
b111 G
#998800000000
0!
0*
09
0>
0C
#998810000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#998820000000
0!
0*
09
0>
0C
#998830000000
1!
1*
b1 6
19
1>
1C
b1 G
#998840000000
0!
0*
09
0>
0C
#998850000000
1!
1*
b10 6
19
1>
1C
b10 G
#998860000000
0!
0*
09
0>
0C
#998870000000
1!
1*
b11 6
19
1>
1C
b11 G
#998880000000
0!
0*
09
0>
0C
#998890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#998900000000
0!
0*
09
0>
0C
#998910000000
1!
1*
b101 6
19
1>
1C
b101 G
#998920000000
0!
0*
09
0>
0C
#998930000000
1!
1*
b110 6
19
1>
1C
b110 G
#998940000000
0!
0*
09
0>
0C
#998950000000
1!
1*
b111 6
19
1>
1C
b111 G
#998960000000
0!
1"
0*
1+
09
1:
0>
0C
#998970000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#998980000000
0!
0*
09
0>
0C
#998990000000
1!
1*
b1 6
19
1>
1C
b1 G
#999000000000
0!
0*
09
0>
0C
#999010000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#999020000000
0!
0*
09
0>
0C
#999030000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#999040000000
0!
0*
09
0>
0C
#999050000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#999060000000
0!
0*
09
0>
0C
#999070000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#999080000000
0!
0#
0*
0,
09
0>
0?
0C
#999090000000
1!
1*
02
19
1>
0@
0A
0B
1C
#999100000000
0!
0*
09
0>
0C
#999110000000
1!
1*
19
1>
1C
#999120000000
0!
0*
09
0>
0C
#999130000000
1!
1*
19
1>
1C
#999140000000
0!
0*
09
0>
0C
#999150000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#999160000000
0!
0*
09
0>
0C
#999170000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#999180000000
0!
0*
09
0>
0C
#999190000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#999200000000
0!
0*
09
0>
0C
#999210000000
1!
1*
b10 6
19
1>
1C
b10 G
#999220000000
0!
0*
09
0>
0C
#999230000000
1!
1*
b11 6
19
1>
1C
b11 G
#999240000000
0!
0*
09
0>
0C
#999250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#999260000000
0!
0*
09
0>
0C
#999270000000
1!
1*
b101 6
19
1>
1C
b101 G
#999280000000
0!
0*
09
0>
0C
#999290000000
1!
1*
b110 6
19
1>
1C
b110 G
#999300000000
0!
0*
09
0>
0C
#999310000000
1!
1*
b111 6
19
1>
1C
b111 G
#999320000000
0!
0*
09
0>
0C
#999330000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#999340000000
0!
0*
09
0>
0C
#999350000000
1!
1*
b1 6
19
1>
1C
b1 G
#999360000000
0!
0*
09
0>
0C
#999370000000
1!
1*
b10 6
19
1>
1C
b10 G
#999380000000
0!
0*
09
0>
0C
#999390000000
1!
1*
b11 6
19
1>
1C
b11 G
#999400000000
0!
0*
09
0>
0C
#999410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#999420000000
0!
0*
09
0>
0C
#999430000000
1!
1*
b101 6
19
1>
1C
b101 G
#999440000000
0!
0*
09
0>
0C
#999450000000
1!
1*
b110 6
19
1>
1C
b110 G
#999460000000
0!
0*
09
0>
0C
#999470000000
1!
1*
b111 6
19
1>
1C
b111 G
#999480000000
0!
0*
09
0>
0C
#999490000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#999500000000
0!
0*
09
0>
0C
#999510000000
1!
1*
b1 6
19
1>
1C
b1 G
#999520000000
0!
0*
09
0>
0C
#999530000000
1!
1*
b10 6
19
1>
1C
b10 G
#999540000000
0!
0*
09
0>
0C
#999550000000
1!
1*
b11 6
19
1>
1C
b11 G
#999560000000
0!
0*
09
0>
0C
#999570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#999580000000
0!
0*
09
0>
0C
#999590000000
1!
1*
b101 6
19
1>
1C
b101 G
#999600000000
0!
0*
09
0>
0C
#999610000000
1!
1*
b110 6
19
1>
1C
b110 G
#999620000000
0!
0*
09
0>
0C
#999630000000
1!
1*
b111 6
19
1>
1C
b111 G
#999640000000
0!
1"
0*
1+
09
1:
0>
0C
#999650000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#999660000000
0!
0*
09
0>
0C
#999670000000
1!
1*
b1 6
19
1>
1C
b1 G
#999680000000
0!
0*
09
0>
0C
#999690000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#999700000000
0!
0*
09
0>
0C
#999710000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#999720000000
0!
0*
09
0>
0C
#999730000000
1!
1&
b1111110 '
1*
1/
b1111110 0
03
14
b0000 5
b100 6
b0 8
19
1>
1C
1D
0E
1F
b100 G
b1111110 H
b0000 I
#999740000000
0!
0*
09
0>
0C
#999750000000
1!
0$
1%
0&
1*
0-
1.
0/
b0 6
19
1>
1C
0F
b0 G
#999760000000
0!
0#
0*
0,
09
0>
0?
0C
#999770000000
1!
1*
02
19
1>
0@
0A
0B
1C
#999780000000
0!
0*
09
0>
0C
#999790000000
1!
1*
19
1>
1C
#999800000000
0!
0*
09
0>
0C
#999810000000
1!
1*
19
1>
1C
#999820000000
0!
0*
09
0>
0C
#999830000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#999840000000
0!
0*
09
0>
0C
#999850000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#999860000000
0!
0*
09
0>
0C
#999870000000
1!
1$
0%
1*
1-
0.
b1 6
19
1>
1C
b1 G
#999880000000
0!
0*
09
0>
0C
#999890000000
1!
1*
b10 6
19
1>
1C
b10 G
#999900000000
0!
0*
09
0>
0C
#999910000000
1!
1*
b11 6
19
1>
1C
b11 G
#999920000000
0!
0*
09
0>
0C
#999930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#999940000000
0!
0*
09
0>
0C
#999950000000
1!
1*
b101 6
19
1>
1C
b101 G
#999960000000
0!
0*
09
0>
0C
#999970000000
1!
1*
b110 6
19
1>
1C
b110 G
#999980000000
0!
0*
09
0>
0C
#999990000000
1!
1*
b111 6
19
1>
1C
b111 G
#1000000000000
0!
0*
09
0>
0C
