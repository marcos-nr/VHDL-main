$date
  Sat May 04 15:23:05 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp2_3 $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 4 # dig3[3:0] $end
$var reg 4 $ dig2[3:0] $end
$var reg 4 % dig1[3:0] $end
$var reg 4 & dig0[3:0] $end
$var reg 4 ' enable_disp[3:0] $end
$var reg 7 ( segmentos[6:0] $end
$scope module uut $end
$var reg 1 ) clk $end
$var reg 1 * reset $end
$var reg 4 + dig3[3:0] $end
$var reg 4 , dig2[3:0] $end
$var reg 4 - dig1[3:0] $end
$var reg 4 . dig0[3:0] $end
$var reg 4 / enable_disp[3:0] $end
$var reg 7 0 segmentos[6:0] $end
$comment state is not handled $end
$var integer 32 1 cuenta $end
$var reg 1 2 debounced_reset $end
$var reg 1 3 enable_conta $end
$var reg 4 4 bcd[3:0] $end
$scope module a $end
$var reg 1 5 clk $end
$var reg 1 6 key $end
$var reg 1 7 debounced_key $end
$var reg 1 8 key_stable $end
$var reg 1 9 last_key $end
$upscope $end
$scope module b $end
$var reg 1 : clk $end
$var reg 1 ; reset $end
$var reg 1 < enable $end
$var reg 1 = cout $end
$var integer 32 > q $end
$upscope $end
$scope module d $end
$var reg 7 ? segmentos[6:0] $end
$var reg 4 @ bcd[3:0] $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
U"
b1000 #
b0110 $
b0100 %
b0010 &
b0001 '
b0000001 (
0)
U*
b1000 +
b0110 ,
b0100 -
b0010 .
b0001 /
b0000001 0
b0 1
U2
13
b0000 4
05
U6
U7
U8
U9
0:
U;
1<
U=
b0 >
b0000001 ?
b0000 @
#10000000
1!
1)
15
1:
0=
#20000000
0!
0)
b1 1
05
0:
b1 >
#30000000
1!
1)
15
1:
#40000000
0!
0)
b10 1
05
0:
b10 >
#50000000
1!
1)
15
1:
#60000000
0!
0)
b11 1
05
0:
b11 >
#70000000
1!
1)
15
1:
1=
#80000000
0!
0)
b100 1
05
0:
b100 >
#90000000
1!
1)
15
1:
#100000000
0!
0)
b101 1
05
0:
b101 >
#110000000
1!
1)
15
1:
#120000000
0!
0)
b110 1
05
0:
b110 >
#130000000
1!
1)
15
1:
#140000000
0!
0)
b111 1
05
0:
b111 >
#150000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
b0100 4
15
1:
0=
b1001100 ?
b0100 @
#160000000
0!
0"
0)
0*
b0 1
05
06
0:
b0 >
#170000000
1!
1)
02
15
07
08
09
1:
0;
#180000000
0!
0)
b1 1
05
0:
b1 >
#190000000
1!
1)
15
1:
#200000000
0!
0)
b10 1
05
0:
b10 >
#210000000
1!
1)
15
1:
#220000000
0!
0)
b11 1
05
0:
b11 >
#230000000
1!
1)
15
1:
1=
#240000000
0!
0)
b100 1
05
0:
b100 >
#250000000
1!
1)
15
1:
#260000000
0!
0)
b101 1
05
0:
b101 >
#270000000
1!
1)
15
1:
#280000000
0!
0)
b110 1
05
0:
b110 >
#290000000
1!
1)
15
1:
#300000000
0!
0)
b111 1
05
0:
b111 >
#310000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
b0110 4
15
1:
0=
b0100000 ?
b0110 @
#320000000
0!
0)
b0 1
05
0:
b0 >
#330000000
1!
1)
15
1:
#340000000
0!
0)
b1 1
05
0:
b1 >
#350000000
1!
1)
15
1:
#360000000
0!
0)
b10 1
05
0:
b10 >
#370000000
1!
1)
15
1:
#380000000
0!
0)
b11 1
05
0:
b11 >
#390000000
1!
1)
15
1:
1=
#400000000
0!
0)
b100 1
05
0:
b100 >
#410000000
1!
1)
15
1:
#420000000
0!
0)
b101 1
05
0:
b101 >
#430000000
1!
1)
15
1:
#440000000
0!
0)
b110 1
05
0:
b110 >
#450000000
1!
1)
15
1:
#460000000
0!
0)
b111 1
05
0:
b111 >
#470000000
1!
b1000 '
b0000000 (
1)
b1000 /
b0000000 0
b1000 4
15
1:
0=
b0000000 ?
b1000 @
#480000000
0!
0)
b0 1
05
0:
b0 >
#490000000
1!
1)
15
1:
#500000000
0!
0)
b1 1
05
0:
b1 >
#510000000
1!
1)
15
1:
#520000000
0!
0)
b10 1
05
0:
b10 >
#530000000
1!
1)
15
1:
#540000000
0!
0)
b11 1
05
0:
b11 >
#550000000
1!
1)
15
1:
1=
#560000000
0!
0)
b100 1
05
0:
b100 >
#570000000
1!
1)
15
1:
#580000000
0!
0)
b101 1
05
0:
b101 >
#590000000
1!
1)
15
1:
#600000000
0!
0)
b110 1
05
0:
b110 >
#610000000
1!
1)
15
1:
#620000000
0!
0)
b111 1
05
0:
b111 >
#630000000
1!
b0001 '
b0010010 (
1)
b0001 /
b0010010 0
b0010 4
15
1:
0=
b0010010 ?
b0010 @
#640000000
0!
0)
b0 1
05
0:
b0 >
#650000000
1!
1)
15
1:
#660000000
0!
0)
b1 1
05
0:
b1 >
#670000000
1!
1)
15
1:
#680000000
0!
0)
b10 1
05
0:
b10 >
#690000000
1!
1)
15
1:
#700000000
0!
0)
b11 1
05
0:
b11 >
#710000000
1!
1)
15
1:
1=
#720000000
0!
0)
b100 1
05
0:
b100 >
#730000000
1!
1)
15
1:
#740000000
0!
0)
b101 1
05
0:
b101 >
#750000000
1!
1)
15
1:
#760000000
0!
0)
b110 1
05
0:
b110 >
#770000000
1!
1)
15
1:
#780000000
0!
0)
b111 1
05
0:
b111 >
#790000000
1!
b0010 '
b1001100 (
1)
b0010 /
b1001100 0
b0100 4
15
1:
0=
b1001100 ?
b0100 @
#800000000
0!
0)
b0 1
05
0:
b0 >
#810000000
1!
1)
15
1:
#820000000
0!
0)
b1 1
05
0:
b1 >
#830000000
1!
1)
15
1:
#840000000
0!
0)
b10 1
05
0:
b10 >
#850000000
1!
1)
15
1:
#860000000
0!
0)
b11 1
05
0:
b11 >
#870000000
1!
1)
15
1:
1=
#880000000
0!
0)
b100 1
05
0:
b100 >
#890000000
1!
1)
15
1:
#900000000
0!
0)
b101 1
05
0:
b101 >
#910000000
1!
1)
15
1:
#920000000
0!
0)
b110 1
05
0:
b110 >
#930000000
1!
1)
15
1:
#940000000
0!
0)
b111 1
05
0:
b111 >
#950000000
1!
b0100 '
b0100000 (
1)
b0100 /
b0100000 0
b0110 4
15
1:
0=
b0100000 ?
b0110 @
#960000000
0!
0)
b0 1
05
0:
b0 >
#970000000
1!
1)
15
1:
#980000000
0!
0)
b1 1
05
0:
b1 >
#990000000
1!
1)
15
1:
#1000000000
0!
0)
b10 1
05
0:
b10 >
