$date
  Mon May 06 00:38:05 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp3_2 $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 1 # up $end
$var reg 1 $ down $end
$var reg 4 % enable_disp[3:0] $end
$var reg 7 & segmentos[6:0] $end
$scope module uut $end
$var reg 1 ' clk $end
$var reg 1 ( reset $end
$var reg 1 ) up $end
$var reg 1 * down $end
$var reg 4 + enable_disp[3:0] $end
$var reg 7 , segmentos[6:0] $end
$var reg 1 - debounced_reset $end
$var reg 1 . debounced_up $end
$var reg 1 / debounced_down $end
$var reg 4 0 dig3[3:0] $end
$var reg 4 1 dig2[3:0] $end
$var reg 4 2 dig1[3:0] $end
$var reg 4 3 dig0[3:0] $end
$scope module a $end
$var reg 1 4 clk $end
$var reg 1 5 key $end
$var reg 1 6 debounced_key $end
$var reg 1 7 key_stable $end
$var reg 1 8 last_key $end
$upscope $end
$scope module b $end
$var reg 1 9 clk $end
$var reg 1 : key $end
$var reg 1 ; debounced_key $end
$var reg 1 < key_stable $end
$var reg 1 = last_key $end
$upscope $end
$scope module c $end
$var reg 1 > clk $end
$var reg 1 ? key $end
$var reg 1 @ debounced_key $end
$var reg 1 A key_stable $end
$var reg 1 B last_key $end
$upscope $end
$scope module d $end
$var reg 1 C clk $end
$var reg 1 D reset $end
$var reg 4 E dig3[3:0] $end
$var reg 4 F dig2[3:0] $end
$var reg 4 G dig1[3:0] $end
$var reg 4 H dig0[3:0] $end
$var reg 4 I enable_disp[3:0] $end
$var reg 7 J segmentos[6:0] $end
$comment state is not handled $end
$var integer 32 K cuenta $end
$var reg 1 L debounced_reset $end
$var reg 1 M clock_reset $end
$var reg 1 N enable_conta $end
$var reg 4 O bcd[3:0] $end
$scope module a $end
$var reg 1 P clk $end
$var reg 1 Q key $end
$var reg 1 R debounced_key $end
$var reg 1 S key_stable $end
$var reg 1 T last_key $end
$upscope $end
$scope module b $end
$var reg 1 U clk $end
$var reg 1 V reset $end
$var reg 1 W enable $end
$var reg 1 X cout $end
$var integer 32 Y q $end
$upscope $end
$scope module d $end
$var reg 7 Z segmentos[6:0] $end
$var reg 4 [ bcd[3:0] $end
$upscope $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
1"
1#
1$
b0001 %
b1000111 &
0'
1(
1)
1*
b0001 +
b1000111 ,
U-
U.
U/
b0000 0
b0000 1
b0000 2
b0000 3
04
15
U6
U7
U8
09
1:
U;
U<
U=
0>
1?
U@
UA
UB
0C
UD
b0000 E
b0000 F
b0000 G
b0000 H
b0001 I
b1000111 J
b0 K
UL
UM
1N
bUUUU O
0P
UQ
UR
US
UT
0U
UV
1W
UX
b0 Y
b1000111 Z
bUUUU [
#10000000
1!
1'
1-
1.
1/
14
16
17
18
19
1;
1<
1=
1>
1@
1A
1B
1C
1D
1P
1Q
1U
0X
#20000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#30000000
1!
1'
14
19
1>
1C
1L
0M
1P
1R
1S
1T
1U
0V
#40000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#50000000
1!
1'
14
19
1>
1C
1P
1U
1X
#60000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#70000000
1!
1'
14
19
1>
1C
1P
1U
#80000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#90000000
1!
1'
14
19
1>
1C
1P
1U
#100000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#110000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#120000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#130000000
1!
1'
14
19
1>
1C
1P
1U
#140000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#150000000
1!
1'
14
19
1>
1C
1P
1U
#160000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#170000000
1!
1'
14
19
1>
1C
1P
1U
1X
#180000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#190000000
1!
1'
14
19
1>
1C
1P
1U
#200000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#210000000
1!
1'
14
19
1>
1C
1P
1U
#220000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#230000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#240000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#250000000
1!
1'
14
19
1>
1C
1P
1U
#260000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#270000000
1!
1'
14
19
1>
1C
1P
1U
#280000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#290000000
1!
1'
14
19
1>
1C
1P
1U
1X
#300000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#310000000
1!
1'
14
19
1>
1C
1P
1U
#320000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#330000000
1!
1'
14
19
1>
1C
1P
1U
#340000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#350000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#360000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#370000000
1!
1'
14
19
1>
1C
1P
1U
#380000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#390000000
1!
1'
14
19
1>
1C
1P
1U
#400000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#410000000
1!
1'
14
19
1>
1C
1P
1U
1X
#420000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#430000000
1!
1'
14
19
1>
1C
1P
1U
#440000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#450000000
1!
1'
14
19
1>
1C
1P
1U
#460000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#470000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#480000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#490000000
1!
1'
14
19
1>
1C
1P
1U
#500000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#510000000
1!
1'
14
19
1>
1C
1P
1U
#520000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#530000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
1X
#540000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#550000000
1!
1'
b0001 3
14
19
1>
1C
b0001 H
1P
1U
#560000000
0!
1#
0'
1)
04
09
1:
0>
0C
b100 K
0P
0U
b100 Y
#570000000
#580000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#590000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#600000000
1!
b0010 %
1'
b0010 +
14
19
1>
1C
b0010 I
1P
1U
0X
#610000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#620000000
1!
1'
14
19
1>
1C
1P
1U
#630000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#640000000
1!
1'
14
19
1>
1C
1P
1U
#650000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#660000000
1!
1'
14
19
1>
1C
1P
1U
1X
#670000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#680000000
1!
1'
14
19
1>
1C
1P
1U
#690000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#700000000
1!
1'
14
19
1>
1C
1P
1U
#710000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#720000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#730000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#740000000
1!
1'
14
19
1>
1C
1P
1U
#750000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#760000000
1!
1'
14
19
1>
1C
1P
1U
#770000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#780000000
1!
1'
14
19
1>
1C
1P
1U
1X
#790000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#800000000
1!
1'
14
19
1>
1C
1P
1U
#810000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#820000000
1!
1'
14
19
1>
1C
1P
1U
#830000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#840000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#850000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#860000000
1!
1'
14
19
1>
1C
1P
1U
#870000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#880000000
1!
1'
14
19
1>
1C
1P
1U
#890000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#900000000
1!
1'
14
19
1>
1C
1P
1U
1X
#910000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#920000000
1!
1'
14
19
1>
1C
1P
1U
#930000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#940000000
1!
1'
14
19
1>
1C
1P
1U
#950000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#960000000
1!
b0001 %
b0110000 &
1'
b0001 +
b0110000 ,
14
19
1>
1C
b0001 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#970000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#980000000
1!
1'
14
19
1>
1C
1P
1U
#990000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#1000000000
1!
1'
14
19
1>
1C
1P
1U
#1010000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#1020000000
1!
1'
14
19
1>
1C
1P
1U
1X
#1030000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#1040000000
1!
1'
14
19
1>
1C
1P
1U
#1050000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#1060000000
1!
1'
14
19
1>
1C
1P
1U
#1070000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#1080000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#1090000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#1100000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#1110000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#1120000000
1!
1'
b0010 3
14
19
1>
1C
b0010 H
1P
1U
#1130000000
0!
1#
0'
1)
04
09
1:
0>
0C
b10 K
0P
0U
b10 Y
#1140000000
#1150000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
1X
#1160000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#1170000000
1!
1'
14
19
1>
1C
1P
1U
#1180000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#1190000000
1!
1'
14
19
1>
1C
1P
1U
#1200000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#1210000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#1220000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#1230000000
1!
1'
14
19
1>
1C
1P
1U
#1240000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#1250000000
1!
1'
14
19
1>
1C
1P
1U
#1260000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#1270000000
1!
1'
14
19
1>
1C
1P
1U
1X
#1280000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#1290000000
1!
1'
14
19
1>
1C
1P
1U
#1300000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#1310000000
1!
1'
14
19
1>
1C
1P
1U
#1320000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#1330000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#1340000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#1350000000
1!
1'
14
19
1>
1C
1P
1U
#1360000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#1370000000
1!
1'
14
19
1>
1C
1P
1U
#1380000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#1390000000
1!
1'
14
19
1>
1C
1P
1U
1X
#1400000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#1410000000
1!
1'
14
19
1>
1C
1P
1U
#1420000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#1430000000
1!
1'
14
19
1>
1C
1P
1U
#1440000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#1450000000
1!
b0001 %
b1101101 &
1'
b0001 +
b1101101 ,
14
19
1>
1C
b0001 I
b1101101 J
b0010 O
1P
1U
0X
b1101101 Z
b0010 [
#1460000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#1470000000
1!
1'
14
19
1>
1C
1P
1U
#1480000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#1490000000
1!
1'
14
19
1>
1C
1P
1U
#1500000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#1510000000
1!
1'
14
19
1>
1C
1P
1U
1X
#1520000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#1530000000
1!
1'
14
19
1>
1C
1P
1U
#1540000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#1550000000
1!
1'
14
19
1>
1C
1P
1U
#1560000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#1570000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#1580000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#1590000000
1!
1'
14
19
1>
1C
1P
1U
#1600000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#1610000000
1!
1'
14
19
1>
1C
1P
1U
#1620000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#1630000000
1!
1'
14
19
1>
1C
1P
1U
1X
#1640000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#1650000000
1!
1'
14
19
1>
1C
1P
1U
#1660000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#1670000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#1680000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#1690000000
1!
b0100 %
1'
b0100 +
b0011 3
14
19
1>
1C
b0011 H
b0100 I
1P
1U
0X
#1700000000
0!
1#
0'
1)
04
09
1:
0>
0C
b0 K
0P
0U
b0 Y
#1710000000
#1720000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#1730000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#1740000000
1!
1'
14
19
1>
1C
1P
1U
#1750000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#1760000000
1!
1'
14
19
1>
1C
1P
1U
1X
#1770000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#1780000000
1!
1'
14
19
1>
1C
1P
1U
#1790000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#1800000000
1!
1'
14
19
1>
1C
1P
1U
#1810000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#1820000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#1830000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#1840000000
1!
1'
14
19
1>
1C
1P
1U
#1850000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#1860000000
1!
1'
14
19
1>
1C
1P
1U
#1870000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#1880000000
1!
1'
14
19
1>
1C
1P
1U
1X
#1890000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#1900000000
1!
1'
14
19
1>
1C
1P
1U
#1910000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#1920000000
1!
1'
14
19
1>
1C
1P
1U
#1930000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#1940000000
1!
b0001 %
b1111001 &
1'
b0001 +
b1111001 ,
14
19
1>
1C
b0001 I
b1111001 J
b0011 O
1P
1U
0X
b1111001 Z
b0011 [
#1950000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#1960000000
1!
1'
14
19
1>
1C
1P
1U
#1970000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#1980000000
1!
1'
14
19
1>
1C
1P
1U
#1990000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#2000000000
1!
1'
14
19
1>
1C
1P
1U
1X
#2010000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#2020000000
1!
1'
14
19
1>
1C
1P
1U
#2030000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#2040000000
1!
1'
14
19
1>
1C
1P
1U
#2050000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#2060000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#2070000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#2080000000
1!
1'
14
19
1>
1C
1P
1U
#2090000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#2100000000
1!
1'
14
19
1>
1C
1P
1U
#2110000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#2120000000
1!
1'
14
19
1>
1C
1P
1U
1X
#2130000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#2140000000
1!
1'
14
19
1>
1C
1P
1U
#2150000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#2160000000
1!
1'
14
19
1>
1C
1P
1U
#2170000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#2180000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#2190000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#2200000000
1!
1'
14
19
1>
1C
1P
1U
#2210000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#2220000000
1!
1'
14
19
1>
1C
1P
1U
#2230000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#2240000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
1X
#2250000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#2260000000
1!
1'
b0100 3
14
19
1>
1C
b0100 H
1P
1U
#2270000000
0!
1#
0'
1)
04
09
1:
0>
0C
b100 K
0P
0U
b100 Y
#2280000000
#2290000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#2300000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#2310000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#2320000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#2330000000
1!
1'
14
19
1>
1C
1P
1U
#2340000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#2350000000
1!
1'
14
19
1>
1C
1P
1U
#2360000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#2370000000
1!
1'
14
19
1>
1C
1P
1U
1X
#2380000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#2390000000
1!
1'
14
19
1>
1C
1P
1U
#2400000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#2410000000
1!
1'
14
19
1>
1C
1P
1U
#2420000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#2430000000
1!
b0001 %
b0110011 &
1'
b0001 +
b0110011 ,
14
19
1>
1C
b0001 I
b0110011 J
b0100 O
1P
1U
0X
b0110011 Z
b0100 [
#2440000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#2450000000
1!
1'
14
19
1>
1C
1P
1U
#2460000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#2470000000
1!
1'
14
19
1>
1C
1P
1U
#2480000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#2490000000
1!
1'
14
19
1>
1C
1P
1U
1X
#2500000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#2510000000
1!
1'
14
19
1>
1C
1P
1U
#2520000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#2530000000
1!
1'
14
19
1>
1C
1P
1U
#2540000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#2550000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#2560000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#2570000000
1!
1'
14
19
1>
1C
1P
1U
#2580000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#2590000000
1!
1'
14
19
1>
1C
1P
1U
#2600000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#2610000000
1!
1'
14
19
1>
1C
1P
1U
1X
#2620000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#2630000000
1!
1'
14
19
1>
1C
1P
1U
#2640000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#2650000000
1!
1'
14
19
1>
1C
1P
1U
#2660000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#2670000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#2680000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#2690000000
1!
1'
14
19
1>
1C
1P
1U
#2700000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#2710000000
1!
1'
14
19
1>
1C
1P
1U
#2720000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#2730000000
1!
1'
14
19
1>
1C
1P
1U
1X
#2740000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#2750000000
1!
1'
14
19
1>
1C
1P
1U
#2760000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#2770000000
1!
1'
14
19
1>
1C
1P
1U
#2780000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#2790000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#2800000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#2810000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#2820000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#2830000000
1!
1'
b0101 3
14
19
1>
1C
b0101 H
1P
1U
#2840000000
0!
1#
0'
1)
04
09
1:
0>
0C
b10 K
0P
0U
b10 Y
#2850000000
#2860000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
1X
#2870000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#2880000000
1!
1'
14
19
1>
1C
1P
1U
#2890000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#2900000000
1!
1'
14
19
1>
1C
1P
1U
#2910000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#2920000000
1!
b0001 %
b1011011 &
1'
b0001 +
b1011011 ,
14
19
1>
1C
b0001 I
b1011011 J
b0101 O
1P
1U
0X
b1011011 Z
b0101 [
#2930000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#2940000000
1!
1'
14
19
1>
1C
1P
1U
#2950000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#2960000000
1!
1'
14
19
1>
1C
1P
1U
#2970000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#2980000000
1!
1'
14
19
1>
1C
1P
1U
1X
#2990000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#3000000000
1!
1'
14
19
1>
1C
1P
1U
#3010000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#3020000000
1!
1'
14
19
1>
1C
1P
1U
#3030000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#3040000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#3050000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#3060000000
1!
1'
14
19
1>
1C
1P
1U
#3070000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#3080000000
1!
1'
14
19
1>
1C
1P
1U
#3090000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#3100000000
1!
1'
14
19
1>
1C
1P
1U
1X
#3110000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#3120000000
1!
1'
14
19
1>
1C
1P
1U
#3130000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#3140000000
1!
1'
14
19
1>
1C
1P
1U
#3150000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#3160000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#3170000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#3180000000
1!
1'
14
19
1>
1C
1P
1U
#3190000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#3200000000
1!
1'
14
19
1>
1C
1P
1U
#3210000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#3220000000
1!
1'
14
19
1>
1C
1P
1U
1X
#3230000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#3240000000
1!
1'
14
19
1>
1C
1P
1U
#3250000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#3260000000
1!
1'
14
19
1>
1C
1P
1U
#3270000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#3280000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#3290000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#3300000000
1!
1'
14
19
1>
1C
1P
1U
#3310000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#3320000000
1!
1'
14
19
1>
1C
1P
1U
#3330000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#3340000000
1!
1'
14
19
1>
1C
1P
1U
1X
#3350000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#3360000000
1!
1'
14
19
1>
1C
1P
1U
#3370000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#3380000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#3390000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#3400000000
1!
b0001 %
b1011111 &
1'
b0001 +
b1011111 ,
b0110 3
14
19
1>
1C
b0110 H
b0001 I
b1011111 J
b0110 O
1P
1U
0X
b1011111 Z
b0110 [
#3410000000
0!
1#
0'
1)
04
09
1:
0>
0C
b0 K
0P
0U
b0 Y
#3420000000
#3430000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#3440000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#3450000000
1!
1'
14
19
1>
1C
1P
1U
#3460000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#3470000000
1!
1'
14
19
1>
1C
1P
1U
1X
#3480000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#3490000000
1!
1'
14
19
1>
1C
1P
1U
#3500000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#3510000000
1!
1'
14
19
1>
1C
1P
1U
#3520000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#3530000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#3540000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#3550000000
1!
1'
14
19
1>
1C
1P
1U
#3560000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#3570000000
1!
1'
14
19
1>
1C
1P
1U
#3580000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#3590000000
1!
1'
14
19
1>
1C
1P
1U
1X
#3600000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#3610000000
1!
1'
14
19
1>
1C
1P
1U
#3620000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#3630000000
1!
1'
14
19
1>
1C
1P
1U
#3640000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#3650000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#3660000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#3670000000
1!
1'
14
19
1>
1C
1P
1U
#3680000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#3690000000
1!
1'
14
19
1>
1C
1P
1U
#3700000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#3710000000
1!
1'
14
19
1>
1C
1P
1U
1X
#3720000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#3730000000
1!
1'
14
19
1>
1C
1P
1U
#3740000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#3750000000
1!
1'
14
19
1>
1C
1P
1U
#3760000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#3770000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#3780000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#3790000000
1!
1'
14
19
1>
1C
1P
1U
#3800000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#3810000000
1!
1'
14
19
1>
1C
1P
1U
#3820000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#3830000000
1!
1'
14
19
1>
1C
1P
1U
1X
#3840000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#3850000000
1!
1'
14
19
1>
1C
1P
1U
#3860000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#3870000000
1!
1'
14
19
1>
1C
1P
1U
#3880000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#3890000000
1!
b0001 %
b1011111 &
1'
b0001 +
b1011111 ,
14
19
1>
1C
b0001 I
b1011111 J
b0110 O
1P
1U
0X
b1011111 Z
b0110 [
#3900000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#3910000000
1!
1'
14
19
1>
1C
1P
1U
#3920000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#3930000000
1!
1'
14
19
1>
1C
1P
1U
#3940000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#3950000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
1X
#3960000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#3970000000
1!
1'
b0111 3
14
19
1>
1C
b0111 H
1P
1U
#3980000000
0!
1#
0'
1)
04
09
1:
0>
0C
b100 K
0P
0U
b100 Y
#3990000000
#4000000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#4010000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#4020000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#4030000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#4040000000
1!
1'
14
19
1>
1C
1P
1U
#4050000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#4060000000
1!
1'
14
19
1>
1C
1P
1U
#4070000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#4080000000
1!
1'
14
19
1>
1C
1P
1U
1X
#4090000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#4100000000
1!
1'
14
19
1>
1C
1P
1U
#4110000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#4120000000
1!
1'
14
19
1>
1C
1P
1U
#4130000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#4140000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#4150000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#4160000000
1!
1'
14
19
1>
1C
1P
1U
#4170000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#4180000000
1!
1'
14
19
1>
1C
1P
1U
#4190000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#4200000000
1!
1'
14
19
1>
1C
1P
1U
1X
#4210000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#4220000000
1!
1'
14
19
1>
1C
1P
1U
#4230000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#4240000000
1!
1'
14
19
1>
1C
1P
1U
#4250000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#4260000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#4270000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#4280000000
1!
1'
14
19
1>
1C
1P
1U
#4290000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#4300000000
1!
1'
14
19
1>
1C
1P
1U
#4310000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#4320000000
1!
1'
14
19
1>
1C
1P
1U
1X
#4330000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#4340000000
1!
1'
14
19
1>
1C
1P
1U
#4350000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#4360000000
1!
1'
14
19
1>
1C
1P
1U
#4370000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#4380000000
1!
b0001 %
b1110000 &
1'
b0001 +
b1110000 ,
14
19
1>
1C
b0001 I
b1110000 J
b0111 O
1P
1U
0X
b1110000 Z
b0111 [
#4390000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#4400000000
1!
1'
14
19
1>
1C
1P
1U
#4410000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#4420000000
1!
1'
14
19
1>
1C
1P
1U
#4430000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#4440000000
1!
1'
14
19
1>
1C
1P
1U
1X
#4450000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#4460000000
1!
1'
14
19
1>
1C
1P
1U
#4470000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#4480000000
1!
1'
14
19
1>
1C
1P
1U
#4490000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#4500000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#4510000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#4520000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#4530000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#4540000000
1!
1'
b1000 3
14
19
1>
1C
b1000 H
1P
1U
#4550000000
0!
1#
0'
1)
04
09
1:
0>
0C
b10 K
0P
0U
b10 Y
#4560000000
#4570000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
1X
#4580000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#4590000000
1!
1'
14
19
1>
1C
1P
1U
#4600000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#4610000000
1!
1'
14
19
1>
1C
1P
1U
#4620000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#4630000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#4640000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#4650000000
1!
1'
14
19
1>
1C
1P
1U
#4660000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#4670000000
1!
1'
14
19
1>
1C
1P
1U
#4680000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#4690000000
1!
1'
14
19
1>
1C
1P
1U
1X
#4700000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#4710000000
1!
1'
14
19
1>
1C
1P
1U
#4720000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#4730000000
1!
1'
14
19
1>
1C
1P
1U
#4740000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#4750000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#4760000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#4770000000
1!
1'
14
19
1>
1C
1P
1U
#4780000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#4790000000
1!
1'
14
19
1>
1C
1P
1U
#4800000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#4810000000
1!
1'
14
19
1>
1C
1P
1U
1X
#4820000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#4830000000
1!
1'
14
19
1>
1C
1P
1U
#4840000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#4850000000
1!
1'
14
19
1>
1C
1P
1U
#4860000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#4870000000
1!
b0001 %
b1111111 &
1'
b0001 +
b1111111 ,
14
19
1>
1C
b0001 I
b1111111 J
b1000 O
1P
1U
0X
b1111111 Z
b1000 [
#4880000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#4890000000
1!
1'
14
19
1>
1C
1P
1U
#4900000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#4910000000
1!
1'
14
19
1>
1C
1P
1U
#4920000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#4930000000
1!
1'
14
19
1>
1C
1P
1U
1X
#4940000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#4950000000
1!
1'
14
19
1>
1C
1P
1U
#4960000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#4970000000
1!
1'
14
19
1>
1C
1P
1U
#4980000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#4990000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#5000000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#5010000000
1!
1'
14
19
1>
1C
1P
1U
#5020000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#5030000000
1!
1'
14
19
1>
1C
1P
1U
#5040000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#5050000000
1!
1'
14
19
1>
1C
1P
1U
1X
#5060000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#5070000000
1!
1'
14
19
1>
1C
1P
1U
#5080000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#5090000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#5100000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#5110000000
1!
b0100 %
1'
b0100 +
b1001 3
14
19
1>
1C
b1001 H
b0100 I
1P
1U
0X
#5120000000
0!
1#
0'
1)
04
09
1:
0>
0C
b0 K
0P
0U
b0 Y
#5130000000
#5140000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#5150000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#5160000000
1!
1'
14
19
1>
1C
1P
1U
#5170000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#5180000000
1!
1'
14
19
1>
1C
1P
1U
1X
#5190000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#5200000000
1!
1'
14
19
1>
1C
1P
1U
#5210000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#5220000000
1!
1'
14
19
1>
1C
1P
1U
#5230000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#5240000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#5250000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#5260000000
1!
1'
14
19
1>
1C
1P
1U
#5270000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#5280000000
1!
1'
14
19
1>
1C
1P
1U
#5290000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#5300000000
1!
1'
14
19
1>
1C
1P
1U
1X
#5310000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#5320000000
1!
1'
14
19
1>
1C
1P
1U
#5330000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#5340000000
1!
1'
14
19
1>
1C
1P
1U
#5350000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#5360000000
1!
b0001 %
b1111011 &
1'
b0001 +
b1111011 ,
14
19
1>
1C
b0001 I
b1111011 J
b1001 O
1P
1U
0X
b1111011 Z
b1001 [
#5370000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#5380000000
1!
1'
14
19
1>
1C
1P
1U
#5390000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#5400000000
1!
1'
14
19
1>
1C
1P
1U
#5410000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#5420000000
1!
1'
14
19
1>
1C
1P
1U
1X
#5430000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#5440000000
1!
1'
14
19
1>
1C
1P
1U
#5450000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#5460000000
1!
1'
14
19
1>
1C
1P
1U
#5470000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#5480000000
1!
b0010 %
b1111110 &
1'
b0010 +
b1111110 ,
14
19
1>
1C
b0010 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#5490000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#5500000000
1!
1'
14
19
1>
1C
1P
1U
#5510000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#5520000000
1!
1'
14
19
1>
1C
1P
1U
#5530000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#5540000000
1!
1'
14
19
1>
1C
1P
1U
1X
#5550000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#5560000000
1!
1'
14
19
1>
1C
1P
1U
#5570000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#5580000000
1!
1'
14
19
1>
1C
1P
1U
#5590000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#5600000000
1!
b0100 %
1'
b0100 +
14
19
1>
1C
b0100 I
1P
1U
0X
#5610000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#5620000000
1!
1'
14
19
1>
1C
1P
1U
#5630000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#5640000000
1!
1'
14
19
1>
1C
1P
1U
#5650000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#5660000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
1X
#5670000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#5680000000
1!
1'
b0001 2
b0000 3
14
19
1>
1C
b0001 G
b0000 H
1P
1U
#5690000000
0!
1#
0'
1)
04
09
1:
0>
0C
b100 K
0P
0U
b100 Y
#5700000000
#5710000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#5720000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#5730000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#5740000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#5750000000
1!
1'
14
19
1>
1C
1P
1U
#5760000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#5770000000
1!
1'
14
19
1>
1C
1P
1U
#5780000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#5790000000
1!
1'
14
19
1>
1C
1P
1U
1X
#5800000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#5810000000
1!
1'
14
19
1>
1C
1P
1U
#5820000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#5830000000
1!
1'
14
19
1>
1C
1P
1U
#5840000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#5850000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#5860000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#5870000000
1!
1'
14
19
1>
1C
1P
1U
#5880000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#5890000000
1!
1'
14
19
1>
1C
1P
1U
#5900000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#5910000000
1!
1'
14
19
1>
1C
1P
1U
1X
#5920000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#5930000000
1!
1'
14
19
1>
1C
1P
1U
#5940000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#5950000000
1!
1'
14
19
1>
1C
1P
1U
#5960000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#5970000000
1!
b0010 %
b0110000 &
1'
b0010 +
b0110000 ,
14
19
1>
1C
b0010 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#5980000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#5990000000
1!
1'
14
19
1>
1C
1P
1U
#6000000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#6010000000
1!
1'
14
19
1>
1C
1P
1U
#6020000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#6030000000
1!
1'
14
19
1>
1C
1P
1U
1X
#6040000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#6050000000
1!
1'
14
19
1>
1C
1P
1U
#6060000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#6070000000
1!
1'
14
19
1>
1C
1P
1U
#6080000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#6090000000
1!
b0100 %
b1111110 &
1'
b0100 +
b1111110 ,
14
19
1>
1C
b0100 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#6100000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#6110000000
1!
1'
14
19
1>
1C
1P
1U
#6120000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#6130000000
1!
1'
14
19
1>
1C
1P
1U
#6140000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#6150000000
1!
1'
14
19
1>
1C
1P
1U
1X
#6160000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#6170000000
1!
1'
14
19
1>
1C
1P
1U
#6180000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#6190000000
1!
1'
14
19
1>
1C
1P
1U
#6200000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#6210000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#6220000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#6230000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#6240000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#6250000000
1!
1'
14
19
1>
1C
1P
1U
#6260000000
0!
1#
0'
1)
04
09
1:
0>
0C
b10 K
0P
0U
b10 Y
#6270000000
#6280000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
1X
#6290000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#6300000000
1!
1'
14
19
1>
1C
1P
1U
#6310000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#6320000000
1!
1'
14
19
1>
1C
1P
1U
#6330000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#6340000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#6350000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#6360000000
1!
1'
14
19
1>
1C
1P
1U
#6370000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#6380000000
1!
1'
14
19
1>
1C
1P
1U
#6390000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#6400000000
1!
1'
14
19
1>
1C
1P
1U
1X
#6410000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#6420000000
1!
1'
14
19
1>
1C
1P
1U
#6430000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#6440000000
1!
1'
14
19
1>
1C
1P
1U
#6450000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#6460000000
1!
b0010 %
b0110000 &
1'
b0010 +
b0110000 ,
14
19
1>
1C
b0010 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#6470000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#6480000000
1!
1'
14
19
1>
1C
1P
1U
#6490000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#6500000000
1!
1'
14
19
1>
1C
1P
1U
#6510000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#6520000000
1!
1'
14
19
1>
1C
1P
1U
1X
#6530000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#6540000000
1!
1'
14
19
1>
1C
1P
1U
#6550000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#6560000000
1!
1'
14
19
1>
1C
1P
1U
#6570000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#6580000000
1!
b0100 %
b1111110 &
1'
b0100 +
b1111110 ,
14
19
1>
1C
b0100 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#6590000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#6600000000
1!
1'
14
19
1>
1C
1P
1U
#6610000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#6620000000
1!
1'
14
19
1>
1C
1P
1U
#6630000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#6640000000
1!
1'
14
19
1>
1C
1P
1U
1X
#6650000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#6660000000
1!
1'
14
19
1>
1C
1P
1U
#6670000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#6680000000
1!
1'
14
19
1>
1C
1P
1U
#6690000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#6700000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#6710000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#6720000000
1!
1'
14
19
1>
1C
1P
1U
#6730000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#6740000000
1!
1'
14
19
1>
1C
1P
1U
#6750000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#6760000000
1!
1'
14
19
1>
1C
1P
1U
1X
#6770000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#6780000000
1!
1'
14
19
1>
1C
1P
1U
#6790000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#6800000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#6810000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#6820000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#6830000000
0!
1#
0'
1)
04
09
1:
0>
0C
b0 K
0P
0U
b0 Y
#6840000000
#6850000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#6860000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#6870000000
1!
1'
14
19
1>
1C
1P
1U
#6880000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#6890000000
1!
1'
14
19
1>
1C
1P
1U
1X
#6900000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#6910000000
1!
1'
14
19
1>
1C
1P
1U
#6920000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#6930000000
1!
1'
14
19
1>
1C
1P
1U
#6940000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#6950000000
1!
b0010 %
b0110000 &
1'
b0010 +
b0110000 ,
14
19
1>
1C
b0010 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#6960000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#6970000000
1!
1'
14
19
1>
1C
1P
1U
#6980000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#6990000000
1!
1'
14
19
1>
1C
1P
1U
#7000000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#7010000000
1!
1'
14
19
1>
1C
1P
1U
1X
#7020000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#7030000000
1!
1'
14
19
1>
1C
1P
1U
#7040000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#7050000000
1!
1'
14
19
1>
1C
1P
1U
#7060000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#7070000000
1!
b0100 %
b1111110 &
1'
b0100 +
b1111110 ,
14
19
1>
1C
b0100 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#7080000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#7090000000
1!
1'
14
19
1>
1C
1P
1U
#7100000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#7110000000
1!
1'
14
19
1>
1C
1P
1U
#7120000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#7130000000
1!
1'
14
19
1>
1C
1P
1U
1X
#7140000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#7150000000
1!
1'
14
19
1>
1C
1P
1U
#7160000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#7170000000
1!
1'
14
19
1>
1C
1P
1U
#7180000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#7190000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#7200000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#7210000000
1!
1'
14
19
1>
1C
1P
1U
#7220000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#7230000000
1!
1'
14
19
1>
1C
1P
1U
#7240000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#7250000000
1!
1'
14
19
1>
1C
1P
1U
1X
#7260000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#7270000000
1!
1'
14
19
1>
1C
1P
1U
#7280000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#7290000000
1!
1'
14
19
1>
1C
1P
1U
#7300000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#7310000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#7320000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#7330000000
1!
1'
14
19
1>
1C
1P
1U
#7340000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#7350000000
1!
1'
14
19
1>
1C
1P
1U
#7360000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#7370000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
1X
#7380000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#7390000000
1!
1'
14
19
1>
1C
1P
1U
#7400000000
0!
1#
0'
1)
04
09
1:
0>
0C
b100 K
0P
0U
b100 Y
#7410000000
#7420000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#7430000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#7440000000
1!
b0010 %
b0110000 &
1'
b0010 +
b0110000 ,
14
19
1>
1C
b0010 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#7450000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#7460000000
1!
1'
14
19
1>
1C
1P
1U
#7470000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#7480000000
1!
1'
14
19
1>
1C
1P
1U
#7490000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#7500000000
1!
1'
14
19
1>
1C
1P
1U
1X
#7510000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#7520000000
1!
1'
14
19
1>
1C
1P
1U
#7530000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#7540000000
1!
1'
14
19
1>
1C
1P
1U
#7550000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#7560000000
1!
b0100 %
b1111110 &
1'
b0100 +
b1111110 ,
14
19
1>
1C
b0100 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#7570000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#7580000000
1!
1'
14
19
1>
1C
1P
1U
#7590000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#7600000000
1!
1'
14
19
1>
1C
1P
1U
#7610000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#7620000000
1!
1'
14
19
1>
1C
1P
1U
1X
#7630000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#7640000000
1!
1'
14
19
1>
1C
1P
1U
#7650000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#7660000000
1!
1'
14
19
1>
1C
1P
1U
#7670000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#7680000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#7690000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#7700000000
1!
1'
14
19
1>
1C
1P
1U
#7710000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#7720000000
1!
1'
14
19
1>
1C
1P
1U
#7730000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#7740000000
1!
1'
14
19
1>
1C
1P
1U
1X
#7750000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#7760000000
1!
1'
14
19
1>
1C
1P
1U
#7770000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#7780000000
1!
1'
14
19
1>
1C
1P
1U
#7790000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#7800000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#7810000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#7820000000
1!
1'
14
19
1>
1C
1P
1U
#7830000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#7840000000
1!
1'
14
19
1>
1C
1P
1U
#7850000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#7860000000
1!
1'
14
19
1>
1C
1P
1U
1X
#7870000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#7880000000
1!
1'
14
19
1>
1C
1P
1U
#7890000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#7900000000
1!
1'
14
19
1>
1C
1P
1U
#7910000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#7920000000
1!
b0010 %
b0110000 &
1'
b0010 +
b0110000 ,
14
19
1>
1C
b0010 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#7930000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#7940000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#7950000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#7960000000
1!
1'
14
19
1>
1C
1P
1U
#7970000000
0!
1#
0'
1)
04
09
1:
0>
0C
b10 K
0P
0U
b10 Y
#7980000000
#7990000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
1X
#8000000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#8010000000
1!
1'
14
19
1>
1C
1P
1U
#8020000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#8030000000
1!
1'
14
19
1>
1C
1P
1U
#8040000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#8050000000
1!
b0100 %
b1111110 &
1'
b0100 +
b1111110 ,
14
19
1>
1C
b0100 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#8060000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#8070000000
1!
1'
14
19
1>
1C
1P
1U
#8080000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#8090000000
1!
1'
14
19
1>
1C
1P
1U
#8100000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#8110000000
1!
1'
14
19
1>
1C
1P
1U
1X
#8120000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#8130000000
1!
1'
14
19
1>
1C
1P
1U
#8140000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#8150000000
1!
1'
14
19
1>
1C
1P
1U
#8160000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#8170000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#8180000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#8190000000
1!
1'
14
19
1>
1C
1P
1U
#8200000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#8210000000
1!
1'
14
19
1>
1C
1P
1U
#8220000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#8230000000
1!
1'
14
19
1>
1C
1P
1U
1X
#8240000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#8250000000
1!
1'
14
19
1>
1C
1P
1U
#8260000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#8270000000
1!
1'
14
19
1>
1C
1P
1U
#8280000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#8290000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#8300000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#8310000000
1!
1'
14
19
1>
1C
1P
1U
#8320000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#8330000000
1!
1'
14
19
1>
1C
1P
1U
#8340000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#8350000000
1!
1'
14
19
1>
1C
1P
1U
1X
#8360000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#8370000000
1!
1'
14
19
1>
1C
1P
1U
#8380000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#8390000000
1!
1'
14
19
1>
1C
1P
1U
#8400000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#8410000000
1!
b0010 %
b0110000 &
1'
b0010 +
b0110000 ,
14
19
1>
1C
b0010 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#8420000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#8430000000
1!
1'
14
19
1>
1C
1P
1U
#8440000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#8450000000
1!
1'
14
19
1>
1C
1P
1U
#8460000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#8470000000
1!
1'
14
19
1>
1C
1P
1U
1X
#8480000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#8490000000
1!
1'
14
19
1>
1C
1P
1U
#8500000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#8510000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#8520000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#8530000000
1!
b0100 %
b1111110 &
1'
b0100 +
b1111110 ,
14
19
1>
1C
b0100 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#8540000000
0!
1#
0'
1)
04
09
1:
0>
0C
b0 K
0P
0U
b0 Y
#8550000000
#8560000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#8570000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#8580000000
1!
1'
14
19
1>
1C
1P
1U
#8590000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#8600000000
1!
1'
14
19
1>
1C
1P
1U
1X
#8610000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#8620000000
1!
1'
14
19
1>
1C
1P
1U
#8630000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#8640000000
1!
1'
14
19
1>
1C
1P
1U
#8650000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#8660000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#8670000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#8680000000
1!
1'
14
19
1>
1C
1P
1U
#8690000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#8700000000
1!
1'
14
19
1>
1C
1P
1U
#8710000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#8720000000
1!
1'
14
19
1>
1C
1P
1U
1X
#8730000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#8740000000
1!
1'
14
19
1>
1C
1P
1U
#8750000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#8760000000
1!
1'
14
19
1>
1C
1P
1U
#8770000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#8780000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#8790000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#8800000000
1!
1'
14
19
1>
1C
1P
1U
#8810000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#8820000000
1!
1'
14
19
1>
1C
1P
1U
#8830000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#8840000000
1!
1'
14
19
1>
1C
1P
1U
1X
#8850000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#8860000000
1!
1'
14
19
1>
1C
1P
1U
#8870000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#8880000000
1!
1'
14
19
1>
1C
1P
1U
#8890000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#8900000000
1!
b0010 %
b0110000 &
1'
b0010 +
b0110000 ,
14
19
1>
1C
b0010 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#8910000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#8920000000
1!
1'
14
19
1>
1C
1P
1U
#8930000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#8940000000
1!
1'
14
19
1>
1C
1P
1U
#8950000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#8960000000
1!
1'
14
19
1>
1C
1P
1U
1X
#8970000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#8980000000
1!
1'
14
19
1>
1C
1P
1U
#8990000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#9000000000
1!
1'
14
19
1>
1C
1P
1U
#9010000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#9020000000
1!
b0100 %
b1111110 &
1'
b0100 +
b1111110 ,
14
19
1>
1C
b0100 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#9030000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#9040000000
1!
1'
14
19
1>
1C
1P
1U
#9050000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#9060000000
1!
1'
14
19
1>
1C
1P
1U
#9070000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#9080000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
1X
#9090000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#9100000000
1!
1'
14
19
1>
1C
1P
1U
#9110000000
0!
1#
0'
1)
04
09
1:
0>
0C
b100 K
0P
0U
b100 Y
#9120000000
#9130000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
#9140000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#9150000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#9160000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#9170000000
1!
1'
14
19
1>
1C
1P
1U
#9180000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#9190000000
1!
1'
14
19
1>
1C
1P
1U
#9200000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#9210000000
1!
1'
14
19
1>
1C
1P
1U
1X
#9220000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#9230000000
1!
1'
14
19
1>
1C
1P
1U
#9240000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#9250000000
1!
1'
14
19
1>
1C
1P
1U
#9260000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#9270000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#9280000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#9290000000
1!
1'
14
19
1>
1C
1P
1U
#9300000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#9310000000
1!
1'
14
19
1>
1C
1P
1U
#9320000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#9330000000
1!
1'
14
19
1>
1C
1P
1U
1X
#9340000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#9350000000
1!
1'
14
19
1>
1C
1P
1U
#9360000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#9370000000
1!
1'
14
19
1>
1C
1P
1U
#9380000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#9390000000
1!
b0010 %
b0110000 &
1'
b0010 +
b0110000 ,
14
19
1>
1C
b0010 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#9400000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#9410000000
1!
1'
14
19
1>
1C
1P
1U
#9420000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#9430000000
1!
1'
14
19
1>
1C
1P
1U
#9440000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#9450000000
1!
1'
14
19
1>
1C
1P
1U
1X
#9460000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#9470000000
1!
1'
14
19
1>
1C
1P
1U
#9480000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#9490000000
1!
1'
14
19
1>
1C
1P
1U
#9500000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#9510000000
1!
b0100 %
b1111110 &
1'
b0100 +
b1111110 ,
14
19
1>
1C
b0100 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
#9520000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#9530000000
1!
1'
14
19
1>
1C
1P
1U
#9540000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#9550000000
1!
1'
14
19
1>
1C
1P
1U
#9560000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#9570000000
1!
1'
14
19
1>
1C
1P
1U
1X
#9580000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#9590000000
1!
1'
14
19
1>
1C
1P
1U
#9600000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#9610000000
1!
1'
14
19
1>
1C
1P
1U
#9620000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#9630000000
1!
b1000 %
1'
b1000 +
14
19
1>
1C
b1000 I
1P
1U
0X
#9640000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#9650000000
1!
0#
1'
0)
0.
14
19
0:
0;
0<
0=
1>
1C
1P
1U
#9660000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#9670000000
1!
1'
14
19
1>
1C
1P
1U
#9680000000
0!
1#
0'
1)
04
09
1:
0>
0C
b10 K
0P
0U
b10 Y
#9690000000
#9700000000
1!
1'
1.
14
19
1;
1<
1=
1>
1C
1P
1U
1X
#9710000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#9720000000
1!
1'
14
19
1>
1C
1P
1U
#9730000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#9740000000
1!
1'
14
19
1>
1C
1P
1U
#9750000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#9760000000
1!
b0001 %
1'
b0001 +
14
19
1>
1C
b0001 I
1P
1U
0X
#9770000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#9780000000
1!
1'
14
19
1>
1C
1P
1U
#9790000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#9800000000
1!
1'
14
19
1>
1C
1P
1U
#9810000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#9820000000
1!
1'
14
19
1>
1C
1P
1U
1X
#9830000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#9840000000
1!
1'
14
19
1>
1C
1P
1U
#9850000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#9860000000
1!
1'
14
19
1>
1C
1P
1U
#9870000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#9880000000
1!
b0010 %
b0110000 &
1'
b0010 +
b0110000 ,
14
19
1>
1C
b0010 I
b0110000 J
b0001 O
1P
1U
0X
b0110000 Z
b0001 [
#9890000000
0!
0'
04
09
0>
0C
b0 K
0P
0U
b0 Y
#9900000000
1!
1'
14
19
1>
1C
1P
1U
#9910000000
0!
0'
04
09
0>
0C
b1 K
0P
0U
b1 Y
#9920000000
1!
1'
14
19
1>
1C
1P
1U
#9930000000
0!
0'
04
09
0>
0C
b10 K
0P
0U
b10 Y
#9940000000
1!
1'
14
19
1>
1C
1P
1U
1X
#9950000000
0!
0'
04
09
0>
0C
b11 K
0P
0U
b11 Y
#9960000000
1!
1'
14
19
1>
1C
1P
1U
#9970000000
0!
0'
04
09
0>
0C
b100 K
0P
0U
b100 Y
#9980000000
1!
1'
14
19
1>
1C
1P
1U
#9990000000
0!
0'
04
09
0>
0C
b101 K
0P
0U
b101 Y
#10000000000
1!
b0100 %
b1111110 &
1'
b0100 +
b1111110 ,
14
19
1>
1C
b0100 I
b1111110 J
b0000 O
1P
1U
0X
b1111110 Z
b0000 [
