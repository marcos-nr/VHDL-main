$date
  Mon Jun 24 21:54:31 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_falso_spi $end
$var reg 1 ! clk $end
$var reg 1 " in1 $end
$var reg 1 # in2 $end
$var reg 1 $ in3 $end
$var reg 1 % pwm_o $end
$scope module uud $end
$var reg 1 & clk $end
$var reg 1 ' in1 $end
$var reg 1 ( in2 $end
$var reg 1 ) in3 $end
$var reg 1 * pwm_o $end
$var integer 32 + duty $end
$scope module inst_pwm0 $end
$var reg 1 , clk $end
$var reg 1 - reset $end
$var reg 1 . enable $end
$var reg 1 / cout $end
$var integer 32 0 q $end
$var integer 32 1 duty $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
U!
1"
U#
U$
U%
U&
1'
U(
U)
U*
b0 +
U,
0-
1.
U/
b0 0
b0 1
#50000000
0"
0'
#60000000
1#
1(
b101111101100100 +
b101111101100100 1
#110000000
0#
0(
#120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#170000000
0$
0)
#180000000
1"
1'
b0 +
b0 1
#230000000
0"
0'
#240000000
1#
1(
b101111101100100 +
b101111101100100 1
#290000000
0#
0(
#300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#350000000
0$
0)
#360000000
1"
1'
b0 +
b0 1
#410000000
0"
0'
#420000000
1#
1(
b101111101100100 +
b101111101100100 1
#470000000
0#
0(
#480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#530000000
0$
0)
#540000000
1"
1'
b0 +
b0 1
#590000000
0"
0'
#600000000
1#
1(
b101111101100100 +
b101111101100100 1
#650000000
0#
0(
#660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#710000000
0$
0)
#720000000
1"
1'
b0 +
b0 1
#770000000
0"
0'
#780000000
1#
1(
b101111101100100 +
b101111101100100 1
#830000000
0#
0(
#840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#890000000
0$
0)
#900000000
1"
1'
b0 +
b0 1
#950000000
0"
0'
#960000000
1#
1(
b101111101100100 +
b101111101100100 1
#1010000000
0#
0(
#1020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#1070000000
0$
0)
#1080000000
1"
1'
b0 +
b0 1
#1130000000
0"
0'
#1140000000
1#
1(
b101111101100100 +
b101111101100100 1
#1190000000
0#
0(
#1200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#1250000000
0$
0)
#1260000000
1"
1'
b0 +
b0 1
#1310000000
0"
0'
#1320000000
1#
1(
b101111101100100 +
b101111101100100 1
#1370000000
0#
0(
#1380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#1430000000
0$
0)
#1440000000
1"
1'
b0 +
b0 1
#1490000000
0"
0'
#1500000000
1#
1(
b101111101100100 +
b101111101100100 1
#1550000000
0#
0(
#1560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#1610000000
0$
0)
#1620000000
1"
1'
b0 +
b0 1
#1670000000
0"
0'
#1680000000
1#
1(
b101111101100100 +
b101111101100100 1
#1730000000
0#
0(
#1740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#1790000000
0$
0)
#1800000000
1"
1'
b0 +
b0 1
#1850000000
0"
0'
#1860000000
1#
1(
b101111101100100 +
b101111101100100 1
#1910000000
0#
0(
#1920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#1970000000
0$
0)
#1980000000
1"
1'
b0 +
b0 1
#2030000000
0"
0'
#2040000000
1#
1(
b101111101100100 +
b101111101100100 1
#2090000000
0#
0(
#2100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#2150000000
0$
0)
#2160000000
1"
1'
b0 +
b0 1
#2210000000
0"
0'
#2220000000
1#
1(
b101111101100100 +
b101111101100100 1
#2270000000
0#
0(
#2280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#2330000000
0$
0)
#2340000000
1"
1'
b0 +
b0 1
#2390000000
0"
0'
#2400000000
1#
1(
b101111101100100 +
b101111101100100 1
#2450000000
0#
0(
#2460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#2510000000
0$
0)
#2520000000
1"
1'
b0 +
b0 1
#2570000000
0"
0'
#2580000000
1#
1(
b101111101100100 +
b101111101100100 1
#2630000000
0#
0(
#2640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#2690000000
0$
0)
#2700000000
1"
1'
b0 +
b0 1
#2750000000
0"
0'
#2760000000
1#
1(
b101111101100100 +
b101111101100100 1
#2810000000
0#
0(
#2820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#2870000000
0$
0)
#2880000000
1"
1'
b0 +
b0 1
#2930000000
0"
0'
#2940000000
1#
1(
b101111101100100 +
b101111101100100 1
#2990000000
0#
0(
#3000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#3050000000
0$
0)
#3060000000
1"
1'
b0 +
b0 1
#3110000000
0"
0'
#3120000000
1#
1(
b101111101100100 +
b101111101100100 1
#3170000000
0#
0(
#3180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#3230000000
0$
0)
#3240000000
1"
1'
b0 +
b0 1
#3290000000
0"
0'
#3300000000
1#
1(
b101111101100100 +
b101111101100100 1
#3350000000
0#
0(
#3360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#3410000000
0$
0)
#3420000000
1"
1'
b0 +
b0 1
#3470000000
0"
0'
#3480000000
1#
1(
b101111101100100 +
b101111101100100 1
#3530000000
0#
0(
#3540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#3590000000
0$
0)
#3600000000
1"
1'
b0 +
b0 1
#3650000000
0"
0'
#3660000000
1#
1(
b101111101100100 +
b101111101100100 1
#3710000000
0#
0(
#3720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#3770000000
0$
0)
#3780000000
1"
1'
b0 +
b0 1
#3830000000
0"
0'
#3840000000
1#
1(
b101111101100100 +
b101111101100100 1
#3890000000
0#
0(
#3900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#3950000000
0$
0)
#3960000000
1"
1'
b0 +
b0 1
#4010000000
0"
0'
#4020000000
1#
1(
b101111101100100 +
b101111101100100 1
#4070000000
0#
0(
#4080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#4130000000
0$
0)
#4140000000
1"
1'
b0 +
b0 1
#4190000000
0"
0'
#4200000000
1#
1(
b101111101100100 +
b101111101100100 1
#4250000000
0#
0(
#4260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#4310000000
0$
0)
#4320000000
1"
1'
b0 +
b0 1
#4370000000
0"
0'
#4380000000
1#
1(
b101111101100100 +
b101111101100100 1
#4430000000
0#
0(
#4440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#4490000000
0$
0)
#4500000000
1"
1'
b0 +
b0 1
#4550000000
0"
0'
#4560000000
1#
1(
b101111101100100 +
b101111101100100 1
#4610000000
0#
0(
#4620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#4670000000
0$
0)
#4680000000
1"
1'
b0 +
b0 1
#4730000000
0"
0'
#4740000000
1#
1(
b101111101100100 +
b101111101100100 1
#4790000000
0#
0(
#4800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#4850000000
0$
0)
#4860000000
1"
1'
b0 +
b0 1
#4910000000
0"
0'
#4920000000
1#
1(
b101111101100100 +
b101111101100100 1
#4970000000
0#
0(
#4980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#5030000000
0$
0)
#5040000000
1"
1'
b0 +
b0 1
#5090000000
0"
0'
#5100000000
1#
1(
b101111101100100 +
b101111101100100 1
#5150000000
0#
0(
#5160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#5210000000
0$
0)
#5220000000
1"
1'
b0 +
b0 1
#5270000000
0"
0'
#5280000000
1#
1(
b101111101100100 +
b101111101100100 1
#5330000000
0#
0(
#5340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#5390000000
0$
0)
#5400000000
1"
1'
b0 +
b0 1
#5450000000
0"
0'
#5460000000
1#
1(
b101111101100100 +
b101111101100100 1
#5510000000
0#
0(
#5520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#5570000000
0$
0)
#5580000000
1"
1'
b0 +
b0 1
#5630000000
0"
0'
#5640000000
1#
1(
b101111101100100 +
b101111101100100 1
#5690000000
0#
0(
#5700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#5750000000
0$
0)
#5760000000
1"
1'
b0 +
b0 1
#5810000000
0"
0'
#5820000000
1#
1(
b101111101100100 +
b101111101100100 1
#5870000000
0#
0(
#5880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#5930000000
0$
0)
#5940000000
1"
1'
b0 +
b0 1
#5990000000
0"
0'
#6000000000
1#
1(
b101111101100100 +
b101111101100100 1
#6050000000
0#
0(
#6060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#6110000000
0$
0)
#6120000000
1"
1'
b0 +
b0 1
#6170000000
0"
0'
#6180000000
1#
1(
b101111101100100 +
b101111101100100 1
#6230000000
0#
0(
#6240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#6290000000
0$
0)
#6300000000
1"
1'
b0 +
b0 1
#6350000000
0"
0'
#6360000000
1#
1(
b101111101100100 +
b101111101100100 1
#6410000000
0#
0(
#6420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#6470000000
0$
0)
#6480000000
1"
1'
b0 +
b0 1
#6530000000
0"
0'
#6540000000
1#
1(
b101111101100100 +
b101111101100100 1
#6590000000
0#
0(
#6600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#6650000000
0$
0)
#6660000000
1"
1'
b0 +
b0 1
#6710000000
0"
0'
#6720000000
1#
1(
b101111101100100 +
b101111101100100 1
#6770000000
0#
0(
#6780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#6830000000
0$
0)
#6840000000
1"
1'
b0 +
b0 1
#6890000000
0"
0'
#6900000000
1#
1(
b101111101100100 +
b101111101100100 1
#6950000000
0#
0(
#6960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#7010000000
0$
0)
#7020000000
1"
1'
b0 +
b0 1
#7070000000
0"
0'
#7080000000
1#
1(
b101111101100100 +
b101111101100100 1
#7130000000
0#
0(
#7140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#7190000000
0$
0)
#7200000000
1"
1'
b0 +
b0 1
#7250000000
0"
0'
#7260000000
1#
1(
b101111101100100 +
b101111101100100 1
#7310000000
0#
0(
#7320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#7370000000
0$
0)
#7380000000
1"
1'
b0 +
b0 1
#7430000000
0"
0'
#7440000000
1#
1(
b101111101100100 +
b101111101100100 1
#7490000000
0#
0(
#7500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#7550000000
0$
0)
#7560000000
1"
1'
b0 +
b0 1
#7610000000
0"
0'
#7620000000
1#
1(
b101111101100100 +
b101111101100100 1
#7670000000
0#
0(
#7680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#7730000000
0$
0)
#7740000000
1"
1'
b0 +
b0 1
#7790000000
0"
0'
#7800000000
1#
1(
b101111101100100 +
b101111101100100 1
#7850000000
0#
0(
#7860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#7910000000
0$
0)
#7920000000
1"
1'
b0 +
b0 1
#7970000000
0"
0'
#7980000000
1#
1(
b101111101100100 +
b101111101100100 1
#8030000000
0#
0(
#8040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#8090000000
0$
0)
#8100000000
1"
1'
b0 +
b0 1
#8150000000
0"
0'
#8160000000
1#
1(
b101111101100100 +
b101111101100100 1
#8210000000
0#
0(
#8220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#8270000000
0$
0)
#8280000000
1"
1'
b0 +
b0 1
#8330000000
0"
0'
#8340000000
1#
1(
b101111101100100 +
b101111101100100 1
#8390000000
0#
0(
#8400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#8450000000
0$
0)
#8460000000
1"
1'
b0 +
b0 1
#8510000000
0"
0'
#8520000000
1#
1(
b101111101100100 +
b101111101100100 1
#8570000000
0#
0(
#8580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#8630000000
0$
0)
#8640000000
1"
1'
b0 +
b0 1
#8690000000
0"
0'
#8700000000
1#
1(
b101111101100100 +
b101111101100100 1
#8750000000
0#
0(
#8760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#8810000000
0$
0)
#8820000000
1"
1'
b0 +
b0 1
#8870000000
0"
0'
#8880000000
1#
1(
b101111101100100 +
b101111101100100 1
#8930000000
0#
0(
#8940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#8990000000
0$
0)
#9000000000
1"
1'
b0 +
b0 1
#9050000000
0"
0'
#9060000000
1#
1(
b101111101100100 +
b101111101100100 1
#9110000000
0#
0(
#9120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#9170000000
0$
0)
#9180000000
1"
1'
b0 +
b0 1
#9230000000
0"
0'
#9240000000
1#
1(
b101111101100100 +
b101111101100100 1
#9290000000
0#
0(
#9300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#9350000000
0$
0)
#9360000000
1"
1'
b0 +
b0 1
#9410000000
0"
0'
#9420000000
1#
1(
b101111101100100 +
b101111101100100 1
#9470000000
0#
0(
#9480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#9530000000
0$
0)
#9540000000
1"
1'
b0 +
b0 1
#9590000000
0"
0'
#9600000000
1#
1(
b101111101100100 +
b101111101100100 1
#9650000000
0#
0(
#9660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#9710000000
0$
0)
#9720000000
1"
1'
b0 +
b0 1
#9770000000
0"
0'
#9780000000
1#
1(
b101111101100100 +
b101111101100100 1
#9830000000
0#
0(
#9840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#9890000000
0$
0)
#9900000000
1"
1'
b0 +
b0 1
#9950000000
0"
0'
#9960000000
1#
1(
b101111101100100 +
b101111101100100 1
#10010000000
0#
0(
#10020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#10070000000
0$
0)
#10080000000
1"
1'
b0 +
b0 1
#10130000000
0"
0'
#10140000000
1#
1(
b101111101100100 +
b101111101100100 1
#10190000000
0#
0(
#10200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#10250000000
0$
0)
#10260000000
1"
1'
b0 +
b0 1
#10310000000
0"
0'
#10320000000
1#
1(
b101111101100100 +
b101111101100100 1
#10370000000
0#
0(
#10380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#10430000000
0$
0)
#10440000000
1"
1'
b0 +
b0 1
#10490000000
0"
0'
#10500000000
1#
1(
b101111101100100 +
b101111101100100 1
#10550000000
0#
0(
#10560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#10610000000
0$
0)
#10620000000
1"
1'
b0 +
b0 1
#10670000000
0"
0'
#10680000000
1#
1(
b101111101100100 +
b101111101100100 1
#10730000000
0#
0(
#10740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#10790000000
0$
0)
#10800000000
1"
1'
b0 +
b0 1
#10850000000
0"
0'
#10860000000
1#
1(
b101111101100100 +
b101111101100100 1
#10910000000
0#
0(
#10920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#10970000000
0$
0)
#10980000000
1"
1'
b0 +
b0 1
#11030000000
0"
0'
#11040000000
1#
1(
b101111101100100 +
b101111101100100 1
#11090000000
0#
0(
#11100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#11150000000
0$
0)
#11160000000
1"
1'
b0 +
b0 1
#11210000000
0"
0'
#11220000000
1#
1(
b101111101100100 +
b101111101100100 1
#11270000000
0#
0(
#11280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#11330000000
0$
0)
#11340000000
1"
1'
b0 +
b0 1
#11390000000
0"
0'
#11400000000
1#
1(
b101111101100100 +
b101111101100100 1
#11450000000
0#
0(
#11460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#11510000000
0$
0)
#11520000000
1"
1'
b0 +
b0 1
#11570000000
0"
0'
#11580000000
1#
1(
b101111101100100 +
b101111101100100 1
#11630000000
0#
0(
#11640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#11690000000
0$
0)
#11700000000
1"
1'
b0 +
b0 1
#11750000000
0"
0'
#11760000000
1#
1(
b101111101100100 +
b101111101100100 1
#11810000000
0#
0(
#11820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#11870000000
0$
0)
#11880000000
1"
1'
b0 +
b0 1
#11930000000
0"
0'
#11940000000
1#
1(
b101111101100100 +
b101111101100100 1
#11990000000
0#
0(
#12000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#12050000000
0$
0)
#12060000000
1"
1'
b0 +
b0 1
#12110000000
0"
0'
#12120000000
1#
1(
b101111101100100 +
b101111101100100 1
#12170000000
0#
0(
#12180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#12230000000
0$
0)
#12240000000
1"
1'
b0 +
b0 1
#12290000000
0"
0'
#12300000000
1#
1(
b101111101100100 +
b101111101100100 1
#12350000000
0#
0(
#12360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#12410000000
0$
0)
#12420000000
1"
1'
b0 +
b0 1
#12470000000
0"
0'
#12480000000
1#
1(
b101111101100100 +
b101111101100100 1
#12530000000
0#
0(
#12540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#12590000000
0$
0)
#12600000000
1"
1'
b0 +
b0 1
#12650000000
0"
0'
#12660000000
1#
1(
b101111101100100 +
b101111101100100 1
#12710000000
0#
0(
#12720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#12770000000
0$
0)
#12780000000
1"
1'
b0 +
b0 1
#12830000000
0"
0'
#12840000000
1#
1(
b101111101100100 +
b101111101100100 1
#12890000000
0#
0(
#12900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#12950000000
0$
0)
#12960000000
1"
1'
b0 +
b0 1
#13010000000
0"
0'
#13020000000
1#
1(
b101111101100100 +
b101111101100100 1
#13070000000
0#
0(
#13080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#13130000000
0$
0)
#13140000000
1"
1'
b0 +
b0 1
#13190000000
0"
0'
#13200000000
1#
1(
b101111101100100 +
b101111101100100 1
#13250000000
0#
0(
#13260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#13310000000
0$
0)
#13320000000
1"
1'
b0 +
b0 1
#13370000000
0"
0'
#13380000000
1#
1(
b101111101100100 +
b101111101100100 1
#13430000000
0#
0(
#13440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#13490000000
0$
0)
#13500000000
1"
1'
b0 +
b0 1
#13550000000
0"
0'
#13560000000
1#
1(
b101111101100100 +
b101111101100100 1
#13610000000
0#
0(
#13620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#13670000000
0$
0)
#13680000000
1"
1'
b0 +
b0 1
#13730000000
0"
0'
#13740000000
1#
1(
b101111101100100 +
b101111101100100 1
#13790000000
0#
0(
#13800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#13850000000
0$
0)
#13860000000
1"
1'
b0 +
b0 1
#13910000000
0"
0'
#13920000000
1#
1(
b101111101100100 +
b101111101100100 1
#13970000000
0#
0(
#13980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#14030000000
0$
0)
#14040000000
1"
1'
b0 +
b0 1
#14090000000
0"
0'
#14100000000
1#
1(
b101111101100100 +
b101111101100100 1
#14150000000
0#
0(
#14160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#14210000000
0$
0)
#14220000000
1"
1'
b0 +
b0 1
#14270000000
0"
0'
#14280000000
1#
1(
b101111101100100 +
b101111101100100 1
#14330000000
0#
0(
#14340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#14390000000
0$
0)
#14400000000
1"
1'
b0 +
b0 1
#14450000000
0"
0'
#14460000000
1#
1(
b101111101100100 +
b101111101100100 1
#14510000000
0#
0(
#14520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#14570000000
0$
0)
#14580000000
1"
1'
b0 +
b0 1
#14630000000
0"
0'
#14640000000
1#
1(
b101111101100100 +
b101111101100100 1
#14690000000
0#
0(
#14700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#14750000000
0$
0)
#14760000000
1"
1'
b0 +
b0 1
#14810000000
0"
0'
#14820000000
1#
1(
b101111101100100 +
b101111101100100 1
#14870000000
0#
0(
#14880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#14930000000
0$
0)
#14940000000
1"
1'
b0 +
b0 1
#14990000000
0"
0'
#15000000000
1#
1(
b101111101100100 +
b101111101100100 1
#15050000000
0#
0(
#15060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#15110000000
0$
0)
#15120000000
1"
1'
b0 +
b0 1
#15170000000
0"
0'
#15180000000
1#
1(
b101111101100100 +
b101111101100100 1
#15230000000
0#
0(
#15240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#15290000000
0$
0)
#15300000000
1"
1'
b0 +
b0 1
#15350000000
0"
0'
#15360000000
1#
1(
b101111101100100 +
b101111101100100 1
#15410000000
0#
0(
#15420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#15470000000
0$
0)
#15480000000
1"
1'
b0 +
b0 1
#15530000000
0"
0'
#15540000000
1#
1(
b101111101100100 +
b101111101100100 1
#15590000000
0#
0(
#15600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#15650000000
0$
0)
#15660000000
1"
1'
b0 +
b0 1
#15710000000
0"
0'
#15720000000
1#
1(
b101111101100100 +
b101111101100100 1
#15770000000
0#
0(
#15780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#15830000000
0$
0)
#15840000000
1"
1'
b0 +
b0 1
#15890000000
0"
0'
#15900000000
1#
1(
b101111101100100 +
b101111101100100 1
#15950000000
0#
0(
#15960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#16010000000
0$
0)
#16020000000
1"
1'
b0 +
b0 1
#16070000000
0"
0'
#16080000000
1#
1(
b101111101100100 +
b101111101100100 1
#16130000000
0#
0(
#16140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#16190000000
0$
0)
#16200000000
1"
1'
b0 +
b0 1
#16250000000
0"
0'
#16260000000
1#
1(
b101111101100100 +
b101111101100100 1
#16310000000
0#
0(
#16320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#16370000000
0$
0)
#16380000000
1"
1'
b0 +
b0 1
#16430000000
0"
0'
#16440000000
1#
1(
b101111101100100 +
b101111101100100 1
#16490000000
0#
0(
#16500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#16550000000
0$
0)
#16560000000
1"
1'
b0 +
b0 1
#16610000000
0"
0'
#16620000000
1#
1(
b101111101100100 +
b101111101100100 1
#16670000000
0#
0(
#16680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#16730000000
0$
0)
#16740000000
1"
1'
b0 +
b0 1
#16790000000
0"
0'
#16800000000
1#
1(
b101111101100100 +
b101111101100100 1
#16850000000
0#
0(
#16860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#16910000000
0$
0)
#16920000000
1"
1'
b0 +
b0 1
#16970000000
0"
0'
#16980000000
1#
1(
b101111101100100 +
b101111101100100 1
#17030000000
0#
0(
#17040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#17090000000
0$
0)
#17100000000
1"
1'
b0 +
b0 1
#17150000000
0"
0'
#17160000000
1#
1(
b101111101100100 +
b101111101100100 1
#17210000000
0#
0(
#17220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#17270000000
0$
0)
#17280000000
1"
1'
b0 +
b0 1
#17330000000
0"
0'
#17340000000
1#
1(
b101111101100100 +
b101111101100100 1
#17390000000
0#
0(
#17400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#17450000000
0$
0)
#17460000000
1"
1'
b0 +
b0 1
#17510000000
0"
0'
#17520000000
1#
1(
b101111101100100 +
b101111101100100 1
#17570000000
0#
0(
#17580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#17630000000
0$
0)
#17640000000
1"
1'
b0 +
b0 1
#17690000000
0"
0'
#17700000000
1#
1(
b101111101100100 +
b101111101100100 1
#17750000000
0#
0(
#17760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#17810000000
0$
0)
#17820000000
1"
1'
b0 +
b0 1
#17870000000
0"
0'
#17880000000
1#
1(
b101111101100100 +
b101111101100100 1
#17930000000
0#
0(
#17940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#17990000000
0$
0)
#18000000000
1"
1'
b0 +
b0 1
#18050000000
0"
0'
#18060000000
1#
1(
b101111101100100 +
b101111101100100 1
#18110000000
0#
0(
#18120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#18170000000
0$
0)
#18180000000
1"
1'
b0 +
b0 1
#18230000000
0"
0'
#18240000000
1#
1(
b101111101100100 +
b101111101100100 1
#18290000000
0#
0(
#18300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#18350000000
0$
0)
#18360000000
1"
1'
b0 +
b0 1
#18410000000
0"
0'
#18420000000
1#
1(
b101111101100100 +
b101111101100100 1
#18470000000
0#
0(
#18480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#18530000000
0$
0)
#18540000000
1"
1'
b0 +
b0 1
#18590000000
0"
0'
#18600000000
1#
1(
b101111101100100 +
b101111101100100 1
#18650000000
0#
0(
#18660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#18710000000
0$
0)
#18720000000
1"
1'
b0 +
b0 1
#18770000000
0"
0'
#18780000000
1#
1(
b101111101100100 +
b101111101100100 1
#18830000000
0#
0(
#18840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#18890000000
0$
0)
#18900000000
1"
1'
b0 +
b0 1
#18950000000
0"
0'
#18960000000
1#
1(
b101111101100100 +
b101111101100100 1
#19010000000
0#
0(
#19020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#19070000000
0$
0)
#19080000000
1"
1'
b0 +
b0 1
#19130000000
0"
0'
#19140000000
1#
1(
b101111101100100 +
b101111101100100 1
#19190000000
0#
0(
#19200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#19250000000
0$
0)
#19260000000
1"
1'
b0 +
b0 1
#19310000000
0"
0'
#19320000000
1#
1(
b101111101100100 +
b101111101100100 1
#19370000000
0#
0(
#19380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#19430000000
0$
0)
#19440000000
1"
1'
b0 +
b0 1
#19490000000
0"
0'
#19500000000
1#
1(
b101111101100100 +
b101111101100100 1
#19550000000
0#
0(
#19560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#19610000000
0$
0)
#19620000000
1"
1'
b0 +
b0 1
#19670000000
0"
0'
#19680000000
1#
1(
b101111101100100 +
b101111101100100 1
#19730000000
0#
0(
#19740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#19790000000
0$
0)
#19800000000
1"
1'
b0 +
b0 1
#19850000000
0"
0'
#19860000000
1#
1(
b101111101100100 +
b101111101100100 1
#19910000000
0#
0(
#19920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#19970000000
0$
0)
#19980000000
1"
1'
b0 +
b0 1
#20030000000
0"
0'
#20040000000
1#
1(
b101111101100100 +
b101111101100100 1
#20090000000
0#
0(
#20100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#20150000000
0$
0)
#20160000000
1"
1'
b0 +
b0 1
#20210000000
0"
0'
#20220000000
1#
1(
b101111101100100 +
b101111101100100 1
#20270000000
0#
0(
#20280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#20330000000
0$
0)
#20340000000
1"
1'
b0 +
b0 1
#20390000000
0"
0'
#20400000000
1#
1(
b101111101100100 +
b101111101100100 1
#20450000000
0#
0(
#20460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#20510000000
0$
0)
#20520000000
1"
1'
b0 +
b0 1
#20570000000
0"
0'
#20580000000
1#
1(
b101111101100100 +
b101111101100100 1
#20630000000
0#
0(
#20640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#20690000000
0$
0)
#20700000000
1"
1'
b0 +
b0 1
#20750000000
0"
0'
#20760000000
1#
1(
b101111101100100 +
b101111101100100 1
#20810000000
0#
0(
#20820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#20870000000
0$
0)
#20880000000
1"
1'
b0 +
b0 1
#20930000000
0"
0'
#20940000000
1#
1(
b101111101100100 +
b101111101100100 1
#20990000000
0#
0(
#21000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#21050000000
0$
0)
#21060000000
1"
1'
b0 +
b0 1
#21110000000
0"
0'
#21120000000
1#
1(
b101111101100100 +
b101111101100100 1
#21170000000
0#
0(
#21180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#21230000000
0$
0)
#21240000000
1"
1'
b0 +
b0 1
#21290000000
0"
0'
#21300000000
1#
1(
b101111101100100 +
b101111101100100 1
#21350000000
0#
0(
#21360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#21410000000
0$
0)
#21420000000
1"
1'
b0 +
b0 1
#21470000000
0"
0'
#21480000000
1#
1(
b101111101100100 +
b101111101100100 1
#21530000000
0#
0(
#21540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#21590000000
0$
0)
#21600000000
1"
1'
b0 +
b0 1
#21650000000
0"
0'
#21660000000
1#
1(
b101111101100100 +
b101111101100100 1
#21710000000
0#
0(
#21720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#21770000000
0$
0)
#21780000000
1"
1'
b0 +
b0 1
#21830000000
0"
0'
#21840000000
1#
1(
b101111101100100 +
b101111101100100 1
#21890000000
0#
0(
#21900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#21950000000
0$
0)
#21960000000
1"
1'
b0 +
b0 1
#22010000000
0"
0'
#22020000000
1#
1(
b101111101100100 +
b101111101100100 1
#22070000000
0#
0(
#22080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#22130000000
0$
0)
#22140000000
1"
1'
b0 +
b0 1
#22190000000
0"
0'
#22200000000
1#
1(
b101111101100100 +
b101111101100100 1
#22250000000
0#
0(
#22260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#22310000000
0$
0)
#22320000000
1"
1'
b0 +
b0 1
#22370000000
0"
0'
#22380000000
1#
1(
b101111101100100 +
b101111101100100 1
#22430000000
0#
0(
#22440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#22490000000
0$
0)
#22500000000
1"
1'
b0 +
b0 1
#22550000000
0"
0'
#22560000000
1#
1(
b101111101100100 +
b101111101100100 1
#22610000000
0#
0(
#22620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#22670000000
0$
0)
#22680000000
1"
1'
b0 +
b0 1
#22730000000
0"
0'
#22740000000
1#
1(
b101111101100100 +
b101111101100100 1
#22790000000
0#
0(
#22800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#22850000000
0$
0)
#22860000000
1"
1'
b0 +
b0 1
#22910000000
0"
0'
#22920000000
1#
1(
b101111101100100 +
b101111101100100 1
#22970000000
0#
0(
#22980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#23030000000
0$
0)
#23040000000
1"
1'
b0 +
b0 1
#23090000000
0"
0'
#23100000000
1#
1(
b101111101100100 +
b101111101100100 1
#23150000000
0#
0(
#23160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#23210000000
0$
0)
#23220000000
1"
1'
b0 +
b0 1
#23270000000
0"
0'
#23280000000
1#
1(
b101111101100100 +
b101111101100100 1
#23330000000
0#
0(
#23340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#23390000000
0$
0)
#23400000000
1"
1'
b0 +
b0 1
#23450000000
0"
0'
#23460000000
1#
1(
b101111101100100 +
b101111101100100 1
#23510000000
0#
0(
#23520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#23570000000
0$
0)
#23580000000
1"
1'
b0 +
b0 1
#23630000000
0"
0'
#23640000000
1#
1(
b101111101100100 +
b101111101100100 1
#23690000000
0#
0(
#23700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#23750000000
0$
0)
#23760000000
1"
1'
b0 +
b0 1
#23810000000
0"
0'
#23820000000
1#
1(
b101111101100100 +
b101111101100100 1
#23870000000
0#
0(
#23880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#23930000000
0$
0)
#23940000000
1"
1'
b0 +
b0 1
#23990000000
0"
0'
#24000000000
1#
1(
b101111101100100 +
b101111101100100 1
#24050000000
0#
0(
#24060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#24110000000
0$
0)
#24120000000
1"
1'
b0 +
b0 1
#24170000000
0"
0'
#24180000000
1#
1(
b101111101100100 +
b101111101100100 1
#24230000000
0#
0(
#24240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#24290000000
0$
0)
#24300000000
1"
1'
b0 +
b0 1
#24350000000
0"
0'
#24360000000
1#
1(
b101111101100100 +
b101111101100100 1
#24410000000
0#
0(
#24420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#24470000000
0$
0)
#24480000000
1"
1'
b0 +
b0 1
#24530000000
0"
0'
#24540000000
1#
1(
b101111101100100 +
b101111101100100 1
#24590000000
0#
0(
#24600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#24650000000
0$
0)
#24660000000
1"
1'
b0 +
b0 1
#24710000000
0"
0'
#24720000000
1#
1(
b101111101100100 +
b101111101100100 1
#24770000000
0#
0(
#24780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#24830000000
0$
0)
#24840000000
1"
1'
b0 +
b0 1
#24890000000
0"
0'
#24900000000
1#
1(
b101111101100100 +
b101111101100100 1
#24950000000
0#
0(
#24960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#25010000000
0$
0)
#25020000000
1"
1'
b0 +
b0 1
#25070000000
0"
0'
#25080000000
1#
1(
b101111101100100 +
b101111101100100 1
#25130000000
0#
0(
#25140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#25190000000
0$
0)
#25200000000
1"
1'
b0 +
b0 1
#25250000000
0"
0'
#25260000000
1#
1(
b101111101100100 +
b101111101100100 1
#25310000000
0#
0(
#25320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#25370000000
0$
0)
#25380000000
1"
1'
b0 +
b0 1
#25430000000
0"
0'
#25440000000
1#
1(
b101111101100100 +
b101111101100100 1
#25490000000
0#
0(
#25500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#25550000000
0$
0)
#25560000000
1"
1'
b0 +
b0 1
#25610000000
0"
0'
#25620000000
1#
1(
b101111101100100 +
b101111101100100 1
#25670000000
0#
0(
#25680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#25730000000
0$
0)
#25740000000
1"
1'
b0 +
b0 1
#25790000000
0"
0'
#25800000000
1#
1(
b101111101100100 +
b101111101100100 1
#25850000000
0#
0(
#25860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#25910000000
0$
0)
#25920000000
1"
1'
b0 +
b0 1
#25970000000
0"
0'
#25980000000
1#
1(
b101111101100100 +
b101111101100100 1
#26030000000
0#
0(
#26040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#26090000000
0$
0)
#26100000000
1"
1'
b0 +
b0 1
#26150000000
0"
0'
#26160000000
1#
1(
b101111101100100 +
b101111101100100 1
#26210000000
0#
0(
#26220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#26270000000
0$
0)
#26280000000
1"
1'
b0 +
b0 1
#26330000000
0"
0'
#26340000000
1#
1(
b101111101100100 +
b101111101100100 1
#26390000000
0#
0(
#26400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#26450000000
0$
0)
#26460000000
1"
1'
b0 +
b0 1
#26510000000
0"
0'
#26520000000
1#
1(
b101111101100100 +
b101111101100100 1
#26570000000
0#
0(
#26580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#26630000000
0$
0)
#26640000000
1"
1'
b0 +
b0 1
#26690000000
0"
0'
#26700000000
1#
1(
b101111101100100 +
b101111101100100 1
#26750000000
0#
0(
#26760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#26810000000
0$
0)
#26820000000
1"
1'
b0 +
b0 1
#26870000000
0"
0'
#26880000000
1#
1(
b101111101100100 +
b101111101100100 1
#26930000000
0#
0(
#26940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#26990000000
0$
0)
#27000000000
1"
1'
b0 +
b0 1
#27050000000
0"
0'
#27060000000
1#
1(
b101111101100100 +
b101111101100100 1
#27110000000
0#
0(
#27120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#27170000000
0$
0)
#27180000000
1"
1'
b0 +
b0 1
#27230000000
0"
0'
#27240000000
1#
1(
b101111101100100 +
b101111101100100 1
#27290000000
0#
0(
#27300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#27350000000
0$
0)
#27360000000
1"
1'
b0 +
b0 1
#27410000000
0"
0'
#27420000000
1#
1(
b101111101100100 +
b101111101100100 1
#27470000000
0#
0(
#27480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#27530000000
0$
0)
#27540000000
1"
1'
b0 +
b0 1
#27590000000
0"
0'
#27600000000
1#
1(
b101111101100100 +
b101111101100100 1
#27650000000
0#
0(
#27660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#27710000000
0$
0)
#27720000000
1"
1'
b0 +
b0 1
#27770000000
0"
0'
#27780000000
1#
1(
b101111101100100 +
b101111101100100 1
#27830000000
0#
0(
#27840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#27890000000
0$
0)
#27900000000
1"
1'
b0 +
b0 1
#27950000000
0"
0'
#27960000000
1#
1(
b101111101100100 +
b101111101100100 1
#28010000000
0#
0(
#28020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#28070000000
0$
0)
#28080000000
1"
1'
b0 +
b0 1
#28130000000
0"
0'
#28140000000
1#
1(
b101111101100100 +
b101111101100100 1
#28190000000
0#
0(
#28200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#28250000000
0$
0)
#28260000000
1"
1'
b0 +
b0 1
#28310000000
0"
0'
#28320000000
1#
1(
b101111101100100 +
b101111101100100 1
#28370000000
0#
0(
#28380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#28430000000
0$
0)
#28440000000
1"
1'
b0 +
b0 1
#28490000000
0"
0'
#28500000000
1#
1(
b101111101100100 +
b101111101100100 1
#28550000000
0#
0(
#28560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#28610000000
0$
0)
#28620000000
1"
1'
b0 +
b0 1
#28670000000
0"
0'
#28680000000
1#
1(
b101111101100100 +
b101111101100100 1
#28730000000
0#
0(
#28740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#28790000000
0$
0)
#28800000000
1"
1'
b0 +
b0 1
#28850000000
0"
0'
#28860000000
1#
1(
b101111101100100 +
b101111101100100 1
#28910000000
0#
0(
#28920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#28970000000
0$
0)
#28980000000
1"
1'
b0 +
b0 1
#29030000000
0"
0'
#29040000000
1#
1(
b101111101100100 +
b101111101100100 1
#29090000000
0#
0(
#29100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#29150000000
0$
0)
#29160000000
1"
1'
b0 +
b0 1
#29210000000
0"
0'
#29220000000
1#
1(
b101111101100100 +
b101111101100100 1
#29270000000
0#
0(
#29280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#29330000000
0$
0)
#29340000000
1"
1'
b0 +
b0 1
#29390000000
0"
0'
#29400000000
1#
1(
b101111101100100 +
b101111101100100 1
#29450000000
0#
0(
#29460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#29510000000
0$
0)
#29520000000
1"
1'
b0 +
b0 1
#29570000000
0"
0'
#29580000000
1#
1(
b101111101100100 +
b101111101100100 1
#29630000000
0#
0(
#29640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#29690000000
0$
0)
#29700000000
1"
1'
b0 +
b0 1
#29750000000
0"
0'
#29760000000
1#
1(
b101111101100100 +
b101111101100100 1
#29810000000
0#
0(
#29820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#29870000000
0$
0)
#29880000000
1"
1'
b0 +
b0 1
#29930000000
0"
0'
#29940000000
1#
1(
b101111101100100 +
b101111101100100 1
#29990000000
0#
0(
#30000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#30050000000
0$
0)
#30060000000
1"
1'
b0 +
b0 1
#30110000000
0"
0'
#30120000000
1#
1(
b101111101100100 +
b101111101100100 1
#30170000000
0#
0(
#30180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#30230000000
0$
0)
#30240000000
1"
1'
b0 +
b0 1
#30290000000
0"
0'
#30300000000
1#
1(
b101111101100100 +
b101111101100100 1
#30350000000
0#
0(
#30360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#30410000000
0$
0)
#30420000000
1"
1'
b0 +
b0 1
#30470000000
0"
0'
#30480000000
1#
1(
b101111101100100 +
b101111101100100 1
#30530000000
0#
0(
#30540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#30590000000
0$
0)
#30600000000
1"
1'
b0 +
b0 1
#30650000000
0"
0'
#30660000000
1#
1(
b101111101100100 +
b101111101100100 1
#30710000000
0#
0(
#30720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#30770000000
0$
0)
#30780000000
1"
1'
b0 +
b0 1
#30830000000
0"
0'
#30840000000
1#
1(
b101111101100100 +
b101111101100100 1
#30890000000
0#
0(
#30900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#30950000000
0$
0)
#30960000000
1"
1'
b0 +
b0 1
#31010000000
0"
0'
#31020000000
1#
1(
b101111101100100 +
b101111101100100 1
#31070000000
0#
0(
#31080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#31130000000
0$
0)
#31140000000
1"
1'
b0 +
b0 1
#31190000000
0"
0'
#31200000000
1#
1(
b101111101100100 +
b101111101100100 1
#31250000000
0#
0(
#31260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#31310000000
0$
0)
#31320000000
1"
1'
b0 +
b0 1
#31370000000
0"
0'
#31380000000
1#
1(
b101111101100100 +
b101111101100100 1
#31430000000
0#
0(
#31440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#31490000000
0$
0)
#31500000000
1"
1'
b0 +
b0 1
#31550000000
0"
0'
#31560000000
1#
1(
b101111101100100 +
b101111101100100 1
#31610000000
0#
0(
#31620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#31670000000
0$
0)
#31680000000
1"
1'
b0 +
b0 1
#31730000000
0"
0'
#31740000000
1#
1(
b101111101100100 +
b101111101100100 1
#31790000000
0#
0(
#31800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#31850000000
0$
0)
#31860000000
1"
1'
b0 +
b0 1
#31910000000
0"
0'
#31920000000
1#
1(
b101111101100100 +
b101111101100100 1
#31970000000
0#
0(
#31980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#32030000000
0$
0)
#32040000000
1"
1'
b0 +
b0 1
#32090000000
0"
0'
#32100000000
1#
1(
b101111101100100 +
b101111101100100 1
#32150000000
0#
0(
#32160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#32210000000
0$
0)
#32220000000
1"
1'
b0 +
b0 1
#32270000000
0"
0'
#32280000000
1#
1(
b101111101100100 +
b101111101100100 1
#32330000000
0#
0(
#32340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#32390000000
0$
0)
#32400000000
1"
1'
b0 +
b0 1
#32450000000
0"
0'
#32460000000
1#
1(
b101111101100100 +
b101111101100100 1
#32510000000
0#
0(
#32520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#32570000000
0$
0)
#32580000000
1"
1'
b0 +
b0 1
#32630000000
0"
0'
#32640000000
1#
1(
b101111101100100 +
b101111101100100 1
#32690000000
0#
0(
#32700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#32750000000
0$
0)
#32760000000
1"
1'
b0 +
b0 1
#32810000000
0"
0'
#32820000000
1#
1(
b101111101100100 +
b101111101100100 1
#32870000000
0#
0(
#32880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#32930000000
0$
0)
#32940000000
1"
1'
b0 +
b0 1
#32990000000
0"
0'
#33000000000
1#
1(
b101111101100100 +
b101111101100100 1
#33050000000
0#
0(
#33060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#33110000000
0$
0)
#33120000000
1"
1'
b0 +
b0 1
#33170000000
0"
0'
#33180000000
1#
1(
b101111101100100 +
b101111101100100 1
#33230000000
0#
0(
#33240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#33290000000
0$
0)
#33300000000
1"
1'
b0 +
b0 1
#33350000000
0"
0'
#33360000000
1#
1(
b101111101100100 +
b101111101100100 1
#33410000000
0#
0(
#33420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#33470000000
0$
0)
#33480000000
1"
1'
b0 +
b0 1
#33530000000
0"
0'
#33540000000
1#
1(
b101111101100100 +
b101111101100100 1
#33590000000
0#
0(
#33600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#33650000000
0$
0)
#33660000000
1"
1'
b0 +
b0 1
#33710000000
0"
0'
#33720000000
1#
1(
b101111101100100 +
b101111101100100 1
#33770000000
0#
0(
#33780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#33830000000
0$
0)
#33840000000
1"
1'
b0 +
b0 1
#33890000000
0"
0'
#33900000000
1#
1(
b101111101100100 +
b101111101100100 1
#33950000000
0#
0(
#33960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#34010000000
0$
0)
#34020000000
1"
1'
b0 +
b0 1
#34070000000
0"
0'
#34080000000
1#
1(
b101111101100100 +
b101111101100100 1
#34130000000
0#
0(
#34140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#34190000000
0$
0)
#34200000000
1"
1'
b0 +
b0 1
#34250000000
0"
0'
#34260000000
1#
1(
b101111101100100 +
b101111101100100 1
#34310000000
0#
0(
#34320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#34370000000
0$
0)
#34380000000
1"
1'
b0 +
b0 1
#34430000000
0"
0'
#34440000000
1#
1(
b101111101100100 +
b101111101100100 1
#34490000000
0#
0(
#34500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#34550000000
0$
0)
#34560000000
1"
1'
b0 +
b0 1
#34610000000
0"
0'
#34620000000
1#
1(
b101111101100100 +
b101111101100100 1
#34670000000
0#
0(
#34680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#34730000000
0$
0)
#34740000000
1"
1'
b0 +
b0 1
#34790000000
0"
0'
#34800000000
1#
1(
b101111101100100 +
b101111101100100 1
#34850000000
0#
0(
#34860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#34910000000
0$
0)
#34920000000
1"
1'
b0 +
b0 1
#34970000000
0"
0'
#34980000000
1#
1(
b101111101100100 +
b101111101100100 1
#35030000000
0#
0(
#35040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#35090000000
0$
0)
#35100000000
1"
1'
b0 +
b0 1
#35150000000
0"
0'
#35160000000
1#
1(
b101111101100100 +
b101111101100100 1
#35210000000
0#
0(
#35220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#35270000000
0$
0)
#35280000000
1"
1'
b0 +
b0 1
#35330000000
0"
0'
#35340000000
1#
1(
b101111101100100 +
b101111101100100 1
#35390000000
0#
0(
#35400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#35450000000
0$
0)
#35460000000
1"
1'
b0 +
b0 1
#35510000000
0"
0'
#35520000000
1#
1(
b101111101100100 +
b101111101100100 1
#35570000000
0#
0(
#35580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#35630000000
0$
0)
#35640000000
1"
1'
b0 +
b0 1
#35690000000
0"
0'
#35700000000
1#
1(
b101111101100100 +
b101111101100100 1
#35750000000
0#
0(
#35760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#35810000000
0$
0)
#35820000000
1"
1'
b0 +
b0 1
#35870000000
0"
0'
#35880000000
1#
1(
b101111101100100 +
b101111101100100 1
#35930000000
0#
0(
#35940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#35990000000
0$
0)
#36000000000
1"
1'
b0 +
b0 1
#36050000000
0"
0'
#36060000000
1#
1(
b101111101100100 +
b101111101100100 1
#36110000000
0#
0(
#36120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#36170000000
0$
0)
#36180000000
1"
1'
b0 +
b0 1
#36230000000
0"
0'
#36240000000
1#
1(
b101111101100100 +
b101111101100100 1
#36290000000
0#
0(
#36300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#36350000000
0$
0)
#36360000000
1"
1'
b0 +
b0 1
#36410000000
0"
0'
#36420000000
1#
1(
b101111101100100 +
b101111101100100 1
#36470000000
0#
0(
#36480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#36530000000
0$
0)
#36540000000
1"
1'
b0 +
b0 1
#36590000000
0"
0'
#36600000000
1#
1(
b101111101100100 +
b101111101100100 1
#36650000000
0#
0(
#36660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#36710000000
0$
0)
#36720000000
1"
1'
b0 +
b0 1
#36770000000
0"
0'
#36780000000
1#
1(
b101111101100100 +
b101111101100100 1
#36830000000
0#
0(
#36840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#36890000000
0$
0)
#36900000000
1"
1'
b0 +
b0 1
#36950000000
0"
0'
#36960000000
1#
1(
b101111101100100 +
b101111101100100 1
#37010000000
0#
0(
#37020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#37070000000
0$
0)
#37080000000
1"
1'
b0 +
b0 1
#37130000000
0"
0'
#37140000000
1#
1(
b101111101100100 +
b101111101100100 1
#37190000000
0#
0(
#37200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#37250000000
0$
0)
#37260000000
1"
1'
b0 +
b0 1
#37310000000
0"
0'
#37320000000
1#
1(
b101111101100100 +
b101111101100100 1
#37370000000
0#
0(
#37380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#37430000000
0$
0)
#37440000000
1"
1'
b0 +
b0 1
#37490000000
0"
0'
#37500000000
1#
1(
b101111101100100 +
b101111101100100 1
#37550000000
0#
0(
#37560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#37610000000
0$
0)
#37620000000
1"
1'
b0 +
b0 1
#37670000000
0"
0'
#37680000000
1#
1(
b101111101100100 +
b101111101100100 1
#37730000000
0#
0(
#37740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#37790000000
0$
0)
#37800000000
1"
1'
b0 +
b0 1
#37850000000
0"
0'
#37860000000
1#
1(
b101111101100100 +
b101111101100100 1
#37910000000
0#
0(
#37920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#37970000000
0$
0)
#37980000000
1"
1'
b0 +
b0 1
#38030000000
0"
0'
#38040000000
1#
1(
b101111101100100 +
b101111101100100 1
#38090000000
0#
0(
#38100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#38150000000
0$
0)
#38160000000
1"
1'
b0 +
b0 1
#38210000000
0"
0'
#38220000000
1#
1(
b101111101100100 +
b101111101100100 1
#38270000000
0#
0(
#38280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#38330000000
0$
0)
#38340000000
1"
1'
b0 +
b0 1
#38390000000
0"
0'
#38400000000
1#
1(
b101111101100100 +
b101111101100100 1
#38450000000
0#
0(
#38460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#38510000000
0$
0)
#38520000000
1"
1'
b0 +
b0 1
#38570000000
0"
0'
#38580000000
1#
1(
b101111101100100 +
b101111101100100 1
#38630000000
0#
0(
#38640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#38690000000
0$
0)
#38700000000
1"
1'
b0 +
b0 1
#38750000000
0"
0'
#38760000000
1#
1(
b101111101100100 +
b101111101100100 1
#38810000000
0#
0(
#38820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#38870000000
0$
0)
#38880000000
1"
1'
b0 +
b0 1
#38930000000
0"
0'
#38940000000
1#
1(
b101111101100100 +
b101111101100100 1
#38990000000
0#
0(
#39000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#39050000000
0$
0)
#39060000000
1"
1'
b0 +
b0 1
#39110000000
0"
0'
#39120000000
1#
1(
b101111101100100 +
b101111101100100 1
#39170000000
0#
0(
#39180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#39230000000
0$
0)
#39240000000
1"
1'
b0 +
b0 1
#39290000000
0"
0'
#39300000000
1#
1(
b101111101100100 +
b101111101100100 1
#39350000000
0#
0(
#39360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#39410000000
0$
0)
#39420000000
1"
1'
b0 +
b0 1
#39470000000
0"
0'
#39480000000
1#
1(
b101111101100100 +
b101111101100100 1
#39530000000
0#
0(
#39540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#39590000000
0$
0)
#39600000000
1"
1'
b0 +
b0 1
#39650000000
0"
0'
#39660000000
1#
1(
b101111101100100 +
b101111101100100 1
#39710000000
0#
0(
#39720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#39770000000
0$
0)
#39780000000
1"
1'
b0 +
b0 1
#39830000000
0"
0'
#39840000000
1#
1(
b101111101100100 +
b101111101100100 1
#39890000000
0#
0(
#39900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#39950000000
0$
0)
#39960000000
1"
1'
b0 +
b0 1
#40010000000
0"
0'
#40020000000
1#
1(
b101111101100100 +
b101111101100100 1
#40070000000
0#
0(
#40080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#40130000000
0$
0)
#40140000000
1"
1'
b0 +
b0 1
#40190000000
0"
0'
#40200000000
1#
1(
b101111101100100 +
b101111101100100 1
#40250000000
0#
0(
#40260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#40310000000
0$
0)
#40320000000
1"
1'
b0 +
b0 1
#40370000000
0"
0'
#40380000000
1#
1(
b101111101100100 +
b101111101100100 1
#40430000000
0#
0(
#40440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#40490000000
0$
0)
#40500000000
1"
1'
b0 +
b0 1
#40550000000
0"
0'
#40560000000
1#
1(
b101111101100100 +
b101111101100100 1
#40610000000
0#
0(
#40620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#40670000000
0$
0)
#40680000000
1"
1'
b0 +
b0 1
#40730000000
0"
0'
#40740000000
1#
1(
b101111101100100 +
b101111101100100 1
#40790000000
0#
0(
#40800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#40850000000
0$
0)
#40860000000
1"
1'
b0 +
b0 1
#40910000000
0"
0'
#40920000000
1#
1(
b101111101100100 +
b101111101100100 1
#40970000000
0#
0(
#40980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#41030000000
0$
0)
#41040000000
1"
1'
b0 +
b0 1
#41090000000
0"
0'
#41100000000
1#
1(
b101111101100100 +
b101111101100100 1
#41150000000
0#
0(
#41160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#41210000000
0$
0)
#41220000000
1"
1'
b0 +
b0 1
#41270000000
0"
0'
#41280000000
1#
1(
b101111101100100 +
b101111101100100 1
#41330000000
0#
0(
#41340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#41390000000
0$
0)
#41400000000
1"
1'
b0 +
b0 1
#41450000000
0"
0'
#41460000000
1#
1(
b101111101100100 +
b101111101100100 1
#41510000000
0#
0(
#41520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#41570000000
0$
0)
#41580000000
1"
1'
b0 +
b0 1
#41630000000
0"
0'
#41640000000
1#
1(
b101111101100100 +
b101111101100100 1
#41690000000
0#
0(
#41700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#41750000000
0$
0)
#41760000000
1"
1'
b0 +
b0 1
#41810000000
0"
0'
#41820000000
1#
1(
b101111101100100 +
b101111101100100 1
#41870000000
0#
0(
#41880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#41930000000
0$
0)
#41940000000
1"
1'
b0 +
b0 1
#41990000000
0"
0'
#42000000000
1#
1(
b101111101100100 +
b101111101100100 1
#42050000000
0#
0(
#42060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#42110000000
0$
0)
#42120000000
1"
1'
b0 +
b0 1
#42170000000
0"
0'
#42180000000
1#
1(
b101111101100100 +
b101111101100100 1
#42230000000
0#
0(
#42240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#42290000000
0$
0)
#42300000000
1"
1'
b0 +
b0 1
#42350000000
0"
0'
#42360000000
1#
1(
b101111101100100 +
b101111101100100 1
#42410000000
0#
0(
#42420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#42470000000
0$
0)
#42480000000
1"
1'
b0 +
b0 1
#42530000000
0"
0'
#42540000000
1#
1(
b101111101100100 +
b101111101100100 1
#42590000000
0#
0(
#42600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#42650000000
0$
0)
#42660000000
1"
1'
b0 +
b0 1
#42710000000
0"
0'
#42720000000
1#
1(
b101111101100100 +
b101111101100100 1
#42770000000
0#
0(
#42780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#42830000000
0$
0)
#42840000000
1"
1'
b0 +
b0 1
#42890000000
0"
0'
#42900000000
1#
1(
b101111101100100 +
b101111101100100 1
#42950000000
0#
0(
#42960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#43010000000
0$
0)
#43020000000
1"
1'
b0 +
b0 1
#43070000000
0"
0'
#43080000000
1#
1(
b101111101100100 +
b101111101100100 1
#43130000000
0#
0(
#43140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#43190000000
0$
0)
#43200000000
1"
1'
b0 +
b0 1
#43250000000
0"
0'
#43260000000
1#
1(
b101111101100100 +
b101111101100100 1
#43310000000
0#
0(
#43320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#43370000000
0$
0)
#43380000000
1"
1'
b0 +
b0 1
#43430000000
0"
0'
#43440000000
1#
1(
b101111101100100 +
b101111101100100 1
#43490000000
0#
0(
#43500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#43550000000
0$
0)
#43560000000
1"
1'
b0 +
b0 1
#43610000000
0"
0'
#43620000000
1#
1(
b101111101100100 +
b101111101100100 1
#43670000000
0#
0(
#43680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#43730000000
0$
0)
#43740000000
1"
1'
b0 +
b0 1
#43790000000
0"
0'
#43800000000
1#
1(
b101111101100100 +
b101111101100100 1
#43850000000
0#
0(
#43860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#43910000000
0$
0)
#43920000000
1"
1'
b0 +
b0 1
#43970000000
0"
0'
#43980000000
1#
1(
b101111101100100 +
b101111101100100 1
#44030000000
0#
0(
#44040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#44090000000
0$
0)
#44100000000
1"
1'
b0 +
b0 1
#44150000000
0"
0'
#44160000000
1#
1(
b101111101100100 +
b101111101100100 1
#44210000000
0#
0(
#44220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#44270000000
0$
0)
#44280000000
1"
1'
b0 +
b0 1
#44330000000
0"
0'
#44340000000
1#
1(
b101111101100100 +
b101111101100100 1
#44390000000
0#
0(
#44400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#44450000000
0$
0)
#44460000000
1"
1'
b0 +
b0 1
#44510000000
0"
0'
#44520000000
1#
1(
b101111101100100 +
b101111101100100 1
#44570000000
0#
0(
#44580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#44630000000
0$
0)
#44640000000
1"
1'
b0 +
b0 1
#44690000000
0"
0'
#44700000000
1#
1(
b101111101100100 +
b101111101100100 1
#44750000000
0#
0(
#44760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#44810000000
0$
0)
#44820000000
1"
1'
b0 +
b0 1
#44870000000
0"
0'
#44880000000
1#
1(
b101111101100100 +
b101111101100100 1
#44930000000
0#
0(
#44940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#44990000000
0$
0)
#45000000000
1"
1'
b0 +
b0 1
#45050000000
0"
0'
#45060000000
1#
1(
b101111101100100 +
b101111101100100 1
#45110000000
0#
0(
#45120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#45170000000
0$
0)
#45180000000
1"
1'
b0 +
b0 1
#45230000000
0"
0'
#45240000000
1#
1(
b101111101100100 +
b101111101100100 1
#45290000000
0#
0(
#45300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#45350000000
0$
0)
#45360000000
1"
1'
b0 +
b0 1
#45410000000
0"
0'
#45420000000
1#
1(
b101111101100100 +
b101111101100100 1
#45470000000
0#
0(
#45480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#45530000000
0$
0)
#45540000000
1"
1'
b0 +
b0 1
#45590000000
0"
0'
#45600000000
1#
1(
b101111101100100 +
b101111101100100 1
#45650000000
0#
0(
#45660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#45710000000
0$
0)
#45720000000
1"
1'
b0 +
b0 1
#45770000000
0"
0'
#45780000000
1#
1(
b101111101100100 +
b101111101100100 1
#45830000000
0#
0(
#45840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#45890000000
0$
0)
#45900000000
1"
1'
b0 +
b0 1
#45950000000
0"
0'
#45960000000
1#
1(
b101111101100100 +
b101111101100100 1
#46010000000
0#
0(
#46020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#46070000000
0$
0)
#46080000000
1"
1'
b0 +
b0 1
#46130000000
0"
0'
#46140000000
1#
1(
b101111101100100 +
b101111101100100 1
#46190000000
0#
0(
#46200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#46250000000
0$
0)
#46260000000
1"
1'
b0 +
b0 1
#46310000000
0"
0'
#46320000000
1#
1(
b101111101100100 +
b101111101100100 1
#46370000000
0#
0(
#46380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#46430000000
0$
0)
#46440000000
1"
1'
b0 +
b0 1
#46490000000
0"
0'
#46500000000
1#
1(
b101111101100100 +
b101111101100100 1
#46550000000
0#
0(
#46560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#46610000000
0$
0)
#46620000000
1"
1'
b0 +
b0 1
#46670000000
0"
0'
#46680000000
1#
1(
b101111101100100 +
b101111101100100 1
#46730000000
0#
0(
#46740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#46790000000
0$
0)
#46800000000
1"
1'
b0 +
b0 1
#46850000000
0"
0'
#46860000000
1#
1(
b101111101100100 +
b101111101100100 1
#46910000000
0#
0(
#46920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#46970000000
0$
0)
#46980000000
1"
1'
b0 +
b0 1
#47030000000
0"
0'
#47040000000
1#
1(
b101111101100100 +
b101111101100100 1
#47090000000
0#
0(
#47100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#47150000000
0$
0)
#47160000000
1"
1'
b0 +
b0 1
#47210000000
0"
0'
#47220000000
1#
1(
b101111101100100 +
b101111101100100 1
#47270000000
0#
0(
#47280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#47330000000
0$
0)
#47340000000
1"
1'
b0 +
b0 1
#47390000000
0"
0'
#47400000000
1#
1(
b101111101100100 +
b101111101100100 1
#47450000000
0#
0(
#47460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#47510000000
0$
0)
#47520000000
1"
1'
b0 +
b0 1
#47570000000
0"
0'
#47580000000
1#
1(
b101111101100100 +
b101111101100100 1
#47630000000
0#
0(
#47640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#47690000000
0$
0)
#47700000000
1"
1'
b0 +
b0 1
#47750000000
0"
0'
#47760000000
1#
1(
b101111101100100 +
b101111101100100 1
#47810000000
0#
0(
#47820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#47870000000
0$
0)
#47880000000
1"
1'
b0 +
b0 1
#47930000000
0"
0'
#47940000000
1#
1(
b101111101100100 +
b101111101100100 1
#47990000000
0#
0(
#48000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#48050000000
0$
0)
#48060000000
1"
1'
b0 +
b0 1
#48110000000
0"
0'
#48120000000
1#
1(
b101111101100100 +
b101111101100100 1
#48170000000
0#
0(
#48180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#48230000000
0$
0)
#48240000000
1"
1'
b0 +
b0 1
#48290000000
0"
0'
#48300000000
1#
1(
b101111101100100 +
b101111101100100 1
#48350000000
0#
0(
#48360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#48410000000
0$
0)
#48420000000
1"
1'
b0 +
b0 1
#48470000000
0"
0'
#48480000000
1#
1(
b101111101100100 +
b101111101100100 1
#48530000000
0#
0(
#48540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#48590000000
0$
0)
#48600000000
1"
1'
b0 +
b0 1
#48650000000
0"
0'
#48660000000
1#
1(
b101111101100100 +
b101111101100100 1
#48710000000
0#
0(
#48720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#48770000000
0$
0)
#48780000000
1"
1'
b0 +
b0 1
#48830000000
0"
0'
#48840000000
1#
1(
b101111101100100 +
b101111101100100 1
#48890000000
0#
0(
#48900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#48950000000
0$
0)
#48960000000
1"
1'
b0 +
b0 1
#49010000000
0"
0'
#49020000000
1#
1(
b101111101100100 +
b101111101100100 1
#49070000000
0#
0(
#49080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#49130000000
0$
0)
#49140000000
1"
1'
b0 +
b0 1
#49190000000
0"
0'
#49200000000
1#
1(
b101111101100100 +
b101111101100100 1
#49250000000
0#
0(
#49260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#49310000000
0$
0)
#49320000000
1"
1'
b0 +
b0 1
#49370000000
0"
0'
#49380000000
1#
1(
b101111101100100 +
b101111101100100 1
#49430000000
0#
0(
#49440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#49490000000
0$
0)
#49500000000
1"
1'
b0 +
b0 1
#49550000000
0"
0'
#49560000000
1#
1(
b101111101100100 +
b101111101100100 1
#49610000000
0#
0(
#49620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#49670000000
0$
0)
#49680000000
1"
1'
b0 +
b0 1
#49730000000
0"
0'
#49740000000
1#
1(
b101111101100100 +
b101111101100100 1
#49790000000
0#
0(
#49800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#49850000000
0$
0)
#49860000000
1"
1'
b0 +
b0 1
#49910000000
0"
0'
#49920000000
1#
1(
b101111101100100 +
b101111101100100 1
#49970000000
0#
0(
#49980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#50030000000
0$
0)
#50040000000
1"
1'
b0 +
b0 1
#50090000000
0"
0'
#50100000000
1#
1(
b101111101100100 +
b101111101100100 1
#50150000000
0#
0(
#50160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#50210000000
0$
0)
#50220000000
1"
1'
b0 +
b0 1
#50270000000
0"
0'
#50280000000
1#
1(
b101111101100100 +
b101111101100100 1
#50330000000
0#
0(
#50340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#50390000000
0$
0)
#50400000000
1"
1'
b0 +
b0 1
#50450000000
0"
0'
#50460000000
1#
1(
b101111101100100 +
b101111101100100 1
#50510000000
0#
0(
#50520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#50570000000
0$
0)
#50580000000
1"
1'
b0 +
b0 1
#50630000000
0"
0'
#50640000000
1#
1(
b101111101100100 +
b101111101100100 1
#50690000000
0#
0(
#50700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#50750000000
0$
0)
#50760000000
1"
1'
b0 +
b0 1
#50810000000
0"
0'
#50820000000
1#
1(
b101111101100100 +
b101111101100100 1
#50870000000
0#
0(
#50880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#50930000000
0$
0)
#50940000000
1"
1'
b0 +
b0 1
#50990000000
0"
0'
#51000000000
1#
1(
b101111101100100 +
b101111101100100 1
#51050000000
0#
0(
#51060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#51110000000
0$
0)
#51120000000
1"
1'
b0 +
b0 1
#51170000000
0"
0'
#51180000000
1#
1(
b101111101100100 +
b101111101100100 1
#51230000000
0#
0(
#51240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#51290000000
0$
0)
#51300000000
1"
1'
b0 +
b0 1
#51350000000
0"
0'
#51360000000
1#
1(
b101111101100100 +
b101111101100100 1
#51410000000
0#
0(
#51420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#51470000000
0$
0)
#51480000000
1"
1'
b0 +
b0 1
#51530000000
0"
0'
#51540000000
1#
1(
b101111101100100 +
b101111101100100 1
#51590000000
0#
0(
#51600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#51650000000
0$
0)
#51660000000
1"
1'
b0 +
b0 1
#51710000000
0"
0'
#51720000000
1#
1(
b101111101100100 +
b101111101100100 1
#51770000000
0#
0(
#51780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#51830000000
0$
0)
#51840000000
1"
1'
b0 +
b0 1
#51890000000
0"
0'
#51900000000
1#
1(
b101111101100100 +
b101111101100100 1
#51950000000
0#
0(
#51960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#52010000000
0$
0)
#52020000000
1"
1'
b0 +
b0 1
#52070000000
0"
0'
#52080000000
1#
1(
b101111101100100 +
b101111101100100 1
#52130000000
0#
0(
#52140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#52190000000
0$
0)
#52200000000
1"
1'
b0 +
b0 1
#52250000000
0"
0'
#52260000000
1#
1(
b101111101100100 +
b101111101100100 1
#52310000000
0#
0(
#52320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#52370000000
0$
0)
#52380000000
1"
1'
b0 +
b0 1
#52430000000
0"
0'
#52440000000
1#
1(
b101111101100100 +
b101111101100100 1
#52490000000
0#
0(
#52500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#52550000000
0$
0)
#52560000000
1"
1'
b0 +
b0 1
#52610000000
0"
0'
#52620000000
1#
1(
b101111101100100 +
b101111101100100 1
#52670000000
0#
0(
#52680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#52730000000
0$
0)
#52740000000
1"
1'
b0 +
b0 1
#52790000000
0"
0'
#52800000000
1#
1(
b101111101100100 +
b101111101100100 1
#52850000000
0#
0(
#52860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#52910000000
0$
0)
#52920000000
1"
1'
b0 +
b0 1
#52970000000
0"
0'
#52980000000
1#
1(
b101111101100100 +
b101111101100100 1
#53030000000
0#
0(
#53040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#53090000000
0$
0)
#53100000000
1"
1'
b0 +
b0 1
#53150000000
0"
0'
#53160000000
1#
1(
b101111101100100 +
b101111101100100 1
#53210000000
0#
0(
#53220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#53270000000
0$
0)
#53280000000
1"
1'
b0 +
b0 1
#53330000000
0"
0'
#53340000000
1#
1(
b101111101100100 +
b101111101100100 1
#53390000000
0#
0(
#53400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#53450000000
0$
0)
#53460000000
1"
1'
b0 +
b0 1
#53510000000
0"
0'
#53520000000
1#
1(
b101111101100100 +
b101111101100100 1
#53570000000
0#
0(
#53580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#53630000000
0$
0)
#53640000000
1"
1'
b0 +
b0 1
#53690000000
0"
0'
#53700000000
1#
1(
b101111101100100 +
b101111101100100 1
#53750000000
0#
0(
#53760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#53810000000
0$
0)
#53820000000
1"
1'
b0 +
b0 1
#53870000000
0"
0'
#53880000000
1#
1(
b101111101100100 +
b101111101100100 1
#53930000000
0#
0(
#53940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#53990000000
0$
0)
#54000000000
1"
1'
b0 +
b0 1
#54050000000
0"
0'
#54060000000
1#
1(
b101111101100100 +
b101111101100100 1
#54110000000
0#
0(
#54120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#54170000000
0$
0)
#54180000000
1"
1'
b0 +
b0 1
#54230000000
0"
0'
#54240000000
1#
1(
b101111101100100 +
b101111101100100 1
#54290000000
0#
0(
#54300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#54350000000
0$
0)
#54360000000
1"
1'
b0 +
b0 1
#54410000000
0"
0'
#54420000000
1#
1(
b101111101100100 +
b101111101100100 1
#54470000000
0#
0(
#54480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#54530000000
0$
0)
#54540000000
1"
1'
b0 +
b0 1
#54590000000
0"
0'
#54600000000
1#
1(
b101111101100100 +
b101111101100100 1
#54650000000
0#
0(
#54660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#54710000000
0$
0)
#54720000000
1"
1'
b0 +
b0 1
#54770000000
0"
0'
#54780000000
1#
1(
b101111101100100 +
b101111101100100 1
#54830000000
0#
0(
#54840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#54890000000
0$
0)
#54900000000
1"
1'
b0 +
b0 1
#54950000000
0"
0'
#54960000000
1#
1(
b101111101100100 +
b101111101100100 1
#55010000000
0#
0(
#55020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#55070000000
0$
0)
#55080000000
1"
1'
b0 +
b0 1
#55130000000
0"
0'
#55140000000
1#
1(
b101111101100100 +
b101111101100100 1
#55190000000
0#
0(
#55200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#55250000000
0$
0)
#55260000000
1"
1'
b0 +
b0 1
#55310000000
0"
0'
#55320000000
1#
1(
b101111101100100 +
b101111101100100 1
#55370000000
0#
0(
#55380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#55430000000
0$
0)
#55440000000
1"
1'
b0 +
b0 1
#55490000000
0"
0'
#55500000000
1#
1(
b101111101100100 +
b101111101100100 1
#55550000000
0#
0(
#55560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#55610000000
0$
0)
#55620000000
1"
1'
b0 +
b0 1
#55670000000
0"
0'
#55680000000
1#
1(
b101111101100100 +
b101111101100100 1
#55730000000
0#
0(
#55740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#55790000000
0$
0)
#55800000000
1"
1'
b0 +
b0 1
#55850000000
0"
0'
#55860000000
1#
1(
b101111101100100 +
b101111101100100 1
#55910000000
0#
0(
#55920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#55970000000
0$
0)
#55980000000
1"
1'
b0 +
b0 1
#56030000000
0"
0'
#56040000000
1#
1(
b101111101100100 +
b101111101100100 1
#56090000000
0#
0(
#56100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#56150000000
0$
0)
#56160000000
1"
1'
b0 +
b0 1
#56210000000
0"
0'
#56220000000
1#
1(
b101111101100100 +
b101111101100100 1
#56270000000
0#
0(
#56280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#56330000000
0$
0)
#56340000000
1"
1'
b0 +
b0 1
#56390000000
0"
0'
#56400000000
1#
1(
b101111101100100 +
b101111101100100 1
#56450000000
0#
0(
#56460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#56510000000
0$
0)
#56520000000
1"
1'
b0 +
b0 1
#56570000000
0"
0'
#56580000000
1#
1(
b101111101100100 +
b101111101100100 1
#56630000000
0#
0(
#56640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#56690000000
0$
0)
#56700000000
1"
1'
b0 +
b0 1
#56750000000
0"
0'
#56760000000
1#
1(
b101111101100100 +
b101111101100100 1
#56810000000
0#
0(
#56820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#56870000000
0$
0)
#56880000000
1"
1'
b0 +
b0 1
#56930000000
0"
0'
#56940000000
1#
1(
b101111101100100 +
b101111101100100 1
#56990000000
0#
0(
#57000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#57050000000
0$
0)
#57060000000
1"
1'
b0 +
b0 1
#57110000000
0"
0'
#57120000000
1#
1(
b101111101100100 +
b101111101100100 1
#57170000000
0#
0(
#57180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#57230000000
0$
0)
#57240000000
1"
1'
b0 +
b0 1
#57290000000
0"
0'
#57300000000
1#
1(
b101111101100100 +
b101111101100100 1
#57350000000
0#
0(
#57360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#57410000000
0$
0)
#57420000000
1"
1'
b0 +
b0 1
#57470000000
0"
0'
#57480000000
1#
1(
b101111101100100 +
b101111101100100 1
#57530000000
0#
0(
#57540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#57590000000
0$
0)
#57600000000
1"
1'
b0 +
b0 1
#57650000000
0"
0'
#57660000000
1#
1(
b101111101100100 +
b101111101100100 1
#57710000000
0#
0(
#57720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#57770000000
0$
0)
#57780000000
1"
1'
b0 +
b0 1
#57830000000
0"
0'
#57840000000
1#
1(
b101111101100100 +
b101111101100100 1
#57890000000
0#
0(
#57900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#57950000000
0$
0)
#57960000000
1"
1'
b0 +
b0 1
#58010000000
0"
0'
#58020000000
1#
1(
b101111101100100 +
b101111101100100 1
#58070000000
0#
0(
#58080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#58130000000
0$
0)
#58140000000
1"
1'
b0 +
b0 1
#58190000000
0"
0'
#58200000000
1#
1(
b101111101100100 +
b101111101100100 1
#58250000000
0#
0(
#58260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#58310000000
0$
0)
#58320000000
1"
1'
b0 +
b0 1
#58370000000
0"
0'
#58380000000
1#
1(
b101111101100100 +
b101111101100100 1
#58430000000
0#
0(
#58440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#58490000000
0$
0)
#58500000000
1"
1'
b0 +
b0 1
#58550000000
0"
0'
#58560000000
1#
1(
b101111101100100 +
b101111101100100 1
#58610000000
0#
0(
#58620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#58670000000
0$
0)
#58680000000
1"
1'
b0 +
b0 1
#58730000000
0"
0'
#58740000000
1#
1(
b101111101100100 +
b101111101100100 1
#58790000000
0#
0(
#58800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#58850000000
0$
0)
#58860000000
1"
1'
b0 +
b0 1
#58910000000
0"
0'
#58920000000
1#
1(
b101111101100100 +
b101111101100100 1
#58970000000
0#
0(
#58980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#59030000000
0$
0)
#59040000000
1"
1'
b0 +
b0 1
#59090000000
0"
0'
#59100000000
1#
1(
b101111101100100 +
b101111101100100 1
#59150000000
0#
0(
#59160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#59210000000
0$
0)
#59220000000
1"
1'
b0 +
b0 1
#59270000000
0"
0'
#59280000000
1#
1(
b101111101100100 +
b101111101100100 1
#59330000000
0#
0(
#59340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#59390000000
0$
0)
#59400000000
1"
1'
b0 +
b0 1
#59450000000
0"
0'
#59460000000
1#
1(
b101111101100100 +
b101111101100100 1
#59510000000
0#
0(
#59520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#59570000000
0$
0)
#59580000000
1"
1'
b0 +
b0 1
#59630000000
0"
0'
#59640000000
1#
1(
b101111101100100 +
b101111101100100 1
#59690000000
0#
0(
#59700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#59750000000
0$
0)
#59760000000
1"
1'
b0 +
b0 1
#59810000000
0"
0'
#59820000000
1#
1(
b101111101100100 +
b101111101100100 1
#59870000000
0#
0(
#59880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#59930000000
0$
0)
#59940000000
1"
1'
b0 +
b0 1
#59990000000
0"
0'
#60000000000
1#
1(
b101111101100100 +
b101111101100100 1
#60050000000
0#
0(
#60060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#60110000000
0$
0)
#60120000000
1"
1'
b0 +
b0 1
#60170000000
0"
0'
#60180000000
1#
1(
b101111101100100 +
b101111101100100 1
#60230000000
0#
0(
#60240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#60290000000
0$
0)
#60300000000
1"
1'
b0 +
b0 1
#60350000000
0"
0'
#60360000000
1#
1(
b101111101100100 +
b101111101100100 1
#60410000000
0#
0(
#60420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#60470000000
0$
0)
#60480000000
1"
1'
b0 +
b0 1
#60530000000
0"
0'
#60540000000
1#
1(
b101111101100100 +
b101111101100100 1
#60590000000
0#
0(
#60600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#60650000000
0$
0)
#60660000000
1"
1'
b0 +
b0 1
#60710000000
0"
0'
#60720000000
1#
1(
b101111101100100 +
b101111101100100 1
#60770000000
0#
0(
#60780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#60830000000
0$
0)
#60840000000
1"
1'
b0 +
b0 1
#60890000000
0"
0'
#60900000000
1#
1(
b101111101100100 +
b101111101100100 1
#60950000000
0#
0(
#60960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#61010000000
0$
0)
#61020000000
1"
1'
b0 +
b0 1
#61070000000
0"
0'
#61080000000
1#
1(
b101111101100100 +
b101111101100100 1
#61130000000
0#
0(
#61140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#61190000000
0$
0)
#61200000000
1"
1'
b0 +
b0 1
#61250000000
0"
0'
#61260000000
1#
1(
b101111101100100 +
b101111101100100 1
#61310000000
0#
0(
#61320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#61370000000
0$
0)
#61380000000
1"
1'
b0 +
b0 1
#61430000000
0"
0'
#61440000000
1#
1(
b101111101100100 +
b101111101100100 1
#61490000000
0#
0(
#61500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#61550000000
0$
0)
#61560000000
1"
1'
b0 +
b0 1
#61610000000
0"
0'
#61620000000
1#
1(
b101111101100100 +
b101111101100100 1
#61670000000
0#
0(
#61680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#61730000000
0$
0)
#61740000000
1"
1'
b0 +
b0 1
#61790000000
0"
0'
#61800000000
1#
1(
b101111101100100 +
b101111101100100 1
#61850000000
0#
0(
#61860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#61910000000
0$
0)
#61920000000
1"
1'
b0 +
b0 1
#61970000000
0"
0'
#61980000000
1#
1(
b101111101100100 +
b101111101100100 1
#62030000000
0#
0(
#62040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#62090000000
0$
0)
#62100000000
1"
1'
b0 +
b0 1
#62150000000
0"
0'
#62160000000
1#
1(
b101111101100100 +
b101111101100100 1
#62210000000
0#
0(
#62220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#62270000000
0$
0)
#62280000000
1"
1'
b0 +
b0 1
#62330000000
0"
0'
#62340000000
1#
1(
b101111101100100 +
b101111101100100 1
#62390000000
0#
0(
#62400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#62450000000
0$
0)
#62460000000
1"
1'
b0 +
b0 1
#62510000000
0"
0'
#62520000000
1#
1(
b101111101100100 +
b101111101100100 1
#62570000000
0#
0(
#62580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#62630000000
0$
0)
#62640000000
1"
1'
b0 +
b0 1
#62690000000
0"
0'
#62700000000
1#
1(
b101111101100100 +
b101111101100100 1
#62750000000
0#
0(
#62760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#62810000000
0$
0)
#62820000000
1"
1'
b0 +
b0 1
#62870000000
0"
0'
#62880000000
1#
1(
b101111101100100 +
b101111101100100 1
#62930000000
0#
0(
#62940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#62990000000
0$
0)
#63000000000
1"
1'
b0 +
b0 1
#63050000000
0"
0'
#63060000000
1#
1(
b101111101100100 +
b101111101100100 1
#63110000000
0#
0(
#63120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#63170000000
0$
0)
#63180000000
1"
1'
b0 +
b0 1
#63230000000
0"
0'
#63240000000
1#
1(
b101111101100100 +
b101111101100100 1
#63290000000
0#
0(
#63300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#63350000000
0$
0)
#63360000000
1"
1'
b0 +
b0 1
#63410000000
0"
0'
#63420000000
1#
1(
b101111101100100 +
b101111101100100 1
#63470000000
0#
0(
#63480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#63530000000
0$
0)
#63540000000
1"
1'
b0 +
b0 1
#63590000000
0"
0'
#63600000000
1#
1(
b101111101100100 +
b101111101100100 1
#63650000000
0#
0(
#63660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#63710000000
0$
0)
#63720000000
1"
1'
b0 +
b0 1
#63770000000
0"
0'
#63780000000
1#
1(
b101111101100100 +
b101111101100100 1
#63830000000
0#
0(
#63840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#63890000000
0$
0)
#63900000000
1"
1'
b0 +
b0 1
#63950000000
0"
0'
#63960000000
1#
1(
b101111101100100 +
b101111101100100 1
#64010000000
0#
0(
#64020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#64070000000
0$
0)
#64080000000
1"
1'
b0 +
b0 1
#64130000000
0"
0'
#64140000000
1#
1(
b101111101100100 +
b101111101100100 1
#64190000000
0#
0(
#64200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#64250000000
0$
0)
#64260000000
1"
1'
b0 +
b0 1
#64310000000
0"
0'
#64320000000
1#
1(
b101111101100100 +
b101111101100100 1
#64370000000
0#
0(
#64380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#64430000000
0$
0)
#64440000000
1"
1'
b0 +
b0 1
#64490000000
0"
0'
#64500000000
1#
1(
b101111101100100 +
b101111101100100 1
#64550000000
0#
0(
#64560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#64610000000
0$
0)
#64620000000
1"
1'
b0 +
b0 1
#64670000000
0"
0'
#64680000000
1#
1(
b101111101100100 +
b101111101100100 1
#64730000000
0#
0(
#64740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#64790000000
0$
0)
#64800000000
1"
1'
b0 +
b0 1
#64850000000
0"
0'
#64860000000
1#
1(
b101111101100100 +
b101111101100100 1
#64910000000
0#
0(
#64920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#64970000000
0$
0)
#64980000000
1"
1'
b0 +
b0 1
#65030000000
0"
0'
#65040000000
1#
1(
b101111101100100 +
b101111101100100 1
#65090000000
0#
0(
#65100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#65150000000
0$
0)
#65160000000
1"
1'
b0 +
b0 1
#65210000000
0"
0'
#65220000000
1#
1(
b101111101100100 +
b101111101100100 1
#65270000000
0#
0(
#65280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#65330000000
0$
0)
#65340000000
1"
1'
b0 +
b0 1
#65390000000
0"
0'
#65400000000
1#
1(
b101111101100100 +
b101111101100100 1
#65450000000
0#
0(
#65460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#65510000000
0$
0)
#65520000000
1"
1'
b0 +
b0 1
#65570000000
0"
0'
#65580000000
1#
1(
b101111101100100 +
b101111101100100 1
#65630000000
0#
0(
#65640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#65690000000
0$
0)
#65700000000
1"
1'
b0 +
b0 1
#65750000000
0"
0'
#65760000000
1#
1(
b101111101100100 +
b101111101100100 1
#65810000000
0#
0(
#65820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#65870000000
0$
0)
#65880000000
1"
1'
b0 +
b0 1
#65930000000
0"
0'
#65940000000
1#
1(
b101111101100100 +
b101111101100100 1
#65990000000
0#
0(
#66000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#66050000000
0$
0)
#66060000000
1"
1'
b0 +
b0 1
#66110000000
0"
0'
#66120000000
1#
1(
b101111101100100 +
b101111101100100 1
#66170000000
0#
0(
#66180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#66230000000
0$
0)
#66240000000
1"
1'
b0 +
b0 1
#66290000000
0"
0'
#66300000000
1#
1(
b101111101100100 +
b101111101100100 1
#66350000000
0#
0(
#66360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#66410000000
0$
0)
#66420000000
1"
1'
b0 +
b0 1
#66470000000
0"
0'
#66480000000
1#
1(
b101111101100100 +
b101111101100100 1
#66530000000
0#
0(
#66540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#66590000000
0$
0)
#66600000000
1"
1'
b0 +
b0 1
#66650000000
0"
0'
#66660000000
1#
1(
b101111101100100 +
b101111101100100 1
#66710000000
0#
0(
#66720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#66770000000
0$
0)
#66780000000
1"
1'
b0 +
b0 1
#66830000000
0"
0'
#66840000000
1#
1(
b101111101100100 +
b101111101100100 1
#66890000000
0#
0(
#66900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#66950000000
0$
0)
#66960000000
1"
1'
b0 +
b0 1
#67010000000
0"
0'
#67020000000
1#
1(
b101111101100100 +
b101111101100100 1
#67070000000
0#
0(
#67080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#67130000000
0$
0)
#67140000000
1"
1'
b0 +
b0 1
#67190000000
0"
0'
#67200000000
1#
1(
b101111101100100 +
b101111101100100 1
#67250000000
0#
0(
#67260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#67310000000
0$
0)
#67320000000
1"
1'
b0 +
b0 1
#67370000000
0"
0'
#67380000000
1#
1(
b101111101100100 +
b101111101100100 1
#67430000000
0#
0(
#67440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#67490000000
0$
0)
#67500000000
1"
1'
b0 +
b0 1
#67550000000
0"
0'
#67560000000
1#
1(
b101111101100100 +
b101111101100100 1
#67610000000
0#
0(
#67620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#67670000000
0$
0)
#67680000000
1"
1'
b0 +
b0 1
#67730000000
0"
0'
#67740000000
1#
1(
b101111101100100 +
b101111101100100 1
#67790000000
0#
0(
#67800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#67850000000
0$
0)
#67860000000
1"
1'
b0 +
b0 1
#67910000000
0"
0'
#67920000000
1#
1(
b101111101100100 +
b101111101100100 1
#67970000000
0#
0(
#67980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#68030000000
0$
0)
#68040000000
1"
1'
b0 +
b0 1
#68090000000
0"
0'
#68100000000
1#
1(
b101111101100100 +
b101111101100100 1
#68150000000
0#
0(
#68160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#68210000000
0$
0)
#68220000000
1"
1'
b0 +
b0 1
#68270000000
0"
0'
#68280000000
1#
1(
b101111101100100 +
b101111101100100 1
#68330000000
0#
0(
#68340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#68390000000
0$
0)
#68400000000
1"
1'
b0 +
b0 1
#68450000000
0"
0'
#68460000000
1#
1(
b101111101100100 +
b101111101100100 1
#68510000000
0#
0(
#68520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#68570000000
0$
0)
#68580000000
1"
1'
b0 +
b0 1
#68630000000
0"
0'
#68640000000
1#
1(
b101111101100100 +
b101111101100100 1
#68690000000
0#
0(
#68700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#68750000000
0$
0)
#68760000000
1"
1'
b0 +
b0 1
#68810000000
0"
0'
#68820000000
1#
1(
b101111101100100 +
b101111101100100 1
#68870000000
0#
0(
#68880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#68930000000
0$
0)
#68940000000
1"
1'
b0 +
b0 1
#68990000000
0"
0'
#69000000000
1#
1(
b101111101100100 +
b101111101100100 1
#69050000000
0#
0(
#69060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#69110000000
0$
0)
#69120000000
1"
1'
b0 +
b0 1
#69170000000
0"
0'
#69180000000
1#
1(
b101111101100100 +
b101111101100100 1
#69230000000
0#
0(
#69240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#69290000000
0$
0)
#69300000000
1"
1'
b0 +
b0 1
#69350000000
0"
0'
#69360000000
1#
1(
b101111101100100 +
b101111101100100 1
#69410000000
0#
0(
#69420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#69470000000
0$
0)
#69480000000
1"
1'
b0 +
b0 1
#69530000000
0"
0'
#69540000000
1#
1(
b101111101100100 +
b101111101100100 1
#69590000000
0#
0(
#69600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#69650000000
0$
0)
#69660000000
1"
1'
b0 +
b0 1
#69710000000
0"
0'
#69720000000
1#
1(
b101111101100100 +
b101111101100100 1
#69770000000
0#
0(
#69780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#69830000000
0$
0)
#69840000000
1"
1'
b0 +
b0 1
#69890000000
0"
0'
#69900000000
1#
1(
b101111101100100 +
b101111101100100 1
#69950000000
0#
0(
#69960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#70010000000
0$
0)
#70020000000
1"
1'
b0 +
b0 1
#70070000000
0"
0'
#70080000000
1#
1(
b101111101100100 +
b101111101100100 1
#70130000000
0#
0(
#70140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#70190000000
0$
0)
#70200000000
1"
1'
b0 +
b0 1
#70250000000
0"
0'
#70260000000
1#
1(
b101111101100100 +
b101111101100100 1
#70310000000
0#
0(
#70320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#70370000000
0$
0)
#70380000000
1"
1'
b0 +
b0 1
#70430000000
0"
0'
#70440000000
1#
1(
b101111101100100 +
b101111101100100 1
#70490000000
0#
0(
#70500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#70550000000
0$
0)
#70560000000
1"
1'
b0 +
b0 1
#70610000000
0"
0'
#70620000000
1#
1(
b101111101100100 +
b101111101100100 1
#70670000000
0#
0(
#70680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#70730000000
0$
0)
#70740000000
1"
1'
b0 +
b0 1
#70790000000
0"
0'
#70800000000
1#
1(
b101111101100100 +
b101111101100100 1
#70850000000
0#
0(
#70860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#70910000000
0$
0)
#70920000000
1"
1'
b0 +
b0 1
#70970000000
0"
0'
#70980000000
1#
1(
b101111101100100 +
b101111101100100 1
#71030000000
0#
0(
#71040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#71090000000
0$
0)
#71100000000
1"
1'
b0 +
b0 1
#71150000000
0"
0'
#71160000000
1#
1(
b101111101100100 +
b101111101100100 1
#71210000000
0#
0(
#71220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#71270000000
0$
0)
#71280000000
1"
1'
b0 +
b0 1
#71330000000
0"
0'
#71340000000
1#
1(
b101111101100100 +
b101111101100100 1
#71390000000
0#
0(
#71400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#71450000000
0$
0)
#71460000000
1"
1'
b0 +
b0 1
#71510000000
0"
0'
#71520000000
1#
1(
b101111101100100 +
b101111101100100 1
#71570000000
0#
0(
#71580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#71630000000
0$
0)
#71640000000
1"
1'
b0 +
b0 1
#71690000000
0"
0'
#71700000000
1#
1(
b101111101100100 +
b101111101100100 1
#71750000000
0#
0(
#71760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#71810000000
0$
0)
#71820000000
1"
1'
b0 +
b0 1
#71870000000
0"
0'
#71880000000
1#
1(
b101111101100100 +
b101111101100100 1
#71930000000
0#
0(
#71940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#71990000000
0$
0)
#72000000000
1"
1'
b0 +
b0 1
#72050000000
0"
0'
#72060000000
1#
1(
b101111101100100 +
b101111101100100 1
#72110000000
0#
0(
#72120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#72170000000
0$
0)
#72180000000
1"
1'
b0 +
b0 1
#72230000000
0"
0'
#72240000000
1#
1(
b101111101100100 +
b101111101100100 1
#72290000000
0#
0(
#72300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#72350000000
0$
0)
#72360000000
1"
1'
b0 +
b0 1
#72410000000
0"
0'
#72420000000
1#
1(
b101111101100100 +
b101111101100100 1
#72470000000
0#
0(
#72480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#72530000000
0$
0)
#72540000000
1"
1'
b0 +
b0 1
#72590000000
0"
0'
#72600000000
1#
1(
b101111101100100 +
b101111101100100 1
#72650000000
0#
0(
#72660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#72710000000
0$
0)
#72720000000
1"
1'
b0 +
b0 1
#72770000000
0"
0'
#72780000000
1#
1(
b101111101100100 +
b101111101100100 1
#72830000000
0#
0(
#72840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#72890000000
0$
0)
#72900000000
1"
1'
b0 +
b0 1
#72950000000
0"
0'
#72960000000
1#
1(
b101111101100100 +
b101111101100100 1
#73010000000
0#
0(
#73020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#73070000000
0$
0)
#73080000000
1"
1'
b0 +
b0 1
#73130000000
0"
0'
#73140000000
1#
1(
b101111101100100 +
b101111101100100 1
#73190000000
0#
0(
#73200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#73250000000
0$
0)
#73260000000
1"
1'
b0 +
b0 1
#73310000000
0"
0'
#73320000000
1#
1(
b101111101100100 +
b101111101100100 1
#73370000000
0#
0(
#73380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#73430000000
0$
0)
#73440000000
1"
1'
b0 +
b0 1
#73490000000
0"
0'
#73500000000
1#
1(
b101111101100100 +
b101111101100100 1
#73550000000
0#
0(
#73560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#73610000000
0$
0)
#73620000000
1"
1'
b0 +
b0 1
#73670000000
0"
0'
#73680000000
1#
1(
b101111101100100 +
b101111101100100 1
#73730000000
0#
0(
#73740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#73790000000
0$
0)
#73800000000
1"
1'
b0 +
b0 1
#73850000000
0"
0'
#73860000000
1#
1(
b101111101100100 +
b101111101100100 1
#73910000000
0#
0(
#73920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#73970000000
0$
0)
#73980000000
1"
1'
b0 +
b0 1
#74030000000
0"
0'
#74040000000
1#
1(
b101111101100100 +
b101111101100100 1
#74090000000
0#
0(
#74100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#74150000000
0$
0)
#74160000000
1"
1'
b0 +
b0 1
#74210000000
0"
0'
#74220000000
1#
1(
b101111101100100 +
b101111101100100 1
#74270000000
0#
0(
#74280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#74330000000
0$
0)
#74340000000
1"
1'
b0 +
b0 1
#74390000000
0"
0'
#74400000000
1#
1(
b101111101100100 +
b101111101100100 1
#74450000000
0#
0(
#74460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#74510000000
0$
0)
#74520000000
1"
1'
b0 +
b0 1
#74570000000
0"
0'
#74580000000
1#
1(
b101111101100100 +
b101111101100100 1
#74630000000
0#
0(
#74640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#74690000000
0$
0)
#74700000000
1"
1'
b0 +
b0 1
#74750000000
0"
0'
#74760000000
1#
1(
b101111101100100 +
b101111101100100 1
#74810000000
0#
0(
#74820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#74870000000
0$
0)
#74880000000
1"
1'
b0 +
b0 1
#74930000000
0"
0'
#74940000000
1#
1(
b101111101100100 +
b101111101100100 1
#74990000000
0#
0(
#75000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#75050000000
0$
0)
#75060000000
1"
1'
b0 +
b0 1
#75110000000
0"
0'
#75120000000
1#
1(
b101111101100100 +
b101111101100100 1
#75170000000
0#
0(
#75180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#75230000000
0$
0)
#75240000000
1"
1'
b0 +
b0 1
#75290000000
0"
0'
#75300000000
1#
1(
b101111101100100 +
b101111101100100 1
#75350000000
0#
0(
#75360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#75410000000
0$
0)
#75420000000
1"
1'
b0 +
b0 1
#75470000000
0"
0'
#75480000000
1#
1(
b101111101100100 +
b101111101100100 1
#75530000000
0#
0(
#75540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#75590000000
0$
0)
#75600000000
1"
1'
b0 +
b0 1
#75650000000
0"
0'
#75660000000
1#
1(
b101111101100100 +
b101111101100100 1
#75710000000
0#
0(
#75720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#75770000000
0$
0)
#75780000000
1"
1'
b0 +
b0 1
#75830000000
0"
0'
#75840000000
1#
1(
b101111101100100 +
b101111101100100 1
#75890000000
0#
0(
#75900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#75950000000
0$
0)
#75960000000
1"
1'
b0 +
b0 1
#76010000000
0"
0'
#76020000000
1#
1(
b101111101100100 +
b101111101100100 1
#76070000000
0#
0(
#76080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#76130000000
0$
0)
#76140000000
1"
1'
b0 +
b0 1
#76190000000
0"
0'
#76200000000
1#
1(
b101111101100100 +
b101111101100100 1
#76250000000
0#
0(
#76260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#76310000000
0$
0)
#76320000000
1"
1'
b0 +
b0 1
#76370000000
0"
0'
#76380000000
1#
1(
b101111101100100 +
b101111101100100 1
#76430000000
0#
0(
#76440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#76490000000
0$
0)
#76500000000
1"
1'
b0 +
b0 1
#76550000000
0"
0'
#76560000000
1#
1(
b101111101100100 +
b101111101100100 1
#76610000000
0#
0(
#76620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#76670000000
0$
0)
#76680000000
1"
1'
b0 +
b0 1
#76730000000
0"
0'
#76740000000
1#
1(
b101111101100100 +
b101111101100100 1
#76790000000
0#
0(
#76800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#76850000000
0$
0)
#76860000000
1"
1'
b0 +
b0 1
#76910000000
0"
0'
#76920000000
1#
1(
b101111101100100 +
b101111101100100 1
#76970000000
0#
0(
#76980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#77030000000
0$
0)
#77040000000
1"
1'
b0 +
b0 1
#77090000000
0"
0'
#77100000000
1#
1(
b101111101100100 +
b101111101100100 1
#77150000000
0#
0(
#77160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#77210000000
0$
0)
#77220000000
1"
1'
b0 +
b0 1
#77270000000
0"
0'
#77280000000
1#
1(
b101111101100100 +
b101111101100100 1
#77330000000
0#
0(
#77340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#77390000000
0$
0)
#77400000000
1"
1'
b0 +
b0 1
#77450000000
0"
0'
#77460000000
1#
1(
b101111101100100 +
b101111101100100 1
#77510000000
0#
0(
#77520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#77570000000
0$
0)
#77580000000
1"
1'
b0 +
b0 1
#77630000000
0"
0'
#77640000000
1#
1(
b101111101100100 +
b101111101100100 1
#77690000000
0#
0(
#77700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#77750000000
0$
0)
#77760000000
1"
1'
b0 +
b0 1
#77810000000
0"
0'
#77820000000
1#
1(
b101111101100100 +
b101111101100100 1
#77870000000
0#
0(
#77880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#77930000000
0$
0)
#77940000000
1"
1'
b0 +
b0 1
#77990000000
0"
0'
#78000000000
1#
1(
b101111101100100 +
b101111101100100 1
#78050000000
0#
0(
#78060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#78110000000
0$
0)
#78120000000
1"
1'
b0 +
b0 1
#78170000000
0"
0'
#78180000000
1#
1(
b101111101100100 +
b101111101100100 1
#78230000000
0#
0(
#78240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#78290000000
0$
0)
#78300000000
1"
1'
b0 +
b0 1
#78350000000
0"
0'
#78360000000
1#
1(
b101111101100100 +
b101111101100100 1
#78410000000
0#
0(
#78420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#78470000000
0$
0)
#78480000000
1"
1'
b0 +
b0 1
#78530000000
0"
0'
#78540000000
1#
1(
b101111101100100 +
b101111101100100 1
#78590000000
0#
0(
#78600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#78650000000
0$
0)
#78660000000
1"
1'
b0 +
b0 1
#78710000000
0"
0'
#78720000000
1#
1(
b101111101100100 +
b101111101100100 1
#78770000000
0#
0(
#78780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#78830000000
0$
0)
#78840000000
1"
1'
b0 +
b0 1
#78890000000
0"
0'
#78900000000
1#
1(
b101111101100100 +
b101111101100100 1
#78950000000
0#
0(
#78960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#79010000000
0$
0)
#79020000000
1"
1'
b0 +
b0 1
#79070000000
0"
0'
#79080000000
1#
1(
b101111101100100 +
b101111101100100 1
#79130000000
0#
0(
#79140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#79190000000
0$
0)
#79200000000
1"
1'
b0 +
b0 1
#79250000000
0"
0'
#79260000000
1#
1(
b101111101100100 +
b101111101100100 1
#79310000000
0#
0(
#79320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#79370000000
0$
0)
#79380000000
1"
1'
b0 +
b0 1
#79430000000
0"
0'
#79440000000
1#
1(
b101111101100100 +
b101111101100100 1
#79490000000
0#
0(
#79500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#79550000000
0$
0)
#79560000000
1"
1'
b0 +
b0 1
#79610000000
0"
0'
#79620000000
1#
1(
b101111101100100 +
b101111101100100 1
#79670000000
0#
0(
#79680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#79730000000
0$
0)
#79740000000
1"
1'
b0 +
b0 1
#79790000000
0"
0'
#79800000000
1#
1(
b101111101100100 +
b101111101100100 1
#79850000000
0#
0(
#79860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#79910000000
0$
0)
#79920000000
1"
1'
b0 +
b0 1
#79970000000
0"
0'
#79980000000
1#
1(
b101111101100100 +
b101111101100100 1
#80030000000
0#
0(
#80040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#80090000000
0$
0)
#80100000000
1"
1'
b0 +
b0 1
#80150000000
0"
0'
#80160000000
1#
1(
b101111101100100 +
b101111101100100 1
#80210000000
0#
0(
#80220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#80270000000
0$
0)
#80280000000
1"
1'
b0 +
b0 1
#80330000000
0"
0'
#80340000000
1#
1(
b101111101100100 +
b101111101100100 1
#80390000000
0#
0(
#80400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#80450000000
0$
0)
#80460000000
1"
1'
b0 +
b0 1
#80510000000
0"
0'
#80520000000
1#
1(
b101111101100100 +
b101111101100100 1
#80570000000
0#
0(
#80580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#80630000000
0$
0)
#80640000000
1"
1'
b0 +
b0 1
#80690000000
0"
0'
#80700000000
1#
1(
b101111101100100 +
b101111101100100 1
#80750000000
0#
0(
#80760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#80810000000
0$
0)
#80820000000
1"
1'
b0 +
b0 1
#80870000000
0"
0'
#80880000000
1#
1(
b101111101100100 +
b101111101100100 1
#80930000000
0#
0(
#80940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#80990000000
0$
0)
#81000000000
1"
1'
b0 +
b0 1
#81050000000
0"
0'
#81060000000
1#
1(
b101111101100100 +
b101111101100100 1
#81110000000
0#
0(
#81120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#81170000000
0$
0)
#81180000000
1"
1'
b0 +
b0 1
#81230000000
0"
0'
#81240000000
1#
1(
b101111101100100 +
b101111101100100 1
#81290000000
0#
0(
#81300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#81350000000
0$
0)
#81360000000
1"
1'
b0 +
b0 1
#81410000000
0"
0'
#81420000000
1#
1(
b101111101100100 +
b101111101100100 1
#81470000000
0#
0(
#81480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#81530000000
0$
0)
#81540000000
1"
1'
b0 +
b0 1
#81590000000
0"
0'
#81600000000
1#
1(
b101111101100100 +
b101111101100100 1
#81650000000
0#
0(
#81660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#81710000000
0$
0)
#81720000000
1"
1'
b0 +
b0 1
#81770000000
0"
0'
#81780000000
1#
1(
b101111101100100 +
b101111101100100 1
#81830000000
0#
0(
#81840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#81890000000
0$
0)
#81900000000
1"
1'
b0 +
b0 1
#81950000000
0"
0'
#81960000000
1#
1(
b101111101100100 +
b101111101100100 1
#82010000000
0#
0(
#82020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#82070000000
0$
0)
#82080000000
1"
1'
b0 +
b0 1
#82130000000
0"
0'
#82140000000
1#
1(
b101111101100100 +
b101111101100100 1
#82190000000
0#
0(
#82200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#82250000000
0$
0)
#82260000000
1"
1'
b0 +
b0 1
#82310000000
0"
0'
#82320000000
1#
1(
b101111101100100 +
b101111101100100 1
#82370000000
0#
0(
#82380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#82430000000
0$
0)
#82440000000
1"
1'
b0 +
b0 1
#82490000000
0"
0'
#82500000000
1#
1(
b101111101100100 +
b101111101100100 1
#82550000000
0#
0(
#82560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#82610000000
0$
0)
#82620000000
1"
1'
b0 +
b0 1
#82670000000
0"
0'
#82680000000
1#
1(
b101111101100100 +
b101111101100100 1
#82730000000
0#
0(
#82740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#82790000000
0$
0)
#82800000000
1"
1'
b0 +
b0 1
#82850000000
0"
0'
#82860000000
1#
1(
b101111101100100 +
b101111101100100 1
#82910000000
0#
0(
#82920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#82970000000
0$
0)
#82980000000
1"
1'
b0 +
b0 1
#83030000000
0"
0'
#83040000000
1#
1(
b101111101100100 +
b101111101100100 1
#83090000000
0#
0(
#83100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#83150000000
0$
0)
#83160000000
1"
1'
b0 +
b0 1
#83210000000
0"
0'
#83220000000
1#
1(
b101111101100100 +
b101111101100100 1
#83270000000
0#
0(
#83280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#83330000000
0$
0)
#83340000000
1"
1'
b0 +
b0 1
#83390000000
0"
0'
#83400000000
1#
1(
b101111101100100 +
b101111101100100 1
#83450000000
0#
0(
#83460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#83510000000
0$
0)
#83520000000
1"
1'
b0 +
b0 1
#83570000000
0"
0'
#83580000000
1#
1(
b101111101100100 +
b101111101100100 1
#83630000000
0#
0(
#83640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#83690000000
0$
0)
#83700000000
1"
1'
b0 +
b0 1
#83750000000
0"
0'
#83760000000
1#
1(
b101111101100100 +
b101111101100100 1
#83810000000
0#
0(
#83820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#83870000000
0$
0)
#83880000000
1"
1'
b0 +
b0 1
#83930000000
0"
0'
#83940000000
1#
1(
b101111101100100 +
b101111101100100 1
#83990000000
0#
0(
#84000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#84050000000
0$
0)
#84060000000
1"
1'
b0 +
b0 1
#84110000000
0"
0'
#84120000000
1#
1(
b101111101100100 +
b101111101100100 1
#84170000000
0#
0(
#84180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#84230000000
0$
0)
#84240000000
1"
1'
b0 +
b0 1
#84290000000
0"
0'
#84300000000
1#
1(
b101111101100100 +
b101111101100100 1
#84350000000
0#
0(
#84360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#84410000000
0$
0)
#84420000000
1"
1'
b0 +
b0 1
#84470000000
0"
0'
#84480000000
1#
1(
b101111101100100 +
b101111101100100 1
#84530000000
0#
0(
#84540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#84590000000
0$
0)
#84600000000
1"
1'
b0 +
b0 1
#84650000000
0"
0'
#84660000000
1#
1(
b101111101100100 +
b101111101100100 1
#84710000000
0#
0(
#84720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#84770000000
0$
0)
#84780000000
1"
1'
b0 +
b0 1
#84830000000
0"
0'
#84840000000
1#
1(
b101111101100100 +
b101111101100100 1
#84890000000
0#
0(
#84900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#84950000000
0$
0)
#84960000000
1"
1'
b0 +
b0 1
#85010000000
0"
0'
#85020000000
1#
1(
b101111101100100 +
b101111101100100 1
#85070000000
0#
0(
#85080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#85130000000
0$
0)
#85140000000
1"
1'
b0 +
b0 1
#85190000000
0"
0'
#85200000000
1#
1(
b101111101100100 +
b101111101100100 1
#85250000000
0#
0(
#85260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#85310000000
0$
0)
#85320000000
1"
1'
b0 +
b0 1
#85370000000
0"
0'
#85380000000
1#
1(
b101111101100100 +
b101111101100100 1
#85430000000
0#
0(
#85440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#85490000000
0$
0)
#85500000000
1"
1'
b0 +
b0 1
#85550000000
0"
0'
#85560000000
1#
1(
b101111101100100 +
b101111101100100 1
#85610000000
0#
0(
#85620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#85670000000
0$
0)
#85680000000
1"
1'
b0 +
b0 1
#85730000000
0"
0'
#85740000000
1#
1(
b101111101100100 +
b101111101100100 1
#85790000000
0#
0(
#85800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#85850000000
0$
0)
#85860000000
1"
1'
b0 +
b0 1
#85910000000
0"
0'
#85920000000
1#
1(
b101111101100100 +
b101111101100100 1
#85970000000
0#
0(
#85980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#86030000000
0$
0)
#86040000000
1"
1'
b0 +
b0 1
#86090000000
0"
0'
#86100000000
1#
1(
b101111101100100 +
b101111101100100 1
#86150000000
0#
0(
#86160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#86210000000
0$
0)
#86220000000
1"
1'
b0 +
b0 1
#86270000000
0"
0'
#86280000000
1#
1(
b101111101100100 +
b101111101100100 1
#86330000000
0#
0(
#86340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#86390000000
0$
0)
#86400000000
1"
1'
b0 +
b0 1
#86450000000
0"
0'
#86460000000
1#
1(
b101111101100100 +
b101111101100100 1
#86510000000
0#
0(
#86520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#86570000000
0$
0)
#86580000000
1"
1'
b0 +
b0 1
#86630000000
0"
0'
#86640000000
1#
1(
b101111101100100 +
b101111101100100 1
#86690000000
0#
0(
#86700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#86750000000
0$
0)
#86760000000
1"
1'
b0 +
b0 1
#86810000000
0"
0'
#86820000000
1#
1(
b101111101100100 +
b101111101100100 1
#86870000000
0#
0(
#86880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#86930000000
0$
0)
#86940000000
1"
1'
b0 +
b0 1
#86990000000
0"
0'
#87000000000
1#
1(
b101111101100100 +
b101111101100100 1
#87050000000
0#
0(
#87060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#87110000000
0$
0)
#87120000000
1"
1'
b0 +
b0 1
#87170000000
0"
0'
#87180000000
1#
1(
b101111101100100 +
b101111101100100 1
#87230000000
0#
0(
#87240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#87290000000
0$
0)
#87300000000
1"
1'
b0 +
b0 1
#87350000000
0"
0'
#87360000000
1#
1(
b101111101100100 +
b101111101100100 1
#87410000000
0#
0(
#87420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#87470000000
0$
0)
#87480000000
1"
1'
b0 +
b0 1
#87530000000
0"
0'
#87540000000
1#
1(
b101111101100100 +
b101111101100100 1
#87590000000
0#
0(
#87600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#87650000000
0$
0)
#87660000000
1"
1'
b0 +
b0 1
#87710000000
0"
0'
#87720000000
1#
1(
b101111101100100 +
b101111101100100 1
#87770000000
0#
0(
#87780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#87830000000
0$
0)
#87840000000
1"
1'
b0 +
b0 1
#87890000000
0"
0'
#87900000000
1#
1(
b101111101100100 +
b101111101100100 1
#87950000000
0#
0(
#87960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#88010000000
0$
0)
#88020000000
1"
1'
b0 +
b0 1
#88070000000
0"
0'
#88080000000
1#
1(
b101111101100100 +
b101111101100100 1
#88130000000
0#
0(
#88140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#88190000000
0$
0)
#88200000000
1"
1'
b0 +
b0 1
#88250000000
0"
0'
#88260000000
1#
1(
b101111101100100 +
b101111101100100 1
#88310000000
0#
0(
#88320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#88370000000
0$
0)
#88380000000
1"
1'
b0 +
b0 1
#88430000000
0"
0'
#88440000000
1#
1(
b101111101100100 +
b101111101100100 1
#88490000000
0#
0(
#88500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#88550000000
0$
0)
#88560000000
1"
1'
b0 +
b0 1
#88610000000
0"
0'
#88620000000
1#
1(
b101111101100100 +
b101111101100100 1
#88670000000
0#
0(
#88680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#88730000000
0$
0)
#88740000000
1"
1'
b0 +
b0 1
#88790000000
0"
0'
#88800000000
1#
1(
b101111101100100 +
b101111101100100 1
#88850000000
0#
0(
#88860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#88910000000
0$
0)
#88920000000
1"
1'
b0 +
b0 1
#88970000000
0"
0'
#88980000000
1#
1(
b101111101100100 +
b101111101100100 1
#89030000000
0#
0(
#89040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#89090000000
0$
0)
#89100000000
1"
1'
b0 +
b0 1
#89150000000
0"
0'
#89160000000
1#
1(
b101111101100100 +
b101111101100100 1
#89210000000
0#
0(
#89220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#89270000000
0$
0)
#89280000000
1"
1'
b0 +
b0 1
#89330000000
0"
0'
#89340000000
1#
1(
b101111101100100 +
b101111101100100 1
#89390000000
0#
0(
#89400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#89450000000
0$
0)
#89460000000
1"
1'
b0 +
b0 1
#89510000000
0"
0'
#89520000000
1#
1(
b101111101100100 +
b101111101100100 1
#89570000000
0#
0(
#89580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#89630000000
0$
0)
#89640000000
1"
1'
b0 +
b0 1
#89690000000
0"
0'
#89700000000
1#
1(
b101111101100100 +
b101111101100100 1
#89750000000
0#
0(
#89760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#89810000000
0$
0)
#89820000000
1"
1'
b0 +
b0 1
#89870000000
0"
0'
#89880000000
1#
1(
b101111101100100 +
b101111101100100 1
#89930000000
0#
0(
#89940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#89990000000
0$
0)
#90000000000
1"
1'
b0 +
b0 1
#90050000000
0"
0'
#90060000000
1#
1(
b101111101100100 +
b101111101100100 1
#90110000000
0#
0(
#90120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#90170000000
0$
0)
#90180000000
1"
1'
b0 +
b0 1
#90230000000
0"
0'
#90240000000
1#
1(
b101111101100100 +
b101111101100100 1
#90290000000
0#
0(
#90300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#90350000000
0$
0)
#90360000000
1"
1'
b0 +
b0 1
#90410000000
0"
0'
#90420000000
1#
1(
b101111101100100 +
b101111101100100 1
#90470000000
0#
0(
#90480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#90530000000
0$
0)
#90540000000
1"
1'
b0 +
b0 1
#90590000000
0"
0'
#90600000000
1#
1(
b101111101100100 +
b101111101100100 1
#90650000000
0#
0(
#90660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#90710000000
0$
0)
#90720000000
1"
1'
b0 +
b0 1
#90770000000
0"
0'
#90780000000
1#
1(
b101111101100100 +
b101111101100100 1
#90830000000
0#
0(
#90840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#90890000000
0$
0)
#90900000000
1"
1'
b0 +
b0 1
#90950000000
0"
0'
#90960000000
1#
1(
b101111101100100 +
b101111101100100 1
#91010000000
0#
0(
#91020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#91070000000
0$
0)
#91080000000
1"
1'
b0 +
b0 1
#91130000000
0"
0'
#91140000000
1#
1(
b101111101100100 +
b101111101100100 1
#91190000000
0#
0(
#91200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#91250000000
0$
0)
#91260000000
1"
1'
b0 +
b0 1
#91310000000
0"
0'
#91320000000
1#
1(
b101111101100100 +
b101111101100100 1
#91370000000
0#
0(
#91380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#91430000000
0$
0)
#91440000000
1"
1'
b0 +
b0 1
#91490000000
0"
0'
#91500000000
1#
1(
b101111101100100 +
b101111101100100 1
#91550000000
0#
0(
#91560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#91610000000
0$
0)
#91620000000
1"
1'
b0 +
b0 1
#91670000000
0"
0'
#91680000000
1#
1(
b101111101100100 +
b101111101100100 1
#91730000000
0#
0(
#91740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#91790000000
0$
0)
#91800000000
1"
1'
b0 +
b0 1
#91850000000
0"
0'
#91860000000
1#
1(
b101111101100100 +
b101111101100100 1
#91910000000
0#
0(
#91920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#91970000000
0$
0)
#91980000000
1"
1'
b0 +
b0 1
#92030000000
0"
0'
#92040000000
1#
1(
b101111101100100 +
b101111101100100 1
#92090000000
0#
0(
#92100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#92150000000
0$
0)
#92160000000
1"
1'
b0 +
b0 1
#92210000000
0"
0'
#92220000000
1#
1(
b101111101100100 +
b101111101100100 1
#92270000000
0#
0(
#92280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#92330000000
0$
0)
#92340000000
1"
1'
b0 +
b0 1
#92390000000
0"
0'
#92400000000
1#
1(
b101111101100100 +
b101111101100100 1
#92450000000
0#
0(
#92460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#92510000000
0$
0)
#92520000000
1"
1'
b0 +
b0 1
#92570000000
0"
0'
#92580000000
1#
1(
b101111101100100 +
b101111101100100 1
#92630000000
0#
0(
#92640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#92690000000
0$
0)
#92700000000
1"
1'
b0 +
b0 1
#92750000000
0"
0'
#92760000000
1#
1(
b101111101100100 +
b101111101100100 1
#92810000000
0#
0(
#92820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#92870000000
0$
0)
#92880000000
1"
1'
b0 +
b0 1
#92930000000
0"
0'
#92940000000
1#
1(
b101111101100100 +
b101111101100100 1
#92990000000
0#
0(
#93000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#93050000000
0$
0)
#93060000000
1"
1'
b0 +
b0 1
#93110000000
0"
0'
#93120000000
1#
1(
b101111101100100 +
b101111101100100 1
#93170000000
0#
0(
#93180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#93230000000
0$
0)
#93240000000
1"
1'
b0 +
b0 1
#93290000000
0"
0'
#93300000000
1#
1(
b101111101100100 +
b101111101100100 1
#93350000000
0#
0(
#93360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#93410000000
0$
0)
#93420000000
1"
1'
b0 +
b0 1
#93470000000
0"
0'
#93480000000
1#
1(
b101111101100100 +
b101111101100100 1
#93530000000
0#
0(
#93540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#93590000000
0$
0)
#93600000000
1"
1'
b0 +
b0 1
#93650000000
0"
0'
#93660000000
1#
1(
b101111101100100 +
b101111101100100 1
#93710000000
0#
0(
#93720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#93770000000
0$
0)
#93780000000
1"
1'
b0 +
b0 1
#93830000000
0"
0'
#93840000000
1#
1(
b101111101100100 +
b101111101100100 1
#93890000000
0#
0(
#93900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#93950000000
0$
0)
#93960000000
1"
1'
b0 +
b0 1
#94010000000
0"
0'
#94020000000
1#
1(
b101111101100100 +
b101111101100100 1
#94070000000
0#
0(
#94080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#94130000000
0$
0)
#94140000000
1"
1'
b0 +
b0 1
#94190000000
0"
0'
#94200000000
1#
1(
b101111101100100 +
b101111101100100 1
#94250000000
0#
0(
#94260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#94310000000
0$
0)
#94320000000
1"
1'
b0 +
b0 1
#94370000000
0"
0'
#94380000000
1#
1(
b101111101100100 +
b101111101100100 1
#94430000000
0#
0(
#94440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#94490000000
0$
0)
#94500000000
1"
1'
b0 +
b0 1
#94550000000
0"
0'
#94560000000
1#
1(
b101111101100100 +
b101111101100100 1
#94610000000
0#
0(
#94620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#94670000000
0$
0)
#94680000000
1"
1'
b0 +
b0 1
#94730000000
0"
0'
#94740000000
1#
1(
b101111101100100 +
b101111101100100 1
#94790000000
0#
0(
#94800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#94850000000
0$
0)
#94860000000
1"
1'
b0 +
b0 1
#94910000000
0"
0'
#94920000000
1#
1(
b101111101100100 +
b101111101100100 1
#94970000000
0#
0(
#94980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#95030000000
0$
0)
#95040000000
1"
1'
b0 +
b0 1
#95090000000
0"
0'
#95100000000
1#
1(
b101111101100100 +
b101111101100100 1
#95150000000
0#
0(
#95160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#95210000000
0$
0)
#95220000000
1"
1'
b0 +
b0 1
#95270000000
0"
0'
#95280000000
1#
1(
b101111101100100 +
b101111101100100 1
#95330000000
0#
0(
#95340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#95390000000
0$
0)
#95400000000
1"
1'
b0 +
b0 1
#95450000000
0"
0'
#95460000000
1#
1(
b101111101100100 +
b101111101100100 1
#95510000000
0#
0(
#95520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#95570000000
0$
0)
#95580000000
1"
1'
b0 +
b0 1
#95630000000
0"
0'
#95640000000
1#
1(
b101111101100100 +
b101111101100100 1
#95690000000
0#
0(
#95700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#95750000000
0$
0)
#95760000000
1"
1'
b0 +
b0 1
#95810000000
0"
0'
#95820000000
1#
1(
b101111101100100 +
b101111101100100 1
#95870000000
0#
0(
#95880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#95930000000
0$
0)
#95940000000
1"
1'
b0 +
b0 1
#95990000000
0"
0'
#96000000000
1#
1(
b101111101100100 +
b101111101100100 1
#96050000000
0#
0(
#96060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#96110000000
0$
0)
#96120000000
1"
1'
b0 +
b0 1
#96170000000
0"
0'
#96180000000
1#
1(
b101111101100100 +
b101111101100100 1
#96230000000
0#
0(
#96240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#96290000000
0$
0)
#96300000000
1"
1'
b0 +
b0 1
#96350000000
0"
0'
#96360000000
1#
1(
b101111101100100 +
b101111101100100 1
#96410000000
0#
0(
#96420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#96470000000
0$
0)
#96480000000
1"
1'
b0 +
b0 1
#96530000000
0"
0'
#96540000000
1#
1(
b101111101100100 +
b101111101100100 1
#96590000000
0#
0(
#96600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#96650000000
0$
0)
#96660000000
1"
1'
b0 +
b0 1
#96710000000
0"
0'
#96720000000
1#
1(
b101111101100100 +
b101111101100100 1
#96770000000
0#
0(
#96780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#96830000000
0$
0)
#96840000000
1"
1'
b0 +
b0 1
#96890000000
0"
0'
#96900000000
1#
1(
b101111101100100 +
b101111101100100 1
#96950000000
0#
0(
#96960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#97010000000
0$
0)
#97020000000
1"
1'
b0 +
b0 1
#97070000000
0"
0'
#97080000000
1#
1(
b101111101100100 +
b101111101100100 1
#97130000000
0#
0(
#97140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#97190000000
0$
0)
#97200000000
1"
1'
b0 +
b0 1
#97250000000
0"
0'
#97260000000
1#
1(
b101111101100100 +
b101111101100100 1
#97310000000
0#
0(
#97320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#97370000000
0$
0)
#97380000000
1"
1'
b0 +
b0 1
#97430000000
0"
0'
#97440000000
1#
1(
b101111101100100 +
b101111101100100 1
#97490000000
0#
0(
#97500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#97550000000
0$
0)
#97560000000
1"
1'
b0 +
b0 1
#97610000000
0"
0'
#97620000000
1#
1(
b101111101100100 +
b101111101100100 1
#97670000000
0#
0(
#97680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#97730000000
0$
0)
#97740000000
1"
1'
b0 +
b0 1
#97790000000
0"
0'
#97800000000
1#
1(
b101111101100100 +
b101111101100100 1
#97850000000
0#
0(
#97860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#97910000000
0$
0)
#97920000000
1"
1'
b0 +
b0 1
#97970000000
0"
0'
#97980000000
1#
1(
b101111101100100 +
b101111101100100 1
#98030000000
0#
0(
#98040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#98090000000
0$
0)
#98100000000
1"
1'
b0 +
b0 1
#98150000000
0"
0'
#98160000000
1#
1(
b101111101100100 +
b101111101100100 1
#98210000000
0#
0(
#98220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#98270000000
0$
0)
#98280000000
1"
1'
b0 +
b0 1
#98330000000
0"
0'
#98340000000
1#
1(
b101111101100100 +
b101111101100100 1
#98390000000
0#
0(
#98400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#98450000000
0$
0)
#98460000000
1"
1'
b0 +
b0 1
#98510000000
0"
0'
#98520000000
1#
1(
b101111101100100 +
b101111101100100 1
#98570000000
0#
0(
#98580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#98630000000
0$
0)
#98640000000
1"
1'
b0 +
b0 1
#98690000000
0"
0'
#98700000000
1#
1(
b101111101100100 +
b101111101100100 1
#98750000000
0#
0(
#98760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#98810000000
0$
0)
#98820000000
1"
1'
b0 +
b0 1
#98870000000
0"
0'
#98880000000
1#
1(
b101111101100100 +
b101111101100100 1
#98930000000
0#
0(
#98940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#98990000000
0$
0)
#99000000000
1"
1'
b0 +
b0 1
#99050000000
0"
0'
#99060000000
1#
1(
b101111101100100 +
b101111101100100 1
#99110000000
0#
0(
#99120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#99170000000
0$
0)
#99180000000
1"
1'
b0 +
b0 1
#99230000000
0"
0'
#99240000000
1#
1(
b101111101100100 +
b101111101100100 1
#99290000000
0#
0(
#99300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#99350000000
0$
0)
#99360000000
1"
1'
b0 +
b0 1
#99410000000
0"
0'
#99420000000
1#
1(
b101111101100100 +
b101111101100100 1
#99470000000
0#
0(
#99480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#99530000000
0$
0)
#99540000000
1"
1'
b0 +
b0 1
#99590000000
0"
0'
#99600000000
1#
1(
b101111101100100 +
b101111101100100 1
#99650000000
0#
0(
#99660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#99710000000
0$
0)
#99720000000
1"
1'
b0 +
b0 1
#99770000000
0"
0'
#99780000000
1#
1(
b101111101100100 +
b101111101100100 1
#99830000000
0#
0(
#99840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#99890000000
0$
0)
#99900000000
1"
1'
b0 +
b0 1
#99950000000
0"
0'
#99960000000
1#
1(
b101111101100100 +
b101111101100100 1
#100010000000
0#
0(
#100020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#100070000000
0$
0)
#100080000000
1"
1'
b0 +
b0 1
#100130000000
0"
0'
#100140000000
1#
1(
b101111101100100 +
b101111101100100 1
#100190000000
0#
0(
#100200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#100250000000
0$
0)
#100260000000
1"
1'
b0 +
b0 1
#100310000000
0"
0'
#100320000000
1#
1(
b101111101100100 +
b101111101100100 1
#100370000000
0#
0(
#100380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#100430000000
0$
0)
#100440000000
1"
1'
b0 +
b0 1
#100490000000
0"
0'
#100500000000
1#
1(
b101111101100100 +
b101111101100100 1
#100550000000
0#
0(
#100560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#100610000000
0$
0)
#100620000000
1"
1'
b0 +
b0 1
#100670000000
0"
0'
#100680000000
1#
1(
b101111101100100 +
b101111101100100 1
#100730000000
0#
0(
#100740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#100790000000
0$
0)
#100800000000
1"
1'
b0 +
b0 1
#100850000000
0"
0'
#100860000000
1#
1(
b101111101100100 +
b101111101100100 1
#100910000000
0#
0(
#100920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#100970000000
0$
0)
#100980000000
1"
1'
b0 +
b0 1
#101030000000
0"
0'
#101040000000
1#
1(
b101111101100100 +
b101111101100100 1
#101090000000
0#
0(
#101100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#101150000000
0$
0)
#101160000000
1"
1'
b0 +
b0 1
#101210000000
0"
0'
#101220000000
1#
1(
b101111101100100 +
b101111101100100 1
#101270000000
0#
0(
#101280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#101330000000
0$
0)
#101340000000
1"
1'
b0 +
b0 1
#101390000000
0"
0'
#101400000000
1#
1(
b101111101100100 +
b101111101100100 1
#101450000000
0#
0(
#101460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#101510000000
0$
0)
#101520000000
1"
1'
b0 +
b0 1
#101570000000
0"
0'
#101580000000
1#
1(
b101111101100100 +
b101111101100100 1
#101630000000
0#
0(
#101640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#101690000000
0$
0)
#101700000000
1"
1'
b0 +
b0 1
#101750000000
0"
0'
#101760000000
1#
1(
b101111101100100 +
b101111101100100 1
#101810000000
0#
0(
#101820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#101870000000
0$
0)
#101880000000
1"
1'
b0 +
b0 1
#101930000000
0"
0'
#101940000000
1#
1(
b101111101100100 +
b101111101100100 1
#101990000000
0#
0(
#102000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#102050000000
0$
0)
#102060000000
1"
1'
b0 +
b0 1
#102110000000
0"
0'
#102120000000
1#
1(
b101111101100100 +
b101111101100100 1
#102170000000
0#
0(
#102180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#102230000000
0$
0)
#102240000000
1"
1'
b0 +
b0 1
#102290000000
0"
0'
#102300000000
1#
1(
b101111101100100 +
b101111101100100 1
#102350000000
0#
0(
#102360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#102410000000
0$
0)
#102420000000
1"
1'
b0 +
b0 1
#102470000000
0"
0'
#102480000000
1#
1(
b101111101100100 +
b101111101100100 1
#102530000000
0#
0(
#102540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#102590000000
0$
0)
#102600000000
1"
1'
b0 +
b0 1
#102650000000
0"
0'
#102660000000
1#
1(
b101111101100100 +
b101111101100100 1
#102710000000
0#
0(
#102720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#102770000000
0$
0)
#102780000000
1"
1'
b0 +
b0 1
#102830000000
0"
0'
#102840000000
1#
1(
b101111101100100 +
b101111101100100 1
#102890000000
0#
0(
#102900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#102950000000
0$
0)
#102960000000
1"
1'
b0 +
b0 1
#103010000000
0"
0'
#103020000000
1#
1(
b101111101100100 +
b101111101100100 1
#103070000000
0#
0(
#103080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#103130000000
0$
0)
#103140000000
1"
1'
b0 +
b0 1
#103190000000
0"
0'
#103200000000
1#
1(
b101111101100100 +
b101111101100100 1
#103250000000
0#
0(
#103260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#103310000000
0$
0)
#103320000000
1"
1'
b0 +
b0 1
#103370000000
0"
0'
#103380000000
1#
1(
b101111101100100 +
b101111101100100 1
#103430000000
0#
0(
#103440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#103490000000
0$
0)
#103500000000
1"
1'
b0 +
b0 1
#103550000000
0"
0'
#103560000000
1#
1(
b101111101100100 +
b101111101100100 1
#103610000000
0#
0(
#103620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#103670000000
0$
0)
#103680000000
1"
1'
b0 +
b0 1
#103730000000
0"
0'
#103740000000
1#
1(
b101111101100100 +
b101111101100100 1
#103790000000
0#
0(
#103800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#103850000000
0$
0)
#103860000000
1"
1'
b0 +
b0 1
#103910000000
0"
0'
#103920000000
1#
1(
b101111101100100 +
b101111101100100 1
#103970000000
0#
0(
#103980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#104030000000
0$
0)
#104040000000
1"
1'
b0 +
b0 1
#104090000000
0"
0'
#104100000000
1#
1(
b101111101100100 +
b101111101100100 1
#104150000000
0#
0(
#104160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#104210000000
0$
0)
#104220000000
1"
1'
b0 +
b0 1
#104270000000
0"
0'
#104280000000
1#
1(
b101111101100100 +
b101111101100100 1
#104330000000
0#
0(
#104340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#104390000000
0$
0)
#104400000000
1"
1'
b0 +
b0 1
#104450000000
0"
0'
#104460000000
1#
1(
b101111101100100 +
b101111101100100 1
#104510000000
0#
0(
#104520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#104570000000
0$
0)
#104580000000
1"
1'
b0 +
b0 1
#104630000000
0"
0'
#104640000000
1#
1(
b101111101100100 +
b101111101100100 1
#104690000000
0#
0(
#104700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#104750000000
0$
0)
#104760000000
1"
1'
b0 +
b0 1
#104810000000
0"
0'
#104820000000
1#
1(
b101111101100100 +
b101111101100100 1
#104870000000
0#
0(
#104880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#104930000000
0$
0)
#104940000000
1"
1'
b0 +
b0 1
#104990000000
0"
0'
#105000000000
1#
1(
b101111101100100 +
b101111101100100 1
#105050000000
0#
0(
#105060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#105110000000
0$
0)
#105120000000
1"
1'
b0 +
b0 1
#105170000000
0"
0'
#105180000000
1#
1(
b101111101100100 +
b101111101100100 1
#105230000000
0#
0(
#105240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#105290000000
0$
0)
#105300000000
1"
1'
b0 +
b0 1
#105350000000
0"
0'
#105360000000
1#
1(
b101111101100100 +
b101111101100100 1
#105410000000
0#
0(
#105420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#105470000000
0$
0)
#105480000000
1"
1'
b0 +
b0 1
#105530000000
0"
0'
#105540000000
1#
1(
b101111101100100 +
b101111101100100 1
#105590000000
0#
0(
#105600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#105650000000
0$
0)
#105660000000
1"
1'
b0 +
b0 1
#105710000000
0"
0'
#105720000000
1#
1(
b101111101100100 +
b101111101100100 1
#105770000000
0#
0(
#105780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#105830000000
0$
0)
#105840000000
1"
1'
b0 +
b0 1
#105890000000
0"
0'
#105900000000
1#
1(
b101111101100100 +
b101111101100100 1
#105950000000
0#
0(
#105960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#106010000000
0$
0)
#106020000000
1"
1'
b0 +
b0 1
#106070000000
0"
0'
#106080000000
1#
1(
b101111101100100 +
b101111101100100 1
#106130000000
0#
0(
#106140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#106190000000
0$
0)
#106200000000
1"
1'
b0 +
b0 1
#106250000000
0"
0'
#106260000000
1#
1(
b101111101100100 +
b101111101100100 1
#106310000000
0#
0(
#106320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#106370000000
0$
0)
#106380000000
1"
1'
b0 +
b0 1
#106430000000
0"
0'
#106440000000
1#
1(
b101111101100100 +
b101111101100100 1
#106490000000
0#
0(
#106500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#106550000000
0$
0)
#106560000000
1"
1'
b0 +
b0 1
#106610000000
0"
0'
#106620000000
1#
1(
b101111101100100 +
b101111101100100 1
#106670000000
0#
0(
#106680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#106730000000
0$
0)
#106740000000
1"
1'
b0 +
b0 1
#106790000000
0"
0'
#106800000000
1#
1(
b101111101100100 +
b101111101100100 1
#106850000000
0#
0(
#106860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#106910000000
0$
0)
#106920000000
1"
1'
b0 +
b0 1
#106970000000
0"
0'
#106980000000
1#
1(
b101111101100100 +
b101111101100100 1
#107030000000
0#
0(
#107040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#107090000000
0$
0)
#107100000000
1"
1'
b0 +
b0 1
#107150000000
0"
0'
#107160000000
1#
1(
b101111101100100 +
b101111101100100 1
#107210000000
0#
0(
#107220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#107270000000
0$
0)
#107280000000
1"
1'
b0 +
b0 1
#107330000000
0"
0'
#107340000000
1#
1(
b101111101100100 +
b101111101100100 1
#107390000000
0#
0(
#107400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#107450000000
0$
0)
#107460000000
1"
1'
b0 +
b0 1
#107510000000
0"
0'
#107520000000
1#
1(
b101111101100100 +
b101111101100100 1
#107570000000
0#
0(
#107580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#107630000000
0$
0)
#107640000000
1"
1'
b0 +
b0 1
#107690000000
0"
0'
#107700000000
1#
1(
b101111101100100 +
b101111101100100 1
#107750000000
0#
0(
#107760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#107810000000
0$
0)
#107820000000
1"
1'
b0 +
b0 1
#107870000000
0"
0'
#107880000000
1#
1(
b101111101100100 +
b101111101100100 1
#107930000000
0#
0(
#107940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#107990000000
0$
0)
#108000000000
1"
1'
b0 +
b0 1
#108050000000
0"
0'
#108060000000
1#
1(
b101111101100100 +
b101111101100100 1
#108110000000
0#
0(
#108120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#108170000000
0$
0)
#108180000000
1"
1'
b0 +
b0 1
#108230000000
0"
0'
#108240000000
1#
1(
b101111101100100 +
b101111101100100 1
#108290000000
0#
0(
#108300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#108350000000
0$
0)
#108360000000
1"
1'
b0 +
b0 1
#108410000000
0"
0'
#108420000000
1#
1(
b101111101100100 +
b101111101100100 1
#108470000000
0#
0(
#108480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#108530000000
0$
0)
#108540000000
1"
1'
b0 +
b0 1
#108590000000
0"
0'
#108600000000
1#
1(
b101111101100100 +
b101111101100100 1
#108650000000
0#
0(
#108660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#108710000000
0$
0)
#108720000000
1"
1'
b0 +
b0 1
#108770000000
0"
0'
#108780000000
1#
1(
b101111101100100 +
b101111101100100 1
#108830000000
0#
0(
#108840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#108890000000
0$
0)
#108900000000
1"
1'
b0 +
b0 1
#108950000000
0"
0'
#108960000000
1#
1(
b101111101100100 +
b101111101100100 1
#109010000000
0#
0(
#109020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#109070000000
0$
0)
#109080000000
1"
1'
b0 +
b0 1
#109130000000
0"
0'
#109140000000
1#
1(
b101111101100100 +
b101111101100100 1
#109190000000
0#
0(
#109200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#109250000000
0$
0)
#109260000000
1"
1'
b0 +
b0 1
#109310000000
0"
0'
#109320000000
1#
1(
b101111101100100 +
b101111101100100 1
#109370000000
0#
0(
#109380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#109430000000
0$
0)
#109440000000
1"
1'
b0 +
b0 1
#109490000000
0"
0'
#109500000000
1#
1(
b101111101100100 +
b101111101100100 1
#109550000000
0#
0(
#109560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#109610000000
0$
0)
#109620000000
1"
1'
b0 +
b0 1
#109670000000
0"
0'
#109680000000
1#
1(
b101111101100100 +
b101111101100100 1
#109730000000
0#
0(
#109740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#109790000000
0$
0)
#109800000000
1"
1'
b0 +
b0 1
#109850000000
0"
0'
#109860000000
1#
1(
b101111101100100 +
b101111101100100 1
#109910000000
0#
0(
#109920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#109970000000
0$
0)
#109980000000
1"
1'
b0 +
b0 1
#110030000000
0"
0'
#110040000000
1#
1(
b101111101100100 +
b101111101100100 1
#110090000000
0#
0(
#110100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#110150000000
0$
0)
#110160000000
1"
1'
b0 +
b0 1
#110210000000
0"
0'
#110220000000
1#
1(
b101111101100100 +
b101111101100100 1
#110270000000
0#
0(
#110280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#110330000000
0$
0)
#110340000000
1"
1'
b0 +
b0 1
#110390000000
0"
0'
#110400000000
1#
1(
b101111101100100 +
b101111101100100 1
#110450000000
0#
0(
#110460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#110510000000
0$
0)
#110520000000
1"
1'
b0 +
b0 1
#110570000000
0"
0'
#110580000000
1#
1(
b101111101100100 +
b101111101100100 1
#110630000000
0#
0(
#110640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#110690000000
0$
0)
#110700000000
1"
1'
b0 +
b0 1
#110750000000
0"
0'
#110760000000
1#
1(
b101111101100100 +
b101111101100100 1
#110810000000
0#
0(
#110820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#110870000000
0$
0)
#110880000000
1"
1'
b0 +
b0 1
#110930000000
0"
0'
#110940000000
1#
1(
b101111101100100 +
b101111101100100 1
#110990000000
0#
0(
#111000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#111050000000
0$
0)
#111060000000
1"
1'
b0 +
b0 1
#111110000000
0"
0'
#111120000000
1#
1(
b101111101100100 +
b101111101100100 1
#111170000000
0#
0(
#111180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#111230000000
0$
0)
#111240000000
1"
1'
b0 +
b0 1
#111290000000
0"
0'
#111300000000
1#
1(
b101111101100100 +
b101111101100100 1
#111350000000
0#
0(
#111360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#111410000000
0$
0)
#111420000000
1"
1'
b0 +
b0 1
#111470000000
0"
0'
#111480000000
1#
1(
b101111101100100 +
b101111101100100 1
#111530000000
0#
0(
#111540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#111590000000
0$
0)
#111600000000
1"
1'
b0 +
b0 1
#111650000000
0"
0'
#111660000000
1#
1(
b101111101100100 +
b101111101100100 1
#111710000000
0#
0(
#111720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#111770000000
0$
0)
#111780000000
1"
1'
b0 +
b0 1
#111830000000
0"
0'
#111840000000
1#
1(
b101111101100100 +
b101111101100100 1
#111890000000
0#
0(
#111900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#111950000000
0$
0)
#111960000000
1"
1'
b0 +
b0 1
#112010000000
0"
0'
#112020000000
1#
1(
b101111101100100 +
b101111101100100 1
#112070000000
0#
0(
#112080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#112130000000
0$
0)
#112140000000
1"
1'
b0 +
b0 1
#112190000000
0"
0'
#112200000000
1#
1(
b101111101100100 +
b101111101100100 1
#112250000000
0#
0(
#112260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#112310000000
0$
0)
#112320000000
1"
1'
b0 +
b0 1
#112370000000
0"
0'
#112380000000
1#
1(
b101111101100100 +
b101111101100100 1
#112430000000
0#
0(
#112440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#112490000000
0$
0)
#112500000000
1"
1'
b0 +
b0 1
#112550000000
0"
0'
#112560000000
1#
1(
b101111101100100 +
b101111101100100 1
#112610000000
0#
0(
#112620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#112670000000
0$
0)
#112680000000
1"
1'
b0 +
b0 1
#112730000000
0"
0'
#112740000000
1#
1(
b101111101100100 +
b101111101100100 1
#112790000000
0#
0(
#112800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#112850000000
0$
0)
#112860000000
1"
1'
b0 +
b0 1
#112910000000
0"
0'
#112920000000
1#
1(
b101111101100100 +
b101111101100100 1
#112970000000
0#
0(
#112980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#113030000000
0$
0)
#113040000000
1"
1'
b0 +
b0 1
#113090000000
0"
0'
#113100000000
1#
1(
b101111101100100 +
b101111101100100 1
#113150000000
0#
0(
#113160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#113210000000
0$
0)
#113220000000
1"
1'
b0 +
b0 1
#113270000000
0"
0'
#113280000000
1#
1(
b101111101100100 +
b101111101100100 1
#113330000000
0#
0(
#113340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#113390000000
0$
0)
#113400000000
1"
1'
b0 +
b0 1
#113450000000
0"
0'
#113460000000
1#
1(
b101111101100100 +
b101111101100100 1
#113510000000
0#
0(
#113520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#113570000000
0$
0)
#113580000000
1"
1'
b0 +
b0 1
#113630000000
0"
0'
#113640000000
1#
1(
b101111101100100 +
b101111101100100 1
#113690000000
0#
0(
#113700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#113750000000
0$
0)
#113760000000
1"
1'
b0 +
b0 1
#113810000000
0"
0'
#113820000000
1#
1(
b101111101100100 +
b101111101100100 1
#113870000000
0#
0(
#113880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#113930000000
0$
0)
#113940000000
1"
1'
b0 +
b0 1
#113990000000
0"
0'
#114000000000
1#
1(
b101111101100100 +
b101111101100100 1
#114050000000
0#
0(
#114060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#114110000000
0$
0)
#114120000000
1"
1'
b0 +
b0 1
#114170000000
0"
0'
#114180000000
1#
1(
b101111101100100 +
b101111101100100 1
#114230000000
0#
0(
#114240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#114290000000
0$
0)
#114300000000
1"
1'
b0 +
b0 1
#114350000000
0"
0'
#114360000000
1#
1(
b101111101100100 +
b101111101100100 1
#114410000000
0#
0(
#114420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#114470000000
0$
0)
#114480000000
1"
1'
b0 +
b0 1
#114530000000
0"
0'
#114540000000
1#
1(
b101111101100100 +
b101111101100100 1
#114590000000
0#
0(
#114600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#114650000000
0$
0)
#114660000000
1"
1'
b0 +
b0 1
#114710000000
0"
0'
#114720000000
1#
1(
b101111101100100 +
b101111101100100 1
#114770000000
0#
0(
#114780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#114830000000
0$
0)
#114840000000
1"
1'
b0 +
b0 1
#114890000000
0"
0'
#114900000000
1#
1(
b101111101100100 +
b101111101100100 1
#114950000000
0#
0(
#114960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#115010000000
0$
0)
#115020000000
1"
1'
b0 +
b0 1
#115070000000
0"
0'
#115080000000
1#
1(
b101111101100100 +
b101111101100100 1
#115130000000
0#
0(
#115140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#115190000000
0$
0)
#115200000000
1"
1'
b0 +
b0 1
#115250000000
0"
0'
#115260000000
1#
1(
b101111101100100 +
b101111101100100 1
#115310000000
0#
0(
#115320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#115370000000
0$
0)
#115380000000
1"
1'
b0 +
b0 1
#115430000000
0"
0'
#115440000000
1#
1(
b101111101100100 +
b101111101100100 1
#115490000000
0#
0(
#115500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#115550000000
0$
0)
#115560000000
1"
1'
b0 +
b0 1
#115610000000
0"
0'
#115620000000
1#
1(
b101111101100100 +
b101111101100100 1
#115670000000
0#
0(
#115680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#115730000000
0$
0)
#115740000000
1"
1'
b0 +
b0 1
#115790000000
0"
0'
#115800000000
1#
1(
b101111101100100 +
b101111101100100 1
#115850000000
0#
0(
#115860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#115910000000
0$
0)
#115920000000
1"
1'
b0 +
b0 1
#115970000000
0"
0'
#115980000000
1#
1(
b101111101100100 +
b101111101100100 1
#116030000000
0#
0(
#116040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#116090000000
0$
0)
#116100000000
1"
1'
b0 +
b0 1
#116150000000
0"
0'
#116160000000
1#
1(
b101111101100100 +
b101111101100100 1
#116210000000
0#
0(
#116220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#116270000000
0$
0)
#116280000000
1"
1'
b0 +
b0 1
#116330000000
0"
0'
#116340000000
1#
1(
b101111101100100 +
b101111101100100 1
#116390000000
0#
0(
#116400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#116450000000
0$
0)
#116460000000
1"
1'
b0 +
b0 1
#116510000000
0"
0'
#116520000000
1#
1(
b101111101100100 +
b101111101100100 1
#116570000000
0#
0(
#116580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#116630000000
0$
0)
#116640000000
1"
1'
b0 +
b0 1
#116690000000
0"
0'
#116700000000
1#
1(
b101111101100100 +
b101111101100100 1
#116750000000
0#
0(
#116760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#116810000000
0$
0)
#116820000000
1"
1'
b0 +
b0 1
#116870000000
0"
0'
#116880000000
1#
1(
b101111101100100 +
b101111101100100 1
#116930000000
0#
0(
#116940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#116990000000
0$
0)
#117000000000
1"
1'
b0 +
b0 1
#117050000000
0"
0'
#117060000000
1#
1(
b101111101100100 +
b101111101100100 1
#117110000000
0#
0(
#117120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#117170000000
0$
0)
#117180000000
1"
1'
b0 +
b0 1
#117230000000
0"
0'
#117240000000
1#
1(
b101111101100100 +
b101111101100100 1
#117290000000
0#
0(
#117300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#117350000000
0$
0)
#117360000000
1"
1'
b0 +
b0 1
#117410000000
0"
0'
#117420000000
1#
1(
b101111101100100 +
b101111101100100 1
#117470000000
0#
0(
#117480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#117530000000
0$
0)
#117540000000
1"
1'
b0 +
b0 1
#117590000000
0"
0'
#117600000000
1#
1(
b101111101100100 +
b101111101100100 1
#117650000000
0#
0(
#117660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#117710000000
0$
0)
#117720000000
1"
1'
b0 +
b0 1
#117770000000
0"
0'
#117780000000
1#
1(
b101111101100100 +
b101111101100100 1
#117830000000
0#
0(
#117840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#117890000000
0$
0)
#117900000000
1"
1'
b0 +
b0 1
#117950000000
0"
0'
#117960000000
1#
1(
b101111101100100 +
b101111101100100 1
#118010000000
0#
0(
#118020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#118070000000
0$
0)
#118080000000
1"
1'
b0 +
b0 1
#118130000000
0"
0'
#118140000000
1#
1(
b101111101100100 +
b101111101100100 1
#118190000000
0#
0(
#118200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#118250000000
0$
0)
#118260000000
1"
1'
b0 +
b0 1
#118310000000
0"
0'
#118320000000
1#
1(
b101111101100100 +
b101111101100100 1
#118370000000
0#
0(
#118380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#118430000000
0$
0)
#118440000000
1"
1'
b0 +
b0 1
#118490000000
0"
0'
#118500000000
1#
1(
b101111101100100 +
b101111101100100 1
#118550000000
0#
0(
#118560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#118610000000
0$
0)
#118620000000
1"
1'
b0 +
b0 1
#118670000000
0"
0'
#118680000000
1#
1(
b101111101100100 +
b101111101100100 1
#118730000000
0#
0(
#118740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#118790000000
0$
0)
#118800000000
1"
1'
b0 +
b0 1
#118850000000
0"
0'
#118860000000
1#
1(
b101111101100100 +
b101111101100100 1
#118910000000
0#
0(
#118920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#118970000000
0$
0)
#118980000000
1"
1'
b0 +
b0 1
#119030000000
0"
0'
#119040000000
1#
1(
b101111101100100 +
b101111101100100 1
#119090000000
0#
0(
#119100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#119150000000
0$
0)
#119160000000
1"
1'
b0 +
b0 1
#119210000000
0"
0'
#119220000000
1#
1(
b101111101100100 +
b101111101100100 1
#119270000000
0#
0(
#119280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#119330000000
0$
0)
#119340000000
1"
1'
b0 +
b0 1
#119390000000
0"
0'
#119400000000
1#
1(
b101111101100100 +
b101111101100100 1
#119450000000
0#
0(
#119460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#119510000000
0$
0)
#119520000000
1"
1'
b0 +
b0 1
#119570000000
0"
0'
#119580000000
1#
1(
b101111101100100 +
b101111101100100 1
#119630000000
0#
0(
#119640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#119690000000
0$
0)
#119700000000
1"
1'
b0 +
b0 1
#119750000000
0"
0'
#119760000000
1#
1(
b101111101100100 +
b101111101100100 1
#119810000000
0#
0(
#119820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#119870000000
0$
0)
#119880000000
1"
1'
b0 +
b0 1
#119930000000
0"
0'
#119940000000
1#
1(
b101111101100100 +
b101111101100100 1
#119990000000
0#
0(
#120000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#120050000000
0$
0)
#120060000000
1"
1'
b0 +
b0 1
#120110000000
0"
0'
#120120000000
1#
1(
b101111101100100 +
b101111101100100 1
#120170000000
0#
0(
#120180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#120230000000
0$
0)
#120240000000
1"
1'
b0 +
b0 1
#120290000000
0"
0'
#120300000000
1#
1(
b101111101100100 +
b101111101100100 1
#120350000000
0#
0(
#120360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#120410000000
0$
0)
#120420000000
1"
1'
b0 +
b0 1
#120470000000
0"
0'
#120480000000
1#
1(
b101111101100100 +
b101111101100100 1
#120530000000
0#
0(
#120540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#120590000000
0$
0)
#120600000000
1"
1'
b0 +
b0 1
#120650000000
0"
0'
#120660000000
1#
1(
b101111101100100 +
b101111101100100 1
#120710000000
0#
0(
#120720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#120770000000
0$
0)
#120780000000
1"
1'
b0 +
b0 1
#120830000000
0"
0'
#120840000000
1#
1(
b101111101100100 +
b101111101100100 1
#120890000000
0#
0(
#120900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#120950000000
0$
0)
#120960000000
1"
1'
b0 +
b0 1
#121010000000
0"
0'
#121020000000
1#
1(
b101111101100100 +
b101111101100100 1
#121070000000
0#
0(
#121080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#121130000000
0$
0)
#121140000000
1"
1'
b0 +
b0 1
#121190000000
0"
0'
#121200000000
1#
1(
b101111101100100 +
b101111101100100 1
#121250000000
0#
0(
#121260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#121310000000
0$
0)
#121320000000
1"
1'
b0 +
b0 1
#121370000000
0"
0'
#121380000000
1#
1(
b101111101100100 +
b101111101100100 1
#121430000000
0#
0(
#121440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#121490000000
0$
0)
#121500000000
1"
1'
b0 +
b0 1
#121550000000
0"
0'
#121560000000
1#
1(
b101111101100100 +
b101111101100100 1
#121610000000
0#
0(
#121620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#121670000000
0$
0)
#121680000000
1"
1'
b0 +
b0 1
#121730000000
0"
0'
#121740000000
1#
1(
b101111101100100 +
b101111101100100 1
#121790000000
0#
0(
#121800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#121850000000
0$
0)
#121860000000
1"
1'
b0 +
b0 1
#121910000000
0"
0'
#121920000000
1#
1(
b101111101100100 +
b101111101100100 1
#121970000000
0#
0(
#121980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#122030000000
0$
0)
#122040000000
1"
1'
b0 +
b0 1
#122090000000
0"
0'
#122100000000
1#
1(
b101111101100100 +
b101111101100100 1
#122150000000
0#
0(
#122160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#122210000000
0$
0)
#122220000000
1"
1'
b0 +
b0 1
#122270000000
0"
0'
#122280000000
1#
1(
b101111101100100 +
b101111101100100 1
#122330000000
0#
0(
#122340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#122390000000
0$
0)
#122400000000
1"
1'
b0 +
b0 1
#122450000000
0"
0'
#122460000000
1#
1(
b101111101100100 +
b101111101100100 1
#122510000000
0#
0(
#122520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#122570000000
0$
0)
#122580000000
1"
1'
b0 +
b0 1
#122630000000
0"
0'
#122640000000
1#
1(
b101111101100100 +
b101111101100100 1
#122690000000
0#
0(
#122700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#122750000000
0$
0)
#122760000000
1"
1'
b0 +
b0 1
#122810000000
0"
0'
#122820000000
1#
1(
b101111101100100 +
b101111101100100 1
#122870000000
0#
0(
#122880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#122930000000
0$
0)
#122940000000
1"
1'
b0 +
b0 1
#122990000000
0"
0'
#123000000000
1#
1(
b101111101100100 +
b101111101100100 1
#123050000000
0#
0(
#123060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#123110000000
0$
0)
#123120000000
1"
1'
b0 +
b0 1
#123170000000
0"
0'
#123180000000
1#
1(
b101111101100100 +
b101111101100100 1
#123230000000
0#
0(
#123240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#123290000000
0$
0)
#123300000000
1"
1'
b0 +
b0 1
#123350000000
0"
0'
#123360000000
1#
1(
b101111101100100 +
b101111101100100 1
#123410000000
0#
0(
#123420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#123470000000
0$
0)
#123480000000
1"
1'
b0 +
b0 1
#123530000000
0"
0'
#123540000000
1#
1(
b101111101100100 +
b101111101100100 1
#123590000000
0#
0(
#123600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#123650000000
0$
0)
#123660000000
1"
1'
b0 +
b0 1
#123710000000
0"
0'
#123720000000
1#
1(
b101111101100100 +
b101111101100100 1
#123770000000
0#
0(
#123780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#123830000000
0$
0)
#123840000000
1"
1'
b0 +
b0 1
#123890000000
0"
0'
#123900000000
1#
1(
b101111101100100 +
b101111101100100 1
#123950000000
0#
0(
#123960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#124010000000
0$
0)
#124020000000
1"
1'
b0 +
b0 1
#124070000000
0"
0'
#124080000000
1#
1(
b101111101100100 +
b101111101100100 1
#124130000000
0#
0(
#124140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#124190000000
0$
0)
#124200000000
1"
1'
b0 +
b0 1
#124250000000
0"
0'
#124260000000
1#
1(
b101111101100100 +
b101111101100100 1
#124310000000
0#
0(
#124320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#124370000000
0$
0)
#124380000000
1"
1'
b0 +
b0 1
#124430000000
0"
0'
#124440000000
1#
1(
b101111101100100 +
b101111101100100 1
#124490000000
0#
0(
#124500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#124550000000
0$
0)
#124560000000
1"
1'
b0 +
b0 1
#124610000000
0"
0'
#124620000000
1#
1(
b101111101100100 +
b101111101100100 1
#124670000000
0#
0(
#124680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#124730000000
0$
0)
#124740000000
1"
1'
b0 +
b0 1
#124790000000
0"
0'
#124800000000
1#
1(
b101111101100100 +
b101111101100100 1
#124850000000
0#
0(
#124860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#124910000000
0$
0)
#124920000000
1"
1'
b0 +
b0 1
#124970000000
0"
0'
#124980000000
1#
1(
b101111101100100 +
b101111101100100 1
#125030000000
0#
0(
#125040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#125090000000
0$
0)
#125100000000
1"
1'
b0 +
b0 1
#125150000000
0"
0'
#125160000000
1#
1(
b101111101100100 +
b101111101100100 1
#125210000000
0#
0(
#125220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#125270000000
0$
0)
#125280000000
1"
1'
b0 +
b0 1
#125330000000
0"
0'
#125340000000
1#
1(
b101111101100100 +
b101111101100100 1
#125390000000
0#
0(
#125400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#125450000000
0$
0)
#125460000000
1"
1'
b0 +
b0 1
#125510000000
0"
0'
#125520000000
1#
1(
b101111101100100 +
b101111101100100 1
#125570000000
0#
0(
#125580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#125630000000
0$
0)
#125640000000
1"
1'
b0 +
b0 1
#125690000000
0"
0'
#125700000000
1#
1(
b101111101100100 +
b101111101100100 1
#125750000000
0#
0(
#125760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#125810000000
0$
0)
#125820000000
1"
1'
b0 +
b0 1
#125870000000
0"
0'
#125880000000
1#
1(
b101111101100100 +
b101111101100100 1
#125930000000
0#
0(
#125940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#125990000000
0$
0)
#126000000000
1"
1'
b0 +
b0 1
#126050000000
0"
0'
#126060000000
1#
1(
b101111101100100 +
b101111101100100 1
#126110000000
0#
0(
#126120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#126170000000
0$
0)
#126180000000
1"
1'
b0 +
b0 1
#126230000000
0"
0'
#126240000000
1#
1(
b101111101100100 +
b101111101100100 1
#126290000000
0#
0(
#126300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#126350000000
0$
0)
#126360000000
1"
1'
b0 +
b0 1
#126410000000
0"
0'
#126420000000
1#
1(
b101111101100100 +
b101111101100100 1
#126470000000
0#
0(
#126480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#126530000000
0$
0)
#126540000000
1"
1'
b0 +
b0 1
#126590000000
0"
0'
#126600000000
1#
1(
b101111101100100 +
b101111101100100 1
#126650000000
0#
0(
#126660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#126710000000
0$
0)
#126720000000
1"
1'
b0 +
b0 1
#126770000000
0"
0'
#126780000000
1#
1(
b101111101100100 +
b101111101100100 1
#126830000000
0#
0(
#126840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#126890000000
0$
0)
#126900000000
1"
1'
b0 +
b0 1
#126950000000
0"
0'
#126960000000
1#
1(
b101111101100100 +
b101111101100100 1
#127010000000
0#
0(
#127020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#127070000000
0$
0)
#127080000000
1"
1'
b0 +
b0 1
#127130000000
0"
0'
#127140000000
1#
1(
b101111101100100 +
b101111101100100 1
#127190000000
0#
0(
#127200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#127250000000
0$
0)
#127260000000
1"
1'
b0 +
b0 1
#127310000000
0"
0'
#127320000000
1#
1(
b101111101100100 +
b101111101100100 1
#127370000000
0#
0(
#127380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#127430000000
0$
0)
#127440000000
1"
1'
b0 +
b0 1
#127490000000
0"
0'
#127500000000
1#
1(
b101111101100100 +
b101111101100100 1
#127550000000
0#
0(
#127560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#127610000000
0$
0)
#127620000000
1"
1'
b0 +
b0 1
#127670000000
0"
0'
#127680000000
1#
1(
b101111101100100 +
b101111101100100 1
#127730000000
0#
0(
#127740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#127790000000
0$
0)
#127800000000
1"
1'
b0 +
b0 1
#127850000000
0"
0'
#127860000000
1#
1(
b101111101100100 +
b101111101100100 1
#127910000000
0#
0(
#127920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#127970000000
0$
0)
#127980000000
1"
1'
b0 +
b0 1
#128030000000
0"
0'
#128040000000
1#
1(
b101111101100100 +
b101111101100100 1
#128090000000
0#
0(
#128100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#128150000000
0$
0)
#128160000000
1"
1'
b0 +
b0 1
#128210000000
0"
0'
#128220000000
1#
1(
b101111101100100 +
b101111101100100 1
#128270000000
0#
0(
#128280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#128330000000
0$
0)
#128340000000
1"
1'
b0 +
b0 1
#128390000000
0"
0'
#128400000000
1#
1(
b101111101100100 +
b101111101100100 1
#128450000000
0#
0(
#128460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#128510000000
0$
0)
#128520000000
1"
1'
b0 +
b0 1
#128570000000
0"
0'
#128580000000
1#
1(
b101111101100100 +
b101111101100100 1
#128630000000
0#
0(
#128640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#128690000000
0$
0)
#128700000000
1"
1'
b0 +
b0 1
#128750000000
0"
0'
#128760000000
1#
1(
b101111101100100 +
b101111101100100 1
#128810000000
0#
0(
#128820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#128870000000
0$
0)
#128880000000
1"
1'
b0 +
b0 1
#128930000000
0"
0'
#128940000000
1#
1(
b101111101100100 +
b101111101100100 1
#128990000000
0#
0(
#129000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#129050000000
0$
0)
#129060000000
1"
1'
b0 +
b0 1
#129110000000
0"
0'
#129120000000
1#
1(
b101111101100100 +
b101111101100100 1
#129170000000
0#
0(
#129180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#129230000000
0$
0)
#129240000000
1"
1'
b0 +
b0 1
#129290000000
0"
0'
#129300000000
1#
1(
b101111101100100 +
b101111101100100 1
#129350000000
0#
0(
#129360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#129410000000
0$
0)
#129420000000
1"
1'
b0 +
b0 1
#129470000000
0"
0'
#129480000000
1#
1(
b101111101100100 +
b101111101100100 1
#129530000000
0#
0(
#129540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#129590000000
0$
0)
#129600000000
1"
1'
b0 +
b0 1
#129650000000
0"
0'
#129660000000
1#
1(
b101111101100100 +
b101111101100100 1
#129710000000
0#
0(
#129720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#129770000000
0$
0)
#129780000000
1"
1'
b0 +
b0 1
#129830000000
0"
0'
#129840000000
1#
1(
b101111101100100 +
b101111101100100 1
#129890000000
0#
0(
#129900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#129950000000
0$
0)
#129960000000
1"
1'
b0 +
b0 1
#130010000000
0"
0'
#130020000000
1#
1(
b101111101100100 +
b101111101100100 1
#130070000000
0#
0(
#130080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#130130000000
0$
0)
#130140000000
1"
1'
b0 +
b0 1
#130190000000
0"
0'
#130200000000
1#
1(
b101111101100100 +
b101111101100100 1
#130250000000
0#
0(
#130260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#130310000000
0$
0)
#130320000000
1"
1'
b0 +
b0 1
#130370000000
0"
0'
#130380000000
1#
1(
b101111101100100 +
b101111101100100 1
#130430000000
0#
0(
#130440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#130490000000
0$
0)
#130500000000
1"
1'
b0 +
b0 1
#130550000000
0"
0'
#130560000000
1#
1(
b101111101100100 +
b101111101100100 1
#130610000000
0#
0(
#130620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#130670000000
0$
0)
#130680000000
1"
1'
b0 +
b0 1
#130730000000
0"
0'
#130740000000
1#
1(
b101111101100100 +
b101111101100100 1
#130790000000
0#
0(
#130800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#130850000000
0$
0)
#130860000000
1"
1'
b0 +
b0 1
#130910000000
0"
0'
#130920000000
1#
1(
b101111101100100 +
b101111101100100 1
#130970000000
0#
0(
#130980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#131030000000
0$
0)
#131040000000
1"
1'
b0 +
b0 1
#131090000000
0"
0'
#131100000000
1#
1(
b101111101100100 +
b101111101100100 1
#131150000000
0#
0(
#131160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#131210000000
0$
0)
#131220000000
1"
1'
b0 +
b0 1
#131270000000
0"
0'
#131280000000
1#
1(
b101111101100100 +
b101111101100100 1
#131330000000
0#
0(
#131340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#131390000000
0$
0)
#131400000000
1"
1'
b0 +
b0 1
#131450000000
0"
0'
#131460000000
1#
1(
b101111101100100 +
b101111101100100 1
#131510000000
0#
0(
#131520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#131570000000
0$
0)
#131580000000
1"
1'
b0 +
b0 1
#131630000000
0"
0'
#131640000000
1#
1(
b101111101100100 +
b101111101100100 1
#131690000000
0#
0(
#131700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#131750000000
0$
0)
#131760000000
1"
1'
b0 +
b0 1
#131810000000
0"
0'
#131820000000
1#
1(
b101111101100100 +
b101111101100100 1
#131870000000
0#
0(
#131880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#131930000000
0$
0)
#131940000000
1"
1'
b0 +
b0 1
#131990000000
0"
0'
#132000000000
1#
1(
b101111101100100 +
b101111101100100 1
#132050000000
0#
0(
#132060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#132110000000
0$
0)
#132120000000
1"
1'
b0 +
b0 1
#132170000000
0"
0'
#132180000000
1#
1(
b101111101100100 +
b101111101100100 1
#132230000000
0#
0(
#132240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#132290000000
0$
0)
#132300000000
1"
1'
b0 +
b0 1
#132350000000
0"
0'
#132360000000
1#
1(
b101111101100100 +
b101111101100100 1
#132410000000
0#
0(
#132420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#132470000000
0$
0)
#132480000000
1"
1'
b0 +
b0 1
#132530000000
0"
0'
#132540000000
1#
1(
b101111101100100 +
b101111101100100 1
#132590000000
0#
0(
#132600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#132650000000
0$
0)
#132660000000
1"
1'
b0 +
b0 1
#132710000000
0"
0'
#132720000000
1#
1(
b101111101100100 +
b101111101100100 1
#132770000000
0#
0(
#132780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#132830000000
0$
0)
#132840000000
1"
1'
b0 +
b0 1
#132890000000
0"
0'
#132900000000
1#
1(
b101111101100100 +
b101111101100100 1
#132950000000
0#
0(
#132960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#133010000000
0$
0)
#133020000000
1"
1'
b0 +
b0 1
#133070000000
0"
0'
#133080000000
1#
1(
b101111101100100 +
b101111101100100 1
#133130000000
0#
0(
#133140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#133190000000
0$
0)
#133200000000
1"
1'
b0 +
b0 1
#133250000000
0"
0'
#133260000000
1#
1(
b101111101100100 +
b101111101100100 1
#133310000000
0#
0(
#133320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#133370000000
0$
0)
#133380000000
1"
1'
b0 +
b0 1
#133430000000
0"
0'
#133440000000
1#
1(
b101111101100100 +
b101111101100100 1
#133490000000
0#
0(
#133500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#133550000000
0$
0)
#133560000000
1"
1'
b0 +
b0 1
#133610000000
0"
0'
#133620000000
1#
1(
b101111101100100 +
b101111101100100 1
#133670000000
0#
0(
#133680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#133730000000
0$
0)
#133740000000
1"
1'
b0 +
b0 1
#133790000000
0"
0'
#133800000000
1#
1(
b101111101100100 +
b101111101100100 1
#133850000000
0#
0(
#133860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#133910000000
0$
0)
#133920000000
1"
1'
b0 +
b0 1
#133970000000
0"
0'
#133980000000
1#
1(
b101111101100100 +
b101111101100100 1
#134030000000
0#
0(
#134040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#134090000000
0$
0)
#134100000000
1"
1'
b0 +
b0 1
#134150000000
0"
0'
#134160000000
1#
1(
b101111101100100 +
b101111101100100 1
#134210000000
0#
0(
#134220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#134270000000
0$
0)
#134280000000
1"
1'
b0 +
b0 1
#134330000000
0"
0'
#134340000000
1#
1(
b101111101100100 +
b101111101100100 1
#134390000000
0#
0(
#134400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#134450000000
0$
0)
#134460000000
1"
1'
b0 +
b0 1
#134510000000
0"
0'
#134520000000
1#
1(
b101111101100100 +
b101111101100100 1
#134570000000
0#
0(
#134580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#134630000000
0$
0)
#134640000000
1"
1'
b0 +
b0 1
#134690000000
0"
0'
#134700000000
1#
1(
b101111101100100 +
b101111101100100 1
#134750000000
0#
0(
#134760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#134810000000
0$
0)
#134820000000
1"
1'
b0 +
b0 1
#134870000000
0"
0'
#134880000000
1#
1(
b101111101100100 +
b101111101100100 1
#134930000000
0#
0(
#134940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#134990000000
0$
0)
#135000000000
1"
1'
b0 +
b0 1
#135050000000
0"
0'
#135060000000
1#
1(
b101111101100100 +
b101111101100100 1
#135110000000
0#
0(
#135120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#135170000000
0$
0)
#135180000000
1"
1'
b0 +
b0 1
#135230000000
0"
0'
#135240000000
1#
1(
b101111101100100 +
b101111101100100 1
#135290000000
0#
0(
#135300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#135350000000
0$
0)
#135360000000
1"
1'
b0 +
b0 1
#135410000000
0"
0'
#135420000000
1#
1(
b101111101100100 +
b101111101100100 1
#135470000000
0#
0(
#135480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#135530000000
0$
0)
#135540000000
1"
1'
b0 +
b0 1
#135590000000
0"
0'
#135600000000
1#
1(
b101111101100100 +
b101111101100100 1
#135650000000
0#
0(
#135660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#135710000000
0$
0)
#135720000000
1"
1'
b0 +
b0 1
#135770000000
0"
0'
#135780000000
1#
1(
b101111101100100 +
b101111101100100 1
#135830000000
0#
0(
#135840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#135890000000
0$
0)
#135900000000
1"
1'
b0 +
b0 1
#135950000000
0"
0'
#135960000000
1#
1(
b101111101100100 +
b101111101100100 1
#136010000000
0#
0(
#136020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#136070000000
0$
0)
#136080000000
1"
1'
b0 +
b0 1
#136130000000
0"
0'
#136140000000
1#
1(
b101111101100100 +
b101111101100100 1
#136190000000
0#
0(
#136200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#136250000000
0$
0)
#136260000000
1"
1'
b0 +
b0 1
#136310000000
0"
0'
#136320000000
1#
1(
b101111101100100 +
b101111101100100 1
#136370000000
0#
0(
#136380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#136430000000
0$
0)
#136440000000
1"
1'
b0 +
b0 1
#136490000000
0"
0'
#136500000000
1#
1(
b101111101100100 +
b101111101100100 1
#136550000000
0#
0(
#136560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#136610000000
0$
0)
#136620000000
1"
1'
b0 +
b0 1
#136670000000
0"
0'
#136680000000
1#
1(
b101111101100100 +
b101111101100100 1
#136730000000
0#
0(
#136740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#136790000000
0$
0)
#136800000000
1"
1'
b0 +
b0 1
#136850000000
0"
0'
#136860000000
1#
1(
b101111101100100 +
b101111101100100 1
#136910000000
0#
0(
#136920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#136970000000
0$
0)
#136980000000
1"
1'
b0 +
b0 1
#137030000000
0"
0'
#137040000000
1#
1(
b101111101100100 +
b101111101100100 1
#137090000000
0#
0(
#137100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#137150000000
0$
0)
#137160000000
1"
1'
b0 +
b0 1
#137210000000
0"
0'
#137220000000
1#
1(
b101111101100100 +
b101111101100100 1
#137270000000
0#
0(
#137280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#137330000000
0$
0)
#137340000000
1"
1'
b0 +
b0 1
#137390000000
0"
0'
#137400000000
1#
1(
b101111101100100 +
b101111101100100 1
#137450000000
0#
0(
#137460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#137510000000
0$
0)
#137520000000
1"
1'
b0 +
b0 1
#137570000000
0"
0'
#137580000000
1#
1(
b101111101100100 +
b101111101100100 1
#137630000000
0#
0(
#137640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#137690000000
0$
0)
#137700000000
1"
1'
b0 +
b0 1
#137750000000
0"
0'
#137760000000
1#
1(
b101111101100100 +
b101111101100100 1
#137810000000
0#
0(
#137820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#137870000000
0$
0)
#137880000000
1"
1'
b0 +
b0 1
#137930000000
0"
0'
#137940000000
1#
1(
b101111101100100 +
b101111101100100 1
#137990000000
0#
0(
#138000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#138050000000
0$
0)
#138060000000
1"
1'
b0 +
b0 1
#138110000000
0"
0'
#138120000000
1#
1(
b101111101100100 +
b101111101100100 1
#138170000000
0#
0(
#138180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#138230000000
0$
0)
#138240000000
1"
1'
b0 +
b0 1
#138290000000
0"
0'
#138300000000
1#
1(
b101111101100100 +
b101111101100100 1
#138350000000
0#
0(
#138360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#138410000000
0$
0)
#138420000000
1"
1'
b0 +
b0 1
#138470000000
0"
0'
#138480000000
1#
1(
b101111101100100 +
b101111101100100 1
#138530000000
0#
0(
#138540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#138590000000
0$
0)
#138600000000
1"
1'
b0 +
b0 1
#138650000000
0"
0'
#138660000000
1#
1(
b101111101100100 +
b101111101100100 1
#138710000000
0#
0(
#138720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#138770000000
0$
0)
#138780000000
1"
1'
b0 +
b0 1
#138830000000
0"
0'
#138840000000
1#
1(
b101111101100100 +
b101111101100100 1
#138890000000
0#
0(
#138900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#138950000000
0$
0)
#138960000000
1"
1'
b0 +
b0 1
#139010000000
0"
0'
#139020000000
1#
1(
b101111101100100 +
b101111101100100 1
#139070000000
0#
0(
#139080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#139130000000
0$
0)
#139140000000
1"
1'
b0 +
b0 1
#139190000000
0"
0'
#139200000000
1#
1(
b101111101100100 +
b101111101100100 1
#139250000000
0#
0(
#139260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#139310000000
0$
0)
#139320000000
1"
1'
b0 +
b0 1
#139370000000
0"
0'
#139380000000
1#
1(
b101111101100100 +
b101111101100100 1
#139430000000
0#
0(
#139440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#139490000000
0$
0)
#139500000000
1"
1'
b0 +
b0 1
#139550000000
0"
0'
#139560000000
1#
1(
b101111101100100 +
b101111101100100 1
#139610000000
0#
0(
#139620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#139670000000
0$
0)
#139680000000
1"
1'
b0 +
b0 1
#139730000000
0"
0'
#139740000000
1#
1(
b101111101100100 +
b101111101100100 1
#139790000000
0#
0(
#139800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#139850000000
0$
0)
#139860000000
1"
1'
b0 +
b0 1
#139910000000
0"
0'
#139920000000
1#
1(
b101111101100100 +
b101111101100100 1
#139970000000
0#
0(
#139980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#140030000000
0$
0)
#140040000000
1"
1'
b0 +
b0 1
#140090000000
0"
0'
#140100000000
1#
1(
b101111101100100 +
b101111101100100 1
#140150000000
0#
0(
#140160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#140210000000
0$
0)
#140220000000
1"
1'
b0 +
b0 1
#140270000000
0"
0'
#140280000000
1#
1(
b101111101100100 +
b101111101100100 1
#140330000000
0#
0(
#140340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#140390000000
0$
0)
#140400000000
1"
1'
b0 +
b0 1
#140450000000
0"
0'
#140460000000
1#
1(
b101111101100100 +
b101111101100100 1
#140510000000
0#
0(
#140520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#140570000000
0$
0)
#140580000000
1"
1'
b0 +
b0 1
#140630000000
0"
0'
#140640000000
1#
1(
b101111101100100 +
b101111101100100 1
#140690000000
0#
0(
#140700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#140750000000
0$
0)
#140760000000
1"
1'
b0 +
b0 1
#140810000000
0"
0'
#140820000000
1#
1(
b101111101100100 +
b101111101100100 1
#140870000000
0#
0(
#140880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#140930000000
0$
0)
#140940000000
1"
1'
b0 +
b0 1
#140990000000
0"
0'
#141000000000
1#
1(
b101111101100100 +
b101111101100100 1
#141050000000
0#
0(
#141060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#141110000000
0$
0)
#141120000000
1"
1'
b0 +
b0 1
#141170000000
0"
0'
#141180000000
1#
1(
b101111101100100 +
b101111101100100 1
#141230000000
0#
0(
#141240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#141290000000
0$
0)
#141300000000
1"
1'
b0 +
b0 1
#141350000000
0"
0'
#141360000000
1#
1(
b101111101100100 +
b101111101100100 1
#141410000000
0#
0(
#141420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#141470000000
0$
0)
#141480000000
1"
1'
b0 +
b0 1
#141530000000
0"
0'
#141540000000
1#
1(
b101111101100100 +
b101111101100100 1
#141590000000
0#
0(
#141600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#141650000000
0$
0)
#141660000000
1"
1'
b0 +
b0 1
#141710000000
0"
0'
#141720000000
1#
1(
b101111101100100 +
b101111101100100 1
#141770000000
0#
0(
#141780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#141830000000
0$
0)
#141840000000
1"
1'
b0 +
b0 1
#141890000000
0"
0'
#141900000000
1#
1(
b101111101100100 +
b101111101100100 1
#141950000000
0#
0(
#141960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#142010000000
0$
0)
#142020000000
1"
1'
b0 +
b0 1
#142070000000
0"
0'
#142080000000
1#
1(
b101111101100100 +
b101111101100100 1
#142130000000
0#
0(
#142140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#142190000000
0$
0)
#142200000000
1"
1'
b0 +
b0 1
#142250000000
0"
0'
#142260000000
1#
1(
b101111101100100 +
b101111101100100 1
#142310000000
0#
0(
#142320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#142370000000
0$
0)
#142380000000
1"
1'
b0 +
b0 1
#142430000000
0"
0'
#142440000000
1#
1(
b101111101100100 +
b101111101100100 1
#142490000000
0#
0(
#142500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#142550000000
0$
0)
#142560000000
1"
1'
b0 +
b0 1
#142610000000
0"
0'
#142620000000
1#
1(
b101111101100100 +
b101111101100100 1
#142670000000
0#
0(
#142680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#142730000000
0$
0)
#142740000000
1"
1'
b0 +
b0 1
#142790000000
0"
0'
#142800000000
1#
1(
b101111101100100 +
b101111101100100 1
#142850000000
0#
0(
#142860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#142910000000
0$
0)
#142920000000
1"
1'
b0 +
b0 1
#142970000000
0"
0'
#142980000000
1#
1(
b101111101100100 +
b101111101100100 1
#143030000000
0#
0(
#143040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#143090000000
0$
0)
#143100000000
1"
1'
b0 +
b0 1
#143150000000
0"
0'
#143160000000
1#
1(
b101111101100100 +
b101111101100100 1
#143210000000
0#
0(
#143220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#143270000000
0$
0)
#143280000000
1"
1'
b0 +
b0 1
#143330000000
0"
0'
#143340000000
1#
1(
b101111101100100 +
b101111101100100 1
#143390000000
0#
0(
#143400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#143450000000
0$
0)
#143460000000
1"
1'
b0 +
b0 1
#143510000000
0"
0'
#143520000000
1#
1(
b101111101100100 +
b101111101100100 1
#143570000000
0#
0(
#143580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#143630000000
0$
0)
#143640000000
1"
1'
b0 +
b0 1
#143690000000
0"
0'
#143700000000
1#
1(
b101111101100100 +
b101111101100100 1
#143750000000
0#
0(
#143760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#143810000000
0$
0)
#143820000000
1"
1'
b0 +
b0 1
#143870000000
0"
0'
#143880000000
1#
1(
b101111101100100 +
b101111101100100 1
#143930000000
0#
0(
#143940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#143990000000
0$
0)
#144000000000
1"
1'
b0 +
b0 1
#144050000000
0"
0'
#144060000000
1#
1(
b101111101100100 +
b101111101100100 1
#144110000000
0#
0(
#144120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#144170000000
0$
0)
#144180000000
1"
1'
b0 +
b0 1
#144230000000
0"
0'
#144240000000
1#
1(
b101111101100100 +
b101111101100100 1
#144290000000
0#
0(
#144300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#144350000000
0$
0)
#144360000000
1"
1'
b0 +
b0 1
#144410000000
0"
0'
#144420000000
1#
1(
b101111101100100 +
b101111101100100 1
#144470000000
0#
0(
#144480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#144530000000
0$
0)
#144540000000
1"
1'
b0 +
b0 1
#144590000000
0"
0'
#144600000000
1#
1(
b101111101100100 +
b101111101100100 1
#144650000000
0#
0(
#144660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#144710000000
0$
0)
#144720000000
1"
1'
b0 +
b0 1
#144770000000
0"
0'
#144780000000
1#
1(
b101111101100100 +
b101111101100100 1
#144830000000
0#
0(
#144840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#144890000000
0$
0)
#144900000000
1"
1'
b0 +
b0 1
#144950000000
0"
0'
#144960000000
1#
1(
b101111101100100 +
b101111101100100 1
#145010000000
0#
0(
#145020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#145070000000
0$
0)
#145080000000
1"
1'
b0 +
b0 1
#145130000000
0"
0'
#145140000000
1#
1(
b101111101100100 +
b101111101100100 1
#145190000000
0#
0(
#145200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#145250000000
0$
0)
#145260000000
1"
1'
b0 +
b0 1
#145310000000
0"
0'
#145320000000
1#
1(
b101111101100100 +
b101111101100100 1
#145370000000
0#
0(
#145380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#145430000000
0$
0)
#145440000000
1"
1'
b0 +
b0 1
#145490000000
0"
0'
#145500000000
1#
1(
b101111101100100 +
b101111101100100 1
#145550000000
0#
0(
#145560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#145610000000
0$
0)
#145620000000
1"
1'
b0 +
b0 1
#145670000000
0"
0'
#145680000000
1#
1(
b101111101100100 +
b101111101100100 1
#145730000000
0#
0(
#145740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#145790000000
0$
0)
#145800000000
1"
1'
b0 +
b0 1
#145850000000
0"
0'
#145860000000
1#
1(
b101111101100100 +
b101111101100100 1
#145910000000
0#
0(
#145920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#145970000000
0$
0)
#145980000000
1"
1'
b0 +
b0 1
#146030000000
0"
0'
#146040000000
1#
1(
b101111101100100 +
b101111101100100 1
#146090000000
0#
0(
#146100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#146150000000
0$
0)
#146160000000
1"
1'
b0 +
b0 1
#146210000000
0"
0'
#146220000000
1#
1(
b101111101100100 +
b101111101100100 1
#146270000000
0#
0(
#146280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#146330000000
0$
0)
#146340000000
1"
1'
b0 +
b0 1
#146390000000
0"
0'
#146400000000
1#
1(
b101111101100100 +
b101111101100100 1
#146450000000
0#
0(
#146460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#146510000000
0$
0)
#146520000000
1"
1'
b0 +
b0 1
#146570000000
0"
0'
#146580000000
1#
1(
b101111101100100 +
b101111101100100 1
#146630000000
0#
0(
#146640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#146690000000
0$
0)
#146700000000
1"
1'
b0 +
b0 1
#146750000000
0"
0'
#146760000000
1#
1(
b101111101100100 +
b101111101100100 1
#146810000000
0#
0(
#146820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#146870000000
0$
0)
#146880000000
1"
1'
b0 +
b0 1
#146930000000
0"
0'
#146940000000
1#
1(
b101111101100100 +
b101111101100100 1
#146990000000
0#
0(
#147000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#147050000000
0$
0)
#147060000000
1"
1'
b0 +
b0 1
#147110000000
0"
0'
#147120000000
1#
1(
b101111101100100 +
b101111101100100 1
#147170000000
0#
0(
#147180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#147230000000
0$
0)
#147240000000
1"
1'
b0 +
b0 1
#147290000000
0"
0'
#147300000000
1#
1(
b101111101100100 +
b101111101100100 1
#147350000000
0#
0(
#147360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#147410000000
0$
0)
#147420000000
1"
1'
b0 +
b0 1
#147470000000
0"
0'
#147480000000
1#
1(
b101111101100100 +
b101111101100100 1
#147530000000
0#
0(
#147540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#147590000000
0$
0)
#147600000000
1"
1'
b0 +
b0 1
#147650000000
0"
0'
#147660000000
1#
1(
b101111101100100 +
b101111101100100 1
#147710000000
0#
0(
#147720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#147770000000
0$
0)
#147780000000
1"
1'
b0 +
b0 1
#147830000000
0"
0'
#147840000000
1#
1(
b101111101100100 +
b101111101100100 1
#147890000000
0#
0(
#147900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#147950000000
0$
0)
#147960000000
1"
1'
b0 +
b0 1
#148010000000
0"
0'
#148020000000
1#
1(
b101111101100100 +
b101111101100100 1
#148070000000
0#
0(
#148080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#148130000000
0$
0)
#148140000000
1"
1'
b0 +
b0 1
#148190000000
0"
0'
#148200000000
1#
1(
b101111101100100 +
b101111101100100 1
#148250000000
0#
0(
#148260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#148310000000
0$
0)
#148320000000
1"
1'
b0 +
b0 1
#148370000000
0"
0'
#148380000000
1#
1(
b101111101100100 +
b101111101100100 1
#148430000000
0#
0(
#148440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#148490000000
0$
0)
#148500000000
1"
1'
b0 +
b0 1
#148550000000
0"
0'
#148560000000
1#
1(
b101111101100100 +
b101111101100100 1
#148610000000
0#
0(
#148620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#148670000000
0$
0)
#148680000000
1"
1'
b0 +
b0 1
#148730000000
0"
0'
#148740000000
1#
1(
b101111101100100 +
b101111101100100 1
#148790000000
0#
0(
#148800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#148850000000
0$
0)
#148860000000
1"
1'
b0 +
b0 1
#148910000000
0"
0'
#148920000000
1#
1(
b101111101100100 +
b101111101100100 1
#148970000000
0#
0(
#148980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#149030000000
0$
0)
#149040000000
1"
1'
b0 +
b0 1
#149090000000
0"
0'
#149100000000
1#
1(
b101111101100100 +
b101111101100100 1
#149150000000
0#
0(
#149160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#149210000000
0$
0)
#149220000000
1"
1'
b0 +
b0 1
#149270000000
0"
0'
#149280000000
1#
1(
b101111101100100 +
b101111101100100 1
#149330000000
0#
0(
#149340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#149390000000
0$
0)
#149400000000
1"
1'
b0 +
b0 1
#149450000000
0"
0'
#149460000000
1#
1(
b101111101100100 +
b101111101100100 1
#149510000000
0#
0(
#149520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#149570000000
0$
0)
#149580000000
1"
1'
b0 +
b0 1
#149630000000
0"
0'
#149640000000
1#
1(
b101111101100100 +
b101111101100100 1
#149690000000
0#
0(
#149700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#149750000000
0$
0)
#149760000000
1"
1'
b0 +
b0 1
#149810000000
0"
0'
#149820000000
1#
1(
b101111101100100 +
b101111101100100 1
#149870000000
0#
0(
#149880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#149930000000
0$
0)
#149940000000
1"
1'
b0 +
b0 1
#149990000000
0"
0'
#150000000000
1#
1(
b101111101100100 +
b101111101100100 1
#150050000000
0#
0(
#150060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#150110000000
0$
0)
#150120000000
1"
1'
b0 +
b0 1
#150170000000
0"
0'
#150180000000
1#
1(
b101111101100100 +
b101111101100100 1
#150230000000
0#
0(
#150240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#150290000000
0$
0)
#150300000000
1"
1'
b0 +
b0 1
#150350000000
0"
0'
#150360000000
1#
1(
b101111101100100 +
b101111101100100 1
#150410000000
0#
0(
#150420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#150470000000
0$
0)
#150480000000
1"
1'
b0 +
b0 1
#150530000000
0"
0'
#150540000000
1#
1(
b101111101100100 +
b101111101100100 1
#150590000000
0#
0(
#150600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#150650000000
0$
0)
#150660000000
1"
1'
b0 +
b0 1
#150710000000
0"
0'
#150720000000
1#
1(
b101111101100100 +
b101111101100100 1
#150770000000
0#
0(
#150780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#150830000000
0$
0)
#150840000000
1"
1'
b0 +
b0 1
#150890000000
0"
0'
#150900000000
1#
1(
b101111101100100 +
b101111101100100 1
#150950000000
0#
0(
#150960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#151010000000
0$
0)
#151020000000
1"
1'
b0 +
b0 1
#151070000000
0"
0'
#151080000000
1#
1(
b101111101100100 +
b101111101100100 1
#151130000000
0#
0(
#151140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#151190000000
0$
0)
#151200000000
1"
1'
b0 +
b0 1
#151250000000
0"
0'
#151260000000
1#
1(
b101111101100100 +
b101111101100100 1
#151310000000
0#
0(
#151320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#151370000000
0$
0)
#151380000000
1"
1'
b0 +
b0 1
#151430000000
0"
0'
#151440000000
1#
1(
b101111101100100 +
b101111101100100 1
#151490000000
0#
0(
#151500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#151550000000
0$
0)
#151560000000
1"
1'
b0 +
b0 1
#151610000000
0"
0'
#151620000000
1#
1(
b101111101100100 +
b101111101100100 1
#151670000000
0#
0(
#151680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#151730000000
0$
0)
#151740000000
1"
1'
b0 +
b0 1
#151790000000
0"
0'
#151800000000
1#
1(
b101111101100100 +
b101111101100100 1
#151850000000
0#
0(
#151860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#151910000000
0$
0)
#151920000000
1"
1'
b0 +
b0 1
#151970000000
0"
0'
#151980000000
1#
1(
b101111101100100 +
b101111101100100 1
#152030000000
0#
0(
#152040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#152090000000
0$
0)
#152100000000
1"
1'
b0 +
b0 1
#152150000000
0"
0'
#152160000000
1#
1(
b101111101100100 +
b101111101100100 1
#152210000000
0#
0(
#152220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#152270000000
0$
0)
#152280000000
1"
1'
b0 +
b0 1
#152330000000
0"
0'
#152340000000
1#
1(
b101111101100100 +
b101111101100100 1
#152390000000
0#
0(
#152400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#152450000000
0$
0)
#152460000000
1"
1'
b0 +
b0 1
#152510000000
0"
0'
#152520000000
1#
1(
b101111101100100 +
b101111101100100 1
#152570000000
0#
0(
#152580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#152630000000
0$
0)
#152640000000
1"
1'
b0 +
b0 1
#152690000000
0"
0'
#152700000000
1#
1(
b101111101100100 +
b101111101100100 1
#152750000000
0#
0(
#152760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#152810000000
0$
0)
#152820000000
1"
1'
b0 +
b0 1
#152870000000
0"
0'
#152880000000
1#
1(
b101111101100100 +
b101111101100100 1
#152930000000
0#
0(
#152940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#152990000000
0$
0)
#153000000000
1"
1'
b0 +
b0 1
#153050000000
0"
0'
#153060000000
1#
1(
b101111101100100 +
b101111101100100 1
#153110000000
0#
0(
#153120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#153170000000
0$
0)
#153180000000
1"
1'
b0 +
b0 1
#153230000000
0"
0'
#153240000000
1#
1(
b101111101100100 +
b101111101100100 1
#153290000000
0#
0(
#153300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#153350000000
0$
0)
#153360000000
1"
1'
b0 +
b0 1
#153410000000
0"
0'
#153420000000
1#
1(
b101111101100100 +
b101111101100100 1
#153470000000
0#
0(
#153480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#153530000000
0$
0)
#153540000000
1"
1'
b0 +
b0 1
#153590000000
0"
0'
#153600000000
1#
1(
b101111101100100 +
b101111101100100 1
#153650000000
0#
0(
#153660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#153710000000
0$
0)
#153720000000
1"
1'
b0 +
b0 1
#153770000000
0"
0'
#153780000000
1#
1(
b101111101100100 +
b101111101100100 1
#153830000000
0#
0(
#153840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#153890000000
0$
0)
#153900000000
1"
1'
b0 +
b0 1
#153950000000
0"
0'
#153960000000
1#
1(
b101111101100100 +
b101111101100100 1
#154010000000
0#
0(
#154020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#154070000000
0$
0)
#154080000000
1"
1'
b0 +
b0 1
#154130000000
0"
0'
#154140000000
1#
1(
b101111101100100 +
b101111101100100 1
#154190000000
0#
0(
#154200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#154250000000
0$
0)
#154260000000
1"
1'
b0 +
b0 1
#154310000000
0"
0'
#154320000000
1#
1(
b101111101100100 +
b101111101100100 1
#154370000000
0#
0(
#154380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#154430000000
0$
0)
#154440000000
1"
1'
b0 +
b0 1
#154490000000
0"
0'
#154500000000
1#
1(
b101111101100100 +
b101111101100100 1
#154550000000
0#
0(
#154560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#154610000000
0$
0)
#154620000000
1"
1'
b0 +
b0 1
#154670000000
0"
0'
#154680000000
1#
1(
b101111101100100 +
b101111101100100 1
#154730000000
0#
0(
#154740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#154790000000
0$
0)
#154800000000
1"
1'
b0 +
b0 1
#154850000000
0"
0'
#154860000000
1#
1(
b101111101100100 +
b101111101100100 1
#154910000000
0#
0(
#154920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#154970000000
0$
0)
#154980000000
1"
1'
b0 +
b0 1
#155030000000
0"
0'
#155040000000
1#
1(
b101111101100100 +
b101111101100100 1
#155090000000
0#
0(
#155100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#155150000000
0$
0)
#155160000000
1"
1'
b0 +
b0 1
#155210000000
0"
0'
#155220000000
1#
1(
b101111101100100 +
b101111101100100 1
#155270000000
0#
0(
#155280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#155330000000
0$
0)
#155340000000
1"
1'
b0 +
b0 1
#155390000000
0"
0'
#155400000000
1#
1(
b101111101100100 +
b101111101100100 1
#155450000000
0#
0(
#155460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#155510000000
0$
0)
#155520000000
1"
1'
b0 +
b0 1
#155570000000
0"
0'
#155580000000
1#
1(
b101111101100100 +
b101111101100100 1
#155630000000
0#
0(
#155640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#155690000000
0$
0)
#155700000000
1"
1'
b0 +
b0 1
#155750000000
0"
0'
#155760000000
1#
1(
b101111101100100 +
b101111101100100 1
#155810000000
0#
0(
#155820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#155870000000
0$
0)
#155880000000
1"
1'
b0 +
b0 1
#155930000000
0"
0'
#155940000000
1#
1(
b101111101100100 +
b101111101100100 1
#155990000000
0#
0(
#156000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#156050000000
0$
0)
#156060000000
1"
1'
b0 +
b0 1
#156110000000
0"
0'
#156120000000
1#
1(
b101111101100100 +
b101111101100100 1
#156170000000
0#
0(
#156180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#156230000000
0$
0)
#156240000000
1"
1'
b0 +
b0 1
#156290000000
0"
0'
#156300000000
1#
1(
b101111101100100 +
b101111101100100 1
#156350000000
0#
0(
#156360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#156410000000
0$
0)
#156420000000
1"
1'
b0 +
b0 1
#156470000000
0"
0'
#156480000000
1#
1(
b101111101100100 +
b101111101100100 1
#156530000000
0#
0(
#156540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#156590000000
0$
0)
#156600000000
1"
1'
b0 +
b0 1
#156650000000
0"
0'
#156660000000
1#
1(
b101111101100100 +
b101111101100100 1
#156710000000
0#
0(
#156720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#156770000000
0$
0)
#156780000000
1"
1'
b0 +
b0 1
#156830000000
0"
0'
#156840000000
1#
1(
b101111101100100 +
b101111101100100 1
#156890000000
0#
0(
#156900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#156950000000
0$
0)
#156960000000
1"
1'
b0 +
b0 1
#157010000000
0"
0'
#157020000000
1#
1(
b101111101100100 +
b101111101100100 1
#157070000000
0#
0(
#157080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#157130000000
0$
0)
#157140000000
1"
1'
b0 +
b0 1
#157190000000
0"
0'
#157200000000
1#
1(
b101111101100100 +
b101111101100100 1
#157250000000
0#
0(
#157260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#157310000000
0$
0)
#157320000000
1"
1'
b0 +
b0 1
#157370000000
0"
0'
#157380000000
1#
1(
b101111101100100 +
b101111101100100 1
#157430000000
0#
0(
#157440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#157490000000
0$
0)
#157500000000
1"
1'
b0 +
b0 1
#157550000000
0"
0'
#157560000000
1#
1(
b101111101100100 +
b101111101100100 1
#157610000000
0#
0(
#157620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#157670000000
0$
0)
#157680000000
1"
1'
b0 +
b0 1
#157730000000
0"
0'
#157740000000
1#
1(
b101111101100100 +
b101111101100100 1
#157790000000
0#
0(
#157800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#157850000000
0$
0)
#157860000000
1"
1'
b0 +
b0 1
#157910000000
0"
0'
#157920000000
1#
1(
b101111101100100 +
b101111101100100 1
#157970000000
0#
0(
#157980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#158030000000
0$
0)
#158040000000
1"
1'
b0 +
b0 1
#158090000000
0"
0'
#158100000000
1#
1(
b101111101100100 +
b101111101100100 1
#158150000000
0#
0(
#158160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#158210000000
0$
0)
#158220000000
1"
1'
b0 +
b0 1
#158270000000
0"
0'
#158280000000
1#
1(
b101111101100100 +
b101111101100100 1
#158330000000
0#
0(
#158340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#158390000000
0$
0)
#158400000000
1"
1'
b0 +
b0 1
#158450000000
0"
0'
#158460000000
1#
1(
b101111101100100 +
b101111101100100 1
#158510000000
0#
0(
#158520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#158570000000
0$
0)
#158580000000
1"
1'
b0 +
b0 1
#158630000000
0"
0'
#158640000000
1#
1(
b101111101100100 +
b101111101100100 1
#158690000000
0#
0(
#158700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#158750000000
0$
0)
#158760000000
1"
1'
b0 +
b0 1
#158810000000
0"
0'
#158820000000
1#
1(
b101111101100100 +
b101111101100100 1
#158870000000
0#
0(
#158880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#158930000000
0$
0)
#158940000000
1"
1'
b0 +
b0 1
#158990000000
0"
0'
#159000000000
1#
1(
b101111101100100 +
b101111101100100 1
#159050000000
0#
0(
#159060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#159110000000
0$
0)
#159120000000
1"
1'
b0 +
b0 1
#159170000000
0"
0'
#159180000000
1#
1(
b101111101100100 +
b101111101100100 1
#159230000000
0#
0(
#159240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#159290000000
0$
0)
#159300000000
1"
1'
b0 +
b0 1
#159350000000
0"
0'
#159360000000
1#
1(
b101111101100100 +
b101111101100100 1
#159410000000
0#
0(
#159420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#159470000000
0$
0)
#159480000000
1"
1'
b0 +
b0 1
#159530000000
0"
0'
#159540000000
1#
1(
b101111101100100 +
b101111101100100 1
#159590000000
0#
0(
#159600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#159650000000
0$
0)
#159660000000
1"
1'
b0 +
b0 1
#159710000000
0"
0'
#159720000000
1#
1(
b101111101100100 +
b101111101100100 1
#159770000000
0#
0(
#159780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#159830000000
0$
0)
#159840000000
1"
1'
b0 +
b0 1
#159890000000
0"
0'
#159900000000
1#
1(
b101111101100100 +
b101111101100100 1
#159950000000
0#
0(
#159960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#160010000000
0$
0)
#160020000000
1"
1'
b0 +
b0 1
#160070000000
0"
0'
#160080000000
1#
1(
b101111101100100 +
b101111101100100 1
#160130000000
0#
0(
#160140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#160190000000
0$
0)
#160200000000
1"
1'
b0 +
b0 1
#160250000000
0"
0'
#160260000000
1#
1(
b101111101100100 +
b101111101100100 1
#160310000000
0#
0(
#160320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#160370000000
0$
0)
#160380000000
1"
1'
b0 +
b0 1
#160430000000
0"
0'
#160440000000
1#
1(
b101111101100100 +
b101111101100100 1
#160490000000
0#
0(
#160500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#160550000000
0$
0)
#160560000000
1"
1'
b0 +
b0 1
#160610000000
0"
0'
#160620000000
1#
1(
b101111101100100 +
b101111101100100 1
#160670000000
0#
0(
#160680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#160730000000
0$
0)
#160740000000
1"
1'
b0 +
b0 1
#160790000000
0"
0'
#160800000000
1#
1(
b101111101100100 +
b101111101100100 1
#160850000000
0#
0(
#160860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#160910000000
0$
0)
#160920000000
1"
1'
b0 +
b0 1
#160970000000
0"
0'
#160980000000
1#
1(
b101111101100100 +
b101111101100100 1
#161030000000
0#
0(
#161040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#161090000000
0$
0)
#161100000000
1"
1'
b0 +
b0 1
#161150000000
0"
0'
#161160000000
1#
1(
b101111101100100 +
b101111101100100 1
#161210000000
0#
0(
#161220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#161270000000
0$
0)
#161280000000
1"
1'
b0 +
b0 1
#161330000000
0"
0'
#161340000000
1#
1(
b101111101100100 +
b101111101100100 1
#161390000000
0#
0(
#161400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#161450000000
0$
0)
#161460000000
1"
1'
b0 +
b0 1
#161510000000
0"
0'
#161520000000
1#
1(
b101111101100100 +
b101111101100100 1
#161570000000
0#
0(
#161580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#161630000000
0$
0)
#161640000000
1"
1'
b0 +
b0 1
#161690000000
0"
0'
#161700000000
1#
1(
b101111101100100 +
b101111101100100 1
#161750000000
0#
0(
#161760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#161810000000
0$
0)
#161820000000
1"
1'
b0 +
b0 1
#161870000000
0"
0'
#161880000000
1#
1(
b101111101100100 +
b101111101100100 1
#161930000000
0#
0(
#161940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#161990000000
0$
0)
#162000000000
1"
1'
b0 +
b0 1
#162050000000
0"
0'
#162060000000
1#
1(
b101111101100100 +
b101111101100100 1
#162110000000
0#
0(
#162120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#162170000000
0$
0)
#162180000000
1"
1'
b0 +
b0 1
#162230000000
0"
0'
#162240000000
1#
1(
b101111101100100 +
b101111101100100 1
#162290000000
0#
0(
#162300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#162350000000
0$
0)
#162360000000
1"
1'
b0 +
b0 1
#162410000000
0"
0'
#162420000000
1#
1(
b101111101100100 +
b101111101100100 1
#162470000000
0#
0(
#162480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#162530000000
0$
0)
#162540000000
1"
1'
b0 +
b0 1
#162590000000
0"
0'
#162600000000
1#
1(
b101111101100100 +
b101111101100100 1
#162650000000
0#
0(
#162660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#162710000000
0$
0)
#162720000000
1"
1'
b0 +
b0 1
#162770000000
0"
0'
#162780000000
1#
1(
b101111101100100 +
b101111101100100 1
#162830000000
0#
0(
#162840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#162890000000
0$
0)
#162900000000
1"
1'
b0 +
b0 1
#162950000000
0"
0'
#162960000000
1#
1(
b101111101100100 +
b101111101100100 1
#163010000000
0#
0(
#163020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#163070000000
0$
0)
#163080000000
1"
1'
b0 +
b0 1
#163130000000
0"
0'
#163140000000
1#
1(
b101111101100100 +
b101111101100100 1
#163190000000
0#
0(
#163200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#163250000000
0$
0)
#163260000000
1"
1'
b0 +
b0 1
#163310000000
0"
0'
#163320000000
1#
1(
b101111101100100 +
b101111101100100 1
#163370000000
0#
0(
#163380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#163430000000
0$
0)
#163440000000
1"
1'
b0 +
b0 1
#163490000000
0"
0'
#163500000000
1#
1(
b101111101100100 +
b101111101100100 1
#163550000000
0#
0(
#163560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#163610000000
0$
0)
#163620000000
1"
1'
b0 +
b0 1
#163670000000
0"
0'
#163680000000
1#
1(
b101111101100100 +
b101111101100100 1
#163730000000
0#
0(
#163740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#163790000000
0$
0)
#163800000000
1"
1'
b0 +
b0 1
#163850000000
0"
0'
#163860000000
1#
1(
b101111101100100 +
b101111101100100 1
#163910000000
0#
0(
#163920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#163970000000
0$
0)
#163980000000
1"
1'
b0 +
b0 1
#164030000000
0"
0'
#164040000000
1#
1(
b101111101100100 +
b101111101100100 1
#164090000000
0#
0(
#164100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#164150000000
0$
0)
#164160000000
1"
1'
b0 +
b0 1
#164210000000
0"
0'
#164220000000
1#
1(
b101111101100100 +
b101111101100100 1
#164270000000
0#
0(
#164280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#164330000000
0$
0)
#164340000000
1"
1'
b0 +
b0 1
#164390000000
0"
0'
#164400000000
1#
1(
b101111101100100 +
b101111101100100 1
#164450000000
0#
0(
#164460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#164510000000
0$
0)
#164520000000
1"
1'
b0 +
b0 1
#164570000000
0"
0'
#164580000000
1#
1(
b101111101100100 +
b101111101100100 1
#164630000000
0#
0(
#164640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#164690000000
0$
0)
#164700000000
1"
1'
b0 +
b0 1
#164750000000
0"
0'
#164760000000
1#
1(
b101111101100100 +
b101111101100100 1
#164810000000
0#
0(
#164820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#164870000000
0$
0)
#164880000000
1"
1'
b0 +
b0 1
#164930000000
0"
0'
#164940000000
1#
1(
b101111101100100 +
b101111101100100 1
#164990000000
0#
0(
#165000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#165050000000
0$
0)
#165060000000
1"
1'
b0 +
b0 1
#165110000000
0"
0'
#165120000000
1#
1(
b101111101100100 +
b101111101100100 1
#165170000000
0#
0(
#165180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#165230000000
0$
0)
#165240000000
1"
1'
b0 +
b0 1
#165290000000
0"
0'
#165300000000
1#
1(
b101111101100100 +
b101111101100100 1
#165350000000
0#
0(
#165360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#165410000000
0$
0)
#165420000000
1"
1'
b0 +
b0 1
#165470000000
0"
0'
#165480000000
1#
1(
b101111101100100 +
b101111101100100 1
#165530000000
0#
0(
#165540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#165590000000
0$
0)
#165600000000
1"
1'
b0 +
b0 1
#165650000000
0"
0'
#165660000000
1#
1(
b101111101100100 +
b101111101100100 1
#165710000000
0#
0(
#165720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#165770000000
0$
0)
#165780000000
1"
1'
b0 +
b0 1
#165830000000
0"
0'
#165840000000
1#
1(
b101111101100100 +
b101111101100100 1
#165890000000
0#
0(
#165900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#165950000000
0$
0)
#165960000000
1"
1'
b0 +
b0 1
#166010000000
0"
0'
#166020000000
1#
1(
b101111101100100 +
b101111101100100 1
#166070000000
0#
0(
#166080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#166130000000
0$
0)
#166140000000
1"
1'
b0 +
b0 1
#166190000000
0"
0'
#166200000000
1#
1(
b101111101100100 +
b101111101100100 1
#166250000000
0#
0(
#166260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#166310000000
0$
0)
#166320000000
1"
1'
b0 +
b0 1
#166370000000
0"
0'
#166380000000
1#
1(
b101111101100100 +
b101111101100100 1
#166430000000
0#
0(
#166440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#166490000000
0$
0)
#166500000000
1"
1'
b0 +
b0 1
#166550000000
0"
0'
#166560000000
1#
1(
b101111101100100 +
b101111101100100 1
#166610000000
0#
0(
#166620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#166670000000
0$
0)
#166680000000
1"
1'
b0 +
b0 1
#166730000000
0"
0'
#166740000000
1#
1(
b101111101100100 +
b101111101100100 1
#166790000000
0#
0(
#166800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#166850000000
0$
0)
#166860000000
1"
1'
b0 +
b0 1
#166910000000
0"
0'
#166920000000
1#
1(
b101111101100100 +
b101111101100100 1
#166970000000
0#
0(
#166980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#167030000000
0$
0)
#167040000000
1"
1'
b0 +
b0 1
#167090000000
0"
0'
#167100000000
1#
1(
b101111101100100 +
b101111101100100 1
#167150000000
0#
0(
#167160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#167210000000
0$
0)
#167220000000
1"
1'
b0 +
b0 1
#167270000000
0"
0'
#167280000000
1#
1(
b101111101100100 +
b101111101100100 1
#167330000000
0#
0(
#167340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#167390000000
0$
0)
#167400000000
1"
1'
b0 +
b0 1
#167450000000
0"
0'
#167460000000
1#
1(
b101111101100100 +
b101111101100100 1
#167510000000
0#
0(
#167520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#167570000000
0$
0)
#167580000000
1"
1'
b0 +
b0 1
#167630000000
0"
0'
#167640000000
1#
1(
b101111101100100 +
b101111101100100 1
#167690000000
0#
0(
#167700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#167750000000
0$
0)
#167760000000
1"
1'
b0 +
b0 1
#167810000000
0"
0'
#167820000000
1#
1(
b101111101100100 +
b101111101100100 1
#167870000000
0#
0(
#167880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#167930000000
0$
0)
#167940000000
1"
1'
b0 +
b0 1
#167990000000
0"
0'
#168000000000
1#
1(
b101111101100100 +
b101111101100100 1
#168050000000
0#
0(
#168060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#168110000000
0$
0)
#168120000000
1"
1'
b0 +
b0 1
#168170000000
0"
0'
#168180000000
1#
1(
b101111101100100 +
b101111101100100 1
#168230000000
0#
0(
#168240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#168290000000
0$
0)
#168300000000
1"
1'
b0 +
b0 1
#168350000000
0"
0'
#168360000000
1#
1(
b101111101100100 +
b101111101100100 1
#168410000000
0#
0(
#168420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#168470000000
0$
0)
#168480000000
1"
1'
b0 +
b0 1
#168530000000
0"
0'
#168540000000
1#
1(
b101111101100100 +
b101111101100100 1
#168590000000
0#
0(
#168600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#168650000000
0$
0)
#168660000000
1"
1'
b0 +
b0 1
#168710000000
0"
0'
#168720000000
1#
1(
b101111101100100 +
b101111101100100 1
#168770000000
0#
0(
#168780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#168830000000
0$
0)
#168840000000
1"
1'
b0 +
b0 1
#168890000000
0"
0'
#168900000000
1#
1(
b101111101100100 +
b101111101100100 1
#168950000000
0#
0(
#168960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#169010000000
0$
0)
#169020000000
1"
1'
b0 +
b0 1
#169070000000
0"
0'
#169080000000
1#
1(
b101111101100100 +
b101111101100100 1
#169130000000
0#
0(
#169140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#169190000000
0$
0)
#169200000000
1"
1'
b0 +
b0 1
#169250000000
0"
0'
#169260000000
1#
1(
b101111101100100 +
b101111101100100 1
#169310000000
0#
0(
#169320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#169370000000
0$
0)
#169380000000
1"
1'
b0 +
b0 1
#169430000000
0"
0'
#169440000000
1#
1(
b101111101100100 +
b101111101100100 1
#169490000000
0#
0(
#169500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#169550000000
0$
0)
#169560000000
1"
1'
b0 +
b0 1
#169610000000
0"
0'
#169620000000
1#
1(
b101111101100100 +
b101111101100100 1
#169670000000
0#
0(
#169680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#169730000000
0$
0)
#169740000000
1"
1'
b0 +
b0 1
#169790000000
0"
0'
#169800000000
1#
1(
b101111101100100 +
b101111101100100 1
#169850000000
0#
0(
#169860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#169910000000
0$
0)
#169920000000
1"
1'
b0 +
b0 1
#169970000000
0"
0'
#169980000000
1#
1(
b101111101100100 +
b101111101100100 1
#170030000000
0#
0(
#170040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#170090000000
0$
0)
#170100000000
1"
1'
b0 +
b0 1
#170150000000
0"
0'
#170160000000
1#
1(
b101111101100100 +
b101111101100100 1
#170210000000
0#
0(
#170220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#170270000000
0$
0)
#170280000000
1"
1'
b0 +
b0 1
#170330000000
0"
0'
#170340000000
1#
1(
b101111101100100 +
b101111101100100 1
#170390000000
0#
0(
#170400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#170450000000
0$
0)
#170460000000
1"
1'
b0 +
b0 1
#170510000000
0"
0'
#170520000000
1#
1(
b101111101100100 +
b101111101100100 1
#170570000000
0#
0(
#170580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#170630000000
0$
0)
#170640000000
1"
1'
b0 +
b0 1
#170690000000
0"
0'
#170700000000
1#
1(
b101111101100100 +
b101111101100100 1
#170750000000
0#
0(
#170760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#170810000000
0$
0)
#170820000000
1"
1'
b0 +
b0 1
#170870000000
0"
0'
#170880000000
1#
1(
b101111101100100 +
b101111101100100 1
#170930000000
0#
0(
#170940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#170990000000
0$
0)
#171000000000
1"
1'
b0 +
b0 1
#171050000000
0"
0'
#171060000000
1#
1(
b101111101100100 +
b101111101100100 1
#171110000000
0#
0(
#171120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#171170000000
0$
0)
#171180000000
1"
1'
b0 +
b0 1
#171230000000
0"
0'
#171240000000
1#
1(
b101111101100100 +
b101111101100100 1
#171290000000
0#
0(
#171300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#171350000000
0$
0)
#171360000000
1"
1'
b0 +
b0 1
#171410000000
0"
0'
#171420000000
1#
1(
b101111101100100 +
b101111101100100 1
#171470000000
0#
0(
#171480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#171530000000
0$
0)
#171540000000
1"
1'
b0 +
b0 1
#171590000000
0"
0'
#171600000000
1#
1(
b101111101100100 +
b101111101100100 1
#171650000000
0#
0(
#171660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#171710000000
0$
0)
#171720000000
1"
1'
b0 +
b0 1
#171770000000
0"
0'
#171780000000
1#
1(
b101111101100100 +
b101111101100100 1
#171830000000
0#
0(
#171840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#171890000000
0$
0)
#171900000000
1"
1'
b0 +
b0 1
#171950000000
0"
0'
#171960000000
1#
1(
b101111101100100 +
b101111101100100 1
#172010000000
0#
0(
#172020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#172070000000
0$
0)
#172080000000
1"
1'
b0 +
b0 1
#172130000000
0"
0'
#172140000000
1#
1(
b101111101100100 +
b101111101100100 1
#172190000000
0#
0(
#172200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#172250000000
0$
0)
#172260000000
1"
1'
b0 +
b0 1
#172310000000
0"
0'
#172320000000
1#
1(
b101111101100100 +
b101111101100100 1
#172370000000
0#
0(
#172380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#172430000000
0$
0)
#172440000000
1"
1'
b0 +
b0 1
#172490000000
0"
0'
#172500000000
1#
1(
b101111101100100 +
b101111101100100 1
#172550000000
0#
0(
#172560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#172610000000
0$
0)
#172620000000
1"
1'
b0 +
b0 1
#172670000000
0"
0'
#172680000000
1#
1(
b101111101100100 +
b101111101100100 1
#172730000000
0#
0(
#172740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#172790000000
0$
0)
#172800000000
1"
1'
b0 +
b0 1
#172850000000
0"
0'
#172860000000
1#
1(
b101111101100100 +
b101111101100100 1
#172910000000
0#
0(
#172920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#172970000000
0$
0)
#172980000000
1"
1'
b0 +
b0 1
#173030000000
0"
0'
#173040000000
1#
1(
b101111101100100 +
b101111101100100 1
#173090000000
0#
0(
#173100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#173150000000
0$
0)
#173160000000
1"
1'
b0 +
b0 1
#173210000000
0"
0'
#173220000000
1#
1(
b101111101100100 +
b101111101100100 1
#173270000000
0#
0(
#173280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#173330000000
0$
0)
#173340000000
1"
1'
b0 +
b0 1
#173390000000
0"
0'
#173400000000
1#
1(
b101111101100100 +
b101111101100100 1
#173450000000
0#
0(
#173460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#173510000000
0$
0)
#173520000000
1"
1'
b0 +
b0 1
#173570000000
0"
0'
#173580000000
1#
1(
b101111101100100 +
b101111101100100 1
#173630000000
0#
0(
#173640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#173690000000
0$
0)
#173700000000
1"
1'
b0 +
b0 1
#173750000000
0"
0'
#173760000000
1#
1(
b101111101100100 +
b101111101100100 1
#173810000000
0#
0(
#173820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#173870000000
0$
0)
#173880000000
1"
1'
b0 +
b0 1
#173930000000
0"
0'
#173940000000
1#
1(
b101111101100100 +
b101111101100100 1
#173990000000
0#
0(
#174000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#174050000000
0$
0)
#174060000000
1"
1'
b0 +
b0 1
#174110000000
0"
0'
#174120000000
1#
1(
b101111101100100 +
b101111101100100 1
#174170000000
0#
0(
#174180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#174230000000
0$
0)
#174240000000
1"
1'
b0 +
b0 1
#174290000000
0"
0'
#174300000000
1#
1(
b101111101100100 +
b101111101100100 1
#174350000000
0#
0(
#174360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#174410000000
0$
0)
#174420000000
1"
1'
b0 +
b0 1
#174470000000
0"
0'
#174480000000
1#
1(
b101111101100100 +
b101111101100100 1
#174530000000
0#
0(
#174540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#174590000000
0$
0)
#174600000000
1"
1'
b0 +
b0 1
#174650000000
0"
0'
#174660000000
1#
1(
b101111101100100 +
b101111101100100 1
#174710000000
0#
0(
#174720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#174770000000
0$
0)
#174780000000
1"
1'
b0 +
b0 1
#174830000000
0"
0'
#174840000000
1#
1(
b101111101100100 +
b101111101100100 1
#174890000000
0#
0(
#174900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#174950000000
0$
0)
#174960000000
1"
1'
b0 +
b0 1
#175010000000
0"
0'
#175020000000
1#
1(
b101111101100100 +
b101111101100100 1
#175070000000
0#
0(
#175080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#175130000000
0$
0)
#175140000000
1"
1'
b0 +
b0 1
#175190000000
0"
0'
#175200000000
1#
1(
b101111101100100 +
b101111101100100 1
#175250000000
0#
0(
#175260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#175310000000
0$
0)
#175320000000
1"
1'
b0 +
b0 1
#175370000000
0"
0'
#175380000000
1#
1(
b101111101100100 +
b101111101100100 1
#175430000000
0#
0(
#175440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#175490000000
0$
0)
#175500000000
1"
1'
b0 +
b0 1
#175550000000
0"
0'
#175560000000
1#
1(
b101111101100100 +
b101111101100100 1
#175610000000
0#
0(
#175620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#175670000000
0$
0)
#175680000000
1"
1'
b0 +
b0 1
#175730000000
0"
0'
#175740000000
1#
1(
b101111101100100 +
b101111101100100 1
#175790000000
0#
0(
#175800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#175850000000
0$
0)
#175860000000
1"
1'
b0 +
b0 1
#175910000000
0"
0'
#175920000000
1#
1(
b101111101100100 +
b101111101100100 1
#175970000000
0#
0(
#175980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#176030000000
0$
0)
#176040000000
1"
1'
b0 +
b0 1
#176090000000
0"
0'
#176100000000
1#
1(
b101111101100100 +
b101111101100100 1
#176150000000
0#
0(
#176160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#176210000000
0$
0)
#176220000000
1"
1'
b0 +
b0 1
#176270000000
0"
0'
#176280000000
1#
1(
b101111101100100 +
b101111101100100 1
#176330000000
0#
0(
#176340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#176390000000
0$
0)
#176400000000
1"
1'
b0 +
b0 1
#176450000000
0"
0'
#176460000000
1#
1(
b101111101100100 +
b101111101100100 1
#176510000000
0#
0(
#176520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#176570000000
0$
0)
#176580000000
1"
1'
b0 +
b0 1
#176630000000
0"
0'
#176640000000
1#
1(
b101111101100100 +
b101111101100100 1
#176690000000
0#
0(
#176700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#176750000000
0$
0)
#176760000000
1"
1'
b0 +
b0 1
#176810000000
0"
0'
#176820000000
1#
1(
b101111101100100 +
b101111101100100 1
#176870000000
0#
0(
#176880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#176930000000
0$
0)
#176940000000
1"
1'
b0 +
b0 1
#176990000000
0"
0'
#177000000000
1#
1(
b101111101100100 +
b101111101100100 1
#177050000000
0#
0(
#177060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#177110000000
0$
0)
#177120000000
1"
1'
b0 +
b0 1
#177170000000
0"
0'
#177180000000
1#
1(
b101111101100100 +
b101111101100100 1
#177230000000
0#
0(
#177240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#177290000000
0$
0)
#177300000000
1"
1'
b0 +
b0 1
#177350000000
0"
0'
#177360000000
1#
1(
b101111101100100 +
b101111101100100 1
#177410000000
0#
0(
#177420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#177470000000
0$
0)
#177480000000
1"
1'
b0 +
b0 1
#177530000000
0"
0'
#177540000000
1#
1(
b101111101100100 +
b101111101100100 1
#177590000000
0#
0(
#177600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#177650000000
0$
0)
#177660000000
1"
1'
b0 +
b0 1
#177710000000
0"
0'
#177720000000
1#
1(
b101111101100100 +
b101111101100100 1
#177770000000
0#
0(
#177780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#177830000000
0$
0)
#177840000000
1"
1'
b0 +
b0 1
#177890000000
0"
0'
#177900000000
1#
1(
b101111101100100 +
b101111101100100 1
#177950000000
0#
0(
#177960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#178010000000
0$
0)
#178020000000
1"
1'
b0 +
b0 1
#178070000000
0"
0'
#178080000000
1#
1(
b101111101100100 +
b101111101100100 1
#178130000000
0#
0(
#178140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#178190000000
0$
0)
#178200000000
1"
1'
b0 +
b0 1
#178250000000
0"
0'
#178260000000
1#
1(
b101111101100100 +
b101111101100100 1
#178310000000
0#
0(
#178320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#178370000000
0$
0)
#178380000000
1"
1'
b0 +
b0 1
#178430000000
0"
0'
#178440000000
1#
1(
b101111101100100 +
b101111101100100 1
#178490000000
0#
0(
#178500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#178550000000
0$
0)
#178560000000
1"
1'
b0 +
b0 1
#178610000000
0"
0'
#178620000000
1#
1(
b101111101100100 +
b101111101100100 1
#178670000000
0#
0(
#178680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#178730000000
0$
0)
#178740000000
1"
1'
b0 +
b0 1
#178790000000
0"
0'
#178800000000
1#
1(
b101111101100100 +
b101111101100100 1
#178850000000
0#
0(
#178860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#178910000000
0$
0)
#178920000000
1"
1'
b0 +
b0 1
#178970000000
0"
0'
#178980000000
1#
1(
b101111101100100 +
b101111101100100 1
#179030000000
0#
0(
#179040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#179090000000
0$
0)
#179100000000
1"
1'
b0 +
b0 1
#179150000000
0"
0'
#179160000000
1#
1(
b101111101100100 +
b101111101100100 1
#179210000000
0#
0(
#179220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#179270000000
0$
0)
#179280000000
1"
1'
b0 +
b0 1
#179330000000
0"
0'
#179340000000
1#
1(
b101111101100100 +
b101111101100100 1
#179390000000
0#
0(
#179400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#179450000000
0$
0)
#179460000000
1"
1'
b0 +
b0 1
#179510000000
0"
0'
#179520000000
1#
1(
b101111101100100 +
b101111101100100 1
#179570000000
0#
0(
#179580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#179630000000
0$
0)
#179640000000
1"
1'
b0 +
b0 1
#179690000000
0"
0'
#179700000000
1#
1(
b101111101100100 +
b101111101100100 1
#179750000000
0#
0(
#179760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#179810000000
0$
0)
#179820000000
1"
1'
b0 +
b0 1
#179870000000
0"
0'
#179880000000
1#
1(
b101111101100100 +
b101111101100100 1
#179930000000
0#
0(
#179940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#179990000000
0$
0)
#180000000000
1"
1'
b0 +
b0 1
#180050000000
0"
0'
#180060000000
1#
1(
b101111101100100 +
b101111101100100 1
#180110000000
0#
0(
#180120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#180170000000
0$
0)
#180180000000
1"
1'
b0 +
b0 1
#180230000000
0"
0'
#180240000000
1#
1(
b101111101100100 +
b101111101100100 1
#180290000000
0#
0(
#180300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#180350000000
0$
0)
#180360000000
1"
1'
b0 +
b0 1
#180410000000
0"
0'
#180420000000
1#
1(
b101111101100100 +
b101111101100100 1
#180470000000
0#
0(
#180480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#180530000000
0$
0)
#180540000000
1"
1'
b0 +
b0 1
#180590000000
0"
0'
#180600000000
1#
1(
b101111101100100 +
b101111101100100 1
#180650000000
0#
0(
#180660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#180710000000
0$
0)
#180720000000
1"
1'
b0 +
b0 1
#180770000000
0"
0'
#180780000000
1#
1(
b101111101100100 +
b101111101100100 1
#180830000000
0#
0(
#180840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#180890000000
0$
0)
#180900000000
1"
1'
b0 +
b0 1
#180950000000
0"
0'
#180960000000
1#
1(
b101111101100100 +
b101111101100100 1
#181010000000
0#
0(
#181020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#181070000000
0$
0)
#181080000000
1"
1'
b0 +
b0 1
#181130000000
0"
0'
#181140000000
1#
1(
b101111101100100 +
b101111101100100 1
#181190000000
0#
0(
#181200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#181250000000
0$
0)
#181260000000
1"
1'
b0 +
b0 1
#181310000000
0"
0'
#181320000000
1#
1(
b101111101100100 +
b101111101100100 1
#181370000000
0#
0(
#181380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#181430000000
0$
0)
#181440000000
1"
1'
b0 +
b0 1
#181490000000
0"
0'
#181500000000
1#
1(
b101111101100100 +
b101111101100100 1
#181550000000
0#
0(
#181560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#181610000000
0$
0)
#181620000000
1"
1'
b0 +
b0 1
#181670000000
0"
0'
#181680000000
1#
1(
b101111101100100 +
b101111101100100 1
#181730000000
0#
0(
#181740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#181790000000
0$
0)
#181800000000
1"
1'
b0 +
b0 1
#181850000000
0"
0'
#181860000000
1#
1(
b101111101100100 +
b101111101100100 1
#181910000000
0#
0(
#181920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#181970000000
0$
0)
#181980000000
1"
1'
b0 +
b0 1
#182030000000
0"
0'
#182040000000
1#
1(
b101111101100100 +
b101111101100100 1
#182090000000
0#
0(
#182100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#182150000000
0$
0)
#182160000000
1"
1'
b0 +
b0 1
#182210000000
0"
0'
#182220000000
1#
1(
b101111101100100 +
b101111101100100 1
#182270000000
0#
0(
#182280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#182330000000
0$
0)
#182340000000
1"
1'
b0 +
b0 1
#182390000000
0"
0'
#182400000000
1#
1(
b101111101100100 +
b101111101100100 1
#182450000000
0#
0(
#182460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#182510000000
0$
0)
#182520000000
1"
1'
b0 +
b0 1
#182570000000
0"
0'
#182580000000
1#
1(
b101111101100100 +
b101111101100100 1
#182630000000
0#
0(
#182640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#182690000000
0$
0)
#182700000000
1"
1'
b0 +
b0 1
#182750000000
0"
0'
#182760000000
1#
1(
b101111101100100 +
b101111101100100 1
#182810000000
0#
0(
#182820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#182870000000
0$
0)
#182880000000
1"
1'
b0 +
b0 1
#182930000000
0"
0'
#182940000000
1#
1(
b101111101100100 +
b101111101100100 1
#182990000000
0#
0(
#183000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#183050000000
0$
0)
#183060000000
1"
1'
b0 +
b0 1
#183110000000
0"
0'
#183120000000
1#
1(
b101111101100100 +
b101111101100100 1
#183170000000
0#
0(
#183180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#183230000000
0$
0)
#183240000000
1"
1'
b0 +
b0 1
#183290000000
0"
0'
#183300000000
1#
1(
b101111101100100 +
b101111101100100 1
#183350000000
0#
0(
#183360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#183410000000
0$
0)
#183420000000
1"
1'
b0 +
b0 1
#183470000000
0"
0'
#183480000000
1#
1(
b101111101100100 +
b101111101100100 1
#183530000000
0#
0(
#183540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#183590000000
0$
0)
#183600000000
1"
1'
b0 +
b0 1
#183650000000
0"
0'
#183660000000
1#
1(
b101111101100100 +
b101111101100100 1
#183710000000
0#
0(
#183720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#183770000000
0$
0)
#183780000000
1"
1'
b0 +
b0 1
#183830000000
0"
0'
#183840000000
1#
1(
b101111101100100 +
b101111101100100 1
#183890000000
0#
0(
#183900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#183950000000
0$
0)
#183960000000
1"
1'
b0 +
b0 1
#184010000000
0"
0'
#184020000000
1#
1(
b101111101100100 +
b101111101100100 1
#184070000000
0#
0(
#184080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#184130000000
0$
0)
#184140000000
1"
1'
b0 +
b0 1
#184190000000
0"
0'
#184200000000
1#
1(
b101111101100100 +
b101111101100100 1
#184250000000
0#
0(
#184260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#184310000000
0$
0)
#184320000000
1"
1'
b0 +
b0 1
#184370000000
0"
0'
#184380000000
1#
1(
b101111101100100 +
b101111101100100 1
#184430000000
0#
0(
#184440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#184490000000
0$
0)
#184500000000
1"
1'
b0 +
b0 1
#184550000000
0"
0'
#184560000000
1#
1(
b101111101100100 +
b101111101100100 1
#184610000000
0#
0(
#184620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#184670000000
0$
0)
#184680000000
1"
1'
b0 +
b0 1
#184730000000
0"
0'
#184740000000
1#
1(
b101111101100100 +
b101111101100100 1
#184790000000
0#
0(
#184800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#184850000000
0$
0)
#184860000000
1"
1'
b0 +
b0 1
#184910000000
0"
0'
#184920000000
1#
1(
b101111101100100 +
b101111101100100 1
#184970000000
0#
0(
#184980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#185030000000
0$
0)
#185040000000
1"
1'
b0 +
b0 1
#185090000000
0"
0'
#185100000000
1#
1(
b101111101100100 +
b101111101100100 1
#185150000000
0#
0(
#185160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#185210000000
0$
0)
#185220000000
1"
1'
b0 +
b0 1
#185270000000
0"
0'
#185280000000
1#
1(
b101111101100100 +
b101111101100100 1
#185330000000
0#
0(
#185340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#185390000000
0$
0)
#185400000000
1"
1'
b0 +
b0 1
#185450000000
0"
0'
#185460000000
1#
1(
b101111101100100 +
b101111101100100 1
#185510000000
0#
0(
#185520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#185570000000
0$
0)
#185580000000
1"
1'
b0 +
b0 1
#185630000000
0"
0'
#185640000000
1#
1(
b101111101100100 +
b101111101100100 1
#185690000000
0#
0(
#185700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#185750000000
0$
0)
#185760000000
1"
1'
b0 +
b0 1
#185810000000
0"
0'
#185820000000
1#
1(
b101111101100100 +
b101111101100100 1
#185870000000
0#
0(
#185880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#185930000000
0$
0)
#185940000000
1"
1'
b0 +
b0 1
#185990000000
0"
0'
#186000000000
1#
1(
b101111101100100 +
b101111101100100 1
#186050000000
0#
0(
#186060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#186110000000
0$
0)
#186120000000
1"
1'
b0 +
b0 1
#186170000000
0"
0'
#186180000000
1#
1(
b101111101100100 +
b101111101100100 1
#186230000000
0#
0(
#186240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#186290000000
0$
0)
#186300000000
1"
1'
b0 +
b0 1
#186350000000
0"
0'
#186360000000
1#
1(
b101111101100100 +
b101111101100100 1
#186410000000
0#
0(
#186420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#186470000000
0$
0)
#186480000000
1"
1'
b0 +
b0 1
#186530000000
0"
0'
#186540000000
1#
1(
b101111101100100 +
b101111101100100 1
#186590000000
0#
0(
#186600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#186650000000
0$
0)
#186660000000
1"
1'
b0 +
b0 1
#186710000000
0"
0'
#186720000000
1#
1(
b101111101100100 +
b101111101100100 1
#186770000000
0#
0(
#186780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#186830000000
0$
0)
#186840000000
1"
1'
b0 +
b0 1
#186890000000
0"
0'
#186900000000
1#
1(
b101111101100100 +
b101111101100100 1
#186950000000
0#
0(
#186960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#187010000000
0$
0)
#187020000000
1"
1'
b0 +
b0 1
#187070000000
0"
0'
#187080000000
1#
1(
b101111101100100 +
b101111101100100 1
#187130000000
0#
0(
#187140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#187190000000
0$
0)
#187200000000
1"
1'
b0 +
b0 1
#187250000000
0"
0'
#187260000000
1#
1(
b101111101100100 +
b101111101100100 1
#187310000000
0#
0(
#187320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#187370000000
0$
0)
#187380000000
1"
1'
b0 +
b0 1
#187430000000
0"
0'
#187440000000
1#
1(
b101111101100100 +
b101111101100100 1
#187490000000
0#
0(
#187500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#187550000000
0$
0)
#187560000000
1"
1'
b0 +
b0 1
#187610000000
0"
0'
#187620000000
1#
1(
b101111101100100 +
b101111101100100 1
#187670000000
0#
0(
#187680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#187730000000
0$
0)
#187740000000
1"
1'
b0 +
b0 1
#187790000000
0"
0'
#187800000000
1#
1(
b101111101100100 +
b101111101100100 1
#187850000000
0#
0(
#187860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#187910000000
0$
0)
#187920000000
1"
1'
b0 +
b0 1
#187970000000
0"
0'
#187980000000
1#
1(
b101111101100100 +
b101111101100100 1
#188030000000
0#
0(
#188040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#188090000000
0$
0)
#188100000000
1"
1'
b0 +
b0 1
#188150000000
0"
0'
#188160000000
1#
1(
b101111101100100 +
b101111101100100 1
#188210000000
0#
0(
#188220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#188270000000
0$
0)
#188280000000
1"
1'
b0 +
b0 1
#188330000000
0"
0'
#188340000000
1#
1(
b101111101100100 +
b101111101100100 1
#188390000000
0#
0(
#188400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#188450000000
0$
0)
#188460000000
1"
1'
b0 +
b0 1
#188510000000
0"
0'
#188520000000
1#
1(
b101111101100100 +
b101111101100100 1
#188570000000
0#
0(
#188580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#188630000000
0$
0)
#188640000000
1"
1'
b0 +
b0 1
#188690000000
0"
0'
#188700000000
1#
1(
b101111101100100 +
b101111101100100 1
#188750000000
0#
0(
#188760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#188810000000
0$
0)
#188820000000
1"
1'
b0 +
b0 1
#188870000000
0"
0'
#188880000000
1#
1(
b101111101100100 +
b101111101100100 1
#188930000000
0#
0(
#188940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#188990000000
0$
0)
#189000000000
1"
1'
b0 +
b0 1
#189050000000
0"
0'
#189060000000
1#
1(
b101111101100100 +
b101111101100100 1
#189110000000
0#
0(
#189120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#189170000000
0$
0)
#189180000000
1"
1'
b0 +
b0 1
#189230000000
0"
0'
#189240000000
1#
1(
b101111101100100 +
b101111101100100 1
#189290000000
0#
0(
#189300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#189350000000
0$
0)
#189360000000
1"
1'
b0 +
b0 1
#189410000000
0"
0'
#189420000000
1#
1(
b101111101100100 +
b101111101100100 1
#189470000000
0#
0(
#189480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#189530000000
0$
0)
#189540000000
1"
1'
b0 +
b0 1
#189590000000
0"
0'
#189600000000
1#
1(
b101111101100100 +
b101111101100100 1
#189650000000
0#
0(
#189660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#189710000000
0$
0)
#189720000000
1"
1'
b0 +
b0 1
#189770000000
0"
0'
#189780000000
1#
1(
b101111101100100 +
b101111101100100 1
#189830000000
0#
0(
#189840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#189890000000
0$
0)
#189900000000
1"
1'
b0 +
b0 1
#189950000000
0"
0'
#189960000000
1#
1(
b101111101100100 +
b101111101100100 1
#190010000000
0#
0(
#190020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#190070000000
0$
0)
#190080000000
1"
1'
b0 +
b0 1
#190130000000
0"
0'
#190140000000
1#
1(
b101111101100100 +
b101111101100100 1
#190190000000
0#
0(
#190200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#190250000000
0$
0)
#190260000000
1"
1'
b0 +
b0 1
#190310000000
0"
0'
#190320000000
1#
1(
b101111101100100 +
b101111101100100 1
#190370000000
0#
0(
#190380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#190430000000
0$
0)
#190440000000
1"
1'
b0 +
b0 1
#190490000000
0"
0'
#190500000000
1#
1(
b101111101100100 +
b101111101100100 1
#190550000000
0#
0(
#190560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#190610000000
0$
0)
#190620000000
1"
1'
b0 +
b0 1
#190670000000
0"
0'
#190680000000
1#
1(
b101111101100100 +
b101111101100100 1
#190730000000
0#
0(
#190740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#190790000000
0$
0)
#190800000000
1"
1'
b0 +
b0 1
#190850000000
0"
0'
#190860000000
1#
1(
b101111101100100 +
b101111101100100 1
#190910000000
0#
0(
#190920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#190970000000
0$
0)
#190980000000
1"
1'
b0 +
b0 1
#191030000000
0"
0'
#191040000000
1#
1(
b101111101100100 +
b101111101100100 1
#191090000000
0#
0(
#191100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#191150000000
0$
0)
#191160000000
1"
1'
b0 +
b0 1
#191210000000
0"
0'
#191220000000
1#
1(
b101111101100100 +
b101111101100100 1
#191270000000
0#
0(
#191280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#191330000000
0$
0)
#191340000000
1"
1'
b0 +
b0 1
#191390000000
0"
0'
#191400000000
1#
1(
b101111101100100 +
b101111101100100 1
#191450000000
0#
0(
#191460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#191510000000
0$
0)
#191520000000
1"
1'
b0 +
b0 1
#191570000000
0"
0'
#191580000000
1#
1(
b101111101100100 +
b101111101100100 1
#191630000000
0#
0(
#191640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#191690000000
0$
0)
#191700000000
1"
1'
b0 +
b0 1
#191750000000
0"
0'
#191760000000
1#
1(
b101111101100100 +
b101111101100100 1
#191810000000
0#
0(
#191820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#191870000000
0$
0)
#191880000000
1"
1'
b0 +
b0 1
#191930000000
0"
0'
#191940000000
1#
1(
b101111101100100 +
b101111101100100 1
#191990000000
0#
0(
#192000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#192050000000
0$
0)
#192060000000
1"
1'
b0 +
b0 1
#192110000000
0"
0'
#192120000000
1#
1(
b101111101100100 +
b101111101100100 1
#192170000000
0#
0(
#192180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#192230000000
0$
0)
#192240000000
1"
1'
b0 +
b0 1
#192290000000
0"
0'
#192300000000
1#
1(
b101111101100100 +
b101111101100100 1
#192350000000
0#
0(
#192360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#192410000000
0$
0)
#192420000000
1"
1'
b0 +
b0 1
#192470000000
0"
0'
#192480000000
1#
1(
b101111101100100 +
b101111101100100 1
#192530000000
0#
0(
#192540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#192590000000
0$
0)
#192600000000
1"
1'
b0 +
b0 1
#192650000000
0"
0'
#192660000000
1#
1(
b101111101100100 +
b101111101100100 1
#192710000000
0#
0(
#192720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#192770000000
0$
0)
#192780000000
1"
1'
b0 +
b0 1
#192830000000
0"
0'
#192840000000
1#
1(
b101111101100100 +
b101111101100100 1
#192890000000
0#
0(
#192900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#192950000000
0$
0)
#192960000000
1"
1'
b0 +
b0 1
#193010000000
0"
0'
#193020000000
1#
1(
b101111101100100 +
b101111101100100 1
#193070000000
0#
0(
#193080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#193130000000
0$
0)
#193140000000
1"
1'
b0 +
b0 1
#193190000000
0"
0'
#193200000000
1#
1(
b101111101100100 +
b101111101100100 1
#193250000000
0#
0(
#193260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#193310000000
0$
0)
#193320000000
1"
1'
b0 +
b0 1
#193370000000
0"
0'
#193380000000
1#
1(
b101111101100100 +
b101111101100100 1
#193430000000
0#
0(
#193440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#193490000000
0$
0)
#193500000000
1"
1'
b0 +
b0 1
#193550000000
0"
0'
#193560000000
1#
1(
b101111101100100 +
b101111101100100 1
#193610000000
0#
0(
#193620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#193670000000
0$
0)
#193680000000
1"
1'
b0 +
b0 1
#193730000000
0"
0'
#193740000000
1#
1(
b101111101100100 +
b101111101100100 1
#193790000000
0#
0(
#193800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#193850000000
0$
0)
#193860000000
1"
1'
b0 +
b0 1
#193910000000
0"
0'
#193920000000
1#
1(
b101111101100100 +
b101111101100100 1
#193970000000
0#
0(
#193980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#194030000000
0$
0)
#194040000000
1"
1'
b0 +
b0 1
#194090000000
0"
0'
#194100000000
1#
1(
b101111101100100 +
b101111101100100 1
#194150000000
0#
0(
#194160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#194210000000
0$
0)
#194220000000
1"
1'
b0 +
b0 1
#194270000000
0"
0'
#194280000000
1#
1(
b101111101100100 +
b101111101100100 1
#194330000000
0#
0(
#194340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#194390000000
0$
0)
#194400000000
1"
1'
b0 +
b0 1
#194450000000
0"
0'
#194460000000
1#
1(
b101111101100100 +
b101111101100100 1
#194510000000
0#
0(
#194520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#194570000000
0$
0)
#194580000000
1"
1'
b0 +
b0 1
#194630000000
0"
0'
#194640000000
1#
1(
b101111101100100 +
b101111101100100 1
#194690000000
0#
0(
#194700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#194750000000
0$
0)
#194760000000
1"
1'
b0 +
b0 1
#194810000000
0"
0'
#194820000000
1#
1(
b101111101100100 +
b101111101100100 1
#194870000000
0#
0(
#194880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#194930000000
0$
0)
#194940000000
1"
1'
b0 +
b0 1
#194990000000
0"
0'
#195000000000
1#
1(
b101111101100100 +
b101111101100100 1
#195050000000
0#
0(
#195060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#195110000000
0$
0)
#195120000000
1"
1'
b0 +
b0 1
#195170000000
0"
0'
#195180000000
1#
1(
b101111101100100 +
b101111101100100 1
#195230000000
0#
0(
#195240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#195290000000
0$
0)
#195300000000
1"
1'
b0 +
b0 1
#195350000000
0"
0'
#195360000000
1#
1(
b101111101100100 +
b101111101100100 1
#195410000000
0#
0(
#195420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#195470000000
0$
0)
#195480000000
1"
1'
b0 +
b0 1
#195530000000
0"
0'
#195540000000
1#
1(
b101111101100100 +
b101111101100100 1
#195590000000
0#
0(
#195600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#195650000000
0$
0)
#195660000000
1"
1'
b0 +
b0 1
#195710000000
0"
0'
#195720000000
1#
1(
b101111101100100 +
b101111101100100 1
#195770000000
0#
0(
#195780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#195830000000
0$
0)
#195840000000
1"
1'
b0 +
b0 1
#195890000000
0"
0'
#195900000000
1#
1(
b101111101100100 +
b101111101100100 1
#195950000000
0#
0(
#195960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#196010000000
0$
0)
#196020000000
1"
1'
b0 +
b0 1
#196070000000
0"
0'
#196080000000
1#
1(
b101111101100100 +
b101111101100100 1
#196130000000
0#
0(
#196140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#196190000000
0$
0)
#196200000000
1"
1'
b0 +
b0 1
#196250000000
0"
0'
#196260000000
1#
1(
b101111101100100 +
b101111101100100 1
#196310000000
0#
0(
#196320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#196370000000
0$
0)
#196380000000
1"
1'
b0 +
b0 1
#196430000000
0"
0'
#196440000000
1#
1(
b101111101100100 +
b101111101100100 1
#196490000000
0#
0(
#196500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#196550000000
0$
0)
#196560000000
1"
1'
b0 +
b0 1
#196610000000
0"
0'
#196620000000
1#
1(
b101111101100100 +
b101111101100100 1
#196670000000
0#
0(
#196680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#196730000000
0$
0)
#196740000000
1"
1'
b0 +
b0 1
#196790000000
0"
0'
#196800000000
1#
1(
b101111101100100 +
b101111101100100 1
#196850000000
0#
0(
#196860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#196910000000
0$
0)
#196920000000
1"
1'
b0 +
b0 1
#196970000000
0"
0'
#196980000000
1#
1(
b101111101100100 +
b101111101100100 1
#197030000000
0#
0(
#197040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#197090000000
0$
0)
#197100000000
1"
1'
b0 +
b0 1
#197150000000
0"
0'
#197160000000
1#
1(
b101111101100100 +
b101111101100100 1
#197210000000
0#
0(
#197220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#197270000000
0$
0)
#197280000000
1"
1'
b0 +
b0 1
#197330000000
0"
0'
#197340000000
1#
1(
b101111101100100 +
b101111101100100 1
#197390000000
0#
0(
#197400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#197450000000
0$
0)
#197460000000
1"
1'
b0 +
b0 1
#197510000000
0"
0'
#197520000000
1#
1(
b101111101100100 +
b101111101100100 1
#197570000000
0#
0(
#197580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#197630000000
0$
0)
#197640000000
1"
1'
b0 +
b0 1
#197690000000
0"
0'
#197700000000
1#
1(
b101111101100100 +
b101111101100100 1
#197750000000
0#
0(
#197760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#197810000000
0$
0)
#197820000000
1"
1'
b0 +
b0 1
#197870000000
0"
0'
#197880000000
1#
1(
b101111101100100 +
b101111101100100 1
#197930000000
0#
0(
#197940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#197990000000
0$
0)
#198000000000
1"
1'
b0 +
b0 1
#198050000000
0"
0'
#198060000000
1#
1(
b101111101100100 +
b101111101100100 1
#198110000000
0#
0(
#198120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#198170000000
0$
0)
#198180000000
1"
1'
b0 +
b0 1
#198230000000
0"
0'
#198240000000
1#
1(
b101111101100100 +
b101111101100100 1
#198290000000
0#
0(
#198300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#198350000000
0$
0)
#198360000000
1"
1'
b0 +
b0 1
#198410000000
0"
0'
#198420000000
1#
1(
b101111101100100 +
b101111101100100 1
#198470000000
0#
0(
#198480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#198530000000
0$
0)
#198540000000
1"
1'
b0 +
b0 1
#198590000000
0"
0'
#198600000000
1#
1(
b101111101100100 +
b101111101100100 1
#198650000000
0#
0(
#198660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#198710000000
0$
0)
#198720000000
1"
1'
b0 +
b0 1
#198770000000
0"
0'
#198780000000
1#
1(
b101111101100100 +
b101111101100100 1
#198830000000
0#
0(
#198840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#198890000000
0$
0)
#198900000000
1"
1'
b0 +
b0 1
#198950000000
0"
0'
#198960000000
1#
1(
b101111101100100 +
b101111101100100 1
#199010000000
0#
0(
#199020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#199070000000
0$
0)
#199080000000
1"
1'
b0 +
b0 1
#199130000000
0"
0'
#199140000000
1#
1(
b101111101100100 +
b101111101100100 1
#199190000000
0#
0(
#199200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#199250000000
0$
0)
#199260000000
1"
1'
b0 +
b0 1
#199310000000
0"
0'
#199320000000
1#
1(
b101111101100100 +
b101111101100100 1
#199370000000
0#
0(
#199380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#199430000000
0$
0)
#199440000000
1"
1'
b0 +
b0 1
#199490000000
0"
0'
#199500000000
1#
1(
b101111101100100 +
b101111101100100 1
#199550000000
0#
0(
#199560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#199610000000
0$
0)
#199620000000
1"
1'
b0 +
b0 1
#199670000000
0"
0'
#199680000000
1#
1(
b101111101100100 +
b101111101100100 1
#199730000000
0#
0(
#199740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#199790000000
0$
0)
#199800000000
1"
1'
b0 +
b0 1
#199850000000
0"
0'
#199860000000
1#
1(
b101111101100100 +
b101111101100100 1
#199910000000
0#
0(
#199920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#199970000000
0$
0)
#199980000000
1"
1'
b0 +
b0 1
#200030000000
0"
0'
#200040000000
1#
1(
b101111101100100 +
b101111101100100 1
#200090000000
0#
0(
#200100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#200150000000
0$
0)
#200160000000
1"
1'
b0 +
b0 1
#200210000000
0"
0'
#200220000000
1#
1(
b101111101100100 +
b101111101100100 1
#200270000000
0#
0(
#200280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#200330000000
0$
0)
#200340000000
1"
1'
b0 +
b0 1
#200390000000
0"
0'
#200400000000
1#
1(
b101111101100100 +
b101111101100100 1
#200450000000
0#
0(
#200460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#200510000000
0$
0)
#200520000000
1"
1'
b0 +
b0 1
#200570000000
0"
0'
#200580000000
1#
1(
b101111101100100 +
b101111101100100 1
#200630000000
0#
0(
#200640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#200690000000
0$
0)
#200700000000
1"
1'
b0 +
b0 1
#200750000000
0"
0'
#200760000000
1#
1(
b101111101100100 +
b101111101100100 1
#200810000000
0#
0(
#200820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#200870000000
0$
0)
#200880000000
1"
1'
b0 +
b0 1
#200930000000
0"
0'
#200940000000
1#
1(
b101111101100100 +
b101111101100100 1
#200990000000
0#
0(
#201000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#201050000000
0$
0)
#201060000000
1"
1'
b0 +
b0 1
#201110000000
0"
0'
#201120000000
1#
1(
b101111101100100 +
b101111101100100 1
#201170000000
0#
0(
#201180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#201230000000
0$
0)
#201240000000
1"
1'
b0 +
b0 1
#201290000000
0"
0'
#201300000000
1#
1(
b101111101100100 +
b101111101100100 1
#201350000000
0#
0(
#201360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#201410000000
0$
0)
#201420000000
1"
1'
b0 +
b0 1
#201470000000
0"
0'
#201480000000
1#
1(
b101111101100100 +
b101111101100100 1
#201530000000
0#
0(
#201540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#201590000000
0$
0)
#201600000000
1"
1'
b0 +
b0 1
#201650000000
0"
0'
#201660000000
1#
1(
b101111101100100 +
b101111101100100 1
#201710000000
0#
0(
#201720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#201770000000
0$
0)
#201780000000
1"
1'
b0 +
b0 1
#201830000000
0"
0'
#201840000000
1#
1(
b101111101100100 +
b101111101100100 1
#201890000000
0#
0(
#201900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#201950000000
0$
0)
#201960000000
1"
1'
b0 +
b0 1
#202010000000
0"
0'
#202020000000
1#
1(
b101111101100100 +
b101111101100100 1
#202070000000
0#
0(
#202080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#202130000000
0$
0)
#202140000000
1"
1'
b0 +
b0 1
#202190000000
0"
0'
#202200000000
1#
1(
b101111101100100 +
b101111101100100 1
#202250000000
0#
0(
#202260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#202310000000
0$
0)
#202320000000
1"
1'
b0 +
b0 1
#202370000000
0"
0'
#202380000000
1#
1(
b101111101100100 +
b101111101100100 1
#202430000000
0#
0(
#202440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#202490000000
0$
0)
#202500000000
1"
1'
b0 +
b0 1
#202550000000
0"
0'
#202560000000
1#
1(
b101111101100100 +
b101111101100100 1
#202610000000
0#
0(
#202620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#202670000000
0$
0)
#202680000000
1"
1'
b0 +
b0 1
#202730000000
0"
0'
#202740000000
1#
1(
b101111101100100 +
b101111101100100 1
#202790000000
0#
0(
#202800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#202850000000
0$
0)
#202860000000
1"
1'
b0 +
b0 1
#202910000000
0"
0'
#202920000000
1#
1(
b101111101100100 +
b101111101100100 1
#202970000000
0#
0(
#202980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#203030000000
0$
0)
#203040000000
1"
1'
b0 +
b0 1
#203090000000
0"
0'
#203100000000
1#
1(
b101111101100100 +
b101111101100100 1
#203150000000
0#
0(
#203160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#203210000000
0$
0)
#203220000000
1"
1'
b0 +
b0 1
#203270000000
0"
0'
#203280000000
1#
1(
b101111101100100 +
b101111101100100 1
#203330000000
0#
0(
#203340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#203390000000
0$
0)
#203400000000
1"
1'
b0 +
b0 1
#203450000000
0"
0'
#203460000000
1#
1(
b101111101100100 +
b101111101100100 1
#203510000000
0#
0(
#203520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#203570000000
0$
0)
#203580000000
1"
1'
b0 +
b0 1
#203630000000
0"
0'
#203640000000
1#
1(
b101111101100100 +
b101111101100100 1
#203690000000
0#
0(
#203700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#203750000000
0$
0)
#203760000000
1"
1'
b0 +
b0 1
#203810000000
0"
0'
#203820000000
1#
1(
b101111101100100 +
b101111101100100 1
#203870000000
0#
0(
#203880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#203930000000
0$
0)
#203940000000
1"
1'
b0 +
b0 1
#203990000000
0"
0'
#204000000000
1#
1(
b101111101100100 +
b101111101100100 1
#204050000000
0#
0(
#204060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#204110000000
0$
0)
#204120000000
1"
1'
b0 +
b0 1
#204170000000
0"
0'
#204180000000
1#
1(
b101111101100100 +
b101111101100100 1
#204230000000
0#
0(
#204240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#204290000000
0$
0)
#204300000000
1"
1'
b0 +
b0 1
#204350000000
0"
0'
#204360000000
1#
1(
b101111101100100 +
b101111101100100 1
#204410000000
0#
0(
#204420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#204470000000
0$
0)
#204480000000
1"
1'
b0 +
b0 1
#204530000000
0"
0'
#204540000000
1#
1(
b101111101100100 +
b101111101100100 1
#204590000000
0#
0(
#204600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#204650000000
0$
0)
#204660000000
1"
1'
b0 +
b0 1
#204710000000
0"
0'
#204720000000
1#
1(
b101111101100100 +
b101111101100100 1
#204770000000
0#
0(
#204780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#204830000000
0$
0)
#204840000000
1"
1'
b0 +
b0 1
#204890000000
0"
0'
#204900000000
1#
1(
b101111101100100 +
b101111101100100 1
#204950000000
0#
0(
#204960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#205010000000
0$
0)
#205020000000
1"
1'
b0 +
b0 1
#205070000000
0"
0'
#205080000000
1#
1(
b101111101100100 +
b101111101100100 1
#205130000000
0#
0(
#205140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#205190000000
0$
0)
#205200000000
1"
1'
b0 +
b0 1
#205250000000
0"
0'
#205260000000
1#
1(
b101111101100100 +
b101111101100100 1
#205310000000
0#
0(
#205320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#205370000000
0$
0)
#205380000000
1"
1'
b0 +
b0 1
#205430000000
0"
0'
#205440000000
1#
1(
b101111101100100 +
b101111101100100 1
#205490000000
0#
0(
#205500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#205550000000
0$
0)
#205560000000
1"
1'
b0 +
b0 1
#205610000000
0"
0'
#205620000000
1#
1(
b101111101100100 +
b101111101100100 1
#205670000000
0#
0(
#205680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#205730000000
0$
0)
#205740000000
1"
1'
b0 +
b0 1
#205790000000
0"
0'
#205800000000
1#
1(
b101111101100100 +
b101111101100100 1
#205850000000
0#
0(
#205860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#205910000000
0$
0)
#205920000000
1"
1'
b0 +
b0 1
#205970000000
0"
0'
#205980000000
1#
1(
b101111101100100 +
b101111101100100 1
#206030000000
0#
0(
#206040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#206090000000
0$
0)
#206100000000
1"
1'
b0 +
b0 1
#206150000000
0"
0'
#206160000000
1#
1(
b101111101100100 +
b101111101100100 1
#206210000000
0#
0(
#206220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#206270000000
0$
0)
#206280000000
1"
1'
b0 +
b0 1
#206330000000
0"
0'
#206340000000
1#
1(
b101111101100100 +
b101111101100100 1
#206390000000
0#
0(
#206400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#206450000000
0$
0)
#206460000000
1"
1'
b0 +
b0 1
#206510000000
0"
0'
#206520000000
1#
1(
b101111101100100 +
b101111101100100 1
#206570000000
0#
0(
#206580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#206630000000
0$
0)
#206640000000
1"
1'
b0 +
b0 1
#206690000000
0"
0'
#206700000000
1#
1(
b101111101100100 +
b101111101100100 1
#206750000000
0#
0(
#206760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#206810000000
0$
0)
#206820000000
1"
1'
b0 +
b0 1
#206870000000
0"
0'
#206880000000
1#
1(
b101111101100100 +
b101111101100100 1
#206930000000
0#
0(
#206940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#206990000000
0$
0)
#207000000000
1"
1'
b0 +
b0 1
#207050000000
0"
0'
#207060000000
1#
1(
b101111101100100 +
b101111101100100 1
#207110000000
0#
0(
#207120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#207170000000
0$
0)
#207180000000
1"
1'
b0 +
b0 1
#207230000000
0"
0'
#207240000000
1#
1(
b101111101100100 +
b101111101100100 1
#207290000000
0#
0(
#207300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#207350000000
0$
0)
#207360000000
1"
1'
b0 +
b0 1
#207410000000
0"
0'
#207420000000
1#
1(
b101111101100100 +
b101111101100100 1
#207470000000
0#
0(
#207480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#207530000000
0$
0)
#207540000000
1"
1'
b0 +
b0 1
#207590000000
0"
0'
#207600000000
1#
1(
b101111101100100 +
b101111101100100 1
#207650000000
0#
0(
#207660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#207710000000
0$
0)
#207720000000
1"
1'
b0 +
b0 1
#207770000000
0"
0'
#207780000000
1#
1(
b101111101100100 +
b101111101100100 1
#207830000000
0#
0(
#207840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#207890000000
0$
0)
#207900000000
1"
1'
b0 +
b0 1
#207950000000
0"
0'
#207960000000
1#
1(
b101111101100100 +
b101111101100100 1
#208010000000
0#
0(
#208020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#208070000000
0$
0)
#208080000000
1"
1'
b0 +
b0 1
#208130000000
0"
0'
#208140000000
1#
1(
b101111101100100 +
b101111101100100 1
#208190000000
0#
0(
#208200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#208250000000
0$
0)
#208260000000
1"
1'
b0 +
b0 1
#208310000000
0"
0'
#208320000000
1#
1(
b101111101100100 +
b101111101100100 1
#208370000000
0#
0(
#208380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#208430000000
0$
0)
#208440000000
1"
1'
b0 +
b0 1
#208490000000
0"
0'
#208500000000
1#
1(
b101111101100100 +
b101111101100100 1
#208550000000
0#
0(
#208560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#208610000000
0$
0)
#208620000000
1"
1'
b0 +
b0 1
#208670000000
0"
0'
#208680000000
1#
1(
b101111101100100 +
b101111101100100 1
#208730000000
0#
0(
#208740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#208790000000
0$
0)
#208800000000
1"
1'
b0 +
b0 1
#208850000000
0"
0'
#208860000000
1#
1(
b101111101100100 +
b101111101100100 1
#208910000000
0#
0(
#208920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#208970000000
0$
0)
#208980000000
1"
1'
b0 +
b0 1
#209030000000
0"
0'
#209040000000
1#
1(
b101111101100100 +
b101111101100100 1
#209090000000
0#
0(
#209100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#209150000000
0$
0)
#209160000000
1"
1'
b0 +
b0 1
#209210000000
0"
0'
#209220000000
1#
1(
b101111101100100 +
b101111101100100 1
#209270000000
0#
0(
#209280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#209330000000
0$
0)
#209340000000
1"
1'
b0 +
b0 1
#209390000000
0"
0'
#209400000000
1#
1(
b101111101100100 +
b101111101100100 1
#209450000000
0#
0(
#209460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#209510000000
0$
0)
#209520000000
1"
1'
b0 +
b0 1
#209570000000
0"
0'
#209580000000
1#
1(
b101111101100100 +
b101111101100100 1
#209630000000
0#
0(
#209640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#209690000000
0$
0)
#209700000000
1"
1'
b0 +
b0 1
#209750000000
0"
0'
#209760000000
1#
1(
b101111101100100 +
b101111101100100 1
#209810000000
0#
0(
#209820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#209870000000
0$
0)
#209880000000
1"
1'
b0 +
b0 1
#209930000000
0"
0'
#209940000000
1#
1(
b101111101100100 +
b101111101100100 1
#209990000000
0#
0(
#210000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#210050000000
0$
0)
#210060000000
1"
1'
b0 +
b0 1
#210110000000
0"
0'
#210120000000
1#
1(
b101111101100100 +
b101111101100100 1
#210170000000
0#
0(
#210180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#210230000000
0$
0)
#210240000000
1"
1'
b0 +
b0 1
#210290000000
0"
0'
#210300000000
1#
1(
b101111101100100 +
b101111101100100 1
#210350000000
0#
0(
#210360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#210410000000
0$
0)
#210420000000
1"
1'
b0 +
b0 1
#210470000000
0"
0'
#210480000000
1#
1(
b101111101100100 +
b101111101100100 1
#210530000000
0#
0(
#210540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#210590000000
0$
0)
#210600000000
1"
1'
b0 +
b0 1
#210650000000
0"
0'
#210660000000
1#
1(
b101111101100100 +
b101111101100100 1
#210710000000
0#
0(
#210720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#210770000000
0$
0)
#210780000000
1"
1'
b0 +
b0 1
#210830000000
0"
0'
#210840000000
1#
1(
b101111101100100 +
b101111101100100 1
#210890000000
0#
0(
#210900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#210950000000
0$
0)
#210960000000
1"
1'
b0 +
b0 1
#211010000000
0"
0'
#211020000000
1#
1(
b101111101100100 +
b101111101100100 1
#211070000000
0#
0(
#211080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#211130000000
0$
0)
#211140000000
1"
1'
b0 +
b0 1
#211190000000
0"
0'
#211200000000
1#
1(
b101111101100100 +
b101111101100100 1
#211250000000
0#
0(
#211260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#211310000000
0$
0)
#211320000000
1"
1'
b0 +
b0 1
#211370000000
0"
0'
#211380000000
1#
1(
b101111101100100 +
b101111101100100 1
#211430000000
0#
0(
#211440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#211490000000
0$
0)
#211500000000
1"
1'
b0 +
b0 1
#211550000000
0"
0'
#211560000000
1#
1(
b101111101100100 +
b101111101100100 1
#211610000000
0#
0(
#211620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#211670000000
0$
0)
#211680000000
1"
1'
b0 +
b0 1
#211730000000
0"
0'
#211740000000
1#
1(
b101111101100100 +
b101111101100100 1
#211790000000
0#
0(
#211800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#211850000000
0$
0)
#211860000000
1"
1'
b0 +
b0 1
#211910000000
0"
0'
#211920000000
1#
1(
b101111101100100 +
b101111101100100 1
#211970000000
0#
0(
#211980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#212030000000
0$
0)
#212040000000
1"
1'
b0 +
b0 1
#212090000000
0"
0'
#212100000000
1#
1(
b101111101100100 +
b101111101100100 1
#212150000000
0#
0(
#212160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#212210000000
0$
0)
#212220000000
1"
1'
b0 +
b0 1
#212270000000
0"
0'
#212280000000
1#
1(
b101111101100100 +
b101111101100100 1
#212330000000
0#
0(
#212340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#212390000000
0$
0)
#212400000000
1"
1'
b0 +
b0 1
#212450000000
0"
0'
#212460000000
1#
1(
b101111101100100 +
b101111101100100 1
#212510000000
0#
0(
#212520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#212570000000
0$
0)
#212580000000
1"
1'
b0 +
b0 1
#212630000000
0"
0'
#212640000000
1#
1(
b101111101100100 +
b101111101100100 1
#212690000000
0#
0(
#212700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#212750000000
0$
0)
#212760000000
1"
1'
b0 +
b0 1
#212810000000
0"
0'
#212820000000
1#
1(
b101111101100100 +
b101111101100100 1
#212870000000
0#
0(
#212880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#212930000000
0$
0)
#212940000000
1"
1'
b0 +
b0 1
#212990000000
0"
0'
#213000000000
1#
1(
b101111101100100 +
b101111101100100 1
#213050000000
0#
0(
#213060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#213110000000
0$
0)
#213120000000
1"
1'
b0 +
b0 1
#213170000000
0"
0'
#213180000000
1#
1(
b101111101100100 +
b101111101100100 1
#213230000000
0#
0(
#213240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#213290000000
0$
0)
#213300000000
1"
1'
b0 +
b0 1
#213350000000
0"
0'
#213360000000
1#
1(
b101111101100100 +
b101111101100100 1
#213410000000
0#
0(
#213420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#213470000000
0$
0)
#213480000000
1"
1'
b0 +
b0 1
#213530000000
0"
0'
#213540000000
1#
1(
b101111101100100 +
b101111101100100 1
#213590000000
0#
0(
#213600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#213650000000
0$
0)
#213660000000
1"
1'
b0 +
b0 1
#213710000000
0"
0'
#213720000000
1#
1(
b101111101100100 +
b101111101100100 1
#213770000000
0#
0(
#213780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#213830000000
0$
0)
#213840000000
1"
1'
b0 +
b0 1
#213890000000
0"
0'
#213900000000
1#
1(
b101111101100100 +
b101111101100100 1
#213950000000
0#
0(
#213960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#214010000000
0$
0)
#214020000000
1"
1'
b0 +
b0 1
#214070000000
0"
0'
#214080000000
1#
1(
b101111101100100 +
b101111101100100 1
#214130000000
0#
0(
#214140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#214190000000
0$
0)
#214200000000
1"
1'
b0 +
b0 1
#214250000000
0"
0'
#214260000000
1#
1(
b101111101100100 +
b101111101100100 1
#214310000000
0#
0(
#214320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#214370000000
0$
0)
#214380000000
1"
1'
b0 +
b0 1
#214430000000
0"
0'
#214440000000
1#
1(
b101111101100100 +
b101111101100100 1
#214490000000
0#
0(
#214500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#214550000000
0$
0)
#214560000000
1"
1'
b0 +
b0 1
#214610000000
0"
0'
#214620000000
1#
1(
b101111101100100 +
b101111101100100 1
#214670000000
0#
0(
#214680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#214730000000
0$
0)
#214740000000
1"
1'
b0 +
b0 1
#214790000000
0"
0'
#214800000000
1#
1(
b101111101100100 +
b101111101100100 1
#214850000000
0#
0(
#214860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#214910000000
0$
0)
#214920000000
1"
1'
b0 +
b0 1
#214970000000
0"
0'
#214980000000
1#
1(
b101111101100100 +
b101111101100100 1
#215030000000
0#
0(
#215040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#215090000000
0$
0)
#215100000000
1"
1'
b0 +
b0 1
#215150000000
0"
0'
#215160000000
1#
1(
b101111101100100 +
b101111101100100 1
#215210000000
0#
0(
#215220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#215270000000
0$
0)
#215280000000
1"
1'
b0 +
b0 1
#215330000000
0"
0'
#215340000000
1#
1(
b101111101100100 +
b101111101100100 1
#215390000000
0#
0(
#215400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#215450000000
0$
0)
#215460000000
1"
1'
b0 +
b0 1
#215510000000
0"
0'
#215520000000
1#
1(
b101111101100100 +
b101111101100100 1
#215570000000
0#
0(
#215580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#215630000000
0$
0)
#215640000000
1"
1'
b0 +
b0 1
#215690000000
0"
0'
#215700000000
1#
1(
b101111101100100 +
b101111101100100 1
#215750000000
0#
0(
#215760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#215810000000
0$
0)
#215820000000
1"
1'
b0 +
b0 1
#215870000000
0"
0'
#215880000000
1#
1(
b101111101100100 +
b101111101100100 1
#215930000000
0#
0(
#215940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#215990000000
0$
0)
#216000000000
1"
1'
b0 +
b0 1
#216050000000
0"
0'
#216060000000
1#
1(
b101111101100100 +
b101111101100100 1
#216110000000
0#
0(
#216120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#216170000000
0$
0)
#216180000000
1"
1'
b0 +
b0 1
#216230000000
0"
0'
#216240000000
1#
1(
b101111101100100 +
b101111101100100 1
#216290000000
0#
0(
#216300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#216350000000
0$
0)
#216360000000
1"
1'
b0 +
b0 1
#216410000000
0"
0'
#216420000000
1#
1(
b101111101100100 +
b101111101100100 1
#216470000000
0#
0(
#216480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#216530000000
0$
0)
#216540000000
1"
1'
b0 +
b0 1
#216590000000
0"
0'
#216600000000
1#
1(
b101111101100100 +
b101111101100100 1
#216650000000
0#
0(
#216660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#216710000000
0$
0)
#216720000000
1"
1'
b0 +
b0 1
#216770000000
0"
0'
#216780000000
1#
1(
b101111101100100 +
b101111101100100 1
#216830000000
0#
0(
#216840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#216890000000
0$
0)
#216900000000
1"
1'
b0 +
b0 1
#216950000000
0"
0'
#216960000000
1#
1(
b101111101100100 +
b101111101100100 1
#217010000000
0#
0(
#217020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#217070000000
0$
0)
#217080000000
1"
1'
b0 +
b0 1
#217130000000
0"
0'
#217140000000
1#
1(
b101111101100100 +
b101111101100100 1
#217190000000
0#
0(
#217200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#217250000000
0$
0)
#217260000000
1"
1'
b0 +
b0 1
#217310000000
0"
0'
#217320000000
1#
1(
b101111101100100 +
b101111101100100 1
#217370000000
0#
0(
#217380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#217430000000
0$
0)
#217440000000
1"
1'
b0 +
b0 1
#217490000000
0"
0'
#217500000000
1#
1(
b101111101100100 +
b101111101100100 1
#217550000000
0#
0(
#217560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#217610000000
0$
0)
#217620000000
1"
1'
b0 +
b0 1
#217670000000
0"
0'
#217680000000
1#
1(
b101111101100100 +
b101111101100100 1
#217730000000
0#
0(
#217740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#217790000000
0$
0)
#217800000000
1"
1'
b0 +
b0 1
#217850000000
0"
0'
#217860000000
1#
1(
b101111101100100 +
b101111101100100 1
#217910000000
0#
0(
#217920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#217970000000
0$
0)
#217980000000
1"
1'
b0 +
b0 1
#218030000000
0"
0'
#218040000000
1#
1(
b101111101100100 +
b101111101100100 1
#218090000000
0#
0(
#218100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#218150000000
0$
0)
#218160000000
1"
1'
b0 +
b0 1
#218210000000
0"
0'
#218220000000
1#
1(
b101111101100100 +
b101111101100100 1
#218270000000
0#
0(
#218280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#218330000000
0$
0)
#218340000000
1"
1'
b0 +
b0 1
#218390000000
0"
0'
#218400000000
1#
1(
b101111101100100 +
b101111101100100 1
#218450000000
0#
0(
#218460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#218510000000
0$
0)
#218520000000
1"
1'
b0 +
b0 1
#218570000000
0"
0'
#218580000000
1#
1(
b101111101100100 +
b101111101100100 1
#218630000000
0#
0(
#218640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#218690000000
0$
0)
#218700000000
1"
1'
b0 +
b0 1
#218750000000
0"
0'
#218760000000
1#
1(
b101111101100100 +
b101111101100100 1
#218810000000
0#
0(
#218820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#218870000000
0$
0)
#218880000000
1"
1'
b0 +
b0 1
#218930000000
0"
0'
#218940000000
1#
1(
b101111101100100 +
b101111101100100 1
#218990000000
0#
0(
#219000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#219050000000
0$
0)
#219060000000
1"
1'
b0 +
b0 1
#219110000000
0"
0'
#219120000000
1#
1(
b101111101100100 +
b101111101100100 1
#219170000000
0#
0(
#219180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#219230000000
0$
0)
#219240000000
1"
1'
b0 +
b0 1
#219290000000
0"
0'
#219300000000
1#
1(
b101111101100100 +
b101111101100100 1
#219350000000
0#
0(
#219360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#219410000000
0$
0)
#219420000000
1"
1'
b0 +
b0 1
#219470000000
0"
0'
#219480000000
1#
1(
b101111101100100 +
b101111101100100 1
#219530000000
0#
0(
#219540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#219590000000
0$
0)
#219600000000
1"
1'
b0 +
b0 1
#219650000000
0"
0'
#219660000000
1#
1(
b101111101100100 +
b101111101100100 1
#219710000000
0#
0(
#219720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#219770000000
0$
0)
#219780000000
1"
1'
b0 +
b0 1
#219830000000
0"
0'
#219840000000
1#
1(
b101111101100100 +
b101111101100100 1
#219890000000
0#
0(
#219900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#219950000000
0$
0)
#219960000000
1"
1'
b0 +
b0 1
#220010000000
0"
0'
#220020000000
1#
1(
b101111101100100 +
b101111101100100 1
#220070000000
0#
0(
#220080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#220130000000
0$
0)
#220140000000
1"
1'
b0 +
b0 1
#220190000000
0"
0'
#220200000000
1#
1(
b101111101100100 +
b101111101100100 1
#220250000000
0#
0(
#220260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#220310000000
0$
0)
#220320000000
1"
1'
b0 +
b0 1
#220370000000
0"
0'
#220380000000
1#
1(
b101111101100100 +
b101111101100100 1
#220430000000
0#
0(
#220440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#220490000000
0$
0)
#220500000000
1"
1'
b0 +
b0 1
#220550000000
0"
0'
#220560000000
1#
1(
b101111101100100 +
b101111101100100 1
#220610000000
0#
0(
#220620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#220670000000
0$
0)
#220680000000
1"
1'
b0 +
b0 1
#220730000000
0"
0'
#220740000000
1#
1(
b101111101100100 +
b101111101100100 1
#220790000000
0#
0(
#220800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#220850000000
0$
0)
#220860000000
1"
1'
b0 +
b0 1
#220910000000
0"
0'
#220920000000
1#
1(
b101111101100100 +
b101111101100100 1
#220970000000
0#
0(
#220980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#221030000000
0$
0)
#221040000000
1"
1'
b0 +
b0 1
#221090000000
0"
0'
#221100000000
1#
1(
b101111101100100 +
b101111101100100 1
#221150000000
0#
0(
#221160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#221210000000
0$
0)
#221220000000
1"
1'
b0 +
b0 1
#221270000000
0"
0'
#221280000000
1#
1(
b101111101100100 +
b101111101100100 1
#221330000000
0#
0(
#221340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#221390000000
0$
0)
#221400000000
1"
1'
b0 +
b0 1
#221450000000
0"
0'
#221460000000
1#
1(
b101111101100100 +
b101111101100100 1
#221510000000
0#
0(
#221520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#221570000000
0$
0)
#221580000000
1"
1'
b0 +
b0 1
#221630000000
0"
0'
#221640000000
1#
1(
b101111101100100 +
b101111101100100 1
#221690000000
0#
0(
#221700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#221750000000
0$
0)
#221760000000
1"
1'
b0 +
b0 1
#221810000000
0"
0'
#221820000000
1#
1(
b101111101100100 +
b101111101100100 1
#221870000000
0#
0(
#221880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#221930000000
0$
0)
#221940000000
1"
1'
b0 +
b0 1
#221990000000
0"
0'
#222000000000
1#
1(
b101111101100100 +
b101111101100100 1
#222050000000
0#
0(
#222060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#222110000000
0$
0)
#222120000000
1"
1'
b0 +
b0 1
#222170000000
0"
0'
#222180000000
1#
1(
b101111101100100 +
b101111101100100 1
#222230000000
0#
0(
#222240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#222290000000
0$
0)
#222300000000
1"
1'
b0 +
b0 1
#222350000000
0"
0'
#222360000000
1#
1(
b101111101100100 +
b101111101100100 1
#222410000000
0#
0(
#222420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#222470000000
0$
0)
#222480000000
1"
1'
b0 +
b0 1
#222530000000
0"
0'
#222540000000
1#
1(
b101111101100100 +
b101111101100100 1
#222590000000
0#
0(
#222600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#222650000000
0$
0)
#222660000000
1"
1'
b0 +
b0 1
#222710000000
0"
0'
#222720000000
1#
1(
b101111101100100 +
b101111101100100 1
#222770000000
0#
0(
#222780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#222830000000
0$
0)
#222840000000
1"
1'
b0 +
b0 1
#222890000000
0"
0'
#222900000000
1#
1(
b101111101100100 +
b101111101100100 1
#222950000000
0#
0(
#222960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#223010000000
0$
0)
#223020000000
1"
1'
b0 +
b0 1
#223070000000
0"
0'
#223080000000
1#
1(
b101111101100100 +
b101111101100100 1
#223130000000
0#
0(
#223140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#223190000000
0$
0)
#223200000000
1"
1'
b0 +
b0 1
#223250000000
0"
0'
#223260000000
1#
1(
b101111101100100 +
b101111101100100 1
#223310000000
0#
0(
#223320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#223370000000
0$
0)
#223380000000
1"
1'
b0 +
b0 1
#223430000000
0"
0'
#223440000000
1#
1(
b101111101100100 +
b101111101100100 1
#223490000000
0#
0(
#223500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#223550000000
0$
0)
#223560000000
1"
1'
b0 +
b0 1
#223610000000
0"
0'
#223620000000
1#
1(
b101111101100100 +
b101111101100100 1
#223670000000
0#
0(
#223680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#223730000000
0$
0)
#223740000000
1"
1'
b0 +
b0 1
#223790000000
0"
0'
#223800000000
1#
1(
b101111101100100 +
b101111101100100 1
#223850000000
0#
0(
#223860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#223910000000
0$
0)
#223920000000
1"
1'
b0 +
b0 1
#223970000000
0"
0'
#223980000000
1#
1(
b101111101100100 +
b101111101100100 1
#224030000000
0#
0(
#224040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#224090000000
0$
0)
#224100000000
1"
1'
b0 +
b0 1
#224150000000
0"
0'
#224160000000
1#
1(
b101111101100100 +
b101111101100100 1
#224210000000
0#
0(
#224220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#224270000000
0$
0)
#224280000000
1"
1'
b0 +
b0 1
#224330000000
0"
0'
#224340000000
1#
1(
b101111101100100 +
b101111101100100 1
#224390000000
0#
0(
#224400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#224450000000
0$
0)
#224460000000
1"
1'
b0 +
b0 1
#224510000000
0"
0'
#224520000000
1#
1(
b101111101100100 +
b101111101100100 1
#224570000000
0#
0(
#224580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#224630000000
0$
0)
#224640000000
1"
1'
b0 +
b0 1
#224690000000
0"
0'
#224700000000
1#
1(
b101111101100100 +
b101111101100100 1
#224750000000
0#
0(
#224760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#224810000000
0$
0)
#224820000000
1"
1'
b0 +
b0 1
#224870000000
0"
0'
#224880000000
1#
1(
b101111101100100 +
b101111101100100 1
#224930000000
0#
0(
#224940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#224990000000
0$
0)
#225000000000
1"
1'
b0 +
b0 1
#225050000000
0"
0'
#225060000000
1#
1(
b101111101100100 +
b101111101100100 1
#225110000000
0#
0(
#225120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#225170000000
0$
0)
#225180000000
1"
1'
b0 +
b0 1
#225230000000
0"
0'
#225240000000
1#
1(
b101111101100100 +
b101111101100100 1
#225290000000
0#
0(
#225300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#225350000000
0$
0)
#225360000000
1"
1'
b0 +
b0 1
#225410000000
0"
0'
#225420000000
1#
1(
b101111101100100 +
b101111101100100 1
#225470000000
0#
0(
#225480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#225530000000
0$
0)
#225540000000
1"
1'
b0 +
b0 1
#225590000000
0"
0'
#225600000000
1#
1(
b101111101100100 +
b101111101100100 1
#225650000000
0#
0(
#225660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#225710000000
0$
0)
#225720000000
1"
1'
b0 +
b0 1
#225770000000
0"
0'
#225780000000
1#
1(
b101111101100100 +
b101111101100100 1
#225830000000
0#
0(
#225840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#225890000000
0$
0)
#225900000000
1"
1'
b0 +
b0 1
#225950000000
0"
0'
#225960000000
1#
1(
b101111101100100 +
b101111101100100 1
#226010000000
0#
0(
#226020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#226070000000
0$
0)
#226080000000
1"
1'
b0 +
b0 1
#226130000000
0"
0'
#226140000000
1#
1(
b101111101100100 +
b101111101100100 1
#226190000000
0#
0(
#226200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#226250000000
0$
0)
#226260000000
1"
1'
b0 +
b0 1
#226310000000
0"
0'
#226320000000
1#
1(
b101111101100100 +
b101111101100100 1
#226370000000
0#
0(
#226380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#226430000000
0$
0)
#226440000000
1"
1'
b0 +
b0 1
#226490000000
0"
0'
#226500000000
1#
1(
b101111101100100 +
b101111101100100 1
#226550000000
0#
0(
#226560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#226610000000
0$
0)
#226620000000
1"
1'
b0 +
b0 1
#226670000000
0"
0'
#226680000000
1#
1(
b101111101100100 +
b101111101100100 1
#226730000000
0#
0(
#226740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#226790000000
0$
0)
#226800000000
1"
1'
b0 +
b0 1
#226850000000
0"
0'
#226860000000
1#
1(
b101111101100100 +
b101111101100100 1
#226910000000
0#
0(
#226920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#226970000000
0$
0)
#226980000000
1"
1'
b0 +
b0 1
#227030000000
0"
0'
#227040000000
1#
1(
b101111101100100 +
b101111101100100 1
#227090000000
0#
0(
#227100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#227150000000
0$
0)
#227160000000
1"
1'
b0 +
b0 1
#227210000000
0"
0'
#227220000000
1#
1(
b101111101100100 +
b101111101100100 1
#227270000000
0#
0(
#227280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#227330000000
0$
0)
#227340000000
1"
1'
b0 +
b0 1
#227390000000
0"
0'
#227400000000
1#
1(
b101111101100100 +
b101111101100100 1
#227450000000
0#
0(
#227460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#227510000000
0$
0)
#227520000000
1"
1'
b0 +
b0 1
#227570000000
0"
0'
#227580000000
1#
1(
b101111101100100 +
b101111101100100 1
#227630000000
0#
0(
#227640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#227690000000
0$
0)
#227700000000
1"
1'
b0 +
b0 1
#227750000000
0"
0'
#227760000000
1#
1(
b101111101100100 +
b101111101100100 1
#227810000000
0#
0(
#227820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#227870000000
0$
0)
#227880000000
1"
1'
b0 +
b0 1
#227930000000
0"
0'
#227940000000
1#
1(
b101111101100100 +
b101111101100100 1
#227990000000
0#
0(
#228000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#228050000000
0$
0)
#228060000000
1"
1'
b0 +
b0 1
#228110000000
0"
0'
#228120000000
1#
1(
b101111101100100 +
b101111101100100 1
#228170000000
0#
0(
#228180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#228230000000
0$
0)
#228240000000
1"
1'
b0 +
b0 1
#228290000000
0"
0'
#228300000000
1#
1(
b101111101100100 +
b101111101100100 1
#228350000000
0#
0(
#228360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#228410000000
0$
0)
#228420000000
1"
1'
b0 +
b0 1
#228470000000
0"
0'
#228480000000
1#
1(
b101111101100100 +
b101111101100100 1
#228530000000
0#
0(
#228540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#228590000000
0$
0)
#228600000000
1"
1'
b0 +
b0 1
#228650000000
0"
0'
#228660000000
1#
1(
b101111101100100 +
b101111101100100 1
#228710000000
0#
0(
#228720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#228770000000
0$
0)
#228780000000
1"
1'
b0 +
b0 1
#228830000000
0"
0'
#228840000000
1#
1(
b101111101100100 +
b101111101100100 1
#228890000000
0#
0(
#228900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#228950000000
0$
0)
#228960000000
1"
1'
b0 +
b0 1
#229010000000
0"
0'
#229020000000
1#
1(
b101111101100100 +
b101111101100100 1
#229070000000
0#
0(
#229080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#229130000000
0$
0)
#229140000000
1"
1'
b0 +
b0 1
#229190000000
0"
0'
#229200000000
1#
1(
b101111101100100 +
b101111101100100 1
#229250000000
0#
0(
#229260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#229310000000
0$
0)
#229320000000
1"
1'
b0 +
b0 1
#229370000000
0"
0'
#229380000000
1#
1(
b101111101100100 +
b101111101100100 1
#229430000000
0#
0(
#229440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#229490000000
0$
0)
#229500000000
1"
1'
b0 +
b0 1
#229550000000
0"
0'
#229560000000
1#
1(
b101111101100100 +
b101111101100100 1
#229610000000
0#
0(
#229620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#229670000000
0$
0)
#229680000000
1"
1'
b0 +
b0 1
#229730000000
0"
0'
#229740000000
1#
1(
b101111101100100 +
b101111101100100 1
#229790000000
0#
0(
#229800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#229850000000
0$
0)
#229860000000
1"
1'
b0 +
b0 1
#229910000000
0"
0'
#229920000000
1#
1(
b101111101100100 +
b101111101100100 1
#229970000000
0#
0(
#229980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#230030000000
0$
0)
#230040000000
1"
1'
b0 +
b0 1
#230090000000
0"
0'
#230100000000
1#
1(
b101111101100100 +
b101111101100100 1
#230150000000
0#
0(
#230160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#230210000000
0$
0)
#230220000000
1"
1'
b0 +
b0 1
#230270000000
0"
0'
#230280000000
1#
1(
b101111101100100 +
b101111101100100 1
#230330000000
0#
0(
#230340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#230390000000
0$
0)
#230400000000
1"
1'
b0 +
b0 1
#230450000000
0"
0'
#230460000000
1#
1(
b101111101100100 +
b101111101100100 1
#230510000000
0#
0(
#230520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#230570000000
0$
0)
#230580000000
1"
1'
b0 +
b0 1
#230630000000
0"
0'
#230640000000
1#
1(
b101111101100100 +
b101111101100100 1
#230690000000
0#
0(
#230700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#230750000000
0$
0)
#230760000000
1"
1'
b0 +
b0 1
#230810000000
0"
0'
#230820000000
1#
1(
b101111101100100 +
b101111101100100 1
#230870000000
0#
0(
#230880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#230930000000
0$
0)
#230940000000
1"
1'
b0 +
b0 1
#230990000000
0"
0'
#231000000000
1#
1(
b101111101100100 +
b101111101100100 1
#231050000000
0#
0(
#231060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#231110000000
0$
0)
#231120000000
1"
1'
b0 +
b0 1
#231170000000
0"
0'
#231180000000
1#
1(
b101111101100100 +
b101111101100100 1
#231230000000
0#
0(
#231240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#231290000000
0$
0)
#231300000000
1"
1'
b0 +
b0 1
#231350000000
0"
0'
#231360000000
1#
1(
b101111101100100 +
b101111101100100 1
#231410000000
0#
0(
#231420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#231470000000
0$
0)
#231480000000
1"
1'
b0 +
b0 1
#231530000000
0"
0'
#231540000000
1#
1(
b101111101100100 +
b101111101100100 1
#231590000000
0#
0(
#231600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#231650000000
0$
0)
#231660000000
1"
1'
b0 +
b0 1
#231710000000
0"
0'
#231720000000
1#
1(
b101111101100100 +
b101111101100100 1
#231770000000
0#
0(
#231780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#231830000000
0$
0)
#231840000000
1"
1'
b0 +
b0 1
#231890000000
0"
0'
#231900000000
1#
1(
b101111101100100 +
b101111101100100 1
#231950000000
0#
0(
#231960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#232010000000
0$
0)
#232020000000
1"
1'
b0 +
b0 1
#232070000000
0"
0'
#232080000000
1#
1(
b101111101100100 +
b101111101100100 1
#232130000000
0#
0(
#232140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#232190000000
0$
0)
#232200000000
1"
1'
b0 +
b0 1
#232250000000
0"
0'
#232260000000
1#
1(
b101111101100100 +
b101111101100100 1
#232310000000
0#
0(
#232320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#232370000000
0$
0)
#232380000000
1"
1'
b0 +
b0 1
#232430000000
0"
0'
#232440000000
1#
1(
b101111101100100 +
b101111101100100 1
#232490000000
0#
0(
#232500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#232550000000
0$
0)
#232560000000
1"
1'
b0 +
b0 1
#232610000000
0"
0'
#232620000000
1#
1(
b101111101100100 +
b101111101100100 1
#232670000000
0#
0(
#232680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#232730000000
0$
0)
#232740000000
1"
1'
b0 +
b0 1
#232790000000
0"
0'
#232800000000
1#
1(
b101111101100100 +
b101111101100100 1
#232850000000
0#
0(
#232860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#232910000000
0$
0)
#232920000000
1"
1'
b0 +
b0 1
#232970000000
0"
0'
#232980000000
1#
1(
b101111101100100 +
b101111101100100 1
#233030000000
0#
0(
#233040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#233090000000
0$
0)
#233100000000
1"
1'
b0 +
b0 1
#233150000000
0"
0'
#233160000000
1#
1(
b101111101100100 +
b101111101100100 1
#233210000000
0#
0(
#233220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#233270000000
0$
0)
#233280000000
1"
1'
b0 +
b0 1
#233330000000
0"
0'
#233340000000
1#
1(
b101111101100100 +
b101111101100100 1
#233390000000
0#
0(
#233400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#233450000000
0$
0)
#233460000000
1"
1'
b0 +
b0 1
#233510000000
0"
0'
#233520000000
1#
1(
b101111101100100 +
b101111101100100 1
#233570000000
0#
0(
#233580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#233630000000
0$
0)
#233640000000
1"
1'
b0 +
b0 1
#233690000000
0"
0'
#233700000000
1#
1(
b101111101100100 +
b101111101100100 1
#233750000000
0#
0(
#233760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#233810000000
0$
0)
#233820000000
1"
1'
b0 +
b0 1
#233870000000
0"
0'
#233880000000
1#
1(
b101111101100100 +
b101111101100100 1
#233930000000
0#
0(
#233940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#233990000000
0$
0)
#234000000000
1"
1'
b0 +
b0 1
#234050000000
0"
0'
#234060000000
1#
1(
b101111101100100 +
b101111101100100 1
#234110000000
0#
0(
#234120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#234170000000
0$
0)
#234180000000
1"
1'
b0 +
b0 1
#234230000000
0"
0'
#234240000000
1#
1(
b101111101100100 +
b101111101100100 1
#234290000000
0#
0(
#234300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#234350000000
0$
0)
#234360000000
1"
1'
b0 +
b0 1
#234410000000
0"
0'
#234420000000
1#
1(
b101111101100100 +
b101111101100100 1
#234470000000
0#
0(
#234480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#234530000000
0$
0)
#234540000000
1"
1'
b0 +
b0 1
#234590000000
0"
0'
#234600000000
1#
1(
b101111101100100 +
b101111101100100 1
#234650000000
0#
0(
#234660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#234710000000
0$
0)
#234720000000
1"
1'
b0 +
b0 1
#234770000000
0"
0'
#234780000000
1#
1(
b101111101100100 +
b101111101100100 1
#234830000000
0#
0(
#234840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#234890000000
0$
0)
#234900000000
1"
1'
b0 +
b0 1
#234950000000
0"
0'
#234960000000
1#
1(
b101111101100100 +
b101111101100100 1
#235010000000
0#
0(
#235020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#235070000000
0$
0)
#235080000000
1"
1'
b0 +
b0 1
#235130000000
0"
0'
#235140000000
1#
1(
b101111101100100 +
b101111101100100 1
#235190000000
0#
0(
#235200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#235250000000
0$
0)
#235260000000
1"
1'
b0 +
b0 1
#235310000000
0"
0'
#235320000000
1#
1(
b101111101100100 +
b101111101100100 1
#235370000000
0#
0(
#235380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#235430000000
0$
0)
#235440000000
1"
1'
b0 +
b0 1
#235490000000
0"
0'
#235500000000
1#
1(
b101111101100100 +
b101111101100100 1
#235550000000
0#
0(
#235560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#235610000000
0$
0)
#235620000000
1"
1'
b0 +
b0 1
#235670000000
0"
0'
#235680000000
1#
1(
b101111101100100 +
b101111101100100 1
#235730000000
0#
0(
#235740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#235790000000
0$
0)
#235800000000
1"
1'
b0 +
b0 1
#235850000000
0"
0'
#235860000000
1#
1(
b101111101100100 +
b101111101100100 1
#235910000000
0#
0(
#235920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#235970000000
0$
0)
#235980000000
1"
1'
b0 +
b0 1
#236030000000
0"
0'
#236040000000
1#
1(
b101111101100100 +
b101111101100100 1
#236090000000
0#
0(
#236100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#236150000000
0$
0)
#236160000000
1"
1'
b0 +
b0 1
#236210000000
0"
0'
#236220000000
1#
1(
b101111101100100 +
b101111101100100 1
#236270000000
0#
0(
#236280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#236330000000
0$
0)
#236340000000
1"
1'
b0 +
b0 1
#236390000000
0"
0'
#236400000000
1#
1(
b101111101100100 +
b101111101100100 1
#236450000000
0#
0(
#236460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#236510000000
0$
0)
#236520000000
1"
1'
b0 +
b0 1
#236570000000
0"
0'
#236580000000
1#
1(
b101111101100100 +
b101111101100100 1
#236630000000
0#
0(
#236640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#236690000000
0$
0)
#236700000000
1"
1'
b0 +
b0 1
#236750000000
0"
0'
#236760000000
1#
1(
b101111101100100 +
b101111101100100 1
#236810000000
0#
0(
#236820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#236870000000
0$
0)
#236880000000
1"
1'
b0 +
b0 1
#236930000000
0"
0'
#236940000000
1#
1(
b101111101100100 +
b101111101100100 1
#236990000000
0#
0(
#237000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#237050000000
0$
0)
#237060000000
1"
1'
b0 +
b0 1
#237110000000
0"
0'
#237120000000
1#
1(
b101111101100100 +
b101111101100100 1
#237170000000
0#
0(
#237180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#237230000000
0$
0)
#237240000000
1"
1'
b0 +
b0 1
#237290000000
0"
0'
#237300000000
1#
1(
b101111101100100 +
b101111101100100 1
#237350000000
0#
0(
#237360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#237410000000
0$
0)
#237420000000
1"
1'
b0 +
b0 1
#237470000000
0"
0'
#237480000000
1#
1(
b101111101100100 +
b101111101100100 1
#237530000000
0#
0(
#237540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#237590000000
0$
0)
#237600000000
1"
1'
b0 +
b0 1
#237650000000
0"
0'
#237660000000
1#
1(
b101111101100100 +
b101111101100100 1
#237710000000
0#
0(
#237720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#237770000000
0$
0)
#237780000000
1"
1'
b0 +
b0 1
#237830000000
0"
0'
#237840000000
1#
1(
b101111101100100 +
b101111101100100 1
#237890000000
0#
0(
#237900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#237950000000
0$
0)
#237960000000
1"
1'
b0 +
b0 1
#238010000000
0"
0'
#238020000000
1#
1(
b101111101100100 +
b101111101100100 1
#238070000000
0#
0(
#238080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#238130000000
0$
0)
#238140000000
1"
1'
b0 +
b0 1
#238190000000
0"
0'
#238200000000
1#
1(
b101111101100100 +
b101111101100100 1
#238250000000
0#
0(
#238260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#238310000000
0$
0)
#238320000000
1"
1'
b0 +
b0 1
#238370000000
0"
0'
#238380000000
1#
1(
b101111101100100 +
b101111101100100 1
#238430000000
0#
0(
#238440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#238490000000
0$
0)
#238500000000
1"
1'
b0 +
b0 1
#238550000000
0"
0'
#238560000000
1#
1(
b101111101100100 +
b101111101100100 1
#238610000000
0#
0(
#238620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#238670000000
0$
0)
#238680000000
1"
1'
b0 +
b0 1
#238730000000
0"
0'
#238740000000
1#
1(
b101111101100100 +
b101111101100100 1
#238790000000
0#
0(
#238800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#238850000000
0$
0)
#238860000000
1"
1'
b0 +
b0 1
#238910000000
0"
0'
#238920000000
1#
1(
b101111101100100 +
b101111101100100 1
#238970000000
0#
0(
#238980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#239030000000
0$
0)
#239040000000
1"
1'
b0 +
b0 1
#239090000000
0"
0'
#239100000000
1#
1(
b101111101100100 +
b101111101100100 1
#239150000000
0#
0(
#239160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#239210000000
0$
0)
#239220000000
1"
1'
b0 +
b0 1
#239270000000
0"
0'
#239280000000
1#
1(
b101111101100100 +
b101111101100100 1
#239330000000
0#
0(
#239340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#239390000000
0$
0)
#239400000000
1"
1'
b0 +
b0 1
#239450000000
0"
0'
#239460000000
1#
1(
b101111101100100 +
b101111101100100 1
#239510000000
0#
0(
#239520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#239570000000
0$
0)
#239580000000
1"
1'
b0 +
b0 1
#239630000000
0"
0'
#239640000000
1#
1(
b101111101100100 +
b101111101100100 1
#239690000000
0#
0(
#239700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#239750000000
0$
0)
#239760000000
1"
1'
b0 +
b0 1
#239810000000
0"
0'
#239820000000
1#
1(
b101111101100100 +
b101111101100100 1
#239870000000
0#
0(
#239880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#239930000000
0$
0)
#239940000000
1"
1'
b0 +
b0 1
#239990000000
0"
0'
#240000000000
1#
1(
b101111101100100 +
b101111101100100 1
#240050000000
0#
0(
#240060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#240110000000
0$
0)
#240120000000
1"
1'
b0 +
b0 1
#240170000000
0"
0'
#240180000000
1#
1(
b101111101100100 +
b101111101100100 1
#240230000000
0#
0(
#240240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#240290000000
0$
0)
#240300000000
1"
1'
b0 +
b0 1
#240350000000
0"
0'
#240360000000
1#
1(
b101111101100100 +
b101111101100100 1
#240410000000
0#
0(
#240420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#240470000000
0$
0)
#240480000000
1"
1'
b0 +
b0 1
#240530000000
0"
0'
#240540000000
1#
1(
b101111101100100 +
b101111101100100 1
#240590000000
0#
0(
#240600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#240650000000
0$
0)
#240660000000
1"
1'
b0 +
b0 1
#240710000000
0"
0'
#240720000000
1#
1(
b101111101100100 +
b101111101100100 1
#240770000000
0#
0(
#240780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#240830000000
0$
0)
#240840000000
1"
1'
b0 +
b0 1
#240890000000
0"
0'
#240900000000
1#
1(
b101111101100100 +
b101111101100100 1
#240950000000
0#
0(
#240960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#241010000000
0$
0)
#241020000000
1"
1'
b0 +
b0 1
#241070000000
0"
0'
#241080000000
1#
1(
b101111101100100 +
b101111101100100 1
#241130000000
0#
0(
#241140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#241190000000
0$
0)
#241200000000
1"
1'
b0 +
b0 1
#241250000000
0"
0'
#241260000000
1#
1(
b101111101100100 +
b101111101100100 1
#241310000000
0#
0(
#241320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#241370000000
0$
0)
#241380000000
1"
1'
b0 +
b0 1
#241430000000
0"
0'
#241440000000
1#
1(
b101111101100100 +
b101111101100100 1
#241490000000
0#
0(
#241500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#241550000000
0$
0)
#241560000000
1"
1'
b0 +
b0 1
#241610000000
0"
0'
#241620000000
1#
1(
b101111101100100 +
b101111101100100 1
#241670000000
0#
0(
#241680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#241730000000
0$
0)
#241740000000
1"
1'
b0 +
b0 1
#241790000000
0"
0'
#241800000000
1#
1(
b101111101100100 +
b101111101100100 1
#241850000000
0#
0(
#241860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#241910000000
0$
0)
#241920000000
1"
1'
b0 +
b0 1
#241970000000
0"
0'
#241980000000
1#
1(
b101111101100100 +
b101111101100100 1
#242030000000
0#
0(
#242040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#242090000000
0$
0)
#242100000000
1"
1'
b0 +
b0 1
#242150000000
0"
0'
#242160000000
1#
1(
b101111101100100 +
b101111101100100 1
#242210000000
0#
0(
#242220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#242270000000
0$
0)
#242280000000
1"
1'
b0 +
b0 1
#242330000000
0"
0'
#242340000000
1#
1(
b101111101100100 +
b101111101100100 1
#242390000000
0#
0(
#242400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#242450000000
0$
0)
#242460000000
1"
1'
b0 +
b0 1
#242510000000
0"
0'
#242520000000
1#
1(
b101111101100100 +
b101111101100100 1
#242570000000
0#
0(
#242580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#242630000000
0$
0)
#242640000000
1"
1'
b0 +
b0 1
#242690000000
0"
0'
#242700000000
1#
1(
b101111101100100 +
b101111101100100 1
#242750000000
0#
0(
#242760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#242810000000
0$
0)
#242820000000
1"
1'
b0 +
b0 1
#242870000000
0"
0'
#242880000000
1#
1(
b101111101100100 +
b101111101100100 1
#242930000000
0#
0(
#242940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#242990000000
0$
0)
#243000000000
1"
1'
b0 +
b0 1
#243050000000
0"
0'
#243060000000
1#
1(
b101111101100100 +
b101111101100100 1
#243110000000
0#
0(
#243120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#243170000000
0$
0)
#243180000000
1"
1'
b0 +
b0 1
#243230000000
0"
0'
#243240000000
1#
1(
b101111101100100 +
b101111101100100 1
#243290000000
0#
0(
#243300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#243350000000
0$
0)
#243360000000
1"
1'
b0 +
b0 1
#243410000000
0"
0'
#243420000000
1#
1(
b101111101100100 +
b101111101100100 1
#243470000000
0#
0(
#243480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#243530000000
0$
0)
#243540000000
1"
1'
b0 +
b0 1
#243590000000
0"
0'
#243600000000
1#
1(
b101111101100100 +
b101111101100100 1
#243650000000
0#
0(
#243660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#243710000000
0$
0)
#243720000000
1"
1'
b0 +
b0 1
#243770000000
0"
0'
#243780000000
1#
1(
b101111101100100 +
b101111101100100 1
#243830000000
0#
0(
#243840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#243890000000
0$
0)
#243900000000
1"
1'
b0 +
b0 1
#243950000000
0"
0'
#243960000000
1#
1(
b101111101100100 +
b101111101100100 1
#244010000000
0#
0(
#244020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#244070000000
0$
0)
#244080000000
1"
1'
b0 +
b0 1
#244130000000
0"
0'
#244140000000
1#
1(
b101111101100100 +
b101111101100100 1
#244190000000
0#
0(
#244200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#244250000000
0$
0)
#244260000000
1"
1'
b0 +
b0 1
#244310000000
0"
0'
#244320000000
1#
1(
b101111101100100 +
b101111101100100 1
#244370000000
0#
0(
#244380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#244430000000
0$
0)
#244440000000
1"
1'
b0 +
b0 1
#244490000000
0"
0'
#244500000000
1#
1(
b101111101100100 +
b101111101100100 1
#244550000000
0#
0(
#244560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#244610000000
0$
0)
#244620000000
1"
1'
b0 +
b0 1
#244670000000
0"
0'
#244680000000
1#
1(
b101111101100100 +
b101111101100100 1
#244730000000
0#
0(
#244740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#244790000000
0$
0)
#244800000000
1"
1'
b0 +
b0 1
#244850000000
0"
0'
#244860000000
1#
1(
b101111101100100 +
b101111101100100 1
#244910000000
0#
0(
#244920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#244970000000
0$
0)
#244980000000
1"
1'
b0 +
b0 1
#245030000000
0"
0'
#245040000000
1#
1(
b101111101100100 +
b101111101100100 1
#245090000000
0#
0(
#245100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#245150000000
0$
0)
#245160000000
1"
1'
b0 +
b0 1
#245210000000
0"
0'
#245220000000
1#
1(
b101111101100100 +
b101111101100100 1
#245270000000
0#
0(
#245280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#245330000000
0$
0)
#245340000000
1"
1'
b0 +
b0 1
#245390000000
0"
0'
#245400000000
1#
1(
b101111101100100 +
b101111101100100 1
#245450000000
0#
0(
#245460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#245510000000
0$
0)
#245520000000
1"
1'
b0 +
b0 1
#245570000000
0"
0'
#245580000000
1#
1(
b101111101100100 +
b101111101100100 1
#245630000000
0#
0(
#245640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#245690000000
0$
0)
#245700000000
1"
1'
b0 +
b0 1
#245750000000
0"
0'
#245760000000
1#
1(
b101111101100100 +
b101111101100100 1
#245810000000
0#
0(
#245820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#245870000000
0$
0)
#245880000000
1"
1'
b0 +
b0 1
#245930000000
0"
0'
#245940000000
1#
1(
b101111101100100 +
b101111101100100 1
#245990000000
0#
0(
#246000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#246050000000
0$
0)
#246060000000
1"
1'
b0 +
b0 1
#246110000000
0"
0'
#246120000000
1#
1(
b101111101100100 +
b101111101100100 1
#246170000000
0#
0(
#246180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#246230000000
0$
0)
#246240000000
1"
1'
b0 +
b0 1
#246290000000
0"
0'
#246300000000
1#
1(
b101111101100100 +
b101111101100100 1
#246350000000
0#
0(
#246360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#246410000000
0$
0)
#246420000000
1"
1'
b0 +
b0 1
#246470000000
0"
0'
#246480000000
1#
1(
b101111101100100 +
b101111101100100 1
#246530000000
0#
0(
#246540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#246590000000
0$
0)
#246600000000
1"
1'
b0 +
b0 1
#246650000000
0"
0'
#246660000000
1#
1(
b101111101100100 +
b101111101100100 1
#246710000000
0#
0(
#246720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#246770000000
0$
0)
#246780000000
1"
1'
b0 +
b0 1
#246830000000
0"
0'
#246840000000
1#
1(
b101111101100100 +
b101111101100100 1
#246890000000
0#
0(
#246900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#246950000000
0$
0)
#246960000000
1"
1'
b0 +
b0 1
#247010000000
0"
0'
#247020000000
1#
1(
b101111101100100 +
b101111101100100 1
#247070000000
0#
0(
#247080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#247130000000
0$
0)
#247140000000
1"
1'
b0 +
b0 1
#247190000000
0"
0'
#247200000000
1#
1(
b101111101100100 +
b101111101100100 1
#247250000000
0#
0(
#247260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#247310000000
0$
0)
#247320000000
1"
1'
b0 +
b0 1
#247370000000
0"
0'
#247380000000
1#
1(
b101111101100100 +
b101111101100100 1
#247430000000
0#
0(
#247440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#247490000000
0$
0)
#247500000000
1"
1'
b0 +
b0 1
#247550000000
0"
0'
#247560000000
1#
1(
b101111101100100 +
b101111101100100 1
#247610000000
0#
0(
#247620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#247670000000
0$
0)
#247680000000
1"
1'
b0 +
b0 1
#247730000000
0"
0'
#247740000000
1#
1(
b101111101100100 +
b101111101100100 1
#247790000000
0#
0(
#247800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#247850000000
0$
0)
#247860000000
1"
1'
b0 +
b0 1
#247910000000
0"
0'
#247920000000
1#
1(
b101111101100100 +
b101111101100100 1
#247970000000
0#
0(
#247980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#248030000000
0$
0)
#248040000000
1"
1'
b0 +
b0 1
#248090000000
0"
0'
#248100000000
1#
1(
b101111101100100 +
b101111101100100 1
#248150000000
0#
0(
#248160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#248210000000
0$
0)
#248220000000
1"
1'
b0 +
b0 1
#248270000000
0"
0'
#248280000000
1#
1(
b101111101100100 +
b101111101100100 1
#248330000000
0#
0(
#248340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#248390000000
0$
0)
#248400000000
1"
1'
b0 +
b0 1
#248450000000
0"
0'
#248460000000
1#
1(
b101111101100100 +
b101111101100100 1
#248510000000
0#
0(
#248520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#248570000000
0$
0)
#248580000000
1"
1'
b0 +
b0 1
#248630000000
0"
0'
#248640000000
1#
1(
b101111101100100 +
b101111101100100 1
#248690000000
0#
0(
#248700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#248750000000
0$
0)
#248760000000
1"
1'
b0 +
b0 1
#248810000000
0"
0'
#248820000000
1#
1(
b101111101100100 +
b101111101100100 1
#248870000000
0#
0(
#248880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#248930000000
0$
0)
#248940000000
1"
1'
b0 +
b0 1
#248990000000
0"
0'
#249000000000
1#
1(
b101111101100100 +
b101111101100100 1
#249050000000
0#
0(
#249060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#249110000000
0$
0)
#249120000000
1"
1'
b0 +
b0 1
#249170000000
0"
0'
#249180000000
1#
1(
b101111101100100 +
b101111101100100 1
#249230000000
0#
0(
#249240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#249290000000
0$
0)
#249300000000
1"
1'
b0 +
b0 1
#249350000000
0"
0'
#249360000000
1#
1(
b101111101100100 +
b101111101100100 1
#249410000000
0#
0(
#249420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#249470000000
0$
0)
#249480000000
1"
1'
b0 +
b0 1
#249530000000
0"
0'
#249540000000
1#
1(
b101111101100100 +
b101111101100100 1
#249590000000
0#
0(
#249600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#249650000000
0$
0)
#249660000000
1"
1'
b0 +
b0 1
#249710000000
0"
0'
#249720000000
1#
1(
b101111101100100 +
b101111101100100 1
#249770000000
0#
0(
#249780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#249830000000
0$
0)
#249840000000
1"
1'
b0 +
b0 1
#249890000000
0"
0'
#249900000000
1#
1(
b101111101100100 +
b101111101100100 1
#249950000000
0#
0(
#249960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#250010000000
0$
0)
#250020000000
1"
1'
b0 +
b0 1
#250070000000
0"
0'
#250080000000
1#
1(
b101111101100100 +
b101111101100100 1
#250130000000
0#
0(
#250140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#250190000000
0$
0)
#250200000000
1"
1'
b0 +
b0 1
#250250000000
0"
0'
#250260000000
1#
1(
b101111101100100 +
b101111101100100 1
#250310000000
0#
0(
#250320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#250370000000
0$
0)
#250380000000
1"
1'
b0 +
b0 1
#250430000000
0"
0'
#250440000000
1#
1(
b101111101100100 +
b101111101100100 1
#250490000000
0#
0(
#250500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#250550000000
0$
0)
#250560000000
1"
1'
b0 +
b0 1
#250610000000
0"
0'
#250620000000
1#
1(
b101111101100100 +
b101111101100100 1
#250670000000
0#
0(
#250680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#250730000000
0$
0)
#250740000000
1"
1'
b0 +
b0 1
#250790000000
0"
0'
#250800000000
1#
1(
b101111101100100 +
b101111101100100 1
#250850000000
0#
0(
#250860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#250910000000
0$
0)
#250920000000
1"
1'
b0 +
b0 1
#250970000000
0"
0'
#250980000000
1#
1(
b101111101100100 +
b101111101100100 1
#251030000000
0#
0(
#251040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#251090000000
0$
0)
#251100000000
1"
1'
b0 +
b0 1
#251150000000
0"
0'
#251160000000
1#
1(
b101111101100100 +
b101111101100100 1
#251210000000
0#
0(
#251220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#251270000000
0$
0)
#251280000000
1"
1'
b0 +
b0 1
#251330000000
0"
0'
#251340000000
1#
1(
b101111101100100 +
b101111101100100 1
#251390000000
0#
0(
#251400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#251450000000
0$
0)
#251460000000
1"
1'
b0 +
b0 1
#251510000000
0"
0'
#251520000000
1#
1(
b101111101100100 +
b101111101100100 1
#251570000000
0#
0(
#251580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#251630000000
0$
0)
#251640000000
1"
1'
b0 +
b0 1
#251690000000
0"
0'
#251700000000
1#
1(
b101111101100100 +
b101111101100100 1
#251750000000
0#
0(
#251760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#251810000000
0$
0)
#251820000000
1"
1'
b0 +
b0 1
#251870000000
0"
0'
#251880000000
1#
1(
b101111101100100 +
b101111101100100 1
#251930000000
0#
0(
#251940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#251990000000
0$
0)
#252000000000
1"
1'
b0 +
b0 1
#252050000000
0"
0'
#252060000000
1#
1(
b101111101100100 +
b101111101100100 1
#252110000000
0#
0(
#252120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#252170000000
0$
0)
#252180000000
1"
1'
b0 +
b0 1
#252230000000
0"
0'
#252240000000
1#
1(
b101111101100100 +
b101111101100100 1
#252290000000
0#
0(
#252300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#252350000000
0$
0)
#252360000000
1"
1'
b0 +
b0 1
#252410000000
0"
0'
#252420000000
1#
1(
b101111101100100 +
b101111101100100 1
#252470000000
0#
0(
#252480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#252530000000
0$
0)
#252540000000
1"
1'
b0 +
b0 1
#252590000000
0"
0'
#252600000000
1#
1(
b101111101100100 +
b101111101100100 1
#252650000000
0#
0(
#252660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#252710000000
0$
0)
#252720000000
1"
1'
b0 +
b0 1
#252770000000
0"
0'
#252780000000
1#
1(
b101111101100100 +
b101111101100100 1
#252830000000
0#
0(
#252840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#252890000000
0$
0)
#252900000000
1"
1'
b0 +
b0 1
#252950000000
0"
0'
#252960000000
1#
1(
b101111101100100 +
b101111101100100 1
#253010000000
0#
0(
#253020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#253070000000
0$
0)
#253080000000
1"
1'
b0 +
b0 1
#253130000000
0"
0'
#253140000000
1#
1(
b101111101100100 +
b101111101100100 1
#253190000000
0#
0(
#253200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#253250000000
0$
0)
#253260000000
1"
1'
b0 +
b0 1
#253310000000
0"
0'
#253320000000
1#
1(
b101111101100100 +
b101111101100100 1
#253370000000
0#
0(
#253380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#253430000000
0$
0)
#253440000000
1"
1'
b0 +
b0 1
#253490000000
0"
0'
#253500000000
1#
1(
b101111101100100 +
b101111101100100 1
#253550000000
0#
0(
#253560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#253610000000
0$
0)
#253620000000
1"
1'
b0 +
b0 1
#253670000000
0"
0'
#253680000000
1#
1(
b101111101100100 +
b101111101100100 1
#253730000000
0#
0(
#253740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#253790000000
0$
0)
#253800000000
1"
1'
b0 +
b0 1
#253850000000
0"
0'
#253860000000
1#
1(
b101111101100100 +
b101111101100100 1
#253910000000
0#
0(
#253920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#253970000000
0$
0)
#253980000000
1"
1'
b0 +
b0 1
#254030000000
0"
0'
#254040000000
1#
1(
b101111101100100 +
b101111101100100 1
#254090000000
0#
0(
#254100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#254150000000
0$
0)
#254160000000
1"
1'
b0 +
b0 1
#254210000000
0"
0'
#254220000000
1#
1(
b101111101100100 +
b101111101100100 1
#254270000000
0#
0(
#254280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#254330000000
0$
0)
#254340000000
1"
1'
b0 +
b0 1
#254390000000
0"
0'
#254400000000
1#
1(
b101111101100100 +
b101111101100100 1
#254450000000
0#
0(
#254460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#254510000000
0$
0)
#254520000000
1"
1'
b0 +
b0 1
#254570000000
0"
0'
#254580000000
1#
1(
b101111101100100 +
b101111101100100 1
#254630000000
0#
0(
#254640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#254690000000
0$
0)
#254700000000
1"
1'
b0 +
b0 1
#254750000000
0"
0'
#254760000000
1#
1(
b101111101100100 +
b101111101100100 1
#254810000000
0#
0(
#254820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#254870000000
0$
0)
#254880000000
1"
1'
b0 +
b0 1
#254930000000
0"
0'
#254940000000
1#
1(
b101111101100100 +
b101111101100100 1
#254990000000
0#
0(
#255000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#255050000000
0$
0)
#255060000000
1"
1'
b0 +
b0 1
#255110000000
0"
0'
#255120000000
1#
1(
b101111101100100 +
b101111101100100 1
#255170000000
0#
0(
#255180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#255230000000
0$
0)
#255240000000
1"
1'
b0 +
b0 1
#255290000000
0"
0'
#255300000000
1#
1(
b101111101100100 +
b101111101100100 1
#255350000000
0#
0(
#255360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#255410000000
0$
0)
#255420000000
1"
1'
b0 +
b0 1
#255470000000
0"
0'
#255480000000
1#
1(
b101111101100100 +
b101111101100100 1
#255530000000
0#
0(
#255540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#255590000000
0$
0)
#255600000000
1"
1'
b0 +
b0 1
#255650000000
0"
0'
#255660000000
1#
1(
b101111101100100 +
b101111101100100 1
#255710000000
0#
0(
#255720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#255770000000
0$
0)
#255780000000
1"
1'
b0 +
b0 1
#255830000000
0"
0'
#255840000000
1#
1(
b101111101100100 +
b101111101100100 1
#255890000000
0#
0(
#255900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#255950000000
0$
0)
#255960000000
1"
1'
b0 +
b0 1
#256010000000
0"
0'
#256020000000
1#
1(
b101111101100100 +
b101111101100100 1
#256070000000
0#
0(
#256080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#256130000000
0$
0)
#256140000000
1"
1'
b0 +
b0 1
#256190000000
0"
0'
#256200000000
1#
1(
b101111101100100 +
b101111101100100 1
#256250000000
0#
0(
#256260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#256310000000
0$
0)
#256320000000
1"
1'
b0 +
b0 1
#256370000000
0"
0'
#256380000000
1#
1(
b101111101100100 +
b101111101100100 1
#256430000000
0#
0(
#256440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#256490000000
0$
0)
#256500000000
1"
1'
b0 +
b0 1
#256550000000
0"
0'
#256560000000
1#
1(
b101111101100100 +
b101111101100100 1
#256610000000
0#
0(
#256620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#256670000000
0$
0)
#256680000000
1"
1'
b0 +
b0 1
#256730000000
0"
0'
#256740000000
1#
1(
b101111101100100 +
b101111101100100 1
#256790000000
0#
0(
#256800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#256850000000
0$
0)
#256860000000
1"
1'
b0 +
b0 1
#256910000000
0"
0'
#256920000000
1#
1(
b101111101100100 +
b101111101100100 1
#256970000000
0#
0(
#256980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#257030000000
0$
0)
#257040000000
1"
1'
b0 +
b0 1
#257090000000
0"
0'
#257100000000
1#
1(
b101111101100100 +
b101111101100100 1
#257150000000
0#
0(
#257160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#257210000000
0$
0)
#257220000000
1"
1'
b0 +
b0 1
#257270000000
0"
0'
#257280000000
1#
1(
b101111101100100 +
b101111101100100 1
#257330000000
0#
0(
#257340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#257390000000
0$
0)
#257400000000
1"
1'
b0 +
b0 1
#257450000000
0"
0'
#257460000000
1#
1(
b101111101100100 +
b101111101100100 1
#257510000000
0#
0(
#257520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#257570000000
0$
0)
#257580000000
1"
1'
b0 +
b0 1
#257630000000
0"
0'
#257640000000
1#
1(
b101111101100100 +
b101111101100100 1
#257690000000
0#
0(
#257700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#257750000000
0$
0)
#257760000000
1"
1'
b0 +
b0 1
#257810000000
0"
0'
#257820000000
1#
1(
b101111101100100 +
b101111101100100 1
#257870000000
0#
0(
#257880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#257930000000
0$
0)
#257940000000
1"
1'
b0 +
b0 1
#257990000000
0"
0'
#258000000000
1#
1(
b101111101100100 +
b101111101100100 1
#258050000000
0#
0(
#258060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#258110000000
0$
0)
#258120000000
1"
1'
b0 +
b0 1
#258170000000
0"
0'
#258180000000
1#
1(
b101111101100100 +
b101111101100100 1
#258230000000
0#
0(
#258240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#258290000000
0$
0)
#258300000000
1"
1'
b0 +
b0 1
#258350000000
0"
0'
#258360000000
1#
1(
b101111101100100 +
b101111101100100 1
#258410000000
0#
0(
#258420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#258470000000
0$
0)
#258480000000
1"
1'
b0 +
b0 1
#258530000000
0"
0'
#258540000000
1#
1(
b101111101100100 +
b101111101100100 1
#258590000000
0#
0(
#258600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#258650000000
0$
0)
#258660000000
1"
1'
b0 +
b0 1
#258710000000
0"
0'
#258720000000
1#
1(
b101111101100100 +
b101111101100100 1
#258770000000
0#
0(
#258780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#258830000000
0$
0)
#258840000000
1"
1'
b0 +
b0 1
#258890000000
0"
0'
#258900000000
1#
1(
b101111101100100 +
b101111101100100 1
#258950000000
0#
0(
#258960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#259010000000
0$
0)
#259020000000
1"
1'
b0 +
b0 1
#259070000000
0"
0'
#259080000000
1#
1(
b101111101100100 +
b101111101100100 1
#259130000000
0#
0(
#259140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#259190000000
0$
0)
#259200000000
1"
1'
b0 +
b0 1
#259250000000
0"
0'
#259260000000
1#
1(
b101111101100100 +
b101111101100100 1
#259310000000
0#
0(
#259320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#259370000000
0$
0)
#259380000000
1"
1'
b0 +
b0 1
#259430000000
0"
0'
#259440000000
1#
1(
b101111101100100 +
b101111101100100 1
#259490000000
0#
0(
#259500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#259550000000
0$
0)
#259560000000
1"
1'
b0 +
b0 1
#259610000000
0"
0'
#259620000000
1#
1(
b101111101100100 +
b101111101100100 1
#259670000000
0#
0(
#259680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#259730000000
0$
0)
#259740000000
1"
1'
b0 +
b0 1
#259790000000
0"
0'
#259800000000
1#
1(
b101111101100100 +
b101111101100100 1
#259850000000
0#
0(
#259860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#259910000000
0$
0)
#259920000000
1"
1'
b0 +
b0 1
#259970000000
0"
0'
#259980000000
1#
1(
b101111101100100 +
b101111101100100 1
#260030000000
0#
0(
#260040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#260090000000
0$
0)
#260100000000
1"
1'
b0 +
b0 1
#260150000000
0"
0'
#260160000000
1#
1(
b101111101100100 +
b101111101100100 1
#260210000000
0#
0(
#260220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#260270000000
0$
0)
#260280000000
1"
1'
b0 +
b0 1
#260330000000
0"
0'
#260340000000
1#
1(
b101111101100100 +
b101111101100100 1
#260390000000
0#
0(
#260400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#260450000000
0$
0)
#260460000000
1"
1'
b0 +
b0 1
#260510000000
0"
0'
#260520000000
1#
1(
b101111101100100 +
b101111101100100 1
#260570000000
0#
0(
#260580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#260630000000
0$
0)
#260640000000
1"
1'
b0 +
b0 1
#260690000000
0"
0'
#260700000000
1#
1(
b101111101100100 +
b101111101100100 1
#260750000000
0#
0(
#260760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#260810000000
0$
0)
#260820000000
1"
1'
b0 +
b0 1
#260870000000
0"
0'
#260880000000
1#
1(
b101111101100100 +
b101111101100100 1
#260930000000
0#
0(
#260940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#260990000000
0$
0)
#261000000000
1"
1'
b0 +
b0 1
#261050000000
0"
0'
#261060000000
1#
1(
b101111101100100 +
b101111101100100 1
#261110000000
0#
0(
#261120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#261170000000
0$
0)
#261180000000
1"
1'
b0 +
b0 1
#261230000000
0"
0'
#261240000000
1#
1(
b101111101100100 +
b101111101100100 1
#261290000000
0#
0(
#261300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#261350000000
0$
0)
#261360000000
1"
1'
b0 +
b0 1
#261410000000
0"
0'
#261420000000
1#
1(
b101111101100100 +
b101111101100100 1
#261470000000
0#
0(
#261480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#261530000000
0$
0)
#261540000000
1"
1'
b0 +
b0 1
#261590000000
0"
0'
#261600000000
1#
1(
b101111101100100 +
b101111101100100 1
#261650000000
0#
0(
#261660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#261710000000
0$
0)
#261720000000
1"
1'
b0 +
b0 1
#261770000000
0"
0'
#261780000000
1#
1(
b101111101100100 +
b101111101100100 1
#261830000000
0#
0(
#261840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#261890000000
0$
0)
#261900000000
1"
1'
b0 +
b0 1
#261950000000
0"
0'
#261960000000
1#
1(
b101111101100100 +
b101111101100100 1
#262010000000
0#
0(
#262020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#262070000000
0$
0)
#262080000000
1"
1'
b0 +
b0 1
#262130000000
0"
0'
#262140000000
1#
1(
b101111101100100 +
b101111101100100 1
#262190000000
0#
0(
#262200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#262250000000
0$
0)
#262260000000
1"
1'
b0 +
b0 1
#262310000000
0"
0'
#262320000000
1#
1(
b101111101100100 +
b101111101100100 1
#262370000000
0#
0(
#262380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#262430000000
0$
0)
#262440000000
1"
1'
b0 +
b0 1
#262490000000
0"
0'
#262500000000
1#
1(
b101111101100100 +
b101111101100100 1
#262550000000
0#
0(
#262560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#262610000000
0$
0)
#262620000000
1"
1'
b0 +
b0 1
#262670000000
0"
0'
#262680000000
1#
1(
b101111101100100 +
b101111101100100 1
#262730000000
0#
0(
#262740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#262790000000
0$
0)
#262800000000
1"
1'
b0 +
b0 1
#262850000000
0"
0'
#262860000000
1#
1(
b101111101100100 +
b101111101100100 1
#262910000000
0#
0(
#262920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#262970000000
0$
0)
#262980000000
1"
1'
b0 +
b0 1
#263030000000
0"
0'
#263040000000
1#
1(
b101111101100100 +
b101111101100100 1
#263090000000
0#
0(
#263100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#263150000000
0$
0)
#263160000000
1"
1'
b0 +
b0 1
#263210000000
0"
0'
#263220000000
1#
1(
b101111101100100 +
b101111101100100 1
#263270000000
0#
0(
#263280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#263330000000
0$
0)
#263340000000
1"
1'
b0 +
b0 1
#263390000000
0"
0'
#263400000000
1#
1(
b101111101100100 +
b101111101100100 1
#263450000000
0#
0(
#263460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#263510000000
0$
0)
#263520000000
1"
1'
b0 +
b0 1
#263570000000
0"
0'
#263580000000
1#
1(
b101111101100100 +
b101111101100100 1
#263630000000
0#
0(
#263640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#263690000000
0$
0)
#263700000000
1"
1'
b0 +
b0 1
#263750000000
0"
0'
#263760000000
1#
1(
b101111101100100 +
b101111101100100 1
#263810000000
0#
0(
#263820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#263870000000
0$
0)
#263880000000
1"
1'
b0 +
b0 1
#263930000000
0"
0'
#263940000000
1#
1(
b101111101100100 +
b101111101100100 1
#263990000000
0#
0(
#264000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#264050000000
0$
0)
#264060000000
1"
1'
b0 +
b0 1
#264110000000
0"
0'
#264120000000
1#
1(
b101111101100100 +
b101111101100100 1
#264170000000
0#
0(
#264180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#264230000000
0$
0)
#264240000000
1"
1'
b0 +
b0 1
#264290000000
0"
0'
#264300000000
1#
1(
b101111101100100 +
b101111101100100 1
#264350000000
0#
0(
#264360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#264410000000
0$
0)
#264420000000
1"
1'
b0 +
b0 1
#264470000000
0"
0'
#264480000000
1#
1(
b101111101100100 +
b101111101100100 1
#264530000000
0#
0(
#264540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#264590000000
0$
0)
#264600000000
1"
1'
b0 +
b0 1
#264650000000
0"
0'
#264660000000
1#
1(
b101111101100100 +
b101111101100100 1
#264710000000
0#
0(
#264720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#264770000000
0$
0)
#264780000000
1"
1'
b0 +
b0 1
#264830000000
0"
0'
#264840000000
1#
1(
b101111101100100 +
b101111101100100 1
#264890000000
0#
0(
#264900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#264950000000
0$
0)
#264960000000
1"
1'
b0 +
b0 1
#265010000000
0"
0'
#265020000000
1#
1(
b101111101100100 +
b101111101100100 1
#265070000000
0#
0(
#265080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#265130000000
0$
0)
#265140000000
1"
1'
b0 +
b0 1
#265190000000
0"
0'
#265200000000
1#
1(
b101111101100100 +
b101111101100100 1
#265250000000
0#
0(
#265260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#265310000000
0$
0)
#265320000000
1"
1'
b0 +
b0 1
#265370000000
0"
0'
#265380000000
1#
1(
b101111101100100 +
b101111101100100 1
#265430000000
0#
0(
#265440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#265490000000
0$
0)
#265500000000
1"
1'
b0 +
b0 1
#265550000000
0"
0'
#265560000000
1#
1(
b101111101100100 +
b101111101100100 1
#265610000000
0#
0(
#265620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#265670000000
0$
0)
#265680000000
1"
1'
b0 +
b0 1
#265730000000
0"
0'
#265740000000
1#
1(
b101111101100100 +
b101111101100100 1
#265790000000
0#
0(
#265800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#265850000000
0$
0)
#265860000000
1"
1'
b0 +
b0 1
#265910000000
0"
0'
#265920000000
1#
1(
b101111101100100 +
b101111101100100 1
#265970000000
0#
0(
#265980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#266030000000
0$
0)
#266040000000
1"
1'
b0 +
b0 1
#266090000000
0"
0'
#266100000000
1#
1(
b101111101100100 +
b101111101100100 1
#266150000000
0#
0(
#266160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#266210000000
0$
0)
#266220000000
1"
1'
b0 +
b0 1
#266270000000
0"
0'
#266280000000
1#
1(
b101111101100100 +
b101111101100100 1
#266330000000
0#
0(
#266340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#266390000000
0$
0)
#266400000000
1"
1'
b0 +
b0 1
#266450000000
0"
0'
#266460000000
1#
1(
b101111101100100 +
b101111101100100 1
#266510000000
0#
0(
#266520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#266570000000
0$
0)
#266580000000
1"
1'
b0 +
b0 1
#266630000000
0"
0'
#266640000000
1#
1(
b101111101100100 +
b101111101100100 1
#266690000000
0#
0(
#266700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#266750000000
0$
0)
#266760000000
1"
1'
b0 +
b0 1
#266810000000
0"
0'
#266820000000
1#
1(
b101111101100100 +
b101111101100100 1
#266870000000
0#
0(
#266880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#266930000000
0$
0)
#266940000000
1"
1'
b0 +
b0 1
#266990000000
0"
0'
#267000000000
1#
1(
b101111101100100 +
b101111101100100 1
#267050000000
0#
0(
#267060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#267110000000
0$
0)
#267120000000
1"
1'
b0 +
b0 1
#267170000000
0"
0'
#267180000000
1#
1(
b101111101100100 +
b101111101100100 1
#267230000000
0#
0(
#267240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#267290000000
0$
0)
#267300000000
1"
1'
b0 +
b0 1
#267350000000
0"
0'
#267360000000
1#
1(
b101111101100100 +
b101111101100100 1
#267410000000
0#
0(
#267420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#267470000000
0$
0)
#267480000000
1"
1'
b0 +
b0 1
#267530000000
0"
0'
#267540000000
1#
1(
b101111101100100 +
b101111101100100 1
#267590000000
0#
0(
#267600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#267650000000
0$
0)
#267660000000
1"
1'
b0 +
b0 1
#267710000000
0"
0'
#267720000000
1#
1(
b101111101100100 +
b101111101100100 1
#267770000000
0#
0(
#267780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#267830000000
0$
0)
#267840000000
1"
1'
b0 +
b0 1
#267890000000
0"
0'
#267900000000
1#
1(
b101111101100100 +
b101111101100100 1
#267950000000
0#
0(
#267960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#268010000000
0$
0)
#268020000000
1"
1'
b0 +
b0 1
#268070000000
0"
0'
#268080000000
1#
1(
b101111101100100 +
b101111101100100 1
#268130000000
0#
0(
#268140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#268190000000
0$
0)
#268200000000
1"
1'
b0 +
b0 1
#268250000000
0"
0'
#268260000000
1#
1(
b101111101100100 +
b101111101100100 1
#268310000000
0#
0(
#268320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#268370000000
0$
0)
#268380000000
1"
1'
b0 +
b0 1
#268430000000
0"
0'
#268440000000
1#
1(
b101111101100100 +
b101111101100100 1
#268490000000
0#
0(
#268500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#268550000000
0$
0)
#268560000000
1"
1'
b0 +
b0 1
#268610000000
0"
0'
#268620000000
1#
1(
b101111101100100 +
b101111101100100 1
#268670000000
0#
0(
#268680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#268730000000
0$
0)
#268740000000
1"
1'
b0 +
b0 1
#268790000000
0"
0'
#268800000000
1#
1(
b101111101100100 +
b101111101100100 1
#268850000000
0#
0(
#268860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#268910000000
0$
0)
#268920000000
1"
1'
b0 +
b0 1
#268970000000
0"
0'
#268980000000
1#
1(
b101111101100100 +
b101111101100100 1
#269030000000
0#
0(
#269040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#269090000000
0$
0)
#269100000000
1"
1'
b0 +
b0 1
#269150000000
0"
0'
#269160000000
1#
1(
b101111101100100 +
b101111101100100 1
#269210000000
0#
0(
#269220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#269270000000
0$
0)
#269280000000
1"
1'
b0 +
b0 1
#269330000000
0"
0'
#269340000000
1#
1(
b101111101100100 +
b101111101100100 1
#269390000000
0#
0(
#269400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#269450000000
0$
0)
#269460000000
1"
1'
b0 +
b0 1
#269510000000
0"
0'
#269520000000
1#
1(
b101111101100100 +
b101111101100100 1
#269570000000
0#
0(
#269580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#269630000000
0$
0)
#269640000000
1"
1'
b0 +
b0 1
#269690000000
0"
0'
#269700000000
1#
1(
b101111101100100 +
b101111101100100 1
#269750000000
0#
0(
#269760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#269810000000
0$
0)
#269820000000
1"
1'
b0 +
b0 1
#269870000000
0"
0'
#269880000000
1#
1(
b101111101100100 +
b101111101100100 1
#269930000000
0#
0(
#269940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#269990000000
0$
0)
#270000000000
1"
1'
b0 +
b0 1
#270050000000
0"
0'
#270060000000
1#
1(
b101111101100100 +
b101111101100100 1
#270110000000
0#
0(
#270120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#270170000000
0$
0)
#270180000000
1"
1'
b0 +
b0 1
#270230000000
0"
0'
#270240000000
1#
1(
b101111101100100 +
b101111101100100 1
#270290000000
0#
0(
#270300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#270350000000
0$
0)
#270360000000
1"
1'
b0 +
b0 1
#270410000000
0"
0'
#270420000000
1#
1(
b101111101100100 +
b101111101100100 1
#270470000000
0#
0(
#270480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#270530000000
0$
0)
#270540000000
1"
1'
b0 +
b0 1
#270590000000
0"
0'
#270600000000
1#
1(
b101111101100100 +
b101111101100100 1
#270650000000
0#
0(
#270660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#270710000000
0$
0)
#270720000000
1"
1'
b0 +
b0 1
#270770000000
0"
0'
#270780000000
1#
1(
b101111101100100 +
b101111101100100 1
#270830000000
0#
0(
#270840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#270890000000
0$
0)
#270900000000
1"
1'
b0 +
b0 1
#270950000000
0"
0'
#270960000000
1#
1(
b101111101100100 +
b101111101100100 1
#271010000000
0#
0(
#271020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#271070000000
0$
0)
#271080000000
1"
1'
b0 +
b0 1
#271130000000
0"
0'
#271140000000
1#
1(
b101111101100100 +
b101111101100100 1
#271190000000
0#
0(
#271200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#271250000000
0$
0)
#271260000000
1"
1'
b0 +
b0 1
#271310000000
0"
0'
#271320000000
1#
1(
b101111101100100 +
b101111101100100 1
#271370000000
0#
0(
#271380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#271430000000
0$
0)
#271440000000
1"
1'
b0 +
b0 1
#271490000000
0"
0'
#271500000000
1#
1(
b101111101100100 +
b101111101100100 1
#271550000000
0#
0(
#271560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#271610000000
0$
0)
#271620000000
1"
1'
b0 +
b0 1
#271670000000
0"
0'
#271680000000
1#
1(
b101111101100100 +
b101111101100100 1
#271730000000
0#
0(
#271740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#271790000000
0$
0)
#271800000000
1"
1'
b0 +
b0 1
#271850000000
0"
0'
#271860000000
1#
1(
b101111101100100 +
b101111101100100 1
#271910000000
0#
0(
#271920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#271970000000
0$
0)
#271980000000
1"
1'
b0 +
b0 1
#272030000000
0"
0'
#272040000000
1#
1(
b101111101100100 +
b101111101100100 1
#272090000000
0#
0(
#272100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#272150000000
0$
0)
#272160000000
1"
1'
b0 +
b0 1
#272210000000
0"
0'
#272220000000
1#
1(
b101111101100100 +
b101111101100100 1
#272270000000
0#
0(
#272280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#272330000000
0$
0)
#272340000000
1"
1'
b0 +
b0 1
#272390000000
0"
0'
#272400000000
1#
1(
b101111101100100 +
b101111101100100 1
#272450000000
0#
0(
#272460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#272510000000
0$
0)
#272520000000
1"
1'
b0 +
b0 1
#272570000000
0"
0'
#272580000000
1#
1(
b101111101100100 +
b101111101100100 1
#272630000000
0#
0(
#272640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#272690000000
0$
0)
#272700000000
1"
1'
b0 +
b0 1
#272750000000
0"
0'
#272760000000
1#
1(
b101111101100100 +
b101111101100100 1
#272810000000
0#
0(
#272820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#272870000000
0$
0)
#272880000000
1"
1'
b0 +
b0 1
#272930000000
0"
0'
#272940000000
1#
1(
b101111101100100 +
b101111101100100 1
#272990000000
0#
0(
#273000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#273050000000
0$
0)
#273060000000
1"
1'
b0 +
b0 1
#273110000000
0"
0'
#273120000000
1#
1(
b101111101100100 +
b101111101100100 1
#273170000000
0#
0(
#273180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#273230000000
0$
0)
#273240000000
1"
1'
b0 +
b0 1
#273290000000
0"
0'
#273300000000
1#
1(
b101111101100100 +
b101111101100100 1
#273350000000
0#
0(
#273360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#273410000000
0$
0)
#273420000000
1"
1'
b0 +
b0 1
#273470000000
0"
0'
#273480000000
1#
1(
b101111101100100 +
b101111101100100 1
#273530000000
0#
0(
#273540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#273590000000
0$
0)
#273600000000
1"
1'
b0 +
b0 1
#273650000000
0"
0'
#273660000000
1#
1(
b101111101100100 +
b101111101100100 1
#273710000000
0#
0(
#273720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#273770000000
0$
0)
#273780000000
1"
1'
b0 +
b0 1
#273830000000
0"
0'
#273840000000
1#
1(
b101111101100100 +
b101111101100100 1
#273890000000
0#
0(
#273900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#273950000000
0$
0)
#273960000000
1"
1'
b0 +
b0 1
#274010000000
0"
0'
#274020000000
1#
1(
b101111101100100 +
b101111101100100 1
#274070000000
0#
0(
#274080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#274130000000
0$
0)
#274140000000
1"
1'
b0 +
b0 1
#274190000000
0"
0'
#274200000000
1#
1(
b101111101100100 +
b101111101100100 1
#274250000000
0#
0(
#274260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#274310000000
0$
0)
#274320000000
1"
1'
b0 +
b0 1
#274370000000
0"
0'
#274380000000
1#
1(
b101111101100100 +
b101111101100100 1
#274430000000
0#
0(
#274440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#274490000000
0$
0)
#274500000000
1"
1'
b0 +
b0 1
#274550000000
0"
0'
#274560000000
1#
1(
b101111101100100 +
b101111101100100 1
#274610000000
0#
0(
#274620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#274670000000
0$
0)
#274680000000
1"
1'
b0 +
b0 1
#274730000000
0"
0'
#274740000000
1#
1(
b101111101100100 +
b101111101100100 1
#274790000000
0#
0(
#274800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#274850000000
0$
0)
#274860000000
1"
1'
b0 +
b0 1
#274910000000
0"
0'
#274920000000
1#
1(
b101111101100100 +
b101111101100100 1
#274970000000
0#
0(
#274980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#275030000000
0$
0)
#275040000000
1"
1'
b0 +
b0 1
#275090000000
0"
0'
#275100000000
1#
1(
b101111101100100 +
b101111101100100 1
#275150000000
0#
0(
#275160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#275210000000
0$
0)
#275220000000
1"
1'
b0 +
b0 1
#275270000000
0"
0'
#275280000000
1#
1(
b101111101100100 +
b101111101100100 1
#275330000000
0#
0(
#275340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#275390000000
0$
0)
#275400000000
1"
1'
b0 +
b0 1
#275450000000
0"
0'
#275460000000
1#
1(
b101111101100100 +
b101111101100100 1
#275510000000
0#
0(
#275520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#275570000000
0$
0)
#275580000000
1"
1'
b0 +
b0 1
#275630000000
0"
0'
#275640000000
1#
1(
b101111101100100 +
b101111101100100 1
#275690000000
0#
0(
#275700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#275750000000
0$
0)
#275760000000
1"
1'
b0 +
b0 1
#275810000000
0"
0'
#275820000000
1#
1(
b101111101100100 +
b101111101100100 1
#275870000000
0#
0(
#275880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#275930000000
0$
0)
#275940000000
1"
1'
b0 +
b0 1
#275990000000
0"
0'
#276000000000
1#
1(
b101111101100100 +
b101111101100100 1
#276050000000
0#
0(
#276060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#276110000000
0$
0)
#276120000000
1"
1'
b0 +
b0 1
#276170000000
0"
0'
#276180000000
1#
1(
b101111101100100 +
b101111101100100 1
#276230000000
0#
0(
#276240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#276290000000
0$
0)
#276300000000
1"
1'
b0 +
b0 1
#276350000000
0"
0'
#276360000000
1#
1(
b101111101100100 +
b101111101100100 1
#276410000000
0#
0(
#276420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#276470000000
0$
0)
#276480000000
1"
1'
b0 +
b0 1
#276530000000
0"
0'
#276540000000
1#
1(
b101111101100100 +
b101111101100100 1
#276590000000
0#
0(
#276600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#276650000000
0$
0)
#276660000000
1"
1'
b0 +
b0 1
#276710000000
0"
0'
#276720000000
1#
1(
b101111101100100 +
b101111101100100 1
#276770000000
0#
0(
#276780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#276830000000
0$
0)
#276840000000
1"
1'
b0 +
b0 1
#276890000000
0"
0'
#276900000000
1#
1(
b101111101100100 +
b101111101100100 1
#276950000000
0#
0(
#276960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#277010000000
0$
0)
#277020000000
1"
1'
b0 +
b0 1
#277070000000
0"
0'
#277080000000
1#
1(
b101111101100100 +
b101111101100100 1
#277130000000
0#
0(
#277140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#277190000000
0$
0)
#277200000000
1"
1'
b0 +
b0 1
#277250000000
0"
0'
#277260000000
1#
1(
b101111101100100 +
b101111101100100 1
#277310000000
0#
0(
#277320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#277370000000
0$
0)
#277380000000
1"
1'
b0 +
b0 1
#277430000000
0"
0'
#277440000000
1#
1(
b101111101100100 +
b101111101100100 1
#277490000000
0#
0(
#277500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#277550000000
0$
0)
#277560000000
1"
1'
b0 +
b0 1
#277610000000
0"
0'
#277620000000
1#
1(
b101111101100100 +
b101111101100100 1
#277670000000
0#
0(
#277680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#277730000000
0$
0)
#277740000000
1"
1'
b0 +
b0 1
#277790000000
0"
0'
#277800000000
1#
1(
b101111101100100 +
b101111101100100 1
#277850000000
0#
0(
#277860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#277910000000
0$
0)
#277920000000
1"
1'
b0 +
b0 1
#277970000000
0"
0'
#277980000000
1#
1(
b101111101100100 +
b101111101100100 1
#278030000000
0#
0(
#278040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#278090000000
0$
0)
#278100000000
1"
1'
b0 +
b0 1
#278150000000
0"
0'
#278160000000
1#
1(
b101111101100100 +
b101111101100100 1
#278210000000
0#
0(
#278220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#278270000000
0$
0)
#278280000000
1"
1'
b0 +
b0 1
#278330000000
0"
0'
#278340000000
1#
1(
b101111101100100 +
b101111101100100 1
#278390000000
0#
0(
#278400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#278450000000
0$
0)
#278460000000
1"
1'
b0 +
b0 1
#278510000000
0"
0'
#278520000000
1#
1(
b101111101100100 +
b101111101100100 1
#278570000000
0#
0(
#278580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#278630000000
0$
0)
#278640000000
1"
1'
b0 +
b0 1
#278690000000
0"
0'
#278700000000
1#
1(
b101111101100100 +
b101111101100100 1
#278750000000
0#
0(
#278760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#278810000000
0$
0)
#278820000000
1"
1'
b0 +
b0 1
#278870000000
0"
0'
#278880000000
1#
1(
b101111101100100 +
b101111101100100 1
#278930000000
0#
0(
#278940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#278990000000
0$
0)
#279000000000
1"
1'
b0 +
b0 1
#279050000000
0"
0'
#279060000000
1#
1(
b101111101100100 +
b101111101100100 1
#279110000000
0#
0(
#279120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#279170000000
0$
0)
#279180000000
1"
1'
b0 +
b0 1
#279230000000
0"
0'
#279240000000
1#
1(
b101111101100100 +
b101111101100100 1
#279290000000
0#
0(
#279300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#279350000000
0$
0)
#279360000000
1"
1'
b0 +
b0 1
#279410000000
0"
0'
#279420000000
1#
1(
b101111101100100 +
b101111101100100 1
#279470000000
0#
0(
#279480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#279530000000
0$
0)
#279540000000
1"
1'
b0 +
b0 1
#279590000000
0"
0'
#279600000000
1#
1(
b101111101100100 +
b101111101100100 1
#279650000000
0#
0(
#279660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#279710000000
0$
0)
#279720000000
1"
1'
b0 +
b0 1
#279770000000
0"
0'
#279780000000
1#
1(
b101111101100100 +
b101111101100100 1
#279830000000
0#
0(
#279840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#279890000000
0$
0)
#279900000000
1"
1'
b0 +
b0 1
#279950000000
0"
0'
#279960000000
1#
1(
b101111101100100 +
b101111101100100 1
#280010000000
0#
0(
#280020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#280070000000
0$
0)
#280080000000
1"
1'
b0 +
b0 1
#280130000000
0"
0'
#280140000000
1#
1(
b101111101100100 +
b101111101100100 1
#280190000000
0#
0(
#280200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#280250000000
0$
0)
#280260000000
1"
1'
b0 +
b0 1
#280310000000
0"
0'
#280320000000
1#
1(
b101111101100100 +
b101111101100100 1
#280370000000
0#
0(
#280380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#280430000000
0$
0)
#280440000000
1"
1'
b0 +
b0 1
#280490000000
0"
0'
#280500000000
1#
1(
b101111101100100 +
b101111101100100 1
#280550000000
0#
0(
#280560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#280610000000
0$
0)
#280620000000
1"
1'
b0 +
b0 1
#280670000000
0"
0'
#280680000000
1#
1(
b101111101100100 +
b101111101100100 1
#280730000000
0#
0(
#280740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#280790000000
0$
0)
#280800000000
1"
1'
b0 +
b0 1
#280850000000
0"
0'
#280860000000
1#
1(
b101111101100100 +
b101111101100100 1
#280910000000
0#
0(
#280920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#280970000000
0$
0)
#280980000000
1"
1'
b0 +
b0 1
#281030000000
0"
0'
#281040000000
1#
1(
b101111101100100 +
b101111101100100 1
#281090000000
0#
0(
#281100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#281150000000
0$
0)
#281160000000
1"
1'
b0 +
b0 1
#281210000000
0"
0'
#281220000000
1#
1(
b101111101100100 +
b101111101100100 1
#281270000000
0#
0(
#281280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#281330000000
0$
0)
#281340000000
1"
1'
b0 +
b0 1
#281390000000
0"
0'
#281400000000
1#
1(
b101111101100100 +
b101111101100100 1
#281450000000
0#
0(
#281460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#281510000000
0$
0)
#281520000000
1"
1'
b0 +
b0 1
#281570000000
0"
0'
#281580000000
1#
1(
b101111101100100 +
b101111101100100 1
#281630000000
0#
0(
#281640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#281690000000
0$
0)
#281700000000
1"
1'
b0 +
b0 1
#281750000000
0"
0'
#281760000000
1#
1(
b101111101100100 +
b101111101100100 1
#281810000000
0#
0(
#281820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#281870000000
0$
0)
#281880000000
1"
1'
b0 +
b0 1
#281930000000
0"
0'
#281940000000
1#
1(
b101111101100100 +
b101111101100100 1
#281990000000
0#
0(
#282000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#282050000000
0$
0)
#282060000000
1"
1'
b0 +
b0 1
#282110000000
0"
0'
#282120000000
1#
1(
b101111101100100 +
b101111101100100 1
#282170000000
0#
0(
#282180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#282230000000
0$
0)
#282240000000
1"
1'
b0 +
b0 1
#282290000000
0"
0'
#282300000000
1#
1(
b101111101100100 +
b101111101100100 1
#282350000000
0#
0(
#282360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#282410000000
0$
0)
#282420000000
1"
1'
b0 +
b0 1
#282470000000
0"
0'
#282480000000
1#
1(
b101111101100100 +
b101111101100100 1
#282530000000
0#
0(
#282540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#282590000000
0$
0)
#282600000000
1"
1'
b0 +
b0 1
#282650000000
0"
0'
#282660000000
1#
1(
b101111101100100 +
b101111101100100 1
#282710000000
0#
0(
#282720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#282770000000
0$
0)
#282780000000
1"
1'
b0 +
b0 1
#282830000000
0"
0'
#282840000000
1#
1(
b101111101100100 +
b101111101100100 1
#282890000000
0#
0(
#282900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#282950000000
0$
0)
#282960000000
1"
1'
b0 +
b0 1
#283010000000
0"
0'
#283020000000
1#
1(
b101111101100100 +
b101111101100100 1
#283070000000
0#
0(
#283080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#283130000000
0$
0)
#283140000000
1"
1'
b0 +
b0 1
#283190000000
0"
0'
#283200000000
1#
1(
b101111101100100 +
b101111101100100 1
#283250000000
0#
0(
#283260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#283310000000
0$
0)
#283320000000
1"
1'
b0 +
b0 1
#283370000000
0"
0'
#283380000000
1#
1(
b101111101100100 +
b101111101100100 1
#283430000000
0#
0(
#283440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#283490000000
0$
0)
#283500000000
1"
1'
b0 +
b0 1
#283550000000
0"
0'
#283560000000
1#
1(
b101111101100100 +
b101111101100100 1
#283610000000
0#
0(
#283620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#283670000000
0$
0)
#283680000000
1"
1'
b0 +
b0 1
#283730000000
0"
0'
#283740000000
1#
1(
b101111101100100 +
b101111101100100 1
#283790000000
0#
0(
#283800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#283850000000
0$
0)
#283860000000
1"
1'
b0 +
b0 1
#283910000000
0"
0'
#283920000000
1#
1(
b101111101100100 +
b101111101100100 1
#283970000000
0#
0(
#283980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#284030000000
0$
0)
#284040000000
1"
1'
b0 +
b0 1
#284090000000
0"
0'
#284100000000
1#
1(
b101111101100100 +
b101111101100100 1
#284150000000
0#
0(
#284160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#284210000000
0$
0)
#284220000000
1"
1'
b0 +
b0 1
#284270000000
0"
0'
#284280000000
1#
1(
b101111101100100 +
b101111101100100 1
#284330000000
0#
0(
#284340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#284390000000
0$
0)
#284400000000
1"
1'
b0 +
b0 1
#284450000000
0"
0'
#284460000000
1#
1(
b101111101100100 +
b101111101100100 1
#284510000000
0#
0(
#284520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#284570000000
0$
0)
#284580000000
1"
1'
b0 +
b0 1
#284630000000
0"
0'
#284640000000
1#
1(
b101111101100100 +
b101111101100100 1
#284690000000
0#
0(
#284700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#284750000000
0$
0)
#284760000000
1"
1'
b0 +
b0 1
#284810000000
0"
0'
#284820000000
1#
1(
b101111101100100 +
b101111101100100 1
#284870000000
0#
0(
#284880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#284930000000
0$
0)
#284940000000
1"
1'
b0 +
b0 1
#284990000000
0"
0'
#285000000000
1#
1(
b101111101100100 +
b101111101100100 1
#285050000000
0#
0(
#285060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#285110000000
0$
0)
#285120000000
1"
1'
b0 +
b0 1
#285170000000
0"
0'
#285180000000
1#
1(
b101111101100100 +
b101111101100100 1
#285230000000
0#
0(
#285240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#285290000000
0$
0)
#285300000000
1"
1'
b0 +
b0 1
#285350000000
0"
0'
#285360000000
1#
1(
b101111101100100 +
b101111101100100 1
#285410000000
0#
0(
#285420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#285470000000
0$
0)
#285480000000
1"
1'
b0 +
b0 1
#285530000000
0"
0'
#285540000000
1#
1(
b101111101100100 +
b101111101100100 1
#285590000000
0#
0(
#285600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#285650000000
0$
0)
#285660000000
1"
1'
b0 +
b0 1
#285710000000
0"
0'
#285720000000
1#
1(
b101111101100100 +
b101111101100100 1
#285770000000
0#
0(
#285780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#285830000000
0$
0)
#285840000000
1"
1'
b0 +
b0 1
#285890000000
0"
0'
#285900000000
1#
1(
b101111101100100 +
b101111101100100 1
#285950000000
0#
0(
#285960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#286010000000
0$
0)
#286020000000
1"
1'
b0 +
b0 1
#286070000000
0"
0'
#286080000000
1#
1(
b101111101100100 +
b101111101100100 1
#286130000000
0#
0(
#286140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#286190000000
0$
0)
#286200000000
1"
1'
b0 +
b0 1
#286250000000
0"
0'
#286260000000
1#
1(
b101111101100100 +
b101111101100100 1
#286310000000
0#
0(
#286320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#286370000000
0$
0)
#286380000000
1"
1'
b0 +
b0 1
#286430000000
0"
0'
#286440000000
1#
1(
b101111101100100 +
b101111101100100 1
#286490000000
0#
0(
#286500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#286550000000
0$
0)
#286560000000
1"
1'
b0 +
b0 1
#286610000000
0"
0'
#286620000000
1#
1(
b101111101100100 +
b101111101100100 1
#286670000000
0#
0(
#286680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#286730000000
0$
0)
#286740000000
1"
1'
b0 +
b0 1
#286790000000
0"
0'
#286800000000
1#
1(
b101111101100100 +
b101111101100100 1
#286850000000
0#
0(
#286860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#286910000000
0$
0)
#286920000000
1"
1'
b0 +
b0 1
#286970000000
0"
0'
#286980000000
1#
1(
b101111101100100 +
b101111101100100 1
#287030000000
0#
0(
#287040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#287090000000
0$
0)
#287100000000
1"
1'
b0 +
b0 1
#287150000000
0"
0'
#287160000000
1#
1(
b101111101100100 +
b101111101100100 1
#287210000000
0#
0(
#287220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#287270000000
0$
0)
#287280000000
1"
1'
b0 +
b0 1
#287330000000
0"
0'
#287340000000
1#
1(
b101111101100100 +
b101111101100100 1
#287390000000
0#
0(
#287400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#287450000000
0$
0)
#287460000000
1"
1'
b0 +
b0 1
#287510000000
0"
0'
#287520000000
1#
1(
b101111101100100 +
b101111101100100 1
#287570000000
0#
0(
#287580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#287630000000
0$
0)
#287640000000
1"
1'
b0 +
b0 1
#287690000000
0"
0'
#287700000000
1#
1(
b101111101100100 +
b101111101100100 1
#287750000000
0#
0(
#287760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#287810000000
0$
0)
#287820000000
1"
1'
b0 +
b0 1
#287870000000
0"
0'
#287880000000
1#
1(
b101111101100100 +
b101111101100100 1
#287930000000
0#
0(
#287940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#287990000000
0$
0)
#288000000000
1"
1'
b0 +
b0 1
#288050000000
0"
0'
#288060000000
1#
1(
b101111101100100 +
b101111101100100 1
#288110000000
0#
0(
#288120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#288170000000
0$
0)
#288180000000
1"
1'
b0 +
b0 1
#288230000000
0"
0'
#288240000000
1#
1(
b101111101100100 +
b101111101100100 1
#288290000000
0#
0(
#288300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#288350000000
0$
0)
#288360000000
1"
1'
b0 +
b0 1
#288410000000
0"
0'
#288420000000
1#
1(
b101111101100100 +
b101111101100100 1
#288470000000
0#
0(
#288480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#288530000000
0$
0)
#288540000000
1"
1'
b0 +
b0 1
#288590000000
0"
0'
#288600000000
1#
1(
b101111101100100 +
b101111101100100 1
#288650000000
0#
0(
#288660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#288710000000
0$
0)
#288720000000
1"
1'
b0 +
b0 1
#288770000000
0"
0'
#288780000000
1#
1(
b101111101100100 +
b101111101100100 1
#288830000000
0#
0(
#288840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#288890000000
0$
0)
#288900000000
1"
1'
b0 +
b0 1
#288950000000
0"
0'
#288960000000
1#
1(
b101111101100100 +
b101111101100100 1
#289010000000
0#
0(
#289020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#289070000000
0$
0)
#289080000000
1"
1'
b0 +
b0 1
#289130000000
0"
0'
#289140000000
1#
1(
b101111101100100 +
b101111101100100 1
#289190000000
0#
0(
#289200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#289250000000
0$
0)
#289260000000
1"
1'
b0 +
b0 1
#289310000000
0"
0'
#289320000000
1#
1(
b101111101100100 +
b101111101100100 1
#289370000000
0#
0(
#289380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#289430000000
0$
0)
#289440000000
1"
1'
b0 +
b0 1
#289490000000
0"
0'
#289500000000
1#
1(
b101111101100100 +
b101111101100100 1
#289550000000
0#
0(
#289560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#289610000000
0$
0)
#289620000000
1"
1'
b0 +
b0 1
#289670000000
0"
0'
#289680000000
1#
1(
b101111101100100 +
b101111101100100 1
#289730000000
0#
0(
#289740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#289790000000
0$
0)
#289800000000
1"
1'
b0 +
b0 1
#289850000000
0"
0'
#289860000000
1#
1(
b101111101100100 +
b101111101100100 1
#289910000000
0#
0(
#289920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#289970000000
0$
0)
#289980000000
1"
1'
b0 +
b0 1
#290030000000
0"
0'
#290040000000
1#
1(
b101111101100100 +
b101111101100100 1
#290090000000
0#
0(
#290100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#290150000000
0$
0)
#290160000000
1"
1'
b0 +
b0 1
#290210000000
0"
0'
#290220000000
1#
1(
b101111101100100 +
b101111101100100 1
#290270000000
0#
0(
#290280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#290330000000
0$
0)
#290340000000
1"
1'
b0 +
b0 1
#290390000000
0"
0'
#290400000000
1#
1(
b101111101100100 +
b101111101100100 1
#290450000000
0#
0(
#290460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#290510000000
0$
0)
#290520000000
1"
1'
b0 +
b0 1
#290570000000
0"
0'
#290580000000
1#
1(
b101111101100100 +
b101111101100100 1
#290630000000
0#
0(
#290640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#290690000000
0$
0)
#290700000000
1"
1'
b0 +
b0 1
#290750000000
0"
0'
#290760000000
1#
1(
b101111101100100 +
b101111101100100 1
#290810000000
0#
0(
#290820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#290870000000
0$
0)
#290880000000
1"
1'
b0 +
b0 1
#290930000000
0"
0'
#290940000000
1#
1(
b101111101100100 +
b101111101100100 1
#290990000000
0#
0(
#291000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#291050000000
0$
0)
#291060000000
1"
1'
b0 +
b0 1
#291110000000
0"
0'
#291120000000
1#
1(
b101111101100100 +
b101111101100100 1
#291170000000
0#
0(
#291180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#291230000000
0$
0)
#291240000000
1"
1'
b0 +
b0 1
#291290000000
0"
0'
#291300000000
1#
1(
b101111101100100 +
b101111101100100 1
#291350000000
0#
0(
#291360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#291410000000
0$
0)
#291420000000
1"
1'
b0 +
b0 1
#291470000000
0"
0'
#291480000000
1#
1(
b101111101100100 +
b101111101100100 1
#291530000000
0#
0(
#291540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#291590000000
0$
0)
#291600000000
1"
1'
b0 +
b0 1
#291650000000
0"
0'
#291660000000
1#
1(
b101111101100100 +
b101111101100100 1
#291710000000
0#
0(
#291720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#291770000000
0$
0)
#291780000000
1"
1'
b0 +
b0 1
#291830000000
0"
0'
#291840000000
1#
1(
b101111101100100 +
b101111101100100 1
#291890000000
0#
0(
#291900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#291950000000
0$
0)
#291960000000
1"
1'
b0 +
b0 1
#292010000000
0"
0'
#292020000000
1#
1(
b101111101100100 +
b101111101100100 1
#292070000000
0#
0(
#292080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#292130000000
0$
0)
#292140000000
1"
1'
b0 +
b0 1
#292190000000
0"
0'
#292200000000
1#
1(
b101111101100100 +
b101111101100100 1
#292250000000
0#
0(
#292260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#292310000000
0$
0)
#292320000000
1"
1'
b0 +
b0 1
#292370000000
0"
0'
#292380000000
1#
1(
b101111101100100 +
b101111101100100 1
#292430000000
0#
0(
#292440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#292490000000
0$
0)
#292500000000
1"
1'
b0 +
b0 1
#292550000000
0"
0'
#292560000000
1#
1(
b101111101100100 +
b101111101100100 1
#292610000000
0#
0(
#292620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#292670000000
0$
0)
#292680000000
1"
1'
b0 +
b0 1
#292730000000
0"
0'
#292740000000
1#
1(
b101111101100100 +
b101111101100100 1
#292790000000
0#
0(
#292800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#292850000000
0$
0)
#292860000000
1"
1'
b0 +
b0 1
#292910000000
0"
0'
#292920000000
1#
1(
b101111101100100 +
b101111101100100 1
#292970000000
0#
0(
#292980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#293030000000
0$
0)
#293040000000
1"
1'
b0 +
b0 1
#293090000000
0"
0'
#293100000000
1#
1(
b101111101100100 +
b101111101100100 1
#293150000000
0#
0(
#293160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#293210000000
0$
0)
#293220000000
1"
1'
b0 +
b0 1
#293270000000
0"
0'
#293280000000
1#
1(
b101111101100100 +
b101111101100100 1
#293330000000
0#
0(
#293340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#293390000000
0$
0)
#293400000000
1"
1'
b0 +
b0 1
#293450000000
0"
0'
#293460000000
1#
1(
b101111101100100 +
b101111101100100 1
#293510000000
0#
0(
#293520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#293570000000
0$
0)
#293580000000
1"
1'
b0 +
b0 1
#293630000000
0"
0'
#293640000000
1#
1(
b101111101100100 +
b101111101100100 1
#293690000000
0#
0(
#293700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#293750000000
0$
0)
#293760000000
1"
1'
b0 +
b0 1
#293810000000
0"
0'
#293820000000
1#
1(
b101111101100100 +
b101111101100100 1
#293870000000
0#
0(
#293880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#293930000000
0$
0)
#293940000000
1"
1'
b0 +
b0 1
#293990000000
0"
0'
#294000000000
1#
1(
b101111101100100 +
b101111101100100 1
#294050000000
0#
0(
#294060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#294110000000
0$
0)
#294120000000
1"
1'
b0 +
b0 1
#294170000000
0"
0'
#294180000000
1#
1(
b101111101100100 +
b101111101100100 1
#294230000000
0#
0(
#294240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#294290000000
0$
0)
#294300000000
1"
1'
b0 +
b0 1
#294350000000
0"
0'
#294360000000
1#
1(
b101111101100100 +
b101111101100100 1
#294410000000
0#
0(
#294420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#294470000000
0$
0)
#294480000000
1"
1'
b0 +
b0 1
#294530000000
0"
0'
#294540000000
1#
1(
b101111101100100 +
b101111101100100 1
#294590000000
0#
0(
#294600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#294650000000
0$
0)
#294660000000
1"
1'
b0 +
b0 1
#294710000000
0"
0'
#294720000000
1#
1(
b101111101100100 +
b101111101100100 1
#294770000000
0#
0(
#294780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#294830000000
0$
0)
#294840000000
1"
1'
b0 +
b0 1
#294890000000
0"
0'
#294900000000
1#
1(
b101111101100100 +
b101111101100100 1
#294950000000
0#
0(
#294960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#295010000000
0$
0)
#295020000000
1"
1'
b0 +
b0 1
#295070000000
0"
0'
#295080000000
1#
1(
b101111101100100 +
b101111101100100 1
#295130000000
0#
0(
#295140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#295190000000
0$
0)
#295200000000
1"
1'
b0 +
b0 1
#295250000000
0"
0'
#295260000000
1#
1(
b101111101100100 +
b101111101100100 1
#295310000000
0#
0(
#295320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#295370000000
0$
0)
#295380000000
1"
1'
b0 +
b0 1
#295430000000
0"
0'
#295440000000
1#
1(
b101111101100100 +
b101111101100100 1
#295490000000
0#
0(
#295500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#295550000000
0$
0)
#295560000000
1"
1'
b0 +
b0 1
#295610000000
0"
0'
#295620000000
1#
1(
b101111101100100 +
b101111101100100 1
#295670000000
0#
0(
#295680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#295730000000
0$
0)
#295740000000
1"
1'
b0 +
b0 1
#295790000000
0"
0'
#295800000000
1#
1(
b101111101100100 +
b101111101100100 1
#295850000000
0#
0(
#295860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#295910000000
0$
0)
#295920000000
1"
1'
b0 +
b0 1
#295970000000
0"
0'
#295980000000
1#
1(
b101111101100100 +
b101111101100100 1
#296030000000
0#
0(
#296040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#296090000000
0$
0)
#296100000000
1"
1'
b0 +
b0 1
#296150000000
0"
0'
#296160000000
1#
1(
b101111101100100 +
b101111101100100 1
#296210000000
0#
0(
#296220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#296270000000
0$
0)
#296280000000
1"
1'
b0 +
b0 1
#296330000000
0"
0'
#296340000000
1#
1(
b101111101100100 +
b101111101100100 1
#296390000000
0#
0(
#296400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#296450000000
0$
0)
#296460000000
1"
1'
b0 +
b0 1
#296510000000
0"
0'
#296520000000
1#
1(
b101111101100100 +
b101111101100100 1
#296570000000
0#
0(
#296580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#296630000000
0$
0)
#296640000000
1"
1'
b0 +
b0 1
#296690000000
0"
0'
#296700000000
1#
1(
b101111101100100 +
b101111101100100 1
#296750000000
0#
0(
#296760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#296810000000
0$
0)
#296820000000
1"
1'
b0 +
b0 1
#296870000000
0"
0'
#296880000000
1#
1(
b101111101100100 +
b101111101100100 1
#296930000000
0#
0(
#296940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#296990000000
0$
0)
#297000000000
1"
1'
b0 +
b0 1
#297050000000
0"
0'
#297060000000
1#
1(
b101111101100100 +
b101111101100100 1
#297110000000
0#
0(
#297120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#297170000000
0$
0)
#297180000000
1"
1'
b0 +
b0 1
#297230000000
0"
0'
#297240000000
1#
1(
b101111101100100 +
b101111101100100 1
#297290000000
0#
0(
#297300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#297350000000
0$
0)
#297360000000
1"
1'
b0 +
b0 1
#297410000000
0"
0'
#297420000000
1#
1(
b101111101100100 +
b101111101100100 1
#297470000000
0#
0(
#297480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#297530000000
0$
0)
#297540000000
1"
1'
b0 +
b0 1
#297590000000
0"
0'
#297600000000
1#
1(
b101111101100100 +
b101111101100100 1
#297650000000
0#
0(
#297660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#297710000000
0$
0)
#297720000000
1"
1'
b0 +
b0 1
#297770000000
0"
0'
#297780000000
1#
1(
b101111101100100 +
b101111101100100 1
#297830000000
0#
0(
#297840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#297890000000
0$
0)
#297900000000
1"
1'
b0 +
b0 1
#297950000000
0"
0'
#297960000000
1#
1(
b101111101100100 +
b101111101100100 1
#298010000000
0#
0(
#298020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#298070000000
0$
0)
#298080000000
1"
1'
b0 +
b0 1
#298130000000
0"
0'
#298140000000
1#
1(
b101111101100100 +
b101111101100100 1
#298190000000
0#
0(
#298200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#298250000000
0$
0)
#298260000000
1"
1'
b0 +
b0 1
#298310000000
0"
0'
#298320000000
1#
1(
b101111101100100 +
b101111101100100 1
#298370000000
0#
0(
#298380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#298430000000
0$
0)
#298440000000
1"
1'
b0 +
b0 1
#298490000000
0"
0'
#298500000000
1#
1(
b101111101100100 +
b101111101100100 1
#298550000000
0#
0(
#298560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#298610000000
0$
0)
#298620000000
1"
1'
b0 +
b0 1
#298670000000
0"
0'
#298680000000
1#
1(
b101111101100100 +
b101111101100100 1
#298730000000
0#
0(
#298740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#298790000000
0$
0)
#298800000000
1"
1'
b0 +
b0 1
#298850000000
0"
0'
#298860000000
1#
1(
b101111101100100 +
b101111101100100 1
#298910000000
0#
0(
#298920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#298970000000
0$
0)
#298980000000
1"
1'
b0 +
b0 1
#299030000000
0"
0'
#299040000000
1#
1(
b101111101100100 +
b101111101100100 1
#299090000000
0#
0(
#299100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#299150000000
0$
0)
#299160000000
1"
1'
b0 +
b0 1
#299210000000
0"
0'
#299220000000
1#
1(
b101111101100100 +
b101111101100100 1
#299270000000
0#
0(
#299280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#299330000000
0$
0)
#299340000000
1"
1'
b0 +
b0 1
#299390000000
0"
0'
#299400000000
1#
1(
b101111101100100 +
b101111101100100 1
#299450000000
0#
0(
#299460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#299510000000
0$
0)
#299520000000
1"
1'
b0 +
b0 1
#299570000000
0"
0'
#299580000000
1#
1(
b101111101100100 +
b101111101100100 1
#299630000000
0#
0(
#299640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#299690000000
0$
0)
#299700000000
1"
1'
b0 +
b0 1
#299750000000
0"
0'
#299760000000
1#
1(
b101111101100100 +
b101111101100100 1
#299810000000
0#
0(
#299820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#299870000000
0$
0)
#299880000000
1"
1'
b0 +
b0 1
#299930000000
0"
0'
#299940000000
1#
1(
b101111101100100 +
b101111101100100 1
#299990000000
0#
0(
#300000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#300050000000
0$
0)
#300060000000
1"
1'
b0 +
b0 1
#300110000000
0"
0'
#300120000000
1#
1(
b101111101100100 +
b101111101100100 1
#300170000000
0#
0(
#300180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#300230000000
0$
0)
#300240000000
1"
1'
b0 +
b0 1
#300290000000
0"
0'
#300300000000
1#
1(
b101111101100100 +
b101111101100100 1
#300350000000
0#
0(
#300360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#300410000000
0$
0)
#300420000000
1"
1'
b0 +
b0 1
#300470000000
0"
0'
#300480000000
1#
1(
b101111101100100 +
b101111101100100 1
#300530000000
0#
0(
#300540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#300590000000
0$
0)
#300600000000
1"
1'
b0 +
b0 1
#300650000000
0"
0'
#300660000000
1#
1(
b101111101100100 +
b101111101100100 1
#300710000000
0#
0(
#300720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#300770000000
0$
0)
#300780000000
1"
1'
b0 +
b0 1
#300830000000
0"
0'
#300840000000
1#
1(
b101111101100100 +
b101111101100100 1
#300890000000
0#
0(
#300900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#300950000000
0$
0)
#300960000000
1"
1'
b0 +
b0 1
#301010000000
0"
0'
#301020000000
1#
1(
b101111101100100 +
b101111101100100 1
#301070000000
0#
0(
#301080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#301130000000
0$
0)
#301140000000
1"
1'
b0 +
b0 1
#301190000000
0"
0'
#301200000000
1#
1(
b101111101100100 +
b101111101100100 1
#301250000000
0#
0(
#301260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#301310000000
0$
0)
#301320000000
1"
1'
b0 +
b0 1
#301370000000
0"
0'
#301380000000
1#
1(
b101111101100100 +
b101111101100100 1
#301430000000
0#
0(
#301440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#301490000000
0$
0)
#301500000000
1"
1'
b0 +
b0 1
#301550000000
0"
0'
#301560000000
1#
1(
b101111101100100 +
b101111101100100 1
#301610000000
0#
0(
#301620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#301670000000
0$
0)
#301680000000
1"
1'
b0 +
b0 1
#301730000000
0"
0'
#301740000000
1#
1(
b101111101100100 +
b101111101100100 1
#301790000000
0#
0(
#301800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#301850000000
0$
0)
#301860000000
1"
1'
b0 +
b0 1
#301910000000
0"
0'
#301920000000
1#
1(
b101111101100100 +
b101111101100100 1
#301970000000
0#
0(
#301980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#302030000000
0$
0)
#302040000000
1"
1'
b0 +
b0 1
#302090000000
0"
0'
#302100000000
1#
1(
b101111101100100 +
b101111101100100 1
#302150000000
0#
0(
#302160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#302210000000
0$
0)
#302220000000
1"
1'
b0 +
b0 1
#302270000000
0"
0'
#302280000000
1#
1(
b101111101100100 +
b101111101100100 1
#302330000000
0#
0(
#302340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#302390000000
0$
0)
#302400000000
1"
1'
b0 +
b0 1
#302450000000
0"
0'
#302460000000
1#
1(
b101111101100100 +
b101111101100100 1
#302510000000
0#
0(
#302520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#302570000000
0$
0)
#302580000000
1"
1'
b0 +
b0 1
#302630000000
0"
0'
#302640000000
1#
1(
b101111101100100 +
b101111101100100 1
#302690000000
0#
0(
#302700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#302750000000
0$
0)
#302760000000
1"
1'
b0 +
b0 1
#302810000000
0"
0'
#302820000000
1#
1(
b101111101100100 +
b101111101100100 1
#302870000000
0#
0(
#302880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#302930000000
0$
0)
#302940000000
1"
1'
b0 +
b0 1
#302990000000
0"
0'
#303000000000
1#
1(
b101111101100100 +
b101111101100100 1
#303050000000
0#
0(
#303060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#303110000000
0$
0)
#303120000000
1"
1'
b0 +
b0 1
#303170000000
0"
0'
#303180000000
1#
1(
b101111101100100 +
b101111101100100 1
#303230000000
0#
0(
#303240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#303290000000
0$
0)
#303300000000
1"
1'
b0 +
b0 1
#303350000000
0"
0'
#303360000000
1#
1(
b101111101100100 +
b101111101100100 1
#303410000000
0#
0(
#303420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#303470000000
0$
0)
#303480000000
1"
1'
b0 +
b0 1
#303530000000
0"
0'
#303540000000
1#
1(
b101111101100100 +
b101111101100100 1
#303590000000
0#
0(
#303600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#303650000000
0$
0)
#303660000000
1"
1'
b0 +
b0 1
#303710000000
0"
0'
#303720000000
1#
1(
b101111101100100 +
b101111101100100 1
#303770000000
0#
0(
#303780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#303830000000
0$
0)
#303840000000
1"
1'
b0 +
b0 1
#303890000000
0"
0'
#303900000000
1#
1(
b101111101100100 +
b101111101100100 1
#303950000000
0#
0(
#303960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#304010000000
0$
0)
#304020000000
1"
1'
b0 +
b0 1
#304070000000
0"
0'
#304080000000
1#
1(
b101111101100100 +
b101111101100100 1
#304130000000
0#
0(
#304140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#304190000000
0$
0)
#304200000000
1"
1'
b0 +
b0 1
#304250000000
0"
0'
#304260000000
1#
1(
b101111101100100 +
b101111101100100 1
#304310000000
0#
0(
#304320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#304370000000
0$
0)
#304380000000
1"
1'
b0 +
b0 1
#304430000000
0"
0'
#304440000000
1#
1(
b101111101100100 +
b101111101100100 1
#304490000000
0#
0(
#304500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#304550000000
0$
0)
#304560000000
1"
1'
b0 +
b0 1
#304610000000
0"
0'
#304620000000
1#
1(
b101111101100100 +
b101111101100100 1
#304670000000
0#
0(
#304680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#304730000000
0$
0)
#304740000000
1"
1'
b0 +
b0 1
#304790000000
0"
0'
#304800000000
1#
1(
b101111101100100 +
b101111101100100 1
#304850000000
0#
0(
#304860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#304910000000
0$
0)
#304920000000
1"
1'
b0 +
b0 1
#304970000000
0"
0'
#304980000000
1#
1(
b101111101100100 +
b101111101100100 1
#305030000000
0#
0(
#305040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#305090000000
0$
0)
#305100000000
1"
1'
b0 +
b0 1
#305150000000
0"
0'
#305160000000
1#
1(
b101111101100100 +
b101111101100100 1
#305210000000
0#
0(
#305220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#305270000000
0$
0)
#305280000000
1"
1'
b0 +
b0 1
#305330000000
0"
0'
#305340000000
1#
1(
b101111101100100 +
b101111101100100 1
#305390000000
0#
0(
#305400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#305450000000
0$
0)
#305460000000
1"
1'
b0 +
b0 1
#305510000000
0"
0'
#305520000000
1#
1(
b101111101100100 +
b101111101100100 1
#305570000000
0#
0(
#305580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#305630000000
0$
0)
#305640000000
1"
1'
b0 +
b0 1
#305690000000
0"
0'
#305700000000
1#
1(
b101111101100100 +
b101111101100100 1
#305750000000
0#
0(
#305760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#305810000000
0$
0)
#305820000000
1"
1'
b0 +
b0 1
#305870000000
0"
0'
#305880000000
1#
1(
b101111101100100 +
b101111101100100 1
#305930000000
0#
0(
#305940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#305990000000
0$
0)
#306000000000
1"
1'
b0 +
b0 1
#306050000000
0"
0'
#306060000000
1#
1(
b101111101100100 +
b101111101100100 1
#306110000000
0#
0(
#306120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#306170000000
0$
0)
#306180000000
1"
1'
b0 +
b0 1
#306230000000
0"
0'
#306240000000
1#
1(
b101111101100100 +
b101111101100100 1
#306290000000
0#
0(
#306300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#306350000000
0$
0)
#306360000000
1"
1'
b0 +
b0 1
#306410000000
0"
0'
#306420000000
1#
1(
b101111101100100 +
b101111101100100 1
#306470000000
0#
0(
#306480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#306530000000
0$
0)
#306540000000
1"
1'
b0 +
b0 1
#306590000000
0"
0'
#306600000000
1#
1(
b101111101100100 +
b101111101100100 1
#306650000000
0#
0(
#306660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#306710000000
0$
0)
#306720000000
1"
1'
b0 +
b0 1
#306770000000
0"
0'
#306780000000
1#
1(
b101111101100100 +
b101111101100100 1
#306830000000
0#
0(
#306840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#306890000000
0$
0)
#306900000000
1"
1'
b0 +
b0 1
#306950000000
0"
0'
#306960000000
1#
1(
b101111101100100 +
b101111101100100 1
#307010000000
0#
0(
#307020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#307070000000
0$
0)
#307080000000
1"
1'
b0 +
b0 1
#307130000000
0"
0'
#307140000000
1#
1(
b101111101100100 +
b101111101100100 1
#307190000000
0#
0(
#307200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#307250000000
0$
0)
#307260000000
1"
1'
b0 +
b0 1
#307310000000
0"
0'
#307320000000
1#
1(
b101111101100100 +
b101111101100100 1
#307370000000
0#
0(
#307380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#307430000000
0$
0)
#307440000000
1"
1'
b0 +
b0 1
#307490000000
0"
0'
#307500000000
1#
1(
b101111101100100 +
b101111101100100 1
#307550000000
0#
0(
#307560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#307610000000
0$
0)
#307620000000
1"
1'
b0 +
b0 1
#307670000000
0"
0'
#307680000000
1#
1(
b101111101100100 +
b101111101100100 1
#307730000000
0#
0(
#307740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#307790000000
0$
0)
#307800000000
1"
1'
b0 +
b0 1
#307850000000
0"
0'
#307860000000
1#
1(
b101111101100100 +
b101111101100100 1
#307910000000
0#
0(
#307920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#307970000000
0$
0)
#307980000000
1"
1'
b0 +
b0 1
#308030000000
0"
0'
#308040000000
1#
1(
b101111101100100 +
b101111101100100 1
#308090000000
0#
0(
#308100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#308150000000
0$
0)
#308160000000
1"
1'
b0 +
b0 1
#308210000000
0"
0'
#308220000000
1#
1(
b101111101100100 +
b101111101100100 1
#308270000000
0#
0(
#308280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#308330000000
0$
0)
#308340000000
1"
1'
b0 +
b0 1
#308390000000
0"
0'
#308400000000
1#
1(
b101111101100100 +
b101111101100100 1
#308450000000
0#
0(
#308460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#308510000000
0$
0)
#308520000000
1"
1'
b0 +
b0 1
#308570000000
0"
0'
#308580000000
1#
1(
b101111101100100 +
b101111101100100 1
#308630000000
0#
0(
#308640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#308690000000
0$
0)
#308700000000
1"
1'
b0 +
b0 1
#308750000000
0"
0'
#308760000000
1#
1(
b101111101100100 +
b101111101100100 1
#308810000000
0#
0(
#308820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#308870000000
0$
0)
#308880000000
1"
1'
b0 +
b0 1
#308930000000
0"
0'
#308940000000
1#
1(
b101111101100100 +
b101111101100100 1
#308990000000
0#
0(
#309000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#309050000000
0$
0)
#309060000000
1"
1'
b0 +
b0 1
#309110000000
0"
0'
#309120000000
1#
1(
b101111101100100 +
b101111101100100 1
#309170000000
0#
0(
#309180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#309230000000
0$
0)
#309240000000
1"
1'
b0 +
b0 1
#309290000000
0"
0'
#309300000000
1#
1(
b101111101100100 +
b101111101100100 1
#309350000000
0#
0(
#309360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#309410000000
0$
0)
#309420000000
1"
1'
b0 +
b0 1
#309470000000
0"
0'
#309480000000
1#
1(
b101111101100100 +
b101111101100100 1
#309530000000
0#
0(
#309540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#309590000000
0$
0)
#309600000000
1"
1'
b0 +
b0 1
#309650000000
0"
0'
#309660000000
1#
1(
b101111101100100 +
b101111101100100 1
#309710000000
0#
0(
#309720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#309770000000
0$
0)
#309780000000
1"
1'
b0 +
b0 1
#309830000000
0"
0'
#309840000000
1#
1(
b101111101100100 +
b101111101100100 1
#309890000000
0#
0(
#309900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#309950000000
0$
0)
#309960000000
1"
1'
b0 +
b0 1
#310010000000
0"
0'
#310020000000
1#
1(
b101111101100100 +
b101111101100100 1
#310070000000
0#
0(
#310080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#310130000000
0$
0)
#310140000000
1"
1'
b0 +
b0 1
#310190000000
0"
0'
#310200000000
1#
1(
b101111101100100 +
b101111101100100 1
#310250000000
0#
0(
#310260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#310310000000
0$
0)
#310320000000
1"
1'
b0 +
b0 1
#310370000000
0"
0'
#310380000000
1#
1(
b101111101100100 +
b101111101100100 1
#310430000000
0#
0(
#310440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#310490000000
0$
0)
#310500000000
1"
1'
b0 +
b0 1
#310550000000
0"
0'
#310560000000
1#
1(
b101111101100100 +
b101111101100100 1
#310610000000
0#
0(
#310620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#310670000000
0$
0)
#310680000000
1"
1'
b0 +
b0 1
#310730000000
0"
0'
#310740000000
1#
1(
b101111101100100 +
b101111101100100 1
#310790000000
0#
0(
#310800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#310850000000
0$
0)
#310860000000
1"
1'
b0 +
b0 1
#310910000000
0"
0'
#310920000000
1#
1(
b101111101100100 +
b101111101100100 1
#310970000000
0#
0(
#310980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#311030000000
0$
0)
#311040000000
1"
1'
b0 +
b0 1
#311090000000
0"
0'
#311100000000
1#
1(
b101111101100100 +
b101111101100100 1
#311150000000
0#
0(
#311160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#311210000000
0$
0)
#311220000000
1"
1'
b0 +
b0 1
#311270000000
0"
0'
#311280000000
1#
1(
b101111101100100 +
b101111101100100 1
#311330000000
0#
0(
#311340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#311390000000
0$
0)
#311400000000
1"
1'
b0 +
b0 1
#311450000000
0"
0'
#311460000000
1#
1(
b101111101100100 +
b101111101100100 1
#311510000000
0#
0(
#311520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#311570000000
0$
0)
#311580000000
1"
1'
b0 +
b0 1
#311630000000
0"
0'
#311640000000
1#
1(
b101111101100100 +
b101111101100100 1
#311690000000
0#
0(
#311700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#311750000000
0$
0)
#311760000000
1"
1'
b0 +
b0 1
#311810000000
0"
0'
#311820000000
1#
1(
b101111101100100 +
b101111101100100 1
#311870000000
0#
0(
#311880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#311930000000
0$
0)
#311940000000
1"
1'
b0 +
b0 1
#311990000000
0"
0'
#312000000000
1#
1(
b101111101100100 +
b101111101100100 1
#312050000000
0#
0(
#312060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#312110000000
0$
0)
#312120000000
1"
1'
b0 +
b0 1
#312170000000
0"
0'
#312180000000
1#
1(
b101111101100100 +
b101111101100100 1
#312230000000
0#
0(
#312240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#312290000000
0$
0)
#312300000000
1"
1'
b0 +
b0 1
#312350000000
0"
0'
#312360000000
1#
1(
b101111101100100 +
b101111101100100 1
#312410000000
0#
0(
#312420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#312470000000
0$
0)
#312480000000
1"
1'
b0 +
b0 1
#312530000000
0"
0'
#312540000000
1#
1(
b101111101100100 +
b101111101100100 1
#312590000000
0#
0(
#312600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#312650000000
0$
0)
#312660000000
1"
1'
b0 +
b0 1
#312710000000
0"
0'
#312720000000
1#
1(
b101111101100100 +
b101111101100100 1
#312770000000
0#
0(
#312780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#312830000000
0$
0)
#312840000000
1"
1'
b0 +
b0 1
#312890000000
0"
0'
#312900000000
1#
1(
b101111101100100 +
b101111101100100 1
#312950000000
0#
0(
#312960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#313010000000
0$
0)
#313020000000
1"
1'
b0 +
b0 1
#313070000000
0"
0'
#313080000000
1#
1(
b101111101100100 +
b101111101100100 1
#313130000000
0#
0(
#313140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#313190000000
0$
0)
#313200000000
1"
1'
b0 +
b0 1
#313250000000
0"
0'
#313260000000
1#
1(
b101111101100100 +
b101111101100100 1
#313310000000
0#
0(
#313320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#313370000000
0$
0)
#313380000000
1"
1'
b0 +
b0 1
#313430000000
0"
0'
#313440000000
1#
1(
b101111101100100 +
b101111101100100 1
#313490000000
0#
0(
#313500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#313550000000
0$
0)
#313560000000
1"
1'
b0 +
b0 1
#313610000000
0"
0'
#313620000000
1#
1(
b101111101100100 +
b101111101100100 1
#313670000000
0#
0(
#313680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#313730000000
0$
0)
#313740000000
1"
1'
b0 +
b0 1
#313790000000
0"
0'
#313800000000
1#
1(
b101111101100100 +
b101111101100100 1
#313850000000
0#
0(
#313860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#313910000000
0$
0)
#313920000000
1"
1'
b0 +
b0 1
#313970000000
0"
0'
#313980000000
1#
1(
b101111101100100 +
b101111101100100 1
#314030000000
0#
0(
#314040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#314090000000
0$
0)
#314100000000
1"
1'
b0 +
b0 1
#314150000000
0"
0'
#314160000000
1#
1(
b101111101100100 +
b101111101100100 1
#314210000000
0#
0(
#314220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#314270000000
0$
0)
#314280000000
1"
1'
b0 +
b0 1
#314330000000
0"
0'
#314340000000
1#
1(
b101111101100100 +
b101111101100100 1
#314390000000
0#
0(
#314400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#314450000000
0$
0)
#314460000000
1"
1'
b0 +
b0 1
#314510000000
0"
0'
#314520000000
1#
1(
b101111101100100 +
b101111101100100 1
#314570000000
0#
0(
#314580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#314630000000
0$
0)
#314640000000
1"
1'
b0 +
b0 1
#314690000000
0"
0'
#314700000000
1#
1(
b101111101100100 +
b101111101100100 1
#314750000000
0#
0(
#314760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#314810000000
0$
0)
#314820000000
1"
1'
b0 +
b0 1
#314870000000
0"
0'
#314880000000
1#
1(
b101111101100100 +
b101111101100100 1
#314930000000
0#
0(
#314940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#314990000000
0$
0)
#315000000000
1"
1'
b0 +
b0 1
#315050000000
0"
0'
#315060000000
1#
1(
b101111101100100 +
b101111101100100 1
#315110000000
0#
0(
#315120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#315170000000
0$
0)
#315180000000
1"
1'
b0 +
b0 1
#315230000000
0"
0'
#315240000000
1#
1(
b101111101100100 +
b101111101100100 1
#315290000000
0#
0(
#315300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#315350000000
0$
0)
#315360000000
1"
1'
b0 +
b0 1
#315410000000
0"
0'
#315420000000
1#
1(
b101111101100100 +
b101111101100100 1
#315470000000
0#
0(
#315480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#315530000000
0$
0)
#315540000000
1"
1'
b0 +
b0 1
#315590000000
0"
0'
#315600000000
1#
1(
b101111101100100 +
b101111101100100 1
#315650000000
0#
0(
#315660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#315710000000
0$
0)
#315720000000
1"
1'
b0 +
b0 1
#315770000000
0"
0'
#315780000000
1#
1(
b101111101100100 +
b101111101100100 1
#315830000000
0#
0(
#315840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#315890000000
0$
0)
#315900000000
1"
1'
b0 +
b0 1
#315950000000
0"
0'
#315960000000
1#
1(
b101111101100100 +
b101111101100100 1
#316010000000
0#
0(
#316020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#316070000000
0$
0)
#316080000000
1"
1'
b0 +
b0 1
#316130000000
0"
0'
#316140000000
1#
1(
b101111101100100 +
b101111101100100 1
#316190000000
0#
0(
#316200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#316250000000
0$
0)
#316260000000
1"
1'
b0 +
b0 1
#316310000000
0"
0'
#316320000000
1#
1(
b101111101100100 +
b101111101100100 1
#316370000000
0#
0(
#316380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#316430000000
0$
0)
#316440000000
1"
1'
b0 +
b0 1
#316490000000
0"
0'
#316500000000
1#
1(
b101111101100100 +
b101111101100100 1
#316550000000
0#
0(
#316560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#316610000000
0$
0)
#316620000000
1"
1'
b0 +
b0 1
#316670000000
0"
0'
#316680000000
1#
1(
b101111101100100 +
b101111101100100 1
#316730000000
0#
0(
#316740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#316790000000
0$
0)
#316800000000
1"
1'
b0 +
b0 1
#316850000000
0"
0'
#316860000000
1#
1(
b101111101100100 +
b101111101100100 1
#316910000000
0#
0(
#316920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#316970000000
0$
0)
#316980000000
1"
1'
b0 +
b0 1
#317030000000
0"
0'
#317040000000
1#
1(
b101111101100100 +
b101111101100100 1
#317090000000
0#
0(
#317100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#317150000000
0$
0)
#317160000000
1"
1'
b0 +
b0 1
#317210000000
0"
0'
#317220000000
1#
1(
b101111101100100 +
b101111101100100 1
#317270000000
0#
0(
#317280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#317330000000
0$
0)
#317340000000
1"
1'
b0 +
b0 1
#317390000000
0"
0'
#317400000000
1#
1(
b101111101100100 +
b101111101100100 1
#317450000000
0#
0(
#317460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#317510000000
0$
0)
#317520000000
1"
1'
b0 +
b0 1
#317570000000
0"
0'
#317580000000
1#
1(
b101111101100100 +
b101111101100100 1
#317630000000
0#
0(
#317640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#317690000000
0$
0)
#317700000000
1"
1'
b0 +
b0 1
#317750000000
0"
0'
#317760000000
1#
1(
b101111101100100 +
b101111101100100 1
#317810000000
0#
0(
#317820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#317870000000
0$
0)
#317880000000
1"
1'
b0 +
b0 1
#317930000000
0"
0'
#317940000000
1#
1(
b101111101100100 +
b101111101100100 1
#317990000000
0#
0(
#318000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#318050000000
0$
0)
#318060000000
1"
1'
b0 +
b0 1
#318110000000
0"
0'
#318120000000
1#
1(
b101111101100100 +
b101111101100100 1
#318170000000
0#
0(
#318180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#318230000000
0$
0)
#318240000000
1"
1'
b0 +
b0 1
#318290000000
0"
0'
#318300000000
1#
1(
b101111101100100 +
b101111101100100 1
#318350000000
0#
0(
#318360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#318410000000
0$
0)
#318420000000
1"
1'
b0 +
b0 1
#318470000000
0"
0'
#318480000000
1#
1(
b101111101100100 +
b101111101100100 1
#318530000000
0#
0(
#318540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#318590000000
0$
0)
#318600000000
1"
1'
b0 +
b0 1
#318650000000
0"
0'
#318660000000
1#
1(
b101111101100100 +
b101111101100100 1
#318710000000
0#
0(
#318720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#318770000000
0$
0)
#318780000000
1"
1'
b0 +
b0 1
#318830000000
0"
0'
#318840000000
1#
1(
b101111101100100 +
b101111101100100 1
#318890000000
0#
0(
#318900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#318950000000
0$
0)
#318960000000
1"
1'
b0 +
b0 1
#319010000000
0"
0'
#319020000000
1#
1(
b101111101100100 +
b101111101100100 1
#319070000000
0#
0(
#319080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#319130000000
0$
0)
#319140000000
1"
1'
b0 +
b0 1
#319190000000
0"
0'
#319200000000
1#
1(
b101111101100100 +
b101111101100100 1
#319250000000
0#
0(
#319260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#319310000000
0$
0)
#319320000000
1"
1'
b0 +
b0 1
#319370000000
0"
0'
#319380000000
1#
1(
b101111101100100 +
b101111101100100 1
#319430000000
0#
0(
#319440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#319490000000
0$
0)
#319500000000
1"
1'
b0 +
b0 1
#319550000000
0"
0'
#319560000000
1#
1(
b101111101100100 +
b101111101100100 1
#319610000000
0#
0(
#319620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#319670000000
0$
0)
#319680000000
1"
1'
b0 +
b0 1
#319730000000
0"
0'
#319740000000
1#
1(
b101111101100100 +
b101111101100100 1
#319790000000
0#
0(
#319800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#319850000000
0$
0)
#319860000000
1"
1'
b0 +
b0 1
#319910000000
0"
0'
#319920000000
1#
1(
b101111101100100 +
b101111101100100 1
#319970000000
0#
0(
#319980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#320030000000
0$
0)
#320040000000
1"
1'
b0 +
b0 1
#320090000000
0"
0'
#320100000000
1#
1(
b101111101100100 +
b101111101100100 1
#320150000000
0#
0(
#320160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#320210000000
0$
0)
#320220000000
1"
1'
b0 +
b0 1
#320270000000
0"
0'
#320280000000
1#
1(
b101111101100100 +
b101111101100100 1
#320330000000
0#
0(
#320340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#320390000000
0$
0)
#320400000000
1"
1'
b0 +
b0 1
#320450000000
0"
0'
#320460000000
1#
1(
b101111101100100 +
b101111101100100 1
#320510000000
0#
0(
#320520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#320570000000
0$
0)
#320580000000
1"
1'
b0 +
b0 1
#320630000000
0"
0'
#320640000000
1#
1(
b101111101100100 +
b101111101100100 1
#320690000000
0#
0(
#320700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#320750000000
0$
0)
#320760000000
1"
1'
b0 +
b0 1
#320810000000
0"
0'
#320820000000
1#
1(
b101111101100100 +
b101111101100100 1
#320870000000
0#
0(
#320880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#320930000000
0$
0)
#320940000000
1"
1'
b0 +
b0 1
#320990000000
0"
0'
#321000000000
1#
1(
b101111101100100 +
b101111101100100 1
#321050000000
0#
0(
#321060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#321110000000
0$
0)
#321120000000
1"
1'
b0 +
b0 1
#321170000000
0"
0'
#321180000000
1#
1(
b101111101100100 +
b101111101100100 1
#321230000000
0#
0(
#321240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#321290000000
0$
0)
#321300000000
1"
1'
b0 +
b0 1
#321350000000
0"
0'
#321360000000
1#
1(
b101111101100100 +
b101111101100100 1
#321410000000
0#
0(
#321420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#321470000000
0$
0)
#321480000000
1"
1'
b0 +
b0 1
#321530000000
0"
0'
#321540000000
1#
1(
b101111101100100 +
b101111101100100 1
#321590000000
0#
0(
#321600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#321650000000
0$
0)
#321660000000
1"
1'
b0 +
b0 1
#321710000000
0"
0'
#321720000000
1#
1(
b101111101100100 +
b101111101100100 1
#321770000000
0#
0(
#321780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#321830000000
0$
0)
#321840000000
1"
1'
b0 +
b0 1
#321890000000
0"
0'
#321900000000
1#
1(
b101111101100100 +
b101111101100100 1
#321950000000
0#
0(
#321960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#322010000000
0$
0)
#322020000000
1"
1'
b0 +
b0 1
#322070000000
0"
0'
#322080000000
1#
1(
b101111101100100 +
b101111101100100 1
#322130000000
0#
0(
#322140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#322190000000
0$
0)
#322200000000
1"
1'
b0 +
b0 1
#322250000000
0"
0'
#322260000000
1#
1(
b101111101100100 +
b101111101100100 1
#322310000000
0#
0(
#322320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#322370000000
0$
0)
#322380000000
1"
1'
b0 +
b0 1
#322430000000
0"
0'
#322440000000
1#
1(
b101111101100100 +
b101111101100100 1
#322490000000
0#
0(
#322500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#322550000000
0$
0)
#322560000000
1"
1'
b0 +
b0 1
#322610000000
0"
0'
#322620000000
1#
1(
b101111101100100 +
b101111101100100 1
#322670000000
0#
0(
#322680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#322730000000
0$
0)
#322740000000
1"
1'
b0 +
b0 1
#322790000000
0"
0'
#322800000000
1#
1(
b101111101100100 +
b101111101100100 1
#322850000000
0#
0(
#322860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#322910000000
0$
0)
#322920000000
1"
1'
b0 +
b0 1
#322970000000
0"
0'
#322980000000
1#
1(
b101111101100100 +
b101111101100100 1
#323030000000
0#
0(
#323040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#323090000000
0$
0)
#323100000000
1"
1'
b0 +
b0 1
#323150000000
0"
0'
#323160000000
1#
1(
b101111101100100 +
b101111101100100 1
#323210000000
0#
0(
#323220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#323270000000
0$
0)
#323280000000
1"
1'
b0 +
b0 1
#323330000000
0"
0'
#323340000000
1#
1(
b101111101100100 +
b101111101100100 1
#323390000000
0#
0(
#323400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#323450000000
0$
0)
#323460000000
1"
1'
b0 +
b0 1
#323510000000
0"
0'
#323520000000
1#
1(
b101111101100100 +
b101111101100100 1
#323570000000
0#
0(
#323580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#323630000000
0$
0)
#323640000000
1"
1'
b0 +
b0 1
#323690000000
0"
0'
#323700000000
1#
1(
b101111101100100 +
b101111101100100 1
#323750000000
0#
0(
#323760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#323810000000
0$
0)
#323820000000
1"
1'
b0 +
b0 1
#323870000000
0"
0'
#323880000000
1#
1(
b101111101100100 +
b101111101100100 1
#323930000000
0#
0(
#323940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#323990000000
0$
0)
#324000000000
1"
1'
b0 +
b0 1
#324050000000
0"
0'
#324060000000
1#
1(
b101111101100100 +
b101111101100100 1
#324110000000
0#
0(
#324120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#324170000000
0$
0)
#324180000000
1"
1'
b0 +
b0 1
#324230000000
0"
0'
#324240000000
1#
1(
b101111101100100 +
b101111101100100 1
#324290000000
0#
0(
#324300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#324350000000
0$
0)
#324360000000
1"
1'
b0 +
b0 1
#324410000000
0"
0'
#324420000000
1#
1(
b101111101100100 +
b101111101100100 1
#324470000000
0#
0(
#324480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#324530000000
0$
0)
#324540000000
1"
1'
b0 +
b0 1
#324590000000
0"
0'
#324600000000
1#
1(
b101111101100100 +
b101111101100100 1
#324650000000
0#
0(
#324660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#324710000000
0$
0)
#324720000000
1"
1'
b0 +
b0 1
#324770000000
0"
0'
#324780000000
1#
1(
b101111101100100 +
b101111101100100 1
#324830000000
0#
0(
#324840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#324890000000
0$
0)
#324900000000
1"
1'
b0 +
b0 1
#324950000000
0"
0'
#324960000000
1#
1(
b101111101100100 +
b101111101100100 1
#325010000000
0#
0(
#325020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#325070000000
0$
0)
#325080000000
1"
1'
b0 +
b0 1
#325130000000
0"
0'
#325140000000
1#
1(
b101111101100100 +
b101111101100100 1
#325190000000
0#
0(
#325200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#325250000000
0$
0)
#325260000000
1"
1'
b0 +
b0 1
#325310000000
0"
0'
#325320000000
1#
1(
b101111101100100 +
b101111101100100 1
#325370000000
0#
0(
#325380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#325430000000
0$
0)
#325440000000
1"
1'
b0 +
b0 1
#325490000000
0"
0'
#325500000000
1#
1(
b101111101100100 +
b101111101100100 1
#325550000000
0#
0(
#325560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#325610000000
0$
0)
#325620000000
1"
1'
b0 +
b0 1
#325670000000
0"
0'
#325680000000
1#
1(
b101111101100100 +
b101111101100100 1
#325730000000
0#
0(
#325740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#325790000000
0$
0)
#325800000000
1"
1'
b0 +
b0 1
#325850000000
0"
0'
#325860000000
1#
1(
b101111101100100 +
b101111101100100 1
#325910000000
0#
0(
#325920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#325970000000
0$
0)
#325980000000
1"
1'
b0 +
b0 1
#326030000000
0"
0'
#326040000000
1#
1(
b101111101100100 +
b101111101100100 1
#326090000000
0#
0(
#326100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#326150000000
0$
0)
#326160000000
1"
1'
b0 +
b0 1
#326210000000
0"
0'
#326220000000
1#
1(
b101111101100100 +
b101111101100100 1
#326270000000
0#
0(
#326280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#326330000000
0$
0)
#326340000000
1"
1'
b0 +
b0 1
#326390000000
0"
0'
#326400000000
1#
1(
b101111101100100 +
b101111101100100 1
#326450000000
0#
0(
#326460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#326510000000
0$
0)
#326520000000
1"
1'
b0 +
b0 1
#326570000000
0"
0'
#326580000000
1#
1(
b101111101100100 +
b101111101100100 1
#326630000000
0#
0(
#326640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#326690000000
0$
0)
#326700000000
1"
1'
b0 +
b0 1
#326750000000
0"
0'
#326760000000
1#
1(
b101111101100100 +
b101111101100100 1
#326810000000
0#
0(
#326820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#326870000000
0$
0)
#326880000000
1"
1'
b0 +
b0 1
#326930000000
0"
0'
#326940000000
1#
1(
b101111101100100 +
b101111101100100 1
#326990000000
0#
0(
#327000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#327050000000
0$
0)
#327060000000
1"
1'
b0 +
b0 1
#327110000000
0"
0'
#327120000000
1#
1(
b101111101100100 +
b101111101100100 1
#327170000000
0#
0(
#327180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#327230000000
0$
0)
#327240000000
1"
1'
b0 +
b0 1
#327290000000
0"
0'
#327300000000
1#
1(
b101111101100100 +
b101111101100100 1
#327350000000
0#
0(
#327360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#327410000000
0$
0)
#327420000000
1"
1'
b0 +
b0 1
#327470000000
0"
0'
#327480000000
1#
1(
b101111101100100 +
b101111101100100 1
#327530000000
0#
0(
#327540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#327590000000
0$
0)
#327600000000
1"
1'
b0 +
b0 1
#327650000000
0"
0'
#327660000000
1#
1(
b101111101100100 +
b101111101100100 1
#327710000000
0#
0(
#327720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#327770000000
0$
0)
#327780000000
1"
1'
b0 +
b0 1
#327830000000
0"
0'
#327840000000
1#
1(
b101111101100100 +
b101111101100100 1
#327890000000
0#
0(
#327900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#327950000000
0$
0)
#327960000000
1"
1'
b0 +
b0 1
#328010000000
0"
0'
#328020000000
1#
1(
b101111101100100 +
b101111101100100 1
#328070000000
0#
0(
#328080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#328130000000
0$
0)
#328140000000
1"
1'
b0 +
b0 1
#328190000000
0"
0'
#328200000000
1#
1(
b101111101100100 +
b101111101100100 1
#328250000000
0#
0(
#328260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#328310000000
0$
0)
#328320000000
1"
1'
b0 +
b0 1
#328370000000
0"
0'
#328380000000
1#
1(
b101111101100100 +
b101111101100100 1
#328430000000
0#
0(
#328440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#328490000000
0$
0)
#328500000000
1"
1'
b0 +
b0 1
#328550000000
0"
0'
#328560000000
1#
1(
b101111101100100 +
b101111101100100 1
#328610000000
0#
0(
#328620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#328670000000
0$
0)
#328680000000
1"
1'
b0 +
b0 1
#328730000000
0"
0'
#328740000000
1#
1(
b101111101100100 +
b101111101100100 1
#328790000000
0#
0(
#328800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#328850000000
0$
0)
#328860000000
1"
1'
b0 +
b0 1
#328910000000
0"
0'
#328920000000
1#
1(
b101111101100100 +
b101111101100100 1
#328970000000
0#
0(
#328980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#329030000000
0$
0)
#329040000000
1"
1'
b0 +
b0 1
#329090000000
0"
0'
#329100000000
1#
1(
b101111101100100 +
b101111101100100 1
#329150000000
0#
0(
#329160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#329210000000
0$
0)
#329220000000
1"
1'
b0 +
b0 1
#329270000000
0"
0'
#329280000000
1#
1(
b101111101100100 +
b101111101100100 1
#329330000000
0#
0(
#329340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#329390000000
0$
0)
#329400000000
1"
1'
b0 +
b0 1
#329450000000
0"
0'
#329460000000
1#
1(
b101111101100100 +
b101111101100100 1
#329510000000
0#
0(
#329520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#329570000000
0$
0)
#329580000000
1"
1'
b0 +
b0 1
#329630000000
0"
0'
#329640000000
1#
1(
b101111101100100 +
b101111101100100 1
#329690000000
0#
0(
#329700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#329750000000
0$
0)
#329760000000
1"
1'
b0 +
b0 1
#329810000000
0"
0'
#329820000000
1#
1(
b101111101100100 +
b101111101100100 1
#329870000000
0#
0(
#329880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#329930000000
0$
0)
#329940000000
1"
1'
b0 +
b0 1
#329990000000
0"
0'
#330000000000
1#
1(
b101111101100100 +
b101111101100100 1
#330050000000
0#
0(
#330060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#330110000000
0$
0)
#330120000000
1"
1'
b0 +
b0 1
#330170000000
0"
0'
#330180000000
1#
1(
b101111101100100 +
b101111101100100 1
#330230000000
0#
0(
#330240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#330290000000
0$
0)
#330300000000
1"
1'
b0 +
b0 1
#330350000000
0"
0'
#330360000000
1#
1(
b101111101100100 +
b101111101100100 1
#330410000000
0#
0(
#330420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#330470000000
0$
0)
#330480000000
1"
1'
b0 +
b0 1
#330530000000
0"
0'
#330540000000
1#
1(
b101111101100100 +
b101111101100100 1
#330590000000
0#
0(
#330600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#330650000000
0$
0)
#330660000000
1"
1'
b0 +
b0 1
#330710000000
0"
0'
#330720000000
1#
1(
b101111101100100 +
b101111101100100 1
#330770000000
0#
0(
#330780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#330830000000
0$
0)
#330840000000
1"
1'
b0 +
b0 1
#330890000000
0"
0'
#330900000000
1#
1(
b101111101100100 +
b101111101100100 1
#330950000000
0#
0(
#330960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#331010000000
0$
0)
#331020000000
1"
1'
b0 +
b0 1
#331070000000
0"
0'
#331080000000
1#
1(
b101111101100100 +
b101111101100100 1
#331130000000
0#
0(
#331140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#331190000000
0$
0)
#331200000000
1"
1'
b0 +
b0 1
#331250000000
0"
0'
#331260000000
1#
1(
b101111101100100 +
b101111101100100 1
#331310000000
0#
0(
#331320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#331370000000
0$
0)
#331380000000
1"
1'
b0 +
b0 1
#331430000000
0"
0'
#331440000000
1#
1(
b101111101100100 +
b101111101100100 1
#331490000000
0#
0(
#331500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#331550000000
0$
0)
#331560000000
1"
1'
b0 +
b0 1
#331610000000
0"
0'
#331620000000
1#
1(
b101111101100100 +
b101111101100100 1
#331670000000
0#
0(
#331680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#331730000000
0$
0)
#331740000000
1"
1'
b0 +
b0 1
#331790000000
0"
0'
#331800000000
1#
1(
b101111101100100 +
b101111101100100 1
#331850000000
0#
0(
#331860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#331910000000
0$
0)
#331920000000
1"
1'
b0 +
b0 1
#331970000000
0"
0'
#331980000000
1#
1(
b101111101100100 +
b101111101100100 1
#332030000000
0#
0(
#332040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#332090000000
0$
0)
#332100000000
1"
1'
b0 +
b0 1
#332150000000
0"
0'
#332160000000
1#
1(
b101111101100100 +
b101111101100100 1
#332210000000
0#
0(
#332220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#332270000000
0$
0)
#332280000000
1"
1'
b0 +
b0 1
#332330000000
0"
0'
#332340000000
1#
1(
b101111101100100 +
b101111101100100 1
#332390000000
0#
0(
#332400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#332450000000
0$
0)
#332460000000
1"
1'
b0 +
b0 1
#332510000000
0"
0'
#332520000000
1#
1(
b101111101100100 +
b101111101100100 1
#332570000000
0#
0(
#332580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#332630000000
0$
0)
#332640000000
1"
1'
b0 +
b0 1
#332690000000
0"
0'
#332700000000
1#
1(
b101111101100100 +
b101111101100100 1
#332750000000
0#
0(
#332760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#332810000000
0$
0)
#332820000000
1"
1'
b0 +
b0 1
#332870000000
0"
0'
#332880000000
1#
1(
b101111101100100 +
b101111101100100 1
#332930000000
0#
0(
#332940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#332990000000
0$
0)
#333000000000
1"
1'
b0 +
b0 1
#333050000000
0"
0'
#333060000000
1#
1(
b101111101100100 +
b101111101100100 1
#333110000000
0#
0(
#333120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#333170000000
0$
0)
#333180000000
1"
1'
b0 +
b0 1
#333230000000
0"
0'
#333240000000
1#
1(
b101111101100100 +
b101111101100100 1
#333290000000
0#
0(
#333300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#333350000000
0$
0)
#333360000000
1"
1'
b0 +
b0 1
#333410000000
0"
0'
#333420000000
1#
1(
b101111101100100 +
b101111101100100 1
#333470000000
0#
0(
#333480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#333530000000
0$
0)
#333540000000
1"
1'
b0 +
b0 1
#333590000000
0"
0'
#333600000000
1#
1(
b101111101100100 +
b101111101100100 1
#333650000000
0#
0(
#333660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#333710000000
0$
0)
#333720000000
1"
1'
b0 +
b0 1
#333770000000
0"
0'
#333780000000
1#
1(
b101111101100100 +
b101111101100100 1
#333830000000
0#
0(
#333840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#333890000000
0$
0)
#333900000000
1"
1'
b0 +
b0 1
#333950000000
0"
0'
#333960000000
1#
1(
b101111101100100 +
b101111101100100 1
#334010000000
0#
0(
#334020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#334070000000
0$
0)
#334080000000
1"
1'
b0 +
b0 1
#334130000000
0"
0'
#334140000000
1#
1(
b101111101100100 +
b101111101100100 1
#334190000000
0#
0(
#334200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#334250000000
0$
0)
#334260000000
1"
1'
b0 +
b0 1
#334310000000
0"
0'
#334320000000
1#
1(
b101111101100100 +
b101111101100100 1
#334370000000
0#
0(
#334380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#334430000000
0$
0)
#334440000000
1"
1'
b0 +
b0 1
#334490000000
0"
0'
#334500000000
1#
1(
b101111101100100 +
b101111101100100 1
#334550000000
0#
0(
#334560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#334610000000
0$
0)
#334620000000
1"
1'
b0 +
b0 1
#334670000000
0"
0'
#334680000000
1#
1(
b101111101100100 +
b101111101100100 1
#334730000000
0#
0(
#334740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#334790000000
0$
0)
#334800000000
1"
1'
b0 +
b0 1
#334850000000
0"
0'
#334860000000
1#
1(
b101111101100100 +
b101111101100100 1
#334910000000
0#
0(
#334920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#334970000000
0$
0)
#334980000000
1"
1'
b0 +
b0 1
#335030000000
0"
0'
#335040000000
1#
1(
b101111101100100 +
b101111101100100 1
#335090000000
0#
0(
#335100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#335150000000
0$
0)
#335160000000
1"
1'
b0 +
b0 1
#335210000000
0"
0'
#335220000000
1#
1(
b101111101100100 +
b101111101100100 1
#335270000000
0#
0(
#335280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#335330000000
0$
0)
#335340000000
1"
1'
b0 +
b0 1
#335390000000
0"
0'
#335400000000
1#
1(
b101111101100100 +
b101111101100100 1
#335450000000
0#
0(
#335460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#335510000000
0$
0)
#335520000000
1"
1'
b0 +
b0 1
#335570000000
0"
0'
#335580000000
1#
1(
b101111101100100 +
b101111101100100 1
#335630000000
0#
0(
#335640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#335690000000
0$
0)
#335700000000
1"
1'
b0 +
b0 1
#335750000000
0"
0'
#335760000000
1#
1(
b101111101100100 +
b101111101100100 1
#335810000000
0#
0(
#335820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#335870000000
0$
0)
#335880000000
1"
1'
b0 +
b0 1
#335930000000
0"
0'
#335940000000
1#
1(
b101111101100100 +
b101111101100100 1
#335990000000
0#
0(
#336000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#336050000000
0$
0)
#336060000000
1"
1'
b0 +
b0 1
#336110000000
0"
0'
#336120000000
1#
1(
b101111101100100 +
b101111101100100 1
#336170000000
0#
0(
#336180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#336230000000
0$
0)
#336240000000
1"
1'
b0 +
b0 1
#336290000000
0"
0'
#336300000000
1#
1(
b101111101100100 +
b101111101100100 1
#336350000000
0#
0(
#336360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#336410000000
0$
0)
#336420000000
1"
1'
b0 +
b0 1
#336470000000
0"
0'
#336480000000
1#
1(
b101111101100100 +
b101111101100100 1
#336530000000
0#
0(
#336540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#336590000000
0$
0)
#336600000000
1"
1'
b0 +
b0 1
#336650000000
0"
0'
#336660000000
1#
1(
b101111101100100 +
b101111101100100 1
#336710000000
0#
0(
#336720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#336770000000
0$
0)
#336780000000
1"
1'
b0 +
b0 1
#336830000000
0"
0'
#336840000000
1#
1(
b101111101100100 +
b101111101100100 1
#336890000000
0#
0(
#336900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#336950000000
0$
0)
#336960000000
1"
1'
b0 +
b0 1
#337010000000
0"
0'
#337020000000
1#
1(
b101111101100100 +
b101111101100100 1
#337070000000
0#
0(
#337080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#337130000000
0$
0)
#337140000000
1"
1'
b0 +
b0 1
#337190000000
0"
0'
#337200000000
1#
1(
b101111101100100 +
b101111101100100 1
#337250000000
0#
0(
#337260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#337310000000
0$
0)
#337320000000
1"
1'
b0 +
b0 1
#337370000000
0"
0'
#337380000000
1#
1(
b101111101100100 +
b101111101100100 1
#337430000000
0#
0(
#337440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#337490000000
0$
0)
#337500000000
1"
1'
b0 +
b0 1
#337550000000
0"
0'
#337560000000
1#
1(
b101111101100100 +
b101111101100100 1
#337610000000
0#
0(
#337620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#337670000000
0$
0)
#337680000000
1"
1'
b0 +
b0 1
#337730000000
0"
0'
#337740000000
1#
1(
b101111101100100 +
b101111101100100 1
#337790000000
0#
0(
#337800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#337850000000
0$
0)
#337860000000
1"
1'
b0 +
b0 1
#337910000000
0"
0'
#337920000000
1#
1(
b101111101100100 +
b101111101100100 1
#337970000000
0#
0(
#337980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#338030000000
0$
0)
#338040000000
1"
1'
b0 +
b0 1
#338090000000
0"
0'
#338100000000
1#
1(
b101111101100100 +
b101111101100100 1
#338150000000
0#
0(
#338160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#338210000000
0$
0)
#338220000000
1"
1'
b0 +
b0 1
#338270000000
0"
0'
#338280000000
1#
1(
b101111101100100 +
b101111101100100 1
#338330000000
0#
0(
#338340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#338390000000
0$
0)
#338400000000
1"
1'
b0 +
b0 1
#338450000000
0"
0'
#338460000000
1#
1(
b101111101100100 +
b101111101100100 1
#338510000000
0#
0(
#338520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#338570000000
0$
0)
#338580000000
1"
1'
b0 +
b0 1
#338630000000
0"
0'
#338640000000
1#
1(
b101111101100100 +
b101111101100100 1
#338690000000
0#
0(
#338700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#338750000000
0$
0)
#338760000000
1"
1'
b0 +
b0 1
#338810000000
0"
0'
#338820000000
1#
1(
b101111101100100 +
b101111101100100 1
#338870000000
0#
0(
#338880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#338930000000
0$
0)
#338940000000
1"
1'
b0 +
b0 1
#338990000000
0"
0'
#339000000000
1#
1(
b101111101100100 +
b101111101100100 1
#339050000000
0#
0(
#339060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#339110000000
0$
0)
#339120000000
1"
1'
b0 +
b0 1
#339170000000
0"
0'
#339180000000
1#
1(
b101111101100100 +
b101111101100100 1
#339230000000
0#
0(
#339240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#339290000000
0$
0)
#339300000000
1"
1'
b0 +
b0 1
#339350000000
0"
0'
#339360000000
1#
1(
b101111101100100 +
b101111101100100 1
#339410000000
0#
0(
#339420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#339470000000
0$
0)
#339480000000
1"
1'
b0 +
b0 1
#339530000000
0"
0'
#339540000000
1#
1(
b101111101100100 +
b101111101100100 1
#339590000000
0#
0(
#339600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#339650000000
0$
0)
#339660000000
1"
1'
b0 +
b0 1
#339710000000
0"
0'
#339720000000
1#
1(
b101111101100100 +
b101111101100100 1
#339770000000
0#
0(
#339780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#339830000000
0$
0)
#339840000000
1"
1'
b0 +
b0 1
#339890000000
0"
0'
#339900000000
1#
1(
b101111101100100 +
b101111101100100 1
#339950000000
0#
0(
#339960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#340010000000
0$
0)
#340020000000
1"
1'
b0 +
b0 1
#340070000000
0"
0'
#340080000000
1#
1(
b101111101100100 +
b101111101100100 1
#340130000000
0#
0(
#340140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#340190000000
0$
0)
#340200000000
1"
1'
b0 +
b0 1
#340250000000
0"
0'
#340260000000
1#
1(
b101111101100100 +
b101111101100100 1
#340310000000
0#
0(
#340320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#340370000000
0$
0)
#340380000000
1"
1'
b0 +
b0 1
#340430000000
0"
0'
#340440000000
1#
1(
b101111101100100 +
b101111101100100 1
#340490000000
0#
0(
#340500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#340550000000
0$
0)
#340560000000
1"
1'
b0 +
b0 1
#340610000000
0"
0'
#340620000000
1#
1(
b101111101100100 +
b101111101100100 1
#340670000000
0#
0(
#340680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#340730000000
0$
0)
#340740000000
1"
1'
b0 +
b0 1
#340790000000
0"
0'
#340800000000
1#
1(
b101111101100100 +
b101111101100100 1
#340850000000
0#
0(
#340860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#340910000000
0$
0)
#340920000000
1"
1'
b0 +
b0 1
#340970000000
0"
0'
#340980000000
1#
1(
b101111101100100 +
b101111101100100 1
#341030000000
0#
0(
#341040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#341090000000
0$
0)
#341100000000
1"
1'
b0 +
b0 1
#341150000000
0"
0'
#341160000000
1#
1(
b101111101100100 +
b101111101100100 1
#341210000000
0#
0(
#341220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#341270000000
0$
0)
#341280000000
1"
1'
b0 +
b0 1
#341330000000
0"
0'
#341340000000
1#
1(
b101111101100100 +
b101111101100100 1
#341390000000
0#
0(
#341400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#341450000000
0$
0)
#341460000000
1"
1'
b0 +
b0 1
#341510000000
0"
0'
#341520000000
1#
1(
b101111101100100 +
b101111101100100 1
#341570000000
0#
0(
#341580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#341630000000
0$
0)
#341640000000
1"
1'
b0 +
b0 1
#341690000000
0"
0'
#341700000000
1#
1(
b101111101100100 +
b101111101100100 1
#341750000000
0#
0(
#341760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#341810000000
0$
0)
#341820000000
1"
1'
b0 +
b0 1
#341870000000
0"
0'
#341880000000
1#
1(
b101111101100100 +
b101111101100100 1
#341930000000
0#
0(
#341940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#341990000000
0$
0)
#342000000000
1"
1'
b0 +
b0 1
#342050000000
0"
0'
#342060000000
1#
1(
b101111101100100 +
b101111101100100 1
#342110000000
0#
0(
#342120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#342170000000
0$
0)
#342180000000
1"
1'
b0 +
b0 1
#342230000000
0"
0'
#342240000000
1#
1(
b101111101100100 +
b101111101100100 1
#342290000000
0#
0(
#342300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#342350000000
0$
0)
#342360000000
1"
1'
b0 +
b0 1
#342410000000
0"
0'
#342420000000
1#
1(
b101111101100100 +
b101111101100100 1
#342470000000
0#
0(
#342480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#342530000000
0$
0)
#342540000000
1"
1'
b0 +
b0 1
#342590000000
0"
0'
#342600000000
1#
1(
b101111101100100 +
b101111101100100 1
#342650000000
0#
0(
#342660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#342710000000
0$
0)
#342720000000
1"
1'
b0 +
b0 1
#342770000000
0"
0'
#342780000000
1#
1(
b101111101100100 +
b101111101100100 1
#342830000000
0#
0(
#342840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#342890000000
0$
0)
#342900000000
1"
1'
b0 +
b0 1
#342950000000
0"
0'
#342960000000
1#
1(
b101111101100100 +
b101111101100100 1
#343010000000
0#
0(
#343020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#343070000000
0$
0)
#343080000000
1"
1'
b0 +
b0 1
#343130000000
0"
0'
#343140000000
1#
1(
b101111101100100 +
b101111101100100 1
#343190000000
0#
0(
#343200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#343250000000
0$
0)
#343260000000
1"
1'
b0 +
b0 1
#343310000000
0"
0'
#343320000000
1#
1(
b101111101100100 +
b101111101100100 1
#343370000000
0#
0(
#343380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#343430000000
0$
0)
#343440000000
1"
1'
b0 +
b0 1
#343490000000
0"
0'
#343500000000
1#
1(
b101111101100100 +
b101111101100100 1
#343550000000
0#
0(
#343560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#343610000000
0$
0)
#343620000000
1"
1'
b0 +
b0 1
#343670000000
0"
0'
#343680000000
1#
1(
b101111101100100 +
b101111101100100 1
#343730000000
0#
0(
#343740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#343790000000
0$
0)
#343800000000
1"
1'
b0 +
b0 1
#343850000000
0"
0'
#343860000000
1#
1(
b101111101100100 +
b101111101100100 1
#343910000000
0#
0(
#343920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#343970000000
0$
0)
#343980000000
1"
1'
b0 +
b0 1
#344030000000
0"
0'
#344040000000
1#
1(
b101111101100100 +
b101111101100100 1
#344090000000
0#
0(
#344100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#344150000000
0$
0)
#344160000000
1"
1'
b0 +
b0 1
#344210000000
0"
0'
#344220000000
1#
1(
b101111101100100 +
b101111101100100 1
#344270000000
0#
0(
#344280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#344330000000
0$
0)
#344340000000
1"
1'
b0 +
b0 1
#344390000000
0"
0'
#344400000000
1#
1(
b101111101100100 +
b101111101100100 1
#344450000000
0#
0(
#344460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#344510000000
0$
0)
#344520000000
1"
1'
b0 +
b0 1
#344570000000
0"
0'
#344580000000
1#
1(
b101111101100100 +
b101111101100100 1
#344630000000
0#
0(
#344640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#344690000000
0$
0)
#344700000000
1"
1'
b0 +
b0 1
#344750000000
0"
0'
#344760000000
1#
1(
b101111101100100 +
b101111101100100 1
#344810000000
0#
0(
#344820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#344870000000
0$
0)
#344880000000
1"
1'
b0 +
b0 1
#344930000000
0"
0'
#344940000000
1#
1(
b101111101100100 +
b101111101100100 1
#344990000000
0#
0(
#345000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#345050000000
0$
0)
#345060000000
1"
1'
b0 +
b0 1
#345110000000
0"
0'
#345120000000
1#
1(
b101111101100100 +
b101111101100100 1
#345170000000
0#
0(
#345180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#345230000000
0$
0)
#345240000000
1"
1'
b0 +
b0 1
#345290000000
0"
0'
#345300000000
1#
1(
b101111101100100 +
b101111101100100 1
#345350000000
0#
0(
#345360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#345410000000
0$
0)
#345420000000
1"
1'
b0 +
b0 1
#345470000000
0"
0'
#345480000000
1#
1(
b101111101100100 +
b101111101100100 1
#345530000000
0#
0(
#345540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#345590000000
0$
0)
#345600000000
1"
1'
b0 +
b0 1
#345650000000
0"
0'
#345660000000
1#
1(
b101111101100100 +
b101111101100100 1
#345710000000
0#
0(
#345720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#345770000000
0$
0)
#345780000000
1"
1'
b0 +
b0 1
#345830000000
0"
0'
#345840000000
1#
1(
b101111101100100 +
b101111101100100 1
#345890000000
0#
0(
#345900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#345950000000
0$
0)
#345960000000
1"
1'
b0 +
b0 1
#346010000000
0"
0'
#346020000000
1#
1(
b101111101100100 +
b101111101100100 1
#346070000000
0#
0(
#346080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#346130000000
0$
0)
#346140000000
1"
1'
b0 +
b0 1
#346190000000
0"
0'
#346200000000
1#
1(
b101111101100100 +
b101111101100100 1
#346250000000
0#
0(
#346260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#346310000000
0$
0)
#346320000000
1"
1'
b0 +
b0 1
#346370000000
0"
0'
#346380000000
1#
1(
b101111101100100 +
b101111101100100 1
#346430000000
0#
0(
#346440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#346490000000
0$
0)
#346500000000
1"
1'
b0 +
b0 1
#346550000000
0"
0'
#346560000000
1#
1(
b101111101100100 +
b101111101100100 1
#346610000000
0#
0(
#346620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#346670000000
0$
0)
#346680000000
1"
1'
b0 +
b0 1
#346730000000
0"
0'
#346740000000
1#
1(
b101111101100100 +
b101111101100100 1
#346790000000
0#
0(
#346800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#346850000000
0$
0)
#346860000000
1"
1'
b0 +
b0 1
#346910000000
0"
0'
#346920000000
1#
1(
b101111101100100 +
b101111101100100 1
#346970000000
0#
0(
#346980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#347030000000
0$
0)
#347040000000
1"
1'
b0 +
b0 1
#347090000000
0"
0'
#347100000000
1#
1(
b101111101100100 +
b101111101100100 1
#347150000000
0#
0(
#347160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#347210000000
0$
0)
#347220000000
1"
1'
b0 +
b0 1
#347270000000
0"
0'
#347280000000
1#
1(
b101111101100100 +
b101111101100100 1
#347330000000
0#
0(
#347340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#347390000000
0$
0)
#347400000000
1"
1'
b0 +
b0 1
#347450000000
0"
0'
#347460000000
1#
1(
b101111101100100 +
b101111101100100 1
#347510000000
0#
0(
#347520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#347570000000
0$
0)
#347580000000
1"
1'
b0 +
b0 1
#347630000000
0"
0'
#347640000000
1#
1(
b101111101100100 +
b101111101100100 1
#347690000000
0#
0(
#347700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#347750000000
0$
0)
#347760000000
1"
1'
b0 +
b0 1
#347810000000
0"
0'
#347820000000
1#
1(
b101111101100100 +
b101111101100100 1
#347870000000
0#
0(
#347880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#347930000000
0$
0)
#347940000000
1"
1'
b0 +
b0 1
#347990000000
0"
0'
#348000000000
1#
1(
b101111101100100 +
b101111101100100 1
#348050000000
0#
0(
#348060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#348110000000
0$
0)
#348120000000
1"
1'
b0 +
b0 1
#348170000000
0"
0'
#348180000000
1#
1(
b101111101100100 +
b101111101100100 1
#348230000000
0#
0(
#348240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#348290000000
0$
0)
#348300000000
1"
1'
b0 +
b0 1
#348350000000
0"
0'
#348360000000
1#
1(
b101111101100100 +
b101111101100100 1
#348410000000
0#
0(
#348420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#348470000000
0$
0)
#348480000000
1"
1'
b0 +
b0 1
#348530000000
0"
0'
#348540000000
1#
1(
b101111101100100 +
b101111101100100 1
#348590000000
0#
0(
#348600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#348650000000
0$
0)
#348660000000
1"
1'
b0 +
b0 1
#348710000000
0"
0'
#348720000000
1#
1(
b101111101100100 +
b101111101100100 1
#348770000000
0#
0(
#348780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#348830000000
0$
0)
#348840000000
1"
1'
b0 +
b0 1
#348890000000
0"
0'
#348900000000
1#
1(
b101111101100100 +
b101111101100100 1
#348950000000
0#
0(
#348960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#349010000000
0$
0)
#349020000000
1"
1'
b0 +
b0 1
#349070000000
0"
0'
#349080000000
1#
1(
b101111101100100 +
b101111101100100 1
#349130000000
0#
0(
#349140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#349190000000
0$
0)
#349200000000
1"
1'
b0 +
b0 1
#349250000000
0"
0'
#349260000000
1#
1(
b101111101100100 +
b101111101100100 1
#349310000000
0#
0(
#349320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#349370000000
0$
0)
#349380000000
1"
1'
b0 +
b0 1
#349430000000
0"
0'
#349440000000
1#
1(
b101111101100100 +
b101111101100100 1
#349490000000
0#
0(
#349500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#349550000000
0$
0)
#349560000000
1"
1'
b0 +
b0 1
#349610000000
0"
0'
#349620000000
1#
1(
b101111101100100 +
b101111101100100 1
#349670000000
0#
0(
#349680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#349730000000
0$
0)
#349740000000
1"
1'
b0 +
b0 1
#349790000000
0"
0'
#349800000000
1#
1(
b101111101100100 +
b101111101100100 1
#349850000000
0#
0(
#349860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#349910000000
0$
0)
#349920000000
1"
1'
b0 +
b0 1
#349970000000
0"
0'
#349980000000
1#
1(
b101111101100100 +
b101111101100100 1
#350030000000
0#
0(
#350040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#350090000000
0$
0)
#350100000000
1"
1'
b0 +
b0 1
#350150000000
0"
0'
#350160000000
1#
1(
b101111101100100 +
b101111101100100 1
#350210000000
0#
0(
#350220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#350270000000
0$
0)
#350280000000
1"
1'
b0 +
b0 1
#350330000000
0"
0'
#350340000000
1#
1(
b101111101100100 +
b101111101100100 1
#350390000000
0#
0(
#350400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#350450000000
0$
0)
#350460000000
1"
1'
b0 +
b0 1
#350510000000
0"
0'
#350520000000
1#
1(
b101111101100100 +
b101111101100100 1
#350570000000
0#
0(
#350580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#350630000000
0$
0)
#350640000000
1"
1'
b0 +
b0 1
#350690000000
0"
0'
#350700000000
1#
1(
b101111101100100 +
b101111101100100 1
#350750000000
0#
0(
#350760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#350810000000
0$
0)
#350820000000
1"
1'
b0 +
b0 1
#350870000000
0"
0'
#350880000000
1#
1(
b101111101100100 +
b101111101100100 1
#350930000000
0#
0(
#350940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#350990000000
0$
0)
#351000000000
1"
1'
b0 +
b0 1
#351050000000
0"
0'
#351060000000
1#
1(
b101111101100100 +
b101111101100100 1
#351110000000
0#
0(
#351120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#351170000000
0$
0)
#351180000000
1"
1'
b0 +
b0 1
#351230000000
0"
0'
#351240000000
1#
1(
b101111101100100 +
b101111101100100 1
#351290000000
0#
0(
#351300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#351350000000
0$
0)
#351360000000
1"
1'
b0 +
b0 1
#351410000000
0"
0'
#351420000000
1#
1(
b101111101100100 +
b101111101100100 1
#351470000000
0#
0(
#351480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#351530000000
0$
0)
#351540000000
1"
1'
b0 +
b0 1
#351590000000
0"
0'
#351600000000
1#
1(
b101111101100100 +
b101111101100100 1
#351650000000
0#
0(
#351660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#351710000000
0$
0)
#351720000000
1"
1'
b0 +
b0 1
#351770000000
0"
0'
#351780000000
1#
1(
b101111101100100 +
b101111101100100 1
#351830000000
0#
0(
#351840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#351890000000
0$
0)
#351900000000
1"
1'
b0 +
b0 1
#351950000000
0"
0'
#351960000000
1#
1(
b101111101100100 +
b101111101100100 1
#352010000000
0#
0(
#352020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#352070000000
0$
0)
#352080000000
1"
1'
b0 +
b0 1
#352130000000
0"
0'
#352140000000
1#
1(
b101111101100100 +
b101111101100100 1
#352190000000
0#
0(
#352200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#352250000000
0$
0)
#352260000000
1"
1'
b0 +
b0 1
#352310000000
0"
0'
#352320000000
1#
1(
b101111101100100 +
b101111101100100 1
#352370000000
0#
0(
#352380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#352430000000
0$
0)
#352440000000
1"
1'
b0 +
b0 1
#352490000000
0"
0'
#352500000000
1#
1(
b101111101100100 +
b101111101100100 1
#352550000000
0#
0(
#352560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#352610000000
0$
0)
#352620000000
1"
1'
b0 +
b0 1
#352670000000
0"
0'
#352680000000
1#
1(
b101111101100100 +
b101111101100100 1
#352730000000
0#
0(
#352740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#352790000000
0$
0)
#352800000000
1"
1'
b0 +
b0 1
#352850000000
0"
0'
#352860000000
1#
1(
b101111101100100 +
b101111101100100 1
#352910000000
0#
0(
#352920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#352970000000
0$
0)
#352980000000
1"
1'
b0 +
b0 1
#353030000000
0"
0'
#353040000000
1#
1(
b101111101100100 +
b101111101100100 1
#353090000000
0#
0(
#353100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#353150000000
0$
0)
#353160000000
1"
1'
b0 +
b0 1
#353210000000
0"
0'
#353220000000
1#
1(
b101111101100100 +
b101111101100100 1
#353270000000
0#
0(
#353280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#353330000000
0$
0)
#353340000000
1"
1'
b0 +
b0 1
#353390000000
0"
0'
#353400000000
1#
1(
b101111101100100 +
b101111101100100 1
#353450000000
0#
0(
#353460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#353510000000
0$
0)
#353520000000
1"
1'
b0 +
b0 1
#353570000000
0"
0'
#353580000000
1#
1(
b101111101100100 +
b101111101100100 1
#353630000000
0#
0(
#353640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#353690000000
0$
0)
#353700000000
1"
1'
b0 +
b0 1
#353750000000
0"
0'
#353760000000
1#
1(
b101111101100100 +
b101111101100100 1
#353810000000
0#
0(
#353820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#353870000000
0$
0)
#353880000000
1"
1'
b0 +
b0 1
#353930000000
0"
0'
#353940000000
1#
1(
b101111101100100 +
b101111101100100 1
#353990000000
0#
0(
#354000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#354050000000
0$
0)
#354060000000
1"
1'
b0 +
b0 1
#354110000000
0"
0'
#354120000000
1#
1(
b101111101100100 +
b101111101100100 1
#354170000000
0#
0(
#354180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#354230000000
0$
0)
#354240000000
1"
1'
b0 +
b0 1
#354290000000
0"
0'
#354300000000
1#
1(
b101111101100100 +
b101111101100100 1
#354350000000
0#
0(
#354360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#354410000000
0$
0)
#354420000000
1"
1'
b0 +
b0 1
#354470000000
0"
0'
#354480000000
1#
1(
b101111101100100 +
b101111101100100 1
#354530000000
0#
0(
#354540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#354590000000
0$
0)
#354600000000
1"
1'
b0 +
b0 1
#354650000000
0"
0'
#354660000000
1#
1(
b101111101100100 +
b101111101100100 1
#354710000000
0#
0(
#354720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#354770000000
0$
0)
#354780000000
1"
1'
b0 +
b0 1
#354830000000
0"
0'
#354840000000
1#
1(
b101111101100100 +
b101111101100100 1
#354890000000
0#
0(
#354900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#354950000000
0$
0)
#354960000000
1"
1'
b0 +
b0 1
#355010000000
0"
0'
#355020000000
1#
1(
b101111101100100 +
b101111101100100 1
#355070000000
0#
0(
#355080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#355130000000
0$
0)
#355140000000
1"
1'
b0 +
b0 1
#355190000000
0"
0'
#355200000000
1#
1(
b101111101100100 +
b101111101100100 1
#355250000000
0#
0(
#355260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#355310000000
0$
0)
#355320000000
1"
1'
b0 +
b0 1
#355370000000
0"
0'
#355380000000
1#
1(
b101111101100100 +
b101111101100100 1
#355430000000
0#
0(
#355440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#355490000000
0$
0)
#355500000000
1"
1'
b0 +
b0 1
#355550000000
0"
0'
#355560000000
1#
1(
b101111101100100 +
b101111101100100 1
#355610000000
0#
0(
#355620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#355670000000
0$
0)
#355680000000
1"
1'
b0 +
b0 1
#355730000000
0"
0'
#355740000000
1#
1(
b101111101100100 +
b101111101100100 1
#355790000000
0#
0(
#355800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#355850000000
0$
0)
#355860000000
1"
1'
b0 +
b0 1
#355910000000
0"
0'
#355920000000
1#
1(
b101111101100100 +
b101111101100100 1
#355970000000
0#
0(
#355980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#356030000000
0$
0)
#356040000000
1"
1'
b0 +
b0 1
#356090000000
0"
0'
#356100000000
1#
1(
b101111101100100 +
b101111101100100 1
#356150000000
0#
0(
#356160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#356210000000
0$
0)
#356220000000
1"
1'
b0 +
b0 1
#356270000000
0"
0'
#356280000000
1#
1(
b101111101100100 +
b101111101100100 1
#356330000000
0#
0(
#356340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#356390000000
0$
0)
#356400000000
1"
1'
b0 +
b0 1
#356450000000
0"
0'
#356460000000
1#
1(
b101111101100100 +
b101111101100100 1
#356510000000
0#
0(
#356520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#356570000000
0$
0)
#356580000000
1"
1'
b0 +
b0 1
#356630000000
0"
0'
#356640000000
1#
1(
b101111101100100 +
b101111101100100 1
#356690000000
0#
0(
#356700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#356750000000
0$
0)
#356760000000
1"
1'
b0 +
b0 1
#356810000000
0"
0'
#356820000000
1#
1(
b101111101100100 +
b101111101100100 1
#356870000000
0#
0(
#356880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#356930000000
0$
0)
#356940000000
1"
1'
b0 +
b0 1
#356990000000
0"
0'
#357000000000
1#
1(
b101111101100100 +
b101111101100100 1
#357050000000
0#
0(
#357060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#357110000000
0$
0)
#357120000000
1"
1'
b0 +
b0 1
#357170000000
0"
0'
#357180000000
1#
1(
b101111101100100 +
b101111101100100 1
#357230000000
0#
0(
#357240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#357290000000
0$
0)
#357300000000
1"
1'
b0 +
b0 1
#357350000000
0"
0'
#357360000000
1#
1(
b101111101100100 +
b101111101100100 1
#357410000000
0#
0(
#357420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#357470000000
0$
0)
#357480000000
1"
1'
b0 +
b0 1
#357530000000
0"
0'
#357540000000
1#
1(
b101111101100100 +
b101111101100100 1
#357590000000
0#
0(
#357600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#357650000000
0$
0)
#357660000000
1"
1'
b0 +
b0 1
#357710000000
0"
0'
#357720000000
1#
1(
b101111101100100 +
b101111101100100 1
#357770000000
0#
0(
#357780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#357830000000
0$
0)
#357840000000
1"
1'
b0 +
b0 1
#357890000000
0"
0'
#357900000000
1#
1(
b101111101100100 +
b101111101100100 1
#357950000000
0#
0(
#357960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#358010000000
0$
0)
#358020000000
1"
1'
b0 +
b0 1
#358070000000
0"
0'
#358080000000
1#
1(
b101111101100100 +
b101111101100100 1
#358130000000
0#
0(
#358140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#358190000000
0$
0)
#358200000000
1"
1'
b0 +
b0 1
#358250000000
0"
0'
#358260000000
1#
1(
b101111101100100 +
b101111101100100 1
#358310000000
0#
0(
#358320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#358370000000
0$
0)
#358380000000
1"
1'
b0 +
b0 1
#358430000000
0"
0'
#358440000000
1#
1(
b101111101100100 +
b101111101100100 1
#358490000000
0#
0(
#358500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#358550000000
0$
0)
#358560000000
1"
1'
b0 +
b0 1
#358610000000
0"
0'
#358620000000
1#
1(
b101111101100100 +
b101111101100100 1
#358670000000
0#
0(
#358680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#358730000000
0$
0)
#358740000000
1"
1'
b0 +
b0 1
#358790000000
0"
0'
#358800000000
1#
1(
b101111101100100 +
b101111101100100 1
#358850000000
0#
0(
#358860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#358910000000
0$
0)
#358920000000
1"
1'
b0 +
b0 1
#358970000000
0"
0'
#358980000000
1#
1(
b101111101100100 +
b101111101100100 1
#359030000000
0#
0(
#359040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#359090000000
0$
0)
#359100000000
1"
1'
b0 +
b0 1
#359150000000
0"
0'
#359160000000
1#
1(
b101111101100100 +
b101111101100100 1
#359210000000
0#
0(
#359220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#359270000000
0$
0)
#359280000000
1"
1'
b0 +
b0 1
#359330000000
0"
0'
#359340000000
1#
1(
b101111101100100 +
b101111101100100 1
#359390000000
0#
0(
#359400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#359450000000
0$
0)
#359460000000
1"
1'
b0 +
b0 1
#359510000000
0"
0'
#359520000000
1#
1(
b101111101100100 +
b101111101100100 1
#359570000000
0#
0(
#359580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#359630000000
0$
0)
#359640000000
1"
1'
b0 +
b0 1
#359690000000
0"
0'
#359700000000
1#
1(
b101111101100100 +
b101111101100100 1
#359750000000
0#
0(
#359760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#359810000000
0$
0)
#359820000000
1"
1'
b0 +
b0 1
#359870000000
0"
0'
#359880000000
1#
1(
b101111101100100 +
b101111101100100 1
#359930000000
0#
0(
#359940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#359990000000
0$
0)
#360000000000
1"
1'
b0 +
b0 1
#360050000000
0"
0'
#360060000000
1#
1(
b101111101100100 +
b101111101100100 1
#360110000000
0#
0(
#360120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#360170000000
0$
0)
#360180000000
1"
1'
b0 +
b0 1
#360230000000
0"
0'
#360240000000
1#
1(
b101111101100100 +
b101111101100100 1
#360290000000
0#
0(
#360300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#360350000000
0$
0)
#360360000000
1"
1'
b0 +
b0 1
#360410000000
0"
0'
#360420000000
1#
1(
b101111101100100 +
b101111101100100 1
#360470000000
0#
0(
#360480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#360530000000
0$
0)
#360540000000
1"
1'
b0 +
b0 1
#360590000000
0"
0'
#360600000000
1#
1(
b101111101100100 +
b101111101100100 1
#360650000000
0#
0(
#360660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#360710000000
0$
0)
#360720000000
1"
1'
b0 +
b0 1
#360770000000
0"
0'
#360780000000
1#
1(
b101111101100100 +
b101111101100100 1
#360830000000
0#
0(
#360840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#360890000000
0$
0)
#360900000000
1"
1'
b0 +
b0 1
#360950000000
0"
0'
#360960000000
1#
1(
b101111101100100 +
b101111101100100 1
#361010000000
0#
0(
#361020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#361070000000
0$
0)
#361080000000
1"
1'
b0 +
b0 1
#361130000000
0"
0'
#361140000000
1#
1(
b101111101100100 +
b101111101100100 1
#361190000000
0#
0(
#361200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#361250000000
0$
0)
#361260000000
1"
1'
b0 +
b0 1
#361310000000
0"
0'
#361320000000
1#
1(
b101111101100100 +
b101111101100100 1
#361370000000
0#
0(
#361380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#361430000000
0$
0)
#361440000000
1"
1'
b0 +
b0 1
#361490000000
0"
0'
#361500000000
1#
1(
b101111101100100 +
b101111101100100 1
#361550000000
0#
0(
#361560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#361610000000
0$
0)
#361620000000
1"
1'
b0 +
b0 1
#361670000000
0"
0'
#361680000000
1#
1(
b101111101100100 +
b101111101100100 1
#361730000000
0#
0(
#361740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#361790000000
0$
0)
#361800000000
1"
1'
b0 +
b0 1
#361850000000
0"
0'
#361860000000
1#
1(
b101111101100100 +
b101111101100100 1
#361910000000
0#
0(
#361920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#361970000000
0$
0)
#361980000000
1"
1'
b0 +
b0 1
#362030000000
0"
0'
#362040000000
1#
1(
b101111101100100 +
b101111101100100 1
#362090000000
0#
0(
#362100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#362150000000
0$
0)
#362160000000
1"
1'
b0 +
b0 1
#362210000000
0"
0'
#362220000000
1#
1(
b101111101100100 +
b101111101100100 1
#362270000000
0#
0(
#362280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#362330000000
0$
0)
#362340000000
1"
1'
b0 +
b0 1
#362390000000
0"
0'
#362400000000
1#
1(
b101111101100100 +
b101111101100100 1
#362450000000
0#
0(
#362460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#362510000000
0$
0)
#362520000000
1"
1'
b0 +
b0 1
#362570000000
0"
0'
#362580000000
1#
1(
b101111101100100 +
b101111101100100 1
#362630000000
0#
0(
#362640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#362690000000
0$
0)
#362700000000
1"
1'
b0 +
b0 1
#362750000000
0"
0'
#362760000000
1#
1(
b101111101100100 +
b101111101100100 1
#362810000000
0#
0(
#362820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#362870000000
0$
0)
#362880000000
1"
1'
b0 +
b0 1
#362930000000
0"
0'
#362940000000
1#
1(
b101111101100100 +
b101111101100100 1
#362990000000
0#
0(
#363000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#363050000000
0$
0)
#363060000000
1"
1'
b0 +
b0 1
#363110000000
0"
0'
#363120000000
1#
1(
b101111101100100 +
b101111101100100 1
#363170000000
0#
0(
#363180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#363230000000
0$
0)
#363240000000
1"
1'
b0 +
b0 1
#363290000000
0"
0'
#363300000000
1#
1(
b101111101100100 +
b101111101100100 1
#363350000000
0#
0(
#363360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#363410000000
0$
0)
#363420000000
1"
1'
b0 +
b0 1
#363470000000
0"
0'
#363480000000
1#
1(
b101111101100100 +
b101111101100100 1
#363530000000
0#
0(
#363540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#363590000000
0$
0)
#363600000000
1"
1'
b0 +
b0 1
#363650000000
0"
0'
#363660000000
1#
1(
b101111101100100 +
b101111101100100 1
#363710000000
0#
0(
#363720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#363770000000
0$
0)
#363780000000
1"
1'
b0 +
b0 1
#363830000000
0"
0'
#363840000000
1#
1(
b101111101100100 +
b101111101100100 1
#363890000000
0#
0(
#363900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#363950000000
0$
0)
#363960000000
1"
1'
b0 +
b0 1
#364010000000
0"
0'
#364020000000
1#
1(
b101111101100100 +
b101111101100100 1
#364070000000
0#
0(
#364080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#364130000000
0$
0)
#364140000000
1"
1'
b0 +
b0 1
#364190000000
0"
0'
#364200000000
1#
1(
b101111101100100 +
b101111101100100 1
#364250000000
0#
0(
#364260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#364310000000
0$
0)
#364320000000
1"
1'
b0 +
b0 1
#364370000000
0"
0'
#364380000000
1#
1(
b101111101100100 +
b101111101100100 1
#364430000000
0#
0(
#364440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#364490000000
0$
0)
#364500000000
1"
1'
b0 +
b0 1
#364550000000
0"
0'
#364560000000
1#
1(
b101111101100100 +
b101111101100100 1
#364610000000
0#
0(
#364620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#364670000000
0$
0)
#364680000000
1"
1'
b0 +
b0 1
#364730000000
0"
0'
#364740000000
1#
1(
b101111101100100 +
b101111101100100 1
#364790000000
0#
0(
#364800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#364850000000
0$
0)
#364860000000
1"
1'
b0 +
b0 1
#364910000000
0"
0'
#364920000000
1#
1(
b101111101100100 +
b101111101100100 1
#364970000000
0#
0(
#364980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#365030000000
0$
0)
#365040000000
1"
1'
b0 +
b0 1
#365090000000
0"
0'
#365100000000
1#
1(
b101111101100100 +
b101111101100100 1
#365150000000
0#
0(
#365160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#365210000000
0$
0)
#365220000000
1"
1'
b0 +
b0 1
#365270000000
0"
0'
#365280000000
1#
1(
b101111101100100 +
b101111101100100 1
#365330000000
0#
0(
#365340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#365390000000
0$
0)
#365400000000
1"
1'
b0 +
b0 1
#365450000000
0"
0'
#365460000000
1#
1(
b101111101100100 +
b101111101100100 1
#365510000000
0#
0(
#365520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#365570000000
0$
0)
#365580000000
1"
1'
b0 +
b0 1
#365630000000
0"
0'
#365640000000
1#
1(
b101111101100100 +
b101111101100100 1
#365690000000
0#
0(
#365700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#365750000000
0$
0)
#365760000000
1"
1'
b0 +
b0 1
#365810000000
0"
0'
#365820000000
1#
1(
b101111101100100 +
b101111101100100 1
#365870000000
0#
0(
#365880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#365930000000
0$
0)
#365940000000
1"
1'
b0 +
b0 1
#365990000000
0"
0'
#366000000000
1#
1(
b101111101100100 +
b101111101100100 1
#366050000000
0#
0(
#366060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#366110000000
0$
0)
#366120000000
1"
1'
b0 +
b0 1
#366170000000
0"
0'
#366180000000
1#
1(
b101111101100100 +
b101111101100100 1
#366230000000
0#
0(
#366240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#366290000000
0$
0)
#366300000000
1"
1'
b0 +
b0 1
#366350000000
0"
0'
#366360000000
1#
1(
b101111101100100 +
b101111101100100 1
#366410000000
0#
0(
#366420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#366470000000
0$
0)
#366480000000
1"
1'
b0 +
b0 1
#366530000000
0"
0'
#366540000000
1#
1(
b101111101100100 +
b101111101100100 1
#366590000000
0#
0(
#366600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#366650000000
0$
0)
#366660000000
1"
1'
b0 +
b0 1
#366710000000
0"
0'
#366720000000
1#
1(
b101111101100100 +
b101111101100100 1
#366770000000
0#
0(
#366780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#366830000000
0$
0)
#366840000000
1"
1'
b0 +
b0 1
#366890000000
0"
0'
#366900000000
1#
1(
b101111101100100 +
b101111101100100 1
#366950000000
0#
0(
#366960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#367010000000
0$
0)
#367020000000
1"
1'
b0 +
b0 1
#367070000000
0"
0'
#367080000000
1#
1(
b101111101100100 +
b101111101100100 1
#367130000000
0#
0(
#367140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#367190000000
0$
0)
#367200000000
1"
1'
b0 +
b0 1
#367250000000
0"
0'
#367260000000
1#
1(
b101111101100100 +
b101111101100100 1
#367310000000
0#
0(
#367320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#367370000000
0$
0)
#367380000000
1"
1'
b0 +
b0 1
#367430000000
0"
0'
#367440000000
1#
1(
b101111101100100 +
b101111101100100 1
#367490000000
0#
0(
#367500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#367550000000
0$
0)
#367560000000
1"
1'
b0 +
b0 1
#367610000000
0"
0'
#367620000000
1#
1(
b101111101100100 +
b101111101100100 1
#367670000000
0#
0(
#367680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#367730000000
0$
0)
#367740000000
1"
1'
b0 +
b0 1
#367790000000
0"
0'
#367800000000
1#
1(
b101111101100100 +
b101111101100100 1
#367850000000
0#
0(
#367860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#367910000000
0$
0)
#367920000000
1"
1'
b0 +
b0 1
#367970000000
0"
0'
#367980000000
1#
1(
b101111101100100 +
b101111101100100 1
#368030000000
0#
0(
#368040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#368090000000
0$
0)
#368100000000
1"
1'
b0 +
b0 1
#368150000000
0"
0'
#368160000000
1#
1(
b101111101100100 +
b101111101100100 1
#368210000000
0#
0(
#368220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#368270000000
0$
0)
#368280000000
1"
1'
b0 +
b0 1
#368330000000
0"
0'
#368340000000
1#
1(
b101111101100100 +
b101111101100100 1
#368390000000
0#
0(
#368400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#368450000000
0$
0)
#368460000000
1"
1'
b0 +
b0 1
#368510000000
0"
0'
#368520000000
1#
1(
b101111101100100 +
b101111101100100 1
#368570000000
0#
0(
#368580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#368630000000
0$
0)
#368640000000
1"
1'
b0 +
b0 1
#368690000000
0"
0'
#368700000000
1#
1(
b101111101100100 +
b101111101100100 1
#368750000000
0#
0(
#368760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#368810000000
0$
0)
#368820000000
1"
1'
b0 +
b0 1
#368870000000
0"
0'
#368880000000
1#
1(
b101111101100100 +
b101111101100100 1
#368930000000
0#
0(
#368940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#368990000000
0$
0)
#369000000000
1"
1'
b0 +
b0 1
#369050000000
0"
0'
#369060000000
1#
1(
b101111101100100 +
b101111101100100 1
#369110000000
0#
0(
#369120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#369170000000
0$
0)
#369180000000
1"
1'
b0 +
b0 1
#369230000000
0"
0'
#369240000000
1#
1(
b101111101100100 +
b101111101100100 1
#369290000000
0#
0(
#369300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#369350000000
0$
0)
#369360000000
1"
1'
b0 +
b0 1
#369410000000
0"
0'
#369420000000
1#
1(
b101111101100100 +
b101111101100100 1
#369470000000
0#
0(
#369480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#369530000000
0$
0)
#369540000000
1"
1'
b0 +
b0 1
#369590000000
0"
0'
#369600000000
1#
1(
b101111101100100 +
b101111101100100 1
#369650000000
0#
0(
#369660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#369710000000
0$
0)
#369720000000
1"
1'
b0 +
b0 1
#369770000000
0"
0'
#369780000000
1#
1(
b101111101100100 +
b101111101100100 1
#369830000000
0#
0(
#369840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#369890000000
0$
0)
#369900000000
1"
1'
b0 +
b0 1
#369950000000
0"
0'
#369960000000
1#
1(
b101111101100100 +
b101111101100100 1
#370010000000
0#
0(
#370020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#370070000000
0$
0)
#370080000000
1"
1'
b0 +
b0 1
#370130000000
0"
0'
#370140000000
1#
1(
b101111101100100 +
b101111101100100 1
#370190000000
0#
0(
#370200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#370250000000
0$
0)
#370260000000
1"
1'
b0 +
b0 1
#370310000000
0"
0'
#370320000000
1#
1(
b101111101100100 +
b101111101100100 1
#370370000000
0#
0(
#370380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#370430000000
0$
0)
#370440000000
1"
1'
b0 +
b0 1
#370490000000
0"
0'
#370500000000
1#
1(
b101111101100100 +
b101111101100100 1
#370550000000
0#
0(
#370560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#370610000000
0$
0)
#370620000000
1"
1'
b0 +
b0 1
#370670000000
0"
0'
#370680000000
1#
1(
b101111101100100 +
b101111101100100 1
#370730000000
0#
0(
#370740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#370790000000
0$
0)
#370800000000
1"
1'
b0 +
b0 1
#370850000000
0"
0'
#370860000000
1#
1(
b101111101100100 +
b101111101100100 1
#370910000000
0#
0(
#370920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#370970000000
0$
0)
#370980000000
1"
1'
b0 +
b0 1
#371030000000
0"
0'
#371040000000
1#
1(
b101111101100100 +
b101111101100100 1
#371090000000
0#
0(
#371100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#371150000000
0$
0)
#371160000000
1"
1'
b0 +
b0 1
#371210000000
0"
0'
#371220000000
1#
1(
b101111101100100 +
b101111101100100 1
#371270000000
0#
0(
#371280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#371330000000
0$
0)
#371340000000
1"
1'
b0 +
b0 1
#371390000000
0"
0'
#371400000000
1#
1(
b101111101100100 +
b101111101100100 1
#371450000000
0#
0(
#371460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#371510000000
0$
0)
#371520000000
1"
1'
b0 +
b0 1
#371570000000
0"
0'
#371580000000
1#
1(
b101111101100100 +
b101111101100100 1
#371630000000
0#
0(
#371640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#371690000000
0$
0)
#371700000000
1"
1'
b0 +
b0 1
#371750000000
0"
0'
#371760000000
1#
1(
b101111101100100 +
b101111101100100 1
#371810000000
0#
0(
#371820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#371870000000
0$
0)
#371880000000
1"
1'
b0 +
b0 1
#371930000000
0"
0'
#371940000000
1#
1(
b101111101100100 +
b101111101100100 1
#371990000000
0#
0(
#372000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#372050000000
0$
0)
#372060000000
1"
1'
b0 +
b0 1
#372110000000
0"
0'
#372120000000
1#
1(
b101111101100100 +
b101111101100100 1
#372170000000
0#
0(
#372180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#372230000000
0$
0)
#372240000000
1"
1'
b0 +
b0 1
#372290000000
0"
0'
#372300000000
1#
1(
b101111101100100 +
b101111101100100 1
#372350000000
0#
0(
#372360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#372410000000
0$
0)
#372420000000
1"
1'
b0 +
b0 1
#372470000000
0"
0'
#372480000000
1#
1(
b101111101100100 +
b101111101100100 1
#372530000000
0#
0(
#372540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#372590000000
0$
0)
#372600000000
1"
1'
b0 +
b0 1
#372650000000
0"
0'
#372660000000
1#
1(
b101111101100100 +
b101111101100100 1
#372710000000
0#
0(
#372720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#372770000000
0$
0)
#372780000000
1"
1'
b0 +
b0 1
#372830000000
0"
0'
#372840000000
1#
1(
b101111101100100 +
b101111101100100 1
#372890000000
0#
0(
#372900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#372950000000
0$
0)
#372960000000
1"
1'
b0 +
b0 1
#373010000000
0"
0'
#373020000000
1#
1(
b101111101100100 +
b101111101100100 1
#373070000000
0#
0(
#373080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#373130000000
0$
0)
#373140000000
1"
1'
b0 +
b0 1
#373190000000
0"
0'
#373200000000
1#
1(
b101111101100100 +
b101111101100100 1
#373250000000
0#
0(
#373260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#373310000000
0$
0)
#373320000000
1"
1'
b0 +
b0 1
#373370000000
0"
0'
#373380000000
1#
1(
b101111101100100 +
b101111101100100 1
#373430000000
0#
0(
#373440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#373490000000
0$
0)
#373500000000
1"
1'
b0 +
b0 1
#373550000000
0"
0'
#373560000000
1#
1(
b101111101100100 +
b101111101100100 1
#373610000000
0#
0(
#373620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#373670000000
0$
0)
#373680000000
1"
1'
b0 +
b0 1
#373730000000
0"
0'
#373740000000
1#
1(
b101111101100100 +
b101111101100100 1
#373790000000
0#
0(
#373800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#373850000000
0$
0)
#373860000000
1"
1'
b0 +
b0 1
#373910000000
0"
0'
#373920000000
1#
1(
b101111101100100 +
b101111101100100 1
#373970000000
0#
0(
#373980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#374030000000
0$
0)
#374040000000
1"
1'
b0 +
b0 1
#374090000000
0"
0'
#374100000000
1#
1(
b101111101100100 +
b101111101100100 1
#374150000000
0#
0(
#374160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#374210000000
0$
0)
#374220000000
1"
1'
b0 +
b0 1
#374270000000
0"
0'
#374280000000
1#
1(
b101111101100100 +
b101111101100100 1
#374330000000
0#
0(
#374340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#374390000000
0$
0)
#374400000000
1"
1'
b0 +
b0 1
#374450000000
0"
0'
#374460000000
1#
1(
b101111101100100 +
b101111101100100 1
#374510000000
0#
0(
#374520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#374570000000
0$
0)
#374580000000
1"
1'
b0 +
b0 1
#374630000000
0"
0'
#374640000000
1#
1(
b101111101100100 +
b101111101100100 1
#374690000000
0#
0(
#374700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#374750000000
0$
0)
#374760000000
1"
1'
b0 +
b0 1
#374810000000
0"
0'
#374820000000
1#
1(
b101111101100100 +
b101111101100100 1
#374870000000
0#
0(
#374880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#374930000000
0$
0)
#374940000000
1"
1'
b0 +
b0 1
#374990000000
0"
0'
#375000000000
1#
1(
b101111101100100 +
b101111101100100 1
#375050000000
0#
0(
#375060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#375110000000
0$
0)
#375120000000
1"
1'
b0 +
b0 1
#375170000000
0"
0'
#375180000000
1#
1(
b101111101100100 +
b101111101100100 1
#375230000000
0#
0(
#375240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#375290000000
0$
0)
#375300000000
1"
1'
b0 +
b0 1
#375350000000
0"
0'
#375360000000
1#
1(
b101111101100100 +
b101111101100100 1
#375410000000
0#
0(
#375420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#375470000000
0$
0)
#375480000000
1"
1'
b0 +
b0 1
#375530000000
0"
0'
#375540000000
1#
1(
b101111101100100 +
b101111101100100 1
#375590000000
0#
0(
#375600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#375650000000
0$
0)
#375660000000
1"
1'
b0 +
b0 1
#375710000000
0"
0'
#375720000000
1#
1(
b101111101100100 +
b101111101100100 1
#375770000000
0#
0(
#375780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#375830000000
0$
0)
#375840000000
1"
1'
b0 +
b0 1
#375890000000
0"
0'
#375900000000
1#
1(
b101111101100100 +
b101111101100100 1
#375950000000
0#
0(
#375960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#376010000000
0$
0)
#376020000000
1"
1'
b0 +
b0 1
#376070000000
0"
0'
#376080000000
1#
1(
b101111101100100 +
b101111101100100 1
#376130000000
0#
0(
#376140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#376190000000
0$
0)
#376200000000
1"
1'
b0 +
b0 1
#376250000000
0"
0'
#376260000000
1#
1(
b101111101100100 +
b101111101100100 1
#376310000000
0#
0(
#376320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#376370000000
0$
0)
#376380000000
1"
1'
b0 +
b0 1
#376430000000
0"
0'
#376440000000
1#
1(
b101111101100100 +
b101111101100100 1
#376490000000
0#
0(
#376500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#376550000000
0$
0)
#376560000000
1"
1'
b0 +
b0 1
#376610000000
0"
0'
#376620000000
1#
1(
b101111101100100 +
b101111101100100 1
#376670000000
0#
0(
#376680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#376730000000
0$
0)
#376740000000
1"
1'
b0 +
b0 1
#376790000000
0"
0'
#376800000000
1#
1(
b101111101100100 +
b101111101100100 1
#376850000000
0#
0(
#376860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#376910000000
0$
0)
#376920000000
1"
1'
b0 +
b0 1
#376970000000
0"
0'
#376980000000
1#
1(
b101111101100100 +
b101111101100100 1
#377030000000
0#
0(
#377040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#377090000000
0$
0)
#377100000000
1"
1'
b0 +
b0 1
#377150000000
0"
0'
#377160000000
1#
1(
b101111101100100 +
b101111101100100 1
#377210000000
0#
0(
#377220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#377270000000
0$
0)
#377280000000
1"
1'
b0 +
b0 1
#377330000000
0"
0'
#377340000000
1#
1(
b101111101100100 +
b101111101100100 1
#377390000000
0#
0(
#377400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#377450000000
0$
0)
#377460000000
1"
1'
b0 +
b0 1
#377510000000
0"
0'
#377520000000
1#
1(
b101111101100100 +
b101111101100100 1
#377570000000
0#
0(
#377580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#377630000000
0$
0)
#377640000000
1"
1'
b0 +
b0 1
#377690000000
0"
0'
#377700000000
1#
1(
b101111101100100 +
b101111101100100 1
#377750000000
0#
0(
#377760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#377810000000
0$
0)
#377820000000
1"
1'
b0 +
b0 1
#377870000000
0"
0'
#377880000000
1#
1(
b101111101100100 +
b101111101100100 1
#377930000000
0#
0(
#377940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#377990000000
0$
0)
#378000000000
1"
1'
b0 +
b0 1
#378050000000
0"
0'
#378060000000
1#
1(
b101111101100100 +
b101111101100100 1
#378110000000
0#
0(
#378120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#378170000000
0$
0)
#378180000000
1"
1'
b0 +
b0 1
#378230000000
0"
0'
#378240000000
1#
1(
b101111101100100 +
b101111101100100 1
#378290000000
0#
0(
#378300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#378350000000
0$
0)
#378360000000
1"
1'
b0 +
b0 1
#378410000000
0"
0'
#378420000000
1#
1(
b101111101100100 +
b101111101100100 1
#378470000000
0#
0(
#378480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#378530000000
0$
0)
#378540000000
1"
1'
b0 +
b0 1
#378590000000
0"
0'
#378600000000
1#
1(
b101111101100100 +
b101111101100100 1
#378650000000
0#
0(
#378660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#378710000000
0$
0)
#378720000000
1"
1'
b0 +
b0 1
#378770000000
0"
0'
#378780000000
1#
1(
b101111101100100 +
b101111101100100 1
#378830000000
0#
0(
#378840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#378890000000
0$
0)
#378900000000
1"
1'
b0 +
b0 1
#378950000000
0"
0'
#378960000000
1#
1(
b101111101100100 +
b101111101100100 1
#379010000000
0#
0(
#379020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#379070000000
0$
0)
#379080000000
1"
1'
b0 +
b0 1
#379130000000
0"
0'
#379140000000
1#
1(
b101111101100100 +
b101111101100100 1
#379190000000
0#
0(
#379200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#379250000000
0$
0)
#379260000000
1"
1'
b0 +
b0 1
#379310000000
0"
0'
#379320000000
1#
1(
b101111101100100 +
b101111101100100 1
#379370000000
0#
0(
#379380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#379430000000
0$
0)
#379440000000
1"
1'
b0 +
b0 1
#379490000000
0"
0'
#379500000000
1#
1(
b101111101100100 +
b101111101100100 1
#379550000000
0#
0(
#379560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#379610000000
0$
0)
#379620000000
1"
1'
b0 +
b0 1
#379670000000
0"
0'
#379680000000
1#
1(
b101111101100100 +
b101111101100100 1
#379730000000
0#
0(
#379740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#379790000000
0$
0)
#379800000000
1"
1'
b0 +
b0 1
#379850000000
0"
0'
#379860000000
1#
1(
b101111101100100 +
b101111101100100 1
#379910000000
0#
0(
#379920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#379970000000
0$
0)
#379980000000
1"
1'
b0 +
b0 1
#380030000000
0"
0'
#380040000000
1#
1(
b101111101100100 +
b101111101100100 1
#380090000000
0#
0(
#380100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#380150000000
0$
0)
#380160000000
1"
1'
b0 +
b0 1
#380210000000
0"
0'
#380220000000
1#
1(
b101111101100100 +
b101111101100100 1
#380270000000
0#
0(
#380280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#380330000000
0$
0)
#380340000000
1"
1'
b0 +
b0 1
#380390000000
0"
0'
#380400000000
1#
1(
b101111101100100 +
b101111101100100 1
#380450000000
0#
0(
#380460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#380510000000
0$
0)
#380520000000
1"
1'
b0 +
b0 1
#380570000000
0"
0'
#380580000000
1#
1(
b101111101100100 +
b101111101100100 1
#380630000000
0#
0(
#380640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#380690000000
0$
0)
#380700000000
1"
1'
b0 +
b0 1
#380750000000
0"
0'
#380760000000
1#
1(
b101111101100100 +
b101111101100100 1
#380810000000
0#
0(
#380820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#380870000000
0$
0)
#380880000000
1"
1'
b0 +
b0 1
#380930000000
0"
0'
#380940000000
1#
1(
b101111101100100 +
b101111101100100 1
#380990000000
0#
0(
#381000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#381050000000
0$
0)
#381060000000
1"
1'
b0 +
b0 1
#381110000000
0"
0'
#381120000000
1#
1(
b101111101100100 +
b101111101100100 1
#381170000000
0#
0(
#381180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#381230000000
0$
0)
#381240000000
1"
1'
b0 +
b0 1
#381290000000
0"
0'
#381300000000
1#
1(
b101111101100100 +
b101111101100100 1
#381350000000
0#
0(
#381360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#381410000000
0$
0)
#381420000000
1"
1'
b0 +
b0 1
#381470000000
0"
0'
#381480000000
1#
1(
b101111101100100 +
b101111101100100 1
#381530000000
0#
0(
#381540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#381590000000
0$
0)
#381600000000
1"
1'
b0 +
b0 1
#381650000000
0"
0'
#381660000000
1#
1(
b101111101100100 +
b101111101100100 1
#381710000000
0#
0(
#381720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#381770000000
0$
0)
#381780000000
1"
1'
b0 +
b0 1
#381830000000
0"
0'
#381840000000
1#
1(
b101111101100100 +
b101111101100100 1
#381890000000
0#
0(
#381900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#381950000000
0$
0)
#381960000000
1"
1'
b0 +
b0 1
#382010000000
0"
0'
#382020000000
1#
1(
b101111101100100 +
b101111101100100 1
#382070000000
0#
0(
#382080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#382130000000
0$
0)
#382140000000
1"
1'
b0 +
b0 1
#382190000000
0"
0'
#382200000000
1#
1(
b101111101100100 +
b101111101100100 1
#382250000000
0#
0(
#382260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#382310000000
0$
0)
#382320000000
1"
1'
b0 +
b0 1
#382370000000
0"
0'
#382380000000
1#
1(
b101111101100100 +
b101111101100100 1
#382430000000
0#
0(
#382440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#382490000000
0$
0)
#382500000000
1"
1'
b0 +
b0 1
#382550000000
0"
0'
#382560000000
1#
1(
b101111101100100 +
b101111101100100 1
#382610000000
0#
0(
#382620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#382670000000
0$
0)
#382680000000
1"
1'
b0 +
b0 1
#382730000000
0"
0'
#382740000000
1#
1(
b101111101100100 +
b101111101100100 1
#382790000000
0#
0(
#382800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#382850000000
0$
0)
#382860000000
1"
1'
b0 +
b0 1
#382910000000
0"
0'
#382920000000
1#
1(
b101111101100100 +
b101111101100100 1
#382970000000
0#
0(
#382980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#383030000000
0$
0)
#383040000000
1"
1'
b0 +
b0 1
#383090000000
0"
0'
#383100000000
1#
1(
b101111101100100 +
b101111101100100 1
#383150000000
0#
0(
#383160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#383210000000
0$
0)
#383220000000
1"
1'
b0 +
b0 1
#383270000000
0"
0'
#383280000000
1#
1(
b101111101100100 +
b101111101100100 1
#383330000000
0#
0(
#383340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#383390000000
0$
0)
#383400000000
1"
1'
b0 +
b0 1
#383450000000
0"
0'
#383460000000
1#
1(
b101111101100100 +
b101111101100100 1
#383510000000
0#
0(
#383520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#383570000000
0$
0)
#383580000000
1"
1'
b0 +
b0 1
#383630000000
0"
0'
#383640000000
1#
1(
b101111101100100 +
b101111101100100 1
#383690000000
0#
0(
#383700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#383750000000
0$
0)
#383760000000
1"
1'
b0 +
b0 1
#383810000000
0"
0'
#383820000000
1#
1(
b101111101100100 +
b101111101100100 1
#383870000000
0#
0(
#383880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#383930000000
0$
0)
#383940000000
1"
1'
b0 +
b0 1
#383990000000
0"
0'
#384000000000
1#
1(
b101111101100100 +
b101111101100100 1
#384050000000
0#
0(
#384060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#384110000000
0$
0)
#384120000000
1"
1'
b0 +
b0 1
#384170000000
0"
0'
#384180000000
1#
1(
b101111101100100 +
b101111101100100 1
#384230000000
0#
0(
#384240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#384290000000
0$
0)
#384300000000
1"
1'
b0 +
b0 1
#384350000000
0"
0'
#384360000000
1#
1(
b101111101100100 +
b101111101100100 1
#384410000000
0#
0(
#384420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#384470000000
0$
0)
#384480000000
1"
1'
b0 +
b0 1
#384530000000
0"
0'
#384540000000
1#
1(
b101111101100100 +
b101111101100100 1
#384590000000
0#
0(
#384600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#384650000000
0$
0)
#384660000000
1"
1'
b0 +
b0 1
#384710000000
0"
0'
#384720000000
1#
1(
b101111101100100 +
b101111101100100 1
#384770000000
0#
0(
#384780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#384830000000
0$
0)
#384840000000
1"
1'
b0 +
b0 1
#384890000000
0"
0'
#384900000000
1#
1(
b101111101100100 +
b101111101100100 1
#384950000000
0#
0(
#384960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#385010000000
0$
0)
#385020000000
1"
1'
b0 +
b0 1
#385070000000
0"
0'
#385080000000
1#
1(
b101111101100100 +
b101111101100100 1
#385130000000
0#
0(
#385140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#385190000000
0$
0)
#385200000000
1"
1'
b0 +
b0 1
#385250000000
0"
0'
#385260000000
1#
1(
b101111101100100 +
b101111101100100 1
#385310000000
0#
0(
#385320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#385370000000
0$
0)
#385380000000
1"
1'
b0 +
b0 1
#385430000000
0"
0'
#385440000000
1#
1(
b101111101100100 +
b101111101100100 1
#385490000000
0#
0(
#385500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#385550000000
0$
0)
#385560000000
1"
1'
b0 +
b0 1
#385610000000
0"
0'
#385620000000
1#
1(
b101111101100100 +
b101111101100100 1
#385670000000
0#
0(
#385680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#385730000000
0$
0)
#385740000000
1"
1'
b0 +
b0 1
#385790000000
0"
0'
#385800000000
1#
1(
b101111101100100 +
b101111101100100 1
#385850000000
0#
0(
#385860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#385910000000
0$
0)
#385920000000
1"
1'
b0 +
b0 1
#385970000000
0"
0'
#385980000000
1#
1(
b101111101100100 +
b101111101100100 1
#386030000000
0#
0(
#386040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#386090000000
0$
0)
#386100000000
1"
1'
b0 +
b0 1
#386150000000
0"
0'
#386160000000
1#
1(
b101111101100100 +
b101111101100100 1
#386210000000
0#
0(
#386220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#386270000000
0$
0)
#386280000000
1"
1'
b0 +
b0 1
#386330000000
0"
0'
#386340000000
1#
1(
b101111101100100 +
b101111101100100 1
#386390000000
0#
0(
#386400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#386450000000
0$
0)
#386460000000
1"
1'
b0 +
b0 1
#386510000000
0"
0'
#386520000000
1#
1(
b101111101100100 +
b101111101100100 1
#386570000000
0#
0(
#386580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#386630000000
0$
0)
#386640000000
1"
1'
b0 +
b0 1
#386690000000
0"
0'
#386700000000
1#
1(
b101111101100100 +
b101111101100100 1
#386750000000
0#
0(
#386760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#386810000000
0$
0)
#386820000000
1"
1'
b0 +
b0 1
#386870000000
0"
0'
#386880000000
1#
1(
b101111101100100 +
b101111101100100 1
#386930000000
0#
0(
#386940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#386990000000
0$
0)
#387000000000
1"
1'
b0 +
b0 1
#387050000000
0"
0'
#387060000000
1#
1(
b101111101100100 +
b101111101100100 1
#387110000000
0#
0(
#387120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#387170000000
0$
0)
#387180000000
1"
1'
b0 +
b0 1
#387230000000
0"
0'
#387240000000
1#
1(
b101111101100100 +
b101111101100100 1
#387290000000
0#
0(
#387300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#387350000000
0$
0)
#387360000000
1"
1'
b0 +
b0 1
#387410000000
0"
0'
#387420000000
1#
1(
b101111101100100 +
b101111101100100 1
#387470000000
0#
0(
#387480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#387530000000
0$
0)
#387540000000
1"
1'
b0 +
b0 1
#387590000000
0"
0'
#387600000000
1#
1(
b101111101100100 +
b101111101100100 1
#387650000000
0#
0(
#387660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#387710000000
0$
0)
#387720000000
1"
1'
b0 +
b0 1
#387770000000
0"
0'
#387780000000
1#
1(
b101111101100100 +
b101111101100100 1
#387830000000
0#
0(
#387840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#387890000000
0$
0)
#387900000000
1"
1'
b0 +
b0 1
#387950000000
0"
0'
#387960000000
1#
1(
b101111101100100 +
b101111101100100 1
#388010000000
0#
0(
#388020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#388070000000
0$
0)
#388080000000
1"
1'
b0 +
b0 1
#388130000000
0"
0'
#388140000000
1#
1(
b101111101100100 +
b101111101100100 1
#388190000000
0#
0(
#388200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#388250000000
0$
0)
#388260000000
1"
1'
b0 +
b0 1
#388310000000
0"
0'
#388320000000
1#
1(
b101111101100100 +
b101111101100100 1
#388370000000
0#
0(
#388380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#388430000000
0$
0)
#388440000000
1"
1'
b0 +
b0 1
#388490000000
0"
0'
#388500000000
1#
1(
b101111101100100 +
b101111101100100 1
#388550000000
0#
0(
#388560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#388610000000
0$
0)
#388620000000
1"
1'
b0 +
b0 1
#388670000000
0"
0'
#388680000000
1#
1(
b101111101100100 +
b101111101100100 1
#388730000000
0#
0(
#388740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#388790000000
0$
0)
#388800000000
1"
1'
b0 +
b0 1
#388850000000
0"
0'
#388860000000
1#
1(
b101111101100100 +
b101111101100100 1
#388910000000
0#
0(
#388920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#388970000000
0$
0)
#388980000000
1"
1'
b0 +
b0 1
#389030000000
0"
0'
#389040000000
1#
1(
b101111101100100 +
b101111101100100 1
#389090000000
0#
0(
#389100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#389150000000
0$
0)
#389160000000
1"
1'
b0 +
b0 1
#389210000000
0"
0'
#389220000000
1#
1(
b101111101100100 +
b101111101100100 1
#389270000000
0#
0(
#389280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#389330000000
0$
0)
#389340000000
1"
1'
b0 +
b0 1
#389390000000
0"
0'
#389400000000
1#
1(
b101111101100100 +
b101111101100100 1
#389450000000
0#
0(
#389460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#389510000000
0$
0)
#389520000000
1"
1'
b0 +
b0 1
#389570000000
0"
0'
#389580000000
1#
1(
b101111101100100 +
b101111101100100 1
#389630000000
0#
0(
#389640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#389690000000
0$
0)
#389700000000
1"
1'
b0 +
b0 1
#389750000000
0"
0'
#389760000000
1#
1(
b101111101100100 +
b101111101100100 1
#389810000000
0#
0(
#389820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#389870000000
0$
0)
#389880000000
1"
1'
b0 +
b0 1
#389930000000
0"
0'
#389940000000
1#
1(
b101111101100100 +
b101111101100100 1
#389990000000
0#
0(
#390000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#390050000000
0$
0)
#390060000000
1"
1'
b0 +
b0 1
#390110000000
0"
0'
#390120000000
1#
1(
b101111101100100 +
b101111101100100 1
#390170000000
0#
0(
#390180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#390230000000
0$
0)
#390240000000
1"
1'
b0 +
b0 1
#390290000000
0"
0'
#390300000000
1#
1(
b101111101100100 +
b101111101100100 1
#390350000000
0#
0(
#390360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#390410000000
0$
0)
#390420000000
1"
1'
b0 +
b0 1
#390470000000
0"
0'
#390480000000
1#
1(
b101111101100100 +
b101111101100100 1
#390530000000
0#
0(
#390540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#390590000000
0$
0)
#390600000000
1"
1'
b0 +
b0 1
#390650000000
0"
0'
#390660000000
1#
1(
b101111101100100 +
b101111101100100 1
#390710000000
0#
0(
#390720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#390770000000
0$
0)
#390780000000
1"
1'
b0 +
b0 1
#390830000000
0"
0'
#390840000000
1#
1(
b101111101100100 +
b101111101100100 1
#390890000000
0#
0(
#390900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#390950000000
0$
0)
#390960000000
1"
1'
b0 +
b0 1
#391010000000
0"
0'
#391020000000
1#
1(
b101111101100100 +
b101111101100100 1
#391070000000
0#
0(
#391080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#391130000000
0$
0)
#391140000000
1"
1'
b0 +
b0 1
#391190000000
0"
0'
#391200000000
1#
1(
b101111101100100 +
b101111101100100 1
#391250000000
0#
0(
#391260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#391310000000
0$
0)
#391320000000
1"
1'
b0 +
b0 1
#391370000000
0"
0'
#391380000000
1#
1(
b101111101100100 +
b101111101100100 1
#391430000000
0#
0(
#391440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#391490000000
0$
0)
#391500000000
1"
1'
b0 +
b0 1
#391550000000
0"
0'
#391560000000
1#
1(
b101111101100100 +
b101111101100100 1
#391610000000
0#
0(
#391620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#391670000000
0$
0)
#391680000000
1"
1'
b0 +
b0 1
#391730000000
0"
0'
#391740000000
1#
1(
b101111101100100 +
b101111101100100 1
#391790000000
0#
0(
#391800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#391850000000
0$
0)
#391860000000
1"
1'
b0 +
b0 1
#391910000000
0"
0'
#391920000000
1#
1(
b101111101100100 +
b101111101100100 1
#391970000000
0#
0(
#391980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#392030000000
0$
0)
#392040000000
1"
1'
b0 +
b0 1
#392090000000
0"
0'
#392100000000
1#
1(
b101111101100100 +
b101111101100100 1
#392150000000
0#
0(
#392160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#392210000000
0$
0)
#392220000000
1"
1'
b0 +
b0 1
#392270000000
0"
0'
#392280000000
1#
1(
b101111101100100 +
b101111101100100 1
#392330000000
0#
0(
#392340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#392390000000
0$
0)
#392400000000
1"
1'
b0 +
b0 1
#392450000000
0"
0'
#392460000000
1#
1(
b101111101100100 +
b101111101100100 1
#392510000000
0#
0(
#392520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#392570000000
0$
0)
#392580000000
1"
1'
b0 +
b0 1
#392630000000
0"
0'
#392640000000
1#
1(
b101111101100100 +
b101111101100100 1
#392690000000
0#
0(
#392700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#392750000000
0$
0)
#392760000000
1"
1'
b0 +
b0 1
#392810000000
0"
0'
#392820000000
1#
1(
b101111101100100 +
b101111101100100 1
#392870000000
0#
0(
#392880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#392930000000
0$
0)
#392940000000
1"
1'
b0 +
b0 1
#392990000000
0"
0'
#393000000000
1#
1(
b101111101100100 +
b101111101100100 1
#393050000000
0#
0(
#393060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#393110000000
0$
0)
#393120000000
1"
1'
b0 +
b0 1
#393170000000
0"
0'
#393180000000
1#
1(
b101111101100100 +
b101111101100100 1
#393230000000
0#
0(
#393240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#393290000000
0$
0)
#393300000000
1"
1'
b0 +
b0 1
#393350000000
0"
0'
#393360000000
1#
1(
b101111101100100 +
b101111101100100 1
#393410000000
0#
0(
#393420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#393470000000
0$
0)
#393480000000
1"
1'
b0 +
b0 1
#393530000000
0"
0'
#393540000000
1#
1(
b101111101100100 +
b101111101100100 1
#393590000000
0#
0(
#393600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#393650000000
0$
0)
#393660000000
1"
1'
b0 +
b0 1
#393710000000
0"
0'
#393720000000
1#
1(
b101111101100100 +
b101111101100100 1
#393770000000
0#
0(
#393780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#393830000000
0$
0)
#393840000000
1"
1'
b0 +
b0 1
#393890000000
0"
0'
#393900000000
1#
1(
b101111101100100 +
b101111101100100 1
#393950000000
0#
0(
#393960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#394010000000
0$
0)
#394020000000
1"
1'
b0 +
b0 1
#394070000000
0"
0'
#394080000000
1#
1(
b101111101100100 +
b101111101100100 1
#394130000000
0#
0(
#394140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#394190000000
0$
0)
#394200000000
1"
1'
b0 +
b0 1
#394250000000
0"
0'
#394260000000
1#
1(
b101111101100100 +
b101111101100100 1
#394310000000
0#
0(
#394320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#394370000000
0$
0)
#394380000000
1"
1'
b0 +
b0 1
#394430000000
0"
0'
#394440000000
1#
1(
b101111101100100 +
b101111101100100 1
#394490000000
0#
0(
#394500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#394550000000
0$
0)
#394560000000
1"
1'
b0 +
b0 1
#394610000000
0"
0'
#394620000000
1#
1(
b101111101100100 +
b101111101100100 1
#394670000000
0#
0(
#394680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#394730000000
0$
0)
#394740000000
1"
1'
b0 +
b0 1
#394790000000
0"
0'
#394800000000
1#
1(
b101111101100100 +
b101111101100100 1
#394850000000
0#
0(
#394860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#394910000000
0$
0)
#394920000000
1"
1'
b0 +
b0 1
#394970000000
0"
0'
#394980000000
1#
1(
b101111101100100 +
b101111101100100 1
#395030000000
0#
0(
#395040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#395090000000
0$
0)
#395100000000
1"
1'
b0 +
b0 1
#395150000000
0"
0'
#395160000000
1#
1(
b101111101100100 +
b101111101100100 1
#395210000000
0#
0(
#395220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#395270000000
0$
0)
#395280000000
1"
1'
b0 +
b0 1
#395330000000
0"
0'
#395340000000
1#
1(
b101111101100100 +
b101111101100100 1
#395390000000
0#
0(
#395400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#395450000000
0$
0)
#395460000000
1"
1'
b0 +
b0 1
#395510000000
0"
0'
#395520000000
1#
1(
b101111101100100 +
b101111101100100 1
#395570000000
0#
0(
#395580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#395630000000
0$
0)
#395640000000
1"
1'
b0 +
b0 1
#395690000000
0"
0'
#395700000000
1#
1(
b101111101100100 +
b101111101100100 1
#395750000000
0#
0(
#395760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#395810000000
0$
0)
#395820000000
1"
1'
b0 +
b0 1
#395870000000
0"
0'
#395880000000
1#
1(
b101111101100100 +
b101111101100100 1
#395930000000
0#
0(
#395940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#395990000000
0$
0)
#396000000000
1"
1'
b0 +
b0 1
#396050000000
0"
0'
#396060000000
1#
1(
b101111101100100 +
b101111101100100 1
#396110000000
0#
0(
#396120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#396170000000
0$
0)
#396180000000
1"
1'
b0 +
b0 1
#396230000000
0"
0'
#396240000000
1#
1(
b101111101100100 +
b101111101100100 1
#396290000000
0#
0(
#396300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#396350000000
0$
0)
#396360000000
1"
1'
b0 +
b0 1
#396410000000
0"
0'
#396420000000
1#
1(
b101111101100100 +
b101111101100100 1
#396470000000
0#
0(
#396480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#396530000000
0$
0)
#396540000000
1"
1'
b0 +
b0 1
#396590000000
0"
0'
#396600000000
1#
1(
b101111101100100 +
b101111101100100 1
#396650000000
0#
0(
#396660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#396710000000
0$
0)
#396720000000
1"
1'
b0 +
b0 1
#396770000000
0"
0'
#396780000000
1#
1(
b101111101100100 +
b101111101100100 1
#396830000000
0#
0(
#396840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#396890000000
0$
0)
#396900000000
1"
1'
b0 +
b0 1
#396950000000
0"
0'
#396960000000
1#
1(
b101111101100100 +
b101111101100100 1
#397010000000
0#
0(
#397020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#397070000000
0$
0)
#397080000000
1"
1'
b0 +
b0 1
#397130000000
0"
0'
#397140000000
1#
1(
b101111101100100 +
b101111101100100 1
#397190000000
0#
0(
#397200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#397250000000
0$
0)
#397260000000
1"
1'
b0 +
b0 1
#397310000000
0"
0'
#397320000000
1#
1(
b101111101100100 +
b101111101100100 1
#397370000000
0#
0(
#397380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#397430000000
0$
0)
#397440000000
1"
1'
b0 +
b0 1
#397490000000
0"
0'
#397500000000
1#
1(
b101111101100100 +
b101111101100100 1
#397550000000
0#
0(
#397560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#397610000000
0$
0)
#397620000000
1"
1'
b0 +
b0 1
#397670000000
0"
0'
#397680000000
1#
1(
b101111101100100 +
b101111101100100 1
#397730000000
0#
0(
#397740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#397790000000
0$
0)
#397800000000
1"
1'
b0 +
b0 1
#397850000000
0"
0'
#397860000000
1#
1(
b101111101100100 +
b101111101100100 1
#397910000000
0#
0(
#397920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#397970000000
0$
0)
#397980000000
1"
1'
b0 +
b0 1
#398030000000
0"
0'
#398040000000
1#
1(
b101111101100100 +
b101111101100100 1
#398090000000
0#
0(
#398100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#398150000000
0$
0)
#398160000000
1"
1'
b0 +
b0 1
#398210000000
0"
0'
#398220000000
1#
1(
b101111101100100 +
b101111101100100 1
#398270000000
0#
0(
#398280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#398330000000
0$
0)
#398340000000
1"
1'
b0 +
b0 1
#398390000000
0"
0'
#398400000000
1#
1(
b101111101100100 +
b101111101100100 1
#398450000000
0#
0(
#398460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#398510000000
0$
0)
#398520000000
1"
1'
b0 +
b0 1
#398570000000
0"
0'
#398580000000
1#
1(
b101111101100100 +
b101111101100100 1
#398630000000
0#
0(
#398640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#398690000000
0$
0)
#398700000000
1"
1'
b0 +
b0 1
#398750000000
0"
0'
#398760000000
1#
1(
b101111101100100 +
b101111101100100 1
#398810000000
0#
0(
#398820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#398870000000
0$
0)
#398880000000
1"
1'
b0 +
b0 1
#398930000000
0"
0'
#398940000000
1#
1(
b101111101100100 +
b101111101100100 1
#398990000000
0#
0(
#399000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#399050000000
0$
0)
#399060000000
1"
1'
b0 +
b0 1
#399110000000
0"
0'
#399120000000
1#
1(
b101111101100100 +
b101111101100100 1
#399170000000
0#
0(
#399180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#399230000000
0$
0)
#399240000000
1"
1'
b0 +
b0 1
#399290000000
0"
0'
#399300000000
1#
1(
b101111101100100 +
b101111101100100 1
#399350000000
0#
0(
#399360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#399410000000
0$
0)
#399420000000
1"
1'
b0 +
b0 1
#399470000000
0"
0'
#399480000000
1#
1(
b101111101100100 +
b101111101100100 1
#399530000000
0#
0(
#399540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#399590000000
0$
0)
#399600000000
1"
1'
b0 +
b0 1
#399650000000
0"
0'
#399660000000
1#
1(
b101111101100100 +
b101111101100100 1
#399710000000
0#
0(
#399720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#399770000000
0$
0)
#399780000000
1"
1'
b0 +
b0 1
#399830000000
0"
0'
#399840000000
1#
1(
b101111101100100 +
b101111101100100 1
#399890000000
0#
0(
#399900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#399950000000
0$
0)
#399960000000
1"
1'
b0 +
b0 1
#400010000000
0"
0'
#400020000000
1#
1(
b101111101100100 +
b101111101100100 1
#400070000000
0#
0(
#400080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#400130000000
0$
0)
#400140000000
1"
1'
b0 +
b0 1
#400190000000
0"
0'
#400200000000
1#
1(
b101111101100100 +
b101111101100100 1
#400250000000
0#
0(
#400260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#400310000000
0$
0)
#400320000000
1"
1'
b0 +
b0 1
#400370000000
0"
0'
#400380000000
1#
1(
b101111101100100 +
b101111101100100 1
#400430000000
0#
0(
#400440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#400490000000
0$
0)
#400500000000
1"
1'
b0 +
b0 1
#400550000000
0"
0'
#400560000000
1#
1(
b101111101100100 +
b101111101100100 1
#400610000000
0#
0(
#400620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#400670000000
0$
0)
#400680000000
1"
1'
b0 +
b0 1
#400730000000
0"
0'
#400740000000
1#
1(
b101111101100100 +
b101111101100100 1
#400790000000
0#
0(
#400800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#400850000000
0$
0)
#400860000000
1"
1'
b0 +
b0 1
#400910000000
0"
0'
#400920000000
1#
1(
b101111101100100 +
b101111101100100 1
#400970000000
0#
0(
#400980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#401030000000
0$
0)
#401040000000
1"
1'
b0 +
b0 1
#401090000000
0"
0'
#401100000000
1#
1(
b101111101100100 +
b101111101100100 1
#401150000000
0#
0(
#401160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#401210000000
0$
0)
#401220000000
1"
1'
b0 +
b0 1
#401270000000
0"
0'
#401280000000
1#
1(
b101111101100100 +
b101111101100100 1
#401330000000
0#
0(
#401340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#401390000000
0$
0)
#401400000000
1"
1'
b0 +
b0 1
#401450000000
0"
0'
#401460000000
1#
1(
b101111101100100 +
b101111101100100 1
#401510000000
0#
0(
#401520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#401570000000
0$
0)
#401580000000
1"
1'
b0 +
b0 1
#401630000000
0"
0'
#401640000000
1#
1(
b101111101100100 +
b101111101100100 1
#401690000000
0#
0(
#401700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#401750000000
0$
0)
#401760000000
1"
1'
b0 +
b0 1
#401810000000
0"
0'
#401820000000
1#
1(
b101111101100100 +
b101111101100100 1
#401870000000
0#
0(
#401880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#401930000000
0$
0)
#401940000000
1"
1'
b0 +
b0 1
#401990000000
0"
0'
#402000000000
1#
1(
b101111101100100 +
b101111101100100 1
#402050000000
0#
0(
#402060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#402110000000
0$
0)
#402120000000
1"
1'
b0 +
b0 1
#402170000000
0"
0'
#402180000000
1#
1(
b101111101100100 +
b101111101100100 1
#402230000000
0#
0(
#402240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#402290000000
0$
0)
#402300000000
1"
1'
b0 +
b0 1
#402350000000
0"
0'
#402360000000
1#
1(
b101111101100100 +
b101111101100100 1
#402410000000
0#
0(
#402420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#402470000000
0$
0)
#402480000000
1"
1'
b0 +
b0 1
#402530000000
0"
0'
#402540000000
1#
1(
b101111101100100 +
b101111101100100 1
#402590000000
0#
0(
#402600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#402650000000
0$
0)
#402660000000
1"
1'
b0 +
b0 1
#402710000000
0"
0'
#402720000000
1#
1(
b101111101100100 +
b101111101100100 1
#402770000000
0#
0(
#402780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#402830000000
0$
0)
#402840000000
1"
1'
b0 +
b0 1
#402890000000
0"
0'
#402900000000
1#
1(
b101111101100100 +
b101111101100100 1
#402950000000
0#
0(
#402960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#403010000000
0$
0)
#403020000000
1"
1'
b0 +
b0 1
#403070000000
0"
0'
#403080000000
1#
1(
b101111101100100 +
b101111101100100 1
#403130000000
0#
0(
#403140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#403190000000
0$
0)
#403200000000
1"
1'
b0 +
b0 1
#403250000000
0"
0'
#403260000000
1#
1(
b101111101100100 +
b101111101100100 1
#403310000000
0#
0(
#403320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#403370000000
0$
0)
#403380000000
1"
1'
b0 +
b0 1
#403430000000
0"
0'
#403440000000
1#
1(
b101111101100100 +
b101111101100100 1
#403490000000
0#
0(
#403500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#403550000000
0$
0)
#403560000000
1"
1'
b0 +
b0 1
#403610000000
0"
0'
#403620000000
1#
1(
b101111101100100 +
b101111101100100 1
#403670000000
0#
0(
#403680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#403730000000
0$
0)
#403740000000
1"
1'
b0 +
b0 1
#403790000000
0"
0'
#403800000000
1#
1(
b101111101100100 +
b101111101100100 1
#403850000000
0#
0(
#403860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#403910000000
0$
0)
#403920000000
1"
1'
b0 +
b0 1
#403970000000
0"
0'
#403980000000
1#
1(
b101111101100100 +
b101111101100100 1
#404030000000
0#
0(
#404040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#404090000000
0$
0)
#404100000000
1"
1'
b0 +
b0 1
#404150000000
0"
0'
#404160000000
1#
1(
b101111101100100 +
b101111101100100 1
#404210000000
0#
0(
#404220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#404270000000
0$
0)
#404280000000
1"
1'
b0 +
b0 1
#404330000000
0"
0'
#404340000000
1#
1(
b101111101100100 +
b101111101100100 1
#404390000000
0#
0(
#404400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#404450000000
0$
0)
#404460000000
1"
1'
b0 +
b0 1
#404510000000
0"
0'
#404520000000
1#
1(
b101111101100100 +
b101111101100100 1
#404570000000
0#
0(
#404580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#404630000000
0$
0)
#404640000000
1"
1'
b0 +
b0 1
#404690000000
0"
0'
#404700000000
1#
1(
b101111101100100 +
b101111101100100 1
#404750000000
0#
0(
#404760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#404810000000
0$
0)
#404820000000
1"
1'
b0 +
b0 1
#404870000000
0"
0'
#404880000000
1#
1(
b101111101100100 +
b101111101100100 1
#404930000000
0#
0(
#404940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#404990000000
0$
0)
#405000000000
1"
1'
b0 +
b0 1
#405050000000
0"
0'
#405060000000
1#
1(
b101111101100100 +
b101111101100100 1
#405110000000
0#
0(
#405120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#405170000000
0$
0)
#405180000000
1"
1'
b0 +
b0 1
#405230000000
0"
0'
#405240000000
1#
1(
b101111101100100 +
b101111101100100 1
#405290000000
0#
0(
#405300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#405350000000
0$
0)
#405360000000
1"
1'
b0 +
b0 1
#405410000000
0"
0'
#405420000000
1#
1(
b101111101100100 +
b101111101100100 1
#405470000000
0#
0(
#405480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#405530000000
0$
0)
#405540000000
1"
1'
b0 +
b0 1
#405590000000
0"
0'
#405600000000
1#
1(
b101111101100100 +
b101111101100100 1
#405650000000
0#
0(
#405660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#405710000000
0$
0)
#405720000000
1"
1'
b0 +
b0 1
#405770000000
0"
0'
#405780000000
1#
1(
b101111101100100 +
b101111101100100 1
#405830000000
0#
0(
#405840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#405890000000
0$
0)
#405900000000
1"
1'
b0 +
b0 1
#405950000000
0"
0'
#405960000000
1#
1(
b101111101100100 +
b101111101100100 1
#406010000000
0#
0(
#406020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#406070000000
0$
0)
#406080000000
1"
1'
b0 +
b0 1
#406130000000
0"
0'
#406140000000
1#
1(
b101111101100100 +
b101111101100100 1
#406190000000
0#
0(
#406200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#406250000000
0$
0)
#406260000000
1"
1'
b0 +
b0 1
#406310000000
0"
0'
#406320000000
1#
1(
b101111101100100 +
b101111101100100 1
#406370000000
0#
0(
#406380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#406430000000
0$
0)
#406440000000
1"
1'
b0 +
b0 1
#406490000000
0"
0'
#406500000000
1#
1(
b101111101100100 +
b101111101100100 1
#406550000000
0#
0(
#406560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#406610000000
0$
0)
#406620000000
1"
1'
b0 +
b0 1
#406670000000
0"
0'
#406680000000
1#
1(
b101111101100100 +
b101111101100100 1
#406730000000
0#
0(
#406740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#406790000000
0$
0)
#406800000000
1"
1'
b0 +
b0 1
#406850000000
0"
0'
#406860000000
1#
1(
b101111101100100 +
b101111101100100 1
#406910000000
0#
0(
#406920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#406970000000
0$
0)
#406980000000
1"
1'
b0 +
b0 1
#407030000000
0"
0'
#407040000000
1#
1(
b101111101100100 +
b101111101100100 1
#407090000000
0#
0(
#407100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#407150000000
0$
0)
#407160000000
1"
1'
b0 +
b0 1
#407210000000
0"
0'
#407220000000
1#
1(
b101111101100100 +
b101111101100100 1
#407270000000
0#
0(
#407280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#407330000000
0$
0)
#407340000000
1"
1'
b0 +
b0 1
#407390000000
0"
0'
#407400000000
1#
1(
b101111101100100 +
b101111101100100 1
#407450000000
0#
0(
#407460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#407510000000
0$
0)
#407520000000
1"
1'
b0 +
b0 1
#407570000000
0"
0'
#407580000000
1#
1(
b101111101100100 +
b101111101100100 1
#407630000000
0#
0(
#407640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#407690000000
0$
0)
#407700000000
1"
1'
b0 +
b0 1
#407750000000
0"
0'
#407760000000
1#
1(
b101111101100100 +
b101111101100100 1
#407810000000
0#
0(
#407820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#407870000000
0$
0)
#407880000000
1"
1'
b0 +
b0 1
#407930000000
0"
0'
#407940000000
1#
1(
b101111101100100 +
b101111101100100 1
#407990000000
0#
0(
#408000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#408050000000
0$
0)
#408060000000
1"
1'
b0 +
b0 1
#408110000000
0"
0'
#408120000000
1#
1(
b101111101100100 +
b101111101100100 1
#408170000000
0#
0(
#408180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#408230000000
0$
0)
#408240000000
1"
1'
b0 +
b0 1
#408290000000
0"
0'
#408300000000
1#
1(
b101111101100100 +
b101111101100100 1
#408350000000
0#
0(
#408360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#408410000000
0$
0)
#408420000000
1"
1'
b0 +
b0 1
#408470000000
0"
0'
#408480000000
1#
1(
b101111101100100 +
b101111101100100 1
#408530000000
0#
0(
#408540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#408590000000
0$
0)
#408600000000
1"
1'
b0 +
b0 1
#408650000000
0"
0'
#408660000000
1#
1(
b101111101100100 +
b101111101100100 1
#408710000000
0#
0(
#408720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#408770000000
0$
0)
#408780000000
1"
1'
b0 +
b0 1
#408830000000
0"
0'
#408840000000
1#
1(
b101111101100100 +
b101111101100100 1
#408890000000
0#
0(
#408900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#408950000000
0$
0)
#408960000000
1"
1'
b0 +
b0 1
#409010000000
0"
0'
#409020000000
1#
1(
b101111101100100 +
b101111101100100 1
#409070000000
0#
0(
#409080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#409130000000
0$
0)
#409140000000
1"
1'
b0 +
b0 1
#409190000000
0"
0'
#409200000000
1#
1(
b101111101100100 +
b101111101100100 1
#409250000000
0#
0(
#409260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#409310000000
0$
0)
#409320000000
1"
1'
b0 +
b0 1
#409370000000
0"
0'
#409380000000
1#
1(
b101111101100100 +
b101111101100100 1
#409430000000
0#
0(
#409440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#409490000000
0$
0)
#409500000000
1"
1'
b0 +
b0 1
#409550000000
0"
0'
#409560000000
1#
1(
b101111101100100 +
b101111101100100 1
#409610000000
0#
0(
#409620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#409670000000
0$
0)
#409680000000
1"
1'
b0 +
b0 1
#409730000000
0"
0'
#409740000000
1#
1(
b101111101100100 +
b101111101100100 1
#409790000000
0#
0(
#409800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#409850000000
0$
0)
#409860000000
1"
1'
b0 +
b0 1
#409910000000
0"
0'
#409920000000
1#
1(
b101111101100100 +
b101111101100100 1
#409970000000
0#
0(
#409980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#410030000000
0$
0)
#410040000000
1"
1'
b0 +
b0 1
#410090000000
0"
0'
#410100000000
1#
1(
b101111101100100 +
b101111101100100 1
#410150000000
0#
0(
#410160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#410210000000
0$
0)
#410220000000
1"
1'
b0 +
b0 1
#410270000000
0"
0'
#410280000000
1#
1(
b101111101100100 +
b101111101100100 1
#410330000000
0#
0(
#410340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#410390000000
0$
0)
#410400000000
1"
1'
b0 +
b0 1
#410450000000
0"
0'
#410460000000
1#
1(
b101111101100100 +
b101111101100100 1
#410510000000
0#
0(
#410520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#410570000000
0$
0)
#410580000000
1"
1'
b0 +
b0 1
#410630000000
0"
0'
#410640000000
1#
1(
b101111101100100 +
b101111101100100 1
#410690000000
0#
0(
#410700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#410750000000
0$
0)
#410760000000
1"
1'
b0 +
b0 1
#410810000000
0"
0'
#410820000000
1#
1(
b101111101100100 +
b101111101100100 1
#410870000000
0#
0(
#410880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#410930000000
0$
0)
#410940000000
1"
1'
b0 +
b0 1
#410990000000
0"
0'
#411000000000
1#
1(
b101111101100100 +
b101111101100100 1
#411050000000
0#
0(
#411060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#411110000000
0$
0)
#411120000000
1"
1'
b0 +
b0 1
#411170000000
0"
0'
#411180000000
1#
1(
b101111101100100 +
b101111101100100 1
#411230000000
0#
0(
#411240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#411290000000
0$
0)
#411300000000
1"
1'
b0 +
b0 1
#411350000000
0"
0'
#411360000000
1#
1(
b101111101100100 +
b101111101100100 1
#411410000000
0#
0(
#411420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#411470000000
0$
0)
#411480000000
1"
1'
b0 +
b0 1
#411530000000
0"
0'
#411540000000
1#
1(
b101111101100100 +
b101111101100100 1
#411590000000
0#
0(
#411600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#411650000000
0$
0)
#411660000000
1"
1'
b0 +
b0 1
#411710000000
0"
0'
#411720000000
1#
1(
b101111101100100 +
b101111101100100 1
#411770000000
0#
0(
#411780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#411830000000
0$
0)
#411840000000
1"
1'
b0 +
b0 1
#411890000000
0"
0'
#411900000000
1#
1(
b101111101100100 +
b101111101100100 1
#411950000000
0#
0(
#411960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#412010000000
0$
0)
#412020000000
1"
1'
b0 +
b0 1
#412070000000
0"
0'
#412080000000
1#
1(
b101111101100100 +
b101111101100100 1
#412130000000
0#
0(
#412140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#412190000000
0$
0)
#412200000000
1"
1'
b0 +
b0 1
#412250000000
0"
0'
#412260000000
1#
1(
b101111101100100 +
b101111101100100 1
#412310000000
0#
0(
#412320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#412370000000
0$
0)
#412380000000
1"
1'
b0 +
b0 1
#412430000000
0"
0'
#412440000000
1#
1(
b101111101100100 +
b101111101100100 1
#412490000000
0#
0(
#412500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#412550000000
0$
0)
#412560000000
1"
1'
b0 +
b0 1
#412610000000
0"
0'
#412620000000
1#
1(
b101111101100100 +
b101111101100100 1
#412670000000
0#
0(
#412680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#412730000000
0$
0)
#412740000000
1"
1'
b0 +
b0 1
#412790000000
0"
0'
#412800000000
1#
1(
b101111101100100 +
b101111101100100 1
#412850000000
0#
0(
#412860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#412910000000
0$
0)
#412920000000
1"
1'
b0 +
b0 1
#412970000000
0"
0'
#412980000000
1#
1(
b101111101100100 +
b101111101100100 1
#413030000000
0#
0(
#413040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#413090000000
0$
0)
#413100000000
1"
1'
b0 +
b0 1
#413150000000
0"
0'
#413160000000
1#
1(
b101111101100100 +
b101111101100100 1
#413210000000
0#
0(
#413220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#413270000000
0$
0)
#413280000000
1"
1'
b0 +
b0 1
#413330000000
0"
0'
#413340000000
1#
1(
b101111101100100 +
b101111101100100 1
#413390000000
0#
0(
#413400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#413450000000
0$
0)
#413460000000
1"
1'
b0 +
b0 1
#413510000000
0"
0'
#413520000000
1#
1(
b101111101100100 +
b101111101100100 1
#413570000000
0#
0(
#413580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#413630000000
0$
0)
#413640000000
1"
1'
b0 +
b0 1
#413690000000
0"
0'
#413700000000
1#
1(
b101111101100100 +
b101111101100100 1
#413750000000
0#
0(
#413760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#413810000000
0$
0)
#413820000000
1"
1'
b0 +
b0 1
#413870000000
0"
0'
#413880000000
1#
1(
b101111101100100 +
b101111101100100 1
#413930000000
0#
0(
#413940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#413990000000
0$
0)
#414000000000
1"
1'
b0 +
b0 1
#414050000000
0"
0'
#414060000000
1#
1(
b101111101100100 +
b101111101100100 1
#414110000000
0#
0(
#414120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#414170000000
0$
0)
#414180000000
1"
1'
b0 +
b0 1
#414230000000
0"
0'
#414240000000
1#
1(
b101111101100100 +
b101111101100100 1
#414290000000
0#
0(
#414300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#414350000000
0$
0)
#414360000000
1"
1'
b0 +
b0 1
#414410000000
0"
0'
#414420000000
1#
1(
b101111101100100 +
b101111101100100 1
#414470000000
0#
0(
#414480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#414530000000
0$
0)
#414540000000
1"
1'
b0 +
b0 1
#414590000000
0"
0'
#414600000000
1#
1(
b101111101100100 +
b101111101100100 1
#414650000000
0#
0(
#414660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#414710000000
0$
0)
#414720000000
1"
1'
b0 +
b0 1
#414770000000
0"
0'
#414780000000
1#
1(
b101111101100100 +
b101111101100100 1
#414830000000
0#
0(
#414840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#414890000000
0$
0)
#414900000000
1"
1'
b0 +
b0 1
#414950000000
0"
0'
#414960000000
1#
1(
b101111101100100 +
b101111101100100 1
#415010000000
0#
0(
#415020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#415070000000
0$
0)
#415080000000
1"
1'
b0 +
b0 1
#415130000000
0"
0'
#415140000000
1#
1(
b101111101100100 +
b101111101100100 1
#415190000000
0#
0(
#415200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#415250000000
0$
0)
#415260000000
1"
1'
b0 +
b0 1
#415310000000
0"
0'
#415320000000
1#
1(
b101111101100100 +
b101111101100100 1
#415370000000
0#
0(
#415380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#415430000000
0$
0)
#415440000000
1"
1'
b0 +
b0 1
#415490000000
0"
0'
#415500000000
1#
1(
b101111101100100 +
b101111101100100 1
#415550000000
0#
0(
#415560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#415610000000
0$
0)
#415620000000
1"
1'
b0 +
b0 1
#415670000000
0"
0'
#415680000000
1#
1(
b101111101100100 +
b101111101100100 1
#415730000000
0#
0(
#415740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#415790000000
0$
0)
#415800000000
1"
1'
b0 +
b0 1
#415850000000
0"
0'
#415860000000
1#
1(
b101111101100100 +
b101111101100100 1
#415910000000
0#
0(
#415920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#415970000000
0$
0)
#415980000000
1"
1'
b0 +
b0 1
#416030000000
0"
0'
#416040000000
1#
1(
b101111101100100 +
b101111101100100 1
#416090000000
0#
0(
#416100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#416150000000
0$
0)
#416160000000
1"
1'
b0 +
b0 1
#416210000000
0"
0'
#416220000000
1#
1(
b101111101100100 +
b101111101100100 1
#416270000000
0#
0(
#416280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#416330000000
0$
0)
#416340000000
1"
1'
b0 +
b0 1
#416390000000
0"
0'
#416400000000
1#
1(
b101111101100100 +
b101111101100100 1
#416450000000
0#
0(
#416460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#416510000000
0$
0)
#416520000000
1"
1'
b0 +
b0 1
#416570000000
0"
0'
#416580000000
1#
1(
b101111101100100 +
b101111101100100 1
#416630000000
0#
0(
#416640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#416690000000
0$
0)
#416700000000
1"
1'
b0 +
b0 1
#416750000000
0"
0'
#416760000000
1#
1(
b101111101100100 +
b101111101100100 1
#416810000000
0#
0(
#416820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#416870000000
0$
0)
#416880000000
1"
1'
b0 +
b0 1
#416930000000
0"
0'
#416940000000
1#
1(
b101111101100100 +
b101111101100100 1
#416990000000
0#
0(
#417000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#417050000000
0$
0)
#417060000000
1"
1'
b0 +
b0 1
#417110000000
0"
0'
#417120000000
1#
1(
b101111101100100 +
b101111101100100 1
#417170000000
0#
0(
#417180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#417230000000
0$
0)
#417240000000
1"
1'
b0 +
b0 1
#417290000000
0"
0'
#417300000000
1#
1(
b101111101100100 +
b101111101100100 1
#417350000000
0#
0(
#417360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#417410000000
0$
0)
#417420000000
1"
1'
b0 +
b0 1
#417470000000
0"
0'
#417480000000
1#
1(
b101111101100100 +
b101111101100100 1
#417530000000
0#
0(
#417540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#417590000000
0$
0)
#417600000000
1"
1'
b0 +
b0 1
#417650000000
0"
0'
#417660000000
1#
1(
b101111101100100 +
b101111101100100 1
#417710000000
0#
0(
#417720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#417770000000
0$
0)
#417780000000
1"
1'
b0 +
b0 1
#417830000000
0"
0'
#417840000000
1#
1(
b101111101100100 +
b101111101100100 1
#417890000000
0#
0(
#417900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#417950000000
0$
0)
#417960000000
1"
1'
b0 +
b0 1
#418010000000
0"
0'
#418020000000
1#
1(
b101111101100100 +
b101111101100100 1
#418070000000
0#
0(
#418080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#418130000000
0$
0)
#418140000000
1"
1'
b0 +
b0 1
#418190000000
0"
0'
#418200000000
1#
1(
b101111101100100 +
b101111101100100 1
#418250000000
0#
0(
#418260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#418310000000
0$
0)
#418320000000
1"
1'
b0 +
b0 1
#418370000000
0"
0'
#418380000000
1#
1(
b101111101100100 +
b101111101100100 1
#418430000000
0#
0(
#418440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#418490000000
0$
0)
#418500000000
1"
1'
b0 +
b0 1
#418550000000
0"
0'
#418560000000
1#
1(
b101111101100100 +
b101111101100100 1
#418610000000
0#
0(
#418620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#418670000000
0$
0)
#418680000000
1"
1'
b0 +
b0 1
#418730000000
0"
0'
#418740000000
1#
1(
b101111101100100 +
b101111101100100 1
#418790000000
0#
0(
#418800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#418850000000
0$
0)
#418860000000
1"
1'
b0 +
b0 1
#418910000000
0"
0'
#418920000000
1#
1(
b101111101100100 +
b101111101100100 1
#418970000000
0#
0(
#418980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#419030000000
0$
0)
#419040000000
1"
1'
b0 +
b0 1
#419090000000
0"
0'
#419100000000
1#
1(
b101111101100100 +
b101111101100100 1
#419150000000
0#
0(
#419160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#419210000000
0$
0)
#419220000000
1"
1'
b0 +
b0 1
#419270000000
0"
0'
#419280000000
1#
1(
b101111101100100 +
b101111101100100 1
#419330000000
0#
0(
#419340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#419390000000
0$
0)
#419400000000
1"
1'
b0 +
b0 1
#419450000000
0"
0'
#419460000000
1#
1(
b101111101100100 +
b101111101100100 1
#419510000000
0#
0(
#419520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#419570000000
0$
0)
#419580000000
1"
1'
b0 +
b0 1
#419630000000
0"
0'
#419640000000
1#
1(
b101111101100100 +
b101111101100100 1
#419690000000
0#
0(
#419700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#419750000000
0$
0)
#419760000000
1"
1'
b0 +
b0 1
#419810000000
0"
0'
#419820000000
1#
1(
b101111101100100 +
b101111101100100 1
#419870000000
0#
0(
#419880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#419930000000
0$
0)
#419940000000
1"
1'
b0 +
b0 1
#419990000000
0"
0'
#420000000000
1#
1(
b101111101100100 +
b101111101100100 1
#420050000000
0#
0(
#420060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#420110000000
0$
0)
#420120000000
1"
1'
b0 +
b0 1
#420170000000
0"
0'
#420180000000
1#
1(
b101111101100100 +
b101111101100100 1
#420230000000
0#
0(
#420240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#420290000000
0$
0)
#420300000000
1"
1'
b0 +
b0 1
#420350000000
0"
0'
#420360000000
1#
1(
b101111101100100 +
b101111101100100 1
#420410000000
0#
0(
#420420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#420470000000
0$
0)
#420480000000
1"
1'
b0 +
b0 1
#420530000000
0"
0'
#420540000000
1#
1(
b101111101100100 +
b101111101100100 1
#420590000000
0#
0(
#420600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#420650000000
0$
0)
#420660000000
1"
1'
b0 +
b0 1
#420710000000
0"
0'
#420720000000
1#
1(
b101111101100100 +
b101111101100100 1
#420770000000
0#
0(
#420780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#420830000000
0$
0)
#420840000000
1"
1'
b0 +
b0 1
#420890000000
0"
0'
#420900000000
1#
1(
b101111101100100 +
b101111101100100 1
#420950000000
0#
0(
#420960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#421010000000
0$
0)
#421020000000
1"
1'
b0 +
b0 1
#421070000000
0"
0'
#421080000000
1#
1(
b101111101100100 +
b101111101100100 1
#421130000000
0#
0(
#421140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#421190000000
0$
0)
#421200000000
1"
1'
b0 +
b0 1
#421250000000
0"
0'
#421260000000
1#
1(
b101111101100100 +
b101111101100100 1
#421310000000
0#
0(
#421320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#421370000000
0$
0)
#421380000000
1"
1'
b0 +
b0 1
#421430000000
0"
0'
#421440000000
1#
1(
b101111101100100 +
b101111101100100 1
#421490000000
0#
0(
#421500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#421550000000
0$
0)
#421560000000
1"
1'
b0 +
b0 1
#421610000000
0"
0'
#421620000000
1#
1(
b101111101100100 +
b101111101100100 1
#421670000000
0#
0(
#421680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#421730000000
0$
0)
#421740000000
1"
1'
b0 +
b0 1
#421790000000
0"
0'
#421800000000
1#
1(
b101111101100100 +
b101111101100100 1
#421850000000
0#
0(
#421860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#421910000000
0$
0)
#421920000000
1"
1'
b0 +
b0 1
#421970000000
0"
0'
#421980000000
1#
1(
b101111101100100 +
b101111101100100 1
#422030000000
0#
0(
#422040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#422090000000
0$
0)
#422100000000
1"
1'
b0 +
b0 1
#422150000000
0"
0'
#422160000000
1#
1(
b101111101100100 +
b101111101100100 1
#422210000000
0#
0(
#422220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#422270000000
0$
0)
#422280000000
1"
1'
b0 +
b0 1
#422330000000
0"
0'
#422340000000
1#
1(
b101111101100100 +
b101111101100100 1
#422390000000
0#
0(
#422400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#422450000000
0$
0)
#422460000000
1"
1'
b0 +
b0 1
#422510000000
0"
0'
#422520000000
1#
1(
b101111101100100 +
b101111101100100 1
#422570000000
0#
0(
#422580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#422630000000
0$
0)
#422640000000
1"
1'
b0 +
b0 1
#422690000000
0"
0'
#422700000000
1#
1(
b101111101100100 +
b101111101100100 1
#422750000000
0#
0(
#422760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#422810000000
0$
0)
#422820000000
1"
1'
b0 +
b0 1
#422870000000
0"
0'
#422880000000
1#
1(
b101111101100100 +
b101111101100100 1
#422930000000
0#
0(
#422940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#422990000000
0$
0)
#423000000000
1"
1'
b0 +
b0 1
#423050000000
0"
0'
#423060000000
1#
1(
b101111101100100 +
b101111101100100 1
#423110000000
0#
0(
#423120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#423170000000
0$
0)
#423180000000
1"
1'
b0 +
b0 1
#423230000000
0"
0'
#423240000000
1#
1(
b101111101100100 +
b101111101100100 1
#423290000000
0#
0(
#423300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#423350000000
0$
0)
#423360000000
1"
1'
b0 +
b0 1
#423410000000
0"
0'
#423420000000
1#
1(
b101111101100100 +
b101111101100100 1
#423470000000
0#
0(
#423480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#423530000000
0$
0)
#423540000000
1"
1'
b0 +
b0 1
#423590000000
0"
0'
#423600000000
1#
1(
b101111101100100 +
b101111101100100 1
#423650000000
0#
0(
#423660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#423710000000
0$
0)
#423720000000
1"
1'
b0 +
b0 1
#423770000000
0"
0'
#423780000000
1#
1(
b101111101100100 +
b101111101100100 1
#423830000000
0#
0(
#423840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#423890000000
0$
0)
#423900000000
1"
1'
b0 +
b0 1
#423950000000
0"
0'
#423960000000
1#
1(
b101111101100100 +
b101111101100100 1
#424010000000
0#
0(
#424020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#424070000000
0$
0)
#424080000000
1"
1'
b0 +
b0 1
#424130000000
0"
0'
#424140000000
1#
1(
b101111101100100 +
b101111101100100 1
#424190000000
0#
0(
#424200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#424250000000
0$
0)
#424260000000
1"
1'
b0 +
b0 1
#424310000000
0"
0'
#424320000000
1#
1(
b101111101100100 +
b101111101100100 1
#424370000000
0#
0(
#424380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#424430000000
0$
0)
#424440000000
1"
1'
b0 +
b0 1
#424490000000
0"
0'
#424500000000
1#
1(
b101111101100100 +
b101111101100100 1
#424550000000
0#
0(
#424560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#424610000000
0$
0)
#424620000000
1"
1'
b0 +
b0 1
#424670000000
0"
0'
#424680000000
1#
1(
b101111101100100 +
b101111101100100 1
#424730000000
0#
0(
#424740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#424790000000
0$
0)
#424800000000
1"
1'
b0 +
b0 1
#424850000000
0"
0'
#424860000000
1#
1(
b101111101100100 +
b101111101100100 1
#424910000000
0#
0(
#424920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#424970000000
0$
0)
#424980000000
1"
1'
b0 +
b0 1
#425030000000
0"
0'
#425040000000
1#
1(
b101111101100100 +
b101111101100100 1
#425090000000
0#
0(
#425100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#425150000000
0$
0)
#425160000000
1"
1'
b0 +
b0 1
#425210000000
0"
0'
#425220000000
1#
1(
b101111101100100 +
b101111101100100 1
#425270000000
0#
0(
#425280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#425330000000
0$
0)
#425340000000
1"
1'
b0 +
b0 1
#425390000000
0"
0'
#425400000000
1#
1(
b101111101100100 +
b101111101100100 1
#425450000000
0#
0(
#425460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#425510000000
0$
0)
#425520000000
1"
1'
b0 +
b0 1
#425570000000
0"
0'
#425580000000
1#
1(
b101111101100100 +
b101111101100100 1
#425630000000
0#
0(
#425640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#425690000000
0$
0)
#425700000000
1"
1'
b0 +
b0 1
#425750000000
0"
0'
#425760000000
1#
1(
b101111101100100 +
b101111101100100 1
#425810000000
0#
0(
#425820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#425870000000
0$
0)
#425880000000
1"
1'
b0 +
b0 1
#425930000000
0"
0'
#425940000000
1#
1(
b101111101100100 +
b101111101100100 1
#425990000000
0#
0(
#426000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#426050000000
0$
0)
#426060000000
1"
1'
b0 +
b0 1
#426110000000
0"
0'
#426120000000
1#
1(
b101111101100100 +
b101111101100100 1
#426170000000
0#
0(
#426180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#426230000000
0$
0)
#426240000000
1"
1'
b0 +
b0 1
#426290000000
0"
0'
#426300000000
1#
1(
b101111101100100 +
b101111101100100 1
#426350000000
0#
0(
#426360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#426410000000
0$
0)
#426420000000
1"
1'
b0 +
b0 1
#426470000000
0"
0'
#426480000000
1#
1(
b101111101100100 +
b101111101100100 1
#426530000000
0#
0(
#426540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#426590000000
0$
0)
#426600000000
1"
1'
b0 +
b0 1
#426650000000
0"
0'
#426660000000
1#
1(
b101111101100100 +
b101111101100100 1
#426710000000
0#
0(
#426720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#426770000000
0$
0)
#426780000000
1"
1'
b0 +
b0 1
#426830000000
0"
0'
#426840000000
1#
1(
b101111101100100 +
b101111101100100 1
#426890000000
0#
0(
#426900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#426950000000
0$
0)
#426960000000
1"
1'
b0 +
b0 1
#427010000000
0"
0'
#427020000000
1#
1(
b101111101100100 +
b101111101100100 1
#427070000000
0#
0(
#427080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#427130000000
0$
0)
#427140000000
1"
1'
b0 +
b0 1
#427190000000
0"
0'
#427200000000
1#
1(
b101111101100100 +
b101111101100100 1
#427250000000
0#
0(
#427260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#427310000000
0$
0)
#427320000000
1"
1'
b0 +
b0 1
#427370000000
0"
0'
#427380000000
1#
1(
b101111101100100 +
b101111101100100 1
#427430000000
0#
0(
#427440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#427490000000
0$
0)
#427500000000
1"
1'
b0 +
b0 1
#427550000000
0"
0'
#427560000000
1#
1(
b101111101100100 +
b101111101100100 1
#427610000000
0#
0(
#427620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#427670000000
0$
0)
#427680000000
1"
1'
b0 +
b0 1
#427730000000
0"
0'
#427740000000
1#
1(
b101111101100100 +
b101111101100100 1
#427790000000
0#
0(
#427800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#427850000000
0$
0)
#427860000000
1"
1'
b0 +
b0 1
#427910000000
0"
0'
#427920000000
1#
1(
b101111101100100 +
b101111101100100 1
#427970000000
0#
0(
#427980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#428030000000
0$
0)
#428040000000
1"
1'
b0 +
b0 1
#428090000000
0"
0'
#428100000000
1#
1(
b101111101100100 +
b101111101100100 1
#428150000000
0#
0(
#428160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#428210000000
0$
0)
#428220000000
1"
1'
b0 +
b0 1
#428270000000
0"
0'
#428280000000
1#
1(
b101111101100100 +
b101111101100100 1
#428330000000
0#
0(
#428340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#428390000000
0$
0)
#428400000000
1"
1'
b0 +
b0 1
#428450000000
0"
0'
#428460000000
1#
1(
b101111101100100 +
b101111101100100 1
#428510000000
0#
0(
#428520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#428570000000
0$
0)
#428580000000
1"
1'
b0 +
b0 1
#428630000000
0"
0'
#428640000000
1#
1(
b101111101100100 +
b101111101100100 1
#428690000000
0#
0(
#428700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#428750000000
0$
0)
#428760000000
1"
1'
b0 +
b0 1
#428810000000
0"
0'
#428820000000
1#
1(
b101111101100100 +
b101111101100100 1
#428870000000
0#
0(
#428880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#428930000000
0$
0)
#428940000000
1"
1'
b0 +
b0 1
#428990000000
0"
0'
#429000000000
1#
1(
b101111101100100 +
b101111101100100 1
#429050000000
0#
0(
#429060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#429110000000
0$
0)
#429120000000
1"
1'
b0 +
b0 1
#429170000000
0"
0'
#429180000000
1#
1(
b101111101100100 +
b101111101100100 1
#429230000000
0#
0(
#429240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#429290000000
0$
0)
#429300000000
1"
1'
b0 +
b0 1
#429350000000
0"
0'
#429360000000
1#
1(
b101111101100100 +
b101111101100100 1
#429410000000
0#
0(
#429420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#429470000000
0$
0)
#429480000000
1"
1'
b0 +
b0 1
#429530000000
0"
0'
#429540000000
1#
1(
b101111101100100 +
b101111101100100 1
#429590000000
0#
0(
#429600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#429650000000
0$
0)
#429660000000
1"
1'
b0 +
b0 1
#429710000000
0"
0'
#429720000000
1#
1(
b101111101100100 +
b101111101100100 1
#429770000000
0#
0(
#429780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#429830000000
0$
0)
#429840000000
1"
1'
b0 +
b0 1
#429890000000
0"
0'
#429900000000
1#
1(
b101111101100100 +
b101111101100100 1
#429950000000
0#
0(
#429960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#430010000000
0$
0)
#430020000000
1"
1'
b0 +
b0 1
#430070000000
0"
0'
#430080000000
1#
1(
b101111101100100 +
b101111101100100 1
#430130000000
0#
0(
#430140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#430190000000
0$
0)
#430200000000
1"
1'
b0 +
b0 1
#430250000000
0"
0'
#430260000000
1#
1(
b101111101100100 +
b101111101100100 1
#430310000000
0#
0(
#430320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#430370000000
0$
0)
#430380000000
1"
1'
b0 +
b0 1
#430430000000
0"
0'
#430440000000
1#
1(
b101111101100100 +
b101111101100100 1
#430490000000
0#
0(
#430500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#430550000000
0$
0)
#430560000000
1"
1'
b0 +
b0 1
#430610000000
0"
0'
#430620000000
1#
1(
b101111101100100 +
b101111101100100 1
#430670000000
0#
0(
#430680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#430730000000
0$
0)
#430740000000
1"
1'
b0 +
b0 1
#430790000000
0"
0'
#430800000000
1#
1(
b101111101100100 +
b101111101100100 1
#430850000000
0#
0(
#430860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#430910000000
0$
0)
#430920000000
1"
1'
b0 +
b0 1
#430970000000
0"
0'
#430980000000
1#
1(
b101111101100100 +
b101111101100100 1
#431030000000
0#
0(
#431040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#431090000000
0$
0)
#431100000000
1"
1'
b0 +
b0 1
#431150000000
0"
0'
#431160000000
1#
1(
b101111101100100 +
b101111101100100 1
#431210000000
0#
0(
#431220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#431270000000
0$
0)
#431280000000
1"
1'
b0 +
b0 1
#431330000000
0"
0'
#431340000000
1#
1(
b101111101100100 +
b101111101100100 1
#431390000000
0#
0(
#431400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#431450000000
0$
0)
#431460000000
1"
1'
b0 +
b0 1
#431510000000
0"
0'
#431520000000
1#
1(
b101111101100100 +
b101111101100100 1
#431570000000
0#
0(
#431580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#431630000000
0$
0)
#431640000000
1"
1'
b0 +
b0 1
#431690000000
0"
0'
#431700000000
1#
1(
b101111101100100 +
b101111101100100 1
#431750000000
0#
0(
#431760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#431810000000
0$
0)
#431820000000
1"
1'
b0 +
b0 1
#431870000000
0"
0'
#431880000000
1#
1(
b101111101100100 +
b101111101100100 1
#431930000000
0#
0(
#431940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#431990000000
0$
0)
#432000000000
1"
1'
b0 +
b0 1
#432050000000
0"
0'
#432060000000
1#
1(
b101111101100100 +
b101111101100100 1
#432110000000
0#
0(
#432120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#432170000000
0$
0)
#432180000000
1"
1'
b0 +
b0 1
#432230000000
0"
0'
#432240000000
1#
1(
b101111101100100 +
b101111101100100 1
#432290000000
0#
0(
#432300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#432350000000
0$
0)
#432360000000
1"
1'
b0 +
b0 1
#432410000000
0"
0'
#432420000000
1#
1(
b101111101100100 +
b101111101100100 1
#432470000000
0#
0(
#432480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#432530000000
0$
0)
#432540000000
1"
1'
b0 +
b0 1
#432590000000
0"
0'
#432600000000
1#
1(
b101111101100100 +
b101111101100100 1
#432650000000
0#
0(
#432660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#432710000000
0$
0)
#432720000000
1"
1'
b0 +
b0 1
#432770000000
0"
0'
#432780000000
1#
1(
b101111101100100 +
b101111101100100 1
#432830000000
0#
0(
#432840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#432890000000
0$
0)
#432900000000
1"
1'
b0 +
b0 1
#432950000000
0"
0'
#432960000000
1#
1(
b101111101100100 +
b101111101100100 1
#433010000000
0#
0(
#433020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#433070000000
0$
0)
#433080000000
1"
1'
b0 +
b0 1
#433130000000
0"
0'
#433140000000
1#
1(
b101111101100100 +
b101111101100100 1
#433190000000
0#
0(
#433200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#433250000000
0$
0)
#433260000000
1"
1'
b0 +
b0 1
#433310000000
0"
0'
#433320000000
1#
1(
b101111101100100 +
b101111101100100 1
#433370000000
0#
0(
#433380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#433430000000
0$
0)
#433440000000
1"
1'
b0 +
b0 1
#433490000000
0"
0'
#433500000000
1#
1(
b101111101100100 +
b101111101100100 1
#433550000000
0#
0(
#433560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#433610000000
0$
0)
#433620000000
1"
1'
b0 +
b0 1
#433670000000
0"
0'
#433680000000
1#
1(
b101111101100100 +
b101111101100100 1
#433730000000
0#
0(
#433740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#433790000000
0$
0)
#433800000000
1"
1'
b0 +
b0 1
#433850000000
0"
0'
#433860000000
1#
1(
b101111101100100 +
b101111101100100 1
#433910000000
0#
0(
#433920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#433970000000
0$
0)
#433980000000
1"
1'
b0 +
b0 1
#434030000000
0"
0'
#434040000000
1#
1(
b101111101100100 +
b101111101100100 1
#434090000000
0#
0(
#434100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#434150000000
0$
0)
#434160000000
1"
1'
b0 +
b0 1
#434210000000
0"
0'
#434220000000
1#
1(
b101111101100100 +
b101111101100100 1
#434270000000
0#
0(
#434280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#434330000000
0$
0)
#434340000000
1"
1'
b0 +
b0 1
#434390000000
0"
0'
#434400000000
1#
1(
b101111101100100 +
b101111101100100 1
#434450000000
0#
0(
#434460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#434510000000
0$
0)
#434520000000
1"
1'
b0 +
b0 1
#434570000000
0"
0'
#434580000000
1#
1(
b101111101100100 +
b101111101100100 1
#434630000000
0#
0(
#434640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#434690000000
0$
0)
#434700000000
1"
1'
b0 +
b0 1
#434750000000
0"
0'
#434760000000
1#
1(
b101111101100100 +
b101111101100100 1
#434810000000
0#
0(
#434820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#434870000000
0$
0)
#434880000000
1"
1'
b0 +
b0 1
#434930000000
0"
0'
#434940000000
1#
1(
b101111101100100 +
b101111101100100 1
#434990000000
0#
0(
#435000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#435050000000
0$
0)
#435060000000
1"
1'
b0 +
b0 1
#435110000000
0"
0'
#435120000000
1#
1(
b101111101100100 +
b101111101100100 1
#435170000000
0#
0(
#435180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#435230000000
0$
0)
#435240000000
1"
1'
b0 +
b0 1
#435290000000
0"
0'
#435300000000
1#
1(
b101111101100100 +
b101111101100100 1
#435350000000
0#
0(
#435360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#435410000000
0$
0)
#435420000000
1"
1'
b0 +
b0 1
#435470000000
0"
0'
#435480000000
1#
1(
b101111101100100 +
b101111101100100 1
#435530000000
0#
0(
#435540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#435590000000
0$
0)
#435600000000
1"
1'
b0 +
b0 1
#435650000000
0"
0'
#435660000000
1#
1(
b101111101100100 +
b101111101100100 1
#435710000000
0#
0(
#435720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#435770000000
0$
0)
#435780000000
1"
1'
b0 +
b0 1
#435830000000
0"
0'
#435840000000
1#
1(
b101111101100100 +
b101111101100100 1
#435890000000
0#
0(
#435900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#435950000000
0$
0)
#435960000000
1"
1'
b0 +
b0 1
#436010000000
0"
0'
#436020000000
1#
1(
b101111101100100 +
b101111101100100 1
#436070000000
0#
0(
#436080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#436130000000
0$
0)
#436140000000
1"
1'
b0 +
b0 1
#436190000000
0"
0'
#436200000000
1#
1(
b101111101100100 +
b101111101100100 1
#436250000000
0#
0(
#436260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#436310000000
0$
0)
#436320000000
1"
1'
b0 +
b0 1
#436370000000
0"
0'
#436380000000
1#
1(
b101111101100100 +
b101111101100100 1
#436430000000
0#
0(
#436440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#436490000000
0$
0)
#436500000000
1"
1'
b0 +
b0 1
#436550000000
0"
0'
#436560000000
1#
1(
b101111101100100 +
b101111101100100 1
#436610000000
0#
0(
#436620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#436670000000
0$
0)
#436680000000
1"
1'
b0 +
b0 1
#436730000000
0"
0'
#436740000000
1#
1(
b101111101100100 +
b101111101100100 1
#436790000000
0#
0(
#436800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#436850000000
0$
0)
#436860000000
1"
1'
b0 +
b0 1
#436910000000
0"
0'
#436920000000
1#
1(
b101111101100100 +
b101111101100100 1
#436970000000
0#
0(
#436980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#437030000000
0$
0)
#437040000000
1"
1'
b0 +
b0 1
#437090000000
0"
0'
#437100000000
1#
1(
b101111101100100 +
b101111101100100 1
#437150000000
0#
0(
#437160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#437210000000
0$
0)
#437220000000
1"
1'
b0 +
b0 1
#437270000000
0"
0'
#437280000000
1#
1(
b101111101100100 +
b101111101100100 1
#437330000000
0#
0(
#437340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#437390000000
0$
0)
#437400000000
1"
1'
b0 +
b0 1
#437450000000
0"
0'
#437460000000
1#
1(
b101111101100100 +
b101111101100100 1
#437510000000
0#
0(
#437520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#437570000000
0$
0)
#437580000000
1"
1'
b0 +
b0 1
#437630000000
0"
0'
#437640000000
1#
1(
b101111101100100 +
b101111101100100 1
#437690000000
0#
0(
#437700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#437750000000
0$
0)
#437760000000
1"
1'
b0 +
b0 1
#437810000000
0"
0'
#437820000000
1#
1(
b101111101100100 +
b101111101100100 1
#437870000000
0#
0(
#437880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#437930000000
0$
0)
#437940000000
1"
1'
b0 +
b0 1
#437990000000
0"
0'
#438000000000
1#
1(
b101111101100100 +
b101111101100100 1
#438050000000
0#
0(
#438060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#438110000000
0$
0)
#438120000000
1"
1'
b0 +
b0 1
#438170000000
0"
0'
#438180000000
1#
1(
b101111101100100 +
b101111101100100 1
#438230000000
0#
0(
#438240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#438290000000
0$
0)
#438300000000
1"
1'
b0 +
b0 1
#438350000000
0"
0'
#438360000000
1#
1(
b101111101100100 +
b101111101100100 1
#438410000000
0#
0(
#438420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#438470000000
0$
0)
#438480000000
1"
1'
b0 +
b0 1
#438530000000
0"
0'
#438540000000
1#
1(
b101111101100100 +
b101111101100100 1
#438590000000
0#
0(
#438600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#438650000000
0$
0)
#438660000000
1"
1'
b0 +
b0 1
#438710000000
0"
0'
#438720000000
1#
1(
b101111101100100 +
b101111101100100 1
#438770000000
0#
0(
#438780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#438830000000
0$
0)
#438840000000
1"
1'
b0 +
b0 1
#438890000000
0"
0'
#438900000000
1#
1(
b101111101100100 +
b101111101100100 1
#438950000000
0#
0(
#438960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#439010000000
0$
0)
#439020000000
1"
1'
b0 +
b0 1
#439070000000
0"
0'
#439080000000
1#
1(
b101111101100100 +
b101111101100100 1
#439130000000
0#
0(
#439140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#439190000000
0$
0)
#439200000000
1"
1'
b0 +
b0 1
#439250000000
0"
0'
#439260000000
1#
1(
b101111101100100 +
b101111101100100 1
#439310000000
0#
0(
#439320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#439370000000
0$
0)
#439380000000
1"
1'
b0 +
b0 1
#439430000000
0"
0'
#439440000000
1#
1(
b101111101100100 +
b101111101100100 1
#439490000000
0#
0(
#439500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#439550000000
0$
0)
#439560000000
1"
1'
b0 +
b0 1
#439610000000
0"
0'
#439620000000
1#
1(
b101111101100100 +
b101111101100100 1
#439670000000
0#
0(
#439680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#439730000000
0$
0)
#439740000000
1"
1'
b0 +
b0 1
#439790000000
0"
0'
#439800000000
1#
1(
b101111101100100 +
b101111101100100 1
#439850000000
0#
0(
#439860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#439910000000
0$
0)
#439920000000
1"
1'
b0 +
b0 1
#439970000000
0"
0'
#439980000000
1#
1(
b101111101100100 +
b101111101100100 1
#440030000000
0#
0(
#440040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#440090000000
0$
0)
#440100000000
1"
1'
b0 +
b0 1
#440150000000
0"
0'
#440160000000
1#
1(
b101111101100100 +
b101111101100100 1
#440210000000
0#
0(
#440220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#440270000000
0$
0)
#440280000000
1"
1'
b0 +
b0 1
#440330000000
0"
0'
#440340000000
1#
1(
b101111101100100 +
b101111101100100 1
#440390000000
0#
0(
#440400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#440450000000
0$
0)
#440460000000
1"
1'
b0 +
b0 1
#440510000000
0"
0'
#440520000000
1#
1(
b101111101100100 +
b101111101100100 1
#440570000000
0#
0(
#440580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#440630000000
0$
0)
#440640000000
1"
1'
b0 +
b0 1
#440690000000
0"
0'
#440700000000
1#
1(
b101111101100100 +
b101111101100100 1
#440750000000
0#
0(
#440760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#440810000000
0$
0)
#440820000000
1"
1'
b0 +
b0 1
#440870000000
0"
0'
#440880000000
1#
1(
b101111101100100 +
b101111101100100 1
#440930000000
0#
0(
#440940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#440990000000
0$
0)
#441000000000
1"
1'
b0 +
b0 1
#441050000000
0"
0'
#441060000000
1#
1(
b101111101100100 +
b101111101100100 1
#441110000000
0#
0(
#441120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#441170000000
0$
0)
#441180000000
1"
1'
b0 +
b0 1
#441230000000
0"
0'
#441240000000
1#
1(
b101111101100100 +
b101111101100100 1
#441290000000
0#
0(
#441300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#441350000000
0$
0)
#441360000000
1"
1'
b0 +
b0 1
#441410000000
0"
0'
#441420000000
1#
1(
b101111101100100 +
b101111101100100 1
#441470000000
0#
0(
#441480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#441530000000
0$
0)
#441540000000
1"
1'
b0 +
b0 1
#441590000000
0"
0'
#441600000000
1#
1(
b101111101100100 +
b101111101100100 1
#441650000000
0#
0(
#441660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#441710000000
0$
0)
#441720000000
1"
1'
b0 +
b0 1
#441770000000
0"
0'
#441780000000
1#
1(
b101111101100100 +
b101111101100100 1
#441830000000
0#
0(
#441840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#441890000000
0$
0)
#441900000000
1"
1'
b0 +
b0 1
#441950000000
0"
0'
#441960000000
1#
1(
b101111101100100 +
b101111101100100 1
#442010000000
0#
0(
#442020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#442070000000
0$
0)
#442080000000
1"
1'
b0 +
b0 1
#442130000000
0"
0'
#442140000000
1#
1(
b101111101100100 +
b101111101100100 1
#442190000000
0#
0(
#442200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#442250000000
0$
0)
#442260000000
1"
1'
b0 +
b0 1
#442310000000
0"
0'
#442320000000
1#
1(
b101111101100100 +
b101111101100100 1
#442370000000
0#
0(
#442380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#442430000000
0$
0)
#442440000000
1"
1'
b0 +
b0 1
#442490000000
0"
0'
#442500000000
1#
1(
b101111101100100 +
b101111101100100 1
#442550000000
0#
0(
#442560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#442610000000
0$
0)
#442620000000
1"
1'
b0 +
b0 1
#442670000000
0"
0'
#442680000000
1#
1(
b101111101100100 +
b101111101100100 1
#442730000000
0#
0(
#442740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#442790000000
0$
0)
#442800000000
1"
1'
b0 +
b0 1
#442850000000
0"
0'
#442860000000
1#
1(
b101111101100100 +
b101111101100100 1
#442910000000
0#
0(
#442920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#442970000000
0$
0)
#442980000000
1"
1'
b0 +
b0 1
#443030000000
0"
0'
#443040000000
1#
1(
b101111101100100 +
b101111101100100 1
#443090000000
0#
0(
#443100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#443150000000
0$
0)
#443160000000
1"
1'
b0 +
b0 1
#443210000000
0"
0'
#443220000000
1#
1(
b101111101100100 +
b101111101100100 1
#443270000000
0#
0(
#443280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#443330000000
0$
0)
#443340000000
1"
1'
b0 +
b0 1
#443390000000
0"
0'
#443400000000
1#
1(
b101111101100100 +
b101111101100100 1
#443450000000
0#
0(
#443460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#443510000000
0$
0)
#443520000000
1"
1'
b0 +
b0 1
#443570000000
0"
0'
#443580000000
1#
1(
b101111101100100 +
b101111101100100 1
#443630000000
0#
0(
#443640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#443690000000
0$
0)
#443700000000
1"
1'
b0 +
b0 1
#443750000000
0"
0'
#443760000000
1#
1(
b101111101100100 +
b101111101100100 1
#443810000000
0#
0(
#443820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#443870000000
0$
0)
#443880000000
1"
1'
b0 +
b0 1
#443930000000
0"
0'
#443940000000
1#
1(
b101111101100100 +
b101111101100100 1
#443990000000
0#
0(
#444000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#444050000000
0$
0)
#444060000000
1"
1'
b0 +
b0 1
#444110000000
0"
0'
#444120000000
1#
1(
b101111101100100 +
b101111101100100 1
#444170000000
0#
0(
#444180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#444230000000
0$
0)
#444240000000
1"
1'
b0 +
b0 1
#444290000000
0"
0'
#444300000000
1#
1(
b101111101100100 +
b101111101100100 1
#444350000000
0#
0(
#444360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#444410000000
0$
0)
#444420000000
1"
1'
b0 +
b0 1
#444470000000
0"
0'
#444480000000
1#
1(
b101111101100100 +
b101111101100100 1
#444530000000
0#
0(
#444540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#444590000000
0$
0)
#444600000000
1"
1'
b0 +
b0 1
#444650000000
0"
0'
#444660000000
1#
1(
b101111101100100 +
b101111101100100 1
#444710000000
0#
0(
#444720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#444770000000
0$
0)
#444780000000
1"
1'
b0 +
b0 1
#444830000000
0"
0'
#444840000000
1#
1(
b101111101100100 +
b101111101100100 1
#444890000000
0#
0(
#444900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#444950000000
0$
0)
#444960000000
1"
1'
b0 +
b0 1
#445010000000
0"
0'
#445020000000
1#
1(
b101111101100100 +
b101111101100100 1
#445070000000
0#
0(
#445080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#445130000000
0$
0)
#445140000000
1"
1'
b0 +
b0 1
#445190000000
0"
0'
#445200000000
1#
1(
b101111101100100 +
b101111101100100 1
#445250000000
0#
0(
#445260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#445310000000
0$
0)
#445320000000
1"
1'
b0 +
b0 1
#445370000000
0"
0'
#445380000000
1#
1(
b101111101100100 +
b101111101100100 1
#445430000000
0#
0(
#445440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#445490000000
0$
0)
#445500000000
1"
1'
b0 +
b0 1
#445550000000
0"
0'
#445560000000
1#
1(
b101111101100100 +
b101111101100100 1
#445610000000
0#
0(
#445620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#445670000000
0$
0)
#445680000000
1"
1'
b0 +
b0 1
#445730000000
0"
0'
#445740000000
1#
1(
b101111101100100 +
b101111101100100 1
#445790000000
0#
0(
#445800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#445850000000
0$
0)
#445860000000
1"
1'
b0 +
b0 1
#445910000000
0"
0'
#445920000000
1#
1(
b101111101100100 +
b101111101100100 1
#445970000000
0#
0(
#445980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#446030000000
0$
0)
#446040000000
1"
1'
b0 +
b0 1
#446090000000
0"
0'
#446100000000
1#
1(
b101111101100100 +
b101111101100100 1
#446150000000
0#
0(
#446160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#446210000000
0$
0)
#446220000000
1"
1'
b0 +
b0 1
#446270000000
0"
0'
#446280000000
1#
1(
b101111101100100 +
b101111101100100 1
#446330000000
0#
0(
#446340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#446390000000
0$
0)
#446400000000
1"
1'
b0 +
b0 1
#446450000000
0"
0'
#446460000000
1#
1(
b101111101100100 +
b101111101100100 1
#446510000000
0#
0(
#446520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#446570000000
0$
0)
#446580000000
1"
1'
b0 +
b0 1
#446630000000
0"
0'
#446640000000
1#
1(
b101111101100100 +
b101111101100100 1
#446690000000
0#
0(
#446700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#446750000000
0$
0)
#446760000000
1"
1'
b0 +
b0 1
#446810000000
0"
0'
#446820000000
1#
1(
b101111101100100 +
b101111101100100 1
#446870000000
0#
0(
#446880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#446930000000
0$
0)
#446940000000
1"
1'
b0 +
b0 1
#446990000000
0"
0'
#447000000000
1#
1(
b101111101100100 +
b101111101100100 1
#447050000000
0#
0(
#447060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#447110000000
0$
0)
#447120000000
1"
1'
b0 +
b0 1
#447170000000
0"
0'
#447180000000
1#
1(
b101111101100100 +
b101111101100100 1
#447230000000
0#
0(
#447240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#447290000000
0$
0)
#447300000000
1"
1'
b0 +
b0 1
#447350000000
0"
0'
#447360000000
1#
1(
b101111101100100 +
b101111101100100 1
#447410000000
0#
0(
#447420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#447470000000
0$
0)
#447480000000
1"
1'
b0 +
b0 1
#447530000000
0"
0'
#447540000000
1#
1(
b101111101100100 +
b101111101100100 1
#447590000000
0#
0(
#447600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#447650000000
0$
0)
#447660000000
1"
1'
b0 +
b0 1
#447710000000
0"
0'
#447720000000
1#
1(
b101111101100100 +
b101111101100100 1
#447770000000
0#
0(
#447780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#447830000000
0$
0)
#447840000000
1"
1'
b0 +
b0 1
#447890000000
0"
0'
#447900000000
1#
1(
b101111101100100 +
b101111101100100 1
#447950000000
0#
0(
#447960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#448010000000
0$
0)
#448020000000
1"
1'
b0 +
b0 1
#448070000000
0"
0'
#448080000000
1#
1(
b101111101100100 +
b101111101100100 1
#448130000000
0#
0(
#448140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#448190000000
0$
0)
#448200000000
1"
1'
b0 +
b0 1
#448250000000
0"
0'
#448260000000
1#
1(
b101111101100100 +
b101111101100100 1
#448310000000
0#
0(
#448320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#448370000000
0$
0)
#448380000000
1"
1'
b0 +
b0 1
#448430000000
0"
0'
#448440000000
1#
1(
b101111101100100 +
b101111101100100 1
#448490000000
0#
0(
#448500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#448550000000
0$
0)
#448560000000
1"
1'
b0 +
b0 1
#448610000000
0"
0'
#448620000000
1#
1(
b101111101100100 +
b101111101100100 1
#448670000000
0#
0(
#448680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#448730000000
0$
0)
#448740000000
1"
1'
b0 +
b0 1
#448790000000
0"
0'
#448800000000
1#
1(
b101111101100100 +
b101111101100100 1
#448850000000
0#
0(
#448860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#448910000000
0$
0)
#448920000000
1"
1'
b0 +
b0 1
#448970000000
0"
0'
#448980000000
1#
1(
b101111101100100 +
b101111101100100 1
#449030000000
0#
0(
#449040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#449090000000
0$
0)
#449100000000
1"
1'
b0 +
b0 1
#449150000000
0"
0'
#449160000000
1#
1(
b101111101100100 +
b101111101100100 1
#449210000000
0#
0(
#449220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#449270000000
0$
0)
#449280000000
1"
1'
b0 +
b0 1
#449330000000
0"
0'
#449340000000
1#
1(
b101111101100100 +
b101111101100100 1
#449390000000
0#
0(
#449400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#449450000000
0$
0)
#449460000000
1"
1'
b0 +
b0 1
#449510000000
0"
0'
#449520000000
1#
1(
b101111101100100 +
b101111101100100 1
#449570000000
0#
0(
#449580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#449630000000
0$
0)
#449640000000
1"
1'
b0 +
b0 1
#449690000000
0"
0'
#449700000000
1#
1(
b101111101100100 +
b101111101100100 1
#449750000000
0#
0(
#449760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#449810000000
0$
0)
#449820000000
1"
1'
b0 +
b0 1
#449870000000
0"
0'
#449880000000
1#
1(
b101111101100100 +
b101111101100100 1
#449930000000
0#
0(
#449940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#449990000000
0$
0)
#450000000000
1"
1'
b0 +
b0 1
#450050000000
0"
0'
#450060000000
1#
1(
b101111101100100 +
b101111101100100 1
#450110000000
0#
0(
#450120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#450170000000
0$
0)
#450180000000
1"
1'
b0 +
b0 1
#450230000000
0"
0'
#450240000000
1#
1(
b101111101100100 +
b101111101100100 1
#450290000000
0#
0(
#450300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#450350000000
0$
0)
#450360000000
1"
1'
b0 +
b0 1
#450410000000
0"
0'
#450420000000
1#
1(
b101111101100100 +
b101111101100100 1
#450470000000
0#
0(
#450480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#450530000000
0$
0)
#450540000000
1"
1'
b0 +
b0 1
#450590000000
0"
0'
#450600000000
1#
1(
b101111101100100 +
b101111101100100 1
#450650000000
0#
0(
#450660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#450710000000
0$
0)
#450720000000
1"
1'
b0 +
b0 1
#450770000000
0"
0'
#450780000000
1#
1(
b101111101100100 +
b101111101100100 1
#450830000000
0#
0(
#450840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#450890000000
0$
0)
#450900000000
1"
1'
b0 +
b0 1
#450950000000
0"
0'
#450960000000
1#
1(
b101111101100100 +
b101111101100100 1
#451010000000
0#
0(
#451020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#451070000000
0$
0)
#451080000000
1"
1'
b0 +
b0 1
#451130000000
0"
0'
#451140000000
1#
1(
b101111101100100 +
b101111101100100 1
#451190000000
0#
0(
#451200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#451250000000
0$
0)
#451260000000
1"
1'
b0 +
b0 1
#451310000000
0"
0'
#451320000000
1#
1(
b101111101100100 +
b101111101100100 1
#451370000000
0#
0(
#451380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#451430000000
0$
0)
#451440000000
1"
1'
b0 +
b0 1
#451490000000
0"
0'
#451500000000
1#
1(
b101111101100100 +
b101111101100100 1
#451550000000
0#
0(
#451560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#451610000000
0$
0)
#451620000000
1"
1'
b0 +
b0 1
#451670000000
0"
0'
#451680000000
1#
1(
b101111101100100 +
b101111101100100 1
#451730000000
0#
0(
#451740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#451790000000
0$
0)
#451800000000
1"
1'
b0 +
b0 1
#451850000000
0"
0'
#451860000000
1#
1(
b101111101100100 +
b101111101100100 1
#451910000000
0#
0(
#451920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#451970000000
0$
0)
#451980000000
1"
1'
b0 +
b0 1
#452030000000
0"
0'
#452040000000
1#
1(
b101111101100100 +
b101111101100100 1
#452090000000
0#
0(
#452100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#452150000000
0$
0)
#452160000000
1"
1'
b0 +
b0 1
#452210000000
0"
0'
#452220000000
1#
1(
b101111101100100 +
b101111101100100 1
#452270000000
0#
0(
#452280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#452330000000
0$
0)
#452340000000
1"
1'
b0 +
b0 1
#452390000000
0"
0'
#452400000000
1#
1(
b101111101100100 +
b101111101100100 1
#452450000000
0#
0(
#452460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#452510000000
0$
0)
#452520000000
1"
1'
b0 +
b0 1
#452570000000
0"
0'
#452580000000
1#
1(
b101111101100100 +
b101111101100100 1
#452630000000
0#
0(
#452640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#452690000000
0$
0)
#452700000000
1"
1'
b0 +
b0 1
#452750000000
0"
0'
#452760000000
1#
1(
b101111101100100 +
b101111101100100 1
#452810000000
0#
0(
#452820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#452870000000
0$
0)
#452880000000
1"
1'
b0 +
b0 1
#452930000000
0"
0'
#452940000000
1#
1(
b101111101100100 +
b101111101100100 1
#452990000000
0#
0(
#453000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#453050000000
0$
0)
#453060000000
1"
1'
b0 +
b0 1
#453110000000
0"
0'
#453120000000
1#
1(
b101111101100100 +
b101111101100100 1
#453170000000
0#
0(
#453180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#453230000000
0$
0)
#453240000000
1"
1'
b0 +
b0 1
#453290000000
0"
0'
#453300000000
1#
1(
b101111101100100 +
b101111101100100 1
#453350000000
0#
0(
#453360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#453410000000
0$
0)
#453420000000
1"
1'
b0 +
b0 1
#453470000000
0"
0'
#453480000000
1#
1(
b101111101100100 +
b101111101100100 1
#453530000000
0#
0(
#453540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#453590000000
0$
0)
#453600000000
1"
1'
b0 +
b0 1
#453650000000
0"
0'
#453660000000
1#
1(
b101111101100100 +
b101111101100100 1
#453710000000
0#
0(
#453720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#453770000000
0$
0)
#453780000000
1"
1'
b0 +
b0 1
#453830000000
0"
0'
#453840000000
1#
1(
b101111101100100 +
b101111101100100 1
#453890000000
0#
0(
#453900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#453950000000
0$
0)
#453960000000
1"
1'
b0 +
b0 1
#454010000000
0"
0'
#454020000000
1#
1(
b101111101100100 +
b101111101100100 1
#454070000000
0#
0(
#454080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#454130000000
0$
0)
#454140000000
1"
1'
b0 +
b0 1
#454190000000
0"
0'
#454200000000
1#
1(
b101111101100100 +
b101111101100100 1
#454250000000
0#
0(
#454260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#454310000000
0$
0)
#454320000000
1"
1'
b0 +
b0 1
#454370000000
0"
0'
#454380000000
1#
1(
b101111101100100 +
b101111101100100 1
#454430000000
0#
0(
#454440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#454490000000
0$
0)
#454500000000
1"
1'
b0 +
b0 1
#454550000000
0"
0'
#454560000000
1#
1(
b101111101100100 +
b101111101100100 1
#454610000000
0#
0(
#454620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#454670000000
0$
0)
#454680000000
1"
1'
b0 +
b0 1
#454730000000
0"
0'
#454740000000
1#
1(
b101111101100100 +
b101111101100100 1
#454790000000
0#
0(
#454800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#454850000000
0$
0)
#454860000000
1"
1'
b0 +
b0 1
#454910000000
0"
0'
#454920000000
1#
1(
b101111101100100 +
b101111101100100 1
#454970000000
0#
0(
#454980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#455030000000
0$
0)
#455040000000
1"
1'
b0 +
b0 1
#455090000000
0"
0'
#455100000000
1#
1(
b101111101100100 +
b101111101100100 1
#455150000000
0#
0(
#455160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#455210000000
0$
0)
#455220000000
1"
1'
b0 +
b0 1
#455270000000
0"
0'
#455280000000
1#
1(
b101111101100100 +
b101111101100100 1
#455330000000
0#
0(
#455340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#455390000000
0$
0)
#455400000000
1"
1'
b0 +
b0 1
#455450000000
0"
0'
#455460000000
1#
1(
b101111101100100 +
b101111101100100 1
#455510000000
0#
0(
#455520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#455570000000
0$
0)
#455580000000
1"
1'
b0 +
b0 1
#455630000000
0"
0'
#455640000000
1#
1(
b101111101100100 +
b101111101100100 1
#455690000000
0#
0(
#455700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#455750000000
0$
0)
#455760000000
1"
1'
b0 +
b0 1
#455810000000
0"
0'
#455820000000
1#
1(
b101111101100100 +
b101111101100100 1
#455870000000
0#
0(
#455880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#455930000000
0$
0)
#455940000000
1"
1'
b0 +
b0 1
#455990000000
0"
0'
#456000000000
1#
1(
b101111101100100 +
b101111101100100 1
#456050000000
0#
0(
#456060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#456110000000
0$
0)
#456120000000
1"
1'
b0 +
b0 1
#456170000000
0"
0'
#456180000000
1#
1(
b101111101100100 +
b101111101100100 1
#456230000000
0#
0(
#456240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#456290000000
0$
0)
#456300000000
1"
1'
b0 +
b0 1
#456350000000
0"
0'
#456360000000
1#
1(
b101111101100100 +
b101111101100100 1
#456410000000
0#
0(
#456420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#456470000000
0$
0)
#456480000000
1"
1'
b0 +
b0 1
#456530000000
0"
0'
#456540000000
1#
1(
b101111101100100 +
b101111101100100 1
#456590000000
0#
0(
#456600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#456650000000
0$
0)
#456660000000
1"
1'
b0 +
b0 1
#456710000000
0"
0'
#456720000000
1#
1(
b101111101100100 +
b101111101100100 1
#456770000000
0#
0(
#456780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#456830000000
0$
0)
#456840000000
1"
1'
b0 +
b0 1
#456890000000
0"
0'
#456900000000
1#
1(
b101111101100100 +
b101111101100100 1
#456950000000
0#
0(
#456960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#457010000000
0$
0)
#457020000000
1"
1'
b0 +
b0 1
#457070000000
0"
0'
#457080000000
1#
1(
b101111101100100 +
b101111101100100 1
#457130000000
0#
0(
#457140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#457190000000
0$
0)
#457200000000
1"
1'
b0 +
b0 1
#457250000000
0"
0'
#457260000000
1#
1(
b101111101100100 +
b101111101100100 1
#457310000000
0#
0(
#457320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#457370000000
0$
0)
#457380000000
1"
1'
b0 +
b0 1
#457430000000
0"
0'
#457440000000
1#
1(
b101111101100100 +
b101111101100100 1
#457490000000
0#
0(
#457500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#457550000000
0$
0)
#457560000000
1"
1'
b0 +
b0 1
#457610000000
0"
0'
#457620000000
1#
1(
b101111101100100 +
b101111101100100 1
#457670000000
0#
0(
#457680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#457730000000
0$
0)
#457740000000
1"
1'
b0 +
b0 1
#457790000000
0"
0'
#457800000000
1#
1(
b101111101100100 +
b101111101100100 1
#457850000000
0#
0(
#457860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#457910000000
0$
0)
#457920000000
1"
1'
b0 +
b0 1
#457970000000
0"
0'
#457980000000
1#
1(
b101111101100100 +
b101111101100100 1
#458030000000
0#
0(
#458040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#458090000000
0$
0)
#458100000000
1"
1'
b0 +
b0 1
#458150000000
0"
0'
#458160000000
1#
1(
b101111101100100 +
b101111101100100 1
#458210000000
0#
0(
#458220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#458270000000
0$
0)
#458280000000
1"
1'
b0 +
b0 1
#458330000000
0"
0'
#458340000000
1#
1(
b101111101100100 +
b101111101100100 1
#458390000000
0#
0(
#458400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#458450000000
0$
0)
#458460000000
1"
1'
b0 +
b0 1
#458510000000
0"
0'
#458520000000
1#
1(
b101111101100100 +
b101111101100100 1
#458570000000
0#
0(
#458580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#458630000000
0$
0)
#458640000000
1"
1'
b0 +
b0 1
#458690000000
0"
0'
#458700000000
1#
1(
b101111101100100 +
b101111101100100 1
#458750000000
0#
0(
#458760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#458810000000
0$
0)
#458820000000
1"
1'
b0 +
b0 1
#458870000000
0"
0'
#458880000000
1#
1(
b101111101100100 +
b101111101100100 1
#458930000000
0#
0(
#458940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#458990000000
0$
0)
#459000000000
1"
1'
b0 +
b0 1
#459050000000
0"
0'
#459060000000
1#
1(
b101111101100100 +
b101111101100100 1
#459110000000
0#
0(
#459120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#459170000000
0$
0)
#459180000000
1"
1'
b0 +
b0 1
#459230000000
0"
0'
#459240000000
1#
1(
b101111101100100 +
b101111101100100 1
#459290000000
0#
0(
#459300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#459350000000
0$
0)
#459360000000
1"
1'
b0 +
b0 1
#459410000000
0"
0'
#459420000000
1#
1(
b101111101100100 +
b101111101100100 1
#459470000000
0#
0(
#459480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#459530000000
0$
0)
#459540000000
1"
1'
b0 +
b0 1
#459590000000
0"
0'
#459600000000
1#
1(
b101111101100100 +
b101111101100100 1
#459650000000
0#
0(
#459660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#459710000000
0$
0)
#459720000000
1"
1'
b0 +
b0 1
#459770000000
0"
0'
#459780000000
1#
1(
b101111101100100 +
b101111101100100 1
#459830000000
0#
0(
#459840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#459890000000
0$
0)
#459900000000
1"
1'
b0 +
b0 1
#459950000000
0"
0'
#459960000000
1#
1(
b101111101100100 +
b101111101100100 1
#460010000000
0#
0(
#460020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#460070000000
0$
0)
#460080000000
1"
1'
b0 +
b0 1
#460130000000
0"
0'
#460140000000
1#
1(
b101111101100100 +
b101111101100100 1
#460190000000
0#
0(
#460200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#460250000000
0$
0)
#460260000000
1"
1'
b0 +
b0 1
#460310000000
0"
0'
#460320000000
1#
1(
b101111101100100 +
b101111101100100 1
#460370000000
0#
0(
#460380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#460430000000
0$
0)
#460440000000
1"
1'
b0 +
b0 1
#460490000000
0"
0'
#460500000000
1#
1(
b101111101100100 +
b101111101100100 1
#460550000000
0#
0(
#460560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#460610000000
0$
0)
#460620000000
1"
1'
b0 +
b0 1
#460670000000
0"
0'
#460680000000
1#
1(
b101111101100100 +
b101111101100100 1
#460730000000
0#
0(
#460740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#460790000000
0$
0)
#460800000000
1"
1'
b0 +
b0 1
#460850000000
0"
0'
#460860000000
1#
1(
b101111101100100 +
b101111101100100 1
#460910000000
0#
0(
#460920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#460970000000
0$
0)
#460980000000
1"
1'
b0 +
b0 1
#461030000000
0"
0'
#461040000000
1#
1(
b101111101100100 +
b101111101100100 1
#461090000000
0#
0(
#461100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#461150000000
0$
0)
#461160000000
1"
1'
b0 +
b0 1
#461210000000
0"
0'
#461220000000
1#
1(
b101111101100100 +
b101111101100100 1
#461270000000
0#
0(
#461280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#461330000000
0$
0)
#461340000000
1"
1'
b0 +
b0 1
#461390000000
0"
0'
#461400000000
1#
1(
b101111101100100 +
b101111101100100 1
#461450000000
0#
0(
#461460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#461510000000
0$
0)
#461520000000
1"
1'
b0 +
b0 1
#461570000000
0"
0'
#461580000000
1#
1(
b101111101100100 +
b101111101100100 1
#461630000000
0#
0(
#461640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#461690000000
0$
0)
#461700000000
1"
1'
b0 +
b0 1
#461750000000
0"
0'
#461760000000
1#
1(
b101111101100100 +
b101111101100100 1
#461810000000
0#
0(
#461820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#461870000000
0$
0)
#461880000000
1"
1'
b0 +
b0 1
#461930000000
0"
0'
#461940000000
1#
1(
b101111101100100 +
b101111101100100 1
#461990000000
0#
0(
#462000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#462050000000
0$
0)
#462060000000
1"
1'
b0 +
b0 1
#462110000000
0"
0'
#462120000000
1#
1(
b101111101100100 +
b101111101100100 1
#462170000000
0#
0(
#462180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#462230000000
0$
0)
#462240000000
1"
1'
b0 +
b0 1
#462290000000
0"
0'
#462300000000
1#
1(
b101111101100100 +
b101111101100100 1
#462350000000
0#
0(
#462360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#462410000000
0$
0)
#462420000000
1"
1'
b0 +
b0 1
#462470000000
0"
0'
#462480000000
1#
1(
b101111101100100 +
b101111101100100 1
#462530000000
0#
0(
#462540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#462590000000
0$
0)
#462600000000
1"
1'
b0 +
b0 1
#462650000000
0"
0'
#462660000000
1#
1(
b101111101100100 +
b101111101100100 1
#462710000000
0#
0(
#462720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#462770000000
0$
0)
#462780000000
1"
1'
b0 +
b0 1
#462830000000
0"
0'
#462840000000
1#
1(
b101111101100100 +
b101111101100100 1
#462890000000
0#
0(
#462900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#462950000000
0$
0)
#462960000000
1"
1'
b0 +
b0 1
#463010000000
0"
0'
#463020000000
1#
1(
b101111101100100 +
b101111101100100 1
#463070000000
0#
0(
#463080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#463130000000
0$
0)
#463140000000
1"
1'
b0 +
b0 1
#463190000000
0"
0'
#463200000000
1#
1(
b101111101100100 +
b101111101100100 1
#463250000000
0#
0(
#463260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#463310000000
0$
0)
#463320000000
1"
1'
b0 +
b0 1
#463370000000
0"
0'
#463380000000
1#
1(
b101111101100100 +
b101111101100100 1
#463430000000
0#
0(
#463440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#463490000000
0$
0)
#463500000000
1"
1'
b0 +
b0 1
#463550000000
0"
0'
#463560000000
1#
1(
b101111101100100 +
b101111101100100 1
#463610000000
0#
0(
#463620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#463670000000
0$
0)
#463680000000
1"
1'
b0 +
b0 1
#463730000000
0"
0'
#463740000000
1#
1(
b101111101100100 +
b101111101100100 1
#463790000000
0#
0(
#463800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#463850000000
0$
0)
#463860000000
1"
1'
b0 +
b0 1
#463910000000
0"
0'
#463920000000
1#
1(
b101111101100100 +
b101111101100100 1
#463970000000
0#
0(
#463980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#464030000000
0$
0)
#464040000000
1"
1'
b0 +
b0 1
#464090000000
0"
0'
#464100000000
1#
1(
b101111101100100 +
b101111101100100 1
#464150000000
0#
0(
#464160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#464210000000
0$
0)
#464220000000
1"
1'
b0 +
b0 1
#464270000000
0"
0'
#464280000000
1#
1(
b101111101100100 +
b101111101100100 1
#464330000000
0#
0(
#464340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#464390000000
0$
0)
#464400000000
1"
1'
b0 +
b0 1
#464450000000
0"
0'
#464460000000
1#
1(
b101111101100100 +
b101111101100100 1
#464510000000
0#
0(
#464520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#464570000000
0$
0)
#464580000000
1"
1'
b0 +
b0 1
#464630000000
0"
0'
#464640000000
1#
1(
b101111101100100 +
b101111101100100 1
#464690000000
0#
0(
#464700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#464750000000
0$
0)
#464760000000
1"
1'
b0 +
b0 1
#464810000000
0"
0'
#464820000000
1#
1(
b101111101100100 +
b101111101100100 1
#464870000000
0#
0(
#464880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#464930000000
0$
0)
#464940000000
1"
1'
b0 +
b0 1
#464990000000
0"
0'
#465000000000
1#
1(
b101111101100100 +
b101111101100100 1
#465050000000
0#
0(
#465060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#465110000000
0$
0)
#465120000000
1"
1'
b0 +
b0 1
#465170000000
0"
0'
#465180000000
1#
1(
b101111101100100 +
b101111101100100 1
#465230000000
0#
0(
#465240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#465290000000
0$
0)
#465300000000
1"
1'
b0 +
b0 1
#465350000000
0"
0'
#465360000000
1#
1(
b101111101100100 +
b101111101100100 1
#465410000000
0#
0(
#465420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#465470000000
0$
0)
#465480000000
1"
1'
b0 +
b0 1
#465530000000
0"
0'
#465540000000
1#
1(
b101111101100100 +
b101111101100100 1
#465590000000
0#
0(
#465600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#465650000000
0$
0)
#465660000000
1"
1'
b0 +
b0 1
#465710000000
0"
0'
#465720000000
1#
1(
b101111101100100 +
b101111101100100 1
#465770000000
0#
0(
#465780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#465830000000
0$
0)
#465840000000
1"
1'
b0 +
b0 1
#465890000000
0"
0'
#465900000000
1#
1(
b101111101100100 +
b101111101100100 1
#465950000000
0#
0(
#465960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#466010000000
0$
0)
#466020000000
1"
1'
b0 +
b0 1
#466070000000
0"
0'
#466080000000
1#
1(
b101111101100100 +
b101111101100100 1
#466130000000
0#
0(
#466140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#466190000000
0$
0)
#466200000000
1"
1'
b0 +
b0 1
#466250000000
0"
0'
#466260000000
1#
1(
b101111101100100 +
b101111101100100 1
#466310000000
0#
0(
#466320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#466370000000
0$
0)
#466380000000
1"
1'
b0 +
b0 1
#466430000000
0"
0'
#466440000000
1#
1(
b101111101100100 +
b101111101100100 1
#466490000000
0#
0(
#466500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#466550000000
0$
0)
#466560000000
1"
1'
b0 +
b0 1
#466610000000
0"
0'
#466620000000
1#
1(
b101111101100100 +
b101111101100100 1
#466670000000
0#
0(
#466680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#466730000000
0$
0)
#466740000000
1"
1'
b0 +
b0 1
#466790000000
0"
0'
#466800000000
1#
1(
b101111101100100 +
b101111101100100 1
#466850000000
0#
0(
#466860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#466910000000
0$
0)
#466920000000
1"
1'
b0 +
b0 1
#466970000000
0"
0'
#466980000000
1#
1(
b101111101100100 +
b101111101100100 1
#467030000000
0#
0(
#467040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#467090000000
0$
0)
#467100000000
1"
1'
b0 +
b0 1
#467150000000
0"
0'
#467160000000
1#
1(
b101111101100100 +
b101111101100100 1
#467210000000
0#
0(
#467220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#467270000000
0$
0)
#467280000000
1"
1'
b0 +
b0 1
#467330000000
0"
0'
#467340000000
1#
1(
b101111101100100 +
b101111101100100 1
#467390000000
0#
0(
#467400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#467450000000
0$
0)
#467460000000
1"
1'
b0 +
b0 1
#467510000000
0"
0'
#467520000000
1#
1(
b101111101100100 +
b101111101100100 1
#467570000000
0#
0(
#467580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#467630000000
0$
0)
#467640000000
1"
1'
b0 +
b0 1
#467690000000
0"
0'
#467700000000
1#
1(
b101111101100100 +
b101111101100100 1
#467750000000
0#
0(
#467760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#467810000000
0$
0)
#467820000000
1"
1'
b0 +
b0 1
#467870000000
0"
0'
#467880000000
1#
1(
b101111101100100 +
b101111101100100 1
#467930000000
0#
0(
#467940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#467990000000
0$
0)
#468000000000
1"
1'
b0 +
b0 1
#468050000000
0"
0'
#468060000000
1#
1(
b101111101100100 +
b101111101100100 1
#468110000000
0#
0(
#468120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#468170000000
0$
0)
#468180000000
1"
1'
b0 +
b0 1
#468230000000
0"
0'
#468240000000
1#
1(
b101111101100100 +
b101111101100100 1
#468290000000
0#
0(
#468300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#468350000000
0$
0)
#468360000000
1"
1'
b0 +
b0 1
#468410000000
0"
0'
#468420000000
1#
1(
b101111101100100 +
b101111101100100 1
#468470000000
0#
0(
#468480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#468530000000
0$
0)
#468540000000
1"
1'
b0 +
b0 1
#468590000000
0"
0'
#468600000000
1#
1(
b101111101100100 +
b101111101100100 1
#468650000000
0#
0(
#468660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#468710000000
0$
0)
#468720000000
1"
1'
b0 +
b0 1
#468770000000
0"
0'
#468780000000
1#
1(
b101111101100100 +
b101111101100100 1
#468830000000
0#
0(
#468840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#468890000000
0$
0)
#468900000000
1"
1'
b0 +
b0 1
#468950000000
0"
0'
#468960000000
1#
1(
b101111101100100 +
b101111101100100 1
#469010000000
0#
0(
#469020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#469070000000
0$
0)
#469080000000
1"
1'
b0 +
b0 1
#469130000000
0"
0'
#469140000000
1#
1(
b101111101100100 +
b101111101100100 1
#469190000000
0#
0(
#469200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#469250000000
0$
0)
#469260000000
1"
1'
b0 +
b0 1
#469310000000
0"
0'
#469320000000
1#
1(
b101111101100100 +
b101111101100100 1
#469370000000
0#
0(
#469380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#469430000000
0$
0)
#469440000000
1"
1'
b0 +
b0 1
#469490000000
0"
0'
#469500000000
1#
1(
b101111101100100 +
b101111101100100 1
#469550000000
0#
0(
#469560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#469610000000
0$
0)
#469620000000
1"
1'
b0 +
b0 1
#469670000000
0"
0'
#469680000000
1#
1(
b101111101100100 +
b101111101100100 1
#469730000000
0#
0(
#469740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#469790000000
0$
0)
#469800000000
1"
1'
b0 +
b0 1
#469850000000
0"
0'
#469860000000
1#
1(
b101111101100100 +
b101111101100100 1
#469910000000
0#
0(
#469920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#469970000000
0$
0)
#469980000000
1"
1'
b0 +
b0 1
#470030000000
0"
0'
#470040000000
1#
1(
b101111101100100 +
b101111101100100 1
#470090000000
0#
0(
#470100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#470150000000
0$
0)
#470160000000
1"
1'
b0 +
b0 1
#470210000000
0"
0'
#470220000000
1#
1(
b101111101100100 +
b101111101100100 1
#470270000000
0#
0(
#470280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#470330000000
0$
0)
#470340000000
1"
1'
b0 +
b0 1
#470390000000
0"
0'
#470400000000
1#
1(
b101111101100100 +
b101111101100100 1
#470450000000
0#
0(
#470460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#470510000000
0$
0)
#470520000000
1"
1'
b0 +
b0 1
#470570000000
0"
0'
#470580000000
1#
1(
b101111101100100 +
b101111101100100 1
#470630000000
0#
0(
#470640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#470690000000
0$
0)
#470700000000
1"
1'
b0 +
b0 1
#470750000000
0"
0'
#470760000000
1#
1(
b101111101100100 +
b101111101100100 1
#470810000000
0#
0(
#470820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#470870000000
0$
0)
#470880000000
1"
1'
b0 +
b0 1
#470930000000
0"
0'
#470940000000
1#
1(
b101111101100100 +
b101111101100100 1
#470990000000
0#
0(
#471000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#471050000000
0$
0)
#471060000000
1"
1'
b0 +
b0 1
#471110000000
0"
0'
#471120000000
1#
1(
b101111101100100 +
b101111101100100 1
#471170000000
0#
0(
#471180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#471230000000
0$
0)
#471240000000
1"
1'
b0 +
b0 1
#471290000000
0"
0'
#471300000000
1#
1(
b101111101100100 +
b101111101100100 1
#471350000000
0#
0(
#471360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#471410000000
0$
0)
#471420000000
1"
1'
b0 +
b0 1
#471470000000
0"
0'
#471480000000
1#
1(
b101111101100100 +
b101111101100100 1
#471530000000
0#
0(
#471540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#471590000000
0$
0)
#471600000000
1"
1'
b0 +
b0 1
#471650000000
0"
0'
#471660000000
1#
1(
b101111101100100 +
b101111101100100 1
#471710000000
0#
0(
#471720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#471770000000
0$
0)
#471780000000
1"
1'
b0 +
b0 1
#471830000000
0"
0'
#471840000000
1#
1(
b101111101100100 +
b101111101100100 1
#471890000000
0#
0(
#471900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#471950000000
0$
0)
#471960000000
1"
1'
b0 +
b0 1
#472010000000
0"
0'
#472020000000
1#
1(
b101111101100100 +
b101111101100100 1
#472070000000
0#
0(
#472080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#472130000000
0$
0)
#472140000000
1"
1'
b0 +
b0 1
#472190000000
0"
0'
#472200000000
1#
1(
b101111101100100 +
b101111101100100 1
#472250000000
0#
0(
#472260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#472310000000
0$
0)
#472320000000
1"
1'
b0 +
b0 1
#472370000000
0"
0'
#472380000000
1#
1(
b101111101100100 +
b101111101100100 1
#472430000000
0#
0(
#472440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#472490000000
0$
0)
#472500000000
1"
1'
b0 +
b0 1
#472550000000
0"
0'
#472560000000
1#
1(
b101111101100100 +
b101111101100100 1
#472610000000
0#
0(
#472620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#472670000000
0$
0)
#472680000000
1"
1'
b0 +
b0 1
#472730000000
0"
0'
#472740000000
1#
1(
b101111101100100 +
b101111101100100 1
#472790000000
0#
0(
#472800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#472850000000
0$
0)
#472860000000
1"
1'
b0 +
b0 1
#472910000000
0"
0'
#472920000000
1#
1(
b101111101100100 +
b101111101100100 1
#472970000000
0#
0(
#472980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#473030000000
0$
0)
#473040000000
1"
1'
b0 +
b0 1
#473090000000
0"
0'
#473100000000
1#
1(
b101111101100100 +
b101111101100100 1
#473150000000
0#
0(
#473160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#473210000000
0$
0)
#473220000000
1"
1'
b0 +
b0 1
#473270000000
0"
0'
#473280000000
1#
1(
b101111101100100 +
b101111101100100 1
#473330000000
0#
0(
#473340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#473390000000
0$
0)
#473400000000
1"
1'
b0 +
b0 1
#473450000000
0"
0'
#473460000000
1#
1(
b101111101100100 +
b101111101100100 1
#473510000000
0#
0(
#473520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#473570000000
0$
0)
#473580000000
1"
1'
b0 +
b0 1
#473630000000
0"
0'
#473640000000
1#
1(
b101111101100100 +
b101111101100100 1
#473690000000
0#
0(
#473700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#473750000000
0$
0)
#473760000000
1"
1'
b0 +
b0 1
#473810000000
0"
0'
#473820000000
1#
1(
b101111101100100 +
b101111101100100 1
#473870000000
0#
0(
#473880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#473930000000
0$
0)
#473940000000
1"
1'
b0 +
b0 1
#473990000000
0"
0'
#474000000000
1#
1(
b101111101100100 +
b101111101100100 1
#474050000000
0#
0(
#474060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#474110000000
0$
0)
#474120000000
1"
1'
b0 +
b0 1
#474170000000
0"
0'
#474180000000
1#
1(
b101111101100100 +
b101111101100100 1
#474230000000
0#
0(
#474240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#474290000000
0$
0)
#474300000000
1"
1'
b0 +
b0 1
#474350000000
0"
0'
#474360000000
1#
1(
b101111101100100 +
b101111101100100 1
#474410000000
0#
0(
#474420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#474470000000
0$
0)
#474480000000
1"
1'
b0 +
b0 1
#474530000000
0"
0'
#474540000000
1#
1(
b101111101100100 +
b101111101100100 1
#474590000000
0#
0(
#474600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#474650000000
0$
0)
#474660000000
1"
1'
b0 +
b0 1
#474710000000
0"
0'
#474720000000
1#
1(
b101111101100100 +
b101111101100100 1
#474770000000
0#
0(
#474780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#474830000000
0$
0)
#474840000000
1"
1'
b0 +
b0 1
#474890000000
0"
0'
#474900000000
1#
1(
b101111101100100 +
b101111101100100 1
#474950000000
0#
0(
#474960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#475010000000
0$
0)
#475020000000
1"
1'
b0 +
b0 1
#475070000000
0"
0'
#475080000000
1#
1(
b101111101100100 +
b101111101100100 1
#475130000000
0#
0(
#475140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#475190000000
0$
0)
#475200000000
1"
1'
b0 +
b0 1
#475250000000
0"
0'
#475260000000
1#
1(
b101111101100100 +
b101111101100100 1
#475310000000
0#
0(
#475320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#475370000000
0$
0)
#475380000000
1"
1'
b0 +
b0 1
#475430000000
0"
0'
#475440000000
1#
1(
b101111101100100 +
b101111101100100 1
#475490000000
0#
0(
#475500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#475550000000
0$
0)
#475560000000
1"
1'
b0 +
b0 1
#475610000000
0"
0'
#475620000000
1#
1(
b101111101100100 +
b101111101100100 1
#475670000000
0#
0(
#475680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#475730000000
0$
0)
#475740000000
1"
1'
b0 +
b0 1
#475790000000
0"
0'
#475800000000
1#
1(
b101111101100100 +
b101111101100100 1
#475850000000
0#
0(
#475860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#475910000000
0$
0)
#475920000000
1"
1'
b0 +
b0 1
#475970000000
0"
0'
#475980000000
1#
1(
b101111101100100 +
b101111101100100 1
#476030000000
0#
0(
#476040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#476090000000
0$
0)
#476100000000
1"
1'
b0 +
b0 1
#476150000000
0"
0'
#476160000000
1#
1(
b101111101100100 +
b101111101100100 1
#476210000000
0#
0(
#476220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#476270000000
0$
0)
#476280000000
1"
1'
b0 +
b0 1
#476330000000
0"
0'
#476340000000
1#
1(
b101111101100100 +
b101111101100100 1
#476390000000
0#
0(
#476400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#476450000000
0$
0)
#476460000000
1"
1'
b0 +
b0 1
#476510000000
0"
0'
#476520000000
1#
1(
b101111101100100 +
b101111101100100 1
#476570000000
0#
0(
#476580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#476630000000
0$
0)
#476640000000
1"
1'
b0 +
b0 1
#476690000000
0"
0'
#476700000000
1#
1(
b101111101100100 +
b101111101100100 1
#476750000000
0#
0(
#476760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#476810000000
0$
0)
#476820000000
1"
1'
b0 +
b0 1
#476870000000
0"
0'
#476880000000
1#
1(
b101111101100100 +
b101111101100100 1
#476930000000
0#
0(
#476940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#476990000000
0$
0)
#477000000000
1"
1'
b0 +
b0 1
#477050000000
0"
0'
#477060000000
1#
1(
b101111101100100 +
b101111101100100 1
#477110000000
0#
0(
#477120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#477170000000
0$
0)
#477180000000
1"
1'
b0 +
b0 1
#477230000000
0"
0'
#477240000000
1#
1(
b101111101100100 +
b101111101100100 1
#477290000000
0#
0(
#477300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#477350000000
0$
0)
#477360000000
1"
1'
b0 +
b0 1
#477410000000
0"
0'
#477420000000
1#
1(
b101111101100100 +
b101111101100100 1
#477470000000
0#
0(
#477480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#477530000000
0$
0)
#477540000000
1"
1'
b0 +
b0 1
#477590000000
0"
0'
#477600000000
1#
1(
b101111101100100 +
b101111101100100 1
#477650000000
0#
0(
#477660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#477710000000
0$
0)
#477720000000
1"
1'
b0 +
b0 1
#477770000000
0"
0'
#477780000000
1#
1(
b101111101100100 +
b101111101100100 1
#477830000000
0#
0(
#477840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#477890000000
0$
0)
#477900000000
1"
1'
b0 +
b0 1
#477950000000
0"
0'
#477960000000
1#
1(
b101111101100100 +
b101111101100100 1
#478010000000
0#
0(
#478020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#478070000000
0$
0)
#478080000000
1"
1'
b0 +
b0 1
#478130000000
0"
0'
#478140000000
1#
1(
b101111101100100 +
b101111101100100 1
#478190000000
0#
0(
#478200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#478250000000
0$
0)
#478260000000
1"
1'
b0 +
b0 1
#478310000000
0"
0'
#478320000000
1#
1(
b101111101100100 +
b101111101100100 1
#478370000000
0#
0(
#478380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#478430000000
0$
0)
#478440000000
1"
1'
b0 +
b0 1
#478490000000
0"
0'
#478500000000
1#
1(
b101111101100100 +
b101111101100100 1
#478550000000
0#
0(
#478560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#478610000000
0$
0)
#478620000000
1"
1'
b0 +
b0 1
#478670000000
0"
0'
#478680000000
1#
1(
b101111101100100 +
b101111101100100 1
#478730000000
0#
0(
#478740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#478790000000
0$
0)
#478800000000
1"
1'
b0 +
b0 1
#478850000000
0"
0'
#478860000000
1#
1(
b101111101100100 +
b101111101100100 1
#478910000000
0#
0(
#478920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#478970000000
0$
0)
#478980000000
1"
1'
b0 +
b0 1
#479030000000
0"
0'
#479040000000
1#
1(
b101111101100100 +
b101111101100100 1
#479090000000
0#
0(
#479100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#479150000000
0$
0)
#479160000000
1"
1'
b0 +
b0 1
#479210000000
0"
0'
#479220000000
1#
1(
b101111101100100 +
b101111101100100 1
#479270000000
0#
0(
#479280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#479330000000
0$
0)
#479340000000
1"
1'
b0 +
b0 1
#479390000000
0"
0'
#479400000000
1#
1(
b101111101100100 +
b101111101100100 1
#479450000000
0#
0(
#479460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#479510000000
0$
0)
#479520000000
1"
1'
b0 +
b0 1
#479570000000
0"
0'
#479580000000
1#
1(
b101111101100100 +
b101111101100100 1
#479630000000
0#
0(
#479640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#479690000000
0$
0)
#479700000000
1"
1'
b0 +
b0 1
#479750000000
0"
0'
#479760000000
1#
1(
b101111101100100 +
b101111101100100 1
#479810000000
0#
0(
#479820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#479870000000
0$
0)
#479880000000
1"
1'
b0 +
b0 1
#479930000000
0"
0'
#479940000000
1#
1(
b101111101100100 +
b101111101100100 1
#479990000000
0#
0(
#480000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#480050000000
0$
0)
#480060000000
1"
1'
b0 +
b0 1
#480110000000
0"
0'
#480120000000
1#
1(
b101111101100100 +
b101111101100100 1
#480170000000
0#
0(
#480180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#480230000000
0$
0)
#480240000000
1"
1'
b0 +
b0 1
#480290000000
0"
0'
#480300000000
1#
1(
b101111101100100 +
b101111101100100 1
#480350000000
0#
0(
#480360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#480410000000
0$
0)
#480420000000
1"
1'
b0 +
b0 1
#480470000000
0"
0'
#480480000000
1#
1(
b101111101100100 +
b101111101100100 1
#480530000000
0#
0(
#480540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#480590000000
0$
0)
#480600000000
1"
1'
b0 +
b0 1
#480650000000
0"
0'
#480660000000
1#
1(
b101111101100100 +
b101111101100100 1
#480710000000
0#
0(
#480720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#480770000000
0$
0)
#480780000000
1"
1'
b0 +
b0 1
#480830000000
0"
0'
#480840000000
1#
1(
b101111101100100 +
b101111101100100 1
#480890000000
0#
0(
#480900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#480950000000
0$
0)
#480960000000
1"
1'
b0 +
b0 1
#481010000000
0"
0'
#481020000000
1#
1(
b101111101100100 +
b101111101100100 1
#481070000000
0#
0(
#481080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#481130000000
0$
0)
#481140000000
1"
1'
b0 +
b0 1
#481190000000
0"
0'
#481200000000
1#
1(
b101111101100100 +
b101111101100100 1
#481250000000
0#
0(
#481260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#481310000000
0$
0)
#481320000000
1"
1'
b0 +
b0 1
#481370000000
0"
0'
#481380000000
1#
1(
b101111101100100 +
b101111101100100 1
#481430000000
0#
0(
#481440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#481490000000
0$
0)
#481500000000
1"
1'
b0 +
b0 1
#481550000000
0"
0'
#481560000000
1#
1(
b101111101100100 +
b101111101100100 1
#481610000000
0#
0(
#481620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#481670000000
0$
0)
#481680000000
1"
1'
b0 +
b0 1
#481730000000
0"
0'
#481740000000
1#
1(
b101111101100100 +
b101111101100100 1
#481790000000
0#
0(
#481800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#481850000000
0$
0)
#481860000000
1"
1'
b0 +
b0 1
#481910000000
0"
0'
#481920000000
1#
1(
b101111101100100 +
b101111101100100 1
#481970000000
0#
0(
#481980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#482030000000
0$
0)
#482040000000
1"
1'
b0 +
b0 1
#482090000000
0"
0'
#482100000000
1#
1(
b101111101100100 +
b101111101100100 1
#482150000000
0#
0(
#482160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#482210000000
0$
0)
#482220000000
1"
1'
b0 +
b0 1
#482270000000
0"
0'
#482280000000
1#
1(
b101111101100100 +
b101111101100100 1
#482330000000
0#
0(
#482340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#482390000000
0$
0)
#482400000000
1"
1'
b0 +
b0 1
#482450000000
0"
0'
#482460000000
1#
1(
b101111101100100 +
b101111101100100 1
#482510000000
0#
0(
#482520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#482570000000
0$
0)
#482580000000
1"
1'
b0 +
b0 1
#482630000000
0"
0'
#482640000000
1#
1(
b101111101100100 +
b101111101100100 1
#482690000000
0#
0(
#482700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#482750000000
0$
0)
#482760000000
1"
1'
b0 +
b0 1
#482810000000
0"
0'
#482820000000
1#
1(
b101111101100100 +
b101111101100100 1
#482870000000
0#
0(
#482880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#482930000000
0$
0)
#482940000000
1"
1'
b0 +
b0 1
#482990000000
0"
0'
#483000000000
1#
1(
b101111101100100 +
b101111101100100 1
#483050000000
0#
0(
#483060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#483110000000
0$
0)
#483120000000
1"
1'
b0 +
b0 1
#483170000000
0"
0'
#483180000000
1#
1(
b101111101100100 +
b101111101100100 1
#483230000000
0#
0(
#483240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#483290000000
0$
0)
#483300000000
1"
1'
b0 +
b0 1
#483350000000
0"
0'
#483360000000
1#
1(
b101111101100100 +
b101111101100100 1
#483410000000
0#
0(
#483420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#483470000000
0$
0)
#483480000000
1"
1'
b0 +
b0 1
#483530000000
0"
0'
#483540000000
1#
1(
b101111101100100 +
b101111101100100 1
#483590000000
0#
0(
#483600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#483650000000
0$
0)
#483660000000
1"
1'
b0 +
b0 1
#483710000000
0"
0'
#483720000000
1#
1(
b101111101100100 +
b101111101100100 1
#483770000000
0#
0(
#483780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#483830000000
0$
0)
#483840000000
1"
1'
b0 +
b0 1
#483890000000
0"
0'
#483900000000
1#
1(
b101111101100100 +
b101111101100100 1
#483950000000
0#
0(
#483960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#484010000000
0$
0)
#484020000000
1"
1'
b0 +
b0 1
#484070000000
0"
0'
#484080000000
1#
1(
b101111101100100 +
b101111101100100 1
#484130000000
0#
0(
#484140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#484190000000
0$
0)
#484200000000
1"
1'
b0 +
b0 1
#484250000000
0"
0'
#484260000000
1#
1(
b101111101100100 +
b101111101100100 1
#484310000000
0#
0(
#484320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#484370000000
0$
0)
#484380000000
1"
1'
b0 +
b0 1
#484430000000
0"
0'
#484440000000
1#
1(
b101111101100100 +
b101111101100100 1
#484490000000
0#
0(
#484500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#484550000000
0$
0)
#484560000000
1"
1'
b0 +
b0 1
#484610000000
0"
0'
#484620000000
1#
1(
b101111101100100 +
b101111101100100 1
#484670000000
0#
0(
#484680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#484730000000
0$
0)
#484740000000
1"
1'
b0 +
b0 1
#484790000000
0"
0'
#484800000000
1#
1(
b101111101100100 +
b101111101100100 1
#484850000000
0#
0(
#484860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#484910000000
0$
0)
#484920000000
1"
1'
b0 +
b0 1
#484970000000
0"
0'
#484980000000
1#
1(
b101111101100100 +
b101111101100100 1
#485030000000
0#
0(
#485040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#485090000000
0$
0)
#485100000000
1"
1'
b0 +
b0 1
#485150000000
0"
0'
#485160000000
1#
1(
b101111101100100 +
b101111101100100 1
#485210000000
0#
0(
#485220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#485270000000
0$
0)
#485280000000
1"
1'
b0 +
b0 1
#485330000000
0"
0'
#485340000000
1#
1(
b101111101100100 +
b101111101100100 1
#485390000000
0#
0(
#485400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#485450000000
0$
0)
#485460000000
1"
1'
b0 +
b0 1
#485510000000
0"
0'
#485520000000
1#
1(
b101111101100100 +
b101111101100100 1
#485570000000
0#
0(
#485580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#485630000000
0$
0)
#485640000000
1"
1'
b0 +
b0 1
#485690000000
0"
0'
#485700000000
1#
1(
b101111101100100 +
b101111101100100 1
#485750000000
0#
0(
#485760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#485810000000
0$
0)
#485820000000
1"
1'
b0 +
b0 1
#485870000000
0"
0'
#485880000000
1#
1(
b101111101100100 +
b101111101100100 1
#485930000000
0#
0(
#485940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#485990000000
0$
0)
#486000000000
1"
1'
b0 +
b0 1
#486050000000
0"
0'
#486060000000
1#
1(
b101111101100100 +
b101111101100100 1
#486110000000
0#
0(
#486120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#486170000000
0$
0)
#486180000000
1"
1'
b0 +
b0 1
#486230000000
0"
0'
#486240000000
1#
1(
b101111101100100 +
b101111101100100 1
#486290000000
0#
0(
#486300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#486350000000
0$
0)
#486360000000
1"
1'
b0 +
b0 1
#486410000000
0"
0'
#486420000000
1#
1(
b101111101100100 +
b101111101100100 1
#486470000000
0#
0(
#486480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#486530000000
0$
0)
#486540000000
1"
1'
b0 +
b0 1
#486590000000
0"
0'
#486600000000
1#
1(
b101111101100100 +
b101111101100100 1
#486650000000
0#
0(
#486660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#486710000000
0$
0)
#486720000000
1"
1'
b0 +
b0 1
#486770000000
0"
0'
#486780000000
1#
1(
b101111101100100 +
b101111101100100 1
#486830000000
0#
0(
#486840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#486890000000
0$
0)
#486900000000
1"
1'
b0 +
b0 1
#486950000000
0"
0'
#486960000000
1#
1(
b101111101100100 +
b101111101100100 1
#487010000000
0#
0(
#487020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#487070000000
0$
0)
#487080000000
1"
1'
b0 +
b0 1
#487130000000
0"
0'
#487140000000
1#
1(
b101111101100100 +
b101111101100100 1
#487190000000
0#
0(
#487200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#487250000000
0$
0)
#487260000000
1"
1'
b0 +
b0 1
#487310000000
0"
0'
#487320000000
1#
1(
b101111101100100 +
b101111101100100 1
#487370000000
0#
0(
#487380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#487430000000
0$
0)
#487440000000
1"
1'
b0 +
b0 1
#487490000000
0"
0'
#487500000000
1#
1(
b101111101100100 +
b101111101100100 1
#487550000000
0#
0(
#487560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#487610000000
0$
0)
#487620000000
1"
1'
b0 +
b0 1
#487670000000
0"
0'
#487680000000
1#
1(
b101111101100100 +
b101111101100100 1
#487730000000
0#
0(
#487740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#487790000000
0$
0)
#487800000000
1"
1'
b0 +
b0 1
#487850000000
0"
0'
#487860000000
1#
1(
b101111101100100 +
b101111101100100 1
#487910000000
0#
0(
#487920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#487970000000
0$
0)
#487980000000
1"
1'
b0 +
b0 1
#488030000000
0"
0'
#488040000000
1#
1(
b101111101100100 +
b101111101100100 1
#488090000000
0#
0(
#488100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#488150000000
0$
0)
#488160000000
1"
1'
b0 +
b0 1
#488210000000
0"
0'
#488220000000
1#
1(
b101111101100100 +
b101111101100100 1
#488270000000
0#
0(
#488280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#488330000000
0$
0)
#488340000000
1"
1'
b0 +
b0 1
#488390000000
0"
0'
#488400000000
1#
1(
b101111101100100 +
b101111101100100 1
#488450000000
0#
0(
#488460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#488510000000
0$
0)
#488520000000
1"
1'
b0 +
b0 1
#488570000000
0"
0'
#488580000000
1#
1(
b101111101100100 +
b101111101100100 1
#488630000000
0#
0(
#488640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#488690000000
0$
0)
#488700000000
1"
1'
b0 +
b0 1
#488750000000
0"
0'
#488760000000
1#
1(
b101111101100100 +
b101111101100100 1
#488810000000
0#
0(
#488820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#488870000000
0$
0)
#488880000000
1"
1'
b0 +
b0 1
#488930000000
0"
0'
#488940000000
1#
1(
b101111101100100 +
b101111101100100 1
#488990000000
0#
0(
#489000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#489050000000
0$
0)
#489060000000
1"
1'
b0 +
b0 1
#489110000000
0"
0'
#489120000000
1#
1(
b101111101100100 +
b101111101100100 1
#489170000000
0#
0(
#489180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#489230000000
0$
0)
#489240000000
1"
1'
b0 +
b0 1
#489290000000
0"
0'
#489300000000
1#
1(
b101111101100100 +
b101111101100100 1
#489350000000
0#
0(
#489360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#489410000000
0$
0)
#489420000000
1"
1'
b0 +
b0 1
#489470000000
0"
0'
#489480000000
1#
1(
b101111101100100 +
b101111101100100 1
#489530000000
0#
0(
#489540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#489590000000
0$
0)
#489600000000
1"
1'
b0 +
b0 1
#489650000000
0"
0'
#489660000000
1#
1(
b101111101100100 +
b101111101100100 1
#489710000000
0#
0(
#489720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#489770000000
0$
0)
#489780000000
1"
1'
b0 +
b0 1
#489830000000
0"
0'
#489840000000
1#
1(
b101111101100100 +
b101111101100100 1
#489890000000
0#
0(
#489900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#489950000000
0$
0)
#489960000000
1"
1'
b0 +
b0 1
#490010000000
0"
0'
#490020000000
1#
1(
b101111101100100 +
b101111101100100 1
#490070000000
0#
0(
#490080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#490130000000
0$
0)
#490140000000
1"
1'
b0 +
b0 1
#490190000000
0"
0'
#490200000000
1#
1(
b101111101100100 +
b101111101100100 1
#490250000000
0#
0(
#490260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#490310000000
0$
0)
#490320000000
1"
1'
b0 +
b0 1
#490370000000
0"
0'
#490380000000
1#
1(
b101111101100100 +
b101111101100100 1
#490430000000
0#
0(
#490440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#490490000000
0$
0)
#490500000000
1"
1'
b0 +
b0 1
#490550000000
0"
0'
#490560000000
1#
1(
b101111101100100 +
b101111101100100 1
#490610000000
0#
0(
#490620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#490670000000
0$
0)
#490680000000
1"
1'
b0 +
b0 1
#490730000000
0"
0'
#490740000000
1#
1(
b101111101100100 +
b101111101100100 1
#490790000000
0#
0(
#490800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#490850000000
0$
0)
#490860000000
1"
1'
b0 +
b0 1
#490910000000
0"
0'
#490920000000
1#
1(
b101111101100100 +
b101111101100100 1
#490970000000
0#
0(
#490980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#491030000000
0$
0)
#491040000000
1"
1'
b0 +
b0 1
#491090000000
0"
0'
#491100000000
1#
1(
b101111101100100 +
b101111101100100 1
#491150000000
0#
0(
#491160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#491210000000
0$
0)
#491220000000
1"
1'
b0 +
b0 1
#491270000000
0"
0'
#491280000000
1#
1(
b101111101100100 +
b101111101100100 1
#491330000000
0#
0(
#491340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#491390000000
0$
0)
#491400000000
1"
1'
b0 +
b0 1
#491450000000
0"
0'
#491460000000
1#
1(
b101111101100100 +
b101111101100100 1
#491510000000
0#
0(
#491520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#491570000000
0$
0)
#491580000000
1"
1'
b0 +
b0 1
#491630000000
0"
0'
#491640000000
1#
1(
b101111101100100 +
b101111101100100 1
#491690000000
0#
0(
#491700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#491750000000
0$
0)
#491760000000
1"
1'
b0 +
b0 1
#491810000000
0"
0'
#491820000000
1#
1(
b101111101100100 +
b101111101100100 1
#491870000000
0#
0(
#491880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#491930000000
0$
0)
#491940000000
1"
1'
b0 +
b0 1
#491990000000
0"
0'
#492000000000
1#
1(
b101111101100100 +
b101111101100100 1
#492050000000
0#
0(
#492060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#492110000000
0$
0)
#492120000000
1"
1'
b0 +
b0 1
#492170000000
0"
0'
#492180000000
1#
1(
b101111101100100 +
b101111101100100 1
#492230000000
0#
0(
#492240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#492290000000
0$
0)
#492300000000
1"
1'
b0 +
b0 1
#492350000000
0"
0'
#492360000000
1#
1(
b101111101100100 +
b101111101100100 1
#492410000000
0#
0(
#492420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#492470000000
0$
0)
#492480000000
1"
1'
b0 +
b0 1
#492530000000
0"
0'
#492540000000
1#
1(
b101111101100100 +
b101111101100100 1
#492590000000
0#
0(
#492600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#492650000000
0$
0)
#492660000000
1"
1'
b0 +
b0 1
#492710000000
0"
0'
#492720000000
1#
1(
b101111101100100 +
b101111101100100 1
#492770000000
0#
0(
#492780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#492830000000
0$
0)
#492840000000
1"
1'
b0 +
b0 1
#492890000000
0"
0'
#492900000000
1#
1(
b101111101100100 +
b101111101100100 1
#492950000000
0#
0(
#492960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#493010000000
0$
0)
#493020000000
1"
1'
b0 +
b0 1
#493070000000
0"
0'
#493080000000
1#
1(
b101111101100100 +
b101111101100100 1
#493130000000
0#
0(
#493140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#493190000000
0$
0)
#493200000000
1"
1'
b0 +
b0 1
#493250000000
0"
0'
#493260000000
1#
1(
b101111101100100 +
b101111101100100 1
#493310000000
0#
0(
#493320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#493370000000
0$
0)
#493380000000
1"
1'
b0 +
b0 1
#493430000000
0"
0'
#493440000000
1#
1(
b101111101100100 +
b101111101100100 1
#493490000000
0#
0(
#493500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#493550000000
0$
0)
#493560000000
1"
1'
b0 +
b0 1
#493610000000
0"
0'
#493620000000
1#
1(
b101111101100100 +
b101111101100100 1
#493670000000
0#
0(
#493680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#493730000000
0$
0)
#493740000000
1"
1'
b0 +
b0 1
#493790000000
0"
0'
#493800000000
1#
1(
b101111101100100 +
b101111101100100 1
#493850000000
0#
0(
#493860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#493910000000
0$
0)
#493920000000
1"
1'
b0 +
b0 1
#493970000000
0"
0'
#493980000000
1#
1(
b101111101100100 +
b101111101100100 1
#494030000000
0#
0(
#494040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#494090000000
0$
0)
#494100000000
1"
1'
b0 +
b0 1
#494150000000
0"
0'
#494160000000
1#
1(
b101111101100100 +
b101111101100100 1
#494210000000
0#
0(
#494220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#494270000000
0$
0)
#494280000000
1"
1'
b0 +
b0 1
#494330000000
0"
0'
#494340000000
1#
1(
b101111101100100 +
b101111101100100 1
#494390000000
0#
0(
#494400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#494450000000
0$
0)
#494460000000
1"
1'
b0 +
b0 1
#494510000000
0"
0'
#494520000000
1#
1(
b101111101100100 +
b101111101100100 1
#494570000000
0#
0(
#494580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#494630000000
0$
0)
#494640000000
1"
1'
b0 +
b0 1
#494690000000
0"
0'
#494700000000
1#
1(
b101111101100100 +
b101111101100100 1
#494750000000
0#
0(
#494760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#494810000000
0$
0)
#494820000000
1"
1'
b0 +
b0 1
#494870000000
0"
0'
#494880000000
1#
1(
b101111101100100 +
b101111101100100 1
#494930000000
0#
0(
#494940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#494990000000
0$
0)
#495000000000
1"
1'
b0 +
b0 1
#495050000000
0"
0'
#495060000000
1#
1(
b101111101100100 +
b101111101100100 1
#495110000000
0#
0(
#495120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#495170000000
0$
0)
#495180000000
1"
1'
b0 +
b0 1
#495230000000
0"
0'
#495240000000
1#
1(
b101111101100100 +
b101111101100100 1
#495290000000
0#
0(
#495300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#495350000000
0$
0)
#495360000000
1"
1'
b0 +
b0 1
#495410000000
0"
0'
#495420000000
1#
1(
b101111101100100 +
b101111101100100 1
#495470000000
0#
0(
#495480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#495530000000
0$
0)
#495540000000
1"
1'
b0 +
b0 1
#495590000000
0"
0'
#495600000000
1#
1(
b101111101100100 +
b101111101100100 1
#495650000000
0#
0(
#495660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#495710000000
0$
0)
#495720000000
1"
1'
b0 +
b0 1
#495770000000
0"
0'
#495780000000
1#
1(
b101111101100100 +
b101111101100100 1
#495830000000
0#
0(
#495840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#495890000000
0$
0)
#495900000000
1"
1'
b0 +
b0 1
#495950000000
0"
0'
#495960000000
1#
1(
b101111101100100 +
b101111101100100 1
#496010000000
0#
0(
#496020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#496070000000
0$
0)
#496080000000
1"
1'
b0 +
b0 1
#496130000000
0"
0'
#496140000000
1#
1(
b101111101100100 +
b101111101100100 1
#496190000000
0#
0(
#496200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#496250000000
0$
0)
#496260000000
1"
1'
b0 +
b0 1
#496310000000
0"
0'
#496320000000
1#
1(
b101111101100100 +
b101111101100100 1
#496370000000
0#
0(
#496380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#496430000000
0$
0)
#496440000000
1"
1'
b0 +
b0 1
#496490000000
0"
0'
#496500000000
1#
1(
b101111101100100 +
b101111101100100 1
#496550000000
0#
0(
#496560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#496610000000
0$
0)
#496620000000
1"
1'
b0 +
b0 1
#496670000000
0"
0'
#496680000000
1#
1(
b101111101100100 +
b101111101100100 1
#496730000000
0#
0(
#496740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#496790000000
0$
0)
#496800000000
1"
1'
b0 +
b0 1
#496850000000
0"
0'
#496860000000
1#
1(
b101111101100100 +
b101111101100100 1
#496910000000
0#
0(
#496920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#496970000000
0$
0)
#496980000000
1"
1'
b0 +
b0 1
#497030000000
0"
0'
#497040000000
1#
1(
b101111101100100 +
b101111101100100 1
#497090000000
0#
0(
#497100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#497150000000
0$
0)
#497160000000
1"
1'
b0 +
b0 1
#497210000000
0"
0'
#497220000000
1#
1(
b101111101100100 +
b101111101100100 1
#497270000000
0#
0(
#497280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#497330000000
0$
0)
#497340000000
1"
1'
b0 +
b0 1
#497390000000
0"
0'
#497400000000
1#
1(
b101111101100100 +
b101111101100100 1
#497450000000
0#
0(
#497460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#497510000000
0$
0)
#497520000000
1"
1'
b0 +
b0 1
#497570000000
0"
0'
#497580000000
1#
1(
b101111101100100 +
b101111101100100 1
#497630000000
0#
0(
#497640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#497690000000
0$
0)
#497700000000
1"
1'
b0 +
b0 1
#497750000000
0"
0'
#497760000000
1#
1(
b101111101100100 +
b101111101100100 1
#497810000000
0#
0(
#497820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#497870000000
0$
0)
#497880000000
1"
1'
b0 +
b0 1
#497930000000
0"
0'
#497940000000
1#
1(
b101111101100100 +
b101111101100100 1
#497990000000
0#
0(
#498000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#498050000000
0$
0)
#498060000000
1"
1'
b0 +
b0 1
#498110000000
0"
0'
#498120000000
1#
1(
b101111101100100 +
b101111101100100 1
#498170000000
0#
0(
#498180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#498230000000
0$
0)
#498240000000
1"
1'
b0 +
b0 1
#498290000000
0"
0'
#498300000000
1#
1(
b101111101100100 +
b101111101100100 1
#498350000000
0#
0(
#498360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#498410000000
0$
0)
#498420000000
1"
1'
b0 +
b0 1
#498470000000
0"
0'
#498480000000
1#
1(
b101111101100100 +
b101111101100100 1
#498530000000
0#
0(
#498540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#498590000000
0$
0)
#498600000000
1"
1'
b0 +
b0 1
#498650000000
0"
0'
#498660000000
1#
1(
b101111101100100 +
b101111101100100 1
#498710000000
0#
0(
#498720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#498770000000
0$
0)
#498780000000
1"
1'
b0 +
b0 1
#498830000000
0"
0'
#498840000000
1#
1(
b101111101100100 +
b101111101100100 1
#498890000000
0#
0(
#498900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#498950000000
0$
0)
#498960000000
1"
1'
b0 +
b0 1
#499010000000
0"
0'
#499020000000
1#
1(
b101111101100100 +
b101111101100100 1
#499070000000
0#
0(
#499080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#499130000000
0$
0)
#499140000000
1"
1'
b0 +
b0 1
#499190000000
0"
0'
#499200000000
1#
1(
b101111101100100 +
b101111101100100 1
#499250000000
0#
0(
#499260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#499310000000
0$
0)
#499320000000
1"
1'
b0 +
b0 1
#499370000000
0"
0'
#499380000000
1#
1(
b101111101100100 +
b101111101100100 1
#499430000000
0#
0(
#499440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#499490000000
0$
0)
#499500000000
1"
1'
b0 +
b0 1
#499550000000
0"
0'
#499560000000
1#
1(
b101111101100100 +
b101111101100100 1
#499610000000
0#
0(
#499620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#499670000000
0$
0)
#499680000000
1"
1'
b0 +
b0 1
#499730000000
0"
0'
#499740000000
1#
1(
b101111101100100 +
b101111101100100 1
#499790000000
0#
0(
#499800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#499850000000
0$
0)
#499860000000
1"
1'
b0 +
b0 1
#499910000000
0"
0'
#499920000000
1#
1(
b101111101100100 +
b101111101100100 1
#499970000000
0#
0(
#499980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#500030000000
0$
0)
#500040000000
1"
1'
b0 +
b0 1
#500090000000
0"
0'
#500100000000
1#
1(
b101111101100100 +
b101111101100100 1
#500150000000
0#
0(
#500160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#500210000000
0$
0)
#500220000000
1"
1'
b0 +
b0 1
#500270000000
0"
0'
#500280000000
1#
1(
b101111101100100 +
b101111101100100 1
#500330000000
0#
0(
#500340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#500390000000
0$
0)
#500400000000
1"
1'
b0 +
b0 1
#500450000000
0"
0'
#500460000000
1#
1(
b101111101100100 +
b101111101100100 1
#500510000000
0#
0(
#500520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#500570000000
0$
0)
#500580000000
1"
1'
b0 +
b0 1
#500630000000
0"
0'
#500640000000
1#
1(
b101111101100100 +
b101111101100100 1
#500690000000
0#
0(
#500700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#500750000000
0$
0)
#500760000000
1"
1'
b0 +
b0 1
#500810000000
0"
0'
#500820000000
1#
1(
b101111101100100 +
b101111101100100 1
#500870000000
0#
0(
#500880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#500930000000
0$
0)
#500940000000
1"
1'
b0 +
b0 1
#500990000000
0"
0'
#501000000000
1#
1(
b101111101100100 +
b101111101100100 1
#501050000000
0#
0(
#501060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#501110000000
0$
0)
#501120000000
1"
1'
b0 +
b0 1
#501170000000
0"
0'
#501180000000
1#
1(
b101111101100100 +
b101111101100100 1
#501230000000
0#
0(
#501240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#501290000000
0$
0)
#501300000000
1"
1'
b0 +
b0 1
#501350000000
0"
0'
#501360000000
1#
1(
b101111101100100 +
b101111101100100 1
#501410000000
0#
0(
#501420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#501470000000
0$
0)
#501480000000
1"
1'
b0 +
b0 1
#501530000000
0"
0'
#501540000000
1#
1(
b101111101100100 +
b101111101100100 1
#501590000000
0#
0(
#501600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#501650000000
0$
0)
#501660000000
1"
1'
b0 +
b0 1
#501710000000
0"
0'
#501720000000
1#
1(
b101111101100100 +
b101111101100100 1
#501770000000
0#
0(
#501780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#501830000000
0$
0)
#501840000000
1"
1'
b0 +
b0 1
#501890000000
0"
0'
#501900000000
1#
1(
b101111101100100 +
b101111101100100 1
#501950000000
0#
0(
#501960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#502010000000
0$
0)
#502020000000
1"
1'
b0 +
b0 1
#502070000000
0"
0'
#502080000000
1#
1(
b101111101100100 +
b101111101100100 1
#502130000000
0#
0(
#502140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#502190000000
0$
0)
#502200000000
1"
1'
b0 +
b0 1
#502250000000
0"
0'
#502260000000
1#
1(
b101111101100100 +
b101111101100100 1
#502310000000
0#
0(
#502320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#502370000000
0$
0)
#502380000000
1"
1'
b0 +
b0 1
#502430000000
0"
0'
#502440000000
1#
1(
b101111101100100 +
b101111101100100 1
#502490000000
0#
0(
#502500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#502550000000
0$
0)
#502560000000
1"
1'
b0 +
b0 1
#502610000000
0"
0'
#502620000000
1#
1(
b101111101100100 +
b101111101100100 1
#502670000000
0#
0(
#502680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#502730000000
0$
0)
#502740000000
1"
1'
b0 +
b0 1
#502790000000
0"
0'
#502800000000
1#
1(
b101111101100100 +
b101111101100100 1
#502850000000
0#
0(
#502860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#502910000000
0$
0)
#502920000000
1"
1'
b0 +
b0 1
#502970000000
0"
0'
#502980000000
1#
1(
b101111101100100 +
b101111101100100 1
#503030000000
0#
0(
#503040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#503090000000
0$
0)
#503100000000
1"
1'
b0 +
b0 1
#503150000000
0"
0'
#503160000000
1#
1(
b101111101100100 +
b101111101100100 1
#503210000000
0#
0(
#503220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#503270000000
0$
0)
#503280000000
1"
1'
b0 +
b0 1
#503330000000
0"
0'
#503340000000
1#
1(
b101111101100100 +
b101111101100100 1
#503390000000
0#
0(
#503400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#503450000000
0$
0)
#503460000000
1"
1'
b0 +
b0 1
#503510000000
0"
0'
#503520000000
1#
1(
b101111101100100 +
b101111101100100 1
#503570000000
0#
0(
#503580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#503630000000
0$
0)
#503640000000
1"
1'
b0 +
b0 1
#503690000000
0"
0'
#503700000000
1#
1(
b101111101100100 +
b101111101100100 1
#503750000000
0#
0(
#503760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#503810000000
0$
0)
#503820000000
1"
1'
b0 +
b0 1
#503870000000
0"
0'
#503880000000
1#
1(
b101111101100100 +
b101111101100100 1
#503930000000
0#
0(
#503940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#503990000000
0$
0)
#504000000000
1"
1'
b0 +
b0 1
#504050000000
0"
0'
#504060000000
1#
1(
b101111101100100 +
b101111101100100 1
#504110000000
0#
0(
#504120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#504170000000
0$
0)
#504180000000
1"
1'
b0 +
b0 1
#504230000000
0"
0'
#504240000000
1#
1(
b101111101100100 +
b101111101100100 1
#504290000000
0#
0(
#504300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#504350000000
0$
0)
#504360000000
1"
1'
b0 +
b0 1
#504410000000
0"
0'
#504420000000
1#
1(
b101111101100100 +
b101111101100100 1
#504470000000
0#
0(
#504480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#504530000000
0$
0)
#504540000000
1"
1'
b0 +
b0 1
#504590000000
0"
0'
#504600000000
1#
1(
b101111101100100 +
b101111101100100 1
#504650000000
0#
0(
#504660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#504710000000
0$
0)
#504720000000
1"
1'
b0 +
b0 1
#504770000000
0"
0'
#504780000000
1#
1(
b101111101100100 +
b101111101100100 1
#504830000000
0#
0(
#504840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#504890000000
0$
0)
#504900000000
1"
1'
b0 +
b0 1
#504950000000
0"
0'
#504960000000
1#
1(
b101111101100100 +
b101111101100100 1
#505010000000
0#
0(
#505020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#505070000000
0$
0)
#505080000000
1"
1'
b0 +
b0 1
#505130000000
0"
0'
#505140000000
1#
1(
b101111101100100 +
b101111101100100 1
#505190000000
0#
0(
#505200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#505250000000
0$
0)
#505260000000
1"
1'
b0 +
b0 1
#505310000000
0"
0'
#505320000000
1#
1(
b101111101100100 +
b101111101100100 1
#505370000000
0#
0(
#505380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#505430000000
0$
0)
#505440000000
1"
1'
b0 +
b0 1
#505490000000
0"
0'
#505500000000
1#
1(
b101111101100100 +
b101111101100100 1
#505550000000
0#
0(
#505560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#505610000000
0$
0)
#505620000000
1"
1'
b0 +
b0 1
#505670000000
0"
0'
#505680000000
1#
1(
b101111101100100 +
b101111101100100 1
#505730000000
0#
0(
#505740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#505790000000
0$
0)
#505800000000
1"
1'
b0 +
b0 1
#505850000000
0"
0'
#505860000000
1#
1(
b101111101100100 +
b101111101100100 1
#505910000000
0#
0(
#505920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#505970000000
0$
0)
#505980000000
1"
1'
b0 +
b0 1
#506030000000
0"
0'
#506040000000
1#
1(
b101111101100100 +
b101111101100100 1
#506090000000
0#
0(
#506100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#506150000000
0$
0)
#506160000000
1"
1'
b0 +
b0 1
#506210000000
0"
0'
#506220000000
1#
1(
b101111101100100 +
b101111101100100 1
#506270000000
0#
0(
#506280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#506330000000
0$
0)
#506340000000
1"
1'
b0 +
b0 1
#506390000000
0"
0'
#506400000000
1#
1(
b101111101100100 +
b101111101100100 1
#506450000000
0#
0(
#506460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#506510000000
0$
0)
#506520000000
1"
1'
b0 +
b0 1
#506570000000
0"
0'
#506580000000
1#
1(
b101111101100100 +
b101111101100100 1
#506630000000
0#
0(
#506640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#506690000000
0$
0)
#506700000000
1"
1'
b0 +
b0 1
#506750000000
0"
0'
#506760000000
1#
1(
b101111101100100 +
b101111101100100 1
#506810000000
0#
0(
#506820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#506870000000
0$
0)
#506880000000
1"
1'
b0 +
b0 1
#506930000000
0"
0'
#506940000000
1#
1(
b101111101100100 +
b101111101100100 1
#506990000000
0#
0(
#507000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#507050000000
0$
0)
#507060000000
1"
1'
b0 +
b0 1
#507110000000
0"
0'
#507120000000
1#
1(
b101111101100100 +
b101111101100100 1
#507170000000
0#
0(
#507180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#507230000000
0$
0)
#507240000000
1"
1'
b0 +
b0 1
#507290000000
0"
0'
#507300000000
1#
1(
b101111101100100 +
b101111101100100 1
#507350000000
0#
0(
#507360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#507410000000
0$
0)
#507420000000
1"
1'
b0 +
b0 1
#507470000000
0"
0'
#507480000000
1#
1(
b101111101100100 +
b101111101100100 1
#507530000000
0#
0(
#507540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#507590000000
0$
0)
#507600000000
1"
1'
b0 +
b0 1
#507650000000
0"
0'
#507660000000
1#
1(
b101111101100100 +
b101111101100100 1
#507710000000
0#
0(
#507720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#507770000000
0$
0)
#507780000000
1"
1'
b0 +
b0 1
#507830000000
0"
0'
#507840000000
1#
1(
b101111101100100 +
b101111101100100 1
#507890000000
0#
0(
#507900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#507950000000
0$
0)
#507960000000
1"
1'
b0 +
b0 1
#508010000000
0"
0'
#508020000000
1#
1(
b101111101100100 +
b101111101100100 1
#508070000000
0#
0(
#508080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#508130000000
0$
0)
#508140000000
1"
1'
b0 +
b0 1
#508190000000
0"
0'
#508200000000
1#
1(
b101111101100100 +
b101111101100100 1
#508250000000
0#
0(
#508260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#508310000000
0$
0)
#508320000000
1"
1'
b0 +
b0 1
#508370000000
0"
0'
#508380000000
1#
1(
b101111101100100 +
b101111101100100 1
#508430000000
0#
0(
#508440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#508490000000
0$
0)
#508500000000
1"
1'
b0 +
b0 1
#508550000000
0"
0'
#508560000000
1#
1(
b101111101100100 +
b101111101100100 1
#508610000000
0#
0(
#508620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#508670000000
0$
0)
#508680000000
1"
1'
b0 +
b0 1
#508730000000
0"
0'
#508740000000
1#
1(
b101111101100100 +
b101111101100100 1
#508790000000
0#
0(
#508800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#508850000000
0$
0)
#508860000000
1"
1'
b0 +
b0 1
#508910000000
0"
0'
#508920000000
1#
1(
b101111101100100 +
b101111101100100 1
#508970000000
0#
0(
#508980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#509030000000
0$
0)
#509040000000
1"
1'
b0 +
b0 1
#509090000000
0"
0'
#509100000000
1#
1(
b101111101100100 +
b101111101100100 1
#509150000000
0#
0(
#509160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#509210000000
0$
0)
#509220000000
1"
1'
b0 +
b0 1
#509270000000
0"
0'
#509280000000
1#
1(
b101111101100100 +
b101111101100100 1
#509330000000
0#
0(
#509340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#509390000000
0$
0)
#509400000000
1"
1'
b0 +
b0 1
#509450000000
0"
0'
#509460000000
1#
1(
b101111101100100 +
b101111101100100 1
#509510000000
0#
0(
#509520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#509570000000
0$
0)
#509580000000
1"
1'
b0 +
b0 1
#509630000000
0"
0'
#509640000000
1#
1(
b101111101100100 +
b101111101100100 1
#509690000000
0#
0(
#509700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#509750000000
0$
0)
#509760000000
1"
1'
b0 +
b0 1
#509810000000
0"
0'
#509820000000
1#
1(
b101111101100100 +
b101111101100100 1
#509870000000
0#
0(
#509880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#509930000000
0$
0)
#509940000000
1"
1'
b0 +
b0 1
#509990000000
0"
0'
#510000000000
1#
1(
b101111101100100 +
b101111101100100 1
#510050000000
0#
0(
#510060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#510110000000
0$
0)
#510120000000
1"
1'
b0 +
b0 1
#510170000000
0"
0'
#510180000000
1#
1(
b101111101100100 +
b101111101100100 1
#510230000000
0#
0(
#510240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#510290000000
0$
0)
#510300000000
1"
1'
b0 +
b0 1
#510350000000
0"
0'
#510360000000
1#
1(
b101111101100100 +
b101111101100100 1
#510410000000
0#
0(
#510420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#510470000000
0$
0)
#510480000000
1"
1'
b0 +
b0 1
#510530000000
0"
0'
#510540000000
1#
1(
b101111101100100 +
b101111101100100 1
#510590000000
0#
0(
#510600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#510650000000
0$
0)
#510660000000
1"
1'
b0 +
b0 1
#510710000000
0"
0'
#510720000000
1#
1(
b101111101100100 +
b101111101100100 1
#510770000000
0#
0(
#510780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#510830000000
0$
0)
#510840000000
1"
1'
b0 +
b0 1
#510890000000
0"
0'
#510900000000
1#
1(
b101111101100100 +
b101111101100100 1
#510950000000
0#
0(
#510960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#511010000000
0$
0)
#511020000000
1"
1'
b0 +
b0 1
#511070000000
0"
0'
#511080000000
1#
1(
b101111101100100 +
b101111101100100 1
#511130000000
0#
0(
#511140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#511190000000
0$
0)
#511200000000
1"
1'
b0 +
b0 1
#511250000000
0"
0'
#511260000000
1#
1(
b101111101100100 +
b101111101100100 1
#511310000000
0#
0(
#511320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#511370000000
0$
0)
#511380000000
1"
1'
b0 +
b0 1
#511430000000
0"
0'
#511440000000
1#
1(
b101111101100100 +
b101111101100100 1
#511490000000
0#
0(
#511500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#511550000000
0$
0)
#511560000000
1"
1'
b0 +
b0 1
#511610000000
0"
0'
#511620000000
1#
1(
b101111101100100 +
b101111101100100 1
#511670000000
0#
0(
#511680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#511730000000
0$
0)
#511740000000
1"
1'
b0 +
b0 1
#511790000000
0"
0'
#511800000000
1#
1(
b101111101100100 +
b101111101100100 1
#511850000000
0#
0(
#511860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#511910000000
0$
0)
#511920000000
1"
1'
b0 +
b0 1
#511970000000
0"
0'
#511980000000
1#
1(
b101111101100100 +
b101111101100100 1
#512030000000
0#
0(
#512040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#512090000000
0$
0)
#512100000000
1"
1'
b0 +
b0 1
#512150000000
0"
0'
#512160000000
1#
1(
b101111101100100 +
b101111101100100 1
#512210000000
0#
0(
#512220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#512270000000
0$
0)
#512280000000
1"
1'
b0 +
b0 1
#512330000000
0"
0'
#512340000000
1#
1(
b101111101100100 +
b101111101100100 1
#512390000000
0#
0(
#512400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#512450000000
0$
0)
#512460000000
1"
1'
b0 +
b0 1
#512510000000
0"
0'
#512520000000
1#
1(
b101111101100100 +
b101111101100100 1
#512570000000
0#
0(
#512580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#512630000000
0$
0)
#512640000000
1"
1'
b0 +
b0 1
#512690000000
0"
0'
#512700000000
1#
1(
b101111101100100 +
b101111101100100 1
#512750000000
0#
0(
#512760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#512810000000
0$
0)
#512820000000
1"
1'
b0 +
b0 1
#512870000000
0"
0'
#512880000000
1#
1(
b101111101100100 +
b101111101100100 1
#512930000000
0#
0(
#512940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#512990000000
0$
0)
#513000000000
1"
1'
b0 +
b0 1
#513050000000
0"
0'
#513060000000
1#
1(
b101111101100100 +
b101111101100100 1
#513110000000
0#
0(
#513120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#513170000000
0$
0)
#513180000000
1"
1'
b0 +
b0 1
#513230000000
0"
0'
#513240000000
1#
1(
b101111101100100 +
b101111101100100 1
#513290000000
0#
0(
#513300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#513350000000
0$
0)
#513360000000
1"
1'
b0 +
b0 1
#513410000000
0"
0'
#513420000000
1#
1(
b101111101100100 +
b101111101100100 1
#513470000000
0#
0(
#513480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#513530000000
0$
0)
#513540000000
1"
1'
b0 +
b0 1
#513590000000
0"
0'
#513600000000
1#
1(
b101111101100100 +
b101111101100100 1
#513650000000
0#
0(
#513660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#513710000000
0$
0)
#513720000000
1"
1'
b0 +
b0 1
#513770000000
0"
0'
#513780000000
1#
1(
b101111101100100 +
b101111101100100 1
#513830000000
0#
0(
#513840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#513890000000
0$
0)
#513900000000
1"
1'
b0 +
b0 1
#513950000000
0"
0'
#513960000000
1#
1(
b101111101100100 +
b101111101100100 1
#514010000000
0#
0(
#514020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#514070000000
0$
0)
#514080000000
1"
1'
b0 +
b0 1
#514130000000
0"
0'
#514140000000
1#
1(
b101111101100100 +
b101111101100100 1
#514190000000
0#
0(
#514200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#514250000000
0$
0)
#514260000000
1"
1'
b0 +
b0 1
#514310000000
0"
0'
#514320000000
1#
1(
b101111101100100 +
b101111101100100 1
#514370000000
0#
0(
#514380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#514430000000
0$
0)
#514440000000
1"
1'
b0 +
b0 1
#514490000000
0"
0'
#514500000000
1#
1(
b101111101100100 +
b101111101100100 1
#514550000000
0#
0(
#514560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#514610000000
0$
0)
#514620000000
1"
1'
b0 +
b0 1
#514670000000
0"
0'
#514680000000
1#
1(
b101111101100100 +
b101111101100100 1
#514730000000
0#
0(
#514740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#514790000000
0$
0)
#514800000000
1"
1'
b0 +
b0 1
#514850000000
0"
0'
#514860000000
1#
1(
b101111101100100 +
b101111101100100 1
#514910000000
0#
0(
#514920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#514970000000
0$
0)
#514980000000
1"
1'
b0 +
b0 1
#515030000000
0"
0'
#515040000000
1#
1(
b101111101100100 +
b101111101100100 1
#515090000000
0#
0(
#515100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#515150000000
0$
0)
#515160000000
1"
1'
b0 +
b0 1
#515210000000
0"
0'
#515220000000
1#
1(
b101111101100100 +
b101111101100100 1
#515270000000
0#
0(
#515280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#515330000000
0$
0)
#515340000000
1"
1'
b0 +
b0 1
#515390000000
0"
0'
#515400000000
1#
1(
b101111101100100 +
b101111101100100 1
#515450000000
0#
0(
#515460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#515510000000
0$
0)
#515520000000
1"
1'
b0 +
b0 1
#515570000000
0"
0'
#515580000000
1#
1(
b101111101100100 +
b101111101100100 1
#515630000000
0#
0(
#515640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#515690000000
0$
0)
#515700000000
1"
1'
b0 +
b0 1
#515750000000
0"
0'
#515760000000
1#
1(
b101111101100100 +
b101111101100100 1
#515810000000
0#
0(
#515820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#515870000000
0$
0)
#515880000000
1"
1'
b0 +
b0 1
#515930000000
0"
0'
#515940000000
1#
1(
b101111101100100 +
b101111101100100 1
#515990000000
0#
0(
#516000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#516050000000
0$
0)
#516060000000
1"
1'
b0 +
b0 1
#516110000000
0"
0'
#516120000000
1#
1(
b101111101100100 +
b101111101100100 1
#516170000000
0#
0(
#516180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#516230000000
0$
0)
#516240000000
1"
1'
b0 +
b0 1
#516290000000
0"
0'
#516300000000
1#
1(
b101111101100100 +
b101111101100100 1
#516350000000
0#
0(
#516360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#516410000000
0$
0)
#516420000000
1"
1'
b0 +
b0 1
#516470000000
0"
0'
#516480000000
1#
1(
b101111101100100 +
b101111101100100 1
#516530000000
0#
0(
#516540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#516590000000
0$
0)
#516600000000
1"
1'
b0 +
b0 1
#516650000000
0"
0'
#516660000000
1#
1(
b101111101100100 +
b101111101100100 1
#516710000000
0#
0(
#516720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#516770000000
0$
0)
#516780000000
1"
1'
b0 +
b0 1
#516830000000
0"
0'
#516840000000
1#
1(
b101111101100100 +
b101111101100100 1
#516890000000
0#
0(
#516900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#516950000000
0$
0)
#516960000000
1"
1'
b0 +
b0 1
#517010000000
0"
0'
#517020000000
1#
1(
b101111101100100 +
b101111101100100 1
#517070000000
0#
0(
#517080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#517130000000
0$
0)
#517140000000
1"
1'
b0 +
b0 1
#517190000000
0"
0'
#517200000000
1#
1(
b101111101100100 +
b101111101100100 1
#517250000000
0#
0(
#517260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#517310000000
0$
0)
#517320000000
1"
1'
b0 +
b0 1
#517370000000
0"
0'
#517380000000
1#
1(
b101111101100100 +
b101111101100100 1
#517430000000
0#
0(
#517440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#517490000000
0$
0)
#517500000000
1"
1'
b0 +
b0 1
#517550000000
0"
0'
#517560000000
1#
1(
b101111101100100 +
b101111101100100 1
#517610000000
0#
0(
#517620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#517670000000
0$
0)
#517680000000
1"
1'
b0 +
b0 1
#517730000000
0"
0'
#517740000000
1#
1(
b101111101100100 +
b101111101100100 1
#517790000000
0#
0(
#517800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#517850000000
0$
0)
#517860000000
1"
1'
b0 +
b0 1
#517910000000
0"
0'
#517920000000
1#
1(
b101111101100100 +
b101111101100100 1
#517970000000
0#
0(
#517980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#518030000000
0$
0)
#518040000000
1"
1'
b0 +
b0 1
#518090000000
0"
0'
#518100000000
1#
1(
b101111101100100 +
b101111101100100 1
#518150000000
0#
0(
#518160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#518210000000
0$
0)
#518220000000
1"
1'
b0 +
b0 1
#518270000000
0"
0'
#518280000000
1#
1(
b101111101100100 +
b101111101100100 1
#518330000000
0#
0(
#518340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#518390000000
0$
0)
#518400000000
1"
1'
b0 +
b0 1
#518450000000
0"
0'
#518460000000
1#
1(
b101111101100100 +
b101111101100100 1
#518510000000
0#
0(
#518520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#518570000000
0$
0)
#518580000000
1"
1'
b0 +
b0 1
#518630000000
0"
0'
#518640000000
1#
1(
b101111101100100 +
b101111101100100 1
#518690000000
0#
0(
#518700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#518750000000
0$
0)
#518760000000
1"
1'
b0 +
b0 1
#518810000000
0"
0'
#518820000000
1#
1(
b101111101100100 +
b101111101100100 1
#518870000000
0#
0(
#518880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#518930000000
0$
0)
#518940000000
1"
1'
b0 +
b0 1
#518990000000
0"
0'
#519000000000
1#
1(
b101111101100100 +
b101111101100100 1
#519050000000
0#
0(
#519060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#519110000000
0$
0)
#519120000000
1"
1'
b0 +
b0 1
#519170000000
0"
0'
#519180000000
1#
1(
b101111101100100 +
b101111101100100 1
#519230000000
0#
0(
#519240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#519290000000
0$
0)
#519300000000
1"
1'
b0 +
b0 1
#519350000000
0"
0'
#519360000000
1#
1(
b101111101100100 +
b101111101100100 1
#519410000000
0#
0(
#519420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#519470000000
0$
0)
#519480000000
1"
1'
b0 +
b0 1
#519530000000
0"
0'
#519540000000
1#
1(
b101111101100100 +
b101111101100100 1
#519590000000
0#
0(
#519600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#519650000000
0$
0)
#519660000000
1"
1'
b0 +
b0 1
#519710000000
0"
0'
#519720000000
1#
1(
b101111101100100 +
b101111101100100 1
#519770000000
0#
0(
#519780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#519830000000
0$
0)
#519840000000
1"
1'
b0 +
b0 1
#519890000000
0"
0'
#519900000000
1#
1(
b101111101100100 +
b101111101100100 1
#519950000000
0#
0(
#519960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#520010000000
0$
0)
#520020000000
1"
1'
b0 +
b0 1
#520070000000
0"
0'
#520080000000
1#
1(
b101111101100100 +
b101111101100100 1
#520130000000
0#
0(
#520140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#520190000000
0$
0)
#520200000000
1"
1'
b0 +
b0 1
#520250000000
0"
0'
#520260000000
1#
1(
b101111101100100 +
b101111101100100 1
#520310000000
0#
0(
#520320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#520370000000
0$
0)
#520380000000
1"
1'
b0 +
b0 1
#520430000000
0"
0'
#520440000000
1#
1(
b101111101100100 +
b101111101100100 1
#520490000000
0#
0(
#520500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#520550000000
0$
0)
#520560000000
1"
1'
b0 +
b0 1
#520610000000
0"
0'
#520620000000
1#
1(
b101111101100100 +
b101111101100100 1
#520670000000
0#
0(
#520680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#520730000000
0$
0)
#520740000000
1"
1'
b0 +
b0 1
#520790000000
0"
0'
#520800000000
1#
1(
b101111101100100 +
b101111101100100 1
#520850000000
0#
0(
#520860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#520910000000
0$
0)
#520920000000
1"
1'
b0 +
b0 1
#520970000000
0"
0'
#520980000000
1#
1(
b101111101100100 +
b101111101100100 1
#521030000000
0#
0(
#521040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#521090000000
0$
0)
#521100000000
1"
1'
b0 +
b0 1
#521150000000
0"
0'
#521160000000
1#
1(
b101111101100100 +
b101111101100100 1
#521210000000
0#
0(
#521220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#521270000000
0$
0)
#521280000000
1"
1'
b0 +
b0 1
#521330000000
0"
0'
#521340000000
1#
1(
b101111101100100 +
b101111101100100 1
#521390000000
0#
0(
#521400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#521450000000
0$
0)
#521460000000
1"
1'
b0 +
b0 1
#521510000000
0"
0'
#521520000000
1#
1(
b101111101100100 +
b101111101100100 1
#521570000000
0#
0(
#521580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#521630000000
0$
0)
#521640000000
1"
1'
b0 +
b0 1
#521690000000
0"
0'
#521700000000
1#
1(
b101111101100100 +
b101111101100100 1
#521750000000
0#
0(
#521760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#521810000000
0$
0)
#521820000000
1"
1'
b0 +
b0 1
#521870000000
0"
0'
#521880000000
1#
1(
b101111101100100 +
b101111101100100 1
#521930000000
0#
0(
#521940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#521990000000
0$
0)
#522000000000
1"
1'
b0 +
b0 1
#522050000000
0"
0'
#522060000000
1#
1(
b101111101100100 +
b101111101100100 1
#522110000000
0#
0(
#522120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#522170000000
0$
0)
#522180000000
1"
1'
b0 +
b0 1
#522230000000
0"
0'
#522240000000
1#
1(
b101111101100100 +
b101111101100100 1
#522290000000
0#
0(
#522300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#522350000000
0$
0)
#522360000000
1"
1'
b0 +
b0 1
#522410000000
0"
0'
#522420000000
1#
1(
b101111101100100 +
b101111101100100 1
#522470000000
0#
0(
#522480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#522530000000
0$
0)
#522540000000
1"
1'
b0 +
b0 1
#522590000000
0"
0'
#522600000000
1#
1(
b101111101100100 +
b101111101100100 1
#522650000000
0#
0(
#522660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#522710000000
0$
0)
#522720000000
1"
1'
b0 +
b0 1
#522770000000
0"
0'
#522780000000
1#
1(
b101111101100100 +
b101111101100100 1
#522830000000
0#
0(
#522840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#522890000000
0$
0)
#522900000000
1"
1'
b0 +
b0 1
#522950000000
0"
0'
#522960000000
1#
1(
b101111101100100 +
b101111101100100 1
#523010000000
0#
0(
#523020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#523070000000
0$
0)
#523080000000
1"
1'
b0 +
b0 1
#523130000000
0"
0'
#523140000000
1#
1(
b101111101100100 +
b101111101100100 1
#523190000000
0#
0(
#523200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#523250000000
0$
0)
#523260000000
1"
1'
b0 +
b0 1
#523310000000
0"
0'
#523320000000
1#
1(
b101111101100100 +
b101111101100100 1
#523370000000
0#
0(
#523380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#523430000000
0$
0)
#523440000000
1"
1'
b0 +
b0 1
#523490000000
0"
0'
#523500000000
1#
1(
b101111101100100 +
b101111101100100 1
#523550000000
0#
0(
#523560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#523610000000
0$
0)
#523620000000
1"
1'
b0 +
b0 1
#523670000000
0"
0'
#523680000000
1#
1(
b101111101100100 +
b101111101100100 1
#523730000000
0#
0(
#523740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#523790000000
0$
0)
#523800000000
1"
1'
b0 +
b0 1
#523850000000
0"
0'
#523860000000
1#
1(
b101111101100100 +
b101111101100100 1
#523910000000
0#
0(
#523920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#523970000000
0$
0)
#523980000000
1"
1'
b0 +
b0 1
#524030000000
0"
0'
#524040000000
1#
1(
b101111101100100 +
b101111101100100 1
#524090000000
0#
0(
#524100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#524150000000
0$
0)
#524160000000
1"
1'
b0 +
b0 1
#524210000000
0"
0'
#524220000000
1#
1(
b101111101100100 +
b101111101100100 1
#524270000000
0#
0(
#524280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#524330000000
0$
0)
#524340000000
1"
1'
b0 +
b0 1
#524390000000
0"
0'
#524400000000
1#
1(
b101111101100100 +
b101111101100100 1
#524450000000
0#
0(
#524460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#524510000000
0$
0)
#524520000000
1"
1'
b0 +
b0 1
#524570000000
0"
0'
#524580000000
1#
1(
b101111101100100 +
b101111101100100 1
#524630000000
0#
0(
#524640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#524690000000
0$
0)
#524700000000
1"
1'
b0 +
b0 1
#524750000000
0"
0'
#524760000000
1#
1(
b101111101100100 +
b101111101100100 1
#524810000000
0#
0(
#524820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#524870000000
0$
0)
#524880000000
1"
1'
b0 +
b0 1
#524930000000
0"
0'
#524940000000
1#
1(
b101111101100100 +
b101111101100100 1
#524990000000
0#
0(
#525000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#525050000000
0$
0)
#525060000000
1"
1'
b0 +
b0 1
#525110000000
0"
0'
#525120000000
1#
1(
b101111101100100 +
b101111101100100 1
#525170000000
0#
0(
#525180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#525230000000
0$
0)
#525240000000
1"
1'
b0 +
b0 1
#525290000000
0"
0'
#525300000000
1#
1(
b101111101100100 +
b101111101100100 1
#525350000000
0#
0(
#525360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#525410000000
0$
0)
#525420000000
1"
1'
b0 +
b0 1
#525470000000
0"
0'
#525480000000
1#
1(
b101111101100100 +
b101111101100100 1
#525530000000
0#
0(
#525540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#525590000000
0$
0)
#525600000000
1"
1'
b0 +
b0 1
#525650000000
0"
0'
#525660000000
1#
1(
b101111101100100 +
b101111101100100 1
#525710000000
0#
0(
#525720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#525770000000
0$
0)
#525780000000
1"
1'
b0 +
b0 1
#525830000000
0"
0'
#525840000000
1#
1(
b101111101100100 +
b101111101100100 1
#525890000000
0#
0(
#525900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#525950000000
0$
0)
#525960000000
1"
1'
b0 +
b0 1
#526010000000
0"
0'
#526020000000
1#
1(
b101111101100100 +
b101111101100100 1
#526070000000
0#
0(
#526080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#526130000000
0$
0)
#526140000000
1"
1'
b0 +
b0 1
#526190000000
0"
0'
#526200000000
1#
1(
b101111101100100 +
b101111101100100 1
#526250000000
0#
0(
#526260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#526310000000
0$
0)
#526320000000
1"
1'
b0 +
b0 1
#526370000000
0"
0'
#526380000000
1#
1(
b101111101100100 +
b101111101100100 1
#526430000000
0#
0(
#526440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#526490000000
0$
0)
#526500000000
1"
1'
b0 +
b0 1
#526550000000
0"
0'
#526560000000
1#
1(
b101111101100100 +
b101111101100100 1
#526610000000
0#
0(
#526620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#526670000000
0$
0)
#526680000000
1"
1'
b0 +
b0 1
#526730000000
0"
0'
#526740000000
1#
1(
b101111101100100 +
b101111101100100 1
#526790000000
0#
0(
#526800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#526850000000
0$
0)
#526860000000
1"
1'
b0 +
b0 1
#526910000000
0"
0'
#526920000000
1#
1(
b101111101100100 +
b101111101100100 1
#526970000000
0#
0(
#526980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#527030000000
0$
0)
#527040000000
1"
1'
b0 +
b0 1
#527090000000
0"
0'
#527100000000
1#
1(
b101111101100100 +
b101111101100100 1
#527150000000
0#
0(
#527160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#527210000000
0$
0)
#527220000000
1"
1'
b0 +
b0 1
#527270000000
0"
0'
#527280000000
1#
1(
b101111101100100 +
b101111101100100 1
#527330000000
0#
0(
#527340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#527390000000
0$
0)
#527400000000
1"
1'
b0 +
b0 1
#527450000000
0"
0'
#527460000000
1#
1(
b101111101100100 +
b101111101100100 1
#527510000000
0#
0(
#527520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#527570000000
0$
0)
#527580000000
1"
1'
b0 +
b0 1
#527630000000
0"
0'
#527640000000
1#
1(
b101111101100100 +
b101111101100100 1
#527690000000
0#
0(
#527700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#527750000000
0$
0)
#527760000000
1"
1'
b0 +
b0 1
#527810000000
0"
0'
#527820000000
1#
1(
b101111101100100 +
b101111101100100 1
#527870000000
0#
0(
#527880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#527930000000
0$
0)
#527940000000
1"
1'
b0 +
b0 1
#527990000000
0"
0'
#528000000000
1#
1(
b101111101100100 +
b101111101100100 1
#528050000000
0#
0(
#528060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#528110000000
0$
0)
#528120000000
1"
1'
b0 +
b0 1
#528170000000
0"
0'
#528180000000
1#
1(
b101111101100100 +
b101111101100100 1
#528230000000
0#
0(
#528240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#528290000000
0$
0)
#528300000000
1"
1'
b0 +
b0 1
#528350000000
0"
0'
#528360000000
1#
1(
b101111101100100 +
b101111101100100 1
#528410000000
0#
0(
#528420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#528470000000
0$
0)
#528480000000
1"
1'
b0 +
b0 1
#528530000000
0"
0'
#528540000000
1#
1(
b101111101100100 +
b101111101100100 1
#528590000000
0#
0(
#528600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#528650000000
0$
0)
#528660000000
1"
1'
b0 +
b0 1
#528710000000
0"
0'
#528720000000
1#
1(
b101111101100100 +
b101111101100100 1
#528770000000
0#
0(
#528780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#528830000000
0$
0)
#528840000000
1"
1'
b0 +
b0 1
#528890000000
0"
0'
#528900000000
1#
1(
b101111101100100 +
b101111101100100 1
#528950000000
0#
0(
#528960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#529010000000
0$
0)
#529020000000
1"
1'
b0 +
b0 1
#529070000000
0"
0'
#529080000000
1#
1(
b101111101100100 +
b101111101100100 1
#529130000000
0#
0(
#529140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#529190000000
0$
0)
#529200000000
1"
1'
b0 +
b0 1
#529250000000
0"
0'
#529260000000
1#
1(
b101111101100100 +
b101111101100100 1
#529310000000
0#
0(
#529320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#529370000000
0$
0)
#529380000000
1"
1'
b0 +
b0 1
#529430000000
0"
0'
#529440000000
1#
1(
b101111101100100 +
b101111101100100 1
#529490000000
0#
0(
#529500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#529550000000
0$
0)
#529560000000
1"
1'
b0 +
b0 1
#529610000000
0"
0'
#529620000000
1#
1(
b101111101100100 +
b101111101100100 1
#529670000000
0#
0(
#529680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#529730000000
0$
0)
#529740000000
1"
1'
b0 +
b0 1
#529790000000
0"
0'
#529800000000
1#
1(
b101111101100100 +
b101111101100100 1
#529850000000
0#
0(
#529860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#529910000000
0$
0)
#529920000000
1"
1'
b0 +
b0 1
#529970000000
0"
0'
#529980000000
1#
1(
b101111101100100 +
b101111101100100 1
#530030000000
0#
0(
#530040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#530090000000
0$
0)
#530100000000
1"
1'
b0 +
b0 1
#530150000000
0"
0'
#530160000000
1#
1(
b101111101100100 +
b101111101100100 1
#530210000000
0#
0(
#530220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#530270000000
0$
0)
#530280000000
1"
1'
b0 +
b0 1
#530330000000
0"
0'
#530340000000
1#
1(
b101111101100100 +
b101111101100100 1
#530390000000
0#
0(
#530400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#530450000000
0$
0)
#530460000000
1"
1'
b0 +
b0 1
#530510000000
0"
0'
#530520000000
1#
1(
b101111101100100 +
b101111101100100 1
#530570000000
0#
0(
#530580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#530630000000
0$
0)
#530640000000
1"
1'
b0 +
b0 1
#530690000000
0"
0'
#530700000000
1#
1(
b101111101100100 +
b101111101100100 1
#530750000000
0#
0(
#530760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#530810000000
0$
0)
#530820000000
1"
1'
b0 +
b0 1
#530870000000
0"
0'
#530880000000
1#
1(
b101111101100100 +
b101111101100100 1
#530930000000
0#
0(
#530940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#530990000000
0$
0)
#531000000000
1"
1'
b0 +
b0 1
#531050000000
0"
0'
#531060000000
1#
1(
b101111101100100 +
b101111101100100 1
#531110000000
0#
0(
#531120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#531170000000
0$
0)
#531180000000
1"
1'
b0 +
b0 1
#531230000000
0"
0'
#531240000000
1#
1(
b101111101100100 +
b101111101100100 1
#531290000000
0#
0(
#531300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#531350000000
0$
0)
#531360000000
1"
1'
b0 +
b0 1
#531410000000
0"
0'
#531420000000
1#
1(
b101111101100100 +
b101111101100100 1
#531470000000
0#
0(
#531480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#531530000000
0$
0)
#531540000000
1"
1'
b0 +
b0 1
#531590000000
0"
0'
#531600000000
1#
1(
b101111101100100 +
b101111101100100 1
#531650000000
0#
0(
#531660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#531710000000
0$
0)
#531720000000
1"
1'
b0 +
b0 1
#531770000000
0"
0'
#531780000000
1#
1(
b101111101100100 +
b101111101100100 1
#531830000000
0#
0(
#531840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#531890000000
0$
0)
#531900000000
1"
1'
b0 +
b0 1
#531950000000
0"
0'
#531960000000
1#
1(
b101111101100100 +
b101111101100100 1
#532010000000
0#
0(
#532020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#532070000000
0$
0)
#532080000000
1"
1'
b0 +
b0 1
#532130000000
0"
0'
#532140000000
1#
1(
b101111101100100 +
b101111101100100 1
#532190000000
0#
0(
#532200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#532250000000
0$
0)
#532260000000
1"
1'
b0 +
b0 1
#532310000000
0"
0'
#532320000000
1#
1(
b101111101100100 +
b101111101100100 1
#532370000000
0#
0(
#532380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#532430000000
0$
0)
#532440000000
1"
1'
b0 +
b0 1
#532490000000
0"
0'
#532500000000
1#
1(
b101111101100100 +
b101111101100100 1
#532550000000
0#
0(
#532560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#532610000000
0$
0)
#532620000000
1"
1'
b0 +
b0 1
#532670000000
0"
0'
#532680000000
1#
1(
b101111101100100 +
b101111101100100 1
#532730000000
0#
0(
#532740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#532790000000
0$
0)
#532800000000
1"
1'
b0 +
b0 1
#532850000000
0"
0'
#532860000000
1#
1(
b101111101100100 +
b101111101100100 1
#532910000000
0#
0(
#532920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#532970000000
0$
0)
#532980000000
1"
1'
b0 +
b0 1
#533030000000
0"
0'
#533040000000
1#
1(
b101111101100100 +
b101111101100100 1
#533090000000
0#
0(
#533100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#533150000000
0$
0)
#533160000000
1"
1'
b0 +
b0 1
#533210000000
0"
0'
#533220000000
1#
1(
b101111101100100 +
b101111101100100 1
#533270000000
0#
0(
#533280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#533330000000
0$
0)
#533340000000
1"
1'
b0 +
b0 1
#533390000000
0"
0'
#533400000000
1#
1(
b101111101100100 +
b101111101100100 1
#533450000000
0#
0(
#533460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#533510000000
0$
0)
#533520000000
1"
1'
b0 +
b0 1
#533570000000
0"
0'
#533580000000
1#
1(
b101111101100100 +
b101111101100100 1
#533630000000
0#
0(
#533640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#533690000000
0$
0)
#533700000000
1"
1'
b0 +
b0 1
#533750000000
0"
0'
#533760000000
1#
1(
b101111101100100 +
b101111101100100 1
#533810000000
0#
0(
#533820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#533870000000
0$
0)
#533880000000
1"
1'
b0 +
b0 1
#533930000000
0"
0'
#533940000000
1#
1(
b101111101100100 +
b101111101100100 1
#533990000000
0#
0(
#534000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#534050000000
0$
0)
#534060000000
1"
1'
b0 +
b0 1
#534110000000
0"
0'
#534120000000
1#
1(
b101111101100100 +
b101111101100100 1
#534170000000
0#
0(
#534180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#534230000000
0$
0)
#534240000000
1"
1'
b0 +
b0 1
#534290000000
0"
0'
#534300000000
1#
1(
b101111101100100 +
b101111101100100 1
#534350000000
0#
0(
#534360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#534410000000
0$
0)
#534420000000
1"
1'
b0 +
b0 1
#534470000000
0"
0'
#534480000000
1#
1(
b101111101100100 +
b101111101100100 1
#534530000000
0#
0(
#534540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#534590000000
0$
0)
#534600000000
1"
1'
b0 +
b0 1
#534650000000
0"
0'
#534660000000
1#
1(
b101111101100100 +
b101111101100100 1
#534710000000
0#
0(
#534720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#534770000000
0$
0)
#534780000000
1"
1'
b0 +
b0 1
#534830000000
0"
0'
#534840000000
1#
1(
b101111101100100 +
b101111101100100 1
#534890000000
0#
0(
#534900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#534950000000
0$
0)
#534960000000
1"
1'
b0 +
b0 1
#535010000000
0"
0'
#535020000000
1#
1(
b101111101100100 +
b101111101100100 1
#535070000000
0#
0(
#535080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#535130000000
0$
0)
#535140000000
1"
1'
b0 +
b0 1
#535190000000
0"
0'
#535200000000
1#
1(
b101111101100100 +
b101111101100100 1
#535250000000
0#
0(
#535260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#535310000000
0$
0)
#535320000000
1"
1'
b0 +
b0 1
#535370000000
0"
0'
#535380000000
1#
1(
b101111101100100 +
b101111101100100 1
#535430000000
0#
0(
#535440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#535490000000
0$
0)
#535500000000
1"
1'
b0 +
b0 1
#535550000000
0"
0'
#535560000000
1#
1(
b101111101100100 +
b101111101100100 1
#535610000000
0#
0(
#535620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#535670000000
0$
0)
#535680000000
1"
1'
b0 +
b0 1
#535730000000
0"
0'
#535740000000
1#
1(
b101111101100100 +
b101111101100100 1
#535790000000
0#
0(
#535800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#535850000000
0$
0)
#535860000000
1"
1'
b0 +
b0 1
#535910000000
0"
0'
#535920000000
1#
1(
b101111101100100 +
b101111101100100 1
#535970000000
0#
0(
#535980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#536030000000
0$
0)
#536040000000
1"
1'
b0 +
b0 1
#536090000000
0"
0'
#536100000000
1#
1(
b101111101100100 +
b101111101100100 1
#536150000000
0#
0(
#536160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#536210000000
0$
0)
#536220000000
1"
1'
b0 +
b0 1
#536270000000
0"
0'
#536280000000
1#
1(
b101111101100100 +
b101111101100100 1
#536330000000
0#
0(
#536340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#536390000000
0$
0)
#536400000000
1"
1'
b0 +
b0 1
#536450000000
0"
0'
#536460000000
1#
1(
b101111101100100 +
b101111101100100 1
#536510000000
0#
0(
#536520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#536570000000
0$
0)
#536580000000
1"
1'
b0 +
b0 1
#536630000000
0"
0'
#536640000000
1#
1(
b101111101100100 +
b101111101100100 1
#536690000000
0#
0(
#536700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#536750000000
0$
0)
#536760000000
1"
1'
b0 +
b0 1
#536810000000
0"
0'
#536820000000
1#
1(
b101111101100100 +
b101111101100100 1
#536870000000
0#
0(
#536880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#536930000000
0$
0)
#536940000000
1"
1'
b0 +
b0 1
#536990000000
0"
0'
#537000000000
1#
1(
b101111101100100 +
b101111101100100 1
#537050000000
0#
0(
#537060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#537110000000
0$
0)
#537120000000
1"
1'
b0 +
b0 1
#537170000000
0"
0'
#537180000000
1#
1(
b101111101100100 +
b101111101100100 1
#537230000000
0#
0(
#537240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#537290000000
0$
0)
#537300000000
1"
1'
b0 +
b0 1
#537350000000
0"
0'
#537360000000
1#
1(
b101111101100100 +
b101111101100100 1
#537410000000
0#
0(
#537420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#537470000000
0$
0)
#537480000000
1"
1'
b0 +
b0 1
#537530000000
0"
0'
#537540000000
1#
1(
b101111101100100 +
b101111101100100 1
#537590000000
0#
0(
#537600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#537650000000
0$
0)
#537660000000
1"
1'
b0 +
b0 1
#537710000000
0"
0'
#537720000000
1#
1(
b101111101100100 +
b101111101100100 1
#537770000000
0#
0(
#537780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#537830000000
0$
0)
#537840000000
1"
1'
b0 +
b0 1
#537890000000
0"
0'
#537900000000
1#
1(
b101111101100100 +
b101111101100100 1
#537950000000
0#
0(
#537960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#538010000000
0$
0)
#538020000000
1"
1'
b0 +
b0 1
#538070000000
0"
0'
#538080000000
1#
1(
b101111101100100 +
b101111101100100 1
#538130000000
0#
0(
#538140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#538190000000
0$
0)
#538200000000
1"
1'
b0 +
b0 1
#538250000000
0"
0'
#538260000000
1#
1(
b101111101100100 +
b101111101100100 1
#538310000000
0#
0(
#538320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#538370000000
0$
0)
#538380000000
1"
1'
b0 +
b0 1
#538430000000
0"
0'
#538440000000
1#
1(
b101111101100100 +
b101111101100100 1
#538490000000
0#
0(
#538500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#538550000000
0$
0)
#538560000000
1"
1'
b0 +
b0 1
#538610000000
0"
0'
#538620000000
1#
1(
b101111101100100 +
b101111101100100 1
#538670000000
0#
0(
#538680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#538730000000
0$
0)
#538740000000
1"
1'
b0 +
b0 1
#538790000000
0"
0'
#538800000000
1#
1(
b101111101100100 +
b101111101100100 1
#538850000000
0#
0(
#538860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#538910000000
0$
0)
#538920000000
1"
1'
b0 +
b0 1
#538970000000
0"
0'
#538980000000
1#
1(
b101111101100100 +
b101111101100100 1
#539030000000
0#
0(
#539040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#539090000000
0$
0)
#539100000000
1"
1'
b0 +
b0 1
#539150000000
0"
0'
#539160000000
1#
1(
b101111101100100 +
b101111101100100 1
#539210000000
0#
0(
#539220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#539270000000
0$
0)
#539280000000
1"
1'
b0 +
b0 1
#539330000000
0"
0'
#539340000000
1#
1(
b101111101100100 +
b101111101100100 1
#539390000000
0#
0(
#539400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#539450000000
0$
0)
#539460000000
1"
1'
b0 +
b0 1
#539510000000
0"
0'
#539520000000
1#
1(
b101111101100100 +
b101111101100100 1
#539570000000
0#
0(
#539580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#539630000000
0$
0)
#539640000000
1"
1'
b0 +
b0 1
#539690000000
0"
0'
#539700000000
1#
1(
b101111101100100 +
b101111101100100 1
#539750000000
0#
0(
#539760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#539810000000
0$
0)
#539820000000
1"
1'
b0 +
b0 1
#539870000000
0"
0'
#539880000000
1#
1(
b101111101100100 +
b101111101100100 1
#539930000000
0#
0(
#539940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#539990000000
0$
0)
#540000000000
1"
1'
b0 +
b0 1
#540050000000
0"
0'
#540060000000
1#
1(
b101111101100100 +
b101111101100100 1
#540110000000
0#
0(
#540120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#540170000000
0$
0)
#540180000000
1"
1'
b0 +
b0 1
#540230000000
0"
0'
#540240000000
1#
1(
b101111101100100 +
b101111101100100 1
#540290000000
0#
0(
#540300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#540350000000
0$
0)
#540360000000
1"
1'
b0 +
b0 1
#540410000000
0"
0'
#540420000000
1#
1(
b101111101100100 +
b101111101100100 1
#540470000000
0#
0(
#540480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#540530000000
0$
0)
#540540000000
1"
1'
b0 +
b0 1
#540590000000
0"
0'
#540600000000
1#
1(
b101111101100100 +
b101111101100100 1
#540650000000
0#
0(
#540660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#540710000000
0$
0)
#540720000000
1"
1'
b0 +
b0 1
#540770000000
0"
0'
#540780000000
1#
1(
b101111101100100 +
b101111101100100 1
#540830000000
0#
0(
#540840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#540890000000
0$
0)
#540900000000
1"
1'
b0 +
b0 1
#540950000000
0"
0'
#540960000000
1#
1(
b101111101100100 +
b101111101100100 1
#541010000000
0#
0(
#541020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#541070000000
0$
0)
#541080000000
1"
1'
b0 +
b0 1
#541130000000
0"
0'
#541140000000
1#
1(
b101111101100100 +
b101111101100100 1
#541190000000
0#
0(
#541200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#541250000000
0$
0)
#541260000000
1"
1'
b0 +
b0 1
#541310000000
0"
0'
#541320000000
1#
1(
b101111101100100 +
b101111101100100 1
#541370000000
0#
0(
#541380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#541430000000
0$
0)
#541440000000
1"
1'
b0 +
b0 1
#541490000000
0"
0'
#541500000000
1#
1(
b101111101100100 +
b101111101100100 1
#541550000000
0#
0(
#541560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#541610000000
0$
0)
#541620000000
1"
1'
b0 +
b0 1
#541670000000
0"
0'
#541680000000
1#
1(
b101111101100100 +
b101111101100100 1
#541730000000
0#
0(
#541740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#541790000000
0$
0)
#541800000000
1"
1'
b0 +
b0 1
#541850000000
0"
0'
#541860000000
1#
1(
b101111101100100 +
b101111101100100 1
#541910000000
0#
0(
#541920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#541970000000
0$
0)
#541980000000
1"
1'
b0 +
b0 1
#542030000000
0"
0'
#542040000000
1#
1(
b101111101100100 +
b101111101100100 1
#542090000000
0#
0(
#542100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#542150000000
0$
0)
#542160000000
1"
1'
b0 +
b0 1
#542210000000
0"
0'
#542220000000
1#
1(
b101111101100100 +
b101111101100100 1
#542270000000
0#
0(
#542280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#542330000000
0$
0)
#542340000000
1"
1'
b0 +
b0 1
#542390000000
0"
0'
#542400000000
1#
1(
b101111101100100 +
b101111101100100 1
#542450000000
0#
0(
#542460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#542510000000
0$
0)
#542520000000
1"
1'
b0 +
b0 1
#542570000000
0"
0'
#542580000000
1#
1(
b101111101100100 +
b101111101100100 1
#542630000000
0#
0(
#542640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#542690000000
0$
0)
#542700000000
1"
1'
b0 +
b0 1
#542750000000
0"
0'
#542760000000
1#
1(
b101111101100100 +
b101111101100100 1
#542810000000
0#
0(
#542820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#542870000000
0$
0)
#542880000000
1"
1'
b0 +
b0 1
#542930000000
0"
0'
#542940000000
1#
1(
b101111101100100 +
b101111101100100 1
#542990000000
0#
0(
#543000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#543050000000
0$
0)
#543060000000
1"
1'
b0 +
b0 1
#543110000000
0"
0'
#543120000000
1#
1(
b101111101100100 +
b101111101100100 1
#543170000000
0#
0(
#543180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#543230000000
0$
0)
#543240000000
1"
1'
b0 +
b0 1
#543290000000
0"
0'
#543300000000
1#
1(
b101111101100100 +
b101111101100100 1
#543350000000
0#
0(
#543360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#543410000000
0$
0)
#543420000000
1"
1'
b0 +
b0 1
#543470000000
0"
0'
#543480000000
1#
1(
b101111101100100 +
b101111101100100 1
#543530000000
0#
0(
#543540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#543590000000
0$
0)
#543600000000
1"
1'
b0 +
b0 1
#543650000000
0"
0'
#543660000000
1#
1(
b101111101100100 +
b101111101100100 1
#543710000000
0#
0(
#543720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#543770000000
0$
0)
#543780000000
1"
1'
b0 +
b0 1
#543830000000
0"
0'
#543840000000
1#
1(
b101111101100100 +
b101111101100100 1
#543890000000
0#
0(
#543900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#543950000000
0$
0)
#543960000000
1"
1'
b0 +
b0 1
#544010000000
0"
0'
#544020000000
1#
1(
b101111101100100 +
b101111101100100 1
#544070000000
0#
0(
#544080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#544130000000
0$
0)
#544140000000
1"
1'
b0 +
b0 1
#544190000000
0"
0'
#544200000000
1#
1(
b101111101100100 +
b101111101100100 1
#544250000000
0#
0(
#544260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#544310000000
0$
0)
#544320000000
1"
1'
b0 +
b0 1
#544370000000
0"
0'
#544380000000
1#
1(
b101111101100100 +
b101111101100100 1
#544430000000
0#
0(
#544440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#544490000000
0$
0)
#544500000000
1"
1'
b0 +
b0 1
#544550000000
0"
0'
#544560000000
1#
1(
b101111101100100 +
b101111101100100 1
#544610000000
0#
0(
#544620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#544670000000
0$
0)
#544680000000
1"
1'
b0 +
b0 1
#544730000000
0"
0'
#544740000000
1#
1(
b101111101100100 +
b101111101100100 1
#544790000000
0#
0(
#544800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#544850000000
0$
0)
#544860000000
1"
1'
b0 +
b0 1
#544910000000
0"
0'
#544920000000
1#
1(
b101111101100100 +
b101111101100100 1
#544970000000
0#
0(
#544980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#545030000000
0$
0)
#545040000000
1"
1'
b0 +
b0 1
#545090000000
0"
0'
#545100000000
1#
1(
b101111101100100 +
b101111101100100 1
#545150000000
0#
0(
#545160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#545210000000
0$
0)
#545220000000
1"
1'
b0 +
b0 1
#545270000000
0"
0'
#545280000000
1#
1(
b101111101100100 +
b101111101100100 1
#545330000000
0#
0(
#545340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#545390000000
0$
0)
#545400000000
1"
1'
b0 +
b0 1
#545450000000
0"
0'
#545460000000
1#
1(
b101111101100100 +
b101111101100100 1
#545510000000
0#
0(
#545520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#545570000000
0$
0)
#545580000000
1"
1'
b0 +
b0 1
#545630000000
0"
0'
#545640000000
1#
1(
b101111101100100 +
b101111101100100 1
#545690000000
0#
0(
#545700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#545750000000
0$
0)
#545760000000
1"
1'
b0 +
b0 1
#545810000000
0"
0'
#545820000000
1#
1(
b101111101100100 +
b101111101100100 1
#545870000000
0#
0(
#545880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#545930000000
0$
0)
#545940000000
1"
1'
b0 +
b0 1
#545990000000
0"
0'
#546000000000
1#
1(
b101111101100100 +
b101111101100100 1
#546050000000
0#
0(
#546060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#546110000000
0$
0)
#546120000000
1"
1'
b0 +
b0 1
#546170000000
0"
0'
#546180000000
1#
1(
b101111101100100 +
b101111101100100 1
#546230000000
0#
0(
#546240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#546290000000
0$
0)
#546300000000
1"
1'
b0 +
b0 1
#546350000000
0"
0'
#546360000000
1#
1(
b101111101100100 +
b101111101100100 1
#546410000000
0#
0(
#546420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#546470000000
0$
0)
#546480000000
1"
1'
b0 +
b0 1
#546530000000
0"
0'
#546540000000
1#
1(
b101111101100100 +
b101111101100100 1
#546590000000
0#
0(
#546600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#546650000000
0$
0)
#546660000000
1"
1'
b0 +
b0 1
#546710000000
0"
0'
#546720000000
1#
1(
b101111101100100 +
b101111101100100 1
#546770000000
0#
0(
#546780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#546830000000
0$
0)
#546840000000
1"
1'
b0 +
b0 1
#546890000000
0"
0'
#546900000000
1#
1(
b101111101100100 +
b101111101100100 1
#546950000000
0#
0(
#546960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#547010000000
0$
0)
#547020000000
1"
1'
b0 +
b0 1
#547070000000
0"
0'
#547080000000
1#
1(
b101111101100100 +
b101111101100100 1
#547130000000
0#
0(
#547140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#547190000000
0$
0)
#547200000000
1"
1'
b0 +
b0 1
#547250000000
0"
0'
#547260000000
1#
1(
b101111101100100 +
b101111101100100 1
#547310000000
0#
0(
#547320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#547370000000
0$
0)
#547380000000
1"
1'
b0 +
b0 1
#547430000000
0"
0'
#547440000000
1#
1(
b101111101100100 +
b101111101100100 1
#547490000000
0#
0(
#547500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#547550000000
0$
0)
#547560000000
1"
1'
b0 +
b0 1
#547610000000
0"
0'
#547620000000
1#
1(
b101111101100100 +
b101111101100100 1
#547670000000
0#
0(
#547680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#547730000000
0$
0)
#547740000000
1"
1'
b0 +
b0 1
#547790000000
0"
0'
#547800000000
1#
1(
b101111101100100 +
b101111101100100 1
#547850000000
0#
0(
#547860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#547910000000
0$
0)
#547920000000
1"
1'
b0 +
b0 1
#547970000000
0"
0'
#547980000000
1#
1(
b101111101100100 +
b101111101100100 1
#548030000000
0#
0(
#548040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#548090000000
0$
0)
#548100000000
1"
1'
b0 +
b0 1
#548150000000
0"
0'
#548160000000
1#
1(
b101111101100100 +
b101111101100100 1
#548210000000
0#
0(
#548220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#548270000000
0$
0)
#548280000000
1"
1'
b0 +
b0 1
#548330000000
0"
0'
#548340000000
1#
1(
b101111101100100 +
b101111101100100 1
#548390000000
0#
0(
#548400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#548450000000
0$
0)
#548460000000
1"
1'
b0 +
b0 1
#548510000000
0"
0'
#548520000000
1#
1(
b101111101100100 +
b101111101100100 1
#548570000000
0#
0(
#548580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#548630000000
0$
0)
#548640000000
1"
1'
b0 +
b0 1
#548690000000
0"
0'
#548700000000
1#
1(
b101111101100100 +
b101111101100100 1
#548750000000
0#
0(
#548760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#548810000000
0$
0)
#548820000000
1"
1'
b0 +
b0 1
#548870000000
0"
0'
#548880000000
1#
1(
b101111101100100 +
b101111101100100 1
#548930000000
0#
0(
#548940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#548990000000
0$
0)
#549000000000
1"
1'
b0 +
b0 1
#549050000000
0"
0'
#549060000000
1#
1(
b101111101100100 +
b101111101100100 1
#549110000000
0#
0(
#549120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#549170000000
0$
0)
#549180000000
1"
1'
b0 +
b0 1
#549230000000
0"
0'
#549240000000
1#
1(
b101111101100100 +
b101111101100100 1
#549290000000
0#
0(
#549300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#549350000000
0$
0)
#549360000000
1"
1'
b0 +
b0 1
#549410000000
0"
0'
#549420000000
1#
1(
b101111101100100 +
b101111101100100 1
#549470000000
0#
0(
#549480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#549530000000
0$
0)
#549540000000
1"
1'
b0 +
b0 1
#549590000000
0"
0'
#549600000000
1#
1(
b101111101100100 +
b101111101100100 1
#549650000000
0#
0(
#549660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#549710000000
0$
0)
#549720000000
1"
1'
b0 +
b0 1
#549770000000
0"
0'
#549780000000
1#
1(
b101111101100100 +
b101111101100100 1
#549830000000
0#
0(
#549840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#549890000000
0$
0)
#549900000000
1"
1'
b0 +
b0 1
#549950000000
0"
0'
#549960000000
1#
1(
b101111101100100 +
b101111101100100 1
#550010000000
0#
0(
#550020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#550070000000
0$
0)
#550080000000
1"
1'
b0 +
b0 1
#550130000000
0"
0'
#550140000000
1#
1(
b101111101100100 +
b101111101100100 1
#550190000000
0#
0(
#550200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#550250000000
0$
0)
#550260000000
1"
1'
b0 +
b0 1
#550310000000
0"
0'
#550320000000
1#
1(
b101111101100100 +
b101111101100100 1
#550370000000
0#
0(
#550380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#550430000000
0$
0)
#550440000000
1"
1'
b0 +
b0 1
#550490000000
0"
0'
#550500000000
1#
1(
b101111101100100 +
b101111101100100 1
#550550000000
0#
0(
#550560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#550610000000
0$
0)
#550620000000
1"
1'
b0 +
b0 1
#550670000000
0"
0'
#550680000000
1#
1(
b101111101100100 +
b101111101100100 1
#550730000000
0#
0(
#550740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#550790000000
0$
0)
#550800000000
1"
1'
b0 +
b0 1
#550850000000
0"
0'
#550860000000
1#
1(
b101111101100100 +
b101111101100100 1
#550910000000
0#
0(
#550920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#550970000000
0$
0)
#550980000000
1"
1'
b0 +
b0 1
#551030000000
0"
0'
#551040000000
1#
1(
b101111101100100 +
b101111101100100 1
#551090000000
0#
0(
#551100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#551150000000
0$
0)
#551160000000
1"
1'
b0 +
b0 1
#551210000000
0"
0'
#551220000000
1#
1(
b101111101100100 +
b101111101100100 1
#551270000000
0#
0(
#551280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#551330000000
0$
0)
#551340000000
1"
1'
b0 +
b0 1
#551390000000
0"
0'
#551400000000
1#
1(
b101111101100100 +
b101111101100100 1
#551450000000
0#
0(
#551460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#551510000000
0$
0)
#551520000000
1"
1'
b0 +
b0 1
#551570000000
0"
0'
#551580000000
1#
1(
b101111101100100 +
b101111101100100 1
#551630000000
0#
0(
#551640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#551690000000
0$
0)
#551700000000
1"
1'
b0 +
b0 1
#551750000000
0"
0'
#551760000000
1#
1(
b101111101100100 +
b101111101100100 1
#551810000000
0#
0(
#551820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#551870000000
0$
0)
#551880000000
1"
1'
b0 +
b0 1
#551930000000
0"
0'
#551940000000
1#
1(
b101111101100100 +
b101111101100100 1
#551990000000
0#
0(
#552000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#552050000000
0$
0)
#552060000000
1"
1'
b0 +
b0 1
#552110000000
0"
0'
#552120000000
1#
1(
b101111101100100 +
b101111101100100 1
#552170000000
0#
0(
#552180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#552230000000
0$
0)
#552240000000
1"
1'
b0 +
b0 1
#552290000000
0"
0'
#552300000000
1#
1(
b101111101100100 +
b101111101100100 1
#552350000000
0#
0(
#552360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#552410000000
0$
0)
#552420000000
1"
1'
b0 +
b0 1
#552470000000
0"
0'
#552480000000
1#
1(
b101111101100100 +
b101111101100100 1
#552530000000
0#
0(
#552540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#552590000000
0$
0)
#552600000000
1"
1'
b0 +
b0 1
#552650000000
0"
0'
#552660000000
1#
1(
b101111101100100 +
b101111101100100 1
#552710000000
0#
0(
#552720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#552770000000
0$
0)
#552780000000
1"
1'
b0 +
b0 1
#552830000000
0"
0'
#552840000000
1#
1(
b101111101100100 +
b101111101100100 1
#552890000000
0#
0(
#552900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#552950000000
0$
0)
#552960000000
1"
1'
b0 +
b0 1
#553010000000
0"
0'
#553020000000
1#
1(
b101111101100100 +
b101111101100100 1
#553070000000
0#
0(
#553080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#553130000000
0$
0)
#553140000000
1"
1'
b0 +
b0 1
#553190000000
0"
0'
#553200000000
1#
1(
b101111101100100 +
b101111101100100 1
#553250000000
0#
0(
#553260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#553310000000
0$
0)
#553320000000
1"
1'
b0 +
b0 1
#553370000000
0"
0'
#553380000000
1#
1(
b101111101100100 +
b101111101100100 1
#553430000000
0#
0(
#553440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#553490000000
0$
0)
#553500000000
1"
1'
b0 +
b0 1
#553550000000
0"
0'
#553560000000
1#
1(
b101111101100100 +
b101111101100100 1
#553610000000
0#
0(
#553620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#553670000000
0$
0)
#553680000000
1"
1'
b0 +
b0 1
#553730000000
0"
0'
#553740000000
1#
1(
b101111101100100 +
b101111101100100 1
#553790000000
0#
0(
#553800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#553850000000
0$
0)
#553860000000
1"
1'
b0 +
b0 1
#553910000000
0"
0'
#553920000000
1#
1(
b101111101100100 +
b101111101100100 1
#553970000000
0#
0(
#553980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#554030000000
0$
0)
#554040000000
1"
1'
b0 +
b0 1
#554090000000
0"
0'
#554100000000
1#
1(
b101111101100100 +
b101111101100100 1
#554150000000
0#
0(
#554160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#554210000000
0$
0)
#554220000000
1"
1'
b0 +
b0 1
#554270000000
0"
0'
#554280000000
1#
1(
b101111101100100 +
b101111101100100 1
#554330000000
0#
0(
#554340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#554390000000
0$
0)
#554400000000
1"
1'
b0 +
b0 1
#554450000000
0"
0'
#554460000000
1#
1(
b101111101100100 +
b101111101100100 1
#554510000000
0#
0(
#554520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#554570000000
0$
0)
#554580000000
1"
1'
b0 +
b0 1
#554630000000
0"
0'
#554640000000
1#
1(
b101111101100100 +
b101111101100100 1
#554690000000
0#
0(
#554700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#554750000000
0$
0)
#554760000000
1"
1'
b0 +
b0 1
#554810000000
0"
0'
#554820000000
1#
1(
b101111101100100 +
b101111101100100 1
#554870000000
0#
0(
#554880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#554930000000
0$
0)
#554940000000
1"
1'
b0 +
b0 1
#554990000000
0"
0'
#555000000000
1#
1(
b101111101100100 +
b101111101100100 1
#555050000000
0#
0(
#555060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#555110000000
0$
0)
#555120000000
1"
1'
b0 +
b0 1
#555170000000
0"
0'
#555180000000
1#
1(
b101111101100100 +
b101111101100100 1
#555230000000
0#
0(
#555240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#555290000000
0$
0)
#555300000000
1"
1'
b0 +
b0 1
#555350000000
0"
0'
#555360000000
1#
1(
b101111101100100 +
b101111101100100 1
#555410000000
0#
0(
#555420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#555470000000
0$
0)
#555480000000
1"
1'
b0 +
b0 1
#555530000000
0"
0'
#555540000000
1#
1(
b101111101100100 +
b101111101100100 1
#555590000000
0#
0(
#555600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#555650000000
0$
0)
#555660000000
1"
1'
b0 +
b0 1
#555710000000
0"
0'
#555720000000
1#
1(
b101111101100100 +
b101111101100100 1
#555770000000
0#
0(
#555780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#555830000000
0$
0)
#555840000000
1"
1'
b0 +
b0 1
#555890000000
0"
0'
#555900000000
1#
1(
b101111101100100 +
b101111101100100 1
#555950000000
0#
0(
#555960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#556010000000
0$
0)
#556020000000
1"
1'
b0 +
b0 1
#556070000000
0"
0'
#556080000000
1#
1(
b101111101100100 +
b101111101100100 1
#556130000000
0#
0(
#556140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#556190000000
0$
0)
#556200000000
1"
1'
b0 +
b0 1
#556250000000
0"
0'
#556260000000
1#
1(
b101111101100100 +
b101111101100100 1
#556310000000
0#
0(
#556320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#556370000000
0$
0)
#556380000000
1"
1'
b0 +
b0 1
#556430000000
0"
0'
#556440000000
1#
1(
b101111101100100 +
b101111101100100 1
#556490000000
0#
0(
#556500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#556550000000
0$
0)
#556560000000
1"
1'
b0 +
b0 1
#556610000000
0"
0'
#556620000000
1#
1(
b101111101100100 +
b101111101100100 1
#556670000000
0#
0(
#556680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#556730000000
0$
0)
#556740000000
1"
1'
b0 +
b0 1
#556790000000
0"
0'
#556800000000
1#
1(
b101111101100100 +
b101111101100100 1
#556850000000
0#
0(
#556860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#556910000000
0$
0)
#556920000000
1"
1'
b0 +
b0 1
#556970000000
0"
0'
#556980000000
1#
1(
b101111101100100 +
b101111101100100 1
#557030000000
0#
0(
#557040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#557090000000
0$
0)
#557100000000
1"
1'
b0 +
b0 1
#557150000000
0"
0'
#557160000000
1#
1(
b101111101100100 +
b101111101100100 1
#557210000000
0#
0(
#557220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#557270000000
0$
0)
#557280000000
1"
1'
b0 +
b0 1
#557330000000
0"
0'
#557340000000
1#
1(
b101111101100100 +
b101111101100100 1
#557390000000
0#
0(
#557400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#557450000000
0$
0)
#557460000000
1"
1'
b0 +
b0 1
#557510000000
0"
0'
#557520000000
1#
1(
b101111101100100 +
b101111101100100 1
#557570000000
0#
0(
#557580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#557630000000
0$
0)
#557640000000
1"
1'
b0 +
b0 1
#557690000000
0"
0'
#557700000000
1#
1(
b101111101100100 +
b101111101100100 1
#557750000000
0#
0(
#557760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#557810000000
0$
0)
#557820000000
1"
1'
b0 +
b0 1
#557870000000
0"
0'
#557880000000
1#
1(
b101111101100100 +
b101111101100100 1
#557930000000
0#
0(
#557940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#557990000000
0$
0)
#558000000000
1"
1'
b0 +
b0 1
#558050000000
0"
0'
#558060000000
1#
1(
b101111101100100 +
b101111101100100 1
#558110000000
0#
0(
#558120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#558170000000
0$
0)
#558180000000
1"
1'
b0 +
b0 1
#558230000000
0"
0'
#558240000000
1#
1(
b101111101100100 +
b101111101100100 1
#558290000000
0#
0(
#558300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#558350000000
0$
0)
#558360000000
1"
1'
b0 +
b0 1
#558410000000
0"
0'
#558420000000
1#
1(
b101111101100100 +
b101111101100100 1
#558470000000
0#
0(
#558480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#558530000000
0$
0)
#558540000000
1"
1'
b0 +
b0 1
#558590000000
0"
0'
#558600000000
1#
1(
b101111101100100 +
b101111101100100 1
#558650000000
0#
0(
#558660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#558710000000
0$
0)
#558720000000
1"
1'
b0 +
b0 1
#558770000000
0"
0'
#558780000000
1#
1(
b101111101100100 +
b101111101100100 1
#558830000000
0#
0(
#558840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#558890000000
0$
0)
#558900000000
1"
1'
b0 +
b0 1
#558950000000
0"
0'
#558960000000
1#
1(
b101111101100100 +
b101111101100100 1
#559010000000
0#
0(
#559020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#559070000000
0$
0)
#559080000000
1"
1'
b0 +
b0 1
#559130000000
0"
0'
#559140000000
1#
1(
b101111101100100 +
b101111101100100 1
#559190000000
0#
0(
#559200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#559250000000
0$
0)
#559260000000
1"
1'
b0 +
b0 1
#559310000000
0"
0'
#559320000000
1#
1(
b101111101100100 +
b101111101100100 1
#559370000000
0#
0(
#559380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#559430000000
0$
0)
#559440000000
1"
1'
b0 +
b0 1
#559490000000
0"
0'
#559500000000
1#
1(
b101111101100100 +
b101111101100100 1
#559550000000
0#
0(
#559560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#559610000000
0$
0)
#559620000000
1"
1'
b0 +
b0 1
#559670000000
0"
0'
#559680000000
1#
1(
b101111101100100 +
b101111101100100 1
#559730000000
0#
0(
#559740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#559790000000
0$
0)
#559800000000
1"
1'
b0 +
b0 1
#559850000000
0"
0'
#559860000000
1#
1(
b101111101100100 +
b101111101100100 1
#559910000000
0#
0(
#559920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#559970000000
0$
0)
#559980000000
1"
1'
b0 +
b0 1
#560030000000
0"
0'
#560040000000
1#
1(
b101111101100100 +
b101111101100100 1
#560090000000
0#
0(
#560100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#560150000000
0$
0)
#560160000000
1"
1'
b0 +
b0 1
#560210000000
0"
0'
#560220000000
1#
1(
b101111101100100 +
b101111101100100 1
#560270000000
0#
0(
#560280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#560330000000
0$
0)
#560340000000
1"
1'
b0 +
b0 1
#560390000000
0"
0'
#560400000000
1#
1(
b101111101100100 +
b101111101100100 1
#560450000000
0#
0(
#560460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#560510000000
0$
0)
#560520000000
1"
1'
b0 +
b0 1
#560570000000
0"
0'
#560580000000
1#
1(
b101111101100100 +
b101111101100100 1
#560630000000
0#
0(
#560640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#560690000000
0$
0)
#560700000000
1"
1'
b0 +
b0 1
#560750000000
0"
0'
#560760000000
1#
1(
b101111101100100 +
b101111101100100 1
#560810000000
0#
0(
#560820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#560870000000
0$
0)
#560880000000
1"
1'
b0 +
b0 1
#560930000000
0"
0'
#560940000000
1#
1(
b101111101100100 +
b101111101100100 1
#560990000000
0#
0(
#561000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#561050000000
0$
0)
#561060000000
1"
1'
b0 +
b0 1
#561110000000
0"
0'
#561120000000
1#
1(
b101111101100100 +
b101111101100100 1
#561170000000
0#
0(
#561180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#561230000000
0$
0)
#561240000000
1"
1'
b0 +
b0 1
#561290000000
0"
0'
#561300000000
1#
1(
b101111101100100 +
b101111101100100 1
#561350000000
0#
0(
#561360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#561410000000
0$
0)
#561420000000
1"
1'
b0 +
b0 1
#561470000000
0"
0'
#561480000000
1#
1(
b101111101100100 +
b101111101100100 1
#561530000000
0#
0(
#561540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#561590000000
0$
0)
#561600000000
1"
1'
b0 +
b0 1
#561650000000
0"
0'
#561660000000
1#
1(
b101111101100100 +
b101111101100100 1
#561710000000
0#
0(
#561720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#561770000000
0$
0)
#561780000000
1"
1'
b0 +
b0 1
#561830000000
0"
0'
#561840000000
1#
1(
b101111101100100 +
b101111101100100 1
#561890000000
0#
0(
#561900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#561950000000
0$
0)
#561960000000
1"
1'
b0 +
b0 1
#562010000000
0"
0'
#562020000000
1#
1(
b101111101100100 +
b101111101100100 1
#562070000000
0#
0(
#562080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#562130000000
0$
0)
#562140000000
1"
1'
b0 +
b0 1
#562190000000
0"
0'
#562200000000
1#
1(
b101111101100100 +
b101111101100100 1
#562250000000
0#
0(
#562260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#562310000000
0$
0)
#562320000000
1"
1'
b0 +
b0 1
#562370000000
0"
0'
#562380000000
1#
1(
b101111101100100 +
b101111101100100 1
#562430000000
0#
0(
#562440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#562490000000
0$
0)
#562500000000
1"
1'
b0 +
b0 1
#562550000000
0"
0'
#562560000000
1#
1(
b101111101100100 +
b101111101100100 1
#562610000000
0#
0(
#562620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#562670000000
0$
0)
#562680000000
1"
1'
b0 +
b0 1
#562730000000
0"
0'
#562740000000
1#
1(
b101111101100100 +
b101111101100100 1
#562790000000
0#
0(
#562800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#562850000000
0$
0)
#562860000000
1"
1'
b0 +
b0 1
#562910000000
0"
0'
#562920000000
1#
1(
b101111101100100 +
b101111101100100 1
#562970000000
0#
0(
#562980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#563030000000
0$
0)
#563040000000
1"
1'
b0 +
b0 1
#563090000000
0"
0'
#563100000000
1#
1(
b101111101100100 +
b101111101100100 1
#563150000000
0#
0(
#563160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#563210000000
0$
0)
#563220000000
1"
1'
b0 +
b0 1
#563270000000
0"
0'
#563280000000
1#
1(
b101111101100100 +
b101111101100100 1
#563330000000
0#
0(
#563340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#563390000000
0$
0)
#563400000000
1"
1'
b0 +
b0 1
#563450000000
0"
0'
#563460000000
1#
1(
b101111101100100 +
b101111101100100 1
#563510000000
0#
0(
#563520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#563570000000
0$
0)
#563580000000
1"
1'
b0 +
b0 1
#563630000000
0"
0'
#563640000000
1#
1(
b101111101100100 +
b101111101100100 1
#563690000000
0#
0(
#563700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#563750000000
0$
0)
#563760000000
1"
1'
b0 +
b0 1
#563810000000
0"
0'
#563820000000
1#
1(
b101111101100100 +
b101111101100100 1
#563870000000
0#
0(
#563880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#563930000000
0$
0)
#563940000000
1"
1'
b0 +
b0 1
#563990000000
0"
0'
#564000000000
1#
1(
b101111101100100 +
b101111101100100 1
#564050000000
0#
0(
#564060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#564110000000
0$
0)
#564120000000
1"
1'
b0 +
b0 1
#564170000000
0"
0'
#564180000000
1#
1(
b101111101100100 +
b101111101100100 1
#564230000000
0#
0(
#564240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#564290000000
0$
0)
#564300000000
1"
1'
b0 +
b0 1
#564350000000
0"
0'
#564360000000
1#
1(
b101111101100100 +
b101111101100100 1
#564410000000
0#
0(
#564420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#564470000000
0$
0)
#564480000000
1"
1'
b0 +
b0 1
#564530000000
0"
0'
#564540000000
1#
1(
b101111101100100 +
b101111101100100 1
#564590000000
0#
0(
#564600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#564650000000
0$
0)
#564660000000
1"
1'
b0 +
b0 1
#564710000000
0"
0'
#564720000000
1#
1(
b101111101100100 +
b101111101100100 1
#564770000000
0#
0(
#564780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#564830000000
0$
0)
#564840000000
1"
1'
b0 +
b0 1
#564890000000
0"
0'
#564900000000
1#
1(
b101111101100100 +
b101111101100100 1
#564950000000
0#
0(
#564960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#565010000000
0$
0)
#565020000000
1"
1'
b0 +
b0 1
#565070000000
0"
0'
#565080000000
1#
1(
b101111101100100 +
b101111101100100 1
#565130000000
0#
0(
#565140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#565190000000
0$
0)
#565200000000
1"
1'
b0 +
b0 1
#565250000000
0"
0'
#565260000000
1#
1(
b101111101100100 +
b101111101100100 1
#565310000000
0#
0(
#565320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#565370000000
0$
0)
#565380000000
1"
1'
b0 +
b0 1
#565430000000
0"
0'
#565440000000
1#
1(
b101111101100100 +
b101111101100100 1
#565490000000
0#
0(
#565500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#565550000000
0$
0)
#565560000000
1"
1'
b0 +
b0 1
#565610000000
0"
0'
#565620000000
1#
1(
b101111101100100 +
b101111101100100 1
#565670000000
0#
0(
#565680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#565730000000
0$
0)
#565740000000
1"
1'
b0 +
b0 1
#565790000000
0"
0'
#565800000000
1#
1(
b101111101100100 +
b101111101100100 1
#565850000000
0#
0(
#565860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#565910000000
0$
0)
#565920000000
1"
1'
b0 +
b0 1
#565970000000
0"
0'
#565980000000
1#
1(
b101111101100100 +
b101111101100100 1
#566030000000
0#
0(
#566040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#566090000000
0$
0)
#566100000000
1"
1'
b0 +
b0 1
#566150000000
0"
0'
#566160000000
1#
1(
b101111101100100 +
b101111101100100 1
#566210000000
0#
0(
#566220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#566270000000
0$
0)
#566280000000
1"
1'
b0 +
b0 1
#566330000000
0"
0'
#566340000000
1#
1(
b101111101100100 +
b101111101100100 1
#566390000000
0#
0(
#566400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#566450000000
0$
0)
#566460000000
1"
1'
b0 +
b0 1
#566510000000
0"
0'
#566520000000
1#
1(
b101111101100100 +
b101111101100100 1
#566570000000
0#
0(
#566580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#566630000000
0$
0)
#566640000000
1"
1'
b0 +
b0 1
#566690000000
0"
0'
#566700000000
1#
1(
b101111101100100 +
b101111101100100 1
#566750000000
0#
0(
#566760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#566810000000
0$
0)
#566820000000
1"
1'
b0 +
b0 1
#566870000000
0"
0'
#566880000000
1#
1(
b101111101100100 +
b101111101100100 1
#566930000000
0#
0(
#566940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#566990000000
0$
0)
#567000000000
1"
1'
b0 +
b0 1
#567050000000
0"
0'
#567060000000
1#
1(
b101111101100100 +
b101111101100100 1
#567110000000
0#
0(
#567120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#567170000000
0$
0)
#567180000000
1"
1'
b0 +
b0 1
#567230000000
0"
0'
#567240000000
1#
1(
b101111101100100 +
b101111101100100 1
#567290000000
0#
0(
#567300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#567350000000
0$
0)
#567360000000
1"
1'
b0 +
b0 1
#567410000000
0"
0'
#567420000000
1#
1(
b101111101100100 +
b101111101100100 1
#567470000000
0#
0(
#567480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#567530000000
0$
0)
#567540000000
1"
1'
b0 +
b0 1
#567590000000
0"
0'
#567600000000
1#
1(
b101111101100100 +
b101111101100100 1
#567650000000
0#
0(
#567660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#567710000000
0$
0)
#567720000000
1"
1'
b0 +
b0 1
#567770000000
0"
0'
#567780000000
1#
1(
b101111101100100 +
b101111101100100 1
#567830000000
0#
0(
#567840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#567890000000
0$
0)
#567900000000
1"
1'
b0 +
b0 1
#567950000000
0"
0'
#567960000000
1#
1(
b101111101100100 +
b101111101100100 1
#568010000000
0#
0(
#568020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#568070000000
0$
0)
#568080000000
1"
1'
b0 +
b0 1
#568130000000
0"
0'
#568140000000
1#
1(
b101111101100100 +
b101111101100100 1
#568190000000
0#
0(
#568200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#568250000000
0$
0)
#568260000000
1"
1'
b0 +
b0 1
#568310000000
0"
0'
#568320000000
1#
1(
b101111101100100 +
b101111101100100 1
#568370000000
0#
0(
#568380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#568430000000
0$
0)
#568440000000
1"
1'
b0 +
b0 1
#568490000000
0"
0'
#568500000000
1#
1(
b101111101100100 +
b101111101100100 1
#568550000000
0#
0(
#568560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#568610000000
0$
0)
#568620000000
1"
1'
b0 +
b0 1
#568670000000
0"
0'
#568680000000
1#
1(
b101111101100100 +
b101111101100100 1
#568730000000
0#
0(
#568740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#568790000000
0$
0)
#568800000000
1"
1'
b0 +
b0 1
#568850000000
0"
0'
#568860000000
1#
1(
b101111101100100 +
b101111101100100 1
#568910000000
0#
0(
#568920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#568970000000
0$
0)
#568980000000
1"
1'
b0 +
b0 1
#569030000000
0"
0'
#569040000000
1#
1(
b101111101100100 +
b101111101100100 1
#569090000000
0#
0(
#569100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#569150000000
0$
0)
#569160000000
1"
1'
b0 +
b0 1
#569210000000
0"
0'
#569220000000
1#
1(
b101111101100100 +
b101111101100100 1
#569270000000
0#
0(
#569280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#569330000000
0$
0)
#569340000000
1"
1'
b0 +
b0 1
#569390000000
0"
0'
#569400000000
1#
1(
b101111101100100 +
b101111101100100 1
#569450000000
0#
0(
#569460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#569510000000
0$
0)
#569520000000
1"
1'
b0 +
b0 1
#569570000000
0"
0'
#569580000000
1#
1(
b101111101100100 +
b101111101100100 1
#569630000000
0#
0(
#569640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#569690000000
0$
0)
#569700000000
1"
1'
b0 +
b0 1
#569750000000
0"
0'
#569760000000
1#
1(
b101111101100100 +
b101111101100100 1
#569810000000
0#
0(
#569820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#569870000000
0$
0)
#569880000000
1"
1'
b0 +
b0 1
#569930000000
0"
0'
#569940000000
1#
1(
b101111101100100 +
b101111101100100 1
#569990000000
0#
0(
#570000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#570050000000
0$
0)
#570060000000
1"
1'
b0 +
b0 1
#570110000000
0"
0'
#570120000000
1#
1(
b101111101100100 +
b101111101100100 1
#570170000000
0#
0(
#570180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#570230000000
0$
0)
#570240000000
1"
1'
b0 +
b0 1
#570290000000
0"
0'
#570300000000
1#
1(
b101111101100100 +
b101111101100100 1
#570350000000
0#
0(
#570360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#570410000000
0$
0)
#570420000000
1"
1'
b0 +
b0 1
#570470000000
0"
0'
#570480000000
1#
1(
b101111101100100 +
b101111101100100 1
#570530000000
0#
0(
#570540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#570590000000
0$
0)
#570600000000
1"
1'
b0 +
b0 1
#570650000000
0"
0'
#570660000000
1#
1(
b101111101100100 +
b101111101100100 1
#570710000000
0#
0(
#570720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#570770000000
0$
0)
#570780000000
1"
1'
b0 +
b0 1
#570830000000
0"
0'
#570840000000
1#
1(
b101111101100100 +
b101111101100100 1
#570890000000
0#
0(
#570900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#570950000000
0$
0)
#570960000000
1"
1'
b0 +
b0 1
#571010000000
0"
0'
#571020000000
1#
1(
b101111101100100 +
b101111101100100 1
#571070000000
0#
0(
#571080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#571130000000
0$
0)
#571140000000
1"
1'
b0 +
b0 1
#571190000000
0"
0'
#571200000000
1#
1(
b101111101100100 +
b101111101100100 1
#571250000000
0#
0(
#571260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#571310000000
0$
0)
#571320000000
1"
1'
b0 +
b0 1
#571370000000
0"
0'
#571380000000
1#
1(
b101111101100100 +
b101111101100100 1
#571430000000
0#
0(
#571440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#571490000000
0$
0)
#571500000000
1"
1'
b0 +
b0 1
#571550000000
0"
0'
#571560000000
1#
1(
b101111101100100 +
b101111101100100 1
#571610000000
0#
0(
#571620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#571670000000
0$
0)
#571680000000
1"
1'
b0 +
b0 1
#571730000000
0"
0'
#571740000000
1#
1(
b101111101100100 +
b101111101100100 1
#571790000000
0#
0(
#571800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#571850000000
0$
0)
#571860000000
1"
1'
b0 +
b0 1
#571910000000
0"
0'
#571920000000
1#
1(
b101111101100100 +
b101111101100100 1
#571970000000
0#
0(
#571980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#572030000000
0$
0)
#572040000000
1"
1'
b0 +
b0 1
#572090000000
0"
0'
#572100000000
1#
1(
b101111101100100 +
b101111101100100 1
#572150000000
0#
0(
#572160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#572210000000
0$
0)
#572220000000
1"
1'
b0 +
b0 1
#572270000000
0"
0'
#572280000000
1#
1(
b101111101100100 +
b101111101100100 1
#572330000000
0#
0(
#572340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#572390000000
0$
0)
#572400000000
1"
1'
b0 +
b0 1
#572450000000
0"
0'
#572460000000
1#
1(
b101111101100100 +
b101111101100100 1
#572510000000
0#
0(
#572520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#572570000000
0$
0)
#572580000000
1"
1'
b0 +
b0 1
#572630000000
0"
0'
#572640000000
1#
1(
b101111101100100 +
b101111101100100 1
#572690000000
0#
0(
#572700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#572750000000
0$
0)
#572760000000
1"
1'
b0 +
b0 1
#572810000000
0"
0'
#572820000000
1#
1(
b101111101100100 +
b101111101100100 1
#572870000000
0#
0(
#572880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#572930000000
0$
0)
#572940000000
1"
1'
b0 +
b0 1
#572990000000
0"
0'
#573000000000
1#
1(
b101111101100100 +
b101111101100100 1
#573050000000
0#
0(
#573060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#573110000000
0$
0)
#573120000000
1"
1'
b0 +
b0 1
#573170000000
0"
0'
#573180000000
1#
1(
b101111101100100 +
b101111101100100 1
#573230000000
0#
0(
#573240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#573290000000
0$
0)
#573300000000
1"
1'
b0 +
b0 1
#573350000000
0"
0'
#573360000000
1#
1(
b101111101100100 +
b101111101100100 1
#573410000000
0#
0(
#573420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#573470000000
0$
0)
#573480000000
1"
1'
b0 +
b0 1
#573530000000
0"
0'
#573540000000
1#
1(
b101111101100100 +
b101111101100100 1
#573590000000
0#
0(
#573600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#573650000000
0$
0)
#573660000000
1"
1'
b0 +
b0 1
#573710000000
0"
0'
#573720000000
1#
1(
b101111101100100 +
b101111101100100 1
#573770000000
0#
0(
#573780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#573830000000
0$
0)
#573840000000
1"
1'
b0 +
b0 1
#573890000000
0"
0'
#573900000000
1#
1(
b101111101100100 +
b101111101100100 1
#573950000000
0#
0(
#573960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#574010000000
0$
0)
#574020000000
1"
1'
b0 +
b0 1
#574070000000
0"
0'
#574080000000
1#
1(
b101111101100100 +
b101111101100100 1
#574130000000
0#
0(
#574140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#574190000000
0$
0)
#574200000000
1"
1'
b0 +
b0 1
#574250000000
0"
0'
#574260000000
1#
1(
b101111101100100 +
b101111101100100 1
#574310000000
0#
0(
#574320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#574370000000
0$
0)
#574380000000
1"
1'
b0 +
b0 1
#574430000000
0"
0'
#574440000000
1#
1(
b101111101100100 +
b101111101100100 1
#574490000000
0#
0(
#574500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#574550000000
0$
0)
#574560000000
1"
1'
b0 +
b0 1
#574610000000
0"
0'
#574620000000
1#
1(
b101111101100100 +
b101111101100100 1
#574670000000
0#
0(
#574680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#574730000000
0$
0)
#574740000000
1"
1'
b0 +
b0 1
#574790000000
0"
0'
#574800000000
1#
1(
b101111101100100 +
b101111101100100 1
#574850000000
0#
0(
#574860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#574910000000
0$
0)
#574920000000
1"
1'
b0 +
b0 1
#574970000000
0"
0'
#574980000000
1#
1(
b101111101100100 +
b101111101100100 1
#575030000000
0#
0(
#575040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#575090000000
0$
0)
#575100000000
1"
1'
b0 +
b0 1
#575150000000
0"
0'
#575160000000
1#
1(
b101111101100100 +
b101111101100100 1
#575210000000
0#
0(
#575220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#575270000000
0$
0)
#575280000000
1"
1'
b0 +
b0 1
#575330000000
0"
0'
#575340000000
1#
1(
b101111101100100 +
b101111101100100 1
#575390000000
0#
0(
#575400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#575450000000
0$
0)
#575460000000
1"
1'
b0 +
b0 1
#575510000000
0"
0'
#575520000000
1#
1(
b101111101100100 +
b101111101100100 1
#575570000000
0#
0(
#575580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#575630000000
0$
0)
#575640000000
1"
1'
b0 +
b0 1
#575690000000
0"
0'
#575700000000
1#
1(
b101111101100100 +
b101111101100100 1
#575750000000
0#
0(
#575760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#575810000000
0$
0)
#575820000000
1"
1'
b0 +
b0 1
#575870000000
0"
0'
#575880000000
1#
1(
b101111101100100 +
b101111101100100 1
#575930000000
0#
0(
#575940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#575990000000
0$
0)
#576000000000
1"
1'
b0 +
b0 1
#576050000000
0"
0'
#576060000000
1#
1(
b101111101100100 +
b101111101100100 1
#576110000000
0#
0(
#576120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#576170000000
0$
0)
#576180000000
1"
1'
b0 +
b0 1
#576230000000
0"
0'
#576240000000
1#
1(
b101111101100100 +
b101111101100100 1
#576290000000
0#
0(
#576300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#576350000000
0$
0)
#576360000000
1"
1'
b0 +
b0 1
#576410000000
0"
0'
#576420000000
1#
1(
b101111101100100 +
b101111101100100 1
#576470000000
0#
0(
#576480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#576530000000
0$
0)
#576540000000
1"
1'
b0 +
b0 1
#576590000000
0"
0'
#576600000000
1#
1(
b101111101100100 +
b101111101100100 1
#576650000000
0#
0(
#576660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#576710000000
0$
0)
#576720000000
1"
1'
b0 +
b0 1
#576770000000
0"
0'
#576780000000
1#
1(
b101111101100100 +
b101111101100100 1
#576830000000
0#
0(
#576840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#576890000000
0$
0)
#576900000000
1"
1'
b0 +
b0 1
#576950000000
0"
0'
#576960000000
1#
1(
b101111101100100 +
b101111101100100 1
#577010000000
0#
0(
#577020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#577070000000
0$
0)
#577080000000
1"
1'
b0 +
b0 1
#577130000000
0"
0'
#577140000000
1#
1(
b101111101100100 +
b101111101100100 1
#577190000000
0#
0(
#577200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#577250000000
0$
0)
#577260000000
1"
1'
b0 +
b0 1
#577310000000
0"
0'
#577320000000
1#
1(
b101111101100100 +
b101111101100100 1
#577370000000
0#
0(
#577380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#577430000000
0$
0)
#577440000000
1"
1'
b0 +
b0 1
#577490000000
0"
0'
#577500000000
1#
1(
b101111101100100 +
b101111101100100 1
#577550000000
0#
0(
#577560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#577610000000
0$
0)
#577620000000
1"
1'
b0 +
b0 1
#577670000000
0"
0'
#577680000000
1#
1(
b101111101100100 +
b101111101100100 1
#577730000000
0#
0(
#577740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#577790000000
0$
0)
#577800000000
1"
1'
b0 +
b0 1
#577850000000
0"
0'
#577860000000
1#
1(
b101111101100100 +
b101111101100100 1
#577910000000
0#
0(
#577920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#577970000000
0$
0)
#577980000000
1"
1'
b0 +
b0 1
#578030000000
0"
0'
#578040000000
1#
1(
b101111101100100 +
b101111101100100 1
#578090000000
0#
0(
#578100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#578150000000
0$
0)
#578160000000
1"
1'
b0 +
b0 1
#578210000000
0"
0'
#578220000000
1#
1(
b101111101100100 +
b101111101100100 1
#578270000000
0#
0(
#578280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#578330000000
0$
0)
#578340000000
1"
1'
b0 +
b0 1
#578390000000
0"
0'
#578400000000
1#
1(
b101111101100100 +
b101111101100100 1
#578450000000
0#
0(
#578460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#578510000000
0$
0)
#578520000000
1"
1'
b0 +
b0 1
#578570000000
0"
0'
#578580000000
1#
1(
b101111101100100 +
b101111101100100 1
#578630000000
0#
0(
#578640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#578690000000
0$
0)
#578700000000
1"
1'
b0 +
b0 1
#578750000000
0"
0'
#578760000000
1#
1(
b101111101100100 +
b101111101100100 1
#578810000000
0#
0(
#578820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#578870000000
0$
0)
#578880000000
1"
1'
b0 +
b0 1
#578930000000
0"
0'
#578940000000
1#
1(
b101111101100100 +
b101111101100100 1
#578990000000
0#
0(
#579000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#579050000000
0$
0)
#579060000000
1"
1'
b0 +
b0 1
#579110000000
0"
0'
#579120000000
1#
1(
b101111101100100 +
b101111101100100 1
#579170000000
0#
0(
#579180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#579230000000
0$
0)
#579240000000
1"
1'
b0 +
b0 1
#579290000000
0"
0'
#579300000000
1#
1(
b101111101100100 +
b101111101100100 1
#579350000000
0#
0(
#579360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#579410000000
0$
0)
#579420000000
1"
1'
b0 +
b0 1
#579470000000
0"
0'
#579480000000
1#
1(
b101111101100100 +
b101111101100100 1
#579530000000
0#
0(
#579540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#579590000000
0$
0)
#579600000000
1"
1'
b0 +
b0 1
#579650000000
0"
0'
#579660000000
1#
1(
b101111101100100 +
b101111101100100 1
#579710000000
0#
0(
#579720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#579770000000
0$
0)
#579780000000
1"
1'
b0 +
b0 1
#579830000000
0"
0'
#579840000000
1#
1(
b101111101100100 +
b101111101100100 1
#579890000000
0#
0(
#579900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#579950000000
0$
0)
#579960000000
1"
1'
b0 +
b0 1
#580010000000
0"
0'
#580020000000
1#
1(
b101111101100100 +
b101111101100100 1
#580070000000
0#
0(
#580080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#580130000000
0$
0)
#580140000000
1"
1'
b0 +
b0 1
#580190000000
0"
0'
#580200000000
1#
1(
b101111101100100 +
b101111101100100 1
#580250000000
0#
0(
#580260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#580310000000
0$
0)
#580320000000
1"
1'
b0 +
b0 1
#580370000000
0"
0'
#580380000000
1#
1(
b101111101100100 +
b101111101100100 1
#580430000000
0#
0(
#580440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#580490000000
0$
0)
#580500000000
1"
1'
b0 +
b0 1
#580550000000
0"
0'
#580560000000
1#
1(
b101111101100100 +
b101111101100100 1
#580610000000
0#
0(
#580620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#580670000000
0$
0)
#580680000000
1"
1'
b0 +
b0 1
#580730000000
0"
0'
#580740000000
1#
1(
b101111101100100 +
b101111101100100 1
#580790000000
0#
0(
#580800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#580850000000
0$
0)
#580860000000
1"
1'
b0 +
b0 1
#580910000000
0"
0'
#580920000000
1#
1(
b101111101100100 +
b101111101100100 1
#580970000000
0#
0(
#580980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#581030000000
0$
0)
#581040000000
1"
1'
b0 +
b0 1
#581090000000
0"
0'
#581100000000
1#
1(
b101111101100100 +
b101111101100100 1
#581150000000
0#
0(
#581160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#581210000000
0$
0)
#581220000000
1"
1'
b0 +
b0 1
#581270000000
0"
0'
#581280000000
1#
1(
b101111101100100 +
b101111101100100 1
#581330000000
0#
0(
#581340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#581390000000
0$
0)
#581400000000
1"
1'
b0 +
b0 1
#581450000000
0"
0'
#581460000000
1#
1(
b101111101100100 +
b101111101100100 1
#581510000000
0#
0(
#581520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#581570000000
0$
0)
#581580000000
1"
1'
b0 +
b0 1
#581630000000
0"
0'
#581640000000
1#
1(
b101111101100100 +
b101111101100100 1
#581690000000
0#
0(
#581700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#581750000000
0$
0)
#581760000000
1"
1'
b0 +
b0 1
#581810000000
0"
0'
#581820000000
1#
1(
b101111101100100 +
b101111101100100 1
#581870000000
0#
0(
#581880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#581930000000
0$
0)
#581940000000
1"
1'
b0 +
b0 1
#581990000000
0"
0'
#582000000000
1#
1(
b101111101100100 +
b101111101100100 1
#582050000000
0#
0(
#582060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#582110000000
0$
0)
#582120000000
1"
1'
b0 +
b0 1
#582170000000
0"
0'
#582180000000
1#
1(
b101111101100100 +
b101111101100100 1
#582230000000
0#
0(
#582240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#582290000000
0$
0)
#582300000000
1"
1'
b0 +
b0 1
#582350000000
0"
0'
#582360000000
1#
1(
b101111101100100 +
b101111101100100 1
#582410000000
0#
0(
#582420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#582470000000
0$
0)
#582480000000
1"
1'
b0 +
b0 1
#582530000000
0"
0'
#582540000000
1#
1(
b101111101100100 +
b101111101100100 1
#582590000000
0#
0(
#582600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#582650000000
0$
0)
#582660000000
1"
1'
b0 +
b0 1
#582710000000
0"
0'
#582720000000
1#
1(
b101111101100100 +
b101111101100100 1
#582770000000
0#
0(
#582780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#582830000000
0$
0)
#582840000000
1"
1'
b0 +
b0 1
#582890000000
0"
0'
#582900000000
1#
1(
b101111101100100 +
b101111101100100 1
#582950000000
0#
0(
#582960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#583010000000
0$
0)
#583020000000
1"
1'
b0 +
b0 1
#583070000000
0"
0'
#583080000000
1#
1(
b101111101100100 +
b101111101100100 1
#583130000000
0#
0(
#583140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#583190000000
0$
0)
#583200000000
1"
1'
b0 +
b0 1
#583250000000
0"
0'
#583260000000
1#
1(
b101111101100100 +
b101111101100100 1
#583310000000
0#
0(
#583320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#583370000000
0$
0)
#583380000000
1"
1'
b0 +
b0 1
#583430000000
0"
0'
#583440000000
1#
1(
b101111101100100 +
b101111101100100 1
#583490000000
0#
0(
#583500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#583550000000
0$
0)
#583560000000
1"
1'
b0 +
b0 1
#583610000000
0"
0'
#583620000000
1#
1(
b101111101100100 +
b101111101100100 1
#583670000000
0#
0(
#583680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#583730000000
0$
0)
#583740000000
1"
1'
b0 +
b0 1
#583790000000
0"
0'
#583800000000
1#
1(
b101111101100100 +
b101111101100100 1
#583850000000
0#
0(
#583860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#583910000000
0$
0)
#583920000000
1"
1'
b0 +
b0 1
#583970000000
0"
0'
#583980000000
1#
1(
b101111101100100 +
b101111101100100 1
#584030000000
0#
0(
#584040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#584090000000
0$
0)
#584100000000
1"
1'
b0 +
b0 1
#584150000000
0"
0'
#584160000000
1#
1(
b101111101100100 +
b101111101100100 1
#584210000000
0#
0(
#584220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#584270000000
0$
0)
#584280000000
1"
1'
b0 +
b0 1
#584330000000
0"
0'
#584340000000
1#
1(
b101111101100100 +
b101111101100100 1
#584390000000
0#
0(
#584400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#584450000000
0$
0)
#584460000000
1"
1'
b0 +
b0 1
#584510000000
0"
0'
#584520000000
1#
1(
b101111101100100 +
b101111101100100 1
#584570000000
0#
0(
#584580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#584630000000
0$
0)
#584640000000
1"
1'
b0 +
b0 1
#584690000000
0"
0'
#584700000000
1#
1(
b101111101100100 +
b101111101100100 1
#584750000000
0#
0(
#584760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#584810000000
0$
0)
#584820000000
1"
1'
b0 +
b0 1
#584870000000
0"
0'
#584880000000
1#
1(
b101111101100100 +
b101111101100100 1
#584930000000
0#
0(
#584940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#584990000000
0$
0)
#585000000000
1"
1'
b0 +
b0 1
#585050000000
0"
0'
#585060000000
1#
1(
b101111101100100 +
b101111101100100 1
#585110000000
0#
0(
#585120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#585170000000
0$
0)
#585180000000
1"
1'
b0 +
b0 1
#585230000000
0"
0'
#585240000000
1#
1(
b101111101100100 +
b101111101100100 1
#585290000000
0#
0(
#585300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#585350000000
0$
0)
#585360000000
1"
1'
b0 +
b0 1
#585410000000
0"
0'
#585420000000
1#
1(
b101111101100100 +
b101111101100100 1
#585470000000
0#
0(
#585480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#585530000000
0$
0)
#585540000000
1"
1'
b0 +
b0 1
#585590000000
0"
0'
#585600000000
1#
1(
b101111101100100 +
b101111101100100 1
#585650000000
0#
0(
#585660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#585710000000
0$
0)
#585720000000
1"
1'
b0 +
b0 1
#585770000000
0"
0'
#585780000000
1#
1(
b101111101100100 +
b101111101100100 1
#585830000000
0#
0(
#585840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#585890000000
0$
0)
#585900000000
1"
1'
b0 +
b0 1
#585950000000
0"
0'
#585960000000
1#
1(
b101111101100100 +
b101111101100100 1
#586010000000
0#
0(
#586020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#586070000000
0$
0)
#586080000000
1"
1'
b0 +
b0 1
#586130000000
0"
0'
#586140000000
1#
1(
b101111101100100 +
b101111101100100 1
#586190000000
0#
0(
#586200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#586250000000
0$
0)
#586260000000
1"
1'
b0 +
b0 1
#586310000000
0"
0'
#586320000000
1#
1(
b101111101100100 +
b101111101100100 1
#586370000000
0#
0(
#586380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#586430000000
0$
0)
#586440000000
1"
1'
b0 +
b0 1
#586490000000
0"
0'
#586500000000
1#
1(
b101111101100100 +
b101111101100100 1
#586550000000
0#
0(
#586560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#586610000000
0$
0)
#586620000000
1"
1'
b0 +
b0 1
#586670000000
0"
0'
#586680000000
1#
1(
b101111101100100 +
b101111101100100 1
#586730000000
0#
0(
#586740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#586790000000
0$
0)
#586800000000
1"
1'
b0 +
b0 1
#586850000000
0"
0'
#586860000000
1#
1(
b101111101100100 +
b101111101100100 1
#586910000000
0#
0(
#586920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#586970000000
0$
0)
#586980000000
1"
1'
b0 +
b0 1
#587030000000
0"
0'
#587040000000
1#
1(
b101111101100100 +
b101111101100100 1
#587090000000
0#
0(
#587100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#587150000000
0$
0)
#587160000000
1"
1'
b0 +
b0 1
#587210000000
0"
0'
#587220000000
1#
1(
b101111101100100 +
b101111101100100 1
#587270000000
0#
0(
#587280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#587330000000
0$
0)
#587340000000
1"
1'
b0 +
b0 1
#587390000000
0"
0'
#587400000000
1#
1(
b101111101100100 +
b101111101100100 1
#587450000000
0#
0(
#587460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#587510000000
0$
0)
#587520000000
1"
1'
b0 +
b0 1
#587570000000
0"
0'
#587580000000
1#
1(
b101111101100100 +
b101111101100100 1
#587630000000
0#
0(
#587640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#587690000000
0$
0)
#587700000000
1"
1'
b0 +
b0 1
#587750000000
0"
0'
#587760000000
1#
1(
b101111101100100 +
b101111101100100 1
#587810000000
0#
0(
#587820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#587870000000
0$
0)
#587880000000
1"
1'
b0 +
b0 1
#587930000000
0"
0'
#587940000000
1#
1(
b101111101100100 +
b101111101100100 1
#587990000000
0#
0(
#588000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#588050000000
0$
0)
#588060000000
1"
1'
b0 +
b0 1
#588110000000
0"
0'
#588120000000
1#
1(
b101111101100100 +
b101111101100100 1
#588170000000
0#
0(
#588180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#588230000000
0$
0)
#588240000000
1"
1'
b0 +
b0 1
#588290000000
0"
0'
#588300000000
1#
1(
b101111101100100 +
b101111101100100 1
#588350000000
0#
0(
#588360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#588410000000
0$
0)
#588420000000
1"
1'
b0 +
b0 1
#588470000000
0"
0'
#588480000000
1#
1(
b101111101100100 +
b101111101100100 1
#588530000000
0#
0(
#588540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#588590000000
0$
0)
#588600000000
1"
1'
b0 +
b0 1
#588650000000
0"
0'
#588660000000
1#
1(
b101111101100100 +
b101111101100100 1
#588710000000
0#
0(
#588720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#588770000000
0$
0)
#588780000000
1"
1'
b0 +
b0 1
#588830000000
0"
0'
#588840000000
1#
1(
b101111101100100 +
b101111101100100 1
#588890000000
0#
0(
#588900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#588950000000
0$
0)
#588960000000
1"
1'
b0 +
b0 1
#589010000000
0"
0'
#589020000000
1#
1(
b101111101100100 +
b101111101100100 1
#589070000000
0#
0(
#589080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#589130000000
0$
0)
#589140000000
1"
1'
b0 +
b0 1
#589190000000
0"
0'
#589200000000
1#
1(
b101111101100100 +
b101111101100100 1
#589250000000
0#
0(
#589260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#589310000000
0$
0)
#589320000000
1"
1'
b0 +
b0 1
#589370000000
0"
0'
#589380000000
1#
1(
b101111101100100 +
b101111101100100 1
#589430000000
0#
0(
#589440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#589490000000
0$
0)
#589500000000
1"
1'
b0 +
b0 1
#589550000000
0"
0'
#589560000000
1#
1(
b101111101100100 +
b101111101100100 1
#589610000000
0#
0(
#589620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#589670000000
0$
0)
#589680000000
1"
1'
b0 +
b0 1
#589730000000
0"
0'
#589740000000
1#
1(
b101111101100100 +
b101111101100100 1
#589790000000
0#
0(
#589800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#589850000000
0$
0)
#589860000000
1"
1'
b0 +
b0 1
#589910000000
0"
0'
#589920000000
1#
1(
b101111101100100 +
b101111101100100 1
#589970000000
0#
0(
#589980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#590030000000
0$
0)
#590040000000
1"
1'
b0 +
b0 1
#590090000000
0"
0'
#590100000000
1#
1(
b101111101100100 +
b101111101100100 1
#590150000000
0#
0(
#590160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#590210000000
0$
0)
#590220000000
1"
1'
b0 +
b0 1
#590270000000
0"
0'
#590280000000
1#
1(
b101111101100100 +
b101111101100100 1
#590330000000
0#
0(
#590340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#590390000000
0$
0)
#590400000000
1"
1'
b0 +
b0 1
#590450000000
0"
0'
#590460000000
1#
1(
b101111101100100 +
b101111101100100 1
#590510000000
0#
0(
#590520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#590570000000
0$
0)
#590580000000
1"
1'
b0 +
b0 1
#590630000000
0"
0'
#590640000000
1#
1(
b101111101100100 +
b101111101100100 1
#590690000000
0#
0(
#590700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#590750000000
0$
0)
#590760000000
1"
1'
b0 +
b0 1
#590810000000
0"
0'
#590820000000
1#
1(
b101111101100100 +
b101111101100100 1
#590870000000
0#
0(
#590880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#590930000000
0$
0)
#590940000000
1"
1'
b0 +
b0 1
#590990000000
0"
0'
#591000000000
1#
1(
b101111101100100 +
b101111101100100 1
#591050000000
0#
0(
#591060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#591110000000
0$
0)
#591120000000
1"
1'
b0 +
b0 1
#591170000000
0"
0'
#591180000000
1#
1(
b101111101100100 +
b101111101100100 1
#591230000000
0#
0(
#591240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#591290000000
0$
0)
#591300000000
1"
1'
b0 +
b0 1
#591350000000
0"
0'
#591360000000
1#
1(
b101111101100100 +
b101111101100100 1
#591410000000
0#
0(
#591420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#591470000000
0$
0)
#591480000000
1"
1'
b0 +
b0 1
#591530000000
0"
0'
#591540000000
1#
1(
b101111101100100 +
b101111101100100 1
#591590000000
0#
0(
#591600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#591650000000
0$
0)
#591660000000
1"
1'
b0 +
b0 1
#591710000000
0"
0'
#591720000000
1#
1(
b101111101100100 +
b101111101100100 1
#591770000000
0#
0(
#591780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#591830000000
0$
0)
#591840000000
1"
1'
b0 +
b0 1
#591890000000
0"
0'
#591900000000
1#
1(
b101111101100100 +
b101111101100100 1
#591950000000
0#
0(
#591960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#592010000000
0$
0)
#592020000000
1"
1'
b0 +
b0 1
#592070000000
0"
0'
#592080000000
1#
1(
b101111101100100 +
b101111101100100 1
#592130000000
0#
0(
#592140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#592190000000
0$
0)
#592200000000
1"
1'
b0 +
b0 1
#592250000000
0"
0'
#592260000000
1#
1(
b101111101100100 +
b101111101100100 1
#592310000000
0#
0(
#592320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#592370000000
0$
0)
#592380000000
1"
1'
b0 +
b0 1
#592430000000
0"
0'
#592440000000
1#
1(
b101111101100100 +
b101111101100100 1
#592490000000
0#
0(
#592500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#592550000000
0$
0)
#592560000000
1"
1'
b0 +
b0 1
#592610000000
0"
0'
#592620000000
1#
1(
b101111101100100 +
b101111101100100 1
#592670000000
0#
0(
#592680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#592730000000
0$
0)
#592740000000
1"
1'
b0 +
b0 1
#592790000000
0"
0'
#592800000000
1#
1(
b101111101100100 +
b101111101100100 1
#592850000000
0#
0(
#592860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#592910000000
0$
0)
#592920000000
1"
1'
b0 +
b0 1
#592970000000
0"
0'
#592980000000
1#
1(
b101111101100100 +
b101111101100100 1
#593030000000
0#
0(
#593040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#593090000000
0$
0)
#593100000000
1"
1'
b0 +
b0 1
#593150000000
0"
0'
#593160000000
1#
1(
b101111101100100 +
b101111101100100 1
#593210000000
0#
0(
#593220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#593270000000
0$
0)
#593280000000
1"
1'
b0 +
b0 1
#593330000000
0"
0'
#593340000000
1#
1(
b101111101100100 +
b101111101100100 1
#593390000000
0#
0(
#593400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#593450000000
0$
0)
#593460000000
1"
1'
b0 +
b0 1
#593510000000
0"
0'
#593520000000
1#
1(
b101111101100100 +
b101111101100100 1
#593570000000
0#
0(
#593580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#593630000000
0$
0)
#593640000000
1"
1'
b0 +
b0 1
#593690000000
0"
0'
#593700000000
1#
1(
b101111101100100 +
b101111101100100 1
#593750000000
0#
0(
#593760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#593810000000
0$
0)
#593820000000
1"
1'
b0 +
b0 1
#593870000000
0"
0'
#593880000000
1#
1(
b101111101100100 +
b101111101100100 1
#593930000000
0#
0(
#593940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#593990000000
0$
0)
#594000000000
1"
1'
b0 +
b0 1
#594050000000
0"
0'
#594060000000
1#
1(
b101111101100100 +
b101111101100100 1
#594110000000
0#
0(
#594120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#594170000000
0$
0)
#594180000000
1"
1'
b0 +
b0 1
#594230000000
0"
0'
#594240000000
1#
1(
b101111101100100 +
b101111101100100 1
#594290000000
0#
0(
#594300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#594350000000
0$
0)
#594360000000
1"
1'
b0 +
b0 1
#594410000000
0"
0'
#594420000000
1#
1(
b101111101100100 +
b101111101100100 1
#594470000000
0#
0(
#594480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#594530000000
0$
0)
#594540000000
1"
1'
b0 +
b0 1
#594590000000
0"
0'
#594600000000
1#
1(
b101111101100100 +
b101111101100100 1
#594650000000
0#
0(
#594660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#594710000000
0$
0)
#594720000000
1"
1'
b0 +
b0 1
#594770000000
0"
0'
#594780000000
1#
1(
b101111101100100 +
b101111101100100 1
#594830000000
0#
0(
#594840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#594890000000
0$
0)
#594900000000
1"
1'
b0 +
b0 1
#594950000000
0"
0'
#594960000000
1#
1(
b101111101100100 +
b101111101100100 1
#595010000000
0#
0(
#595020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#595070000000
0$
0)
#595080000000
1"
1'
b0 +
b0 1
#595130000000
0"
0'
#595140000000
1#
1(
b101111101100100 +
b101111101100100 1
#595190000000
0#
0(
#595200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#595250000000
0$
0)
#595260000000
1"
1'
b0 +
b0 1
#595310000000
0"
0'
#595320000000
1#
1(
b101111101100100 +
b101111101100100 1
#595370000000
0#
0(
#595380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#595430000000
0$
0)
#595440000000
1"
1'
b0 +
b0 1
#595490000000
0"
0'
#595500000000
1#
1(
b101111101100100 +
b101111101100100 1
#595550000000
0#
0(
#595560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#595610000000
0$
0)
#595620000000
1"
1'
b0 +
b0 1
#595670000000
0"
0'
#595680000000
1#
1(
b101111101100100 +
b101111101100100 1
#595730000000
0#
0(
#595740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#595790000000
0$
0)
#595800000000
1"
1'
b0 +
b0 1
#595850000000
0"
0'
#595860000000
1#
1(
b101111101100100 +
b101111101100100 1
#595910000000
0#
0(
#595920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#595970000000
0$
0)
#595980000000
1"
1'
b0 +
b0 1
#596030000000
0"
0'
#596040000000
1#
1(
b101111101100100 +
b101111101100100 1
#596090000000
0#
0(
#596100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#596150000000
0$
0)
#596160000000
1"
1'
b0 +
b0 1
#596210000000
0"
0'
#596220000000
1#
1(
b101111101100100 +
b101111101100100 1
#596270000000
0#
0(
#596280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#596330000000
0$
0)
#596340000000
1"
1'
b0 +
b0 1
#596390000000
0"
0'
#596400000000
1#
1(
b101111101100100 +
b101111101100100 1
#596450000000
0#
0(
#596460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#596510000000
0$
0)
#596520000000
1"
1'
b0 +
b0 1
#596570000000
0"
0'
#596580000000
1#
1(
b101111101100100 +
b101111101100100 1
#596630000000
0#
0(
#596640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#596690000000
0$
0)
#596700000000
1"
1'
b0 +
b0 1
#596750000000
0"
0'
#596760000000
1#
1(
b101111101100100 +
b101111101100100 1
#596810000000
0#
0(
#596820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#596870000000
0$
0)
#596880000000
1"
1'
b0 +
b0 1
#596930000000
0"
0'
#596940000000
1#
1(
b101111101100100 +
b101111101100100 1
#596990000000
0#
0(
#597000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#597050000000
0$
0)
#597060000000
1"
1'
b0 +
b0 1
#597110000000
0"
0'
#597120000000
1#
1(
b101111101100100 +
b101111101100100 1
#597170000000
0#
0(
#597180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#597230000000
0$
0)
#597240000000
1"
1'
b0 +
b0 1
#597290000000
0"
0'
#597300000000
1#
1(
b101111101100100 +
b101111101100100 1
#597350000000
0#
0(
#597360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#597410000000
0$
0)
#597420000000
1"
1'
b0 +
b0 1
#597470000000
0"
0'
#597480000000
1#
1(
b101111101100100 +
b101111101100100 1
#597530000000
0#
0(
#597540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#597590000000
0$
0)
#597600000000
1"
1'
b0 +
b0 1
#597650000000
0"
0'
#597660000000
1#
1(
b101111101100100 +
b101111101100100 1
#597710000000
0#
0(
#597720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#597770000000
0$
0)
#597780000000
1"
1'
b0 +
b0 1
#597830000000
0"
0'
#597840000000
1#
1(
b101111101100100 +
b101111101100100 1
#597890000000
0#
0(
#597900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#597950000000
0$
0)
#597960000000
1"
1'
b0 +
b0 1
#598010000000
0"
0'
#598020000000
1#
1(
b101111101100100 +
b101111101100100 1
#598070000000
0#
0(
#598080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#598130000000
0$
0)
#598140000000
1"
1'
b0 +
b0 1
#598190000000
0"
0'
#598200000000
1#
1(
b101111101100100 +
b101111101100100 1
#598250000000
0#
0(
#598260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#598310000000
0$
0)
#598320000000
1"
1'
b0 +
b0 1
#598370000000
0"
0'
#598380000000
1#
1(
b101111101100100 +
b101111101100100 1
#598430000000
0#
0(
#598440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#598490000000
0$
0)
#598500000000
1"
1'
b0 +
b0 1
#598550000000
0"
0'
#598560000000
1#
1(
b101111101100100 +
b101111101100100 1
#598610000000
0#
0(
#598620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#598670000000
0$
0)
#598680000000
1"
1'
b0 +
b0 1
#598730000000
0"
0'
#598740000000
1#
1(
b101111101100100 +
b101111101100100 1
#598790000000
0#
0(
#598800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#598850000000
0$
0)
#598860000000
1"
1'
b0 +
b0 1
#598910000000
0"
0'
#598920000000
1#
1(
b101111101100100 +
b101111101100100 1
#598970000000
0#
0(
#598980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#599030000000
0$
0)
#599040000000
1"
1'
b0 +
b0 1
#599090000000
0"
0'
#599100000000
1#
1(
b101111101100100 +
b101111101100100 1
#599150000000
0#
0(
#599160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#599210000000
0$
0)
#599220000000
1"
1'
b0 +
b0 1
#599270000000
0"
0'
#599280000000
1#
1(
b101111101100100 +
b101111101100100 1
#599330000000
0#
0(
#599340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#599390000000
0$
0)
#599400000000
1"
1'
b0 +
b0 1
#599450000000
0"
0'
#599460000000
1#
1(
b101111101100100 +
b101111101100100 1
#599510000000
0#
0(
#599520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#599570000000
0$
0)
#599580000000
1"
1'
b0 +
b0 1
#599630000000
0"
0'
#599640000000
1#
1(
b101111101100100 +
b101111101100100 1
#599690000000
0#
0(
#599700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#599750000000
0$
0)
#599760000000
1"
1'
b0 +
b0 1
#599810000000
0"
0'
#599820000000
1#
1(
b101111101100100 +
b101111101100100 1
#599870000000
0#
0(
#599880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#599930000000
0$
0)
#599940000000
1"
1'
b0 +
b0 1
#599990000000
0"
0'
#600000000000
1#
1(
b101111101100100 +
b101111101100100 1
#600050000000
0#
0(
#600060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#600110000000
0$
0)
#600120000000
1"
1'
b0 +
b0 1
#600170000000
0"
0'
#600180000000
1#
1(
b101111101100100 +
b101111101100100 1
#600230000000
0#
0(
#600240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#600290000000
0$
0)
#600300000000
1"
1'
b0 +
b0 1
#600350000000
0"
0'
#600360000000
1#
1(
b101111101100100 +
b101111101100100 1
#600410000000
0#
0(
#600420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#600470000000
0$
0)
#600480000000
1"
1'
b0 +
b0 1
#600530000000
0"
0'
#600540000000
1#
1(
b101111101100100 +
b101111101100100 1
#600590000000
0#
0(
#600600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#600650000000
0$
0)
#600660000000
1"
1'
b0 +
b0 1
#600710000000
0"
0'
#600720000000
1#
1(
b101111101100100 +
b101111101100100 1
#600770000000
0#
0(
#600780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#600830000000
0$
0)
#600840000000
1"
1'
b0 +
b0 1
#600890000000
0"
0'
#600900000000
1#
1(
b101111101100100 +
b101111101100100 1
#600950000000
0#
0(
#600960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#601010000000
0$
0)
#601020000000
1"
1'
b0 +
b0 1
#601070000000
0"
0'
#601080000000
1#
1(
b101111101100100 +
b101111101100100 1
#601130000000
0#
0(
#601140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#601190000000
0$
0)
#601200000000
1"
1'
b0 +
b0 1
#601250000000
0"
0'
#601260000000
1#
1(
b101111101100100 +
b101111101100100 1
#601310000000
0#
0(
#601320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#601370000000
0$
0)
#601380000000
1"
1'
b0 +
b0 1
#601430000000
0"
0'
#601440000000
1#
1(
b101111101100100 +
b101111101100100 1
#601490000000
0#
0(
#601500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#601550000000
0$
0)
#601560000000
1"
1'
b0 +
b0 1
#601610000000
0"
0'
#601620000000
1#
1(
b101111101100100 +
b101111101100100 1
#601670000000
0#
0(
#601680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#601730000000
0$
0)
#601740000000
1"
1'
b0 +
b0 1
#601790000000
0"
0'
#601800000000
1#
1(
b101111101100100 +
b101111101100100 1
#601850000000
0#
0(
#601860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#601910000000
0$
0)
#601920000000
1"
1'
b0 +
b0 1
#601970000000
0"
0'
#601980000000
1#
1(
b101111101100100 +
b101111101100100 1
#602030000000
0#
0(
#602040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#602090000000
0$
0)
#602100000000
1"
1'
b0 +
b0 1
#602150000000
0"
0'
#602160000000
1#
1(
b101111101100100 +
b101111101100100 1
#602210000000
0#
0(
#602220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#602270000000
0$
0)
#602280000000
1"
1'
b0 +
b0 1
#602330000000
0"
0'
#602340000000
1#
1(
b101111101100100 +
b101111101100100 1
#602390000000
0#
0(
#602400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#602450000000
0$
0)
#602460000000
1"
1'
b0 +
b0 1
#602510000000
0"
0'
#602520000000
1#
1(
b101111101100100 +
b101111101100100 1
#602570000000
0#
0(
#602580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#602630000000
0$
0)
#602640000000
1"
1'
b0 +
b0 1
#602690000000
0"
0'
#602700000000
1#
1(
b101111101100100 +
b101111101100100 1
#602750000000
0#
0(
#602760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#602810000000
0$
0)
#602820000000
1"
1'
b0 +
b0 1
#602870000000
0"
0'
#602880000000
1#
1(
b101111101100100 +
b101111101100100 1
#602930000000
0#
0(
#602940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#602990000000
0$
0)
#603000000000
1"
1'
b0 +
b0 1
#603050000000
0"
0'
#603060000000
1#
1(
b101111101100100 +
b101111101100100 1
#603110000000
0#
0(
#603120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#603170000000
0$
0)
#603180000000
1"
1'
b0 +
b0 1
#603230000000
0"
0'
#603240000000
1#
1(
b101111101100100 +
b101111101100100 1
#603290000000
0#
0(
#603300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#603350000000
0$
0)
#603360000000
1"
1'
b0 +
b0 1
#603410000000
0"
0'
#603420000000
1#
1(
b101111101100100 +
b101111101100100 1
#603470000000
0#
0(
#603480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#603530000000
0$
0)
#603540000000
1"
1'
b0 +
b0 1
#603590000000
0"
0'
#603600000000
1#
1(
b101111101100100 +
b101111101100100 1
#603650000000
0#
0(
#603660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#603710000000
0$
0)
#603720000000
1"
1'
b0 +
b0 1
#603770000000
0"
0'
#603780000000
1#
1(
b101111101100100 +
b101111101100100 1
#603830000000
0#
0(
#603840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#603890000000
0$
0)
#603900000000
1"
1'
b0 +
b0 1
#603950000000
0"
0'
#603960000000
1#
1(
b101111101100100 +
b101111101100100 1
#604010000000
0#
0(
#604020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#604070000000
0$
0)
#604080000000
1"
1'
b0 +
b0 1
#604130000000
0"
0'
#604140000000
1#
1(
b101111101100100 +
b101111101100100 1
#604190000000
0#
0(
#604200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#604250000000
0$
0)
#604260000000
1"
1'
b0 +
b0 1
#604310000000
0"
0'
#604320000000
1#
1(
b101111101100100 +
b101111101100100 1
#604370000000
0#
0(
#604380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#604430000000
0$
0)
#604440000000
1"
1'
b0 +
b0 1
#604490000000
0"
0'
#604500000000
1#
1(
b101111101100100 +
b101111101100100 1
#604550000000
0#
0(
#604560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#604610000000
0$
0)
#604620000000
1"
1'
b0 +
b0 1
#604670000000
0"
0'
#604680000000
1#
1(
b101111101100100 +
b101111101100100 1
#604730000000
0#
0(
#604740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#604790000000
0$
0)
#604800000000
1"
1'
b0 +
b0 1
#604850000000
0"
0'
#604860000000
1#
1(
b101111101100100 +
b101111101100100 1
#604910000000
0#
0(
#604920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#604970000000
0$
0)
#604980000000
1"
1'
b0 +
b0 1
#605030000000
0"
0'
#605040000000
1#
1(
b101111101100100 +
b101111101100100 1
#605090000000
0#
0(
#605100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#605150000000
0$
0)
#605160000000
1"
1'
b0 +
b0 1
#605210000000
0"
0'
#605220000000
1#
1(
b101111101100100 +
b101111101100100 1
#605270000000
0#
0(
#605280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#605330000000
0$
0)
#605340000000
1"
1'
b0 +
b0 1
#605390000000
0"
0'
#605400000000
1#
1(
b101111101100100 +
b101111101100100 1
#605450000000
0#
0(
#605460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#605510000000
0$
0)
#605520000000
1"
1'
b0 +
b0 1
#605570000000
0"
0'
#605580000000
1#
1(
b101111101100100 +
b101111101100100 1
#605630000000
0#
0(
#605640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#605690000000
0$
0)
#605700000000
1"
1'
b0 +
b0 1
#605750000000
0"
0'
#605760000000
1#
1(
b101111101100100 +
b101111101100100 1
#605810000000
0#
0(
#605820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#605870000000
0$
0)
#605880000000
1"
1'
b0 +
b0 1
#605930000000
0"
0'
#605940000000
1#
1(
b101111101100100 +
b101111101100100 1
#605990000000
0#
0(
#606000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#606050000000
0$
0)
#606060000000
1"
1'
b0 +
b0 1
#606110000000
0"
0'
#606120000000
1#
1(
b101111101100100 +
b101111101100100 1
#606170000000
0#
0(
#606180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#606230000000
0$
0)
#606240000000
1"
1'
b0 +
b0 1
#606290000000
0"
0'
#606300000000
1#
1(
b101111101100100 +
b101111101100100 1
#606350000000
0#
0(
#606360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#606410000000
0$
0)
#606420000000
1"
1'
b0 +
b0 1
#606470000000
0"
0'
#606480000000
1#
1(
b101111101100100 +
b101111101100100 1
#606530000000
0#
0(
#606540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#606590000000
0$
0)
#606600000000
1"
1'
b0 +
b0 1
#606650000000
0"
0'
#606660000000
1#
1(
b101111101100100 +
b101111101100100 1
#606710000000
0#
0(
#606720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#606770000000
0$
0)
#606780000000
1"
1'
b0 +
b0 1
#606830000000
0"
0'
#606840000000
1#
1(
b101111101100100 +
b101111101100100 1
#606890000000
0#
0(
#606900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#606950000000
0$
0)
#606960000000
1"
1'
b0 +
b0 1
#607010000000
0"
0'
#607020000000
1#
1(
b101111101100100 +
b101111101100100 1
#607070000000
0#
0(
#607080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#607130000000
0$
0)
#607140000000
1"
1'
b0 +
b0 1
#607190000000
0"
0'
#607200000000
1#
1(
b101111101100100 +
b101111101100100 1
#607250000000
0#
0(
#607260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#607310000000
0$
0)
#607320000000
1"
1'
b0 +
b0 1
#607370000000
0"
0'
#607380000000
1#
1(
b101111101100100 +
b101111101100100 1
#607430000000
0#
0(
#607440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#607490000000
0$
0)
#607500000000
1"
1'
b0 +
b0 1
#607550000000
0"
0'
#607560000000
1#
1(
b101111101100100 +
b101111101100100 1
#607610000000
0#
0(
#607620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#607670000000
0$
0)
#607680000000
1"
1'
b0 +
b0 1
#607730000000
0"
0'
#607740000000
1#
1(
b101111101100100 +
b101111101100100 1
#607790000000
0#
0(
#607800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#607850000000
0$
0)
#607860000000
1"
1'
b0 +
b0 1
#607910000000
0"
0'
#607920000000
1#
1(
b101111101100100 +
b101111101100100 1
#607970000000
0#
0(
#607980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#608030000000
0$
0)
#608040000000
1"
1'
b0 +
b0 1
#608090000000
0"
0'
#608100000000
1#
1(
b101111101100100 +
b101111101100100 1
#608150000000
0#
0(
#608160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#608210000000
0$
0)
#608220000000
1"
1'
b0 +
b0 1
#608270000000
0"
0'
#608280000000
1#
1(
b101111101100100 +
b101111101100100 1
#608330000000
0#
0(
#608340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#608390000000
0$
0)
#608400000000
1"
1'
b0 +
b0 1
#608450000000
0"
0'
#608460000000
1#
1(
b101111101100100 +
b101111101100100 1
#608510000000
0#
0(
#608520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#608570000000
0$
0)
#608580000000
1"
1'
b0 +
b0 1
#608630000000
0"
0'
#608640000000
1#
1(
b101111101100100 +
b101111101100100 1
#608690000000
0#
0(
#608700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#608750000000
0$
0)
#608760000000
1"
1'
b0 +
b0 1
#608810000000
0"
0'
#608820000000
1#
1(
b101111101100100 +
b101111101100100 1
#608870000000
0#
0(
#608880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#608930000000
0$
0)
#608940000000
1"
1'
b0 +
b0 1
#608990000000
0"
0'
#609000000000
1#
1(
b101111101100100 +
b101111101100100 1
#609050000000
0#
0(
#609060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#609110000000
0$
0)
#609120000000
1"
1'
b0 +
b0 1
#609170000000
0"
0'
#609180000000
1#
1(
b101111101100100 +
b101111101100100 1
#609230000000
0#
0(
#609240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#609290000000
0$
0)
#609300000000
1"
1'
b0 +
b0 1
#609350000000
0"
0'
#609360000000
1#
1(
b101111101100100 +
b101111101100100 1
#609410000000
0#
0(
#609420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#609470000000
0$
0)
#609480000000
1"
1'
b0 +
b0 1
#609530000000
0"
0'
#609540000000
1#
1(
b101111101100100 +
b101111101100100 1
#609590000000
0#
0(
#609600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#609650000000
0$
0)
#609660000000
1"
1'
b0 +
b0 1
#609710000000
0"
0'
#609720000000
1#
1(
b101111101100100 +
b101111101100100 1
#609770000000
0#
0(
#609780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#609830000000
0$
0)
#609840000000
1"
1'
b0 +
b0 1
#609890000000
0"
0'
#609900000000
1#
1(
b101111101100100 +
b101111101100100 1
#609950000000
0#
0(
#609960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#610010000000
0$
0)
#610020000000
1"
1'
b0 +
b0 1
#610070000000
0"
0'
#610080000000
1#
1(
b101111101100100 +
b101111101100100 1
#610130000000
0#
0(
#610140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#610190000000
0$
0)
#610200000000
1"
1'
b0 +
b0 1
#610250000000
0"
0'
#610260000000
1#
1(
b101111101100100 +
b101111101100100 1
#610310000000
0#
0(
#610320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#610370000000
0$
0)
#610380000000
1"
1'
b0 +
b0 1
#610430000000
0"
0'
#610440000000
1#
1(
b101111101100100 +
b101111101100100 1
#610490000000
0#
0(
#610500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#610550000000
0$
0)
#610560000000
1"
1'
b0 +
b0 1
#610610000000
0"
0'
#610620000000
1#
1(
b101111101100100 +
b101111101100100 1
#610670000000
0#
0(
#610680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#610730000000
0$
0)
#610740000000
1"
1'
b0 +
b0 1
#610790000000
0"
0'
#610800000000
1#
1(
b101111101100100 +
b101111101100100 1
#610850000000
0#
0(
#610860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#610910000000
0$
0)
#610920000000
1"
1'
b0 +
b0 1
#610970000000
0"
0'
#610980000000
1#
1(
b101111101100100 +
b101111101100100 1
#611030000000
0#
0(
#611040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#611090000000
0$
0)
#611100000000
1"
1'
b0 +
b0 1
#611150000000
0"
0'
#611160000000
1#
1(
b101111101100100 +
b101111101100100 1
#611210000000
0#
0(
#611220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#611270000000
0$
0)
#611280000000
1"
1'
b0 +
b0 1
#611330000000
0"
0'
#611340000000
1#
1(
b101111101100100 +
b101111101100100 1
#611390000000
0#
0(
#611400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#611450000000
0$
0)
#611460000000
1"
1'
b0 +
b0 1
#611510000000
0"
0'
#611520000000
1#
1(
b101111101100100 +
b101111101100100 1
#611570000000
0#
0(
#611580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#611630000000
0$
0)
#611640000000
1"
1'
b0 +
b0 1
#611690000000
0"
0'
#611700000000
1#
1(
b101111101100100 +
b101111101100100 1
#611750000000
0#
0(
#611760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#611810000000
0$
0)
#611820000000
1"
1'
b0 +
b0 1
#611870000000
0"
0'
#611880000000
1#
1(
b101111101100100 +
b101111101100100 1
#611930000000
0#
0(
#611940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#611990000000
0$
0)
#612000000000
1"
1'
b0 +
b0 1
#612050000000
0"
0'
#612060000000
1#
1(
b101111101100100 +
b101111101100100 1
#612110000000
0#
0(
#612120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#612170000000
0$
0)
#612180000000
1"
1'
b0 +
b0 1
#612230000000
0"
0'
#612240000000
1#
1(
b101111101100100 +
b101111101100100 1
#612290000000
0#
0(
#612300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#612350000000
0$
0)
#612360000000
1"
1'
b0 +
b0 1
#612410000000
0"
0'
#612420000000
1#
1(
b101111101100100 +
b101111101100100 1
#612470000000
0#
0(
#612480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#612530000000
0$
0)
#612540000000
1"
1'
b0 +
b0 1
#612590000000
0"
0'
#612600000000
1#
1(
b101111101100100 +
b101111101100100 1
#612650000000
0#
0(
#612660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#612710000000
0$
0)
#612720000000
1"
1'
b0 +
b0 1
#612770000000
0"
0'
#612780000000
1#
1(
b101111101100100 +
b101111101100100 1
#612830000000
0#
0(
#612840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#612890000000
0$
0)
#612900000000
1"
1'
b0 +
b0 1
#612950000000
0"
0'
#612960000000
1#
1(
b101111101100100 +
b101111101100100 1
#613010000000
0#
0(
#613020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#613070000000
0$
0)
#613080000000
1"
1'
b0 +
b0 1
#613130000000
0"
0'
#613140000000
1#
1(
b101111101100100 +
b101111101100100 1
#613190000000
0#
0(
#613200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#613250000000
0$
0)
#613260000000
1"
1'
b0 +
b0 1
#613310000000
0"
0'
#613320000000
1#
1(
b101111101100100 +
b101111101100100 1
#613370000000
0#
0(
#613380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#613430000000
0$
0)
#613440000000
1"
1'
b0 +
b0 1
#613490000000
0"
0'
#613500000000
1#
1(
b101111101100100 +
b101111101100100 1
#613550000000
0#
0(
#613560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#613610000000
0$
0)
#613620000000
1"
1'
b0 +
b0 1
#613670000000
0"
0'
#613680000000
1#
1(
b101111101100100 +
b101111101100100 1
#613730000000
0#
0(
#613740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#613790000000
0$
0)
#613800000000
1"
1'
b0 +
b0 1
#613850000000
0"
0'
#613860000000
1#
1(
b101111101100100 +
b101111101100100 1
#613910000000
0#
0(
#613920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#613970000000
0$
0)
#613980000000
1"
1'
b0 +
b0 1
#614030000000
0"
0'
#614040000000
1#
1(
b101111101100100 +
b101111101100100 1
#614090000000
0#
0(
#614100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#614150000000
0$
0)
#614160000000
1"
1'
b0 +
b0 1
#614210000000
0"
0'
#614220000000
1#
1(
b101111101100100 +
b101111101100100 1
#614270000000
0#
0(
#614280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#614330000000
0$
0)
#614340000000
1"
1'
b0 +
b0 1
#614390000000
0"
0'
#614400000000
1#
1(
b101111101100100 +
b101111101100100 1
#614450000000
0#
0(
#614460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#614510000000
0$
0)
#614520000000
1"
1'
b0 +
b0 1
#614570000000
0"
0'
#614580000000
1#
1(
b101111101100100 +
b101111101100100 1
#614630000000
0#
0(
#614640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#614690000000
0$
0)
#614700000000
1"
1'
b0 +
b0 1
#614750000000
0"
0'
#614760000000
1#
1(
b101111101100100 +
b101111101100100 1
#614810000000
0#
0(
#614820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#614870000000
0$
0)
#614880000000
1"
1'
b0 +
b0 1
#614930000000
0"
0'
#614940000000
1#
1(
b101111101100100 +
b101111101100100 1
#614990000000
0#
0(
#615000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#615050000000
0$
0)
#615060000000
1"
1'
b0 +
b0 1
#615110000000
0"
0'
#615120000000
1#
1(
b101111101100100 +
b101111101100100 1
#615170000000
0#
0(
#615180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#615230000000
0$
0)
#615240000000
1"
1'
b0 +
b0 1
#615290000000
0"
0'
#615300000000
1#
1(
b101111101100100 +
b101111101100100 1
#615350000000
0#
0(
#615360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#615410000000
0$
0)
#615420000000
1"
1'
b0 +
b0 1
#615470000000
0"
0'
#615480000000
1#
1(
b101111101100100 +
b101111101100100 1
#615530000000
0#
0(
#615540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#615590000000
0$
0)
#615600000000
1"
1'
b0 +
b0 1
#615650000000
0"
0'
#615660000000
1#
1(
b101111101100100 +
b101111101100100 1
#615710000000
0#
0(
#615720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#615770000000
0$
0)
#615780000000
1"
1'
b0 +
b0 1
#615830000000
0"
0'
#615840000000
1#
1(
b101111101100100 +
b101111101100100 1
#615890000000
0#
0(
#615900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#615950000000
0$
0)
#615960000000
1"
1'
b0 +
b0 1
#616010000000
0"
0'
#616020000000
1#
1(
b101111101100100 +
b101111101100100 1
#616070000000
0#
0(
#616080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#616130000000
0$
0)
#616140000000
1"
1'
b0 +
b0 1
#616190000000
0"
0'
#616200000000
1#
1(
b101111101100100 +
b101111101100100 1
#616250000000
0#
0(
#616260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#616310000000
0$
0)
#616320000000
1"
1'
b0 +
b0 1
#616370000000
0"
0'
#616380000000
1#
1(
b101111101100100 +
b101111101100100 1
#616430000000
0#
0(
#616440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#616490000000
0$
0)
#616500000000
1"
1'
b0 +
b0 1
#616550000000
0"
0'
#616560000000
1#
1(
b101111101100100 +
b101111101100100 1
#616610000000
0#
0(
#616620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#616670000000
0$
0)
#616680000000
1"
1'
b0 +
b0 1
#616730000000
0"
0'
#616740000000
1#
1(
b101111101100100 +
b101111101100100 1
#616790000000
0#
0(
#616800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#616850000000
0$
0)
#616860000000
1"
1'
b0 +
b0 1
#616910000000
0"
0'
#616920000000
1#
1(
b101111101100100 +
b101111101100100 1
#616970000000
0#
0(
#616980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#617030000000
0$
0)
#617040000000
1"
1'
b0 +
b0 1
#617090000000
0"
0'
#617100000000
1#
1(
b101111101100100 +
b101111101100100 1
#617150000000
0#
0(
#617160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#617210000000
0$
0)
#617220000000
1"
1'
b0 +
b0 1
#617270000000
0"
0'
#617280000000
1#
1(
b101111101100100 +
b101111101100100 1
#617330000000
0#
0(
#617340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#617390000000
0$
0)
#617400000000
1"
1'
b0 +
b0 1
#617450000000
0"
0'
#617460000000
1#
1(
b101111101100100 +
b101111101100100 1
#617510000000
0#
0(
#617520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#617570000000
0$
0)
#617580000000
1"
1'
b0 +
b0 1
#617630000000
0"
0'
#617640000000
1#
1(
b101111101100100 +
b101111101100100 1
#617690000000
0#
0(
#617700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#617750000000
0$
0)
#617760000000
1"
1'
b0 +
b0 1
#617810000000
0"
0'
#617820000000
1#
1(
b101111101100100 +
b101111101100100 1
#617870000000
0#
0(
#617880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#617930000000
0$
0)
#617940000000
1"
1'
b0 +
b0 1
#617990000000
0"
0'
#618000000000
1#
1(
b101111101100100 +
b101111101100100 1
#618050000000
0#
0(
#618060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#618110000000
0$
0)
#618120000000
1"
1'
b0 +
b0 1
#618170000000
0"
0'
#618180000000
1#
1(
b101111101100100 +
b101111101100100 1
#618230000000
0#
0(
#618240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#618290000000
0$
0)
#618300000000
1"
1'
b0 +
b0 1
#618350000000
0"
0'
#618360000000
1#
1(
b101111101100100 +
b101111101100100 1
#618410000000
0#
0(
#618420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#618470000000
0$
0)
#618480000000
1"
1'
b0 +
b0 1
#618530000000
0"
0'
#618540000000
1#
1(
b101111101100100 +
b101111101100100 1
#618590000000
0#
0(
#618600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#618650000000
0$
0)
#618660000000
1"
1'
b0 +
b0 1
#618710000000
0"
0'
#618720000000
1#
1(
b101111101100100 +
b101111101100100 1
#618770000000
0#
0(
#618780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#618830000000
0$
0)
#618840000000
1"
1'
b0 +
b0 1
#618890000000
0"
0'
#618900000000
1#
1(
b101111101100100 +
b101111101100100 1
#618950000000
0#
0(
#618960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#619010000000
0$
0)
#619020000000
1"
1'
b0 +
b0 1
#619070000000
0"
0'
#619080000000
1#
1(
b101111101100100 +
b101111101100100 1
#619130000000
0#
0(
#619140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#619190000000
0$
0)
#619200000000
1"
1'
b0 +
b0 1
#619250000000
0"
0'
#619260000000
1#
1(
b101111101100100 +
b101111101100100 1
#619310000000
0#
0(
#619320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#619370000000
0$
0)
#619380000000
1"
1'
b0 +
b0 1
#619430000000
0"
0'
#619440000000
1#
1(
b101111101100100 +
b101111101100100 1
#619490000000
0#
0(
#619500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#619550000000
0$
0)
#619560000000
1"
1'
b0 +
b0 1
#619610000000
0"
0'
#619620000000
1#
1(
b101111101100100 +
b101111101100100 1
#619670000000
0#
0(
#619680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#619730000000
0$
0)
#619740000000
1"
1'
b0 +
b0 1
#619790000000
0"
0'
#619800000000
1#
1(
b101111101100100 +
b101111101100100 1
#619850000000
0#
0(
#619860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#619910000000
0$
0)
#619920000000
1"
1'
b0 +
b0 1
#619970000000
0"
0'
#619980000000
1#
1(
b101111101100100 +
b101111101100100 1
#620030000000
0#
0(
#620040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#620090000000
0$
0)
#620100000000
1"
1'
b0 +
b0 1
#620150000000
0"
0'
#620160000000
1#
1(
b101111101100100 +
b101111101100100 1
#620210000000
0#
0(
#620220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#620270000000
0$
0)
#620280000000
1"
1'
b0 +
b0 1
#620330000000
0"
0'
#620340000000
1#
1(
b101111101100100 +
b101111101100100 1
#620390000000
0#
0(
#620400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#620450000000
0$
0)
#620460000000
1"
1'
b0 +
b0 1
#620510000000
0"
0'
#620520000000
1#
1(
b101111101100100 +
b101111101100100 1
#620570000000
0#
0(
#620580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#620630000000
0$
0)
#620640000000
1"
1'
b0 +
b0 1
#620690000000
0"
0'
#620700000000
1#
1(
b101111101100100 +
b101111101100100 1
#620750000000
0#
0(
#620760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#620810000000
0$
0)
#620820000000
1"
1'
b0 +
b0 1
#620870000000
0"
0'
#620880000000
1#
1(
b101111101100100 +
b101111101100100 1
#620930000000
0#
0(
#620940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#620990000000
0$
0)
#621000000000
1"
1'
b0 +
b0 1
#621050000000
0"
0'
#621060000000
1#
1(
b101111101100100 +
b101111101100100 1
#621110000000
0#
0(
#621120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#621170000000
0$
0)
#621180000000
1"
1'
b0 +
b0 1
#621230000000
0"
0'
#621240000000
1#
1(
b101111101100100 +
b101111101100100 1
#621290000000
0#
0(
#621300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#621350000000
0$
0)
#621360000000
1"
1'
b0 +
b0 1
#621410000000
0"
0'
#621420000000
1#
1(
b101111101100100 +
b101111101100100 1
#621470000000
0#
0(
#621480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#621530000000
0$
0)
#621540000000
1"
1'
b0 +
b0 1
#621590000000
0"
0'
#621600000000
1#
1(
b101111101100100 +
b101111101100100 1
#621650000000
0#
0(
#621660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#621710000000
0$
0)
#621720000000
1"
1'
b0 +
b0 1
#621770000000
0"
0'
#621780000000
1#
1(
b101111101100100 +
b101111101100100 1
#621830000000
0#
0(
#621840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#621890000000
0$
0)
#621900000000
1"
1'
b0 +
b0 1
#621950000000
0"
0'
#621960000000
1#
1(
b101111101100100 +
b101111101100100 1
#622010000000
0#
0(
#622020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#622070000000
0$
0)
#622080000000
1"
1'
b0 +
b0 1
#622130000000
0"
0'
#622140000000
1#
1(
b101111101100100 +
b101111101100100 1
#622190000000
0#
0(
#622200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#622250000000
0$
0)
#622260000000
1"
1'
b0 +
b0 1
#622310000000
0"
0'
#622320000000
1#
1(
b101111101100100 +
b101111101100100 1
#622370000000
0#
0(
#622380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#622430000000
0$
0)
#622440000000
1"
1'
b0 +
b0 1
#622490000000
0"
0'
#622500000000
1#
1(
b101111101100100 +
b101111101100100 1
#622550000000
0#
0(
#622560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#622610000000
0$
0)
#622620000000
1"
1'
b0 +
b0 1
#622670000000
0"
0'
#622680000000
1#
1(
b101111101100100 +
b101111101100100 1
#622730000000
0#
0(
#622740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#622790000000
0$
0)
#622800000000
1"
1'
b0 +
b0 1
#622850000000
0"
0'
#622860000000
1#
1(
b101111101100100 +
b101111101100100 1
#622910000000
0#
0(
#622920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#622970000000
0$
0)
#622980000000
1"
1'
b0 +
b0 1
#623030000000
0"
0'
#623040000000
1#
1(
b101111101100100 +
b101111101100100 1
#623090000000
0#
0(
#623100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#623150000000
0$
0)
#623160000000
1"
1'
b0 +
b0 1
#623210000000
0"
0'
#623220000000
1#
1(
b101111101100100 +
b101111101100100 1
#623270000000
0#
0(
#623280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#623330000000
0$
0)
#623340000000
1"
1'
b0 +
b0 1
#623390000000
0"
0'
#623400000000
1#
1(
b101111101100100 +
b101111101100100 1
#623450000000
0#
0(
#623460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#623510000000
0$
0)
#623520000000
1"
1'
b0 +
b0 1
#623570000000
0"
0'
#623580000000
1#
1(
b101111101100100 +
b101111101100100 1
#623630000000
0#
0(
#623640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#623690000000
0$
0)
#623700000000
1"
1'
b0 +
b0 1
#623750000000
0"
0'
#623760000000
1#
1(
b101111101100100 +
b101111101100100 1
#623810000000
0#
0(
#623820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#623870000000
0$
0)
#623880000000
1"
1'
b0 +
b0 1
#623930000000
0"
0'
#623940000000
1#
1(
b101111101100100 +
b101111101100100 1
#623990000000
0#
0(
#624000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#624050000000
0$
0)
#624060000000
1"
1'
b0 +
b0 1
#624110000000
0"
0'
#624120000000
1#
1(
b101111101100100 +
b101111101100100 1
#624170000000
0#
0(
#624180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#624230000000
0$
0)
#624240000000
1"
1'
b0 +
b0 1
#624290000000
0"
0'
#624300000000
1#
1(
b101111101100100 +
b101111101100100 1
#624350000000
0#
0(
#624360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#624410000000
0$
0)
#624420000000
1"
1'
b0 +
b0 1
#624470000000
0"
0'
#624480000000
1#
1(
b101111101100100 +
b101111101100100 1
#624530000000
0#
0(
#624540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#624590000000
0$
0)
#624600000000
1"
1'
b0 +
b0 1
#624650000000
0"
0'
#624660000000
1#
1(
b101111101100100 +
b101111101100100 1
#624710000000
0#
0(
#624720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#624770000000
0$
0)
#624780000000
1"
1'
b0 +
b0 1
#624830000000
0"
0'
#624840000000
1#
1(
b101111101100100 +
b101111101100100 1
#624890000000
0#
0(
#624900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#624950000000
0$
0)
#624960000000
1"
1'
b0 +
b0 1
#625010000000
0"
0'
#625020000000
1#
1(
b101111101100100 +
b101111101100100 1
#625070000000
0#
0(
#625080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#625130000000
0$
0)
#625140000000
1"
1'
b0 +
b0 1
#625190000000
0"
0'
#625200000000
1#
1(
b101111101100100 +
b101111101100100 1
#625250000000
0#
0(
#625260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#625310000000
0$
0)
#625320000000
1"
1'
b0 +
b0 1
#625370000000
0"
0'
#625380000000
1#
1(
b101111101100100 +
b101111101100100 1
#625430000000
0#
0(
#625440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#625490000000
0$
0)
#625500000000
1"
1'
b0 +
b0 1
#625550000000
0"
0'
#625560000000
1#
1(
b101111101100100 +
b101111101100100 1
#625610000000
0#
0(
#625620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#625670000000
0$
0)
#625680000000
1"
1'
b0 +
b0 1
#625730000000
0"
0'
#625740000000
1#
1(
b101111101100100 +
b101111101100100 1
#625790000000
0#
0(
#625800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#625850000000
0$
0)
#625860000000
1"
1'
b0 +
b0 1
#625910000000
0"
0'
#625920000000
1#
1(
b101111101100100 +
b101111101100100 1
#625970000000
0#
0(
#625980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#626030000000
0$
0)
#626040000000
1"
1'
b0 +
b0 1
#626090000000
0"
0'
#626100000000
1#
1(
b101111101100100 +
b101111101100100 1
#626150000000
0#
0(
#626160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#626210000000
0$
0)
#626220000000
1"
1'
b0 +
b0 1
#626270000000
0"
0'
#626280000000
1#
1(
b101111101100100 +
b101111101100100 1
#626330000000
0#
0(
#626340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#626390000000
0$
0)
#626400000000
1"
1'
b0 +
b0 1
#626450000000
0"
0'
#626460000000
1#
1(
b101111101100100 +
b101111101100100 1
#626510000000
0#
0(
#626520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#626570000000
0$
0)
#626580000000
1"
1'
b0 +
b0 1
#626630000000
0"
0'
#626640000000
1#
1(
b101111101100100 +
b101111101100100 1
#626690000000
0#
0(
#626700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#626750000000
0$
0)
#626760000000
1"
1'
b0 +
b0 1
#626810000000
0"
0'
#626820000000
1#
1(
b101111101100100 +
b101111101100100 1
#626870000000
0#
0(
#626880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#626930000000
0$
0)
#626940000000
1"
1'
b0 +
b0 1
#626990000000
0"
0'
#627000000000
1#
1(
b101111101100100 +
b101111101100100 1
#627050000000
0#
0(
#627060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#627110000000
0$
0)
#627120000000
1"
1'
b0 +
b0 1
#627170000000
0"
0'
#627180000000
1#
1(
b101111101100100 +
b101111101100100 1
#627230000000
0#
0(
#627240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#627290000000
0$
0)
#627300000000
1"
1'
b0 +
b0 1
#627350000000
0"
0'
#627360000000
1#
1(
b101111101100100 +
b101111101100100 1
#627410000000
0#
0(
#627420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#627470000000
0$
0)
#627480000000
1"
1'
b0 +
b0 1
#627530000000
0"
0'
#627540000000
1#
1(
b101111101100100 +
b101111101100100 1
#627590000000
0#
0(
#627600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#627650000000
0$
0)
#627660000000
1"
1'
b0 +
b0 1
#627710000000
0"
0'
#627720000000
1#
1(
b101111101100100 +
b101111101100100 1
#627770000000
0#
0(
#627780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#627830000000
0$
0)
#627840000000
1"
1'
b0 +
b0 1
#627890000000
0"
0'
#627900000000
1#
1(
b101111101100100 +
b101111101100100 1
#627950000000
0#
0(
#627960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#628010000000
0$
0)
#628020000000
1"
1'
b0 +
b0 1
#628070000000
0"
0'
#628080000000
1#
1(
b101111101100100 +
b101111101100100 1
#628130000000
0#
0(
#628140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#628190000000
0$
0)
#628200000000
1"
1'
b0 +
b0 1
#628250000000
0"
0'
#628260000000
1#
1(
b101111101100100 +
b101111101100100 1
#628310000000
0#
0(
#628320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#628370000000
0$
0)
#628380000000
1"
1'
b0 +
b0 1
#628430000000
0"
0'
#628440000000
1#
1(
b101111101100100 +
b101111101100100 1
#628490000000
0#
0(
#628500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#628550000000
0$
0)
#628560000000
1"
1'
b0 +
b0 1
#628610000000
0"
0'
#628620000000
1#
1(
b101111101100100 +
b101111101100100 1
#628670000000
0#
0(
#628680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#628730000000
0$
0)
#628740000000
1"
1'
b0 +
b0 1
#628790000000
0"
0'
#628800000000
1#
1(
b101111101100100 +
b101111101100100 1
#628850000000
0#
0(
#628860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#628910000000
0$
0)
#628920000000
1"
1'
b0 +
b0 1
#628970000000
0"
0'
#628980000000
1#
1(
b101111101100100 +
b101111101100100 1
#629030000000
0#
0(
#629040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#629090000000
0$
0)
#629100000000
1"
1'
b0 +
b0 1
#629150000000
0"
0'
#629160000000
1#
1(
b101111101100100 +
b101111101100100 1
#629210000000
0#
0(
#629220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#629270000000
0$
0)
#629280000000
1"
1'
b0 +
b0 1
#629330000000
0"
0'
#629340000000
1#
1(
b101111101100100 +
b101111101100100 1
#629390000000
0#
0(
#629400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#629450000000
0$
0)
#629460000000
1"
1'
b0 +
b0 1
#629510000000
0"
0'
#629520000000
1#
1(
b101111101100100 +
b101111101100100 1
#629570000000
0#
0(
#629580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#629630000000
0$
0)
#629640000000
1"
1'
b0 +
b0 1
#629690000000
0"
0'
#629700000000
1#
1(
b101111101100100 +
b101111101100100 1
#629750000000
0#
0(
#629760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#629810000000
0$
0)
#629820000000
1"
1'
b0 +
b0 1
#629870000000
0"
0'
#629880000000
1#
1(
b101111101100100 +
b101111101100100 1
#629930000000
0#
0(
#629940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#629990000000
0$
0)
#630000000000
1"
1'
b0 +
b0 1
#630050000000
0"
0'
#630060000000
1#
1(
b101111101100100 +
b101111101100100 1
#630110000000
0#
0(
#630120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#630170000000
0$
0)
#630180000000
1"
1'
b0 +
b0 1
#630230000000
0"
0'
#630240000000
1#
1(
b101111101100100 +
b101111101100100 1
#630290000000
0#
0(
#630300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#630350000000
0$
0)
#630360000000
1"
1'
b0 +
b0 1
#630410000000
0"
0'
#630420000000
1#
1(
b101111101100100 +
b101111101100100 1
#630470000000
0#
0(
#630480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#630530000000
0$
0)
#630540000000
1"
1'
b0 +
b0 1
#630590000000
0"
0'
#630600000000
1#
1(
b101111101100100 +
b101111101100100 1
#630650000000
0#
0(
#630660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#630710000000
0$
0)
#630720000000
1"
1'
b0 +
b0 1
#630770000000
0"
0'
#630780000000
1#
1(
b101111101100100 +
b101111101100100 1
#630830000000
0#
0(
#630840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#630890000000
0$
0)
#630900000000
1"
1'
b0 +
b0 1
#630950000000
0"
0'
#630960000000
1#
1(
b101111101100100 +
b101111101100100 1
#631010000000
0#
0(
#631020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#631070000000
0$
0)
#631080000000
1"
1'
b0 +
b0 1
#631130000000
0"
0'
#631140000000
1#
1(
b101111101100100 +
b101111101100100 1
#631190000000
0#
0(
#631200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#631250000000
0$
0)
#631260000000
1"
1'
b0 +
b0 1
#631310000000
0"
0'
#631320000000
1#
1(
b101111101100100 +
b101111101100100 1
#631370000000
0#
0(
#631380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#631430000000
0$
0)
#631440000000
1"
1'
b0 +
b0 1
#631490000000
0"
0'
#631500000000
1#
1(
b101111101100100 +
b101111101100100 1
#631550000000
0#
0(
#631560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#631610000000
0$
0)
#631620000000
1"
1'
b0 +
b0 1
#631670000000
0"
0'
#631680000000
1#
1(
b101111101100100 +
b101111101100100 1
#631730000000
0#
0(
#631740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#631790000000
0$
0)
#631800000000
1"
1'
b0 +
b0 1
#631850000000
0"
0'
#631860000000
1#
1(
b101111101100100 +
b101111101100100 1
#631910000000
0#
0(
#631920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#631970000000
0$
0)
#631980000000
1"
1'
b0 +
b0 1
#632030000000
0"
0'
#632040000000
1#
1(
b101111101100100 +
b101111101100100 1
#632090000000
0#
0(
#632100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#632150000000
0$
0)
#632160000000
1"
1'
b0 +
b0 1
#632210000000
0"
0'
#632220000000
1#
1(
b101111101100100 +
b101111101100100 1
#632270000000
0#
0(
#632280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#632330000000
0$
0)
#632340000000
1"
1'
b0 +
b0 1
#632390000000
0"
0'
#632400000000
1#
1(
b101111101100100 +
b101111101100100 1
#632450000000
0#
0(
#632460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#632510000000
0$
0)
#632520000000
1"
1'
b0 +
b0 1
#632570000000
0"
0'
#632580000000
1#
1(
b101111101100100 +
b101111101100100 1
#632630000000
0#
0(
#632640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#632690000000
0$
0)
#632700000000
1"
1'
b0 +
b0 1
#632750000000
0"
0'
#632760000000
1#
1(
b101111101100100 +
b101111101100100 1
#632810000000
0#
0(
#632820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#632870000000
0$
0)
#632880000000
1"
1'
b0 +
b0 1
#632930000000
0"
0'
#632940000000
1#
1(
b101111101100100 +
b101111101100100 1
#632990000000
0#
0(
#633000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#633050000000
0$
0)
#633060000000
1"
1'
b0 +
b0 1
#633110000000
0"
0'
#633120000000
1#
1(
b101111101100100 +
b101111101100100 1
#633170000000
0#
0(
#633180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#633230000000
0$
0)
#633240000000
1"
1'
b0 +
b0 1
#633290000000
0"
0'
#633300000000
1#
1(
b101111101100100 +
b101111101100100 1
#633350000000
0#
0(
#633360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#633410000000
0$
0)
#633420000000
1"
1'
b0 +
b0 1
#633470000000
0"
0'
#633480000000
1#
1(
b101111101100100 +
b101111101100100 1
#633530000000
0#
0(
#633540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#633590000000
0$
0)
#633600000000
1"
1'
b0 +
b0 1
#633650000000
0"
0'
#633660000000
1#
1(
b101111101100100 +
b101111101100100 1
#633710000000
0#
0(
#633720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#633770000000
0$
0)
#633780000000
1"
1'
b0 +
b0 1
#633830000000
0"
0'
#633840000000
1#
1(
b101111101100100 +
b101111101100100 1
#633890000000
0#
0(
#633900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#633950000000
0$
0)
#633960000000
1"
1'
b0 +
b0 1
#634010000000
0"
0'
#634020000000
1#
1(
b101111101100100 +
b101111101100100 1
#634070000000
0#
0(
#634080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#634130000000
0$
0)
#634140000000
1"
1'
b0 +
b0 1
#634190000000
0"
0'
#634200000000
1#
1(
b101111101100100 +
b101111101100100 1
#634250000000
0#
0(
#634260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#634310000000
0$
0)
#634320000000
1"
1'
b0 +
b0 1
#634370000000
0"
0'
#634380000000
1#
1(
b101111101100100 +
b101111101100100 1
#634430000000
0#
0(
#634440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#634490000000
0$
0)
#634500000000
1"
1'
b0 +
b0 1
#634550000000
0"
0'
#634560000000
1#
1(
b101111101100100 +
b101111101100100 1
#634610000000
0#
0(
#634620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#634670000000
0$
0)
#634680000000
1"
1'
b0 +
b0 1
#634730000000
0"
0'
#634740000000
1#
1(
b101111101100100 +
b101111101100100 1
#634790000000
0#
0(
#634800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#634850000000
0$
0)
#634860000000
1"
1'
b0 +
b0 1
#634910000000
0"
0'
#634920000000
1#
1(
b101111101100100 +
b101111101100100 1
#634970000000
0#
0(
#634980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#635030000000
0$
0)
#635040000000
1"
1'
b0 +
b0 1
#635090000000
0"
0'
#635100000000
1#
1(
b101111101100100 +
b101111101100100 1
#635150000000
0#
0(
#635160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#635210000000
0$
0)
#635220000000
1"
1'
b0 +
b0 1
#635270000000
0"
0'
#635280000000
1#
1(
b101111101100100 +
b101111101100100 1
#635330000000
0#
0(
#635340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#635390000000
0$
0)
#635400000000
1"
1'
b0 +
b0 1
#635450000000
0"
0'
#635460000000
1#
1(
b101111101100100 +
b101111101100100 1
#635510000000
0#
0(
#635520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#635570000000
0$
0)
#635580000000
1"
1'
b0 +
b0 1
#635630000000
0"
0'
#635640000000
1#
1(
b101111101100100 +
b101111101100100 1
#635690000000
0#
0(
#635700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#635750000000
0$
0)
#635760000000
1"
1'
b0 +
b0 1
#635810000000
0"
0'
#635820000000
1#
1(
b101111101100100 +
b101111101100100 1
#635870000000
0#
0(
#635880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#635930000000
0$
0)
#635940000000
1"
1'
b0 +
b0 1
#635990000000
0"
0'
#636000000000
1#
1(
b101111101100100 +
b101111101100100 1
#636050000000
0#
0(
#636060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#636110000000
0$
0)
#636120000000
1"
1'
b0 +
b0 1
#636170000000
0"
0'
#636180000000
1#
1(
b101111101100100 +
b101111101100100 1
#636230000000
0#
0(
#636240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#636290000000
0$
0)
#636300000000
1"
1'
b0 +
b0 1
#636350000000
0"
0'
#636360000000
1#
1(
b101111101100100 +
b101111101100100 1
#636410000000
0#
0(
#636420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#636470000000
0$
0)
#636480000000
1"
1'
b0 +
b0 1
#636530000000
0"
0'
#636540000000
1#
1(
b101111101100100 +
b101111101100100 1
#636590000000
0#
0(
#636600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#636650000000
0$
0)
#636660000000
1"
1'
b0 +
b0 1
#636710000000
0"
0'
#636720000000
1#
1(
b101111101100100 +
b101111101100100 1
#636770000000
0#
0(
#636780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#636830000000
0$
0)
#636840000000
1"
1'
b0 +
b0 1
#636890000000
0"
0'
#636900000000
1#
1(
b101111101100100 +
b101111101100100 1
#636950000000
0#
0(
#636960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#637010000000
0$
0)
#637020000000
1"
1'
b0 +
b0 1
#637070000000
0"
0'
#637080000000
1#
1(
b101111101100100 +
b101111101100100 1
#637130000000
0#
0(
#637140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#637190000000
0$
0)
#637200000000
1"
1'
b0 +
b0 1
#637250000000
0"
0'
#637260000000
1#
1(
b101111101100100 +
b101111101100100 1
#637310000000
0#
0(
#637320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#637370000000
0$
0)
#637380000000
1"
1'
b0 +
b0 1
#637430000000
0"
0'
#637440000000
1#
1(
b101111101100100 +
b101111101100100 1
#637490000000
0#
0(
#637500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#637550000000
0$
0)
#637560000000
1"
1'
b0 +
b0 1
#637610000000
0"
0'
#637620000000
1#
1(
b101111101100100 +
b101111101100100 1
#637670000000
0#
0(
#637680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#637730000000
0$
0)
#637740000000
1"
1'
b0 +
b0 1
#637790000000
0"
0'
#637800000000
1#
1(
b101111101100100 +
b101111101100100 1
#637850000000
0#
0(
#637860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#637910000000
0$
0)
#637920000000
1"
1'
b0 +
b0 1
#637970000000
0"
0'
#637980000000
1#
1(
b101111101100100 +
b101111101100100 1
#638030000000
0#
0(
#638040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#638090000000
0$
0)
#638100000000
1"
1'
b0 +
b0 1
#638150000000
0"
0'
#638160000000
1#
1(
b101111101100100 +
b101111101100100 1
#638210000000
0#
0(
#638220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#638270000000
0$
0)
#638280000000
1"
1'
b0 +
b0 1
#638330000000
0"
0'
#638340000000
1#
1(
b101111101100100 +
b101111101100100 1
#638390000000
0#
0(
#638400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#638450000000
0$
0)
#638460000000
1"
1'
b0 +
b0 1
#638510000000
0"
0'
#638520000000
1#
1(
b101111101100100 +
b101111101100100 1
#638570000000
0#
0(
#638580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#638630000000
0$
0)
#638640000000
1"
1'
b0 +
b0 1
#638690000000
0"
0'
#638700000000
1#
1(
b101111101100100 +
b101111101100100 1
#638750000000
0#
0(
#638760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#638810000000
0$
0)
#638820000000
1"
1'
b0 +
b0 1
#638870000000
0"
0'
#638880000000
1#
1(
b101111101100100 +
b101111101100100 1
#638930000000
0#
0(
#638940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#638990000000
0$
0)
#639000000000
1"
1'
b0 +
b0 1
#639050000000
0"
0'
#639060000000
1#
1(
b101111101100100 +
b101111101100100 1
#639110000000
0#
0(
#639120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#639170000000
0$
0)
#639180000000
1"
1'
b0 +
b0 1
#639230000000
0"
0'
#639240000000
1#
1(
b101111101100100 +
b101111101100100 1
#639290000000
0#
0(
#639300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#639350000000
0$
0)
#639360000000
1"
1'
b0 +
b0 1
#639410000000
0"
0'
#639420000000
1#
1(
b101111101100100 +
b101111101100100 1
#639470000000
0#
0(
#639480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#639530000000
0$
0)
#639540000000
1"
1'
b0 +
b0 1
#639590000000
0"
0'
#639600000000
1#
1(
b101111101100100 +
b101111101100100 1
#639650000000
0#
0(
#639660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#639710000000
0$
0)
#639720000000
1"
1'
b0 +
b0 1
#639770000000
0"
0'
#639780000000
1#
1(
b101111101100100 +
b101111101100100 1
#639830000000
0#
0(
#639840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#639890000000
0$
0)
#639900000000
1"
1'
b0 +
b0 1
#639950000000
0"
0'
#639960000000
1#
1(
b101111101100100 +
b101111101100100 1
#640010000000
0#
0(
#640020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#640070000000
0$
0)
#640080000000
1"
1'
b0 +
b0 1
#640130000000
0"
0'
#640140000000
1#
1(
b101111101100100 +
b101111101100100 1
#640190000000
0#
0(
#640200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#640250000000
0$
0)
#640260000000
1"
1'
b0 +
b0 1
#640310000000
0"
0'
#640320000000
1#
1(
b101111101100100 +
b101111101100100 1
#640370000000
0#
0(
#640380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#640430000000
0$
0)
#640440000000
1"
1'
b0 +
b0 1
#640490000000
0"
0'
#640500000000
1#
1(
b101111101100100 +
b101111101100100 1
#640550000000
0#
0(
#640560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#640610000000
0$
0)
#640620000000
1"
1'
b0 +
b0 1
#640670000000
0"
0'
#640680000000
1#
1(
b101111101100100 +
b101111101100100 1
#640730000000
0#
0(
#640740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#640790000000
0$
0)
#640800000000
1"
1'
b0 +
b0 1
#640850000000
0"
0'
#640860000000
1#
1(
b101111101100100 +
b101111101100100 1
#640910000000
0#
0(
#640920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#640970000000
0$
0)
#640980000000
1"
1'
b0 +
b0 1
#641030000000
0"
0'
#641040000000
1#
1(
b101111101100100 +
b101111101100100 1
#641090000000
0#
0(
#641100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#641150000000
0$
0)
#641160000000
1"
1'
b0 +
b0 1
#641210000000
0"
0'
#641220000000
1#
1(
b101111101100100 +
b101111101100100 1
#641270000000
0#
0(
#641280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#641330000000
0$
0)
#641340000000
1"
1'
b0 +
b0 1
#641390000000
0"
0'
#641400000000
1#
1(
b101111101100100 +
b101111101100100 1
#641450000000
0#
0(
#641460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#641510000000
0$
0)
#641520000000
1"
1'
b0 +
b0 1
#641570000000
0"
0'
#641580000000
1#
1(
b101111101100100 +
b101111101100100 1
#641630000000
0#
0(
#641640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#641690000000
0$
0)
#641700000000
1"
1'
b0 +
b0 1
#641750000000
0"
0'
#641760000000
1#
1(
b101111101100100 +
b101111101100100 1
#641810000000
0#
0(
#641820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#641870000000
0$
0)
#641880000000
1"
1'
b0 +
b0 1
#641930000000
0"
0'
#641940000000
1#
1(
b101111101100100 +
b101111101100100 1
#641990000000
0#
0(
#642000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#642050000000
0$
0)
#642060000000
1"
1'
b0 +
b0 1
#642110000000
0"
0'
#642120000000
1#
1(
b101111101100100 +
b101111101100100 1
#642170000000
0#
0(
#642180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#642230000000
0$
0)
#642240000000
1"
1'
b0 +
b0 1
#642290000000
0"
0'
#642300000000
1#
1(
b101111101100100 +
b101111101100100 1
#642350000000
0#
0(
#642360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#642410000000
0$
0)
#642420000000
1"
1'
b0 +
b0 1
#642470000000
0"
0'
#642480000000
1#
1(
b101111101100100 +
b101111101100100 1
#642530000000
0#
0(
#642540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#642590000000
0$
0)
#642600000000
1"
1'
b0 +
b0 1
#642650000000
0"
0'
#642660000000
1#
1(
b101111101100100 +
b101111101100100 1
#642710000000
0#
0(
#642720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#642770000000
0$
0)
#642780000000
1"
1'
b0 +
b0 1
#642830000000
0"
0'
#642840000000
1#
1(
b101111101100100 +
b101111101100100 1
#642890000000
0#
0(
#642900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#642950000000
0$
0)
#642960000000
1"
1'
b0 +
b0 1
#643010000000
0"
0'
#643020000000
1#
1(
b101111101100100 +
b101111101100100 1
#643070000000
0#
0(
#643080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#643130000000
0$
0)
#643140000000
1"
1'
b0 +
b0 1
#643190000000
0"
0'
#643200000000
1#
1(
b101111101100100 +
b101111101100100 1
#643250000000
0#
0(
#643260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#643310000000
0$
0)
#643320000000
1"
1'
b0 +
b0 1
#643370000000
0"
0'
#643380000000
1#
1(
b101111101100100 +
b101111101100100 1
#643430000000
0#
0(
#643440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#643490000000
0$
0)
#643500000000
1"
1'
b0 +
b0 1
#643550000000
0"
0'
#643560000000
1#
1(
b101111101100100 +
b101111101100100 1
#643610000000
0#
0(
#643620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#643670000000
0$
0)
#643680000000
1"
1'
b0 +
b0 1
#643730000000
0"
0'
#643740000000
1#
1(
b101111101100100 +
b101111101100100 1
#643790000000
0#
0(
#643800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#643850000000
0$
0)
#643860000000
1"
1'
b0 +
b0 1
#643910000000
0"
0'
#643920000000
1#
1(
b101111101100100 +
b101111101100100 1
#643970000000
0#
0(
#643980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#644030000000
0$
0)
#644040000000
1"
1'
b0 +
b0 1
#644090000000
0"
0'
#644100000000
1#
1(
b101111101100100 +
b101111101100100 1
#644150000000
0#
0(
#644160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#644210000000
0$
0)
#644220000000
1"
1'
b0 +
b0 1
#644270000000
0"
0'
#644280000000
1#
1(
b101111101100100 +
b101111101100100 1
#644330000000
0#
0(
#644340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#644390000000
0$
0)
#644400000000
1"
1'
b0 +
b0 1
#644450000000
0"
0'
#644460000000
1#
1(
b101111101100100 +
b101111101100100 1
#644510000000
0#
0(
#644520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#644570000000
0$
0)
#644580000000
1"
1'
b0 +
b0 1
#644630000000
0"
0'
#644640000000
1#
1(
b101111101100100 +
b101111101100100 1
#644690000000
0#
0(
#644700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#644750000000
0$
0)
#644760000000
1"
1'
b0 +
b0 1
#644810000000
0"
0'
#644820000000
1#
1(
b101111101100100 +
b101111101100100 1
#644870000000
0#
0(
#644880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#644930000000
0$
0)
#644940000000
1"
1'
b0 +
b0 1
#644990000000
0"
0'
#645000000000
1#
1(
b101111101100100 +
b101111101100100 1
#645050000000
0#
0(
#645060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#645110000000
0$
0)
#645120000000
1"
1'
b0 +
b0 1
#645170000000
0"
0'
#645180000000
1#
1(
b101111101100100 +
b101111101100100 1
#645230000000
0#
0(
#645240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#645290000000
0$
0)
#645300000000
1"
1'
b0 +
b0 1
#645350000000
0"
0'
#645360000000
1#
1(
b101111101100100 +
b101111101100100 1
#645410000000
0#
0(
#645420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#645470000000
0$
0)
#645480000000
1"
1'
b0 +
b0 1
#645530000000
0"
0'
#645540000000
1#
1(
b101111101100100 +
b101111101100100 1
#645590000000
0#
0(
#645600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#645650000000
0$
0)
#645660000000
1"
1'
b0 +
b0 1
#645710000000
0"
0'
#645720000000
1#
1(
b101111101100100 +
b101111101100100 1
#645770000000
0#
0(
#645780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#645830000000
0$
0)
#645840000000
1"
1'
b0 +
b0 1
#645890000000
0"
0'
#645900000000
1#
1(
b101111101100100 +
b101111101100100 1
#645950000000
0#
0(
#645960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#646010000000
0$
0)
#646020000000
1"
1'
b0 +
b0 1
#646070000000
0"
0'
#646080000000
1#
1(
b101111101100100 +
b101111101100100 1
#646130000000
0#
0(
#646140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#646190000000
0$
0)
#646200000000
1"
1'
b0 +
b0 1
#646250000000
0"
0'
#646260000000
1#
1(
b101111101100100 +
b101111101100100 1
#646310000000
0#
0(
#646320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#646370000000
0$
0)
#646380000000
1"
1'
b0 +
b0 1
#646430000000
0"
0'
#646440000000
1#
1(
b101111101100100 +
b101111101100100 1
#646490000000
0#
0(
#646500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#646550000000
0$
0)
#646560000000
1"
1'
b0 +
b0 1
#646610000000
0"
0'
#646620000000
1#
1(
b101111101100100 +
b101111101100100 1
#646670000000
0#
0(
#646680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#646730000000
0$
0)
#646740000000
1"
1'
b0 +
b0 1
#646790000000
0"
0'
#646800000000
1#
1(
b101111101100100 +
b101111101100100 1
#646850000000
0#
0(
#646860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#646910000000
0$
0)
#646920000000
1"
1'
b0 +
b0 1
#646970000000
0"
0'
#646980000000
1#
1(
b101111101100100 +
b101111101100100 1
#647030000000
0#
0(
#647040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#647090000000
0$
0)
#647100000000
1"
1'
b0 +
b0 1
#647150000000
0"
0'
#647160000000
1#
1(
b101111101100100 +
b101111101100100 1
#647210000000
0#
0(
#647220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#647270000000
0$
0)
#647280000000
1"
1'
b0 +
b0 1
#647330000000
0"
0'
#647340000000
1#
1(
b101111101100100 +
b101111101100100 1
#647390000000
0#
0(
#647400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#647450000000
0$
0)
#647460000000
1"
1'
b0 +
b0 1
#647510000000
0"
0'
#647520000000
1#
1(
b101111101100100 +
b101111101100100 1
#647570000000
0#
0(
#647580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#647630000000
0$
0)
#647640000000
1"
1'
b0 +
b0 1
#647690000000
0"
0'
#647700000000
1#
1(
b101111101100100 +
b101111101100100 1
#647750000000
0#
0(
#647760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#647810000000
0$
0)
#647820000000
1"
1'
b0 +
b0 1
#647870000000
0"
0'
#647880000000
1#
1(
b101111101100100 +
b101111101100100 1
#647930000000
0#
0(
#647940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#647990000000
0$
0)
#648000000000
1"
1'
b0 +
b0 1
#648050000000
0"
0'
#648060000000
1#
1(
b101111101100100 +
b101111101100100 1
#648110000000
0#
0(
#648120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#648170000000
0$
0)
#648180000000
1"
1'
b0 +
b0 1
#648230000000
0"
0'
#648240000000
1#
1(
b101111101100100 +
b101111101100100 1
#648290000000
0#
0(
#648300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#648350000000
0$
0)
#648360000000
1"
1'
b0 +
b0 1
#648410000000
0"
0'
#648420000000
1#
1(
b101111101100100 +
b101111101100100 1
#648470000000
0#
0(
#648480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#648530000000
0$
0)
#648540000000
1"
1'
b0 +
b0 1
#648590000000
0"
0'
#648600000000
1#
1(
b101111101100100 +
b101111101100100 1
#648650000000
0#
0(
#648660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#648710000000
0$
0)
#648720000000
1"
1'
b0 +
b0 1
#648770000000
0"
0'
#648780000000
1#
1(
b101111101100100 +
b101111101100100 1
#648830000000
0#
0(
#648840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#648890000000
0$
0)
#648900000000
1"
1'
b0 +
b0 1
#648950000000
0"
0'
#648960000000
1#
1(
b101111101100100 +
b101111101100100 1
#649010000000
0#
0(
#649020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#649070000000
0$
0)
#649080000000
1"
1'
b0 +
b0 1
#649130000000
0"
0'
#649140000000
1#
1(
b101111101100100 +
b101111101100100 1
#649190000000
0#
0(
#649200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#649250000000
0$
0)
#649260000000
1"
1'
b0 +
b0 1
#649310000000
0"
0'
#649320000000
1#
1(
b101111101100100 +
b101111101100100 1
#649370000000
0#
0(
#649380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#649430000000
0$
0)
#649440000000
1"
1'
b0 +
b0 1
#649490000000
0"
0'
#649500000000
1#
1(
b101111101100100 +
b101111101100100 1
#649550000000
0#
0(
#649560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#649610000000
0$
0)
#649620000000
1"
1'
b0 +
b0 1
#649670000000
0"
0'
#649680000000
1#
1(
b101111101100100 +
b101111101100100 1
#649730000000
0#
0(
#649740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#649790000000
0$
0)
#649800000000
1"
1'
b0 +
b0 1
#649850000000
0"
0'
#649860000000
1#
1(
b101111101100100 +
b101111101100100 1
#649910000000
0#
0(
#649920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#649970000000
0$
0)
#649980000000
1"
1'
b0 +
b0 1
#650030000000
0"
0'
#650040000000
1#
1(
b101111101100100 +
b101111101100100 1
#650090000000
0#
0(
#650100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#650150000000
0$
0)
#650160000000
1"
1'
b0 +
b0 1
#650210000000
0"
0'
#650220000000
1#
1(
b101111101100100 +
b101111101100100 1
#650270000000
0#
0(
#650280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#650330000000
0$
0)
#650340000000
1"
1'
b0 +
b0 1
#650390000000
0"
0'
#650400000000
1#
1(
b101111101100100 +
b101111101100100 1
#650450000000
0#
0(
#650460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#650510000000
0$
0)
#650520000000
1"
1'
b0 +
b0 1
#650570000000
0"
0'
#650580000000
1#
1(
b101111101100100 +
b101111101100100 1
#650630000000
0#
0(
#650640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#650690000000
0$
0)
#650700000000
1"
1'
b0 +
b0 1
#650750000000
0"
0'
#650760000000
1#
1(
b101111101100100 +
b101111101100100 1
#650810000000
0#
0(
#650820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#650870000000
0$
0)
#650880000000
1"
1'
b0 +
b0 1
#650930000000
0"
0'
#650940000000
1#
1(
b101111101100100 +
b101111101100100 1
#650990000000
0#
0(
#651000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#651050000000
0$
0)
#651060000000
1"
1'
b0 +
b0 1
#651110000000
0"
0'
#651120000000
1#
1(
b101111101100100 +
b101111101100100 1
#651170000000
0#
0(
#651180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#651230000000
0$
0)
#651240000000
1"
1'
b0 +
b0 1
#651290000000
0"
0'
#651300000000
1#
1(
b101111101100100 +
b101111101100100 1
#651350000000
0#
0(
#651360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#651410000000
0$
0)
#651420000000
1"
1'
b0 +
b0 1
#651470000000
0"
0'
#651480000000
1#
1(
b101111101100100 +
b101111101100100 1
#651530000000
0#
0(
#651540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#651590000000
0$
0)
#651600000000
1"
1'
b0 +
b0 1
#651650000000
0"
0'
#651660000000
1#
1(
b101111101100100 +
b101111101100100 1
#651710000000
0#
0(
#651720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#651770000000
0$
0)
#651780000000
1"
1'
b0 +
b0 1
#651830000000
0"
0'
#651840000000
1#
1(
b101111101100100 +
b101111101100100 1
#651890000000
0#
0(
#651900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#651950000000
0$
0)
#651960000000
1"
1'
b0 +
b0 1
#652010000000
0"
0'
#652020000000
1#
1(
b101111101100100 +
b101111101100100 1
#652070000000
0#
0(
#652080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#652130000000
0$
0)
#652140000000
1"
1'
b0 +
b0 1
#652190000000
0"
0'
#652200000000
1#
1(
b101111101100100 +
b101111101100100 1
#652250000000
0#
0(
#652260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#652310000000
0$
0)
#652320000000
1"
1'
b0 +
b0 1
#652370000000
0"
0'
#652380000000
1#
1(
b101111101100100 +
b101111101100100 1
#652430000000
0#
0(
#652440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#652490000000
0$
0)
#652500000000
1"
1'
b0 +
b0 1
#652550000000
0"
0'
#652560000000
1#
1(
b101111101100100 +
b101111101100100 1
#652610000000
0#
0(
#652620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#652670000000
0$
0)
#652680000000
1"
1'
b0 +
b0 1
#652730000000
0"
0'
#652740000000
1#
1(
b101111101100100 +
b101111101100100 1
#652790000000
0#
0(
#652800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#652850000000
0$
0)
#652860000000
1"
1'
b0 +
b0 1
#652910000000
0"
0'
#652920000000
1#
1(
b101111101100100 +
b101111101100100 1
#652970000000
0#
0(
#652980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#653030000000
0$
0)
#653040000000
1"
1'
b0 +
b0 1
#653090000000
0"
0'
#653100000000
1#
1(
b101111101100100 +
b101111101100100 1
#653150000000
0#
0(
#653160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#653210000000
0$
0)
#653220000000
1"
1'
b0 +
b0 1
#653270000000
0"
0'
#653280000000
1#
1(
b101111101100100 +
b101111101100100 1
#653330000000
0#
0(
#653340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#653390000000
0$
0)
#653400000000
1"
1'
b0 +
b0 1
#653450000000
0"
0'
#653460000000
1#
1(
b101111101100100 +
b101111101100100 1
#653510000000
0#
0(
#653520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#653570000000
0$
0)
#653580000000
1"
1'
b0 +
b0 1
#653630000000
0"
0'
#653640000000
1#
1(
b101111101100100 +
b101111101100100 1
#653690000000
0#
0(
#653700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#653750000000
0$
0)
#653760000000
1"
1'
b0 +
b0 1
#653810000000
0"
0'
#653820000000
1#
1(
b101111101100100 +
b101111101100100 1
#653870000000
0#
0(
#653880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#653930000000
0$
0)
#653940000000
1"
1'
b0 +
b0 1
#653990000000
0"
0'
#654000000000
1#
1(
b101111101100100 +
b101111101100100 1
#654050000000
0#
0(
#654060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#654110000000
0$
0)
#654120000000
1"
1'
b0 +
b0 1
#654170000000
0"
0'
#654180000000
1#
1(
b101111101100100 +
b101111101100100 1
#654230000000
0#
0(
#654240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#654290000000
0$
0)
#654300000000
1"
1'
b0 +
b0 1
#654350000000
0"
0'
#654360000000
1#
1(
b101111101100100 +
b101111101100100 1
#654410000000
0#
0(
#654420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#654470000000
0$
0)
#654480000000
1"
1'
b0 +
b0 1
#654530000000
0"
0'
#654540000000
1#
1(
b101111101100100 +
b101111101100100 1
#654590000000
0#
0(
#654600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#654650000000
0$
0)
#654660000000
1"
1'
b0 +
b0 1
#654710000000
0"
0'
#654720000000
1#
1(
b101111101100100 +
b101111101100100 1
#654770000000
0#
0(
#654780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#654830000000
0$
0)
#654840000000
1"
1'
b0 +
b0 1
#654890000000
0"
0'
#654900000000
1#
1(
b101111101100100 +
b101111101100100 1
#654950000000
0#
0(
#654960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#655010000000
0$
0)
#655020000000
1"
1'
b0 +
b0 1
#655070000000
0"
0'
#655080000000
1#
1(
b101111101100100 +
b101111101100100 1
#655130000000
0#
0(
#655140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#655190000000
0$
0)
#655200000000
1"
1'
b0 +
b0 1
#655250000000
0"
0'
#655260000000
1#
1(
b101111101100100 +
b101111101100100 1
#655310000000
0#
0(
#655320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#655370000000
0$
0)
#655380000000
1"
1'
b0 +
b0 1
#655430000000
0"
0'
#655440000000
1#
1(
b101111101100100 +
b101111101100100 1
#655490000000
0#
0(
#655500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#655550000000
0$
0)
#655560000000
1"
1'
b0 +
b0 1
#655610000000
0"
0'
#655620000000
1#
1(
b101111101100100 +
b101111101100100 1
#655670000000
0#
0(
#655680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#655730000000
0$
0)
#655740000000
1"
1'
b0 +
b0 1
#655790000000
0"
0'
#655800000000
1#
1(
b101111101100100 +
b101111101100100 1
#655850000000
0#
0(
#655860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#655910000000
0$
0)
#655920000000
1"
1'
b0 +
b0 1
#655970000000
0"
0'
#655980000000
1#
1(
b101111101100100 +
b101111101100100 1
#656030000000
0#
0(
#656040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#656090000000
0$
0)
#656100000000
1"
1'
b0 +
b0 1
#656150000000
0"
0'
#656160000000
1#
1(
b101111101100100 +
b101111101100100 1
#656210000000
0#
0(
#656220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#656270000000
0$
0)
#656280000000
1"
1'
b0 +
b0 1
#656330000000
0"
0'
#656340000000
1#
1(
b101111101100100 +
b101111101100100 1
#656390000000
0#
0(
#656400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#656450000000
0$
0)
#656460000000
1"
1'
b0 +
b0 1
#656510000000
0"
0'
#656520000000
1#
1(
b101111101100100 +
b101111101100100 1
#656570000000
0#
0(
#656580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#656630000000
0$
0)
#656640000000
1"
1'
b0 +
b0 1
#656690000000
0"
0'
#656700000000
1#
1(
b101111101100100 +
b101111101100100 1
#656750000000
0#
0(
#656760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#656810000000
0$
0)
#656820000000
1"
1'
b0 +
b0 1
#656870000000
0"
0'
#656880000000
1#
1(
b101111101100100 +
b101111101100100 1
#656930000000
0#
0(
#656940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#656990000000
0$
0)
#657000000000
1"
1'
b0 +
b0 1
#657050000000
0"
0'
#657060000000
1#
1(
b101111101100100 +
b101111101100100 1
#657110000000
0#
0(
#657120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#657170000000
0$
0)
#657180000000
1"
1'
b0 +
b0 1
#657230000000
0"
0'
#657240000000
1#
1(
b101111101100100 +
b101111101100100 1
#657290000000
0#
0(
#657300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#657350000000
0$
0)
#657360000000
1"
1'
b0 +
b0 1
#657410000000
0"
0'
#657420000000
1#
1(
b101111101100100 +
b101111101100100 1
#657470000000
0#
0(
#657480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#657530000000
0$
0)
#657540000000
1"
1'
b0 +
b0 1
#657590000000
0"
0'
#657600000000
1#
1(
b101111101100100 +
b101111101100100 1
#657650000000
0#
0(
#657660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#657710000000
0$
0)
#657720000000
1"
1'
b0 +
b0 1
#657770000000
0"
0'
#657780000000
1#
1(
b101111101100100 +
b101111101100100 1
#657830000000
0#
0(
#657840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#657890000000
0$
0)
#657900000000
1"
1'
b0 +
b0 1
#657950000000
0"
0'
#657960000000
1#
1(
b101111101100100 +
b101111101100100 1
#658010000000
0#
0(
#658020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#658070000000
0$
0)
#658080000000
1"
1'
b0 +
b0 1
#658130000000
0"
0'
#658140000000
1#
1(
b101111101100100 +
b101111101100100 1
#658190000000
0#
0(
#658200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#658250000000
0$
0)
#658260000000
1"
1'
b0 +
b0 1
#658310000000
0"
0'
#658320000000
1#
1(
b101111101100100 +
b101111101100100 1
#658370000000
0#
0(
#658380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#658430000000
0$
0)
#658440000000
1"
1'
b0 +
b0 1
#658490000000
0"
0'
#658500000000
1#
1(
b101111101100100 +
b101111101100100 1
#658550000000
0#
0(
#658560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#658610000000
0$
0)
#658620000000
1"
1'
b0 +
b0 1
#658670000000
0"
0'
#658680000000
1#
1(
b101111101100100 +
b101111101100100 1
#658730000000
0#
0(
#658740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#658790000000
0$
0)
#658800000000
1"
1'
b0 +
b0 1
#658850000000
0"
0'
#658860000000
1#
1(
b101111101100100 +
b101111101100100 1
#658910000000
0#
0(
#658920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#658970000000
0$
0)
#658980000000
1"
1'
b0 +
b0 1
#659030000000
0"
0'
#659040000000
1#
1(
b101111101100100 +
b101111101100100 1
#659090000000
0#
0(
#659100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#659150000000
0$
0)
#659160000000
1"
1'
b0 +
b0 1
#659210000000
0"
0'
#659220000000
1#
1(
b101111101100100 +
b101111101100100 1
#659270000000
0#
0(
#659280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#659330000000
0$
0)
#659340000000
1"
1'
b0 +
b0 1
#659390000000
0"
0'
#659400000000
1#
1(
b101111101100100 +
b101111101100100 1
#659450000000
0#
0(
#659460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#659510000000
0$
0)
#659520000000
1"
1'
b0 +
b0 1
#659570000000
0"
0'
#659580000000
1#
1(
b101111101100100 +
b101111101100100 1
#659630000000
0#
0(
#659640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#659690000000
0$
0)
#659700000000
1"
1'
b0 +
b0 1
#659750000000
0"
0'
#659760000000
1#
1(
b101111101100100 +
b101111101100100 1
#659810000000
0#
0(
#659820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#659870000000
0$
0)
#659880000000
1"
1'
b0 +
b0 1
#659930000000
0"
0'
#659940000000
1#
1(
b101111101100100 +
b101111101100100 1
#659990000000
0#
0(
#660000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#660050000000
0$
0)
#660060000000
1"
1'
b0 +
b0 1
#660110000000
0"
0'
#660120000000
1#
1(
b101111101100100 +
b101111101100100 1
#660170000000
0#
0(
#660180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#660230000000
0$
0)
#660240000000
1"
1'
b0 +
b0 1
#660290000000
0"
0'
#660300000000
1#
1(
b101111101100100 +
b101111101100100 1
#660350000000
0#
0(
#660360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#660410000000
0$
0)
#660420000000
1"
1'
b0 +
b0 1
#660470000000
0"
0'
#660480000000
1#
1(
b101111101100100 +
b101111101100100 1
#660530000000
0#
0(
#660540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#660590000000
0$
0)
#660600000000
1"
1'
b0 +
b0 1
#660650000000
0"
0'
#660660000000
1#
1(
b101111101100100 +
b101111101100100 1
#660710000000
0#
0(
#660720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#660770000000
0$
0)
#660780000000
1"
1'
b0 +
b0 1
#660830000000
0"
0'
#660840000000
1#
1(
b101111101100100 +
b101111101100100 1
#660890000000
0#
0(
#660900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#660950000000
0$
0)
#660960000000
1"
1'
b0 +
b0 1
#661010000000
0"
0'
#661020000000
1#
1(
b101111101100100 +
b101111101100100 1
#661070000000
0#
0(
#661080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#661130000000
0$
0)
#661140000000
1"
1'
b0 +
b0 1
#661190000000
0"
0'
#661200000000
1#
1(
b101111101100100 +
b101111101100100 1
#661250000000
0#
0(
#661260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#661310000000
0$
0)
#661320000000
1"
1'
b0 +
b0 1
#661370000000
0"
0'
#661380000000
1#
1(
b101111101100100 +
b101111101100100 1
#661430000000
0#
0(
#661440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#661490000000
0$
0)
#661500000000
1"
1'
b0 +
b0 1
#661550000000
0"
0'
#661560000000
1#
1(
b101111101100100 +
b101111101100100 1
#661610000000
0#
0(
#661620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#661670000000
0$
0)
#661680000000
1"
1'
b0 +
b0 1
#661730000000
0"
0'
#661740000000
1#
1(
b101111101100100 +
b101111101100100 1
#661790000000
0#
0(
#661800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#661850000000
0$
0)
#661860000000
1"
1'
b0 +
b0 1
#661910000000
0"
0'
#661920000000
1#
1(
b101111101100100 +
b101111101100100 1
#661970000000
0#
0(
#661980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#662030000000
0$
0)
#662040000000
1"
1'
b0 +
b0 1
#662090000000
0"
0'
#662100000000
1#
1(
b101111101100100 +
b101111101100100 1
#662150000000
0#
0(
#662160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#662210000000
0$
0)
#662220000000
1"
1'
b0 +
b0 1
#662270000000
0"
0'
#662280000000
1#
1(
b101111101100100 +
b101111101100100 1
#662330000000
0#
0(
#662340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#662390000000
0$
0)
#662400000000
1"
1'
b0 +
b0 1
#662450000000
0"
0'
#662460000000
1#
1(
b101111101100100 +
b101111101100100 1
#662510000000
0#
0(
#662520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#662570000000
0$
0)
#662580000000
1"
1'
b0 +
b0 1
#662630000000
0"
0'
#662640000000
1#
1(
b101111101100100 +
b101111101100100 1
#662690000000
0#
0(
#662700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#662750000000
0$
0)
#662760000000
1"
1'
b0 +
b0 1
#662810000000
0"
0'
#662820000000
1#
1(
b101111101100100 +
b101111101100100 1
#662870000000
0#
0(
#662880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#662930000000
0$
0)
#662940000000
1"
1'
b0 +
b0 1
#662990000000
0"
0'
#663000000000
1#
1(
b101111101100100 +
b101111101100100 1
#663050000000
0#
0(
#663060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#663110000000
0$
0)
#663120000000
1"
1'
b0 +
b0 1
#663170000000
0"
0'
#663180000000
1#
1(
b101111101100100 +
b101111101100100 1
#663230000000
0#
0(
#663240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#663290000000
0$
0)
#663300000000
1"
1'
b0 +
b0 1
#663350000000
0"
0'
#663360000000
1#
1(
b101111101100100 +
b101111101100100 1
#663410000000
0#
0(
#663420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#663470000000
0$
0)
#663480000000
1"
1'
b0 +
b0 1
#663530000000
0"
0'
#663540000000
1#
1(
b101111101100100 +
b101111101100100 1
#663590000000
0#
0(
#663600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#663650000000
0$
0)
#663660000000
1"
1'
b0 +
b0 1
#663710000000
0"
0'
#663720000000
1#
1(
b101111101100100 +
b101111101100100 1
#663770000000
0#
0(
#663780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#663830000000
0$
0)
#663840000000
1"
1'
b0 +
b0 1
#663890000000
0"
0'
#663900000000
1#
1(
b101111101100100 +
b101111101100100 1
#663950000000
0#
0(
#663960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#664010000000
0$
0)
#664020000000
1"
1'
b0 +
b0 1
#664070000000
0"
0'
#664080000000
1#
1(
b101111101100100 +
b101111101100100 1
#664130000000
0#
0(
#664140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#664190000000
0$
0)
#664200000000
1"
1'
b0 +
b0 1
#664250000000
0"
0'
#664260000000
1#
1(
b101111101100100 +
b101111101100100 1
#664310000000
0#
0(
#664320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#664370000000
0$
0)
#664380000000
1"
1'
b0 +
b0 1
#664430000000
0"
0'
#664440000000
1#
1(
b101111101100100 +
b101111101100100 1
#664490000000
0#
0(
#664500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#664550000000
0$
0)
#664560000000
1"
1'
b0 +
b0 1
#664610000000
0"
0'
#664620000000
1#
1(
b101111101100100 +
b101111101100100 1
#664670000000
0#
0(
#664680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#664730000000
0$
0)
#664740000000
1"
1'
b0 +
b0 1
#664790000000
0"
0'
#664800000000
1#
1(
b101111101100100 +
b101111101100100 1
#664850000000
0#
0(
#664860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#664910000000
0$
0)
#664920000000
1"
1'
b0 +
b0 1
#664970000000
0"
0'
#664980000000
1#
1(
b101111101100100 +
b101111101100100 1
#665030000000
0#
0(
#665040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#665090000000
0$
0)
#665100000000
1"
1'
b0 +
b0 1
#665150000000
0"
0'
#665160000000
1#
1(
b101111101100100 +
b101111101100100 1
#665210000000
0#
0(
#665220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#665270000000
0$
0)
#665280000000
1"
1'
b0 +
b0 1
#665330000000
0"
0'
#665340000000
1#
1(
b101111101100100 +
b101111101100100 1
#665390000000
0#
0(
#665400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#665450000000
0$
0)
#665460000000
1"
1'
b0 +
b0 1
#665510000000
0"
0'
#665520000000
1#
1(
b101111101100100 +
b101111101100100 1
#665570000000
0#
0(
#665580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#665630000000
0$
0)
#665640000000
1"
1'
b0 +
b0 1
#665690000000
0"
0'
#665700000000
1#
1(
b101111101100100 +
b101111101100100 1
#665750000000
0#
0(
#665760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#665810000000
0$
0)
#665820000000
1"
1'
b0 +
b0 1
#665870000000
0"
0'
#665880000000
1#
1(
b101111101100100 +
b101111101100100 1
#665930000000
0#
0(
#665940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#665990000000
0$
0)
#666000000000
1"
1'
b0 +
b0 1
#666050000000
0"
0'
#666060000000
1#
1(
b101111101100100 +
b101111101100100 1
#666110000000
0#
0(
#666120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#666170000000
0$
0)
#666180000000
1"
1'
b0 +
b0 1
#666230000000
0"
0'
#666240000000
1#
1(
b101111101100100 +
b101111101100100 1
#666290000000
0#
0(
#666300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#666350000000
0$
0)
#666360000000
1"
1'
b0 +
b0 1
#666410000000
0"
0'
#666420000000
1#
1(
b101111101100100 +
b101111101100100 1
#666470000000
0#
0(
#666480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#666530000000
0$
0)
#666540000000
1"
1'
b0 +
b0 1
#666590000000
0"
0'
#666600000000
1#
1(
b101111101100100 +
b101111101100100 1
#666650000000
0#
0(
#666660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#666710000000
0$
0)
#666720000000
1"
1'
b0 +
b0 1
#666770000000
0"
0'
#666780000000
1#
1(
b101111101100100 +
b101111101100100 1
#666830000000
0#
0(
#666840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#666890000000
0$
0)
#666900000000
1"
1'
b0 +
b0 1
#666950000000
0"
0'
#666960000000
1#
1(
b101111101100100 +
b101111101100100 1
#667010000000
0#
0(
#667020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#667070000000
0$
0)
#667080000000
1"
1'
b0 +
b0 1
#667130000000
0"
0'
#667140000000
1#
1(
b101111101100100 +
b101111101100100 1
#667190000000
0#
0(
#667200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#667250000000
0$
0)
#667260000000
1"
1'
b0 +
b0 1
#667310000000
0"
0'
#667320000000
1#
1(
b101111101100100 +
b101111101100100 1
#667370000000
0#
0(
#667380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#667430000000
0$
0)
#667440000000
1"
1'
b0 +
b0 1
#667490000000
0"
0'
#667500000000
1#
1(
b101111101100100 +
b101111101100100 1
#667550000000
0#
0(
#667560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#667610000000
0$
0)
#667620000000
1"
1'
b0 +
b0 1
#667670000000
0"
0'
#667680000000
1#
1(
b101111101100100 +
b101111101100100 1
#667730000000
0#
0(
#667740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#667790000000
0$
0)
#667800000000
1"
1'
b0 +
b0 1
#667850000000
0"
0'
#667860000000
1#
1(
b101111101100100 +
b101111101100100 1
#667910000000
0#
0(
#667920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#667970000000
0$
0)
#667980000000
1"
1'
b0 +
b0 1
#668030000000
0"
0'
#668040000000
1#
1(
b101111101100100 +
b101111101100100 1
#668090000000
0#
0(
#668100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#668150000000
0$
0)
#668160000000
1"
1'
b0 +
b0 1
#668210000000
0"
0'
#668220000000
1#
1(
b101111101100100 +
b101111101100100 1
#668270000000
0#
0(
#668280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#668330000000
0$
0)
#668340000000
1"
1'
b0 +
b0 1
#668390000000
0"
0'
#668400000000
1#
1(
b101111101100100 +
b101111101100100 1
#668450000000
0#
0(
#668460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#668510000000
0$
0)
#668520000000
1"
1'
b0 +
b0 1
#668570000000
0"
0'
#668580000000
1#
1(
b101111101100100 +
b101111101100100 1
#668630000000
0#
0(
#668640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#668690000000
0$
0)
#668700000000
1"
1'
b0 +
b0 1
#668750000000
0"
0'
#668760000000
1#
1(
b101111101100100 +
b101111101100100 1
#668810000000
0#
0(
#668820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#668870000000
0$
0)
#668880000000
1"
1'
b0 +
b0 1
#668930000000
0"
0'
#668940000000
1#
1(
b101111101100100 +
b101111101100100 1
#668990000000
0#
0(
#669000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#669050000000
0$
0)
#669060000000
1"
1'
b0 +
b0 1
#669110000000
0"
0'
#669120000000
1#
1(
b101111101100100 +
b101111101100100 1
#669170000000
0#
0(
#669180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#669230000000
0$
0)
#669240000000
1"
1'
b0 +
b0 1
#669290000000
0"
0'
#669300000000
1#
1(
b101111101100100 +
b101111101100100 1
#669350000000
0#
0(
#669360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#669410000000
0$
0)
#669420000000
1"
1'
b0 +
b0 1
#669470000000
0"
0'
#669480000000
1#
1(
b101111101100100 +
b101111101100100 1
#669530000000
0#
0(
#669540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#669590000000
0$
0)
#669600000000
1"
1'
b0 +
b0 1
#669650000000
0"
0'
#669660000000
1#
1(
b101111101100100 +
b101111101100100 1
#669710000000
0#
0(
#669720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#669770000000
0$
0)
#669780000000
1"
1'
b0 +
b0 1
#669830000000
0"
0'
#669840000000
1#
1(
b101111101100100 +
b101111101100100 1
#669890000000
0#
0(
#669900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#669950000000
0$
0)
#669960000000
1"
1'
b0 +
b0 1
#670010000000
0"
0'
#670020000000
1#
1(
b101111101100100 +
b101111101100100 1
#670070000000
0#
0(
#670080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#670130000000
0$
0)
#670140000000
1"
1'
b0 +
b0 1
#670190000000
0"
0'
#670200000000
1#
1(
b101111101100100 +
b101111101100100 1
#670250000000
0#
0(
#670260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#670310000000
0$
0)
#670320000000
1"
1'
b0 +
b0 1
#670370000000
0"
0'
#670380000000
1#
1(
b101111101100100 +
b101111101100100 1
#670430000000
0#
0(
#670440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#670490000000
0$
0)
#670500000000
1"
1'
b0 +
b0 1
#670550000000
0"
0'
#670560000000
1#
1(
b101111101100100 +
b101111101100100 1
#670610000000
0#
0(
#670620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#670670000000
0$
0)
#670680000000
1"
1'
b0 +
b0 1
#670730000000
0"
0'
#670740000000
1#
1(
b101111101100100 +
b101111101100100 1
#670790000000
0#
0(
#670800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#670850000000
0$
0)
#670860000000
1"
1'
b0 +
b0 1
#670910000000
0"
0'
#670920000000
1#
1(
b101111101100100 +
b101111101100100 1
#670970000000
0#
0(
#670980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#671030000000
0$
0)
#671040000000
1"
1'
b0 +
b0 1
#671090000000
0"
0'
#671100000000
1#
1(
b101111101100100 +
b101111101100100 1
#671150000000
0#
0(
#671160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#671210000000
0$
0)
#671220000000
1"
1'
b0 +
b0 1
#671270000000
0"
0'
#671280000000
1#
1(
b101111101100100 +
b101111101100100 1
#671330000000
0#
0(
#671340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#671390000000
0$
0)
#671400000000
1"
1'
b0 +
b0 1
#671450000000
0"
0'
#671460000000
1#
1(
b101111101100100 +
b101111101100100 1
#671510000000
0#
0(
#671520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#671570000000
0$
0)
#671580000000
1"
1'
b0 +
b0 1
#671630000000
0"
0'
#671640000000
1#
1(
b101111101100100 +
b101111101100100 1
#671690000000
0#
0(
#671700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#671750000000
0$
0)
#671760000000
1"
1'
b0 +
b0 1
#671810000000
0"
0'
#671820000000
1#
1(
b101111101100100 +
b101111101100100 1
#671870000000
0#
0(
#671880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#671930000000
0$
0)
#671940000000
1"
1'
b0 +
b0 1
#671990000000
0"
0'
#672000000000
1#
1(
b101111101100100 +
b101111101100100 1
#672050000000
0#
0(
#672060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#672110000000
0$
0)
#672120000000
1"
1'
b0 +
b0 1
#672170000000
0"
0'
#672180000000
1#
1(
b101111101100100 +
b101111101100100 1
#672230000000
0#
0(
#672240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#672290000000
0$
0)
#672300000000
1"
1'
b0 +
b0 1
#672350000000
0"
0'
#672360000000
1#
1(
b101111101100100 +
b101111101100100 1
#672410000000
0#
0(
#672420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#672470000000
0$
0)
#672480000000
1"
1'
b0 +
b0 1
#672530000000
0"
0'
#672540000000
1#
1(
b101111101100100 +
b101111101100100 1
#672590000000
0#
0(
#672600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#672650000000
0$
0)
#672660000000
1"
1'
b0 +
b0 1
#672710000000
0"
0'
#672720000000
1#
1(
b101111101100100 +
b101111101100100 1
#672770000000
0#
0(
#672780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#672830000000
0$
0)
#672840000000
1"
1'
b0 +
b0 1
#672890000000
0"
0'
#672900000000
1#
1(
b101111101100100 +
b101111101100100 1
#672950000000
0#
0(
#672960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#673010000000
0$
0)
#673020000000
1"
1'
b0 +
b0 1
#673070000000
0"
0'
#673080000000
1#
1(
b101111101100100 +
b101111101100100 1
#673130000000
0#
0(
#673140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#673190000000
0$
0)
#673200000000
1"
1'
b0 +
b0 1
#673250000000
0"
0'
#673260000000
1#
1(
b101111101100100 +
b101111101100100 1
#673310000000
0#
0(
#673320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#673370000000
0$
0)
#673380000000
1"
1'
b0 +
b0 1
#673430000000
0"
0'
#673440000000
1#
1(
b101111101100100 +
b101111101100100 1
#673490000000
0#
0(
#673500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#673550000000
0$
0)
#673560000000
1"
1'
b0 +
b0 1
#673610000000
0"
0'
#673620000000
1#
1(
b101111101100100 +
b101111101100100 1
#673670000000
0#
0(
#673680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#673730000000
0$
0)
#673740000000
1"
1'
b0 +
b0 1
#673790000000
0"
0'
#673800000000
1#
1(
b101111101100100 +
b101111101100100 1
#673850000000
0#
0(
#673860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#673910000000
0$
0)
#673920000000
1"
1'
b0 +
b0 1
#673970000000
0"
0'
#673980000000
1#
1(
b101111101100100 +
b101111101100100 1
#674030000000
0#
0(
#674040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#674090000000
0$
0)
#674100000000
1"
1'
b0 +
b0 1
#674150000000
0"
0'
#674160000000
1#
1(
b101111101100100 +
b101111101100100 1
#674210000000
0#
0(
#674220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#674270000000
0$
0)
#674280000000
1"
1'
b0 +
b0 1
#674330000000
0"
0'
#674340000000
1#
1(
b101111101100100 +
b101111101100100 1
#674390000000
0#
0(
#674400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#674450000000
0$
0)
#674460000000
1"
1'
b0 +
b0 1
#674510000000
0"
0'
#674520000000
1#
1(
b101111101100100 +
b101111101100100 1
#674570000000
0#
0(
#674580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#674630000000
0$
0)
#674640000000
1"
1'
b0 +
b0 1
#674690000000
0"
0'
#674700000000
1#
1(
b101111101100100 +
b101111101100100 1
#674750000000
0#
0(
#674760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#674810000000
0$
0)
#674820000000
1"
1'
b0 +
b0 1
#674870000000
0"
0'
#674880000000
1#
1(
b101111101100100 +
b101111101100100 1
#674930000000
0#
0(
#674940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#674990000000
0$
0)
#675000000000
1"
1'
b0 +
b0 1
#675050000000
0"
0'
#675060000000
1#
1(
b101111101100100 +
b101111101100100 1
#675110000000
0#
0(
#675120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#675170000000
0$
0)
#675180000000
1"
1'
b0 +
b0 1
#675230000000
0"
0'
#675240000000
1#
1(
b101111101100100 +
b101111101100100 1
#675290000000
0#
0(
#675300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#675350000000
0$
0)
#675360000000
1"
1'
b0 +
b0 1
#675410000000
0"
0'
#675420000000
1#
1(
b101111101100100 +
b101111101100100 1
#675470000000
0#
0(
#675480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#675530000000
0$
0)
#675540000000
1"
1'
b0 +
b0 1
#675590000000
0"
0'
#675600000000
1#
1(
b101111101100100 +
b101111101100100 1
#675650000000
0#
0(
#675660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#675710000000
0$
0)
#675720000000
1"
1'
b0 +
b0 1
#675770000000
0"
0'
#675780000000
1#
1(
b101111101100100 +
b101111101100100 1
#675830000000
0#
0(
#675840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#675890000000
0$
0)
#675900000000
1"
1'
b0 +
b0 1
#675950000000
0"
0'
#675960000000
1#
1(
b101111101100100 +
b101111101100100 1
#676010000000
0#
0(
#676020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#676070000000
0$
0)
#676080000000
1"
1'
b0 +
b0 1
#676130000000
0"
0'
#676140000000
1#
1(
b101111101100100 +
b101111101100100 1
#676190000000
0#
0(
#676200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#676250000000
0$
0)
#676260000000
1"
1'
b0 +
b0 1
#676310000000
0"
0'
#676320000000
1#
1(
b101111101100100 +
b101111101100100 1
#676370000000
0#
0(
#676380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#676430000000
0$
0)
#676440000000
1"
1'
b0 +
b0 1
#676490000000
0"
0'
#676500000000
1#
1(
b101111101100100 +
b101111101100100 1
#676550000000
0#
0(
#676560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#676610000000
0$
0)
#676620000000
1"
1'
b0 +
b0 1
#676670000000
0"
0'
#676680000000
1#
1(
b101111101100100 +
b101111101100100 1
#676730000000
0#
0(
#676740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#676790000000
0$
0)
#676800000000
1"
1'
b0 +
b0 1
#676850000000
0"
0'
#676860000000
1#
1(
b101111101100100 +
b101111101100100 1
#676910000000
0#
0(
#676920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#676970000000
0$
0)
#676980000000
1"
1'
b0 +
b0 1
#677030000000
0"
0'
#677040000000
1#
1(
b101111101100100 +
b101111101100100 1
#677090000000
0#
0(
#677100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#677150000000
0$
0)
#677160000000
1"
1'
b0 +
b0 1
#677210000000
0"
0'
#677220000000
1#
1(
b101111101100100 +
b101111101100100 1
#677270000000
0#
0(
#677280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#677330000000
0$
0)
#677340000000
1"
1'
b0 +
b0 1
#677390000000
0"
0'
#677400000000
1#
1(
b101111101100100 +
b101111101100100 1
#677450000000
0#
0(
#677460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#677510000000
0$
0)
#677520000000
1"
1'
b0 +
b0 1
#677570000000
0"
0'
#677580000000
1#
1(
b101111101100100 +
b101111101100100 1
#677630000000
0#
0(
#677640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#677690000000
0$
0)
#677700000000
1"
1'
b0 +
b0 1
#677750000000
0"
0'
#677760000000
1#
1(
b101111101100100 +
b101111101100100 1
#677810000000
0#
0(
#677820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#677870000000
0$
0)
#677880000000
1"
1'
b0 +
b0 1
#677930000000
0"
0'
#677940000000
1#
1(
b101111101100100 +
b101111101100100 1
#677990000000
0#
0(
#678000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#678050000000
0$
0)
#678060000000
1"
1'
b0 +
b0 1
#678110000000
0"
0'
#678120000000
1#
1(
b101111101100100 +
b101111101100100 1
#678170000000
0#
0(
#678180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#678230000000
0$
0)
#678240000000
1"
1'
b0 +
b0 1
#678290000000
0"
0'
#678300000000
1#
1(
b101111101100100 +
b101111101100100 1
#678350000000
0#
0(
#678360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#678410000000
0$
0)
#678420000000
1"
1'
b0 +
b0 1
#678470000000
0"
0'
#678480000000
1#
1(
b101111101100100 +
b101111101100100 1
#678530000000
0#
0(
#678540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#678590000000
0$
0)
#678600000000
1"
1'
b0 +
b0 1
#678650000000
0"
0'
#678660000000
1#
1(
b101111101100100 +
b101111101100100 1
#678710000000
0#
0(
#678720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#678770000000
0$
0)
#678780000000
1"
1'
b0 +
b0 1
#678830000000
0"
0'
#678840000000
1#
1(
b101111101100100 +
b101111101100100 1
#678890000000
0#
0(
#678900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#678950000000
0$
0)
#678960000000
1"
1'
b0 +
b0 1
#679010000000
0"
0'
#679020000000
1#
1(
b101111101100100 +
b101111101100100 1
#679070000000
0#
0(
#679080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#679130000000
0$
0)
#679140000000
1"
1'
b0 +
b0 1
#679190000000
0"
0'
#679200000000
1#
1(
b101111101100100 +
b101111101100100 1
#679250000000
0#
0(
#679260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#679310000000
0$
0)
#679320000000
1"
1'
b0 +
b0 1
#679370000000
0"
0'
#679380000000
1#
1(
b101111101100100 +
b101111101100100 1
#679430000000
0#
0(
#679440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#679490000000
0$
0)
#679500000000
1"
1'
b0 +
b0 1
#679550000000
0"
0'
#679560000000
1#
1(
b101111101100100 +
b101111101100100 1
#679610000000
0#
0(
#679620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#679670000000
0$
0)
#679680000000
1"
1'
b0 +
b0 1
#679730000000
0"
0'
#679740000000
1#
1(
b101111101100100 +
b101111101100100 1
#679790000000
0#
0(
#679800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#679850000000
0$
0)
#679860000000
1"
1'
b0 +
b0 1
#679910000000
0"
0'
#679920000000
1#
1(
b101111101100100 +
b101111101100100 1
#679970000000
0#
0(
#679980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#680030000000
0$
0)
#680040000000
1"
1'
b0 +
b0 1
#680090000000
0"
0'
#680100000000
1#
1(
b101111101100100 +
b101111101100100 1
#680150000000
0#
0(
#680160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#680210000000
0$
0)
#680220000000
1"
1'
b0 +
b0 1
#680270000000
0"
0'
#680280000000
1#
1(
b101111101100100 +
b101111101100100 1
#680330000000
0#
0(
#680340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#680390000000
0$
0)
#680400000000
1"
1'
b0 +
b0 1
#680450000000
0"
0'
#680460000000
1#
1(
b101111101100100 +
b101111101100100 1
#680510000000
0#
0(
#680520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#680570000000
0$
0)
#680580000000
1"
1'
b0 +
b0 1
#680630000000
0"
0'
#680640000000
1#
1(
b101111101100100 +
b101111101100100 1
#680690000000
0#
0(
#680700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#680750000000
0$
0)
#680760000000
1"
1'
b0 +
b0 1
#680810000000
0"
0'
#680820000000
1#
1(
b101111101100100 +
b101111101100100 1
#680870000000
0#
0(
#680880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#680930000000
0$
0)
#680940000000
1"
1'
b0 +
b0 1
#680990000000
0"
0'
#681000000000
1#
1(
b101111101100100 +
b101111101100100 1
#681050000000
0#
0(
#681060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#681110000000
0$
0)
#681120000000
1"
1'
b0 +
b0 1
#681170000000
0"
0'
#681180000000
1#
1(
b101111101100100 +
b101111101100100 1
#681230000000
0#
0(
#681240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#681290000000
0$
0)
#681300000000
1"
1'
b0 +
b0 1
#681350000000
0"
0'
#681360000000
1#
1(
b101111101100100 +
b101111101100100 1
#681410000000
0#
0(
#681420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#681470000000
0$
0)
#681480000000
1"
1'
b0 +
b0 1
#681530000000
0"
0'
#681540000000
1#
1(
b101111101100100 +
b101111101100100 1
#681590000000
0#
0(
#681600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#681650000000
0$
0)
#681660000000
1"
1'
b0 +
b0 1
#681710000000
0"
0'
#681720000000
1#
1(
b101111101100100 +
b101111101100100 1
#681770000000
0#
0(
#681780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#681830000000
0$
0)
#681840000000
1"
1'
b0 +
b0 1
#681890000000
0"
0'
#681900000000
1#
1(
b101111101100100 +
b101111101100100 1
#681950000000
0#
0(
#681960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#682010000000
0$
0)
#682020000000
1"
1'
b0 +
b0 1
#682070000000
0"
0'
#682080000000
1#
1(
b101111101100100 +
b101111101100100 1
#682130000000
0#
0(
#682140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#682190000000
0$
0)
#682200000000
1"
1'
b0 +
b0 1
#682250000000
0"
0'
#682260000000
1#
1(
b101111101100100 +
b101111101100100 1
#682310000000
0#
0(
#682320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#682370000000
0$
0)
#682380000000
1"
1'
b0 +
b0 1
#682430000000
0"
0'
#682440000000
1#
1(
b101111101100100 +
b101111101100100 1
#682490000000
0#
0(
#682500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#682550000000
0$
0)
#682560000000
1"
1'
b0 +
b0 1
#682610000000
0"
0'
#682620000000
1#
1(
b101111101100100 +
b101111101100100 1
#682670000000
0#
0(
#682680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#682730000000
0$
0)
#682740000000
1"
1'
b0 +
b0 1
#682790000000
0"
0'
#682800000000
1#
1(
b101111101100100 +
b101111101100100 1
#682850000000
0#
0(
#682860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#682910000000
0$
0)
#682920000000
1"
1'
b0 +
b0 1
#682970000000
0"
0'
#682980000000
1#
1(
b101111101100100 +
b101111101100100 1
#683030000000
0#
0(
#683040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#683090000000
0$
0)
#683100000000
1"
1'
b0 +
b0 1
#683150000000
0"
0'
#683160000000
1#
1(
b101111101100100 +
b101111101100100 1
#683210000000
0#
0(
#683220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#683270000000
0$
0)
#683280000000
1"
1'
b0 +
b0 1
#683330000000
0"
0'
#683340000000
1#
1(
b101111101100100 +
b101111101100100 1
#683390000000
0#
0(
#683400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#683450000000
0$
0)
#683460000000
1"
1'
b0 +
b0 1
#683510000000
0"
0'
#683520000000
1#
1(
b101111101100100 +
b101111101100100 1
#683570000000
0#
0(
#683580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#683630000000
0$
0)
#683640000000
1"
1'
b0 +
b0 1
#683690000000
0"
0'
#683700000000
1#
1(
b101111101100100 +
b101111101100100 1
#683750000000
0#
0(
#683760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#683810000000
0$
0)
#683820000000
1"
1'
b0 +
b0 1
#683870000000
0"
0'
#683880000000
1#
1(
b101111101100100 +
b101111101100100 1
#683930000000
0#
0(
#683940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#683990000000
0$
0)
#684000000000
1"
1'
b0 +
b0 1
#684050000000
0"
0'
#684060000000
1#
1(
b101111101100100 +
b101111101100100 1
#684110000000
0#
0(
#684120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#684170000000
0$
0)
#684180000000
1"
1'
b0 +
b0 1
#684230000000
0"
0'
#684240000000
1#
1(
b101111101100100 +
b101111101100100 1
#684290000000
0#
0(
#684300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#684350000000
0$
0)
#684360000000
1"
1'
b0 +
b0 1
#684410000000
0"
0'
#684420000000
1#
1(
b101111101100100 +
b101111101100100 1
#684470000000
0#
0(
#684480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#684530000000
0$
0)
#684540000000
1"
1'
b0 +
b0 1
#684590000000
0"
0'
#684600000000
1#
1(
b101111101100100 +
b101111101100100 1
#684650000000
0#
0(
#684660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#684710000000
0$
0)
#684720000000
1"
1'
b0 +
b0 1
#684770000000
0"
0'
#684780000000
1#
1(
b101111101100100 +
b101111101100100 1
#684830000000
0#
0(
#684840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#684890000000
0$
0)
#684900000000
1"
1'
b0 +
b0 1
#684950000000
0"
0'
#684960000000
1#
1(
b101111101100100 +
b101111101100100 1
#685010000000
0#
0(
#685020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#685070000000
0$
0)
#685080000000
1"
1'
b0 +
b0 1
#685130000000
0"
0'
#685140000000
1#
1(
b101111101100100 +
b101111101100100 1
#685190000000
0#
0(
#685200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#685250000000
0$
0)
#685260000000
1"
1'
b0 +
b0 1
#685310000000
0"
0'
#685320000000
1#
1(
b101111101100100 +
b101111101100100 1
#685370000000
0#
0(
#685380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#685430000000
0$
0)
#685440000000
1"
1'
b0 +
b0 1
#685490000000
0"
0'
#685500000000
1#
1(
b101111101100100 +
b101111101100100 1
#685550000000
0#
0(
#685560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#685610000000
0$
0)
#685620000000
1"
1'
b0 +
b0 1
#685670000000
0"
0'
#685680000000
1#
1(
b101111101100100 +
b101111101100100 1
#685730000000
0#
0(
#685740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#685790000000
0$
0)
#685800000000
1"
1'
b0 +
b0 1
#685850000000
0"
0'
#685860000000
1#
1(
b101111101100100 +
b101111101100100 1
#685910000000
0#
0(
#685920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#685970000000
0$
0)
#685980000000
1"
1'
b0 +
b0 1
#686030000000
0"
0'
#686040000000
1#
1(
b101111101100100 +
b101111101100100 1
#686090000000
0#
0(
#686100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#686150000000
0$
0)
#686160000000
1"
1'
b0 +
b0 1
#686210000000
0"
0'
#686220000000
1#
1(
b101111101100100 +
b101111101100100 1
#686270000000
0#
0(
#686280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#686330000000
0$
0)
#686340000000
1"
1'
b0 +
b0 1
#686390000000
0"
0'
#686400000000
1#
1(
b101111101100100 +
b101111101100100 1
#686450000000
0#
0(
#686460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#686510000000
0$
0)
#686520000000
1"
1'
b0 +
b0 1
#686570000000
0"
0'
#686580000000
1#
1(
b101111101100100 +
b101111101100100 1
#686630000000
0#
0(
#686640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#686690000000
0$
0)
#686700000000
1"
1'
b0 +
b0 1
#686750000000
0"
0'
#686760000000
1#
1(
b101111101100100 +
b101111101100100 1
#686810000000
0#
0(
#686820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#686870000000
0$
0)
#686880000000
1"
1'
b0 +
b0 1
#686930000000
0"
0'
#686940000000
1#
1(
b101111101100100 +
b101111101100100 1
#686990000000
0#
0(
#687000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#687050000000
0$
0)
#687060000000
1"
1'
b0 +
b0 1
#687110000000
0"
0'
#687120000000
1#
1(
b101111101100100 +
b101111101100100 1
#687170000000
0#
0(
#687180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#687230000000
0$
0)
#687240000000
1"
1'
b0 +
b0 1
#687290000000
0"
0'
#687300000000
1#
1(
b101111101100100 +
b101111101100100 1
#687350000000
0#
0(
#687360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#687410000000
0$
0)
#687420000000
1"
1'
b0 +
b0 1
#687470000000
0"
0'
#687480000000
1#
1(
b101111101100100 +
b101111101100100 1
#687530000000
0#
0(
#687540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#687590000000
0$
0)
#687600000000
1"
1'
b0 +
b0 1
#687650000000
0"
0'
#687660000000
1#
1(
b101111101100100 +
b101111101100100 1
#687710000000
0#
0(
#687720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#687770000000
0$
0)
#687780000000
1"
1'
b0 +
b0 1
#687830000000
0"
0'
#687840000000
1#
1(
b101111101100100 +
b101111101100100 1
#687890000000
0#
0(
#687900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#687950000000
0$
0)
#687960000000
1"
1'
b0 +
b0 1
#688010000000
0"
0'
#688020000000
1#
1(
b101111101100100 +
b101111101100100 1
#688070000000
0#
0(
#688080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#688130000000
0$
0)
#688140000000
1"
1'
b0 +
b0 1
#688190000000
0"
0'
#688200000000
1#
1(
b101111101100100 +
b101111101100100 1
#688250000000
0#
0(
#688260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#688310000000
0$
0)
#688320000000
1"
1'
b0 +
b0 1
#688370000000
0"
0'
#688380000000
1#
1(
b101111101100100 +
b101111101100100 1
#688430000000
0#
0(
#688440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#688490000000
0$
0)
#688500000000
1"
1'
b0 +
b0 1
#688550000000
0"
0'
#688560000000
1#
1(
b101111101100100 +
b101111101100100 1
#688610000000
0#
0(
#688620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#688670000000
0$
0)
#688680000000
1"
1'
b0 +
b0 1
#688730000000
0"
0'
#688740000000
1#
1(
b101111101100100 +
b101111101100100 1
#688790000000
0#
0(
#688800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#688850000000
0$
0)
#688860000000
1"
1'
b0 +
b0 1
#688910000000
0"
0'
#688920000000
1#
1(
b101111101100100 +
b101111101100100 1
#688970000000
0#
0(
#688980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#689030000000
0$
0)
#689040000000
1"
1'
b0 +
b0 1
#689090000000
0"
0'
#689100000000
1#
1(
b101111101100100 +
b101111101100100 1
#689150000000
0#
0(
#689160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#689210000000
0$
0)
#689220000000
1"
1'
b0 +
b0 1
#689270000000
0"
0'
#689280000000
1#
1(
b101111101100100 +
b101111101100100 1
#689330000000
0#
0(
#689340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#689390000000
0$
0)
#689400000000
1"
1'
b0 +
b0 1
#689450000000
0"
0'
#689460000000
1#
1(
b101111101100100 +
b101111101100100 1
#689510000000
0#
0(
#689520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#689570000000
0$
0)
#689580000000
1"
1'
b0 +
b0 1
#689630000000
0"
0'
#689640000000
1#
1(
b101111101100100 +
b101111101100100 1
#689690000000
0#
0(
#689700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#689750000000
0$
0)
#689760000000
1"
1'
b0 +
b0 1
#689810000000
0"
0'
#689820000000
1#
1(
b101111101100100 +
b101111101100100 1
#689870000000
0#
0(
#689880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#689930000000
0$
0)
#689940000000
1"
1'
b0 +
b0 1
#689990000000
0"
0'
#690000000000
1#
1(
b101111101100100 +
b101111101100100 1
#690050000000
0#
0(
#690060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#690110000000
0$
0)
#690120000000
1"
1'
b0 +
b0 1
#690170000000
0"
0'
#690180000000
1#
1(
b101111101100100 +
b101111101100100 1
#690230000000
0#
0(
#690240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#690290000000
0$
0)
#690300000000
1"
1'
b0 +
b0 1
#690350000000
0"
0'
#690360000000
1#
1(
b101111101100100 +
b101111101100100 1
#690410000000
0#
0(
#690420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#690470000000
0$
0)
#690480000000
1"
1'
b0 +
b0 1
#690530000000
0"
0'
#690540000000
1#
1(
b101111101100100 +
b101111101100100 1
#690590000000
0#
0(
#690600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#690650000000
0$
0)
#690660000000
1"
1'
b0 +
b0 1
#690710000000
0"
0'
#690720000000
1#
1(
b101111101100100 +
b101111101100100 1
#690770000000
0#
0(
#690780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#690830000000
0$
0)
#690840000000
1"
1'
b0 +
b0 1
#690890000000
0"
0'
#690900000000
1#
1(
b101111101100100 +
b101111101100100 1
#690950000000
0#
0(
#690960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#691010000000
0$
0)
#691020000000
1"
1'
b0 +
b0 1
#691070000000
0"
0'
#691080000000
1#
1(
b101111101100100 +
b101111101100100 1
#691130000000
0#
0(
#691140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#691190000000
0$
0)
#691200000000
1"
1'
b0 +
b0 1
#691250000000
0"
0'
#691260000000
1#
1(
b101111101100100 +
b101111101100100 1
#691310000000
0#
0(
#691320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#691370000000
0$
0)
#691380000000
1"
1'
b0 +
b0 1
#691430000000
0"
0'
#691440000000
1#
1(
b101111101100100 +
b101111101100100 1
#691490000000
0#
0(
#691500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#691550000000
0$
0)
#691560000000
1"
1'
b0 +
b0 1
#691610000000
0"
0'
#691620000000
1#
1(
b101111101100100 +
b101111101100100 1
#691670000000
0#
0(
#691680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#691730000000
0$
0)
#691740000000
1"
1'
b0 +
b0 1
#691790000000
0"
0'
#691800000000
1#
1(
b101111101100100 +
b101111101100100 1
#691850000000
0#
0(
#691860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#691910000000
0$
0)
#691920000000
1"
1'
b0 +
b0 1
#691970000000
0"
0'
#691980000000
1#
1(
b101111101100100 +
b101111101100100 1
#692030000000
0#
0(
#692040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#692090000000
0$
0)
#692100000000
1"
1'
b0 +
b0 1
#692150000000
0"
0'
#692160000000
1#
1(
b101111101100100 +
b101111101100100 1
#692210000000
0#
0(
#692220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#692270000000
0$
0)
#692280000000
1"
1'
b0 +
b0 1
#692330000000
0"
0'
#692340000000
1#
1(
b101111101100100 +
b101111101100100 1
#692390000000
0#
0(
#692400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#692450000000
0$
0)
#692460000000
1"
1'
b0 +
b0 1
#692510000000
0"
0'
#692520000000
1#
1(
b101111101100100 +
b101111101100100 1
#692570000000
0#
0(
#692580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#692630000000
0$
0)
#692640000000
1"
1'
b0 +
b0 1
#692690000000
0"
0'
#692700000000
1#
1(
b101111101100100 +
b101111101100100 1
#692750000000
0#
0(
#692760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#692810000000
0$
0)
#692820000000
1"
1'
b0 +
b0 1
#692870000000
0"
0'
#692880000000
1#
1(
b101111101100100 +
b101111101100100 1
#692930000000
0#
0(
#692940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#692990000000
0$
0)
#693000000000
1"
1'
b0 +
b0 1
#693050000000
0"
0'
#693060000000
1#
1(
b101111101100100 +
b101111101100100 1
#693110000000
0#
0(
#693120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#693170000000
0$
0)
#693180000000
1"
1'
b0 +
b0 1
#693230000000
0"
0'
#693240000000
1#
1(
b101111101100100 +
b101111101100100 1
#693290000000
0#
0(
#693300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#693350000000
0$
0)
#693360000000
1"
1'
b0 +
b0 1
#693410000000
0"
0'
#693420000000
1#
1(
b101111101100100 +
b101111101100100 1
#693470000000
0#
0(
#693480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#693530000000
0$
0)
#693540000000
1"
1'
b0 +
b0 1
#693590000000
0"
0'
#693600000000
1#
1(
b101111101100100 +
b101111101100100 1
#693650000000
0#
0(
#693660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#693710000000
0$
0)
#693720000000
1"
1'
b0 +
b0 1
#693770000000
0"
0'
#693780000000
1#
1(
b101111101100100 +
b101111101100100 1
#693830000000
0#
0(
#693840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#693890000000
0$
0)
#693900000000
1"
1'
b0 +
b0 1
#693950000000
0"
0'
#693960000000
1#
1(
b101111101100100 +
b101111101100100 1
#694010000000
0#
0(
#694020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#694070000000
0$
0)
#694080000000
1"
1'
b0 +
b0 1
#694130000000
0"
0'
#694140000000
1#
1(
b101111101100100 +
b101111101100100 1
#694190000000
0#
0(
#694200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#694250000000
0$
0)
#694260000000
1"
1'
b0 +
b0 1
#694310000000
0"
0'
#694320000000
1#
1(
b101111101100100 +
b101111101100100 1
#694370000000
0#
0(
#694380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#694430000000
0$
0)
#694440000000
1"
1'
b0 +
b0 1
#694490000000
0"
0'
#694500000000
1#
1(
b101111101100100 +
b101111101100100 1
#694550000000
0#
0(
#694560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#694610000000
0$
0)
#694620000000
1"
1'
b0 +
b0 1
#694670000000
0"
0'
#694680000000
1#
1(
b101111101100100 +
b101111101100100 1
#694730000000
0#
0(
#694740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#694790000000
0$
0)
#694800000000
1"
1'
b0 +
b0 1
#694850000000
0"
0'
#694860000000
1#
1(
b101111101100100 +
b101111101100100 1
#694910000000
0#
0(
#694920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#694970000000
0$
0)
#694980000000
1"
1'
b0 +
b0 1
#695030000000
0"
0'
#695040000000
1#
1(
b101111101100100 +
b101111101100100 1
#695090000000
0#
0(
#695100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#695150000000
0$
0)
#695160000000
1"
1'
b0 +
b0 1
#695210000000
0"
0'
#695220000000
1#
1(
b101111101100100 +
b101111101100100 1
#695270000000
0#
0(
#695280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#695330000000
0$
0)
#695340000000
1"
1'
b0 +
b0 1
#695390000000
0"
0'
#695400000000
1#
1(
b101111101100100 +
b101111101100100 1
#695450000000
0#
0(
#695460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#695510000000
0$
0)
#695520000000
1"
1'
b0 +
b0 1
#695570000000
0"
0'
#695580000000
1#
1(
b101111101100100 +
b101111101100100 1
#695630000000
0#
0(
#695640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#695690000000
0$
0)
#695700000000
1"
1'
b0 +
b0 1
#695750000000
0"
0'
#695760000000
1#
1(
b101111101100100 +
b101111101100100 1
#695810000000
0#
0(
#695820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#695870000000
0$
0)
#695880000000
1"
1'
b0 +
b0 1
#695930000000
0"
0'
#695940000000
1#
1(
b101111101100100 +
b101111101100100 1
#695990000000
0#
0(
#696000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#696050000000
0$
0)
#696060000000
1"
1'
b0 +
b0 1
#696110000000
0"
0'
#696120000000
1#
1(
b101111101100100 +
b101111101100100 1
#696170000000
0#
0(
#696180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#696230000000
0$
0)
#696240000000
1"
1'
b0 +
b0 1
#696290000000
0"
0'
#696300000000
1#
1(
b101111101100100 +
b101111101100100 1
#696350000000
0#
0(
#696360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#696410000000
0$
0)
#696420000000
1"
1'
b0 +
b0 1
#696470000000
0"
0'
#696480000000
1#
1(
b101111101100100 +
b101111101100100 1
#696530000000
0#
0(
#696540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#696590000000
0$
0)
#696600000000
1"
1'
b0 +
b0 1
#696650000000
0"
0'
#696660000000
1#
1(
b101111101100100 +
b101111101100100 1
#696710000000
0#
0(
#696720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#696770000000
0$
0)
#696780000000
1"
1'
b0 +
b0 1
#696830000000
0"
0'
#696840000000
1#
1(
b101111101100100 +
b101111101100100 1
#696890000000
0#
0(
#696900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#696950000000
0$
0)
#696960000000
1"
1'
b0 +
b0 1
#697010000000
0"
0'
#697020000000
1#
1(
b101111101100100 +
b101111101100100 1
#697070000000
0#
0(
#697080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#697130000000
0$
0)
#697140000000
1"
1'
b0 +
b0 1
#697190000000
0"
0'
#697200000000
1#
1(
b101111101100100 +
b101111101100100 1
#697250000000
0#
0(
#697260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#697310000000
0$
0)
#697320000000
1"
1'
b0 +
b0 1
#697370000000
0"
0'
#697380000000
1#
1(
b101111101100100 +
b101111101100100 1
#697430000000
0#
0(
#697440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#697490000000
0$
0)
#697500000000
1"
1'
b0 +
b0 1
#697550000000
0"
0'
#697560000000
1#
1(
b101111101100100 +
b101111101100100 1
#697610000000
0#
0(
#697620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#697670000000
0$
0)
#697680000000
1"
1'
b0 +
b0 1
#697730000000
0"
0'
#697740000000
1#
1(
b101111101100100 +
b101111101100100 1
#697790000000
0#
0(
#697800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#697850000000
0$
0)
#697860000000
1"
1'
b0 +
b0 1
#697910000000
0"
0'
#697920000000
1#
1(
b101111101100100 +
b101111101100100 1
#697970000000
0#
0(
#697980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#698030000000
0$
0)
#698040000000
1"
1'
b0 +
b0 1
#698090000000
0"
0'
#698100000000
1#
1(
b101111101100100 +
b101111101100100 1
#698150000000
0#
0(
#698160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#698210000000
0$
0)
#698220000000
1"
1'
b0 +
b0 1
#698270000000
0"
0'
#698280000000
1#
1(
b101111101100100 +
b101111101100100 1
#698330000000
0#
0(
#698340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#698390000000
0$
0)
#698400000000
1"
1'
b0 +
b0 1
#698450000000
0"
0'
#698460000000
1#
1(
b101111101100100 +
b101111101100100 1
#698510000000
0#
0(
#698520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#698570000000
0$
0)
#698580000000
1"
1'
b0 +
b0 1
#698630000000
0"
0'
#698640000000
1#
1(
b101111101100100 +
b101111101100100 1
#698690000000
0#
0(
#698700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#698750000000
0$
0)
#698760000000
1"
1'
b0 +
b0 1
#698810000000
0"
0'
#698820000000
1#
1(
b101111101100100 +
b101111101100100 1
#698870000000
0#
0(
#698880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#698930000000
0$
0)
#698940000000
1"
1'
b0 +
b0 1
#698990000000
0"
0'
#699000000000
1#
1(
b101111101100100 +
b101111101100100 1
#699050000000
0#
0(
#699060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#699110000000
0$
0)
#699120000000
1"
1'
b0 +
b0 1
#699170000000
0"
0'
#699180000000
1#
1(
b101111101100100 +
b101111101100100 1
#699230000000
0#
0(
#699240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#699290000000
0$
0)
#699300000000
1"
1'
b0 +
b0 1
#699350000000
0"
0'
#699360000000
1#
1(
b101111101100100 +
b101111101100100 1
#699410000000
0#
0(
#699420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#699470000000
0$
0)
#699480000000
1"
1'
b0 +
b0 1
#699530000000
0"
0'
#699540000000
1#
1(
b101111101100100 +
b101111101100100 1
#699590000000
0#
0(
#699600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#699650000000
0$
0)
#699660000000
1"
1'
b0 +
b0 1
#699710000000
0"
0'
#699720000000
1#
1(
b101111101100100 +
b101111101100100 1
#699770000000
0#
0(
#699780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#699830000000
0$
0)
#699840000000
1"
1'
b0 +
b0 1
#699890000000
0"
0'
#699900000000
1#
1(
b101111101100100 +
b101111101100100 1
#699950000000
0#
0(
#699960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#700010000000
0$
0)
#700020000000
1"
1'
b0 +
b0 1
#700070000000
0"
0'
#700080000000
1#
1(
b101111101100100 +
b101111101100100 1
#700130000000
0#
0(
#700140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#700190000000
0$
0)
#700200000000
1"
1'
b0 +
b0 1
#700250000000
0"
0'
#700260000000
1#
1(
b101111101100100 +
b101111101100100 1
#700310000000
0#
0(
#700320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#700370000000
0$
0)
#700380000000
1"
1'
b0 +
b0 1
#700430000000
0"
0'
#700440000000
1#
1(
b101111101100100 +
b101111101100100 1
#700490000000
0#
0(
#700500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#700550000000
0$
0)
#700560000000
1"
1'
b0 +
b0 1
#700610000000
0"
0'
#700620000000
1#
1(
b101111101100100 +
b101111101100100 1
#700670000000
0#
0(
#700680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#700730000000
0$
0)
#700740000000
1"
1'
b0 +
b0 1
#700790000000
0"
0'
#700800000000
1#
1(
b101111101100100 +
b101111101100100 1
#700850000000
0#
0(
#700860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#700910000000
0$
0)
#700920000000
1"
1'
b0 +
b0 1
#700970000000
0"
0'
#700980000000
1#
1(
b101111101100100 +
b101111101100100 1
#701030000000
0#
0(
#701040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#701090000000
0$
0)
#701100000000
1"
1'
b0 +
b0 1
#701150000000
0"
0'
#701160000000
1#
1(
b101111101100100 +
b101111101100100 1
#701210000000
0#
0(
#701220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#701270000000
0$
0)
#701280000000
1"
1'
b0 +
b0 1
#701330000000
0"
0'
#701340000000
1#
1(
b101111101100100 +
b101111101100100 1
#701390000000
0#
0(
#701400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#701450000000
0$
0)
#701460000000
1"
1'
b0 +
b0 1
#701510000000
0"
0'
#701520000000
1#
1(
b101111101100100 +
b101111101100100 1
#701570000000
0#
0(
#701580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#701630000000
0$
0)
#701640000000
1"
1'
b0 +
b0 1
#701690000000
0"
0'
#701700000000
1#
1(
b101111101100100 +
b101111101100100 1
#701750000000
0#
0(
#701760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#701810000000
0$
0)
#701820000000
1"
1'
b0 +
b0 1
#701870000000
0"
0'
#701880000000
1#
1(
b101111101100100 +
b101111101100100 1
#701930000000
0#
0(
#701940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#701990000000
0$
0)
#702000000000
1"
1'
b0 +
b0 1
#702050000000
0"
0'
#702060000000
1#
1(
b101111101100100 +
b101111101100100 1
#702110000000
0#
0(
#702120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#702170000000
0$
0)
#702180000000
1"
1'
b0 +
b0 1
#702230000000
0"
0'
#702240000000
1#
1(
b101111101100100 +
b101111101100100 1
#702290000000
0#
0(
#702300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#702350000000
0$
0)
#702360000000
1"
1'
b0 +
b0 1
#702410000000
0"
0'
#702420000000
1#
1(
b101111101100100 +
b101111101100100 1
#702470000000
0#
0(
#702480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#702530000000
0$
0)
#702540000000
1"
1'
b0 +
b0 1
#702590000000
0"
0'
#702600000000
1#
1(
b101111101100100 +
b101111101100100 1
#702650000000
0#
0(
#702660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#702710000000
0$
0)
#702720000000
1"
1'
b0 +
b0 1
#702770000000
0"
0'
#702780000000
1#
1(
b101111101100100 +
b101111101100100 1
#702830000000
0#
0(
#702840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#702890000000
0$
0)
#702900000000
1"
1'
b0 +
b0 1
#702950000000
0"
0'
#702960000000
1#
1(
b101111101100100 +
b101111101100100 1
#703010000000
0#
0(
#703020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#703070000000
0$
0)
#703080000000
1"
1'
b0 +
b0 1
#703130000000
0"
0'
#703140000000
1#
1(
b101111101100100 +
b101111101100100 1
#703190000000
0#
0(
#703200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#703250000000
0$
0)
#703260000000
1"
1'
b0 +
b0 1
#703310000000
0"
0'
#703320000000
1#
1(
b101111101100100 +
b101111101100100 1
#703370000000
0#
0(
#703380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#703430000000
0$
0)
#703440000000
1"
1'
b0 +
b0 1
#703490000000
0"
0'
#703500000000
1#
1(
b101111101100100 +
b101111101100100 1
#703550000000
0#
0(
#703560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#703610000000
0$
0)
#703620000000
1"
1'
b0 +
b0 1
#703670000000
0"
0'
#703680000000
1#
1(
b101111101100100 +
b101111101100100 1
#703730000000
0#
0(
#703740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#703790000000
0$
0)
#703800000000
1"
1'
b0 +
b0 1
#703850000000
0"
0'
#703860000000
1#
1(
b101111101100100 +
b101111101100100 1
#703910000000
0#
0(
#703920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#703970000000
0$
0)
#703980000000
1"
1'
b0 +
b0 1
#704030000000
0"
0'
#704040000000
1#
1(
b101111101100100 +
b101111101100100 1
#704090000000
0#
0(
#704100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#704150000000
0$
0)
#704160000000
1"
1'
b0 +
b0 1
#704210000000
0"
0'
#704220000000
1#
1(
b101111101100100 +
b101111101100100 1
#704270000000
0#
0(
#704280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#704330000000
0$
0)
#704340000000
1"
1'
b0 +
b0 1
#704390000000
0"
0'
#704400000000
1#
1(
b101111101100100 +
b101111101100100 1
#704450000000
0#
0(
#704460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#704510000000
0$
0)
#704520000000
1"
1'
b0 +
b0 1
#704570000000
0"
0'
#704580000000
1#
1(
b101111101100100 +
b101111101100100 1
#704630000000
0#
0(
#704640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#704690000000
0$
0)
#704700000000
1"
1'
b0 +
b0 1
#704750000000
0"
0'
#704760000000
1#
1(
b101111101100100 +
b101111101100100 1
#704810000000
0#
0(
#704820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#704870000000
0$
0)
#704880000000
1"
1'
b0 +
b0 1
#704930000000
0"
0'
#704940000000
1#
1(
b101111101100100 +
b101111101100100 1
#704990000000
0#
0(
#705000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#705050000000
0$
0)
#705060000000
1"
1'
b0 +
b0 1
#705110000000
0"
0'
#705120000000
1#
1(
b101111101100100 +
b101111101100100 1
#705170000000
0#
0(
#705180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#705230000000
0$
0)
#705240000000
1"
1'
b0 +
b0 1
#705290000000
0"
0'
#705300000000
1#
1(
b101111101100100 +
b101111101100100 1
#705350000000
0#
0(
#705360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#705410000000
0$
0)
#705420000000
1"
1'
b0 +
b0 1
#705470000000
0"
0'
#705480000000
1#
1(
b101111101100100 +
b101111101100100 1
#705530000000
0#
0(
#705540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#705590000000
0$
0)
#705600000000
1"
1'
b0 +
b0 1
#705650000000
0"
0'
#705660000000
1#
1(
b101111101100100 +
b101111101100100 1
#705710000000
0#
0(
#705720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#705770000000
0$
0)
#705780000000
1"
1'
b0 +
b0 1
#705830000000
0"
0'
#705840000000
1#
1(
b101111101100100 +
b101111101100100 1
#705890000000
0#
0(
#705900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#705950000000
0$
0)
#705960000000
1"
1'
b0 +
b0 1
#706010000000
0"
0'
#706020000000
1#
1(
b101111101100100 +
b101111101100100 1
#706070000000
0#
0(
#706080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#706130000000
0$
0)
#706140000000
1"
1'
b0 +
b0 1
#706190000000
0"
0'
#706200000000
1#
1(
b101111101100100 +
b101111101100100 1
#706250000000
0#
0(
#706260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#706310000000
0$
0)
#706320000000
1"
1'
b0 +
b0 1
#706370000000
0"
0'
#706380000000
1#
1(
b101111101100100 +
b101111101100100 1
#706430000000
0#
0(
#706440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#706490000000
0$
0)
#706500000000
1"
1'
b0 +
b0 1
#706550000000
0"
0'
#706560000000
1#
1(
b101111101100100 +
b101111101100100 1
#706610000000
0#
0(
#706620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#706670000000
0$
0)
#706680000000
1"
1'
b0 +
b0 1
#706730000000
0"
0'
#706740000000
1#
1(
b101111101100100 +
b101111101100100 1
#706790000000
0#
0(
#706800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#706850000000
0$
0)
#706860000000
1"
1'
b0 +
b0 1
#706910000000
0"
0'
#706920000000
1#
1(
b101111101100100 +
b101111101100100 1
#706970000000
0#
0(
#706980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#707030000000
0$
0)
#707040000000
1"
1'
b0 +
b0 1
#707090000000
0"
0'
#707100000000
1#
1(
b101111101100100 +
b101111101100100 1
#707150000000
0#
0(
#707160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#707210000000
0$
0)
#707220000000
1"
1'
b0 +
b0 1
#707270000000
0"
0'
#707280000000
1#
1(
b101111101100100 +
b101111101100100 1
#707330000000
0#
0(
#707340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#707390000000
0$
0)
#707400000000
1"
1'
b0 +
b0 1
#707450000000
0"
0'
#707460000000
1#
1(
b101111101100100 +
b101111101100100 1
#707510000000
0#
0(
#707520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#707570000000
0$
0)
#707580000000
1"
1'
b0 +
b0 1
#707630000000
0"
0'
#707640000000
1#
1(
b101111101100100 +
b101111101100100 1
#707690000000
0#
0(
#707700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#707750000000
0$
0)
#707760000000
1"
1'
b0 +
b0 1
#707810000000
0"
0'
#707820000000
1#
1(
b101111101100100 +
b101111101100100 1
#707870000000
0#
0(
#707880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#707930000000
0$
0)
#707940000000
1"
1'
b0 +
b0 1
#707990000000
0"
0'
#708000000000
1#
1(
b101111101100100 +
b101111101100100 1
#708050000000
0#
0(
#708060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#708110000000
0$
0)
#708120000000
1"
1'
b0 +
b0 1
#708170000000
0"
0'
#708180000000
1#
1(
b101111101100100 +
b101111101100100 1
#708230000000
0#
0(
#708240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#708290000000
0$
0)
#708300000000
1"
1'
b0 +
b0 1
#708350000000
0"
0'
#708360000000
1#
1(
b101111101100100 +
b101111101100100 1
#708410000000
0#
0(
#708420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#708470000000
0$
0)
#708480000000
1"
1'
b0 +
b0 1
#708530000000
0"
0'
#708540000000
1#
1(
b101111101100100 +
b101111101100100 1
#708590000000
0#
0(
#708600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#708650000000
0$
0)
#708660000000
1"
1'
b0 +
b0 1
#708710000000
0"
0'
#708720000000
1#
1(
b101111101100100 +
b101111101100100 1
#708770000000
0#
0(
#708780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#708830000000
0$
0)
#708840000000
1"
1'
b0 +
b0 1
#708890000000
0"
0'
#708900000000
1#
1(
b101111101100100 +
b101111101100100 1
#708950000000
0#
0(
#708960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#709010000000
0$
0)
#709020000000
1"
1'
b0 +
b0 1
#709070000000
0"
0'
#709080000000
1#
1(
b101111101100100 +
b101111101100100 1
#709130000000
0#
0(
#709140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#709190000000
0$
0)
#709200000000
1"
1'
b0 +
b0 1
#709250000000
0"
0'
#709260000000
1#
1(
b101111101100100 +
b101111101100100 1
#709310000000
0#
0(
#709320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#709370000000
0$
0)
#709380000000
1"
1'
b0 +
b0 1
#709430000000
0"
0'
#709440000000
1#
1(
b101111101100100 +
b101111101100100 1
#709490000000
0#
0(
#709500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#709550000000
0$
0)
#709560000000
1"
1'
b0 +
b0 1
#709610000000
0"
0'
#709620000000
1#
1(
b101111101100100 +
b101111101100100 1
#709670000000
0#
0(
#709680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#709730000000
0$
0)
#709740000000
1"
1'
b0 +
b0 1
#709790000000
0"
0'
#709800000000
1#
1(
b101111101100100 +
b101111101100100 1
#709850000000
0#
0(
#709860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#709910000000
0$
0)
#709920000000
1"
1'
b0 +
b0 1
#709970000000
0"
0'
#709980000000
1#
1(
b101111101100100 +
b101111101100100 1
#710030000000
0#
0(
#710040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#710090000000
0$
0)
#710100000000
1"
1'
b0 +
b0 1
#710150000000
0"
0'
#710160000000
1#
1(
b101111101100100 +
b101111101100100 1
#710210000000
0#
0(
#710220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#710270000000
0$
0)
#710280000000
1"
1'
b0 +
b0 1
#710330000000
0"
0'
#710340000000
1#
1(
b101111101100100 +
b101111101100100 1
#710390000000
0#
0(
#710400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#710450000000
0$
0)
#710460000000
1"
1'
b0 +
b0 1
#710510000000
0"
0'
#710520000000
1#
1(
b101111101100100 +
b101111101100100 1
#710570000000
0#
0(
#710580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#710630000000
0$
0)
#710640000000
1"
1'
b0 +
b0 1
#710690000000
0"
0'
#710700000000
1#
1(
b101111101100100 +
b101111101100100 1
#710750000000
0#
0(
#710760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#710810000000
0$
0)
#710820000000
1"
1'
b0 +
b0 1
#710870000000
0"
0'
#710880000000
1#
1(
b101111101100100 +
b101111101100100 1
#710930000000
0#
0(
#710940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#710990000000
0$
0)
#711000000000
1"
1'
b0 +
b0 1
#711050000000
0"
0'
#711060000000
1#
1(
b101111101100100 +
b101111101100100 1
#711110000000
0#
0(
#711120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#711170000000
0$
0)
#711180000000
1"
1'
b0 +
b0 1
#711230000000
0"
0'
#711240000000
1#
1(
b101111101100100 +
b101111101100100 1
#711290000000
0#
0(
#711300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#711350000000
0$
0)
#711360000000
1"
1'
b0 +
b0 1
#711410000000
0"
0'
#711420000000
1#
1(
b101111101100100 +
b101111101100100 1
#711470000000
0#
0(
#711480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#711530000000
0$
0)
#711540000000
1"
1'
b0 +
b0 1
#711590000000
0"
0'
#711600000000
1#
1(
b101111101100100 +
b101111101100100 1
#711650000000
0#
0(
#711660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#711710000000
0$
0)
#711720000000
1"
1'
b0 +
b0 1
#711770000000
0"
0'
#711780000000
1#
1(
b101111101100100 +
b101111101100100 1
#711830000000
0#
0(
#711840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#711890000000
0$
0)
#711900000000
1"
1'
b0 +
b0 1
#711950000000
0"
0'
#711960000000
1#
1(
b101111101100100 +
b101111101100100 1
#712010000000
0#
0(
#712020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#712070000000
0$
0)
#712080000000
1"
1'
b0 +
b0 1
#712130000000
0"
0'
#712140000000
1#
1(
b101111101100100 +
b101111101100100 1
#712190000000
0#
0(
#712200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#712250000000
0$
0)
#712260000000
1"
1'
b0 +
b0 1
#712310000000
0"
0'
#712320000000
1#
1(
b101111101100100 +
b101111101100100 1
#712370000000
0#
0(
#712380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#712430000000
0$
0)
#712440000000
1"
1'
b0 +
b0 1
#712490000000
0"
0'
#712500000000
1#
1(
b101111101100100 +
b101111101100100 1
#712550000000
0#
0(
#712560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#712610000000
0$
0)
#712620000000
1"
1'
b0 +
b0 1
#712670000000
0"
0'
#712680000000
1#
1(
b101111101100100 +
b101111101100100 1
#712730000000
0#
0(
#712740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#712790000000
0$
0)
#712800000000
1"
1'
b0 +
b0 1
#712850000000
0"
0'
#712860000000
1#
1(
b101111101100100 +
b101111101100100 1
#712910000000
0#
0(
#712920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#712970000000
0$
0)
#712980000000
1"
1'
b0 +
b0 1
#713030000000
0"
0'
#713040000000
1#
1(
b101111101100100 +
b101111101100100 1
#713090000000
0#
0(
#713100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#713150000000
0$
0)
#713160000000
1"
1'
b0 +
b0 1
#713210000000
0"
0'
#713220000000
1#
1(
b101111101100100 +
b101111101100100 1
#713270000000
0#
0(
#713280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#713330000000
0$
0)
#713340000000
1"
1'
b0 +
b0 1
#713390000000
0"
0'
#713400000000
1#
1(
b101111101100100 +
b101111101100100 1
#713450000000
0#
0(
#713460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#713510000000
0$
0)
#713520000000
1"
1'
b0 +
b0 1
#713570000000
0"
0'
#713580000000
1#
1(
b101111101100100 +
b101111101100100 1
#713630000000
0#
0(
#713640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#713690000000
0$
0)
#713700000000
1"
1'
b0 +
b0 1
#713750000000
0"
0'
#713760000000
1#
1(
b101111101100100 +
b101111101100100 1
#713810000000
0#
0(
#713820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#713870000000
0$
0)
#713880000000
1"
1'
b0 +
b0 1
#713930000000
0"
0'
#713940000000
1#
1(
b101111101100100 +
b101111101100100 1
#713990000000
0#
0(
#714000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#714050000000
0$
0)
#714060000000
1"
1'
b0 +
b0 1
#714110000000
0"
0'
#714120000000
1#
1(
b101111101100100 +
b101111101100100 1
#714170000000
0#
0(
#714180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#714230000000
0$
0)
#714240000000
1"
1'
b0 +
b0 1
#714290000000
0"
0'
#714300000000
1#
1(
b101111101100100 +
b101111101100100 1
#714350000000
0#
0(
#714360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#714410000000
0$
0)
#714420000000
1"
1'
b0 +
b0 1
#714470000000
0"
0'
#714480000000
1#
1(
b101111101100100 +
b101111101100100 1
#714530000000
0#
0(
#714540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#714590000000
0$
0)
#714600000000
1"
1'
b0 +
b0 1
#714650000000
0"
0'
#714660000000
1#
1(
b101111101100100 +
b101111101100100 1
#714710000000
0#
0(
#714720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#714770000000
0$
0)
#714780000000
1"
1'
b0 +
b0 1
#714830000000
0"
0'
#714840000000
1#
1(
b101111101100100 +
b101111101100100 1
#714890000000
0#
0(
#714900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#714950000000
0$
0)
#714960000000
1"
1'
b0 +
b0 1
#715010000000
0"
0'
#715020000000
1#
1(
b101111101100100 +
b101111101100100 1
#715070000000
0#
0(
#715080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#715130000000
0$
0)
#715140000000
1"
1'
b0 +
b0 1
#715190000000
0"
0'
#715200000000
1#
1(
b101111101100100 +
b101111101100100 1
#715250000000
0#
0(
#715260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#715310000000
0$
0)
#715320000000
1"
1'
b0 +
b0 1
#715370000000
0"
0'
#715380000000
1#
1(
b101111101100100 +
b101111101100100 1
#715430000000
0#
0(
#715440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#715490000000
0$
0)
#715500000000
1"
1'
b0 +
b0 1
#715550000000
0"
0'
#715560000000
1#
1(
b101111101100100 +
b101111101100100 1
#715610000000
0#
0(
#715620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#715670000000
0$
0)
#715680000000
1"
1'
b0 +
b0 1
#715730000000
0"
0'
#715740000000
1#
1(
b101111101100100 +
b101111101100100 1
#715790000000
0#
0(
#715800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#715850000000
0$
0)
#715860000000
1"
1'
b0 +
b0 1
#715910000000
0"
0'
#715920000000
1#
1(
b101111101100100 +
b101111101100100 1
#715970000000
0#
0(
#715980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#716030000000
0$
0)
#716040000000
1"
1'
b0 +
b0 1
#716090000000
0"
0'
#716100000000
1#
1(
b101111101100100 +
b101111101100100 1
#716150000000
0#
0(
#716160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#716210000000
0$
0)
#716220000000
1"
1'
b0 +
b0 1
#716270000000
0"
0'
#716280000000
1#
1(
b101111101100100 +
b101111101100100 1
#716330000000
0#
0(
#716340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#716390000000
0$
0)
#716400000000
1"
1'
b0 +
b0 1
#716450000000
0"
0'
#716460000000
1#
1(
b101111101100100 +
b101111101100100 1
#716510000000
0#
0(
#716520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#716570000000
0$
0)
#716580000000
1"
1'
b0 +
b0 1
#716630000000
0"
0'
#716640000000
1#
1(
b101111101100100 +
b101111101100100 1
#716690000000
0#
0(
#716700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#716750000000
0$
0)
#716760000000
1"
1'
b0 +
b0 1
#716810000000
0"
0'
#716820000000
1#
1(
b101111101100100 +
b101111101100100 1
#716870000000
0#
0(
#716880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#716930000000
0$
0)
#716940000000
1"
1'
b0 +
b0 1
#716990000000
0"
0'
#717000000000
1#
1(
b101111101100100 +
b101111101100100 1
#717050000000
0#
0(
#717060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#717110000000
0$
0)
#717120000000
1"
1'
b0 +
b0 1
#717170000000
0"
0'
#717180000000
1#
1(
b101111101100100 +
b101111101100100 1
#717230000000
0#
0(
#717240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#717290000000
0$
0)
#717300000000
1"
1'
b0 +
b0 1
#717350000000
0"
0'
#717360000000
1#
1(
b101111101100100 +
b101111101100100 1
#717410000000
0#
0(
#717420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#717470000000
0$
0)
#717480000000
1"
1'
b0 +
b0 1
#717530000000
0"
0'
#717540000000
1#
1(
b101111101100100 +
b101111101100100 1
#717590000000
0#
0(
#717600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#717650000000
0$
0)
#717660000000
1"
1'
b0 +
b0 1
#717710000000
0"
0'
#717720000000
1#
1(
b101111101100100 +
b101111101100100 1
#717770000000
0#
0(
#717780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#717830000000
0$
0)
#717840000000
1"
1'
b0 +
b0 1
#717890000000
0"
0'
#717900000000
1#
1(
b101111101100100 +
b101111101100100 1
#717950000000
0#
0(
#717960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#718010000000
0$
0)
#718020000000
1"
1'
b0 +
b0 1
#718070000000
0"
0'
#718080000000
1#
1(
b101111101100100 +
b101111101100100 1
#718130000000
0#
0(
#718140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#718190000000
0$
0)
#718200000000
1"
1'
b0 +
b0 1
#718250000000
0"
0'
#718260000000
1#
1(
b101111101100100 +
b101111101100100 1
#718310000000
0#
0(
#718320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#718370000000
0$
0)
#718380000000
1"
1'
b0 +
b0 1
#718430000000
0"
0'
#718440000000
1#
1(
b101111101100100 +
b101111101100100 1
#718490000000
0#
0(
#718500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#718550000000
0$
0)
#718560000000
1"
1'
b0 +
b0 1
#718610000000
0"
0'
#718620000000
1#
1(
b101111101100100 +
b101111101100100 1
#718670000000
0#
0(
#718680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#718730000000
0$
0)
#718740000000
1"
1'
b0 +
b0 1
#718790000000
0"
0'
#718800000000
1#
1(
b101111101100100 +
b101111101100100 1
#718850000000
0#
0(
#718860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#718910000000
0$
0)
#718920000000
1"
1'
b0 +
b0 1
#718970000000
0"
0'
#718980000000
1#
1(
b101111101100100 +
b101111101100100 1
#719030000000
0#
0(
#719040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#719090000000
0$
0)
#719100000000
1"
1'
b0 +
b0 1
#719150000000
0"
0'
#719160000000
1#
1(
b101111101100100 +
b101111101100100 1
#719210000000
0#
0(
#719220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#719270000000
0$
0)
#719280000000
1"
1'
b0 +
b0 1
#719330000000
0"
0'
#719340000000
1#
1(
b101111101100100 +
b101111101100100 1
#719390000000
0#
0(
#719400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#719450000000
0$
0)
#719460000000
1"
1'
b0 +
b0 1
#719510000000
0"
0'
#719520000000
1#
1(
b101111101100100 +
b101111101100100 1
#719570000000
0#
0(
#719580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#719630000000
0$
0)
#719640000000
1"
1'
b0 +
b0 1
#719690000000
0"
0'
#719700000000
1#
1(
b101111101100100 +
b101111101100100 1
#719750000000
0#
0(
#719760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#719810000000
0$
0)
#719820000000
1"
1'
b0 +
b0 1
#719870000000
0"
0'
#719880000000
1#
1(
b101111101100100 +
b101111101100100 1
#719930000000
0#
0(
#719940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#719990000000
0$
0)
#720000000000
1"
1'
b0 +
b0 1
#720050000000
0"
0'
#720060000000
1#
1(
b101111101100100 +
b101111101100100 1
#720110000000
0#
0(
#720120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#720170000000
0$
0)
#720180000000
1"
1'
b0 +
b0 1
#720230000000
0"
0'
#720240000000
1#
1(
b101111101100100 +
b101111101100100 1
#720290000000
0#
0(
#720300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#720350000000
0$
0)
#720360000000
1"
1'
b0 +
b0 1
#720410000000
0"
0'
#720420000000
1#
1(
b101111101100100 +
b101111101100100 1
#720470000000
0#
0(
#720480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#720530000000
0$
0)
#720540000000
1"
1'
b0 +
b0 1
#720590000000
0"
0'
#720600000000
1#
1(
b101111101100100 +
b101111101100100 1
#720650000000
0#
0(
#720660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#720710000000
0$
0)
#720720000000
1"
1'
b0 +
b0 1
#720770000000
0"
0'
#720780000000
1#
1(
b101111101100100 +
b101111101100100 1
#720830000000
0#
0(
#720840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#720890000000
0$
0)
#720900000000
1"
1'
b0 +
b0 1
#720950000000
0"
0'
#720960000000
1#
1(
b101111101100100 +
b101111101100100 1
#721010000000
0#
0(
#721020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#721070000000
0$
0)
#721080000000
1"
1'
b0 +
b0 1
#721130000000
0"
0'
#721140000000
1#
1(
b101111101100100 +
b101111101100100 1
#721190000000
0#
0(
#721200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#721250000000
0$
0)
#721260000000
1"
1'
b0 +
b0 1
#721310000000
0"
0'
#721320000000
1#
1(
b101111101100100 +
b101111101100100 1
#721370000000
0#
0(
#721380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#721430000000
0$
0)
#721440000000
1"
1'
b0 +
b0 1
#721490000000
0"
0'
#721500000000
1#
1(
b101111101100100 +
b101111101100100 1
#721550000000
0#
0(
#721560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#721610000000
0$
0)
#721620000000
1"
1'
b0 +
b0 1
#721670000000
0"
0'
#721680000000
1#
1(
b101111101100100 +
b101111101100100 1
#721730000000
0#
0(
#721740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#721790000000
0$
0)
#721800000000
1"
1'
b0 +
b0 1
#721850000000
0"
0'
#721860000000
1#
1(
b101111101100100 +
b101111101100100 1
#721910000000
0#
0(
#721920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#721970000000
0$
0)
#721980000000
1"
1'
b0 +
b0 1
#722030000000
0"
0'
#722040000000
1#
1(
b101111101100100 +
b101111101100100 1
#722090000000
0#
0(
#722100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#722150000000
0$
0)
#722160000000
1"
1'
b0 +
b0 1
#722210000000
0"
0'
#722220000000
1#
1(
b101111101100100 +
b101111101100100 1
#722270000000
0#
0(
#722280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#722330000000
0$
0)
#722340000000
1"
1'
b0 +
b0 1
#722390000000
0"
0'
#722400000000
1#
1(
b101111101100100 +
b101111101100100 1
#722450000000
0#
0(
#722460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#722510000000
0$
0)
#722520000000
1"
1'
b0 +
b0 1
#722570000000
0"
0'
#722580000000
1#
1(
b101111101100100 +
b101111101100100 1
#722630000000
0#
0(
#722640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#722690000000
0$
0)
#722700000000
1"
1'
b0 +
b0 1
#722750000000
0"
0'
#722760000000
1#
1(
b101111101100100 +
b101111101100100 1
#722810000000
0#
0(
#722820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#722870000000
0$
0)
#722880000000
1"
1'
b0 +
b0 1
#722930000000
0"
0'
#722940000000
1#
1(
b101111101100100 +
b101111101100100 1
#722990000000
0#
0(
#723000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#723050000000
0$
0)
#723060000000
1"
1'
b0 +
b0 1
#723110000000
0"
0'
#723120000000
1#
1(
b101111101100100 +
b101111101100100 1
#723170000000
0#
0(
#723180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#723230000000
0$
0)
#723240000000
1"
1'
b0 +
b0 1
#723290000000
0"
0'
#723300000000
1#
1(
b101111101100100 +
b101111101100100 1
#723350000000
0#
0(
#723360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#723410000000
0$
0)
#723420000000
1"
1'
b0 +
b0 1
#723470000000
0"
0'
#723480000000
1#
1(
b101111101100100 +
b101111101100100 1
#723530000000
0#
0(
#723540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#723590000000
0$
0)
#723600000000
1"
1'
b0 +
b0 1
#723650000000
0"
0'
#723660000000
1#
1(
b101111101100100 +
b101111101100100 1
#723710000000
0#
0(
#723720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#723770000000
0$
0)
#723780000000
1"
1'
b0 +
b0 1
#723830000000
0"
0'
#723840000000
1#
1(
b101111101100100 +
b101111101100100 1
#723890000000
0#
0(
#723900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#723950000000
0$
0)
#723960000000
1"
1'
b0 +
b0 1
#724010000000
0"
0'
#724020000000
1#
1(
b101111101100100 +
b101111101100100 1
#724070000000
0#
0(
#724080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#724130000000
0$
0)
#724140000000
1"
1'
b0 +
b0 1
#724190000000
0"
0'
#724200000000
1#
1(
b101111101100100 +
b101111101100100 1
#724250000000
0#
0(
#724260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#724310000000
0$
0)
#724320000000
1"
1'
b0 +
b0 1
#724370000000
0"
0'
#724380000000
1#
1(
b101111101100100 +
b101111101100100 1
#724430000000
0#
0(
#724440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#724490000000
0$
0)
#724500000000
1"
1'
b0 +
b0 1
#724550000000
0"
0'
#724560000000
1#
1(
b101111101100100 +
b101111101100100 1
#724610000000
0#
0(
#724620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#724670000000
0$
0)
#724680000000
1"
1'
b0 +
b0 1
#724730000000
0"
0'
#724740000000
1#
1(
b101111101100100 +
b101111101100100 1
#724790000000
0#
0(
#724800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#724850000000
0$
0)
#724860000000
1"
1'
b0 +
b0 1
#724910000000
0"
0'
#724920000000
1#
1(
b101111101100100 +
b101111101100100 1
#724970000000
0#
0(
#724980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#725030000000
0$
0)
#725040000000
1"
1'
b0 +
b0 1
#725090000000
0"
0'
#725100000000
1#
1(
b101111101100100 +
b101111101100100 1
#725150000000
0#
0(
#725160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#725210000000
0$
0)
#725220000000
1"
1'
b0 +
b0 1
#725270000000
0"
0'
#725280000000
1#
1(
b101111101100100 +
b101111101100100 1
#725330000000
0#
0(
#725340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#725390000000
0$
0)
#725400000000
1"
1'
b0 +
b0 1
#725450000000
0"
0'
#725460000000
1#
1(
b101111101100100 +
b101111101100100 1
#725510000000
0#
0(
#725520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#725570000000
0$
0)
#725580000000
1"
1'
b0 +
b0 1
#725630000000
0"
0'
#725640000000
1#
1(
b101111101100100 +
b101111101100100 1
#725690000000
0#
0(
#725700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#725750000000
0$
0)
#725760000000
1"
1'
b0 +
b0 1
#725810000000
0"
0'
#725820000000
1#
1(
b101111101100100 +
b101111101100100 1
#725870000000
0#
0(
#725880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#725930000000
0$
0)
#725940000000
1"
1'
b0 +
b0 1
#725990000000
0"
0'
#726000000000
1#
1(
b101111101100100 +
b101111101100100 1
#726050000000
0#
0(
#726060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#726110000000
0$
0)
#726120000000
1"
1'
b0 +
b0 1
#726170000000
0"
0'
#726180000000
1#
1(
b101111101100100 +
b101111101100100 1
#726230000000
0#
0(
#726240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#726290000000
0$
0)
#726300000000
1"
1'
b0 +
b0 1
#726350000000
0"
0'
#726360000000
1#
1(
b101111101100100 +
b101111101100100 1
#726410000000
0#
0(
#726420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#726470000000
0$
0)
#726480000000
1"
1'
b0 +
b0 1
#726530000000
0"
0'
#726540000000
1#
1(
b101111101100100 +
b101111101100100 1
#726590000000
0#
0(
#726600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#726650000000
0$
0)
#726660000000
1"
1'
b0 +
b0 1
#726710000000
0"
0'
#726720000000
1#
1(
b101111101100100 +
b101111101100100 1
#726770000000
0#
0(
#726780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#726830000000
0$
0)
#726840000000
1"
1'
b0 +
b0 1
#726890000000
0"
0'
#726900000000
1#
1(
b101111101100100 +
b101111101100100 1
#726950000000
0#
0(
#726960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#727010000000
0$
0)
#727020000000
1"
1'
b0 +
b0 1
#727070000000
0"
0'
#727080000000
1#
1(
b101111101100100 +
b101111101100100 1
#727130000000
0#
0(
#727140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#727190000000
0$
0)
#727200000000
1"
1'
b0 +
b0 1
#727250000000
0"
0'
#727260000000
1#
1(
b101111101100100 +
b101111101100100 1
#727310000000
0#
0(
#727320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#727370000000
0$
0)
#727380000000
1"
1'
b0 +
b0 1
#727430000000
0"
0'
#727440000000
1#
1(
b101111101100100 +
b101111101100100 1
#727490000000
0#
0(
#727500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#727550000000
0$
0)
#727560000000
1"
1'
b0 +
b0 1
#727610000000
0"
0'
#727620000000
1#
1(
b101111101100100 +
b101111101100100 1
#727670000000
0#
0(
#727680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#727730000000
0$
0)
#727740000000
1"
1'
b0 +
b0 1
#727790000000
0"
0'
#727800000000
1#
1(
b101111101100100 +
b101111101100100 1
#727850000000
0#
0(
#727860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#727910000000
0$
0)
#727920000000
1"
1'
b0 +
b0 1
#727970000000
0"
0'
#727980000000
1#
1(
b101111101100100 +
b101111101100100 1
#728030000000
0#
0(
#728040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#728090000000
0$
0)
#728100000000
1"
1'
b0 +
b0 1
#728150000000
0"
0'
#728160000000
1#
1(
b101111101100100 +
b101111101100100 1
#728210000000
0#
0(
#728220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#728270000000
0$
0)
#728280000000
1"
1'
b0 +
b0 1
#728330000000
0"
0'
#728340000000
1#
1(
b101111101100100 +
b101111101100100 1
#728390000000
0#
0(
#728400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#728450000000
0$
0)
#728460000000
1"
1'
b0 +
b0 1
#728510000000
0"
0'
#728520000000
1#
1(
b101111101100100 +
b101111101100100 1
#728570000000
0#
0(
#728580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#728630000000
0$
0)
#728640000000
1"
1'
b0 +
b0 1
#728690000000
0"
0'
#728700000000
1#
1(
b101111101100100 +
b101111101100100 1
#728750000000
0#
0(
#728760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#728810000000
0$
0)
#728820000000
1"
1'
b0 +
b0 1
#728870000000
0"
0'
#728880000000
1#
1(
b101111101100100 +
b101111101100100 1
#728930000000
0#
0(
#728940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#728990000000
0$
0)
#729000000000
1"
1'
b0 +
b0 1
#729050000000
0"
0'
#729060000000
1#
1(
b101111101100100 +
b101111101100100 1
#729110000000
0#
0(
#729120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#729170000000
0$
0)
#729180000000
1"
1'
b0 +
b0 1
#729230000000
0"
0'
#729240000000
1#
1(
b101111101100100 +
b101111101100100 1
#729290000000
0#
0(
#729300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#729350000000
0$
0)
#729360000000
1"
1'
b0 +
b0 1
#729410000000
0"
0'
#729420000000
1#
1(
b101111101100100 +
b101111101100100 1
#729470000000
0#
0(
#729480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#729530000000
0$
0)
#729540000000
1"
1'
b0 +
b0 1
#729590000000
0"
0'
#729600000000
1#
1(
b101111101100100 +
b101111101100100 1
#729650000000
0#
0(
#729660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#729710000000
0$
0)
#729720000000
1"
1'
b0 +
b0 1
#729770000000
0"
0'
#729780000000
1#
1(
b101111101100100 +
b101111101100100 1
#729830000000
0#
0(
#729840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#729890000000
0$
0)
#729900000000
1"
1'
b0 +
b0 1
#729950000000
0"
0'
#729960000000
1#
1(
b101111101100100 +
b101111101100100 1
#730010000000
0#
0(
#730020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#730070000000
0$
0)
#730080000000
1"
1'
b0 +
b0 1
#730130000000
0"
0'
#730140000000
1#
1(
b101111101100100 +
b101111101100100 1
#730190000000
0#
0(
#730200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#730250000000
0$
0)
#730260000000
1"
1'
b0 +
b0 1
#730310000000
0"
0'
#730320000000
1#
1(
b101111101100100 +
b101111101100100 1
#730370000000
0#
0(
#730380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#730430000000
0$
0)
#730440000000
1"
1'
b0 +
b0 1
#730490000000
0"
0'
#730500000000
1#
1(
b101111101100100 +
b101111101100100 1
#730550000000
0#
0(
#730560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#730610000000
0$
0)
#730620000000
1"
1'
b0 +
b0 1
#730670000000
0"
0'
#730680000000
1#
1(
b101111101100100 +
b101111101100100 1
#730730000000
0#
0(
#730740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#730790000000
0$
0)
#730800000000
1"
1'
b0 +
b0 1
#730850000000
0"
0'
#730860000000
1#
1(
b101111101100100 +
b101111101100100 1
#730910000000
0#
0(
#730920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#730970000000
0$
0)
#730980000000
1"
1'
b0 +
b0 1
#731030000000
0"
0'
#731040000000
1#
1(
b101111101100100 +
b101111101100100 1
#731090000000
0#
0(
#731100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#731150000000
0$
0)
#731160000000
1"
1'
b0 +
b0 1
#731210000000
0"
0'
#731220000000
1#
1(
b101111101100100 +
b101111101100100 1
#731270000000
0#
0(
#731280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#731330000000
0$
0)
#731340000000
1"
1'
b0 +
b0 1
#731390000000
0"
0'
#731400000000
1#
1(
b101111101100100 +
b101111101100100 1
#731450000000
0#
0(
#731460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#731510000000
0$
0)
#731520000000
1"
1'
b0 +
b0 1
#731570000000
0"
0'
#731580000000
1#
1(
b101111101100100 +
b101111101100100 1
#731630000000
0#
0(
#731640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#731690000000
0$
0)
#731700000000
1"
1'
b0 +
b0 1
#731750000000
0"
0'
#731760000000
1#
1(
b101111101100100 +
b101111101100100 1
#731810000000
0#
0(
#731820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#731870000000
0$
0)
#731880000000
1"
1'
b0 +
b0 1
#731930000000
0"
0'
#731940000000
1#
1(
b101111101100100 +
b101111101100100 1
#731990000000
0#
0(
#732000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#732050000000
0$
0)
#732060000000
1"
1'
b0 +
b0 1
#732110000000
0"
0'
#732120000000
1#
1(
b101111101100100 +
b101111101100100 1
#732170000000
0#
0(
#732180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#732230000000
0$
0)
#732240000000
1"
1'
b0 +
b0 1
#732290000000
0"
0'
#732300000000
1#
1(
b101111101100100 +
b101111101100100 1
#732350000000
0#
0(
#732360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#732410000000
0$
0)
#732420000000
1"
1'
b0 +
b0 1
#732470000000
0"
0'
#732480000000
1#
1(
b101111101100100 +
b101111101100100 1
#732530000000
0#
0(
#732540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#732590000000
0$
0)
#732600000000
1"
1'
b0 +
b0 1
#732650000000
0"
0'
#732660000000
1#
1(
b101111101100100 +
b101111101100100 1
#732710000000
0#
0(
#732720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#732770000000
0$
0)
#732780000000
1"
1'
b0 +
b0 1
#732830000000
0"
0'
#732840000000
1#
1(
b101111101100100 +
b101111101100100 1
#732890000000
0#
0(
#732900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#732950000000
0$
0)
#732960000000
1"
1'
b0 +
b0 1
#733010000000
0"
0'
#733020000000
1#
1(
b101111101100100 +
b101111101100100 1
#733070000000
0#
0(
#733080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#733130000000
0$
0)
#733140000000
1"
1'
b0 +
b0 1
#733190000000
0"
0'
#733200000000
1#
1(
b101111101100100 +
b101111101100100 1
#733250000000
0#
0(
#733260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#733310000000
0$
0)
#733320000000
1"
1'
b0 +
b0 1
#733370000000
0"
0'
#733380000000
1#
1(
b101111101100100 +
b101111101100100 1
#733430000000
0#
0(
#733440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#733490000000
0$
0)
#733500000000
1"
1'
b0 +
b0 1
#733550000000
0"
0'
#733560000000
1#
1(
b101111101100100 +
b101111101100100 1
#733610000000
0#
0(
#733620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#733670000000
0$
0)
#733680000000
1"
1'
b0 +
b0 1
#733730000000
0"
0'
#733740000000
1#
1(
b101111101100100 +
b101111101100100 1
#733790000000
0#
0(
#733800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#733850000000
0$
0)
#733860000000
1"
1'
b0 +
b0 1
#733910000000
0"
0'
#733920000000
1#
1(
b101111101100100 +
b101111101100100 1
#733970000000
0#
0(
#733980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#734030000000
0$
0)
#734040000000
1"
1'
b0 +
b0 1
#734090000000
0"
0'
#734100000000
1#
1(
b101111101100100 +
b101111101100100 1
#734150000000
0#
0(
#734160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#734210000000
0$
0)
#734220000000
1"
1'
b0 +
b0 1
#734270000000
0"
0'
#734280000000
1#
1(
b101111101100100 +
b101111101100100 1
#734330000000
0#
0(
#734340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#734390000000
0$
0)
#734400000000
1"
1'
b0 +
b0 1
#734450000000
0"
0'
#734460000000
1#
1(
b101111101100100 +
b101111101100100 1
#734510000000
0#
0(
#734520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#734570000000
0$
0)
#734580000000
1"
1'
b0 +
b0 1
#734630000000
0"
0'
#734640000000
1#
1(
b101111101100100 +
b101111101100100 1
#734690000000
0#
0(
#734700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#734750000000
0$
0)
#734760000000
1"
1'
b0 +
b0 1
#734810000000
0"
0'
#734820000000
1#
1(
b101111101100100 +
b101111101100100 1
#734870000000
0#
0(
#734880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#734930000000
0$
0)
#734940000000
1"
1'
b0 +
b0 1
#734990000000
0"
0'
#735000000000
1#
1(
b101111101100100 +
b101111101100100 1
#735050000000
0#
0(
#735060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#735110000000
0$
0)
#735120000000
1"
1'
b0 +
b0 1
#735170000000
0"
0'
#735180000000
1#
1(
b101111101100100 +
b101111101100100 1
#735230000000
0#
0(
#735240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#735290000000
0$
0)
#735300000000
1"
1'
b0 +
b0 1
#735350000000
0"
0'
#735360000000
1#
1(
b101111101100100 +
b101111101100100 1
#735410000000
0#
0(
#735420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#735470000000
0$
0)
#735480000000
1"
1'
b0 +
b0 1
#735530000000
0"
0'
#735540000000
1#
1(
b101111101100100 +
b101111101100100 1
#735590000000
0#
0(
#735600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#735650000000
0$
0)
#735660000000
1"
1'
b0 +
b0 1
#735710000000
0"
0'
#735720000000
1#
1(
b101111101100100 +
b101111101100100 1
#735770000000
0#
0(
#735780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#735830000000
0$
0)
#735840000000
1"
1'
b0 +
b0 1
#735890000000
0"
0'
#735900000000
1#
1(
b101111101100100 +
b101111101100100 1
#735950000000
0#
0(
#735960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#736010000000
0$
0)
#736020000000
1"
1'
b0 +
b0 1
#736070000000
0"
0'
#736080000000
1#
1(
b101111101100100 +
b101111101100100 1
#736130000000
0#
0(
#736140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#736190000000
0$
0)
#736200000000
1"
1'
b0 +
b0 1
#736250000000
0"
0'
#736260000000
1#
1(
b101111101100100 +
b101111101100100 1
#736310000000
0#
0(
#736320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#736370000000
0$
0)
#736380000000
1"
1'
b0 +
b0 1
#736430000000
0"
0'
#736440000000
1#
1(
b101111101100100 +
b101111101100100 1
#736490000000
0#
0(
#736500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#736550000000
0$
0)
#736560000000
1"
1'
b0 +
b0 1
#736610000000
0"
0'
#736620000000
1#
1(
b101111101100100 +
b101111101100100 1
#736670000000
0#
0(
#736680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#736730000000
0$
0)
#736740000000
1"
1'
b0 +
b0 1
#736790000000
0"
0'
#736800000000
1#
1(
b101111101100100 +
b101111101100100 1
#736850000000
0#
0(
#736860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#736910000000
0$
0)
#736920000000
1"
1'
b0 +
b0 1
#736970000000
0"
0'
#736980000000
1#
1(
b101111101100100 +
b101111101100100 1
#737030000000
0#
0(
#737040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#737090000000
0$
0)
#737100000000
1"
1'
b0 +
b0 1
#737150000000
0"
0'
#737160000000
1#
1(
b101111101100100 +
b101111101100100 1
#737210000000
0#
0(
#737220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#737270000000
0$
0)
#737280000000
1"
1'
b0 +
b0 1
#737330000000
0"
0'
#737340000000
1#
1(
b101111101100100 +
b101111101100100 1
#737390000000
0#
0(
#737400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#737450000000
0$
0)
#737460000000
1"
1'
b0 +
b0 1
#737510000000
0"
0'
#737520000000
1#
1(
b101111101100100 +
b101111101100100 1
#737570000000
0#
0(
#737580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#737630000000
0$
0)
#737640000000
1"
1'
b0 +
b0 1
#737690000000
0"
0'
#737700000000
1#
1(
b101111101100100 +
b101111101100100 1
#737750000000
0#
0(
#737760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#737810000000
0$
0)
#737820000000
1"
1'
b0 +
b0 1
#737870000000
0"
0'
#737880000000
1#
1(
b101111101100100 +
b101111101100100 1
#737930000000
0#
0(
#737940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#737990000000
0$
0)
#738000000000
1"
1'
b0 +
b0 1
#738050000000
0"
0'
#738060000000
1#
1(
b101111101100100 +
b101111101100100 1
#738110000000
0#
0(
#738120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#738170000000
0$
0)
#738180000000
1"
1'
b0 +
b0 1
#738230000000
0"
0'
#738240000000
1#
1(
b101111101100100 +
b101111101100100 1
#738290000000
0#
0(
#738300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#738350000000
0$
0)
#738360000000
1"
1'
b0 +
b0 1
#738410000000
0"
0'
#738420000000
1#
1(
b101111101100100 +
b101111101100100 1
#738470000000
0#
0(
#738480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#738530000000
0$
0)
#738540000000
1"
1'
b0 +
b0 1
#738590000000
0"
0'
#738600000000
1#
1(
b101111101100100 +
b101111101100100 1
#738650000000
0#
0(
#738660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#738710000000
0$
0)
#738720000000
1"
1'
b0 +
b0 1
#738770000000
0"
0'
#738780000000
1#
1(
b101111101100100 +
b101111101100100 1
#738830000000
0#
0(
#738840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#738890000000
0$
0)
#738900000000
1"
1'
b0 +
b0 1
#738950000000
0"
0'
#738960000000
1#
1(
b101111101100100 +
b101111101100100 1
#739010000000
0#
0(
#739020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#739070000000
0$
0)
#739080000000
1"
1'
b0 +
b0 1
#739130000000
0"
0'
#739140000000
1#
1(
b101111101100100 +
b101111101100100 1
#739190000000
0#
0(
#739200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#739250000000
0$
0)
#739260000000
1"
1'
b0 +
b0 1
#739310000000
0"
0'
#739320000000
1#
1(
b101111101100100 +
b101111101100100 1
#739370000000
0#
0(
#739380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#739430000000
0$
0)
#739440000000
1"
1'
b0 +
b0 1
#739490000000
0"
0'
#739500000000
1#
1(
b101111101100100 +
b101111101100100 1
#739550000000
0#
0(
#739560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#739610000000
0$
0)
#739620000000
1"
1'
b0 +
b0 1
#739670000000
0"
0'
#739680000000
1#
1(
b101111101100100 +
b101111101100100 1
#739730000000
0#
0(
#739740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#739790000000
0$
0)
#739800000000
1"
1'
b0 +
b0 1
#739850000000
0"
0'
#739860000000
1#
1(
b101111101100100 +
b101111101100100 1
#739910000000
0#
0(
#739920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#739970000000
0$
0)
#739980000000
1"
1'
b0 +
b0 1
#740030000000
0"
0'
#740040000000
1#
1(
b101111101100100 +
b101111101100100 1
#740090000000
0#
0(
#740100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#740150000000
0$
0)
#740160000000
1"
1'
b0 +
b0 1
#740210000000
0"
0'
#740220000000
1#
1(
b101111101100100 +
b101111101100100 1
#740270000000
0#
0(
#740280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#740330000000
0$
0)
#740340000000
1"
1'
b0 +
b0 1
#740390000000
0"
0'
#740400000000
1#
1(
b101111101100100 +
b101111101100100 1
#740450000000
0#
0(
#740460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#740510000000
0$
0)
#740520000000
1"
1'
b0 +
b0 1
#740570000000
0"
0'
#740580000000
1#
1(
b101111101100100 +
b101111101100100 1
#740630000000
0#
0(
#740640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#740690000000
0$
0)
#740700000000
1"
1'
b0 +
b0 1
#740750000000
0"
0'
#740760000000
1#
1(
b101111101100100 +
b101111101100100 1
#740810000000
0#
0(
#740820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#740870000000
0$
0)
#740880000000
1"
1'
b0 +
b0 1
#740930000000
0"
0'
#740940000000
1#
1(
b101111101100100 +
b101111101100100 1
#740990000000
0#
0(
#741000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#741050000000
0$
0)
#741060000000
1"
1'
b0 +
b0 1
#741110000000
0"
0'
#741120000000
1#
1(
b101111101100100 +
b101111101100100 1
#741170000000
0#
0(
#741180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#741230000000
0$
0)
#741240000000
1"
1'
b0 +
b0 1
#741290000000
0"
0'
#741300000000
1#
1(
b101111101100100 +
b101111101100100 1
#741350000000
0#
0(
#741360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#741410000000
0$
0)
#741420000000
1"
1'
b0 +
b0 1
#741470000000
0"
0'
#741480000000
1#
1(
b101111101100100 +
b101111101100100 1
#741530000000
0#
0(
#741540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#741590000000
0$
0)
#741600000000
1"
1'
b0 +
b0 1
#741650000000
0"
0'
#741660000000
1#
1(
b101111101100100 +
b101111101100100 1
#741710000000
0#
0(
#741720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#741770000000
0$
0)
#741780000000
1"
1'
b0 +
b0 1
#741830000000
0"
0'
#741840000000
1#
1(
b101111101100100 +
b101111101100100 1
#741890000000
0#
0(
#741900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#741950000000
0$
0)
#741960000000
1"
1'
b0 +
b0 1
#742010000000
0"
0'
#742020000000
1#
1(
b101111101100100 +
b101111101100100 1
#742070000000
0#
0(
#742080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#742130000000
0$
0)
#742140000000
1"
1'
b0 +
b0 1
#742190000000
0"
0'
#742200000000
1#
1(
b101111101100100 +
b101111101100100 1
#742250000000
0#
0(
#742260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#742310000000
0$
0)
#742320000000
1"
1'
b0 +
b0 1
#742370000000
0"
0'
#742380000000
1#
1(
b101111101100100 +
b101111101100100 1
#742430000000
0#
0(
#742440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#742490000000
0$
0)
#742500000000
1"
1'
b0 +
b0 1
#742550000000
0"
0'
#742560000000
1#
1(
b101111101100100 +
b101111101100100 1
#742610000000
0#
0(
#742620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#742670000000
0$
0)
#742680000000
1"
1'
b0 +
b0 1
#742730000000
0"
0'
#742740000000
1#
1(
b101111101100100 +
b101111101100100 1
#742790000000
0#
0(
#742800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#742850000000
0$
0)
#742860000000
1"
1'
b0 +
b0 1
#742910000000
0"
0'
#742920000000
1#
1(
b101111101100100 +
b101111101100100 1
#742970000000
0#
0(
#742980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#743030000000
0$
0)
#743040000000
1"
1'
b0 +
b0 1
#743090000000
0"
0'
#743100000000
1#
1(
b101111101100100 +
b101111101100100 1
#743150000000
0#
0(
#743160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#743210000000
0$
0)
#743220000000
1"
1'
b0 +
b0 1
#743270000000
0"
0'
#743280000000
1#
1(
b101111101100100 +
b101111101100100 1
#743330000000
0#
0(
#743340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#743390000000
0$
0)
#743400000000
1"
1'
b0 +
b0 1
#743450000000
0"
0'
#743460000000
1#
1(
b101111101100100 +
b101111101100100 1
#743510000000
0#
0(
#743520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#743570000000
0$
0)
#743580000000
1"
1'
b0 +
b0 1
#743630000000
0"
0'
#743640000000
1#
1(
b101111101100100 +
b101111101100100 1
#743690000000
0#
0(
#743700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#743750000000
0$
0)
#743760000000
1"
1'
b0 +
b0 1
#743810000000
0"
0'
#743820000000
1#
1(
b101111101100100 +
b101111101100100 1
#743870000000
0#
0(
#743880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#743930000000
0$
0)
#743940000000
1"
1'
b0 +
b0 1
#743990000000
0"
0'
#744000000000
1#
1(
b101111101100100 +
b101111101100100 1
#744050000000
0#
0(
#744060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#744110000000
0$
0)
#744120000000
1"
1'
b0 +
b0 1
#744170000000
0"
0'
#744180000000
1#
1(
b101111101100100 +
b101111101100100 1
#744230000000
0#
0(
#744240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#744290000000
0$
0)
#744300000000
1"
1'
b0 +
b0 1
#744350000000
0"
0'
#744360000000
1#
1(
b101111101100100 +
b101111101100100 1
#744410000000
0#
0(
#744420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#744470000000
0$
0)
#744480000000
1"
1'
b0 +
b0 1
#744530000000
0"
0'
#744540000000
1#
1(
b101111101100100 +
b101111101100100 1
#744590000000
0#
0(
#744600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#744650000000
0$
0)
#744660000000
1"
1'
b0 +
b0 1
#744710000000
0"
0'
#744720000000
1#
1(
b101111101100100 +
b101111101100100 1
#744770000000
0#
0(
#744780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#744830000000
0$
0)
#744840000000
1"
1'
b0 +
b0 1
#744890000000
0"
0'
#744900000000
1#
1(
b101111101100100 +
b101111101100100 1
#744950000000
0#
0(
#744960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#745010000000
0$
0)
#745020000000
1"
1'
b0 +
b0 1
#745070000000
0"
0'
#745080000000
1#
1(
b101111101100100 +
b101111101100100 1
#745130000000
0#
0(
#745140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#745190000000
0$
0)
#745200000000
1"
1'
b0 +
b0 1
#745250000000
0"
0'
#745260000000
1#
1(
b101111101100100 +
b101111101100100 1
#745310000000
0#
0(
#745320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#745370000000
0$
0)
#745380000000
1"
1'
b0 +
b0 1
#745430000000
0"
0'
#745440000000
1#
1(
b101111101100100 +
b101111101100100 1
#745490000000
0#
0(
#745500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#745550000000
0$
0)
#745560000000
1"
1'
b0 +
b0 1
#745610000000
0"
0'
#745620000000
1#
1(
b101111101100100 +
b101111101100100 1
#745670000000
0#
0(
#745680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#745730000000
0$
0)
#745740000000
1"
1'
b0 +
b0 1
#745790000000
0"
0'
#745800000000
1#
1(
b101111101100100 +
b101111101100100 1
#745850000000
0#
0(
#745860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#745910000000
0$
0)
#745920000000
1"
1'
b0 +
b0 1
#745970000000
0"
0'
#745980000000
1#
1(
b101111101100100 +
b101111101100100 1
#746030000000
0#
0(
#746040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#746090000000
0$
0)
#746100000000
1"
1'
b0 +
b0 1
#746150000000
0"
0'
#746160000000
1#
1(
b101111101100100 +
b101111101100100 1
#746210000000
0#
0(
#746220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#746270000000
0$
0)
#746280000000
1"
1'
b0 +
b0 1
#746330000000
0"
0'
#746340000000
1#
1(
b101111101100100 +
b101111101100100 1
#746390000000
0#
0(
#746400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#746450000000
0$
0)
#746460000000
1"
1'
b0 +
b0 1
#746510000000
0"
0'
#746520000000
1#
1(
b101111101100100 +
b101111101100100 1
#746570000000
0#
0(
#746580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#746630000000
0$
0)
#746640000000
1"
1'
b0 +
b0 1
#746690000000
0"
0'
#746700000000
1#
1(
b101111101100100 +
b101111101100100 1
#746750000000
0#
0(
#746760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#746810000000
0$
0)
#746820000000
1"
1'
b0 +
b0 1
#746870000000
0"
0'
#746880000000
1#
1(
b101111101100100 +
b101111101100100 1
#746930000000
0#
0(
#746940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#746990000000
0$
0)
#747000000000
1"
1'
b0 +
b0 1
#747050000000
0"
0'
#747060000000
1#
1(
b101111101100100 +
b101111101100100 1
#747110000000
0#
0(
#747120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#747170000000
0$
0)
#747180000000
1"
1'
b0 +
b0 1
#747230000000
0"
0'
#747240000000
1#
1(
b101111101100100 +
b101111101100100 1
#747290000000
0#
0(
#747300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#747350000000
0$
0)
#747360000000
1"
1'
b0 +
b0 1
#747410000000
0"
0'
#747420000000
1#
1(
b101111101100100 +
b101111101100100 1
#747470000000
0#
0(
#747480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#747530000000
0$
0)
#747540000000
1"
1'
b0 +
b0 1
#747590000000
0"
0'
#747600000000
1#
1(
b101111101100100 +
b101111101100100 1
#747650000000
0#
0(
#747660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#747710000000
0$
0)
#747720000000
1"
1'
b0 +
b0 1
#747770000000
0"
0'
#747780000000
1#
1(
b101111101100100 +
b101111101100100 1
#747830000000
0#
0(
#747840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#747890000000
0$
0)
#747900000000
1"
1'
b0 +
b0 1
#747950000000
0"
0'
#747960000000
1#
1(
b101111101100100 +
b101111101100100 1
#748010000000
0#
0(
#748020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#748070000000
0$
0)
#748080000000
1"
1'
b0 +
b0 1
#748130000000
0"
0'
#748140000000
1#
1(
b101111101100100 +
b101111101100100 1
#748190000000
0#
0(
#748200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#748250000000
0$
0)
#748260000000
1"
1'
b0 +
b0 1
#748310000000
0"
0'
#748320000000
1#
1(
b101111101100100 +
b101111101100100 1
#748370000000
0#
0(
#748380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#748430000000
0$
0)
#748440000000
1"
1'
b0 +
b0 1
#748490000000
0"
0'
#748500000000
1#
1(
b101111101100100 +
b101111101100100 1
#748550000000
0#
0(
#748560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#748610000000
0$
0)
#748620000000
1"
1'
b0 +
b0 1
#748670000000
0"
0'
#748680000000
1#
1(
b101111101100100 +
b101111101100100 1
#748730000000
0#
0(
#748740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#748790000000
0$
0)
#748800000000
1"
1'
b0 +
b0 1
#748850000000
0"
0'
#748860000000
1#
1(
b101111101100100 +
b101111101100100 1
#748910000000
0#
0(
#748920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#748970000000
0$
0)
#748980000000
1"
1'
b0 +
b0 1
#749030000000
0"
0'
#749040000000
1#
1(
b101111101100100 +
b101111101100100 1
#749090000000
0#
0(
#749100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#749150000000
0$
0)
#749160000000
1"
1'
b0 +
b0 1
#749210000000
0"
0'
#749220000000
1#
1(
b101111101100100 +
b101111101100100 1
#749270000000
0#
0(
#749280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#749330000000
0$
0)
#749340000000
1"
1'
b0 +
b0 1
#749390000000
0"
0'
#749400000000
1#
1(
b101111101100100 +
b101111101100100 1
#749450000000
0#
0(
#749460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#749510000000
0$
0)
#749520000000
1"
1'
b0 +
b0 1
#749570000000
0"
0'
#749580000000
1#
1(
b101111101100100 +
b101111101100100 1
#749630000000
0#
0(
#749640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#749690000000
0$
0)
#749700000000
1"
1'
b0 +
b0 1
#749750000000
0"
0'
#749760000000
1#
1(
b101111101100100 +
b101111101100100 1
#749810000000
0#
0(
#749820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#749870000000
0$
0)
#749880000000
1"
1'
b0 +
b0 1
#749930000000
0"
0'
#749940000000
1#
1(
b101111101100100 +
b101111101100100 1
#749990000000
0#
0(
#750000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#750050000000
0$
0)
#750060000000
1"
1'
b0 +
b0 1
#750110000000
0"
0'
#750120000000
1#
1(
b101111101100100 +
b101111101100100 1
#750170000000
0#
0(
#750180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#750230000000
0$
0)
#750240000000
1"
1'
b0 +
b0 1
#750290000000
0"
0'
#750300000000
1#
1(
b101111101100100 +
b101111101100100 1
#750350000000
0#
0(
#750360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#750410000000
0$
0)
#750420000000
1"
1'
b0 +
b0 1
#750470000000
0"
0'
#750480000000
1#
1(
b101111101100100 +
b101111101100100 1
#750530000000
0#
0(
#750540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#750590000000
0$
0)
#750600000000
1"
1'
b0 +
b0 1
#750650000000
0"
0'
#750660000000
1#
1(
b101111101100100 +
b101111101100100 1
#750710000000
0#
0(
#750720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#750770000000
0$
0)
#750780000000
1"
1'
b0 +
b0 1
#750830000000
0"
0'
#750840000000
1#
1(
b101111101100100 +
b101111101100100 1
#750890000000
0#
0(
#750900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#750950000000
0$
0)
#750960000000
1"
1'
b0 +
b0 1
#751010000000
0"
0'
#751020000000
1#
1(
b101111101100100 +
b101111101100100 1
#751070000000
0#
0(
#751080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#751130000000
0$
0)
#751140000000
1"
1'
b0 +
b0 1
#751190000000
0"
0'
#751200000000
1#
1(
b101111101100100 +
b101111101100100 1
#751250000000
0#
0(
#751260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#751310000000
0$
0)
#751320000000
1"
1'
b0 +
b0 1
#751370000000
0"
0'
#751380000000
1#
1(
b101111101100100 +
b101111101100100 1
#751430000000
0#
0(
#751440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#751490000000
0$
0)
#751500000000
1"
1'
b0 +
b0 1
#751550000000
0"
0'
#751560000000
1#
1(
b101111101100100 +
b101111101100100 1
#751610000000
0#
0(
#751620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#751670000000
0$
0)
#751680000000
1"
1'
b0 +
b0 1
#751730000000
0"
0'
#751740000000
1#
1(
b101111101100100 +
b101111101100100 1
#751790000000
0#
0(
#751800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#751850000000
0$
0)
#751860000000
1"
1'
b0 +
b0 1
#751910000000
0"
0'
#751920000000
1#
1(
b101111101100100 +
b101111101100100 1
#751970000000
0#
0(
#751980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#752030000000
0$
0)
#752040000000
1"
1'
b0 +
b0 1
#752090000000
0"
0'
#752100000000
1#
1(
b101111101100100 +
b101111101100100 1
#752150000000
0#
0(
#752160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#752210000000
0$
0)
#752220000000
1"
1'
b0 +
b0 1
#752270000000
0"
0'
#752280000000
1#
1(
b101111101100100 +
b101111101100100 1
#752330000000
0#
0(
#752340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#752390000000
0$
0)
#752400000000
1"
1'
b0 +
b0 1
#752450000000
0"
0'
#752460000000
1#
1(
b101111101100100 +
b101111101100100 1
#752510000000
0#
0(
#752520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#752570000000
0$
0)
#752580000000
1"
1'
b0 +
b0 1
#752630000000
0"
0'
#752640000000
1#
1(
b101111101100100 +
b101111101100100 1
#752690000000
0#
0(
#752700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#752750000000
0$
0)
#752760000000
1"
1'
b0 +
b0 1
#752810000000
0"
0'
#752820000000
1#
1(
b101111101100100 +
b101111101100100 1
#752870000000
0#
0(
#752880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#752930000000
0$
0)
#752940000000
1"
1'
b0 +
b0 1
#752990000000
0"
0'
#753000000000
1#
1(
b101111101100100 +
b101111101100100 1
#753050000000
0#
0(
#753060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#753110000000
0$
0)
#753120000000
1"
1'
b0 +
b0 1
#753170000000
0"
0'
#753180000000
1#
1(
b101111101100100 +
b101111101100100 1
#753230000000
0#
0(
#753240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#753290000000
0$
0)
#753300000000
1"
1'
b0 +
b0 1
#753350000000
0"
0'
#753360000000
1#
1(
b101111101100100 +
b101111101100100 1
#753410000000
0#
0(
#753420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#753470000000
0$
0)
#753480000000
1"
1'
b0 +
b0 1
#753530000000
0"
0'
#753540000000
1#
1(
b101111101100100 +
b101111101100100 1
#753590000000
0#
0(
#753600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#753650000000
0$
0)
#753660000000
1"
1'
b0 +
b0 1
#753710000000
0"
0'
#753720000000
1#
1(
b101111101100100 +
b101111101100100 1
#753770000000
0#
0(
#753780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#753830000000
0$
0)
#753840000000
1"
1'
b0 +
b0 1
#753890000000
0"
0'
#753900000000
1#
1(
b101111101100100 +
b101111101100100 1
#753950000000
0#
0(
#753960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#754010000000
0$
0)
#754020000000
1"
1'
b0 +
b0 1
#754070000000
0"
0'
#754080000000
1#
1(
b101111101100100 +
b101111101100100 1
#754130000000
0#
0(
#754140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#754190000000
0$
0)
#754200000000
1"
1'
b0 +
b0 1
#754250000000
0"
0'
#754260000000
1#
1(
b101111101100100 +
b101111101100100 1
#754310000000
0#
0(
#754320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#754370000000
0$
0)
#754380000000
1"
1'
b0 +
b0 1
#754430000000
0"
0'
#754440000000
1#
1(
b101111101100100 +
b101111101100100 1
#754490000000
0#
0(
#754500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#754550000000
0$
0)
#754560000000
1"
1'
b0 +
b0 1
#754610000000
0"
0'
#754620000000
1#
1(
b101111101100100 +
b101111101100100 1
#754670000000
0#
0(
#754680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#754730000000
0$
0)
#754740000000
1"
1'
b0 +
b0 1
#754790000000
0"
0'
#754800000000
1#
1(
b101111101100100 +
b101111101100100 1
#754850000000
0#
0(
#754860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#754910000000
0$
0)
#754920000000
1"
1'
b0 +
b0 1
#754970000000
0"
0'
#754980000000
1#
1(
b101111101100100 +
b101111101100100 1
#755030000000
0#
0(
#755040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#755090000000
0$
0)
#755100000000
1"
1'
b0 +
b0 1
#755150000000
0"
0'
#755160000000
1#
1(
b101111101100100 +
b101111101100100 1
#755210000000
0#
0(
#755220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#755270000000
0$
0)
#755280000000
1"
1'
b0 +
b0 1
#755330000000
0"
0'
#755340000000
1#
1(
b101111101100100 +
b101111101100100 1
#755390000000
0#
0(
#755400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#755450000000
0$
0)
#755460000000
1"
1'
b0 +
b0 1
#755510000000
0"
0'
#755520000000
1#
1(
b101111101100100 +
b101111101100100 1
#755570000000
0#
0(
#755580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#755630000000
0$
0)
#755640000000
1"
1'
b0 +
b0 1
#755690000000
0"
0'
#755700000000
1#
1(
b101111101100100 +
b101111101100100 1
#755750000000
0#
0(
#755760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#755810000000
0$
0)
#755820000000
1"
1'
b0 +
b0 1
#755870000000
0"
0'
#755880000000
1#
1(
b101111101100100 +
b101111101100100 1
#755930000000
0#
0(
#755940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#755990000000
0$
0)
#756000000000
1"
1'
b0 +
b0 1
#756050000000
0"
0'
#756060000000
1#
1(
b101111101100100 +
b101111101100100 1
#756110000000
0#
0(
#756120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#756170000000
0$
0)
#756180000000
1"
1'
b0 +
b0 1
#756230000000
0"
0'
#756240000000
1#
1(
b101111101100100 +
b101111101100100 1
#756290000000
0#
0(
#756300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#756350000000
0$
0)
#756360000000
1"
1'
b0 +
b0 1
#756410000000
0"
0'
#756420000000
1#
1(
b101111101100100 +
b101111101100100 1
#756470000000
0#
0(
#756480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#756530000000
0$
0)
#756540000000
1"
1'
b0 +
b0 1
#756590000000
0"
0'
#756600000000
1#
1(
b101111101100100 +
b101111101100100 1
#756650000000
0#
0(
#756660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#756710000000
0$
0)
#756720000000
1"
1'
b0 +
b0 1
#756770000000
0"
0'
#756780000000
1#
1(
b101111101100100 +
b101111101100100 1
#756830000000
0#
0(
#756840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#756890000000
0$
0)
#756900000000
1"
1'
b0 +
b0 1
#756950000000
0"
0'
#756960000000
1#
1(
b101111101100100 +
b101111101100100 1
#757010000000
0#
0(
#757020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#757070000000
0$
0)
#757080000000
1"
1'
b0 +
b0 1
#757130000000
0"
0'
#757140000000
1#
1(
b101111101100100 +
b101111101100100 1
#757190000000
0#
0(
#757200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#757250000000
0$
0)
#757260000000
1"
1'
b0 +
b0 1
#757310000000
0"
0'
#757320000000
1#
1(
b101111101100100 +
b101111101100100 1
#757370000000
0#
0(
#757380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#757430000000
0$
0)
#757440000000
1"
1'
b0 +
b0 1
#757490000000
0"
0'
#757500000000
1#
1(
b101111101100100 +
b101111101100100 1
#757550000000
0#
0(
#757560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#757610000000
0$
0)
#757620000000
1"
1'
b0 +
b0 1
#757670000000
0"
0'
#757680000000
1#
1(
b101111101100100 +
b101111101100100 1
#757730000000
0#
0(
#757740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#757790000000
0$
0)
#757800000000
1"
1'
b0 +
b0 1
#757850000000
0"
0'
#757860000000
1#
1(
b101111101100100 +
b101111101100100 1
#757910000000
0#
0(
#757920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#757970000000
0$
0)
#757980000000
1"
1'
b0 +
b0 1
#758030000000
0"
0'
#758040000000
1#
1(
b101111101100100 +
b101111101100100 1
#758090000000
0#
0(
#758100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#758150000000
0$
0)
#758160000000
1"
1'
b0 +
b0 1
#758210000000
0"
0'
#758220000000
1#
1(
b101111101100100 +
b101111101100100 1
#758270000000
0#
0(
#758280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#758330000000
0$
0)
#758340000000
1"
1'
b0 +
b0 1
#758390000000
0"
0'
#758400000000
1#
1(
b101111101100100 +
b101111101100100 1
#758450000000
0#
0(
#758460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#758510000000
0$
0)
#758520000000
1"
1'
b0 +
b0 1
#758570000000
0"
0'
#758580000000
1#
1(
b101111101100100 +
b101111101100100 1
#758630000000
0#
0(
#758640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#758690000000
0$
0)
#758700000000
1"
1'
b0 +
b0 1
#758750000000
0"
0'
#758760000000
1#
1(
b101111101100100 +
b101111101100100 1
#758810000000
0#
0(
#758820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#758870000000
0$
0)
#758880000000
1"
1'
b0 +
b0 1
#758930000000
0"
0'
#758940000000
1#
1(
b101111101100100 +
b101111101100100 1
#758990000000
0#
0(
#759000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#759050000000
0$
0)
#759060000000
1"
1'
b0 +
b0 1
#759110000000
0"
0'
#759120000000
1#
1(
b101111101100100 +
b101111101100100 1
#759170000000
0#
0(
#759180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#759230000000
0$
0)
#759240000000
1"
1'
b0 +
b0 1
#759290000000
0"
0'
#759300000000
1#
1(
b101111101100100 +
b101111101100100 1
#759350000000
0#
0(
#759360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#759410000000
0$
0)
#759420000000
1"
1'
b0 +
b0 1
#759470000000
0"
0'
#759480000000
1#
1(
b101111101100100 +
b101111101100100 1
#759530000000
0#
0(
#759540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#759590000000
0$
0)
#759600000000
1"
1'
b0 +
b0 1
#759650000000
0"
0'
#759660000000
1#
1(
b101111101100100 +
b101111101100100 1
#759710000000
0#
0(
#759720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#759770000000
0$
0)
#759780000000
1"
1'
b0 +
b0 1
#759830000000
0"
0'
#759840000000
1#
1(
b101111101100100 +
b101111101100100 1
#759890000000
0#
0(
#759900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#759950000000
0$
0)
#759960000000
1"
1'
b0 +
b0 1
#760010000000
0"
0'
#760020000000
1#
1(
b101111101100100 +
b101111101100100 1
#760070000000
0#
0(
#760080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#760130000000
0$
0)
#760140000000
1"
1'
b0 +
b0 1
#760190000000
0"
0'
#760200000000
1#
1(
b101111101100100 +
b101111101100100 1
#760250000000
0#
0(
#760260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#760310000000
0$
0)
#760320000000
1"
1'
b0 +
b0 1
#760370000000
0"
0'
#760380000000
1#
1(
b101111101100100 +
b101111101100100 1
#760430000000
0#
0(
#760440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#760490000000
0$
0)
#760500000000
1"
1'
b0 +
b0 1
#760550000000
0"
0'
#760560000000
1#
1(
b101111101100100 +
b101111101100100 1
#760610000000
0#
0(
#760620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#760670000000
0$
0)
#760680000000
1"
1'
b0 +
b0 1
#760730000000
0"
0'
#760740000000
1#
1(
b101111101100100 +
b101111101100100 1
#760790000000
0#
0(
#760800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#760850000000
0$
0)
#760860000000
1"
1'
b0 +
b0 1
#760910000000
0"
0'
#760920000000
1#
1(
b101111101100100 +
b101111101100100 1
#760970000000
0#
0(
#760980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#761030000000
0$
0)
#761040000000
1"
1'
b0 +
b0 1
#761090000000
0"
0'
#761100000000
1#
1(
b101111101100100 +
b101111101100100 1
#761150000000
0#
0(
#761160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#761210000000
0$
0)
#761220000000
1"
1'
b0 +
b0 1
#761270000000
0"
0'
#761280000000
1#
1(
b101111101100100 +
b101111101100100 1
#761330000000
0#
0(
#761340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#761390000000
0$
0)
#761400000000
1"
1'
b0 +
b0 1
#761450000000
0"
0'
#761460000000
1#
1(
b101111101100100 +
b101111101100100 1
#761510000000
0#
0(
#761520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#761570000000
0$
0)
#761580000000
1"
1'
b0 +
b0 1
#761630000000
0"
0'
#761640000000
1#
1(
b101111101100100 +
b101111101100100 1
#761690000000
0#
0(
#761700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#761750000000
0$
0)
#761760000000
1"
1'
b0 +
b0 1
#761810000000
0"
0'
#761820000000
1#
1(
b101111101100100 +
b101111101100100 1
#761870000000
0#
0(
#761880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#761930000000
0$
0)
#761940000000
1"
1'
b0 +
b0 1
#761990000000
0"
0'
#762000000000
1#
1(
b101111101100100 +
b101111101100100 1
#762050000000
0#
0(
#762060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#762110000000
0$
0)
#762120000000
1"
1'
b0 +
b0 1
#762170000000
0"
0'
#762180000000
1#
1(
b101111101100100 +
b101111101100100 1
#762230000000
0#
0(
#762240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#762290000000
0$
0)
#762300000000
1"
1'
b0 +
b0 1
#762350000000
0"
0'
#762360000000
1#
1(
b101111101100100 +
b101111101100100 1
#762410000000
0#
0(
#762420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#762470000000
0$
0)
#762480000000
1"
1'
b0 +
b0 1
#762530000000
0"
0'
#762540000000
1#
1(
b101111101100100 +
b101111101100100 1
#762590000000
0#
0(
#762600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#762650000000
0$
0)
#762660000000
1"
1'
b0 +
b0 1
#762710000000
0"
0'
#762720000000
1#
1(
b101111101100100 +
b101111101100100 1
#762770000000
0#
0(
#762780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#762830000000
0$
0)
#762840000000
1"
1'
b0 +
b0 1
#762890000000
0"
0'
#762900000000
1#
1(
b101111101100100 +
b101111101100100 1
#762950000000
0#
0(
#762960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#763010000000
0$
0)
#763020000000
1"
1'
b0 +
b0 1
#763070000000
0"
0'
#763080000000
1#
1(
b101111101100100 +
b101111101100100 1
#763130000000
0#
0(
#763140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#763190000000
0$
0)
#763200000000
1"
1'
b0 +
b0 1
#763250000000
0"
0'
#763260000000
1#
1(
b101111101100100 +
b101111101100100 1
#763310000000
0#
0(
#763320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#763370000000
0$
0)
#763380000000
1"
1'
b0 +
b0 1
#763430000000
0"
0'
#763440000000
1#
1(
b101111101100100 +
b101111101100100 1
#763490000000
0#
0(
#763500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#763550000000
0$
0)
#763560000000
1"
1'
b0 +
b0 1
#763610000000
0"
0'
#763620000000
1#
1(
b101111101100100 +
b101111101100100 1
#763670000000
0#
0(
#763680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#763730000000
0$
0)
#763740000000
1"
1'
b0 +
b0 1
#763790000000
0"
0'
#763800000000
1#
1(
b101111101100100 +
b101111101100100 1
#763850000000
0#
0(
#763860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#763910000000
0$
0)
#763920000000
1"
1'
b0 +
b0 1
#763970000000
0"
0'
#763980000000
1#
1(
b101111101100100 +
b101111101100100 1
#764030000000
0#
0(
#764040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#764090000000
0$
0)
#764100000000
1"
1'
b0 +
b0 1
#764150000000
0"
0'
#764160000000
1#
1(
b101111101100100 +
b101111101100100 1
#764210000000
0#
0(
#764220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#764270000000
0$
0)
#764280000000
1"
1'
b0 +
b0 1
#764330000000
0"
0'
#764340000000
1#
1(
b101111101100100 +
b101111101100100 1
#764390000000
0#
0(
#764400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#764450000000
0$
0)
#764460000000
1"
1'
b0 +
b0 1
#764510000000
0"
0'
#764520000000
1#
1(
b101111101100100 +
b101111101100100 1
#764570000000
0#
0(
#764580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#764630000000
0$
0)
#764640000000
1"
1'
b0 +
b0 1
#764690000000
0"
0'
#764700000000
1#
1(
b101111101100100 +
b101111101100100 1
#764750000000
0#
0(
#764760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#764810000000
0$
0)
#764820000000
1"
1'
b0 +
b0 1
#764870000000
0"
0'
#764880000000
1#
1(
b101111101100100 +
b101111101100100 1
#764930000000
0#
0(
#764940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#764990000000
0$
0)
#765000000000
1"
1'
b0 +
b0 1
#765050000000
0"
0'
#765060000000
1#
1(
b101111101100100 +
b101111101100100 1
#765110000000
0#
0(
#765120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#765170000000
0$
0)
#765180000000
1"
1'
b0 +
b0 1
#765230000000
0"
0'
#765240000000
1#
1(
b101111101100100 +
b101111101100100 1
#765290000000
0#
0(
#765300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#765350000000
0$
0)
#765360000000
1"
1'
b0 +
b0 1
#765410000000
0"
0'
#765420000000
1#
1(
b101111101100100 +
b101111101100100 1
#765470000000
0#
0(
#765480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#765530000000
0$
0)
#765540000000
1"
1'
b0 +
b0 1
#765590000000
0"
0'
#765600000000
1#
1(
b101111101100100 +
b101111101100100 1
#765650000000
0#
0(
#765660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#765710000000
0$
0)
#765720000000
1"
1'
b0 +
b0 1
#765770000000
0"
0'
#765780000000
1#
1(
b101111101100100 +
b101111101100100 1
#765830000000
0#
0(
#765840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#765890000000
0$
0)
#765900000000
1"
1'
b0 +
b0 1
#765950000000
0"
0'
#765960000000
1#
1(
b101111101100100 +
b101111101100100 1
#766010000000
0#
0(
#766020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#766070000000
0$
0)
#766080000000
1"
1'
b0 +
b0 1
#766130000000
0"
0'
#766140000000
1#
1(
b101111101100100 +
b101111101100100 1
#766190000000
0#
0(
#766200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#766250000000
0$
0)
#766260000000
1"
1'
b0 +
b0 1
#766310000000
0"
0'
#766320000000
1#
1(
b101111101100100 +
b101111101100100 1
#766370000000
0#
0(
#766380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#766430000000
0$
0)
#766440000000
1"
1'
b0 +
b0 1
#766490000000
0"
0'
#766500000000
1#
1(
b101111101100100 +
b101111101100100 1
#766550000000
0#
0(
#766560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#766610000000
0$
0)
#766620000000
1"
1'
b0 +
b0 1
#766670000000
0"
0'
#766680000000
1#
1(
b101111101100100 +
b101111101100100 1
#766730000000
0#
0(
#766740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#766790000000
0$
0)
#766800000000
1"
1'
b0 +
b0 1
#766850000000
0"
0'
#766860000000
1#
1(
b101111101100100 +
b101111101100100 1
#766910000000
0#
0(
#766920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#766970000000
0$
0)
#766980000000
1"
1'
b0 +
b0 1
#767030000000
0"
0'
#767040000000
1#
1(
b101111101100100 +
b101111101100100 1
#767090000000
0#
0(
#767100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#767150000000
0$
0)
#767160000000
1"
1'
b0 +
b0 1
#767210000000
0"
0'
#767220000000
1#
1(
b101111101100100 +
b101111101100100 1
#767270000000
0#
0(
#767280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#767330000000
0$
0)
#767340000000
1"
1'
b0 +
b0 1
#767390000000
0"
0'
#767400000000
1#
1(
b101111101100100 +
b101111101100100 1
#767450000000
0#
0(
#767460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#767510000000
0$
0)
#767520000000
1"
1'
b0 +
b0 1
#767570000000
0"
0'
#767580000000
1#
1(
b101111101100100 +
b101111101100100 1
#767630000000
0#
0(
#767640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#767690000000
0$
0)
#767700000000
1"
1'
b0 +
b0 1
#767750000000
0"
0'
#767760000000
1#
1(
b101111101100100 +
b101111101100100 1
#767810000000
0#
0(
#767820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#767870000000
0$
0)
#767880000000
1"
1'
b0 +
b0 1
#767930000000
0"
0'
#767940000000
1#
1(
b101111101100100 +
b101111101100100 1
#767990000000
0#
0(
#768000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#768050000000
0$
0)
#768060000000
1"
1'
b0 +
b0 1
#768110000000
0"
0'
#768120000000
1#
1(
b101111101100100 +
b101111101100100 1
#768170000000
0#
0(
#768180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#768230000000
0$
0)
#768240000000
1"
1'
b0 +
b0 1
#768290000000
0"
0'
#768300000000
1#
1(
b101111101100100 +
b101111101100100 1
#768350000000
0#
0(
#768360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#768410000000
0$
0)
#768420000000
1"
1'
b0 +
b0 1
#768470000000
0"
0'
#768480000000
1#
1(
b101111101100100 +
b101111101100100 1
#768530000000
0#
0(
#768540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#768590000000
0$
0)
#768600000000
1"
1'
b0 +
b0 1
#768650000000
0"
0'
#768660000000
1#
1(
b101111101100100 +
b101111101100100 1
#768710000000
0#
0(
#768720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#768770000000
0$
0)
#768780000000
1"
1'
b0 +
b0 1
#768830000000
0"
0'
#768840000000
1#
1(
b101111101100100 +
b101111101100100 1
#768890000000
0#
0(
#768900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#768950000000
0$
0)
#768960000000
1"
1'
b0 +
b0 1
#769010000000
0"
0'
#769020000000
1#
1(
b101111101100100 +
b101111101100100 1
#769070000000
0#
0(
#769080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#769130000000
0$
0)
#769140000000
1"
1'
b0 +
b0 1
#769190000000
0"
0'
#769200000000
1#
1(
b101111101100100 +
b101111101100100 1
#769250000000
0#
0(
#769260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#769310000000
0$
0)
#769320000000
1"
1'
b0 +
b0 1
#769370000000
0"
0'
#769380000000
1#
1(
b101111101100100 +
b101111101100100 1
#769430000000
0#
0(
#769440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#769490000000
0$
0)
#769500000000
1"
1'
b0 +
b0 1
#769550000000
0"
0'
#769560000000
1#
1(
b101111101100100 +
b101111101100100 1
#769610000000
0#
0(
#769620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#769670000000
0$
0)
#769680000000
1"
1'
b0 +
b0 1
#769730000000
0"
0'
#769740000000
1#
1(
b101111101100100 +
b101111101100100 1
#769790000000
0#
0(
#769800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#769850000000
0$
0)
#769860000000
1"
1'
b0 +
b0 1
#769910000000
0"
0'
#769920000000
1#
1(
b101111101100100 +
b101111101100100 1
#769970000000
0#
0(
#769980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#770030000000
0$
0)
#770040000000
1"
1'
b0 +
b0 1
#770090000000
0"
0'
#770100000000
1#
1(
b101111101100100 +
b101111101100100 1
#770150000000
0#
0(
#770160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#770210000000
0$
0)
#770220000000
1"
1'
b0 +
b0 1
#770270000000
0"
0'
#770280000000
1#
1(
b101111101100100 +
b101111101100100 1
#770330000000
0#
0(
#770340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#770390000000
0$
0)
#770400000000
1"
1'
b0 +
b0 1
#770450000000
0"
0'
#770460000000
1#
1(
b101111101100100 +
b101111101100100 1
#770510000000
0#
0(
#770520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#770570000000
0$
0)
#770580000000
1"
1'
b0 +
b0 1
#770630000000
0"
0'
#770640000000
1#
1(
b101111101100100 +
b101111101100100 1
#770690000000
0#
0(
#770700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#770750000000
0$
0)
#770760000000
1"
1'
b0 +
b0 1
#770810000000
0"
0'
#770820000000
1#
1(
b101111101100100 +
b101111101100100 1
#770870000000
0#
0(
#770880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#770930000000
0$
0)
#770940000000
1"
1'
b0 +
b0 1
#770990000000
0"
0'
#771000000000
1#
1(
b101111101100100 +
b101111101100100 1
#771050000000
0#
0(
#771060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#771110000000
0$
0)
#771120000000
1"
1'
b0 +
b0 1
#771170000000
0"
0'
#771180000000
1#
1(
b101111101100100 +
b101111101100100 1
#771230000000
0#
0(
#771240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#771290000000
0$
0)
#771300000000
1"
1'
b0 +
b0 1
#771350000000
0"
0'
#771360000000
1#
1(
b101111101100100 +
b101111101100100 1
#771410000000
0#
0(
#771420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#771470000000
0$
0)
#771480000000
1"
1'
b0 +
b0 1
#771530000000
0"
0'
#771540000000
1#
1(
b101111101100100 +
b101111101100100 1
#771590000000
0#
0(
#771600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#771650000000
0$
0)
#771660000000
1"
1'
b0 +
b0 1
#771710000000
0"
0'
#771720000000
1#
1(
b101111101100100 +
b101111101100100 1
#771770000000
0#
0(
#771780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#771830000000
0$
0)
#771840000000
1"
1'
b0 +
b0 1
#771890000000
0"
0'
#771900000000
1#
1(
b101111101100100 +
b101111101100100 1
#771950000000
0#
0(
#771960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#772010000000
0$
0)
#772020000000
1"
1'
b0 +
b0 1
#772070000000
0"
0'
#772080000000
1#
1(
b101111101100100 +
b101111101100100 1
#772130000000
0#
0(
#772140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#772190000000
0$
0)
#772200000000
1"
1'
b0 +
b0 1
#772250000000
0"
0'
#772260000000
1#
1(
b101111101100100 +
b101111101100100 1
#772310000000
0#
0(
#772320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#772370000000
0$
0)
#772380000000
1"
1'
b0 +
b0 1
#772430000000
0"
0'
#772440000000
1#
1(
b101111101100100 +
b101111101100100 1
#772490000000
0#
0(
#772500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#772550000000
0$
0)
#772560000000
1"
1'
b0 +
b0 1
#772610000000
0"
0'
#772620000000
1#
1(
b101111101100100 +
b101111101100100 1
#772670000000
0#
0(
#772680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#772730000000
0$
0)
#772740000000
1"
1'
b0 +
b0 1
#772790000000
0"
0'
#772800000000
1#
1(
b101111101100100 +
b101111101100100 1
#772850000000
0#
0(
#772860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#772910000000
0$
0)
#772920000000
1"
1'
b0 +
b0 1
#772970000000
0"
0'
#772980000000
1#
1(
b101111101100100 +
b101111101100100 1
#773030000000
0#
0(
#773040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#773090000000
0$
0)
#773100000000
1"
1'
b0 +
b0 1
#773150000000
0"
0'
#773160000000
1#
1(
b101111101100100 +
b101111101100100 1
#773210000000
0#
0(
#773220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#773270000000
0$
0)
#773280000000
1"
1'
b0 +
b0 1
#773330000000
0"
0'
#773340000000
1#
1(
b101111101100100 +
b101111101100100 1
#773390000000
0#
0(
#773400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#773450000000
0$
0)
#773460000000
1"
1'
b0 +
b0 1
#773510000000
0"
0'
#773520000000
1#
1(
b101111101100100 +
b101111101100100 1
#773570000000
0#
0(
#773580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#773630000000
0$
0)
#773640000000
1"
1'
b0 +
b0 1
#773690000000
0"
0'
#773700000000
1#
1(
b101111101100100 +
b101111101100100 1
#773750000000
0#
0(
#773760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#773810000000
0$
0)
#773820000000
1"
1'
b0 +
b0 1
#773870000000
0"
0'
#773880000000
1#
1(
b101111101100100 +
b101111101100100 1
#773930000000
0#
0(
#773940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#773990000000
0$
0)
#774000000000
1"
1'
b0 +
b0 1
#774050000000
0"
0'
#774060000000
1#
1(
b101111101100100 +
b101111101100100 1
#774110000000
0#
0(
#774120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#774170000000
0$
0)
#774180000000
1"
1'
b0 +
b0 1
#774230000000
0"
0'
#774240000000
1#
1(
b101111101100100 +
b101111101100100 1
#774290000000
0#
0(
#774300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#774350000000
0$
0)
#774360000000
1"
1'
b0 +
b0 1
#774410000000
0"
0'
#774420000000
1#
1(
b101111101100100 +
b101111101100100 1
#774470000000
0#
0(
#774480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#774530000000
0$
0)
#774540000000
1"
1'
b0 +
b0 1
#774590000000
0"
0'
#774600000000
1#
1(
b101111101100100 +
b101111101100100 1
#774650000000
0#
0(
#774660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#774710000000
0$
0)
#774720000000
1"
1'
b0 +
b0 1
#774770000000
0"
0'
#774780000000
1#
1(
b101111101100100 +
b101111101100100 1
#774830000000
0#
0(
#774840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#774890000000
0$
0)
#774900000000
1"
1'
b0 +
b0 1
#774950000000
0"
0'
#774960000000
1#
1(
b101111101100100 +
b101111101100100 1
#775010000000
0#
0(
#775020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#775070000000
0$
0)
#775080000000
1"
1'
b0 +
b0 1
#775130000000
0"
0'
#775140000000
1#
1(
b101111101100100 +
b101111101100100 1
#775190000000
0#
0(
#775200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#775250000000
0$
0)
#775260000000
1"
1'
b0 +
b0 1
#775310000000
0"
0'
#775320000000
1#
1(
b101111101100100 +
b101111101100100 1
#775370000000
0#
0(
#775380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#775430000000
0$
0)
#775440000000
1"
1'
b0 +
b0 1
#775490000000
0"
0'
#775500000000
1#
1(
b101111101100100 +
b101111101100100 1
#775550000000
0#
0(
#775560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#775610000000
0$
0)
#775620000000
1"
1'
b0 +
b0 1
#775670000000
0"
0'
#775680000000
1#
1(
b101111101100100 +
b101111101100100 1
#775730000000
0#
0(
#775740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#775790000000
0$
0)
#775800000000
1"
1'
b0 +
b0 1
#775850000000
0"
0'
#775860000000
1#
1(
b101111101100100 +
b101111101100100 1
#775910000000
0#
0(
#775920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#775970000000
0$
0)
#775980000000
1"
1'
b0 +
b0 1
#776030000000
0"
0'
#776040000000
1#
1(
b101111101100100 +
b101111101100100 1
#776090000000
0#
0(
#776100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#776150000000
0$
0)
#776160000000
1"
1'
b0 +
b0 1
#776210000000
0"
0'
#776220000000
1#
1(
b101111101100100 +
b101111101100100 1
#776270000000
0#
0(
#776280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#776330000000
0$
0)
#776340000000
1"
1'
b0 +
b0 1
#776390000000
0"
0'
#776400000000
1#
1(
b101111101100100 +
b101111101100100 1
#776450000000
0#
0(
#776460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#776510000000
0$
0)
#776520000000
1"
1'
b0 +
b0 1
#776570000000
0"
0'
#776580000000
1#
1(
b101111101100100 +
b101111101100100 1
#776630000000
0#
0(
#776640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#776690000000
0$
0)
#776700000000
1"
1'
b0 +
b0 1
#776750000000
0"
0'
#776760000000
1#
1(
b101111101100100 +
b101111101100100 1
#776810000000
0#
0(
#776820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#776870000000
0$
0)
#776880000000
1"
1'
b0 +
b0 1
#776930000000
0"
0'
#776940000000
1#
1(
b101111101100100 +
b101111101100100 1
#776990000000
0#
0(
#777000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#777050000000
0$
0)
#777060000000
1"
1'
b0 +
b0 1
#777110000000
0"
0'
#777120000000
1#
1(
b101111101100100 +
b101111101100100 1
#777170000000
0#
0(
#777180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#777230000000
0$
0)
#777240000000
1"
1'
b0 +
b0 1
#777290000000
0"
0'
#777300000000
1#
1(
b101111101100100 +
b101111101100100 1
#777350000000
0#
0(
#777360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#777410000000
0$
0)
#777420000000
1"
1'
b0 +
b0 1
#777470000000
0"
0'
#777480000000
1#
1(
b101111101100100 +
b101111101100100 1
#777530000000
0#
0(
#777540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#777590000000
0$
0)
#777600000000
1"
1'
b0 +
b0 1
#777650000000
0"
0'
#777660000000
1#
1(
b101111101100100 +
b101111101100100 1
#777710000000
0#
0(
#777720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#777770000000
0$
0)
#777780000000
1"
1'
b0 +
b0 1
#777830000000
0"
0'
#777840000000
1#
1(
b101111101100100 +
b101111101100100 1
#777890000000
0#
0(
#777900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#777950000000
0$
0)
#777960000000
1"
1'
b0 +
b0 1
#778010000000
0"
0'
#778020000000
1#
1(
b101111101100100 +
b101111101100100 1
#778070000000
0#
0(
#778080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#778130000000
0$
0)
#778140000000
1"
1'
b0 +
b0 1
#778190000000
0"
0'
#778200000000
1#
1(
b101111101100100 +
b101111101100100 1
#778250000000
0#
0(
#778260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#778310000000
0$
0)
#778320000000
1"
1'
b0 +
b0 1
#778370000000
0"
0'
#778380000000
1#
1(
b101111101100100 +
b101111101100100 1
#778430000000
0#
0(
#778440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#778490000000
0$
0)
#778500000000
1"
1'
b0 +
b0 1
#778550000000
0"
0'
#778560000000
1#
1(
b101111101100100 +
b101111101100100 1
#778610000000
0#
0(
#778620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#778670000000
0$
0)
#778680000000
1"
1'
b0 +
b0 1
#778730000000
0"
0'
#778740000000
1#
1(
b101111101100100 +
b101111101100100 1
#778790000000
0#
0(
#778800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#778850000000
0$
0)
#778860000000
1"
1'
b0 +
b0 1
#778910000000
0"
0'
#778920000000
1#
1(
b101111101100100 +
b101111101100100 1
#778970000000
0#
0(
#778980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#779030000000
0$
0)
#779040000000
1"
1'
b0 +
b0 1
#779090000000
0"
0'
#779100000000
1#
1(
b101111101100100 +
b101111101100100 1
#779150000000
0#
0(
#779160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#779210000000
0$
0)
#779220000000
1"
1'
b0 +
b0 1
#779270000000
0"
0'
#779280000000
1#
1(
b101111101100100 +
b101111101100100 1
#779330000000
0#
0(
#779340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#779390000000
0$
0)
#779400000000
1"
1'
b0 +
b0 1
#779450000000
0"
0'
#779460000000
1#
1(
b101111101100100 +
b101111101100100 1
#779510000000
0#
0(
#779520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#779570000000
0$
0)
#779580000000
1"
1'
b0 +
b0 1
#779630000000
0"
0'
#779640000000
1#
1(
b101111101100100 +
b101111101100100 1
#779690000000
0#
0(
#779700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#779750000000
0$
0)
#779760000000
1"
1'
b0 +
b0 1
#779810000000
0"
0'
#779820000000
1#
1(
b101111101100100 +
b101111101100100 1
#779870000000
0#
0(
#779880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#779930000000
0$
0)
#779940000000
1"
1'
b0 +
b0 1
#779990000000
0"
0'
#780000000000
1#
1(
b101111101100100 +
b101111101100100 1
#780050000000
0#
0(
#780060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#780110000000
0$
0)
#780120000000
1"
1'
b0 +
b0 1
#780170000000
0"
0'
#780180000000
1#
1(
b101111101100100 +
b101111101100100 1
#780230000000
0#
0(
#780240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#780290000000
0$
0)
#780300000000
1"
1'
b0 +
b0 1
#780350000000
0"
0'
#780360000000
1#
1(
b101111101100100 +
b101111101100100 1
#780410000000
0#
0(
#780420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#780470000000
0$
0)
#780480000000
1"
1'
b0 +
b0 1
#780530000000
0"
0'
#780540000000
1#
1(
b101111101100100 +
b101111101100100 1
#780590000000
0#
0(
#780600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#780650000000
0$
0)
#780660000000
1"
1'
b0 +
b0 1
#780710000000
0"
0'
#780720000000
1#
1(
b101111101100100 +
b101111101100100 1
#780770000000
0#
0(
#780780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#780830000000
0$
0)
#780840000000
1"
1'
b0 +
b0 1
#780890000000
0"
0'
#780900000000
1#
1(
b101111101100100 +
b101111101100100 1
#780950000000
0#
0(
#780960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#781010000000
0$
0)
#781020000000
1"
1'
b0 +
b0 1
#781070000000
0"
0'
#781080000000
1#
1(
b101111101100100 +
b101111101100100 1
#781130000000
0#
0(
#781140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#781190000000
0$
0)
#781200000000
1"
1'
b0 +
b0 1
#781250000000
0"
0'
#781260000000
1#
1(
b101111101100100 +
b101111101100100 1
#781310000000
0#
0(
#781320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#781370000000
0$
0)
#781380000000
1"
1'
b0 +
b0 1
#781430000000
0"
0'
#781440000000
1#
1(
b101111101100100 +
b101111101100100 1
#781490000000
0#
0(
#781500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#781550000000
0$
0)
#781560000000
1"
1'
b0 +
b0 1
#781610000000
0"
0'
#781620000000
1#
1(
b101111101100100 +
b101111101100100 1
#781670000000
0#
0(
#781680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#781730000000
0$
0)
#781740000000
1"
1'
b0 +
b0 1
#781790000000
0"
0'
#781800000000
1#
1(
b101111101100100 +
b101111101100100 1
#781850000000
0#
0(
#781860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#781910000000
0$
0)
#781920000000
1"
1'
b0 +
b0 1
#781970000000
0"
0'
#781980000000
1#
1(
b101111101100100 +
b101111101100100 1
#782030000000
0#
0(
#782040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#782090000000
0$
0)
#782100000000
1"
1'
b0 +
b0 1
#782150000000
0"
0'
#782160000000
1#
1(
b101111101100100 +
b101111101100100 1
#782210000000
0#
0(
#782220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#782270000000
0$
0)
#782280000000
1"
1'
b0 +
b0 1
#782330000000
0"
0'
#782340000000
1#
1(
b101111101100100 +
b101111101100100 1
#782390000000
0#
0(
#782400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#782450000000
0$
0)
#782460000000
1"
1'
b0 +
b0 1
#782510000000
0"
0'
#782520000000
1#
1(
b101111101100100 +
b101111101100100 1
#782570000000
0#
0(
#782580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#782630000000
0$
0)
#782640000000
1"
1'
b0 +
b0 1
#782690000000
0"
0'
#782700000000
1#
1(
b101111101100100 +
b101111101100100 1
#782750000000
0#
0(
#782760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#782810000000
0$
0)
#782820000000
1"
1'
b0 +
b0 1
#782870000000
0"
0'
#782880000000
1#
1(
b101111101100100 +
b101111101100100 1
#782930000000
0#
0(
#782940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#782990000000
0$
0)
#783000000000
1"
1'
b0 +
b0 1
#783050000000
0"
0'
#783060000000
1#
1(
b101111101100100 +
b101111101100100 1
#783110000000
0#
0(
#783120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#783170000000
0$
0)
#783180000000
1"
1'
b0 +
b0 1
#783230000000
0"
0'
#783240000000
1#
1(
b101111101100100 +
b101111101100100 1
#783290000000
0#
0(
#783300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#783350000000
0$
0)
#783360000000
1"
1'
b0 +
b0 1
#783410000000
0"
0'
#783420000000
1#
1(
b101111101100100 +
b101111101100100 1
#783470000000
0#
0(
#783480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#783530000000
0$
0)
#783540000000
1"
1'
b0 +
b0 1
#783590000000
0"
0'
#783600000000
1#
1(
b101111101100100 +
b101111101100100 1
#783650000000
0#
0(
#783660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#783710000000
0$
0)
#783720000000
1"
1'
b0 +
b0 1
#783770000000
0"
0'
#783780000000
1#
1(
b101111101100100 +
b101111101100100 1
#783830000000
0#
0(
#783840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#783890000000
0$
0)
#783900000000
1"
1'
b0 +
b0 1
#783950000000
0"
0'
#783960000000
1#
1(
b101111101100100 +
b101111101100100 1
#784010000000
0#
0(
#784020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#784070000000
0$
0)
#784080000000
1"
1'
b0 +
b0 1
#784130000000
0"
0'
#784140000000
1#
1(
b101111101100100 +
b101111101100100 1
#784190000000
0#
0(
#784200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#784250000000
0$
0)
#784260000000
1"
1'
b0 +
b0 1
#784310000000
0"
0'
#784320000000
1#
1(
b101111101100100 +
b101111101100100 1
#784370000000
0#
0(
#784380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#784430000000
0$
0)
#784440000000
1"
1'
b0 +
b0 1
#784490000000
0"
0'
#784500000000
1#
1(
b101111101100100 +
b101111101100100 1
#784550000000
0#
0(
#784560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#784610000000
0$
0)
#784620000000
1"
1'
b0 +
b0 1
#784670000000
0"
0'
#784680000000
1#
1(
b101111101100100 +
b101111101100100 1
#784730000000
0#
0(
#784740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#784790000000
0$
0)
#784800000000
1"
1'
b0 +
b0 1
#784850000000
0"
0'
#784860000000
1#
1(
b101111101100100 +
b101111101100100 1
#784910000000
0#
0(
#784920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#784970000000
0$
0)
#784980000000
1"
1'
b0 +
b0 1
#785030000000
0"
0'
#785040000000
1#
1(
b101111101100100 +
b101111101100100 1
#785090000000
0#
0(
#785100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#785150000000
0$
0)
#785160000000
1"
1'
b0 +
b0 1
#785210000000
0"
0'
#785220000000
1#
1(
b101111101100100 +
b101111101100100 1
#785270000000
0#
0(
#785280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#785330000000
0$
0)
#785340000000
1"
1'
b0 +
b0 1
#785390000000
0"
0'
#785400000000
1#
1(
b101111101100100 +
b101111101100100 1
#785450000000
0#
0(
#785460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#785510000000
0$
0)
#785520000000
1"
1'
b0 +
b0 1
#785570000000
0"
0'
#785580000000
1#
1(
b101111101100100 +
b101111101100100 1
#785630000000
0#
0(
#785640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#785690000000
0$
0)
#785700000000
1"
1'
b0 +
b0 1
#785750000000
0"
0'
#785760000000
1#
1(
b101111101100100 +
b101111101100100 1
#785810000000
0#
0(
#785820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#785870000000
0$
0)
#785880000000
1"
1'
b0 +
b0 1
#785930000000
0"
0'
#785940000000
1#
1(
b101111101100100 +
b101111101100100 1
#785990000000
0#
0(
#786000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#786050000000
0$
0)
#786060000000
1"
1'
b0 +
b0 1
#786110000000
0"
0'
#786120000000
1#
1(
b101111101100100 +
b101111101100100 1
#786170000000
0#
0(
#786180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#786230000000
0$
0)
#786240000000
1"
1'
b0 +
b0 1
#786290000000
0"
0'
#786300000000
1#
1(
b101111101100100 +
b101111101100100 1
#786350000000
0#
0(
#786360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#786410000000
0$
0)
#786420000000
1"
1'
b0 +
b0 1
#786470000000
0"
0'
#786480000000
1#
1(
b101111101100100 +
b101111101100100 1
#786530000000
0#
0(
#786540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#786590000000
0$
0)
#786600000000
1"
1'
b0 +
b0 1
#786650000000
0"
0'
#786660000000
1#
1(
b101111101100100 +
b101111101100100 1
#786710000000
0#
0(
#786720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#786770000000
0$
0)
#786780000000
1"
1'
b0 +
b0 1
#786830000000
0"
0'
#786840000000
1#
1(
b101111101100100 +
b101111101100100 1
#786890000000
0#
0(
#786900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#786950000000
0$
0)
#786960000000
1"
1'
b0 +
b0 1
#787010000000
0"
0'
#787020000000
1#
1(
b101111101100100 +
b101111101100100 1
#787070000000
0#
0(
#787080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#787130000000
0$
0)
#787140000000
1"
1'
b0 +
b0 1
#787190000000
0"
0'
#787200000000
1#
1(
b101111101100100 +
b101111101100100 1
#787250000000
0#
0(
#787260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#787310000000
0$
0)
#787320000000
1"
1'
b0 +
b0 1
#787370000000
0"
0'
#787380000000
1#
1(
b101111101100100 +
b101111101100100 1
#787430000000
0#
0(
#787440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#787490000000
0$
0)
#787500000000
1"
1'
b0 +
b0 1
#787550000000
0"
0'
#787560000000
1#
1(
b101111101100100 +
b101111101100100 1
#787610000000
0#
0(
#787620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#787670000000
0$
0)
#787680000000
1"
1'
b0 +
b0 1
#787730000000
0"
0'
#787740000000
1#
1(
b101111101100100 +
b101111101100100 1
#787790000000
0#
0(
#787800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#787850000000
0$
0)
#787860000000
1"
1'
b0 +
b0 1
#787910000000
0"
0'
#787920000000
1#
1(
b101111101100100 +
b101111101100100 1
#787970000000
0#
0(
#787980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#788030000000
0$
0)
#788040000000
1"
1'
b0 +
b0 1
#788090000000
0"
0'
#788100000000
1#
1(
b101111101100100 +
b101111101100100 1
#788150000000
0#
0(
#788160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#788210000000
0$
0)
#788220000000
1"
1'
b0 +
b0 1
#788270000000
0"
0'
#788280000000
1#
1(
b101111101100100 +
b101111101100100 1
#788330000000
0#
0(
#788340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#788390000000
0$
0)
#788400000000
1"
1'
b0 +
b0 1
#788450000000
0"
0'
#788460000000
1#
1(
b101111101100100 +
b101111101100100 1
#788510000000
0#
0(
#788520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#788570000000
0$
0)
#788580000000
1"
1'
b0 +
b0 1
#788630000000
0"
0'
#788640000000
1#
1(
b101111101100100 +
b101111101100100 1
#788690000000
0#
0(
#788700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#788750000000
0$
0)
#788760000000
1"
1'
b0 +
b0 1
#788810000000
0"
0'
#788820000000
1#
1(
b101111101100100 +
b101111101100100 1
#788870000000
0#
0(
#788880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#788930000000
0$
0)
#788940000000
1"
1'
b0 +
b0 1
#788990000000
0"
0'
#789000000000
1#
1(
b101111101100100 +
b101111101100100 1
#789050000000
0#
0(
#789060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#789110000000
0$
0)
#789120000000
1"
1'
b0 +
b0 1
#789170000000
0"
0'
#789180000000
1#
1(
b101111101100100 +
b101111101100100 1
#789230000000
0#
0(
#789240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#789290000000
0$
0)
#789300000000
1"
1'
b0 +
b0 1
#789350000000
0"
0'
#789360000000
1#
1(
b101111101100100 +
b101111101100100 1
#789410000000
0#
0(
#789420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#789470000000
0$
0)
#789480000000
1"
1'
b0 +
b0 1
#789530000000
0"
0'
#789540000000
1#
1(
b101111101100100 +
b101111101100100 1
#789590000000
0#
0(
#789600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#789650000000
0$
0)
#789660000000
1"
1'
b0 +
b0 1
#789710000000
0"
0'
#789720000000
1#
1(
b101111101100100 +
b101111101100100 1
#789770000000
0#
0(
#789780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#789830000000
0$
0)
#789840000000
1"
1'
b0 +
b0 1
#789890000000
0"
0'
#789900000000
1#
1(
b101111101100100 +
b101111101100100 1
#789950000000
0#
0(
#789960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#790010000000
0$
0)
#790020000000
1"
1'
b0 +
b0 1
#790070000000
0"
0'
#790080000000
1#
1(
b101111101100100 +
b101111101100100 1
#790130000000
0#
0(
#790140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#790190000000
0$
0)
#790200000000
1"
1'
b0 +
b0 1
#790250000000
0"
0'
#790260000000
1#
1(
b101111101100100 +
b101111101100100 1
#790310000000
0#
0(
#790320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#790370000000
0$
0)
#790380000000
1"
1'
b0 +
b0 1
#790430000000
0"
0'
#790440000000
1#
1(
b101111101100100 +
b101111101100100 1
#790490000000
0#
0(
#790500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#790550000000
0$
0)
#790560000000
1"
1'
b0 +
b0 1
#790610000000
0"
0'
#790620000000
1#
1(
b101111101100100 +
b101111101100100 1
#790670000000
0#
0(
#790680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#790730000000
0$
0)
#790740000000
1"
1'
b0 +
b0 1
#790790000000
0"
0'
#790800000000
1#
1(
b101111101100100 +
b101111101100100 1
#790850000000
0#
0(
#790860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#790910000000
0$
0)
#790920000000
1"
1'
b0 +
b0 1
#790970000000
0"
0'
#790980000000
1#
1(
b101111101100100 +
b101111101100100 1
#791030000000
0#
0(
#791040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#791090000000
0$
0)
#791100000000
1"
1'
b0 +
b0 1
#791150000000
0"
0'
#791160000000
1#
1(
b101111101100100 +
b101111101100100 1
#791210000000
0#
0(
#791220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#791270000000
0$
0)
#791280000000
1"
1'
b0 +
b0 1
#791330000000
0"
0'
#791340000000
1#
1(
b101111101100100 +
b101111101100100 1
#791390000000
0#
0(
#791400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#791450000000
0$
0)
#791460000000
1"
1'
b0 +
b0 1
#791510000000
0"
0'
#791520000000
1#
1(
b101111101100100 +
b101111101100100 1
#791570000000
0#
0(
#791580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#791630000000
0$
0)
#791640000000
1"
1'
b0 +
b0 1
#791690000000
0"
0'
#791700000000
1#
1(
b101111101100100 +
b101111101100100 1
#791750000000
0#
0(
#791760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#791810000000
0$
0)
#791820000000
1"
1'
b0 +
b0 1
#791870000000
0"
0'
#791880000000
1#
1(
b101111101100100 +
b101111101100100 1
#791930000000
0#
0(
#791940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#791990000000
0$
0)
#792000000000
1"
1'
b0 +
b0 1
#792050000000
0"
0'
#792060000000
1#
1(
b101111101100100 +
b101111101100100 1
#792110000000
0#
0(
#792120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#792170000000
0$
0)
#792180000000
1"
1'
b0 +
b0 1
#792230000000
0"
0'
#792240000000
1#
1(
b101111101100100 +
b101111101100100 1
#792290000000
0#
0(
#792300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#792350000000
0$
0)
#792360000000
1"
1'
b0 +
b0 1
#792410000000
0"
0'
#792420000000
1#
1(
b101111101100100 +
b101111101100100 1
#792470000000
0#
0(
#792480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#792530000000
0$
0)
#792540000000
1"
1'
b0 +
b0 1
#792590000000
0"
0'
#792600000000
1#
1(
b101111101100100 +
b101111101100100 1
#792650000000
0#
0(
#792660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#792710000000
0$
0)
#792720000000
1"
1'
b0 +
b0 1
#792770000000
0"
0'
#792780000000
1#
1(
b101111101100100 +
b101111101100100 1
#792830000000
0#
0(
#792840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#792890000000
0$
0)
#792900000000
1"
1'
b0 +
b0 1
#792950000000
0"
0'
#792960000000
1#
1(
b101111101100100 +
b101111101100100 1
#793010000000
0#
0(
#793020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#793070000000
0$
0)
#793080000000
1"
1'
b0 +
b0 1
#793130000000
0"
0'
#793140000000
1#
1(
b101111101100100 +
b101111101100100 1
#793190000000
0#
0(
#793200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#793250000000
0$
0)
#793260000000
1"
1'
b0 +
b0 1
#793310000000
0"
0'
#793320000000
1#
1(
b101111101100100 +
b101111101100100 1
#793370000000
0#
0(
#793380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#793430000000
0$
0)
#793440000000
1"
1'
b0 +
b0 1
#793490000000
0"
0'
#793500000000
1#
1(
b101111101100100 +
b101111101100100 1
#793550000000
0#
0(
#793560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#793610000000
0$
0)
#793620000000
1"
1'
b0 +
b0 1
#793670000000
0"
0'
#793680000000
1#
1(
b101111101100100 +
b101111101100100 1
#793730000000
0#
0(
#793740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#793790000000
0$
0)
#793800000000
1"
1'
b0 +
b0 1
#793850000000
0"
0'
#793860000000
1#
1(
b101111101100100 +
b101111101100100 1
#793910000000
0#
0(
#793920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#793970000000
0$
0)
#793980000000
1"
1'
b0 +
b0 1
#794030000000
0"
0'
#794040000000
1#
1(
b101111101100100 +
b101111101100100 1
#794090000000
0#
0(
#794100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#794150000000
0$
0)
#794160000000
1"
1'
b0 +
b0 1
#794210000000
0"
0'
#794220000000
1#
1(
b101111101100100 +
b101111101100100 1
#794270000000
0#
0(
#794280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#794330000000
0$
0)
#794340000000
1"
1'
b0 +
b0 1
#794390000000
0"
0'
#794400000000
1#
1(
b101111101100100 +
b101111101100100 1
#794450000000
0#
0(
#794460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#794510000000
0$
0)
#794520000000
1"
1'
b0 +
b0 1
#794570000000
0"
0'
#794580000000
1#
1(
b101111101100100 +
b101111101100100 1
#794630000000
0#
0(
#794640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#794690000000
0$
0)
#794700000000
1"
1'
b0 +
b0 1
#794750000000
0"
0'
#794760000000
1#
1(
b101111101100100 +
b101111101100100 1
#794810000000
0#
0(
#794820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#794870000000
0$
0)
#794880000000
1"
1'
b0 +
b0 1
#794930000000
0"
0'
#794940000000
1#
1(
b101111101100100 +
b101111101100100 1
#794990000000
0#
0(
#795000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#795050000000
0$
0)
#795060000000
1"
1'
b0 +
b0 1
#795110000000
0"
0'
#795120000000
1#
1(
b101111101100100 +
b101111101100100 1
#795170000000
0#
0(
#795180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#795230000000
0$
0)
#795240000000
1"
1'
b0 +
b0 1
#795290000000
0"
0'
#795300000000
1#
1(
b101111101100100 +
b101111101100100 1
#795350000000
0#
0(
#795360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#795410000000
0$
0)
#795420000000
1"
1'
b0 +
b0 1
#795470000000
0"
0'
#795480000000
1#
1(
b101111101100100 +
b101111101100100 1
#795530000000
0#
0(
#795540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#795590000000
0$
0)
#795600000000
1"
1'
b0 +
b0 1
#795650000000
0"
0'
#795660000000
1#
1(
b101111101100100 +
b101111101100100 1
#795710000000
0#
0(
#795720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#795770000000
0$
0)
#795780000000
1"
1'
b0 +
b0 1
#795830000000
0"
0'
#795840000000
1#
1(
b101111101100100 +
b101111101100100 1
#795890000000
0#
0(
#795900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#795950000000
0$
0)
#795960000000
1"
1'
b0 +
b0 1
#796010000000
0"
0'
#796020000000
1#
1(
b101111101100100 +
b101111101100100 1
#796070000000
0#
0(
#796080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#796130000000
0$
0)
#796140000000
1"
1'
b0 +
b0 1
#796190000000
0"
0'
#796200000000
1#
1(
b101111101100100 +
b101111101100100 1
#796250000000
0#
0(
#796260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#796310000000
0$
0)
#796320000000
1"
1'
b0 +
b0 1
#796370000000
0"
0'
#796380000000
1#
1(
b101111101100100 +
b101111101100100 1
#796430000000
0#
0(
#796440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#796490000000
0$
0)
#796500000000
1"
1'
b0 +
b0 1
#796550000000
0"
0'
#796560000000
1#
1(
b101111101100100 +
b101111101100100 1
#796610000000
0#
0(
#796620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#796670000000
0$
0)
#796680000000
1"
1'
b0 +
b0 1
#796730000000
0"
0'
#796740000000
1#
1(
b101111101100100 +
b101111101100100 1
#796790000000
0#
0(
#796800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#796850000000
0$
0)
#796860000000
1"
1'
b0 +
b0 1
#796910000000
0"
0'
#796920000000
1#
1(
b101111101100100 +
b101111101100100 1
#796970000000
0#
0(
#796980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#797030000000
0$
0)
#797040000000
1"
1'
b0 +
b0 1
#797090000000
0"
0'
#797100000000
1#
1(
b101111101100100 +
b101111101100100 1
#797150000000
0#
0(
#797160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#797210000000
0$
0)
#797220000000
1"
1'
b0 +
b0 1
#797270000000
0"
0'
#797280000000
1#
1(
b101111101100100 +
b101111101100100 1
#797330000000
0#
0(
#797340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#797390000000
0$
0)
#797400000000
1"
1'
b0 +
b0 1
#797450000000
0"
0'
#797460000000
1#
1(
b101111101100100 +
b101111101100100 1
#797510000000
0#
0(
#797520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#797570000000
0$
0)
#797580000000
1"
1'
b0 +
b0 1
#797630000000
0"
0'
#797640000000
1#
1(
b101111101100100 +
b101111101100100 1
#797690000000
0#
0(
#797700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#797750000000
0$
0)
#797760000000
1"
1'
b0 +
b0 1
#797810000000
0"
0'
#797820000000
1#
1(
b101111101100100 +
b101111101100100 1
#797870000000
0#
0(
#797880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#797930000000
0$
0)
#797940000000
1"
1'
b0 +
b0 1
#797990000000
0"
0'
#798000000000
1#
1(
b101111101100100 +
b101111101100100 1
#798050000000
0#
0(
#798060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#798110000000
0$
0)
#798120000000
1"
1'
b0 +
b0 1
#798170000000
0"
0'
#798180000000
1#
1(
b101111101100100 +
b101111101100100 1
#798230000000
0#
0(
#798240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#798290000000
0$
0)
#798300000000
1"
1'
b0 +
b0 1
#798350000000
0"
0'
#798360000000
1#
1(
b101111101100100 +
b101111101100100 1
#798410000000
0#
0(
#798420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#798470000000
0$
0)
#798480000000
1"
1'
b0 +
b0 1
#798530000000
0"
0'
#798540000000
1#
1(
b101111101100100 +
b101111101100100 1
#798590000000
0#
0(
#798600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#798650000000
0$
0)
#798660000000
1"
1'
b0 +
b0 1
#798710000000
0"
0'
#798720000000
1#
1(
b101111101100100 +
b101111101100100 1
#798770000000
0#
0(
#798780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#798830000000
0$
0)
#798840000000
1"
1'
b0 +
b0 1
#798890000000
0"
0'
#798900000000
1#
1(
b101111101100100 +
b101111101100100 1
#798950000000
0#
0(
#798960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#799010000000
0$
0)
#799020000000
1"
1'
b0 +
b0 1
#799070000000
0"
0'
#799080000000
1#
1(
b101111101100100 +
b101111101100100 1
#799130000000
0#
0(
#799140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#799190000000
0$
0)
#799200000000
1"
1'
b0 +
b0 1
#799250000000
0"
0'
#799260000000
1#
1(
b101111101100100 +
b101111101100100 1
#799310000000
0#
0(
#799320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#799370000000
0$
0)
#799380000000
1"
1'
b0 +
b0 1
#799430000000
0"
0'
#799440000000
1#
1(
b101111101100100 +
b101111101100100 1
#799490000000
0#
0(
#799500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#799550000000
0$
0)
#799560000000
1"
1'
b0 +
b0 1
#799610000000
0"
0'
#799620000000
1#
1(
b101111101100100 +
b101111101100100 1
#799670000000
0#
0(
#799680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#799730000000
0$
0)
#799740000000
1"
1'
b0 +
b0 1
#799790000000
0"
0'
#799800000000
1#
1(
b101111101100100 +
b101111101100100 1
#799850000000
0#
0(
#799860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#799910000000
0$
0)
#799920000000
1"
1'
b0 +
b0 1
#799970000000
0"
0'
#799980000000
1#
1(
b101111101100100 +
b101111101100100 1
#800030000000
0#
0(
#800040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#800090000000
0$
0)
#800100000000
1"
1'
b0 +
b0 1
#800150000000
0"
0'
#800160000000
1#
1(
b101111101100100 +
b101111101100100 1
#800210000000
0#
0(
#800220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#800270000000
0$
0)
#800280000000
1"
1'
b0 +
b0 1
#800330000000
0"
0'
#800340000000
1#
1(
b101111101100100 +
b101111101100100 1
#800390000000
0#
0(
#800400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#800450000000
0$
0)
#800460000000
1"
1'
b0 +
b0 1
#800510000000
0"
0'
#800520000000
1#
1(
b101111101100100 +
b101111101100100 1
#800570000000
0#
0(
#800580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#800630000000
0$
0)
#800640000000
1"
1'
b0 +
b0 1
#800690000000
0"
0'
#800700000000
1#
1(
b101111101100100 +
b101111101100100 1
#800750000000
0#
0(
#800760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#800810000000
0$
0)
#800820000000
1"
1'
b0 +
b0 1
#800870000000
0"
0'
#800880000000
1#
1(
b101111101100100 +
b101111101100100 1
#800930000000
0#
0(
#800940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#800990000000
0$
0)
#801000000000
1"
1'
b0 +
b0 1
#801050000000
0"
0'
#801060000000
1#
1(
b101111101100100 +
b101111101100100 1
#801110000000
0#
0(
#801120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#801170000000
0$
0)
#801180000000
1"
1'
b0 +
b0 1
#801230000000
0"
0'
#801240000000
1#
1(
b101111101100100 +
b101111101100100 1
#801290000000
0#
0(
#801300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#801350000000
0$
0)
#801360000000
1"
1'
b0 +
b0 1
#801410000000
0"
0'
#801420000000
1#
1(
b101111101100100 +
b101111101100100 1
#801470000000
0#
0(
#801480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#801530000000
0$
0)
#801540000000
1"
1'
b0 +
b0 1
#801590000000
0"
0'
#801600000000
1#
1(
b101111101100100 +
b101111101100100 1
#801650000000
0#
0(
#801660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#801710000000
0$
0)
#801720000000
1"
1'
b0 +
b0 1
#801770000000
0"
0'
#801780000000
1#
1(
b101111101100100 +
b101111101100100 1
#801830000000
0#
0(
#801840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#801890000000
0$
0)
#801900000000
1"
1'
b0 +
b0 1
#801950000000
0"
0'
#801960000000
1#
1(
b101111101100100 +
b101111101100100 1
#802010000000
0#
0(
#802020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#802070000000
0$
0)
#802080000000
1"
1'
b0 +
b0 1
#802130000000
0"
0'
#802140000000
1#
1(
b101111101100100 +
b101111101100100 1
#802190000000
0#
0(
#802200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#802250000000
0$
0)
#802260000000
1"
1'
b0 +
b0 1
#802310000000
0"
0'
#802320000000
1#
1(
b101111101100100 +
b101111101100100 1
#802370000000
0#
0(
#802380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#802430000000
0$
0)
#802440000000
1"
1'
b0 +
b0 1
#802490000000
0"
0'
#802500000000
1#
1(
b101111101100100 +
b101111101100100 1
#802550000000
0#
0(
#802560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#802610000000
0$
0)
#802620000000
1"
1'
b0 +
b0 1
#802670000000
0"
0'
#802680000000
1#
1(
b101111101100100 +
b101111101100100 1
#802730000000
0#
0(
#802740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#802790000000
0$
0)
#802800000000
1"
1'
b0 +
b0 1
#802850000000
0"
0'
#802860000000
1#
1(
b101111101100100 +
b101111101100100 1
#802910000000
0#
0(
#802920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#802970000000
0$
0)
#802980000000
1"
1'
b0 +
b0 1
#803030000000
0"
0'
#803040000000
1#
1(
b101111101100100 +
b101111101100100 1
#803090000000
0#
0(
#803100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#803150000000
0$
0)
#803160000000
1"
1'
b0 +
b0 1
#803210000000
0"
0'
#803220000000
1#
1(
b101111101100100 +
b101111101100100 1
#803270000000
0#
0(
#803280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#803330000000
0$
0)
#803340000000
1"
1'
b0 +
b0 1
#803390000000
0"
0'
#803400000000
1#
1(
b101111101100100 +
b101111101100100 1
#803450000000
0#
0(
#803460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#803510000000
0$
0)
#803520000000
1"
1'
b0 +
b0 1
#803570000000
0"
0'
#803580000000
1#
1(
b101111101100100 +
b101111101100100 1
#803630000000
0#
0(
#803640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#803690000000
0$
0)
#803700000000
1"
1'
b0 +
b0 1
#803750000000
0"
0'
#803760000000
1#
1(
b101111101100100 +
b101111101100100 1
#803810000000
0#
0(
#803820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#803870000000
0$
0)
#803880000000
1"
1'
b0 +
b0 1
#803930000000
0"
0'
#803940000000
1#
1(
b101111101100100 +
b101111101100100 1
#803990000000
0#
0(
#804000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#804050000000
0$
0)
#804060000000
1"
1'
b0 +
b0 1
#804110000000
0"
0'
#804120000000
1#
1(
b101111101100100 +
b101111101100100 1
#804170000000
0#
0(
#804180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#804230000000
0$
0)
#804240000000
1"
1'
b0 +
b0 1
#804290000000
0"
0'
#804300000000
1#
1(
b101111101100100 +
b101111101100100 1
#804350000000
0#
0(
#804360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#804410000000
0$
0)
#804420000000
1"
1'
b0 +
b0 1
#804470000000
0"
0'
#804480000000
1#
1(
b101111101100100 +
b101111101100100 1
#804530000000
0#
0(
#804540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#804590000000
0$
0)
#804600000000
1"
1'
b0 +
b0 1
#804650000000
0"
0'
#804660000000
1#
1(
b101111101100100 +
b101111101100100 1
#804710000000
0#
0(
#804720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#804770000000
0$
0)
#804780000000
1"
1'
b0 +
b0 1
#804830000000
0"
0'
#804840000000
1#
1(
b101111101100100 +
b101111101100100 1
#804890000000
0#
0(
#804900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#804950000000
0$
0)
#804960000000
1"
1'
b0 +
b0 1
#805010000000
0"
0'
#805020000000
1#
1(
b101111101100100 +
b101111101100100 1
#805070000000
0#
0(
#805080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#805130000000
0$
0)
#805140000000
1"
1'
b0 +
b0 1
#805190000000
0"
0'
#805200000000
1#
1(
b101111101100100 +
b101111101100100 1
#805250000000
0#
0(
#805260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#805310000000
0$
0)
#805320000000
1"
1'
b0 +
b0 1
#805370000000
0"
0'
#805380000000
1#
1(
b101111101100100 +
b101111101100100 1
#805430000000
0#
0(
#805440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#805490000000
0$
0)
#805500000000
1"
1'
b0 +
b0 1
#805550000000
0"
0'
#805560000000
1#
1(
b101111101100100 +
b101111101100100 1
#805610000000
0#
0(
#805620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#805670000000
0$
0)
#805680000000
1"
1'
b0 +
b0 1
#805730000000
0"
0'
#805740000000
1#
1(
b101111101100100 +
b101111101100100 1
#805790000000
0#
0(
#805800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#805850000000
0$
0)
#805860000000
1"
1'
b0 +
b0 1
#805910000000
0"
0'
#805920000000
1#
1(
b101111101100100 +
b101111101100100 1
#805970000000
0#
0(
#805980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#806030000000
0$
0)
#806040000000
1"
1'
b0 +
b0 1
#806090000000
0"
0'
#806100000000
1#
1(
b101111101100100 +
b101111101100100 1
#806150000000
0#
0(
#806160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#806210000000
0$
0)
#806220000000
1"
1'
b0 +
b0 1
#806270000000
0"
0'
#806280000000
1#
1(
b101111101100100 +
b101111101100100 1
#806330000000
0#
0(
#806340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#806390000000
0$
0)
#806400000000
1"
1'
b0 +
b0 1
#806450000000
0"
0'
#806460000000
1#
1(
b101111101100100 +
b101111101100100 1
#806510000000
0#
0(
#806520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#806570000000
0$
0)
#806580000000
1"
1'
b0 +
b0 1
#806630000000
0"
0'
#806640000000
1#
1(
b101111101100100 +
b101111101100100 1
#806690000000
0#
0(
#806700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#806750000000
0$
0)
#806760000000
1"
1'
b0 +
b0 1
#806810000000
0"
0'
#806820000000
1#
1(
b101111101100100 +
b101111101100100 1
#806870000000
0#
0(
#806880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#806930000000
0$
0)
#806940000000
1"
1'
b0 +
b0 1
#806990000000
0"
0'
#807000000000
1#
1(
b101111101100100 +
b101111101100100 1
#807050000000
0#
0(
#807060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#807110000000
0$
0)
#807120000000
1"
1'
b0 +
b0 1
#807170000000
0"
0'
#807180000000
1#
1(
b101111101100100 +
b101111101100100 1
#807230000000
0#
0(
#807240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#807290000000
0$
0)
#807300000000
1"
1'
b0 +
b0 1
#807350000000
0"
0'
#807360000000
1#
1(
b101111101100100 +
b101111101100100 1
#807410000000
0#
0(
#807420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#807470000000
0$
0)
#807480000000
1"
1'
b0 +
b0 1
#807530000000
0"
0'
#807540000000
1#
1(
b101111101100100 +
b101111101100100 1
#807590000000
0#
0(
#807600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#807650000000
0$
0)
#807660000000
1"
1'
b0 +
b0 1
#807710000000
0"
0'
#807720000000
1#
1(
b101111101100100 +
b101111101100100 1
#807770000000
0#
0(
#807780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#807830000000
0$
0)
#807840000000
1"
1'
b0 +
b0 1
#807890000000
0"
0'
#807900000000
1#
1(
b101111101100100 +
b101111101100100 1
#807950000000
0#
0(
#807960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#808010000000
0$
0)
#808020000000
1"
1'
b0 +
b0 1
#808070000000
0"
0'
#808080000000
1#
1(
b101111101100100 +
b101111101100100 1
#808130000000
0#
0(
#808140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#808190000000
0$
0)
#808200000000
1"
1'
b0 +
b0 1
#808250000000
0"
0'
#808260000000
1#
1(
b101111101100100 +
b101111101100100 1
#808310000000
0#
0(
#808320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#808370000000
0$
0)
#808380000000
1"
1'
b0 +
b0 1
#808430000000
0"
0'
#808440000000
1#
1(
b101111101100100 +
b101111101100100 1
#808490000000
0#
0(
#808500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#808550000000
0$
0)
#808560000000
1"
1'
b0 +
b0 1
#808610000000
0"
0'
#808620000000
1#
1(
b101111101100100 +
b101111101100100 1
#808670000000
0#
0(
#808680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#808730000000
0$
0)
#808740000000
1"
1'
b0 +
b0 1
#808790000000
0"
0'
#808800000000
1#
1(
b101111101100100 +
b101111101100100 1
#808850000000
0#
0(
#808860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#808910000000
0$
0)
#808920000000
1"
1'
b0 +
b0 1
#808970000000
0"
0'
#808980000000
1#
1(
b101111101100100 +
b101111101100100 1
#809030000000
0#
0(
#809040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#809090000000
0$
0)
#809100000000
1"
1'
b0 +
b0 1
#809150000000
0"
0'
#809160000000
1#
1(
b101111101100100 +
b101111101100100 1
#809210000000
0#
0(
#809220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#809270000000
0$
0)
#809280000000
1"
1'
b0 +
b0 1
#809330000000
0"
0'
#809340000000
1#
1(
b101111101100100 +
b101111101100100 1
#809390000000
0#
0(
#809400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#809450000000
0$
0)
#809460000000
1"
1'
b0 +
b0 1
#809510000000
0"
0'
#809520000000
1#
1(
b101111101100100 +
b101111101100100 1
#809570000000
0#
0(
#809580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#809630000000
0$
0)
#809640000000
1"
1'
b0 +
b0 1
#809690000000
0"
0'
#809700000000
1#
1(
b101111101100100 +
b101111101100100 1
#809750000000
0#
0(
#809760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#809810000000
0$
0)
#809820000000
1"
1'
b0 +
b0 1
#809870000000
0"
0'
#809880000000
1#
1(
b101111101100100 +
b101111101100100 1
#809930000000
0#
0(
#809940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#809990000000
0$
0)
#810000000000
1"
1'
b0 +
b0 1
#810050000000
0"
0'
#810060000000
1#
1(
b101111101100100 +
b101111101100100 1
#810110000000
0#
0(
#810120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#810170000000
0$
0)
#810180000000
1"
1'
b0 +
b0 1
#810230000000
0"
0'
#810240000000
1#
1(
b101111101100100 +
b101111101100100 1
#810290000000
0#
0(
#810300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#810350000000
0$
0)
#810360000000
1"
1'
b0 +
b0 1
#810410000000
0"
0'
#810420000000
1#
1(
b101111101100100 +
b101111101100100 1
#810470000000
0#
0(
#810480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#810530000000
0$
0)
#810540000000
1"
1'
b0 +
b0 1
#810590000000
0"
0'
#810600000000
1#
1(
b101111101100100 +
b101111101100100 1
#810650000000
0#
0(
#810660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#810710000000
0$
0)
#810720000000
1"
1'
b0 +
b0 1
#810770000000
0"
0'
#810780000000
1#
1(
b101111101100100 +
b101111101100100 1
#810830000000
0#
0(
#810840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#810890000000
0$
0)
#810900000000
1"
1'
b0 +
b0 1
#810950000000
0"
0'
#810960000000
1#
1(
b101111101100100 +
b101111101100100 1
#811010000000
0#
0(
#811020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#811070000000
0$
0)
#811080000000
1"
1'
b0 +
b0 1
#811130000000
0"
0'
#811140000000
1#
1(
b101111101100100 +
b101111101100100 1
#811190000000
0#
0(
#811200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#811250000000
0$
0)
#811260000000
1"
1'
b0 +
b0 1
#811310000000
0"
0'
#811320000000
1#
1(
b101111101100100 +
b101111101100100 1
#811370000000
0#
0(
#811380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#811430000000
0$
0)
#811440000000
1"
1'
b0 +
b0 1
#811490000000
0"
0'
#811500000000
1#
1(
b101111101100100 +
b101111101100100 1
#811550000000
0#
0(
#811560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#811610000000
0$
0)
#811620000000
1"
1'
b0 +
b0 1
#811670000000
0"
0'
#811680000000
1#
1(
b101111101100100 +
b101111101100100 1
#811730000000
0#
0(
#811740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#811790000000
0$
0)
#811800000000
1"
1'
b0 +
b0 1
#811850000000
0"
0'
#811860000000
1#
1(
b101111101100100 +
b101111101100100 1
#811910000000
0#
0(
#811920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#811970000000
0$
0)
#811980000000
1"
1'
b0 +
b0 1
#812030000000
0"
0'
#812040000000
1#
1(
b101111101100100 +
b101111101100100 1
#812090000000
0#
0(
#812100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#812150000000
0$
0)
#812160000000
1"
1'
b0 +
b0 1
#812210000000
0"
0'
#812220000000
1#
1(
b101111101100100 +
b101111101100100 1
#812270000000
0#
0(
#812280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#812330000000
0$
0)
#812340000000
1"
1'
b0 +
b0 1
#812390000000
0"
0'
#812400000000
1#
1(
b101111101100100 +
b101111101100100 1
#812450000000
0#
0(
#812460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#812510000000
0$
0)
#812520000000
1"
1'
b0 +
b0 1
#812570000000
0"
0'
#812580000000
1#
1(
b101111101100100 +
b101111101100100 1
#812630000000
0#
0(
#812640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#812690000000
0$
0)
#812700000000
1"
1'
b0 +
b0 1
#812750000000
0"
0'
#812760000000
1#
1(
b101111101100100 +
b101111101100100 1
#812810000000
0#
0(
#812820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#812870000000
0$
0)
#812880000000
1"
1'
b0 +
b0 1
#812930000000
0"
0'
#812940000000
1#
1(
b101111101100100 +
b101111101100100 1
#812990000000
0#
0(
#813000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#813050000000
0$
0)
#813060000000
1"
1'
b0 +
b0 1
#813110000000
0"
0'
#813120000000
1#
1(
b101111101100100 +
b101111101100100 1
#813170000000
0#
0(
#813180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#813230000000
0$
0)
#813240000000
1"
1'
b0 +
b0 1
#813290000000
0"
0'
#813300000000
1#
1(
b101111101100100 +
b101111101100100 1
#813350000000
0#
0(
#813360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#813410000000
0$
0)
#813420000000
1"
1'
b0 +
b0 1
#813470000000
0"
0'
#813480000000
1#
1(
b101111101100100 +
b101111101100100 1
#813530000000
0#
0(
#813540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#813590000000
0$
0)
#813600000000
1"
1'
b0 +
b0 1
#813650000000
0"
0'
#813660000000
1#
1(
b101111101100100 +
b101111101100100 1
#813710000000
0#
0(
#813720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#813770000000
0$
0)
#813780000000
1"
1'
b0 +
b0 1
#813830000000
0"
0'
#813840000000
1#
1(
b101111101100100 +
b101111101100100 1
#813890000000
0#
0(
#813900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#813950000000
0$
0)
#813960000000
1"
1'
b0 +
b0 1
#814010000000
0"
0'
#814020000000
1#
1(
b101111101100100 +
b101111101100100 1
#814070000000
0#
0(
#814080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#814130000000
0$
0)
#814140000000
1"
1'
b0 +
b0 1
#814190000000
0"
0'
#814200000000
1#
1(
b101111101100100 +
b101111101100100 1
#814250000000
0#
0(
#814260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#814310000000
0$
0)
#814320000000
1"
1'
b0 +
b0 1
#814370000000
0"
0'
#814380000000
1#
1(
b101111101100100 +
b101111101100100 1
#814430000000
0#
0(
#814440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#814490000000
0$
0)
#814500000000
1"
1'
b0 +
b0 1
#814550000000
0"
0'
#814560000000
1#
1(
b101111101100100 +
b101111101100100 1
#814610000000
0#
0(
#814620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#814670000000
0$
0)
#814680000000
1"
1'
b0 +
b0 1
#814730000000
0"
0'
#814740000000
1#
1(
b101111101100100 +
b101111101100100 1
#814790000000
0#
0(
#814800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#814850000000
0$
0)
#814860000000
1"
1'
b0 +
b0 1
#814910000000
0"
0'
#814920000000
1#
1(
b101111101100100 +
b101111101100100 1
#814970000000
0#
0(
#814980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#815030000000
0$
0)
#815040000000
1"
1'
b0 +
b0 1
#815090000000
0"
0'
#815100000000
1#
1(
b101111101100100 +
b101111101100100 1
#815150000000
0#
0(
#815160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#815210000000
0$
0)
#815220000000
1"
1'
b0 +
b0 1
#815270000000
0"
0'
#815280000000
1#
1(
b101111101100100 +
b101111101100100 1
#815330000000
0#
0(
#815340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#815390000000
0$
0)
#815400000000
1"
1'
b0 +
b0 1
#815450000000
0"
0'
#815460000000
1#
1(
b101111101100100 +
b101111101100100 1
#815510000000
0#
0(
#815520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#815570000000
0$
0)
#815580000000
1"
1'
b0 +
b0 1
#815630000000
0"
0'
#815640000000
1#
1(
b101111101100100 +
b101111101100100 1
#815690000000
0#
0(
#815700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#815750000000
0$
0)
#815760000000
1"
1'
b0 +
b0 1
#815810000000
0"
0'
#815820000000
1#
1(
b101111101100100 +
b101111101100100 1
#815870000000
0#
0(
#815880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#815930000000
0$
0)
#815940000000
1"
1'
b0 +
b0 1
#815990000000
0"
0'
#816000000000
1#
1(
b101111101100100 +
b101111101100100 1
#816050000000
0#
0(
#816060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#816110000000
0$
0)
#816120000000
1"
1'
b0 +
b0 1
#816170000000
0"
0'
#816180000000
1#
1(
b101111101100100 +
b101111101100100 1
#816230000000
0#
0(
#816240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#816290000000
0$
0)
#816300000000
1"
1'
b0 +
b0 1
#816350000000
0"
0'
#816360000000
1#
1(
b101111101100100 +
b101111101100100 1
#816410000000
0#
0(
#816420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#816470000000
0$
0)
#816480000000
1"
1'
b0 +
b0 1
#816530000000
0"
0'
#816540000000
1#
1(
b101111101100100 +
b101111101100100 1
#816590000000
0#
0(
#816600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#816650000000
0$
0)
#816660000000
1"
1'
b0 +
b0 1
#816710000000
0"
0'
#816720000000
1#
1(
b101111101100100 +
b101111101100100 1
#816770000000
0#
0(
#816780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#816830000000
0$
0)
#816840000000
1"
1'
b0 +
b0 1
#816890000000
0"
0'
#816900000000
1#
1(
b101111101100100 +
b101111101100100 1
#816950000000
0#
0(
#816960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#817010000000
0$
0)
#817020000000
1"
1'
b0 +
b0 1
#817070000000
0"
0'
#817080000000
1#
1(
b101111101100100 +
b101111101100100 1
#817130000000
0#
0(
#817140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#817190000000
0$
0)
#817200000000
1"
1'
b0 +
b0 1
#817250000000
0"
0'
#817260000000
1#
1(
b101111101100100 +
b101111101100100 1
#817310000000
0#
0(
#817320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#817370000000
0$
0)
#817380000000
1"
1'
b0 +
b0 1
#817430000000
0"
0'
#817440000000
1#
1(
b101111101100100 +
b101111101100100 1
#817490000000
0#
0(
#817500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#817550000000
0$
0)
#817560000000
1"
1'
b0 +
b0 1
#817610000000
0"
0'
#817620000000
1#
1(
b101111101100100 +
b101111101100100 1
#817670000000
0#
0(
#817680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#817730000000
0$
0)
#817740000000
1"
1'
b0 +
b0 1
#817790000000
0"
0'
#817800000000
1#
1(
b101111101100100 +
b101111101100100 1
#817850000000
0#
0(
#817860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#817910000000
0$
0)
#817920000000
1"
1'
b0 +
b0 1
#817970000000
0"
0'
#817980000000
1#
1(
b101111101100100 +
b101111101100100 1
#818030000000
0#
0(
#818040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#818090000000
0$
0)
#818100000000
1"
1'
b0 +
b0 1
#818150000000
0"
0'
#818160000000
1#
1(
b101111101100100 +
b101111101100100 1
#818210000000
0#
0(
#818220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#818270000000
0$
0)
#818280000000
1"
1'
b0 +
b0 1
#818330000000
0"
0'
#818340000000
1#
1(
b101111101100100 +
b101111101100100 1
#818390000000
0#
0(
#818400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#818450000000
0$
0)
#818460000000
1"
1'
b0 +
b0 1
#818510000000
0"
0'
#818520000000
1#
1(
b101111101100100 +
b101111101100100 1
#818570000000
0#
0(
#818580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#818630000000
0$
0)
#818640000000
1"
1'
b0 +
b0 1
#818690000000
0"
0'
#818700000000
1#
1(
b101111101100100 +
b101111101100100 1
#818750000000
0#
0(
#818760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#818810000000
0$
0)
#818820000000
1"
1'
b0 +
b0 1
#818870000000
0"
0'
#818880000000
1#
1(
b101111101100100 +
b101111101100100 1
#818930000000
0#
0(
#818940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#818990000000
0$
0)
#819000000000
1"
1'
b0 +
b0 1
#819050000000
0"
0'
#819060000000
1#
1(
b101111101100100 +
b101111101100100 1
#819110000000
0#
0(
#819120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#819170000000
0$
0)
#819180000000
1"
1'
b0 +
b0 1
#819230000000
0"
0'
#819240000000
1#
1(
b101111101100100 +
b101111101100100 1
#819290000000
0#
0(
#819300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#819350000000
0$
0)
#819360000000
1"
1'
b0 +
b0 1
#819410000000
0"
0'
#819420000000
1#
1(
b101111101100100 +
b101111101100100 1
#819470000000
0#
0(
#819480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#819530000000
0$
0)
#819540000000
1"
1'
b0 +
b0 1
#819590000000
0"
0'
#819600000000
1#
1(
b101111101100100 +
b101111101100100 1
#819650000000
0#
0(
#819660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#819710000000
0$
0)
#819720000000
1"
1'
b0 +
b0 1
#819770000000
0"
0'
#819780000000
1#
1(
b101111101100100 +
b101111101100100 1
#819830000000
0#
0(
#819840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#819890000000
0$
0)
#819900000000
1"
1'
b0 +
b0 1
#819950000000
0"
0'
#819960000000
1#
1(
b101111101100100 +
b101111101100100 1
#820010000000
0#
0(
#820020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#820070000000
0$
0)
#820080000000
1"
1'
b0 +
b0 1
#820130000000
0"
0'
#820140000000
1#
1(
b101111101100100 +
b101111101100100 1
#820190000000
0#
0(
#820200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#820250000000
0$
0)
#820260000000
1"
1'
b0 +
b0 1
#820310000000
0"
0'
#820320000000
1#
1(
b101111101100100 +
b101111101100100 1
#820370000000
0#
0(
#820380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#820430000000
0$
0)
#820440000000
1"
1'
b0 +
b0 1
#820490000000
0"
0'
#820500000000
1#
1(
b101111101100100 +
b101111101100100 1
#820550000000
0#
0(
#820560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#820610000000
0$
0)
#820620000000
1"
1'
b0 +
b0 1
#820670000000
0"
0'
#820680000000
1#
1(
b101111101100100 +
b101111101100100 1
#820730000000
0#
0(
#820740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#820790000000
0$
0)
#820800000000
1"
1'
b0 +
b0 1
#820850000000
0"
0'
#820860000000
1#
1(
b101111101100100 +
b101111101100100 1
#820910000000
0#
0(
#820920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#820970000000
0$
0)
#820980000000
1"
1'
b0 +
b0 1
#821030000000
0"
0'
#821040000000
1#
1(
b101111101100100 +
b101111101100100 1
#821090000000
0#
0(
#821100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#821150000000
0$
0)
#821160000000
1"
1'
b0 +
b0 1
#821210000000
0"
0'
#821220000000
1#
1(
b101111101100100 +
b101111101100100 1
#821270000000
0#
0(
#821280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#821330000000
0$
0)
#821340000000
1"
1'
b0 +
b0 1
#821390000000
0"
0'
#821400000000
1#
1(
b101111101100100 +
b101111101100100 1
#821450000000
0#
0(
#821460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#821510000000
0$
0)
#821520000000
1"
1'
b0 +
b0 1
#821570000000
0"
0'
#821580000000
1#
1(
b101111101100100 +
b101111101100100 1
#821630000000
0#
0(
#821640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#821690000000
0$
0)
#821700000000
1"
1'
b0 +
b0 1
#821750000000
0"
0'
#821760000000
1#
1(
b101111101100100 +
b101111101100100 1
#821810000000
0#
0(
#821820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#821870000000
0$
0)
#821880000000
1"
1'
b0 +
b0 1
#821930000000
0"
0'
#821940000000
1#
1(
b101111101100100 +
b101111101100100 1
#821990000000
0#
0(
#822000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#822050000000
0$
0)
#822060000000
1"
1'
b0 +
b0 1
#822110000000
0"
0'
#822120000000
1#
1(
b101111101100100 +
b101111101100100 1
#822170000000
0#
0(
#822180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#822230000000
0$
0)
#822240000000
1"
1'
b0 +
b0 1
#822290000000
0"
0'
#822300000000
1#
1(
b101111101100100 +
b101111101100100 1
#822350000000
0#
0(
#822360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#822410000000
0$
0)
#822420000000
1"
1'
b0 +
b0 1
#822470000000
0"
0'
#822480000000
1#
1(
b101111101100100 +
b101111101100100 1
#822530000000
0#
0(
#822540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#822590000000
0$
0)
#822600000000
1"
1'
b0 +
b0 1
#822650000000
0"
0'
#822660000000
1#
1(
b101111101100100 +
b101111101100100 1
#822710000000
0#
0(
#822720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#822770000000
0$
0)
#822780000000
1"
1'
b0 +
b0 1
#822830000000
0"
0'
#822840000000
1#
1(
b101111101100100 +
b101111101100100 1
#822890000000
0#
0(
#822900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#822950000000
0$
0)
#822960000000
1"
1'
b0 +
b0 1
#823010000000
0"
0'
#823020000000
1#
1(
b101111101100100 +
b101111101100100 1
#823070000000
0#
0(
#823080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#823130000000
0$
0)
#823140000000
1"
1'
b0 +
b0 1
#823190000000
0"
0'
#823200000000
1#
1(
b101111101100100 +
b101111101100100 1
#823250000000
0#
0(
#823260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#823310000000
0$
0)
#823320000000
1"
1'
b0 +
b0 1
#823370000000
0"
0'
#823380000000
1#
1(
b101111101100100 +
b101111101100100 1
#823430000000
0#
0(
#823440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#823490000000
0$
0)
#823500000000
1"
1'
b0 +
b0 1
#823550000000
0"
0'
#823560000000
1#
1(
b101111101100100 +
b101111101100100 1
#823610000000
0#
0(
#823620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#823670000000
0$
0)
#823680000000
1"
1'
b0 +
b0 1
#823730000000
0"
0'
#823740000000
1#
1(
b101111101100100 +
b101111101100100 1
#823790000000
0#
0(
#823800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#823850000000
0$
0)
#823860000000
1"
1'
b0 +
b0 1
#823910000000
0"
0'
#823920000000
1#
1(
b101111101100100 +
b101111101100100 1
#823970000000
0#
0(
#823980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#824030000000
0$
0)
#824040000000
1"
1'
b0 +
b0 1
#824090000000
0"
0'
#824100000000
1#
1(
b101111101100100 +
b101111101100100 1
#824150000000
0#
0(
#824160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#824210000000
0$
0)
#824220000000
1"
1'
b0 +
b0 1
#824270000000
0"
0'
#824280000000
1#
1(
b101111101100100 +
b101111101100100 1
#824330000000
0#
0(
#824340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#824390000000
0$
0)
#824400000000
1"
1'
b0 +
b0 1
#824450000000
0"
0'
#824460000000
1#
1(
b101111101100100 +
b101111101100100 1
#824510000000
0#
0(
#824520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#824570000000
0$
0)
#824580000000
1"
1'
b0 +
b0 1
#824630000000
0"
0'
#824640000000
1#
1(
b101111101100100 +
b101111101100100 1
#824690000000
0#
0(
#824700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#824750000000
0$
0)
#824760000000
1"
1'
b0 +
b0 1
#824810000000
0"
0'
#824820000000
1#
1(
b101111101100100 +
b101111101100100 1
#824870000000
0#
0(
#824880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#824930000000
0$
0)
#824940000000
1"
1'
b0 +
b0 1
#824990000000
0"
0'
#825000000000
1#
1(
b101111101100100 +
b101111101100100 1
#825050000000
0#
0(
#825060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#825110000000
0$
0)
#825120000000
1"
1'
b0 +
b0 1
#825170000000
0"
0'
#825180000000
1#
1(
b101111101100100 +
b101111101100100 1
#825230000000
0#
0(
#825240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#825290000000
0$
0)
#825300000000
1"
1'
b0 +
b0 1
#825350000000
0"
0'
#825360000000
1#
1(
b101111101100100 +
b101111101100100 1
#825410000000
0#
0(
#825420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#825470000000
0$
0)
#825480000000
1"
1'
b0 +
b0 1
#825530000000
0"
0'
#825540000000
1#
1(
b101111101100100 +
b101111101100100 1
#825590000000
0#
0(
#825600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#825650000000
0$
0)
#825660000000
1"
1'
b0 +
b0 1
#825710000000
0"
0'
#825720000000
1#
1(
b101111101100100 +
b101111101100100 1
#825770000000
0#
0(
#825780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#825830000000
0$
0)
#825840000000
1"
1'
b0 +
b0 1
#825890000000
0"
0'
#825900000000
1#
1(
b101111101100100 +
b101111101100100 1
#825950000000
0#
0(
#825960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#826010000000
0$
0)
#826020000000
1"
1'
b0 +
b0 1
#826070000000
0"
0'
#826080000000
1#
1(
b101111101100100 +
b101111101100100 1
#826130000000
0#
0(
#826140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#826190000000
0$
0)
#826200000000
1"
1'
b0 +
b0 1
#826250000000
0"
0'
#826260000000
1#
1(
b101111101100100 +
b101111101100100 1
#826310000000
0#
0(
#826320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#826370000000
0$
0)
#826380000000
1"
1'
b0 +
b0 1
#826430000000
0"
0'
#826440000000
1#
1(
b101111101100100 +
b101111101100100 1
#826490000000
0#
0(
#826500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#826550000000
0$
0)
#826560000000
1"
1'
b0 +
b0 1
#826610000000
0"
0'
#826620000000
1#
1(
b101111101100100 +
b101111101100100 1
#826670000000
0#
0(
#826680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#826730000000
0$
0)
#826740000000
1"
1'
b0 +
b0 1
#826790000000
0"
0'
#826800000000
1#
1(
b101111101100100 +
b101111101100100 1
#826850000000
0#
0(
#826860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#826910000000
0$
0)
#826920000000
1"
1'
b0 +
b0 1
#826970000000
0"
0'
#826980000000
1#
1(
b101111101100100 +
b101111101100100 1
#827030000000
0#
0(
#827040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#827090000000
0$
0)
#827100000000
1"
1'
b0 +
b0 1
#827150000000
0"
0'
#827160000000
1#
1(
b101111101100100 +
b101111101100100 1
#827210000000
0#
0(
#827220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#827270000000
0$
0)
#827280000000
1"
1'
b0 +
b0 1
#827330000000
0"
0'
#827340000000
1#
1(
b101111101100100 +
b101111101100100 1
#827390000000
0#
0(
#827400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#827450000000
0$
0)
#827460000000
1"
1'
b0 +
b0 1
#827510000000
0"
0'
#827520000000
1#
1(
b101111101100100 +
b101111101100100 1
#827570000000
0#
0(
#827580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#827630000000
0$
0)
#827640000000
1"
1'
b0 +
b0 1
#827690000000
0"
0'
#827700000000
1#
1(
b101111101100100 +
b101111101100100 1
#827750000000
0#
0(
#827760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#827810000000
0$
0)
#827820000000
1"
1'
b0 +
b0 1
#827870000000
0"
0'
#827880000000
1#
1(
b101111101100100 +
b101111101100100 1
#827930000000
0#
0(
#827940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#827990000000
0$
0)
#828000000000
1"
1'
b0 +
b0 1
#828050000000
0"
0'
#828060000000
1#
1(
b101111101100100 +
b101111101100100 1
#828110000000
0#
0(
#828120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#828170000000
0$
0)
#828180000000
1"
1'
b0 +
b0 1
#828230000000
0"
0'
#828240000000
1#
1(
b101111101100100 +
b101111101100100 1
#828290000000
0#
0(
#828300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#828350000000
0$
0)
#828360000000
1"
1'
b0 +
b0 1
#828410000000
0"
0'
#828420000000
1#
1(
b101111101100100 +
b101111101100100 1
#828470000000
0#
0(
#828480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#828530000000
0$
0)
#828540000000
1"
1'
b0 +
b0 1
#828590000000
0"
0'
#828600000000
1#
1(
b101111101100100 +
b101111101100100 1
#828650000000
0#
0(
#828660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#828710000000
0$
0)
#828720000000
1"
1'
b0 +
b0 1
#828770000000
0"
0'
#828780000000
1#
1(
b101111101100100 +
b101111101100100 1
#828830000000
0#
0(
#828840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#828890000000
0$
0)
#828900000000
1"
1'
b0 +
b0 1
#828950000000
0"
0'
#828960000000
1#
1(
b101111101100100 +
b101111101100100 1
#829010000000
0#
0(
#829020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#829070000000
0$
0)
#829080000000
1"
1'
b0 +
b0 1
#829130000000
0"
0'
#829140000000
1#
1(
b101111101100100 +
b101111101100100 1
#829190000000
0#
0(
#829200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#829250000000
0$
0)
#829260000000
1"
1'
b0 +
b0 1
#829310000000
0"
0'
#829320000000
1#
1(
b101111101100100 +
b101111101100100 1
#829370000000
0#
0(
#829380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#829430000000
0$
0)
#829440000000
1"
1'
b0 +
b0 1
#829490000000
0"
0'
#829500000000
1#
1(
b101111101100100 +
b101111101100100 1
#829550000000
0#
0(
#829560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#829610000000
0$
0)
#829620000000
1"
1'
b0 +
b0 1
#829670000000
0"
0'
#829680000000
1#
1(
b101111101100100 +
b101111101100100 1
#829730000000
0#
0(
#829740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#829790000000
0$
0)
#829800000000
1"
1'
b0 +
b0 1
#829850000000
0"
0'
#829860000000
1#
1(
b101111101100100 +
b101111101100100 1
#829910000000
0#
0(
#829920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#829970000000
0$
0)
#829980000000
1"
1'
b0 +
b0 1
#830030000000
0"
0'
#830040000000
1#
1(
b101111101100100 +
b101111101100100 1
#830090000000
0#
0(
#830100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#830150000000
0$
0)
#830160000000
1"
1'
b0 +
b0 1
#830210000000
0"
0'
#830220000000
1#
1(
b101111101100100 +
b101111101100100 1
#830270000000
0#
0(
#830280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#830330000000
0$
0)
#830340000000
1"
1'
b0 +
b0 1
#830390000000
0"
0'
#830400000000
1#
1(
b101111101100100 +
b101111101100100 1
#830450000000
0#
0(
#830460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#830510000000
0$
0)
#830520000000
1"
1'
b0 +
b0 1
#830570000000
0"
0'
#830580000000
1#
1(
b101111101100100 +
b101111101100100 1
#830630000000
0#
0(
#830640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#830690000000
0$
0)
#830700000000
1"
1'
b0 +
b0 1
#830750000000
0"
0'
#830760000000
1#
1(
b101111101100100 +
b101111101100100 1
#830810000000
0#
0(
#830820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#830870000000
0$
0)
#830880000000
1"
1'
b0 +
b0 1
#830930000000
0"
0'
#830940000000
1#
1(
b101111101100100 +
b101111101100100 1
#830990000000
0#
0(
#831000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#831050000000
0$
0)
#831060000000
1"
1'
b0 +
b0 1
#831110000000
0"
0'
#831120000000
1#
1(
b101111101100100 +
b101111101100100 1
#831170000000
0#
0(
#831180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#831230000000
0$
0)
#831240000000
1"
1'
b0 +
b0 1
#831290000000
0"
0'
#831300000000
1#
1(
b101111101100100 +
b101111101100100 1
#831350000000
0#
0(
#831360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#831410000000
0$
0)
#831420000000
1"
1'
b0 +
b0 1
#831470000000
0"
0'
#831480000000
1#
1(
b101111101100100 +
b101111101100100 1
#831530000000
0#
0(
#831540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#831590000000
0$
0)
#831600000000
1"
1'
b0 +
b0 1
#831650000000
0"
0'
#831660000000
1#
1(
b101111101100100 +
b101111101100100 1
#831710000000
0#
0(
#831720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#831770000000
0$
0)
#831780000000
1"
1'
b0 +
b0 1
#831830000000
0"
0'
#831840000000
1#
1(
b101111101100100 +
b101111101100100 1
#831890000000
0#
0(
#831900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#831950000000
0$
0)
#831960000000
1"
1'
b0 +
b0 1
#832010000000
0"
0'
#832020000000
1#
1(
b101111101100100 +
b101111101100100 1
#832070000000
0#
0(
#832080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#832130000000
0$
0)
#832140000000
1"
1'
b0 +
b0 1
#832190000000
0"
0'
#832200000000
1#
1(
b101111101100100 +
b101111101100100 1
#832250000000
0#
0(
#832260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#832310000000
0$
0)
#832320000000
1"
1'
b0 +
b0 1
#832370000000
0"
0'
#832380000000
1#
1(
b101111101100100 +
b101111101100100 1
#832430000000
0#
0(
#832440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#832490000000
0$
0)
#832500000000
1"
1'
b0 +
b0 1
#832550000000
0"
0'
#832560000000
1#
1(
b101111101100100 +
b101111101100100 1
#832610000000
0#
0(
#832620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#832670000000
0$
0)
#832680000000
1"
1'
b0 +
b0 1
#832730000000
0"
0'
#832740000000
1#
1(
b101111101100100 +
b101111101100100 1
#832790000000
0#
0(
#832800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#832850000000
0$
0)
#832860000000
1"
1'
b0 +
b0 1
#832910000000
0"
0'
#832920000000
1#
1(
b101111101100100 +
b101111101100100 1
#832970000000
0#
0(
#832980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#833030000000
0$
0)
#833040000000
1"
1'
b0 +
b0 1
#833090000000
0"
0'
#833100000000
1#
1(
b101111101100100 +
b101111101100100 1
#833150000000
0#
0(
#833160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#833210000000
0$
0)
#833220000000
1"
1'
b0 +
b0 1
#833270000000
0"
0'
#833280000000
1#
1(
b101111101100100 +
b101111101100100 1
#833330000000
0#
0(
#833340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#833390000000
0$
0)
#833400000000
1"
1'
b0 +
b0 1
#833450000000
0"
0'
#833460000000
1#
1(
b101111101100100 +
b101111101100100 1
#833510000000
0#
0(
#833520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#833570000000
0$
0)
#833580000000
1"
1'
b0 +
b0 1
#833630000000
0"
0'
#833640000000
1#
1(
b101111101100100 +
b101111101100100 1
#833690000000
0#
0(
#833700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#833750000000
0$
0)
#833760000000
1"
1'
b0 +
b0 1
#833810000000
0"
0'
#833820000000
1#
1(
b101111101100100 +
b101111101100100 1
#833870000000
0#
0(
#833880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#833930000000
0$
0)
#833940000000
1"
1'
b0 +
b0 1
#833990000000
0"
0'
#834000000000
1#
1(
b101111101100100 +
b101111101100100 1
#834050000000
0#
0(
#834060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#834110000000
0$
0)
#834120000000
1"
1'
b0 +
b0 1
#834170000000
0"
0'
#834180000000
1#
1(
b101111101100100 +
b101111101100100 1
#834230000000
0#
0(
#834240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#834290000000
0$
0)
#834300000000
1"
1'
b0 +
b0 1
#834350000000
0"
0'
#834360000000
1#
1(
b101111101100100 +
b101111101100100 1
#834410000000
0#
0(
#834420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#834470000000
0$
0)
#834480000000
1"
1'
b0 +
b0 1
#834530000000
0"
0'
#834540000000
1#
1(
b101111101100100 +
b101111101100100 1
#834590000000
0#
0(
#834600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#834650000000
0$
0)
#834660000000
1"
1'
b0 +
b0 1
#834710000000
0"
0'
#834720000000
1#
1(
b101111101100100 +
b101111101100100 1
#834770000000
0#
0(
#834780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#834830000000
0$
0)
#834840000000
1"
1'
b0 +
b0 1
#834890000000
0"
0'
#834900000000
1#
1(
b101111101100100 +
b101111101100100 1
#834950000000
0#
0(
#834960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#835010000000
0$
0)
#835020000000
1"
1'
b0 +
b0 1
#835070000000
0"
0'
#835080000000
1#
1(
b101111101100100 +
b101111101100100 1
#835130000000
0#
0(
#835140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#835190000000
0$
0)
#835200000000
1"
1'
b0 +
b0 1
#835250000000
0"
0'
#835260000000
1#
1(
b101111101100100 +
b101111101100100 1
#835310000000
0#
0(
#835320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#835370000000
0$
0)
#835380000000
1"
1'
b0 +
b0 1
#835430000000
0"
0'
#835440000000
1#
1(
b101111101100100 +
b101111101100100 1
#835490000000
0#
0(
#835500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#835550000000
0$
0)
#835560000000
1"
1'
b0 +
b0 1
#835610000000
0"
0'
#835620000000
1#
1(
b101111101100100 +
b101111101100100 1
#835670000000
0#
0(
#835680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#835730000000
0$
0)
#835740000000
1"
1'
b0 +
b0 1
#835790000000
0"
0'
#835800000000
1#
1(
b101111101100100 +
b101111101100100 1
#835850000000
0#
0(
#835860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#835910000000
0$
0)
#835920000000
1"
1'
b0 +
b0 1
#835970000000
0"
0'
#835980000000
1#
1(
b101111101100100 +
b101111101100100 1
#836030000000
0#
0(
#836040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#836090000000
0$
0)
#836100000000
1"
1'
b0 +
b0 1
#836150000000
0"
0'
#836160000000
1#
1(
b101111101100100 +
b101111101100100 1
#836210000000
0#
0(
#836220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#836270000000
0$
0)
#836280000000
1"
1'
b0 +
b0 1
#836330000000
0"
0'
#836340000000
1#
1(
b101111101100100 +
b101111101100100 1
#836390000000
0#
0(
#836400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#836450000000
0$
0)
#836460000000
1"
1'
b0 +
b0 1
#836510000000
0"
0'
#836520000000
1#
1(
b101111101100100 +
b101111101100100 1
#836570000000
0#
0(
#836580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#836630000000
0$
0)
#836640000000
1"
1'
b0 +
b0 1
#836690000000
0"
0'
#836700000000
1#
1(
b101111101100100 +
b101111101100100 1
#836750000000
0#
0(
#836760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#836810000000
0$
0)
#836820000000
1"
1'
b0 +
b0 1
#836870000000
0"
0'
#836880000000
1#
1(
b101111101100100 +
b101111101100100 1
#836930000000
0#
0(
#836940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#836990000000
0$
0)
#837000000000
1"
1'
b0 +
b0 1
#837050000000
0"
0'
#837060000000
1#
1(
b101111101100100 +
b101111101100100 1
#837110000000
0#
0(
#837120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#837170000000
0$
0)
#837180000000
1"
1'
b0 +
b0 1
#837230000000
0"
0'
#837240000000
1#
1(
b101111101100100 +
b101111101100100 1
#837290000000
0#
0(
#837300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#837350000000
0$
0)
#837360000000
1"
1'
b0 +
b0 1
#837410000000
0"
0'
#837420000000
1#
1(
b101111101100100 +
b101111101100100 1
#837470000000
0#
0(
#837480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#837530000000
0$
0)
#837540000000
1"
1'
b0 +
b0 1
#837590000000
0"
0'
#837600000000
1#
1(
b101111101100100 +
b101111101100100 1
#837650000000
0#
0(
#837660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#837710000000
0$
0)
#837720000000
1"
1'
b0 +
b0 1
#837770000000
0"
0'
#837780000000
1#
1(
b101111101100100 +
b101111101100100 1
#837830000000
0#
0(
#837840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#837890000000
0$
0)
#837900000000
1"
1'
b0 +
b0 1
#837950000000
0"
0'
#837960000000
1#
1(
b101111101100100 +
b101111101100100 1
#838010000000
0#
0(
#838020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#838070000000
0$
0)
#838080000000
1"
1'
b0 +
b0 1
#838130000000
0"
0'
#838140000000
1#
1(
b101111101100100 +
b101111101100100 1
#838190000000
0#
0(
#838200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#838250000000
0$
0)
#838260000000
1"
1'
b0 +
b0 1
#838310000000
0"
0'
#838320000000
1#
1(
b101111101100100 +
b101111101100100 1
#838370000000
0#
0(
#838380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#838430000000
0$
0)
#838440000000
1"
1'
b0 +
b0 1
#838490000000
0"
0'
#838500000000
1#
1(
b101111101100100 +
b101111101100100 1
#838550000000
0#
0(
#838560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#838610000000
0$
0)
#838620000000
1"
1'
b0 +
b0 1
#838670000000
0"
0'
#838680000000
1#
1(
b101111101100100 +
b101111101100100 1
#838730000000
0#
0(
#838740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#838790000000
0$
0)
#838800000000
1"
1'
b0 +
b0 1
#838850000000
0"
0'
#838860000000
1#
1(
b101111101100100 +
b101111101100100 1
#838910000000
0#
0(
#838920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#838970000000
0$
0)
#838980000000
1"
1'
b0 +
b0 1
#839030000000
0"
0'
#839040000000
1#
1(
b101111101100100 +
b101111101100100 1
#839090000000
0#
0(
#839100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#839150000000
0$
0)
#839160000000
1"
1'
b0 +
b0 1
#839210000000
0"
0'
#839220000000
1#
1(
b101111101100100 +
b101111101100100 1
#839270000000
0#
0(
#839280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#839330000000
0$
0)
#839340000000
1"
1'
b0 +
b0 1
#839390000000
0"
0'
#839400000000
1#
1(
b101111101100100 +
b101111101100100 1
#839450000000
0#
0(
#839460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#839510000000
0$
0)
#839520000000
1"
1'
b0 +
b0 1
#839570000000
0"
0'
#839580000000
1#
1(
b101111101100100 +
b101111101100100 1
#839630000000
0#
0(
#839640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#839690000000
0$
0)
#839700000000
1"
1'
b0 +
b0 1
#839750000000
0"
0'
#839760000000
1#
1(
b101111101100100 +
b101111101100100 1
#839810000000
0#
0(
#839820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#839870000000
0$
0)
#839880000000
1"
1'
b0 +
b0 1
#839930000000
0"
0'
#839940000000
1#
1(
b101111101100100 +
b101111101100100 1
#839990000000
0#
0(
#840000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#840050000000
0$
0)
#840060000000
1"
1'
b0 +
b0 1
#840110000000
0"
0'
#840120000000
1#
1(
b101111101100100 +
b101111101100100 1
#840170000000
0#
0(
#840180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#840230000000
0$
0)
#840240000000
1"
1'
b0 +
b0 1
#840290000000
0"
0'
#840300000000
1#
1(
b101111101100100 +
b101111101100100 1
#840350000000
0#
0(
#840360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#840410000000
0$
0)
#840420000000
1"
1'
b0 +
b0 1
#840470000000
0"
0'
#840480000000
1#
1(
b101111101100100 +
b101111101100100 1
#840530000000
0#
0(
#840540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#840590000000
0$
0)
#840600000000
1"
1'
b0 +
b0 1
#840650000000
0"
0'
#840660000000
1#
1(
b101111101100100 +
b101111101100100 1
#840710000000
0#
0(
#840720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#840770000000
0$
0)
#840780000000
1"
1'
b0 +
b0 1
#840830000000
0"
0'
#840840000000
1#
1(
b101111101100100 +
b101111101100100 1
#840890000000
0#
0(
#840900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#840950000000
0$
0)
#840960000000
1"
1'
b0 +
b0 1
#841010000000
0"
0'
#841020000000
1#
1(
b101111101100100 +
b101111101100100 1
#841070000000
0#
0(
#841080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#841130000000
0$
0)
#841140000000
1"
1'
b0 +
b0 1
#841190000000
0"
0'
#841200000000
1#
1(
b101111101100100 +
b101111101100100 1
#841250000000
0#
0(
#841260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#841310000000
0$
0)
#841320000000
1"
1'
b0 +
b0 1
#841370000000
0"
0'
#841380000000
1#
1(
b101111101100100 +
b101111101100100 1
#841430000000
0#
0(
#841440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#841490000000
0$
0)
#841500000000
1"
1'
b0 +
b0 1
#841550000000
0"
0'
#841560000000
1#
1(
b101111101100100 +
b101111101100100 1
#841610000000
0#
0(
#841620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#841670000000
0$
0)
#841680000000
1"
1'
b0 +
b0 1
#841730000000
0"
0'
#841740000000
1#
1(
b101111101100100 +
b101111101100100 1
#841790000000
0#
0(
#841800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#841850000000
0$
0)
#841860000000
1"
1'
b0 +
b0 1
#841910000000
0"
0'
#841920000000
1#
1(
b101111101100100 +
b101111101100100 1
#841970000000
0#
0(
#841980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#842030000000
0$
0)
#842040000000
1"
1'
b0 +
b0 1
#842090000000
0"
0'
#842100000000
1#
1(
b101111101100100 +
b101111101100100 1
#842150000000
0#
0(
#842160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#842210000000
0$
0)
#842220000000
1"
1'
b0 +
b0 1
#842270000000
0"
0'
#842280000000
1#
1(
b101111101100100 +
b101111101100100 1
#842330000000
0#
0(
#842340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#842390000000
0$
0)
#842400000000
1"
1'
b0 +
b0 1
#842450000000
0"
0'
#842460000000
1#
1(
b101111101100100 +
b101111101100100 1
#842510000000
0#
0(
#842520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#842570000000
0$
0)
#842580000000
1"
1'
b0 +
b0 1
#842630000000
0"
0'
#842640000000
1#
1(
b101111101100100 +
b101111101100100 1
#842690000000
0#
0(
#842700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#842750000000
0$
0)
#842760000000
1"
1'
b0 +
b0 1
#842810000000
0"
0'
#842820000000
1#
1(
b101111101100100 +
b101111101100100 1
#842870000000
0#
0(
#842880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#842930000000
0$
0)
#842940000000
1"
1'
b0 +
b0 1
#842990000000
0"
0'
#843000000000
1#
1(
b101111101100100 +
b101111101100100 1
#843050000000
0#
0(
#843060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#843110000000
0$
0)
#843120000000
1"
1'
b0 +
b0 1
#843170000000
0"
0'
#843180000000
1#
1(
b101111101100100 +
b101111101100100 1
#843230000000
0#
0(
#843240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#843290000000
0$
0)
#843300000000
1"
1'
b0 +
b0 1
#843350000000
0"
0'
#843360000000
1#
1(
b101111101100100 +
b101111101100100 1
#843410000000
0#
0(
#843420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#843470000000
0$
0)
#843480000000
1"
1'
b0 +
b0 1
#843530000000
0"
0'
#843540000000
1#
1(
b101111101100100 +
b101111101100100 1
#843590000000
0#
0(
#843600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#843650000000
0$
0)
#843660000000
1"
1'
b0 +
b0 1
#843710000000
0"
0'
#843720000000
1#
1(
b101111101100100 +
b101111101100100 1
#843770000000
0#
0(
#843780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#843830000000
0$
0)
#843840000000
1"
1'
b0 +
b0 1
#843890000000
0"
0'
#843900000000
1#
1(
b101111101100100 +
b101111101100100 1
#843950000000
0#
0(
#843960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#844010000000
0$
0)
#844020000000
1"
1'
b0 +
b0 1
#844070000000
0"
0'
#844080000000
1#
1(
b101111101100100 +
b101111101100100 1
#844130000000
0#
0(
#844140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#844190000000
0$
0)
#844200000000
1"
1'
b0 +
b0 1
#844250000000
0"
0'
#844260000000
1#
1(
b101111101100100 +
b101111101100100 1
#844310000000
0#
0(
#844320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#844370000000
0$
0)
#844380000000
1"
1'
b0 +
b0 1
#844430000000
0"
0'
#844440000000
1#
1(
b101111101100100 +
b101111101100100 1
#844490000000
0#
0(
#844500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#844550000000
0$
0)
#844560000000
1"
1'
b0 +
b0 1
#844610000000
0"
0'
#844620000000
1#
1(
b101111101100100 +
b101111101100100 1
#844670000000
0#
0(
#844680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#844730000000
0$
0)
#844740000000
1"
1'
b0 +
b0 1
#844790000000
0"
0'
#844800000000
1#
1(
b101111101100100 +
b101111101100100 1
#844850000000
0#
0(
#844860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#844910000000
0$
0)
#844920000000
1"
1'
b0 +
b0 1
#844970000000
0"
0'
#844980000000
1#
1(
b101111101100100 +
b101111101100100 1
#845030000000
0#
0(
#845040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#845090000000
0$
0)
#845100000000
1"
1'
b0 +
b0 1
#845150000000
0"
0'
#845160000000
1#
1(
b101111101100100 +
b101111101100100 1
#845210000000
0#
0(
#845220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#845270000000
0$
0)
#845280000000
1"
1'
b0 +
b0 1
#845330000000
0"
0'
#845340000000
1#
1(
b101111101100100 +
b101111101100100 1
#845390000000
0#
0(
#845400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#845450000000
0$
0)
#845460000000
1"
1'
b0 +
b0 1
#845510000000
0"
0'
#845520000000
1#
1(
b101111101100100 +
b101111101100100 1
#845570000000
0#
0(
#845580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#845630000000
0$
0)
#845640000000
1"
1'
b0 +
b0 1
#845690000000
0"
0'
#845700000000
1#
1(
b101111101100100 +
b101111101100100 1
#845750000000
0#
0(
#845760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#845810000000
0$
0)
#845820000000
1"
1'
b0 +
b0 1
#845870000000
0"
0'
#845880000000
1#
1(
b101111101100100 +
b101111101100100 1
#845930000000
0#
0(
#845940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#845990000000
0$
0)
#846000000000
1"
1'
b0 +
b0 1
#846050000000
0"
0'
#846060000000
1#
1(
b101111101100100 +
b101111101100100 1
#846110000000
0#
0(
#846120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#846170000000
0$
0)
#846180000000
1"
1'
b0 +
b0 1
#846230000000
0"
0'
#846240000000
1#
1(
b101111101100100 +
b101111101100100 1
#846290000000
0#
0(
#846300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#846350000000
0$
0)
#846360000000
1"
1'
b0 +
b0 1
#846410000000
0"
0'
#846420000000
1#
1(
b101111101100100 +
b101111101100100 1
#846470000000
0#
0(
#846480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#846530000000
0$
0)
#846540000000
1"
1'
b0 +
b0 1
#846590000000
0"
0'
#846600000000
1#
1(
b101111101100100 +
b101111101100100 1
#846650000000
0#
0(
#846660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#846710000000
0$
0)
#846720000000
1"
1'
b0 +
b0 1
#846770000000
0"
0'
#846780000000
1#
1(
b101111101100100 +
b101111101100100 1
#846830000000
0#
0(
#846840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#846890000000
0$
0)
#846900000000
1"
1'
b0 +
b0 1
#846950000000
0"
0'
#846960000000
1#
1(
b101111101100100 +
b101111101100100 1
#847010000000
0#
0(
#847020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#847070000000
0$
0)
#847080000000
1"
1'
b0 +
b0 1
#847130000000
0"
0'
#847140000000
1#
1(
b101111101100100 +
b101111101100100 1
#847190000000
0#
0(
#847200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#847250000000
0$
0)
#847260000000
1"
1'
b0 +
b0 1
#847310000000
0"
0'
#847320000000
1#
1(
b101111101100100 +
b101111101100100 1
#847370000000
0#
0(
#847380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#847430000000
0$
0)
#847440000000
1"
1'
b0 +
b0 1
#847490000000
0"
0'
#847500000000
1#
1(
b101111101100100 +
b101111101100100 1
#847550000000
0#
0(
#847560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#847610000000
0$
0)
#847620000000
1"
1'
b0 +
b0 1
#847670000000
0"
0'
#847680000000
1#
1(
b101111101100100 +
b101111101100100 1
#847730000000
0#
0(
#847740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#847790000000
0$
0)
#847800000000
1"
1'
b0 +
b0 1
#847850000000
0"
0'
#847860000000
1#
1(
b101111101100100 +
b101111101100100 1
#847910000000
0#
0(
#847920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#847970000000
0$
0)
#847980000000
1"
1'
b0 +
b0 1
#848030000000
0"
0'
#848040000000
1#
1(
b101111101100100 +
b101111101100100 1
#848090000000
0#
0(
#848100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#848150000000
0$
0)
#848160000000
1"
1'
b0 +
b0 1
#848210000000
0"
0'
#848220000000
1#
1(
b101111101100100 +
b101111101100100 1
#848270000000
0#
0(
#848280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#848330000000
0$
0)
#848340000000
1"
1'
b0 +
b0 1
#848390000000
0"
0'
#848400000000
1#
1(
b101111101100100 +
b101111101100100 1
#848450000000
0#
0(
#848460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#848510000000
0$
0)
#848520000000
1"
1'
b0 +
b0 1
#848570000000
0"
0'
#848580000000
1#
1(
b101111101100100 +
b101111101100100 1
#848630000000
0#
0(
#848640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#848690000000
0$
0)
#848700000000
1"
1'
b0 +
b0 1
#848750000000
0"
0'
#848760000000
1#
1(
b101111101100100 +
b101111101100100 1
#848810000000
0#
0(
#848820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#848870000000
0$
0)
#848880000000
1"
1'
b0 +
b0 1
#848930000000
0"
0'
#848940000000
1#
1(
b101111101100100 +
b101111101100100 1
#848990000000
0#
0(
#849000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#849050000000
0$
0)
#849060000000
1"
1'
b0 +
b0 1
#849110000000
0"
0'
#849120000000
1#
1(
b101111101100100 +
b101111101100100 1
#849170000000
0#
0(
#849180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#849230000000
0$
0)
#849240000000
1"
1'
b0 +
b0 1
#849290000000
0"
0'
#849300000000
1#
1(
b101111101100100 +
b101111101100100 1
#849350000000
0#
0(
#849360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#849410000000
0$
0)
#849420000000
1"
1'
b0 +
b0 1
#849470000000
0"
0'
#849480000000
1#
1(
b101111101100100 +
b101111101100100 1
#849530000000
0#
0(
#849540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#849590000000
0$
0)
#849600000000
1"
1'
b0 +
b0 1
#849650000000
0"
0'
#849660000000
1#
1(
b101111101100100 +
b101111101100100 1
#849710000000
0#
0(
#849720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#849770000000
0$
0)
#849780000000
1"
1'
b0 +
b0 1
#849830000000
0"
0'
#849840000000
1#
1(
b101111101100100 +
b101111101100100 1
#849890000000
0#
0(
#849900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#849950000000
0$
0)
#849960000000
1"
1'
b0 +
b0 1
#850010000000
0"
0'
#850020000000
1#
1(
b101111101100100 +
b101111101100100 1
#850070000000
0#
0(
#850080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#850130000000
0$
0)
#850140000000
1"
1'
b0 +
b0 1
#850190000000
0"
0'
#850200000000
1#
1(
b101111101100100 +
b101111101100100 1
#850250000000
0#
0(
#850260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#850310000000
0$
0)
#850320000000
1"
1'
b0 +
b0 1
#850370000000
0"
0'
#850380000000
1#
1(
b101111101100100 +
b101111101100100 1
#850430000000
0#
0(
#850440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#850490000000
0$
0)
#850500000000
1"
1'
b0 +
b0 1
#850550000000
0"
0'
#850560000000
1#
1(
b101111101100100 +
b101111101100100 1
#850610000000
0#
0(
#850620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#850670000000
0$
0)
#850680000000
1"
1'
b0 +
b0 1
#850730000000
0"
0'
#850740000000
1#
1(
b101111101100100 +
b101111101100100 1
#850790000000
0#
0(
#850800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#850850000000
0$
0)
#850860000000
1"
1'
b0 +
b0 1
#850910000000
0"
0'
#850920000000
1#
1(
b101111101100100 +
b101111101100100 1
#850970000000
0#
0(
#850980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#851030000000
0$
0)
#851040000000
1"
1'
b0 +
b0 1
#851090000000
0"
0'
#851100000000
1#
1(
b101111101100100 +
b101111101100100 1
#851150000000
0#
0(
#851160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#851210000000
0$
0)
#851220000000
1"
1'
b0 +
b0 1
#851270000000
0"
0'
#851280000000
1#
1(
b101111101100100 +
b101111101100100 1
#851330000000
0#
0(
#851340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#851390000000
0$
0)
#851400000000
1"
1'
b0 +
b0 1
#851450000000
0"
0'
#851460000000
1#
1(
b101111101100100 +
b101111101100100 1
#851510000000
0#
0(
#851520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#851570000000
0$
0)
#851580000000
1"
1'
b0 +
b0 1
#851630000000
0"
0'
#851640000000
1#
1(
b101111101100100 +
b101111101100100 1
#851690000000
0#
0(
#851700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#851750000000
0$
0)
#851760000000
1"
1'
b0 +
b0 1
#851810000000
0"
0'
#851820000000
1#
1(
b101111101100100 +
b101111101100100 1
#851870000000
0#
0(
#851880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#851930000000
0$
0)
#851940000000
1"
1'
b0 +
b0 1
#851990000000
0"
0'
#852000000000
1#
1(
b101111101100100 +
b101111101100100 1
#852050000000
0#
0(
#852060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#852110000000
0$
0)
#852120000000
1"
1'
b0 +
b0 1
#852170000000
0"
0'
#852180000000
1#
1(
b101111101100100 +
b101111101100100 1
#852230000000
0#
0(
#852240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#852290000000
0$
0)
#852300000000
1"
1'
b0 +
b0 1
#852350000000
0"
0'
#852360000000
1#
1(
b101111101100100 +
b101111101100100 1
#852410000000
0#
0(
#852420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#852470000000
0$
0)
#852480000000
1"
1'
b0 +
b0 1
#852530000000
0"
0'
#852540000000
1#
1(
b101111101100100 +
b101111101100100 1
#852590000000
0#
0(
#852600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#852650000000
0$
0)
#852660000000
1"
1'
b0 +
b0 1
#852710000000
0"
0'
#852720000000
1#
1(
b101111101100100 +
b101111101100100 1
#852770000000
0#
0(
#852780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#852830000000
0$
0)
#852840000000
1"
1'
b0 +
b0 1
#852890000000
0"
0'
#852900000000
1#
1(
b101111101100100 +
b101111101100100 1
#852950000000
0#
0(
#852960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#853010000000
0$
0)
#853020000000
1"
1'
b0 +
b0 1
#853070000000
0"
0'
#853080000000
1#
1(
b101111101100100 +
b101111101100100 1
#853130000000
0#
0(
#853140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#853190000000
0$
0)
#853200000000
1"
1'
b0 +
b0 1
#853250000000
0"
0'
#853260000000
1#
1(
b101111101100100 +
b101111101100100 1
#853310000000
0#
0(
#853320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#853370000000
0$
0)
#853380000000
1"
1'
b0 +
b0 1
#853430000000
0"
0'
#853440000000
1#
1(
b101111101100100 +
b101111101100100 1
#853490000000
0#
0(
#853500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#853550000000
0$
0)
#853560000000
1"
1'
b0 +
b0 1
#853610000000
0"
0'
#853620000000
1#
1(
b101111101100100 +
b101111101100100 1
#853670000000
0#
0(
#853680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#853730000000
0$
0)
#853740000000
1"
1'
b0 +
b0 1
#853790000000
0"
0'
#853800000000
1#
1(
b101111101100100 +
b101111101100100 1
#853850000000
0#
0(
#853860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#853910000000
0$
0)
#853920000000
1"
1'
b0 +
b0 1
#853970000000
0"
0'
#853980000000
1#
1(
b101111101100100 +
b101111101100100 1
#854030000000
0#
0(
#854040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#854090000000
0$
0)
#854100000000
1"
1'
b0 +
b0 1
#854150000000
0"
0'
#854160000000
1#
1(
b101111101100100 +
b101111101100100 1
#854210000000
0#
0(
#854220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#854270000000
0$
0)
#854280000000
1"
1'
b0 +
b0 1
#854330000000
0"
0'
#854340000000
1#
1(
b101111101100100 +
b101111101100100 1
#854390000000
0#
0(
#854400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#854450000000
0$
0)
#854460000000
1"
1'
b0 +
b0 1
#854510000000
0"
0'
#854520000000
1#
1(
b101111101100100 +
b101111101100100 1
#854570000000
0#
0(
#854580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#854630000000
0$
0)
#854640000000
1"
1'
b0 +
b0 1
#854690000000
0"
0'
#854700000000
1#
1(
b101111101100100 +
b101111101100100 1
#854750000000
0#
0(
#854760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#854810000000
0$
0)
#854820000000
1"
1'
b0 +
b0 1
#854870000000
0"
0'
#854880000000
1#
1(
b101111101100100 +
b101111101100100 1
#854930000000
0#
0(
#854940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#854990000000
0$
0)
#855000000000
1"
1'
b0 +
b0 1
#855050000000
0"
0'
#855060000000
1#
1(
b101111101100100 +
b101111101100100 1
#855110000000
0#
0(
#855120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#855170000000
0$
0)
#855180000000
1"
1'
b0 +
b0 1
#855230000000
0"
0'
#855240000000
1#
1(
b101111101100100 +
b101111101100100 1
#855290000000
0#
0(
#855300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#855350000000
0$
0)
#855360000000
1"
1'
b0 +
b0 1
#855410000000
0"
0'
#855420000000
1#
1(
b101111101100100 +
b101111101100100 1
#855470000000
0#
0(
#855480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#855530000000
0$
0)
#855540000000
1"
1'
b0 +
b0 1
#855590000000
0"
0'
#855600000000
1#
1(
b101111101100100 +
b101111101100100 1
#855650000000
0#
0(
#855660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#855710000000
0$
0)
#855720000000
1"
1'
b0 +
b0 1
#855770000000
0"
0'
#855780000000
1#
1(
b101111101100100 +
b101111101100100 1
#855830000000
0#
0(
#855840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#855890000000
0$
0)
#855900000000
1"
1'
b0 +
b0 1
#855950000000
0"
0'
#855960000000
1#
1(
b101111101100100 +
b101111101100100 1
#856010000000
0#
0(
#856020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#856070000000
0$
0)
#856080000000
1"
1'
b0 +
b0 1
#856130000000
0"
0'
#856140000000
1#
1(
b101111101100100 +
b101111101100100 1
#856190000000
0#
0(
#856200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#856250000000
0$
0)
#856260000000
1"
1'
b0 +
b0 1
#856310000000
0"
0'
#856320000000
1#
1(
b101111101100100 +
b101111101100100 1
#856370000000
0#
0(
#856380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#856430000000
0$
0)
#856440000000
1"
1'
b0 +
b0 1
#856490000000
0"
0'
#856500000000
1#
1(
b101111101100100 +
b101111101100100 1
#856550000000
0#
0(
#856560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#856610000000
0$
0)
#856620000000
1"
1'
b0 +
b0 1
#856670000000
0"
0'
#856680000000
1#
1(
b101111101100100 +
b101111101100100 1
#856730000000
0#
0(
#856740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#856790000000
0$
0)
#856800000000
1"
1'
b0 +
b0 1
#856850000000
0"
0'
#856860000000
1#
1(
b101111101100100 +
b101111101100100 1
#856910000000
0#
0(
#856920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#856970000000
0$
0)
#856980000000
1"
1'
b0 +
b0 1
#857030000000
0"
0'
#857040000000
1#
1(
b101111101100100 +
b101111101100100 1
#857090000000
0#
0(
#857100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#857150000000
0$
0)
#857160000000
1"
1'
b0 +
b0 1
#857210000000
0"
0'
#857220000000
1#
1(
b101111101100100 +
b101111101100100 1
#857270000000
0#
0(
#857280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#857330000000
0$
0)
#857340000000
1"
1'
b0 +
b0 1
#857390000000
0"
0'
#857400000000
1#
1(
b101111101100100 +
b101111101100100 1
#857450000000
0#
0(
#857460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#857510000000
0$
0)
#857520000000
1"
1'
b0 +
b0 1
#857570000000
0"
0'
#857580000000
1#
1(
b101111101100100 +
b101111101100100 1
#857630000000
0#
0(
#857640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#857690000000
0$
0)
#857700000000
1"
1'
b0 +
b0 1
#857750000000
0"
0'
#857760000000
1#
1(
b101111101100100 +
b101111101100100 1
#857810000000
0#
0(
#857820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#857870000000
0$
0)
#857880000000
1"
1'
b0 +
b0 1
#857930000000
0"
0'
#857940000000
1#
1(
b101111101100100 +
b101111101100100 1
#857990000000
0#
0(
#858000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#858050000000
0$
0)
#858060000000
1"
1'
b0 +
b0 1
#858110000000
0"
0'
#858120000000
1#
1(
b101111101100100 +
b101111101100100 1
#858170000000
0#
0(
#858180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#858230000000
0$
0)
#858240000000
1"
1'
b0 +
b0 1
#858290000000
0"
0'
#858300000000
1#
1(
b101111101100100 +
b101111101100100 1
#858350000000
0#
0(
#858360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#858410000000
0$
0)
#858420000000
1"
1'
b0 +
b0 1
#858470000000
0"
0'
#858480000000
1#
1(
b101111101100100 +
b101111101100100 1
#858530000000
0#
0(
#858540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#858590000000
0$
0)
#858600000000
1"
1'
b0 +
b0 1
#858650000000
0"
0'
#858660000000
1#
1(
b101111101100100 +
b101111101100100 1
#858710000000
0#
0(
#858720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#858770000000
0$
0)
#858780000000
1"
1'
b0 +
b0 1
#858830000000
0"
0'
#858840000000
1#
1(
b101111101100100 +
b101111101100100 1
#858890000000
0#
0(
#858900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#858950000000
0$
0)
#858960000000
1"
1'
b0 +
b0 1
#859010000000
0"
0'
#859020000000
1#
1(
b101111101100100 +
b101111101100100 1
#859070000000
0#
0(
#859080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#859130000000
0$
0)
#859140000000
1"
1'
b0 +
b0 1
#859190000000
0"
0'
#859200000000
1#
1(
b101111101100100 +
b101111101100100 1
#859250000000
0#
0(
#859260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#859310000000
0$
0)
#859320000000
1"
1'
b0 +
b0 1
#859370000000
0"
0'
#859380000000
1#
1(
b101111101100100 +
b101111101100100 1
#859430000000
0#
0(
#859440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#859490000000
0$
0)
#859500000000
1"
1'
b0 +
b0 1
#859550000000
0"
0'
#859560000000
1#
1(
b101111101100100 +
b101111101100100 1
#859610000000
0#
0(
#859620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#859670000000
0$
0)
#859680000000
1"
1'
b0 +
b0 1
#859730000000
0"
0'
#859740000000
1#
1(
b101111101100100 +
b101111101100100 1
#859790000000
0#
0(
#859800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#859850000000
0$
0)
#859860000000
1"
1'
b0 +
b0 1
#859910000000
0"
0'
#859920000000
1#
1(
b101111101100100 +
b101111101100100 1
#859970000000
0#
0(
#859980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#860030000000
0$
0)
#860040000000
1"
1'
b0 +
b0 1
#860090000000
0"
0'
#860100000000
1#
1(
b101111101100100 +
b101111101100100 1
#860150000000
0#
0(
#860160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#860210000000
0$
0)
#860220000000
1"
1'
b0 +
b0 1
#860270000000
0"
0'
#860280000000
1#
1(
b101111101100100 +
b101111101100100 1
#860330000000
0#
0(
#860340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#860390000000
0$
0)
#860400000000
1"
1'
b0 +
b0 1
#860450000000
0"
0'
#860460000000
1#
1(
b101111101100100 +
b101111101100100 1
#860510000000
0#
0(
#860520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#860570000000
0$
0)
#860580000000
1"
1'
b0 +
b0 1
#860630000000
0"
0'
#860640000000
1#
1(
b101111101100100 +
b101111101100100 1
#860690000000
0#
0(
#860700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#860750000000
0$
0)
#860760000000
1"
1'
b0 +
b0 1
#860810000000
0"
0'
#860820000000
1#
1(
b101111101100100 +
b101111101100100 1
#860870000000
0#
0(
#860880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#860930000000
0$
0)
#860940000000
1"
1'
b0 +
b0 1
#860990000000
0"
0'
#861000000000
1#
1(
b101111101100100 +
b101111101100100 1
#861050000000
0#
0(
#861060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#861110000000
0$
0)
#861120000000
1"
1'
b0 +
b0 1
#861170000000
0"
0'
#861180000000
1#
1(
b101111101100100 +
b101111101100100 1
#861230000000
0#
0(
#861240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#861290000000
0$
0)
#861300000000
1"
1'
b0 +
b0 1
#861350000000
0"
0'
#861360000000
1#
1(
b101111101100100 +
b101111101100100 1
#861410000000
0#
0(
#861420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#861470000000
0$
0)
#861480000000
1"
1'
b0 +
b0 1
#861530000000
0"
0'
#861540000000
1#
1(
b101111101100100 +
b101111101100100 1
#861590000000
0#
0(
#861600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#861650000000
0$
0)
#861660000000
1"
1'
b0 +
b0 1
#861710000000
0"
0'
#861720000000
1#
1(
b101111101100100 +
b101111101100100 1
#861770000000
0#
0(
#861780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#861830000000
0$
0)
#861840000000
1"
1'
b0 +
b0 1
#861890000000
0"
0'
#861900000000
1#
1(
b101111101100100 +
b101111101100100 1
#861950000000
0#
0(
#861960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#862010000000
0$
0)
#862020000000
1"
1'
b0 +
b0 1
#862070000000
0"
0'
#862080000000
1#
1(
b101111101100100 +
b101111101100100 1
#862130000000
0#
0(
#862140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#862190000000
0$
0)
#862200000000
1"
1'
b0 +
b0 1
#862250000000
0"
0'
#862260000000
1#
1(
b101111101100100 +
b101111101100100 1
#862310000000
0#
0(
#862320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#862370000000
0$
0)
#862380000000
1"
1'
b0 +
b0 1
#862430000000
0"
0'
#862440000000
1#
1(
b101111101100100 +
b101111101100100 1
#862490000000
0#
0(
#862500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#862550000000
0$
0)
#862560000000
1"
1'
b0 +
b0 1
#862610000000
0"
0'
#862620000000
1#
1(
b101111101100100 +
b101111101100100 1
#862670000000
0#
0(
#862680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#862730000000
0$
0)
#862740000000
1"
1'
b0 +
b0 1
#862790000000
0"
0'
#862800000000
1#
1(
b101111101100100 +
b101111101100100 1
#862850000000
0#
0(
#862860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#862910000000
0$
0)
#862920000000
1"
1'
b0 +
b0 1
#862970000000
0"
0'
#862980000000
1#
1(
b101111101100100 +
b101111101100100 1
#863030000000
0#
0(
#863040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#863090000000
0$
0)
#863100000000
1"
1'
b0 +
b0 1
#863150000000
0"
0'
#863160000000
1#
1(
b101111101100100 +
b101111101100100 1
#863210000000
0#
0(
#863220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#863270000000
0$
0)
#863280000000
1"
1'
b0 +
b0 1
#863330000000
0"
0'
#863340000000
1#
1(
b101111101100100 +
b101111101100100 1
#863390000000
0#
0(
#863400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#863450000000
0$
0)
#863460000000
1"
1'
b0 +
b0 1
#863510000000
0"
0'
#863520000000
1#
1(
b101111101100100 +
b101111101100100 1
#863570000000
0#
0(
#863580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#863630000000
0$
0)
#863640000000
1"
1'
b0 +
b0 1
#863690000000
0"
0'
#863700000000
1#
1(
b101111101100100 +
b101111101100100 1
#863750000000
0#
0(
#863760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#863810000000
0$
0)
#863820000000
1"
1'
b0 +
b0 1
#863870000000
0"
0'
#863880000000
1#
1(
b101111101100100 +
b101111101100100 1
#863930000000
0#
0(
#863940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#863990000000
0$
0)
#864000000000
1"
1'
b0 +
b0 1
#864050000000
0"
0'
#864060000000
1#
1(
b101111101100100 +
b101111101100100 1
#864110000000
0#
0(
#864120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#864170000000
0$
0)
#864180000000
1"
1'
b0 +
b0 1
#864230000000
0"
0'
#864240000000
1#
1(
b101111101100100 +
b101111101100100 1
#864290000000
0#
0(
#864300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#864350000000
0$
0)
#864360000000
1"
1'
b0 +
b0 1
#864410000000
0"
0'
#864420000000
1#
1(
b101111101100100 +
b101111101100100 1
#864470000000
0#
0(
#864480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#864530000000
0$
0)
#864540000000
1"
1'
b0 +
b0 1
#864590000000
0"
0'
#864600000000
1#
1(
b101111101100100 +
b101111101100100 1
#864650000000
0#
0(
#864660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#864710000000
0$
0)
#864720000000
1"
1'
b0 +
b0 1
#864770000000
0"
0'
#864780000000
1#
1(
b101111101100100 +
b101111101100100 1
#864830000000
0#
0(
#864840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#864890000000
0$
0)
#864900000000
1"
1'
b0 +
b0 1
#864950000000
0"
0'
#864960000000
1#
1(
b101111101100100 +
b101111101100100 1
#865010000000
0#
0(
#865020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#865070000000
0$
0)
#865080000000
1"
1'
b0 +
b0 1
#865130000000
0"
0'
#865140000000
1#
1(
b101111101100100 +
b101111101100100 1
#865190000000
0#
0(
#865200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#865250000000
0$
0)
#865260000000
1"
1'
b0 +
b0 1
#865310000000
0"
0'
#865320000000
1#
1(
b101111101100100 +
b101111101100100 1
#865370000000
0#
0(
#865380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#865430000000
0$
0)
#865440000000
1"
1'
b0 +
b0 1
#865490000000
0"
0'
#865500000000
1#
1(
b101111101100100 +
b101111101100100 1
#865550000000
0#
0(
#865560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#865610000000
0$
0)
#865620000000
1"
1'
b0 +
b0 1
#865670000000
0"
0'
#865680000000
1#
1(
b101111101100100 +
b101111101100100 1
#865730000000
0#
0(
#865740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#865790000000
0$
0)
#865800000000
1"
1'
b0 +
b0 1
#865850000000
0"
0'
#865860000000
1#
1(
b101111101100100 +
b101111101100100 1
#865910000000
0#
0(
#865920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#865970000000
0$
0)
#865980000000
1"
1'
b0 +
b0 1
#866030000000
0"
0'
#866040000000
1#
1(
b101111101100100 +
b101111101100100 1
#866090000000
0#
0(
#866100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#866150000000
0$
0)
#866160000000
1"
1'
b0 +
b0 1
#866210000000
0"
0'
#866220000000
1#
1(
b101111101100100 +
b101111101100100 1
#866270000000
0#
0(
#866280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#866330000000
0$
0)
#866340000000
1"
1'
b0 +
b0 1
#866390000000
0"
0'
#866400000000
1#
1(
b101111101100100 +
b101111101100100 1
#866450000000
0#
0(
#866460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#866510000000
0$
0)
#866520000000
1"
1'
b0 +
b0 1
#866570000000
0"
0'
#866580000000
1#
1(
b101111101100100 +
b101111101100100 1
#866630000000
0#
0(
#866640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#866690000000
0$
0)
#866700000000
1"
1'
b0 +
b0 1
#866750000000
0"
0'
#866760000000
1#
1(
b101111101100100 +
b101111101100100 1
#866810000000
0#
0(
#866820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#866870000000
0$
0)
#866880000000
1"
1'
b0 +
b0 1
#866930000000
0"
0'
#866940000000
1#
1(
b101111101100100 +
b101111101100100 1
#866990000000
0#
0(
#867000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#867050000000
0$
0)
#867060000000
1"
1'
b0 +
b0 1
#867110000000
0"
0'
#867120000000
1#
1(
b101111101100100 +
b101111101100100 1
#867170000000
0#
0(
#867180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#867230000000
0$
0)
#867240000000
1"
1'
b0 +
b0 1
#867290000000
0"
0'
#867300000000
1#
1(
b101111101100100 +
b101111101100100 1
#867350000000
0#
0(
#867360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#867410000000
0$
0)
#867420000000
1"
1'
b0 +
b0 1
#867470000000
0"
0'
#867480000000
1#
1(
b101111101100100 +
b101111101100100 1
#867530000000
0#
0(
#867540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#867590000000
0$
0)
#867600000000
1"
1'
b0 +
b0 1
#867650000000
0"
0'
#867660000000
1#
1(
b101111101100100 +
b101111101100100 1
#867710000000
0#
0(
#867720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#867770000000
0$
0)
#867780000000
1"
1'
b0 +
b0 1
#867830000000
0"
0'
#867840000000
1#
1(
b101111101100100 +
b101111101100100 1
#867890000000
0#
0(
#867900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#867950000000
0$
0)
#867960000000
1"
1'
b0 +
b0 1
#868010000000
0"
0'
#868020000000
1#
1(
b101111101100100 +
b101111101100100 1
#868070000000
0#
0(
#868080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#868130000000
0$
0)
#868140000000
1"
1'
b0 +
b0 1
#868190000000
0"
0'
#868200000000
1#
1(
b101111101100100 +
b101111101100100 1
#868250000000
0#
0(
#868260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#868310000000
0$
0)
#868320000000
1"
1'
b0 +
b0 1
#868370000000
0"
0'
#868380000000
1#
1(
b101111101100100 +
b101111101100100 1
#868430000000
0#
0(
#868440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#868490000000
0$
0)
#868500000000
1"
1'
b0 +
b0 1
#868550000000
0"
0'
#868560000000
1#
1(
b101111101100100 +
b101111101100100 1
#868610000000
0#
0(
#868620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#868670000000
0$
0)
#868680000000
1"
1'
b0 +
b0 1
#868730000000
0"
0'
#868740000000
1#
1(
b101111101100100 +
b101111101100100 1
#868790000000
0#
0(
#868800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#868850000000
0$
0)
#868860000000
1"
1'
b0 +
b0 1
#868910000000
0"
0'
#868920000000
1#
1(
b101111101100100 +
b101111101100100 1
#868970000000
0#
0(
#868980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#869030000000
0$
0)
#869040000000
1"
1'
b0 +
b0 1
#869090000000
0"
0'
#869100000000
1#
1(
b101111101100100 +
b101111101100100 1
#869150000000
0#
0(
#869160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#869210000000
0$
0)
#869220000000
1"
1'
b0 +
b0 1
#869270000000
0"
0'
#869280000000
1#
1(
b101111101100100 +
b101111101100100 1
#869330000000
0#
0(
#869340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#869390000000
0$
0)
#869400000000
1"
1'
b0 +
b0 1
#869450000000
0"
0'
#869460000000
1#
1(
b101111101100100 +
b101111101100100 1
#869510000000
0#
0(
#869520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#869570000000
0$
0)
#869580000000
1"
1'
b0 +
b0 1
#869630000000
0"
0'
#869640000000
1#
1(
b101111101100100 +
b101111101100100 1
#869690000000
0#
0(
#869700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#869750000000
0$
0)
#869760000000
1"
1'
b0 +
b0 1
#869810000000
0"
0'
#869820000000
1#
1(
b101111101100100 +
b101111101100100 1
#869870000000
0#
0(
#869880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#869930000000
0$
0)
#869940000000
1"
1'
b0 +
b0 1
#869990000000
0"
0'
#870000000000
1#
1(
b101111101100100 +
b101111101100100 1
#870050000000
0#
0(
#870060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#870110000000
0$
0)
#870120000000
1"
1'
b0 +
b0 1
#870170000000
0"
0'
#870180000000
1#
1(
b101111101100100 +
b101111101100100 1
#870230000000
0#
0(
#870240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#870290000000
0$
0)
#870300000000
1"
1'
b0 +
b0 1
#870350000000
0"
0'
#870360000000
1#
1(
b101111101100100 +
b101111101100100 1
#870410000000
0#
0(
#870420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#870470000000
0$
0)
#870480000000
1"
1'
b0 +
b0 1
#870530000000
0"
0'
#870540000000
1#
1(
b101111101100100 +
b101111101100100 1
#870590000000
0#
0(
#870600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#870650000000
0$
0)
#870660000000
1"
1'
b0 +
b0 1
#870710000000
0"
0'
#870720000000
1#
1(
b101111101100100 +
b101111101100100 1
#870770000000
0#
0(
#870780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#870830000000
0$
0)
#870840000000
1"
1'
b0 +
b0 1
#870890000000
0"
0'
#870900000000
1#
1(
b101111101100100 +
b101111101100100 1
#870950000000
0#
0(
#870960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#871010000000
0$
0)
#871020000000
1"
1'
b0 +
b0 1
#871070000000
0"
0'
#871080000000
1#
1(
b101111101100100 +
b101111101100100 1
#871130000000
0#
0(
#871140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#871190000000
0$
0)
#871200000000
1"
1'
b0 +
b0 1
#871250000000
0"
0'
#871260000000
1#
1(
b101111101100100 +
b101111101100100 1
#871310000000
0#
0(
#871320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#871370000000
0$
0)
#871380000000
1"
1'
b0 +
b0 1
#871430000000
0"
0'
#871440000000
1#
1(
b101111101100100 +
b101111101100100 1
#871490000000
0#
0(
#871500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#871550000000
0$
0)
#871560000000
1"
1'
b0 +
b0 1
#871610000000
0"
0'
#871620000000
1#
1(
b101111101100100 +
b101111101100100 1
#871670000000
0#
0(
#871680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#871730000000
0$
0)
#871740000000
1"
1'
b0 +
b0 1
#871790000000
0"
0'
#871800000000
1#
1(
b101111101100100 +
b101111101100100 1
#871850000000
0#
0(
#871860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#871910000000
0$
0)
#871920000000
1"
1'
b0 +
b0 1
#871970000000
0"
0'
#871980000000
1#
1(
b101111101100100 +
b101111101100100 1
#872030000000
0#
0(
#872040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#872090000000
0$
0)
#872100000000
1"
1'
b0 +
b0 1
#872150000000
0"
0'
#872160000000
1#
1(
b101111101100100 +
b101111101100100 1
#872210000000
0#
0(
#872220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#872270000000
0$
0)
#872280000000
1"
1'
b0 +
b0 1
#872330000000
0"
0'
#872340000000
1#
1(
b101111101100100 +
b101111101100100 1
#872390000000
0#
0(
#872400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#872450000000
0$
0)
#872460000000
1"
1'
b0 +
b0 1
#872510000000
0"
0'
#872520000000
1#
1(
b101111101100100 +
b101111101100100 1
#872570000000
0#
0(
#872580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#872630000000
0$
0)
#872640000000
1"
1'
b0 +
b0 1
#872690000000
0"
0'
#872700000000
1#
1(
b101111101100100 +
b101111101100100 1
#872750000000
0#
0(
#872760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#872810000000
0$
0)
#872820000000
1"
1'
b0 +
b0 1
#872870000000
0"
0'
#872880000000
1#
1(
b101111101100100 +
b101111101100100 1
#872930000000
0#
0(
#872940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#872990000000
0$
0)
#873000000000
1"
1'
b0 +
b0 1
#873050000000
0"
0'
#873060000000
1#
1(
b101111101100100 +
b101111101100100 1
#873110000000
0#
0(
#873120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#873170000000
0$
0)
#873180000000
1"
1'
b0 +
b0 1
#873230000000
0"
0'
#873240000000
1#
1(
b101111101100100 +
b101111101100100 1
#873290000000
0#
0(
#873300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#873350000000
0$
0)
#873360000000
1"
1'
b0 +
b0 1
#873410000000
0"
0'
#873420000000
1#
1(
b101111101100100 +
b101111101100100 1
#873470000000
0#
0(
#873480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#873530000000
0$
0)
#873540000000
1"
1'
b0 +
b0 1
#873590000000
0"
0'
#873600000000
1#
1(
b101111101100100 +
b101111101100100 1
#873650000000
0#
0(
#873660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#873710000000
0$
0)
#873720000000
1"
1'
b0 +
b0 1
#873770000000
0"
0'
#873780000000
1#
1(
b101111101100100 +
b101111101100100 1
#873830000000
0#
0(
#873840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#873890000000
0$
0)
#873900000000
1"
1'
b0 +
b0 1
#873950000000
0"
0'
#873960000000
1#
1(
b101111101100100 +
b101111101100100 1
#874010000000
0#
0(
#874020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#874070000000
0$
0)
#874080000000
1"
1'
b0 +
b0 1
#874130000000
0"
0'
#874140000000
1#
1(
b101111101100100 +
b101111101100100 1
#874190000000
0#
0(
#874200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#874250000000
0$
0)
#874260000000
1"
1'
b0 +
b0 1
#874310000000
0"
0'
#874320000000
1#
1(
b101111101100100 +
b101111101100100 1
#874370000000
0#
0(
#874380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#874430000000
0$
0)
#874440000000
1"
1'
b0 +
b0 1
#874490000000
0"
0'
#874500000000
1#
1(
b101111101100100 +
b101111101100100 1
#874550000000
0#
0(
#874560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#874610000000
0$
0)
#874620000000
1"
1'
b0 +
b0 1
#874670000000
0"
0'
#874680000000
1#
1(
b101111101100100 +
b101111101100100 1
#874730000000
0#
0(
#874740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#874790000000
0$
0)
#874800000000
1"
1'
b0 +
b0 1
#874850000000
0"
0'
#874860000000
1#
1(
b101111101100100 +
b101111101100100 1
#874910000000
0#
0(
#874920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#874970000000
0$
0)
#874980000000
1"
1'
b0 +
b0 1
#875030000000
0"
0'
#875040000000
1#
1(
b101111101100100 +
b101111101100100 1
#875090000000
0#
0(
#875100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#875150000000
0$
0)
#875160000000
1"
1'
b0 +
b0 1
#875210000000
0"
0'
#875220000000
1#
1(
b101111101100100 +
b101111101100100 1
#875270000000
0#
0(
#875280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#875330000000
0$
0)
#875340000000
1"
1'
b0 +
b0 1
#875390000000
0"
0'
#875400000000
1#
1(
b101111101100100 +
b101111101100100 1
#875450000000
0#
0(
#875460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#875510000000
0$
0)
#875520000000
1"
1'
b0 +
b0 1
#875570000000
0"
0'
#875580000000
1#
1(
b101111101100100 +
b101111101100100 1
#875630000000
0#
0(
#875640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#875690000000
0$
0)
#875700000000
1"
1'
b0 +
b0 1
#875750000000
0"
0'
#875760000000
1#
1(
b101111101100100 +
b101111101100100 1
#875810000000
0#
0(
#875820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#875870000000
0$
0)
#875880000000
1"
1'
b0 +
b0 1
#875930000000
0"
0'
#875940000000
1#
1(
b101111101100100 +
b101111101100100 1
#875990000000
0#
0(
#876000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#876050000000
0$
0)
#876060000000
1"
1'
b0 +
b0 1
#876110000000
0"
0'
#876120000000
1#
1(
b101111101100100 +
b101111101100100 1
#876170000000
0#
0(
#876180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#876230000000
0$
0)
#876240000000
1"
1'
b0 +
b0 1
#876290000000
0"
0'
#876300000000
1#
1(
b101111101100100 +
b101111101100100 1
#876350000000
0#
0(
#876360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#876410000000
0$
0)
#876420000000
1"
1'
b0 +
b0 1
#876470000000
0"
0'
#876480000000
1#
1(
b101111101100100 +
b101111101100100 1
#876530000000
0#
0(
#876540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#876590000000
0$
0)
#876600000000
1"
1'
b0 +
b0 1
#876650000000
0"
0'
#876660000000
1#
1(
b101111101100100 +
b101111101100100 1
#876710000000
0#
0(
#876720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#876770000000
0$
0)
#876780000000
1"
1'
b0 +
b0 1
#876830000000
0"
0'
#876840000000
1#
1(
b101111101100100 +
b101111101100100 1
#876890000000
0#
0(
#876900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#876950000000
0$
0)
#876960000000
1"
1'
b0 +
b0 1
#877010000000
0"
0'
#877020000000
1#
1(
b101111101100100 +
b101111101100100 1
#877070000000
0#
0(
#877080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#877130000000
0$
0)
#877140000000
1"
1'
b0 +
b0 1
#877190000000
0"
0'
#877200000000
1#
1(
b101111101100100 +
b101111101100100 1
#877250000000
0#
0(
#877260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#877310000000
0$
0)
#877320000000
1"
1'
b0 +
b0 1
#877370000000
0"
0'
#877380000000
1#
1(
b101111101100100 +
b101111101100100 1
#877430000000
0#
0(
#877440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#877490000000
0$
0)
#877500000000
1"
1'
b0 +
b0 1
#877550000000
0"
0'
#877560000000
1#
1(
b101111101100100 +
b101111101100100 1
#877610000000
0#
0(
#877620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#877670000000
0$
0)
#877680000000
1"
1'
b0 +
b0 1
#877730000000
0"
0'
#877740000000
1#
1(
b101111101100100 +
b101111101100100 1
#877790000000
0#
0(
#877800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#877850000000
0$
0)
#877860000000
1"
1'
b0 +
b0 1
#877910000000
0"
0'
#877920000000
1#
1(
b101111101100100 +
b101111101100100 1
#877970000000
0#
0(
#877980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#878030000000
0$
0)
#878040000000
1"
1'
b0 +
b0 1
#878090000000
0"
0'
#878100000000
1#
1(
b101111101100100 +
b101111101100100 1
#878150000000
0#
0(
#878160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#878210000000
0$
0)
#878220000000
1"
1'
b0 +
b0 1
#878270000000
0"
0'
#878280000000
1#
1(
b101111101100100 +
b101111101100100 1
#878330000000
0#
0(
#878340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#878390000000
0$
0)
#878400000000
1"
1'
b0 +
b0 1
#878450000000
0"
0'
#878460000000
1#
1(
b101111101100100 +
b101111101100100 1
#878510000000
0#
0(
#878520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#878570000000
0$
0)
#878580000000
1"
1'
b0 +
b0 1
#878630000000
0"
0'
#878640000000
1#
1(
b101111101100100 +
b101111101100100 1
#878690000000
0#
0(
#878700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#878750000000
0$
0)
#878760000000
1"
1'
b0 +
b0 1
#878810000000
0"
0'
#878820000000
1#
1(
b101111101100100 +
b101111101100100 1
#878870000000
0#
0(
#878880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#878930000000
0$
0)
#878940000000
1"
1'
b0 +
b0 1
#878990000000
0"
0'
#879000000000
1#
1(
b101111101100100 +
b101111101100100 1
#879050000000
0#
0(
#879060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#879110000000
0$
0)
#879120000000
1"
1'
b0 +
b0 1
#879170000000
0"
0'
#879180000000
1#
1(
b101111101100100 +
b101111101100100 1
#879230000000
0#
0(
#879240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#879290000000
0$
0)
#879300000000
1"
1'
b0 +
b0 1
#879350000000
0"
0'
#879360000000
1#
1(
b101111101100100 +
b101111101100100 1
#879410000000
0#
0(
#879420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#879470000000
0$
0)
#879480000000
1"
1'
b0 +
b0 1
#879530000000
0"
0'
#879540000000
1#
1(
b101111101100100 +
b101111101100100 1
#879590000000
0#
0(
#879600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#879650000000
0$
0)
#879660000000
1"
1'
b0 +
b0 1
#879710000000
0"
0'
#879720000000
1#
1(
b101111101100100 +
b101111101100100 1
#879770000000
0#
0(
#879780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#879830000000
0$
0)
#879840000000
1"
1'
b0 +
b0 1
#879890000000
0"
0'
#879900000000
1#
1(
b101111101100100 +
b101111101100100 1
#879950000000
0#
0(
#879960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#880010000000
0$
0)
#880020000000
1"
1'
b0 +
b0 1
#880070000000
0"
0'
#880080000000
1#
1(
b101111101100100 +
b101111101100100 1
#880130000000
0#
0(
#880140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#880190000000
0$
0)
#880200000000
1"
1'
b0 +
b0 1
#880250000000
0"
0'
#880260000000
1#
1(
b101111101100100 +
b101111101100100 1
#880310000000
0#
0(
#880320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#880370000000
0$
0)
#880380000000
1"
1'
b0 +
b0 1
#880430000000
0"
0'
#880440000000
1#
1(
b101111101100100 +
b101111101100100 1
#880490000000
0#
0(
#880500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#880550000000
0$
0)
#880560000000
1"
1'
b0 +
b0 1
#880610000000
0"
0'
#880620000000
1#
1(
b101111101100100 +
b101111101100100 1
#880670000000
0#
0(
#880680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#880730000000
0$
0)
#880740000000
1"
1'
b0 +
b0 1
#880790000000
0"
0'
#880800000000
1#
1(
b101111101100100 +
b101111101100100 1
#880850000000
0#
0(
#880860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#880910000000
0$
0)
#880920000000
1"
1'
b0 +
b0 1
#880970000000
0"
0'
#880980000000
1#
1(
b101111101100100 +
b101111101100100 1
#881030000000
0#
0(
#881040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#881090000000
0$
0)
#881100000000
1"
1'
b0 +
b0 1
#881150000000
0"
0'
#881160000000
1#
1(
b101111101100100 +
b101111101100100 1
#881210000000
0#
0(
#881220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#881270000000
0$
0)
#881280000000
1"
1'
b0 +
b0 1
#881330000000
0"
0'
#881340000000
1#
1(
b101111101100100 +
b101111101100100 1
#881390000000
0#
0(
#881400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#881450000000
0$
0)
#881460000000
1"
1'
b0 +
b0 1
#881510000000
0"
0'
#881520000000
1#
1(
b101111101100100 +
b101111101100100 1
#881570000000
0#
0(
#881580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#881630000000
0$
0)
#881640000000
1"
1'
b0 +
b0 1
#881690000000
0"
0'
#881700000000
1#
1(
b101111101100100 +
b101111101100100 1
#881750000000
0#
0(
#881760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#881810000000
0$
0)
#881820000000
1"
1'
b0 +
b0 1
#881870000000
0"
0'
#881880000000
1#
1(
b101111101100100 +
b101111101100100 1
#881930000000
0#
0(
#881940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#881990000000
0$
0)
#882000000000
1"
1'
b0 +
b0 1
#882050000000
0"
0'
#882060000000
1#
1(
b101111101100100 +
b101111101100100 1
#882110000000
0#
0(
#882120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#882170000000
0$
0)
#882180000000
1"
1'
b0 +
b0 1
#882230000000
0"
0'
#882240000000
1#
1(
b101111101100100 +
b101111101100100 1
#882290000000
0#
0(
#882300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#882350000000
0$
0)
#882360000000
1"
1'
b0 +
b0 1
#882410000000
0"
0'
#882420000000
1#
1(
b101111101100100 +
b101111101100100 1
#882470000000
0#
0(
#882480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#882530000000
0$
0)
#882540000000
1"
1'
b0 +
b0 1
#882590000000
0"
0'
#882600000000
1#
1(
b101111101100100 +
b101111101100100 1
#882650000000
0#
0(
#882660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#882710000000
0$
0)
#882720000000
1"
1'
b0 +
b0 1
#882770000000
0"
0'
#882780000000
1#
1(
b101111101100100 +
b101111101100100 1
#882830000000
0#
0(
#882840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#882890000000
0$
0)
#882900000000
1"
1'
b0 +
b0 1
#882950000000
0"
0'
#882960000000
1#
1(
b101111101100100 +
b101111101100100 1
#883010000000
0#
0(
#883020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#883070000000
0$
0)
#883080000000
1"
1'
b0 +
b0 1
#883130000000
0"
0'
#883140000000
1#
1(
b101111101100100 +
b101111101100100 1
#883190000000
0#
0(
#883200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#883250000000
0$
0)
#883260000000
1"
1'
b0 +
b0 1
#883310000000
0"
0'
#883320000000
1#
1(
b101111101100100 +
b101111101100100 1
#883370000000
0#
0(
#883380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#883430000000
0$
0)
#883440000000
1"
1'
b0 +
b0 1
#883490000000
0"
0'
#883500000000
1#
1(
b101111101100100 +
b101111101100100 1
#883550000000
0#
0(
#883560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#883610000000
0$
0)
#883620000000
1"
1'
b0 +
b0 1
#883670000000
0"
0'
#883680000000
1#
1(
b101111101100100 +
b101111101100100 1
#883730000000
0#
0(
#883740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#883790000000
0$
0)
#883800000000
1"
1'
b0 +
b0 1
#883850000000
0"
0'
#883860000000
1#
1(
b101111101100100 +
b101111101100100 1
#883910000000
0#
0(
#883920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#883970000000
0$
0)
#883980000000
1"
1'
b0 +
b0 1
#884030000000
0"
0'
#884040000000
1#
1(
b101111101100100 +
b101111101100100 1
#884090000000
0#
0(
#884100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#884150000000
0$
0)
#884160000000
1"
1'
b0 +
b0 1
#884210000000
0"
0'
#884220000000
1#
1(
b101111101100100 +
b101111101100100 1
#884270000000
0#
0(
#884280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#884330000000
0$
0)
#884340000000
1"
1'
b0 +
b0 1
#884390000000
0"
0'
#884400000000
1#
1(
b101111101100100 +
b101111101100100 1
#884450000000
0#
0(
#884460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#884510000000
0$
0)
#884520000000
1"
1'
b0 +
b0 1
#884570000000
0"
0'
#884580000000
1#
1(
b101111101100100 +
b101111101100100 1
#884630000000
0#
0(
#884640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#884690000000
0$
0)
#884700000000
1"
1'
b0 +
b0 1
#884750000000
0"
0'
#884760000000
1#
1(
b101111101100100 +
b101111101100100 1
#884810000000
0#
0(
#884820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#884870000000
0$
0)
#884880000000
1"
1'
b0 +
b0 1
#884930000000
0"
0'
#884940000000
1#
1(
b101111101100100 +
b101111101100100 1
#884990000000
0#
0(
#885000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#885050000000
0$
0)
#885060000000
1"
1'
b0 +
b0 1
#885110000000
0"
0'
#885120000000
1#
1(
b101111101100100 +
b101111101100100 1
#885170000000
0#
0(
#885180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#885230000000
0$
0)
#885240000000
1"
1'
b0 +
b0 1
#885290000000
0"
0'
#885300000000
1#
1(
b101111101100100 +
b101111101100100 1
#885350000000
0#
0(
#885360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#885410000000
0$
0)
#885420000000
1"
1'
b0 +
b0 1
#885470000000
0"
0'
#885480000000
1#
1(
b101111101100100 +
b101111101100100 1
#885530000000
0#
0(
#885540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#885590000000
0$
0)
#885600000000
1"
1'
b0 +
b0 1
#885650000000
0"
0'
#885660000000
1#
1(
b101111101100100 +
b101111101100100 1
#885710000000
0#
0(
#885720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#885770000000
0$
0)
#885780000000
1"
1'
b0 +
b0 1
#885830000000
0"
0'
#885840000000
1#
1(
b101111101100100 +
b101111101100100 1
#885890000000
0#
0(
#885900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#885950000000
0$
0)
#885960000000
1"
1'
b0 +
b0 1
#886010000000
0"
0'
#886020000000
1#
1(
b101111101100100 +
b101111101100100 1
#886070000000
0#
0(
#886080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#886130000000
0$
0)
#886140000000
1"
1'
b0 +
b0 1
#886190000000
0"
0'
#886200000000
1#
1(
b101111101100100 +
b101111101100100 1
#886250000000
0#
0(
#886260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#886310000000
0$
0)
#886320000000
1"
1'
b0 +
b0 1
#886370000000
0"
0'
#886380000000
1#
1(
b101111101100100 +
b101111101100100 1
#886430000000
0#
0(
#886440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#886490000000
0$
0)
#886500000000
1"
1'
b0 +
b0 1
#886550000000
0"
0'
#886560000000
1#
1(
b101111101100100 +
b101111101100100 1
#886610000000
0#
0(
#886620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#886670000000
0$
0)
#886680000000
1"
1'
b0 +
b0 1
#886730000000
0"
0'
#886740000000
1#
1(
b101111101100100 +
b101111101100100 1
#886790000000
0#
0(
#886800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#886850000000
0$
0)
#886860000000
1"
1'
b0 +
b0 1
#886910000000
0"
0'
#886920000000
1#
1(
b101111101100100 +
b101111101100100 1
#886970000000
0#
0(
#886980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#887030000000
0$
0)
#887040000000
1"
1'
b0 +
b0 1
#887090000000
0"
0'
#887100000000
1#
1(
b101111101100100 +
b101111101100100 1
#887150000000
0#
0(
#887160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#887210000000
0$
0)
#887220000000
1"
1'
b0 +
b0 1
#887270000000
0"
0'
#887280000000
1#
1(
b101111101100100 +
b101111101100100 1
#887330000000
0#
0(
#887340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#887390000000
0$
0)
#887400000000
1"
1'
b0 +
b0 1
#887450000000
0"
0'
#887460000000
1#
1(
b101111101100100 +
b101111101100100 1
#887510000000
0#
0(
#887520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#887570000000
0$
0)
#887580000000
1"
1'
b0 +
b0 1
#887630000000
0"
0'
#887640000000
1#
1(
b101111101100100 +
b101111101100100 1
#887690000000
0#
0(
#887700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#887750000000
0$
0)
#887760000000
1"
1'
b0 +
b0 1
#887810000000
0"
0'
#887820000000
1#
1(
b101111101100100 +
b101111101100100 1
#887870000000
0#
0(
#887880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#887930000000
0$
0)
#887940000000
1"
1'
b0 +
b0 1
#887990000000
0"
0'
#888000000000
1#
1(
b101111101100100 +
b101111101100100 1
#888050000000
0#
0(
#888060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#888110000000
0$
0)
#888120000000
1"
1'
b0 +
b0 1
#888170000000
0"
0'
#888180000000
1#
1(
b101111101100100 +
b101111101100100 1
#888230000000
0#
0(
#888240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#888290000000
0$
0)
#888300000000
1"
1'
b0 +
b0 1
#888350000000
0"
0'
#888360000000
1#
1(
b101111101100100 +
b101111101100100 1
#888410000000
0#
0(
#888420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#888470000000
0$
0)
#888480000000
1"
1'
b0 +
b0 1
#888530000000
0"
0'
#888540000000
1#
1(
b101111101100100 +
b101111101100100 1
#888590000000
0#
0(
#888600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#888650000000
0$
0)
#888660000000
1"
1'
b0 +
b0 1
#888710000000
0"
0'
#888720000000
1#
1(
b101111101100100 +
b101111101100100 1
#888770000000
0#
0(
#888780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#888830000000
0$
0)
#888840000000
1"
1'
b0 +
b0 1
#888890000000
0"
0'
#888900000000
1#
1(
b101111101100100 +
b101111101100100 1
#888950000000
0#
0(
#888960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#889010000000
0$
0)
#889020000000
1"
1'
b0 +
b0 1
#889070000000
0"
0'
#889080000000
1#
1(
b101111101100100 +
b101111101100100 1
#889130000000
0#
0(
#889140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#889190000000
0$
0)
#889200000000
1"
1'
b0 +
b0 1
#889250000000
0"
0'
#889260000000
1#
1(
b101111101100100 +
b101111101100100 1
#889310000000
0#
0(
#889320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#889370000000
0$
0)
#889380000000
1"
1'
b0 +
b0 1
#889430000000
0"
0'
#889440000000
1#
1(
b101111101100100 +
b101111101100100 1
#889490000000
0#
0(
#889500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#889550000000
0$
0)
#889560000000
1"
1'
b0 +
b0 1
#889610000000
0"
0'
#889620000000
1#
1(
b101111101100100 +
b101111101100100 1
#889670000000
0#
0(
#889680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#889730000000
0$
0)
#889740000000
1"
1'
b0 +
b0 1
#889790000000
0"
0'
#889800000000
1#
1(
b101111101100100 +
b101111101100100 1
#889850000000
0#
0(
#889860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#889910000000
0$
0)
#889920000000
1"
1'
b0 +
b0 1
#889970000000
0"
0'
#889980000000
1#
1(
b101111101100100 +
b101111101100100 1
#890030000000
0#
0(
#890040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#890090000000
0$
0)
#890100000000
1"
1'
b0 +
b0 1
#890150000000
0"
0'
#890160000000
1#
1(
b101111101100100 +
b101111101100100 1
#890210000000
0#
0(
#890220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#890270000000
0$
0)
#890280000000
1"
1'
b0 +
b0 1
#890330000000
0"
0'
#890340000000
1#
1(
b101111101100100 +
b101111101100100 1
#890390000000
0#
0(
#890400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#890450000000
0$
0)
#890460000000
1"
1'
b0 +
b0 1
#890510000000
0"
0'
#890520000000
1#
1(
b101111101100100 +
b101111101100100 1
#890570000000
0#
0(
#890580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#890630000000
0$
0)
#890640000000
1"
1'
b0 +
b0 1
#890690000000
0"
0'
#890700000000
1#
1(
b101111101100100 +
b101111101100100 1
#890750000000
0#
0(
#890760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#890810000000
0$
0)
#890820000000
1"
1'
b0 +
b0 1
#890870000000
0"
0'
#890880000000
1#
1(
b101111101100100 +
b101111101100100 1
#890930000000
0#
0(
#890940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#890990000000
0$
0)
#891000000000
1"
1'
b0 +
b0 1
#891050000000
0"
0'
#891060000000
1#
1(
b101111101100100 +
b101111101100100 1
#891110000000
0#
0(
#891120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#891170000000
0$
0)
#891180000000
1"
1'
b0 +
b0 1
#891230000000
0"
0'
#891240000000
1#
1(
b101111101100100 +
b101111101100100 1
#891290000000
0#
0(
#891300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#891350000000
0$
0)
#891360000000
1"
1'
b0 +
b0 1
#891410000000
0"
0'
#891420000000
1#
1(
b101111101100100 +
b101111101100100 1
#891470000000
0#
0(
#891480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#891530000000
0$
0)
#891540000000
1"
1'
b0 +
b0 1
#891590000000
0"
0'
#891600000000
1#
1(
b101111101100100 +
b101111101100100 1
#891650000000
0#
0(
#891660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#891710000000
0$
0)
#891720000000
1"
1'
b0 +
b0 1
#891770000000
0"
0'
#891780000000
1#
1(
b101111101100100 +
b101111101100100 1
#891830000000
0#
0(
#891840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#891890000000
0$
0)
#891900000000
1"
1'
b0 +
b0 1
#891950000000
0"
0'
#891960000000
1#
1(
b101111101100100 +
b101111101100100 1
#892010000000
0#
0(
#892020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#892070000000
0$
0)
#892080000000
1"
1'
b0 +
b0 1
#892130000000
0"
0'
#892140000000
1#
1(
b101111101100100 +
b101111101100100 1
#892190000000
0#
0(
#892200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#892250000000
0$
0)
#892260000000
1"
1'
b0 +
b0 1
#892310000000
0"
0'
#892320000000
1#
1(
b101111101100100 +
b101111101100100 1
#892370000000
0#
0(
#892380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#892430000000
0$
0)
#892440000000
1"
1'
b0 +
b0 1
#892490000000
0"
0'
#892500000000
1#
1(
b101111101100100 +
b101111101100100 1
#892550000000
0#
0(
#892560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#892610000000
0$
0)
#892620000000
1"
1'
b0 +
b0 1
#892670000000
0"
0'
#892680000000
1#
1(
b101111101100100 +
b101111101100100 1
#892730000000
0#
0(
#892740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#892790000000
0$
0)
#892800000000
1"
1'
b0 +
b0 1
#892850000000
0"
0'
#892860000000
1#
1(
b101111101100100 +
b101111101100100 1
#892910000000
0#
0(
#892920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#892970000000
0$
0)
#892980000000
1"
1'
b0 +
b0 1
#893030000000
0"
0'
#893040000000
1#
1(
b101111101100100 +
b101111101100100 1
#893090000000
0#
0(
#893100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#893150000000
0$
0)
#893160000000
1"
1'
b0 +
b0 1
#893210000000
0"
0'
#893220000000
1#
1(
b101111101100100 +
b101111101100100 1
#893270000000
0#
0(
#893280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#893330000000
0$
0)
#893340000000
1"
1'
b0 +
b0 1
#893390000000
0"
0'
#893400000000
1#
1(
b101111101100100 +
b101111101100100 1
#893450000000
0#
0(
#893460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#893510000000
0$
0)
#893520000000
1"
1'
b0 +
b0 1
#893570000000
0"
0'
#893580000000
1#
1(
b101111101100100 +
b101111101100100 1
#893630000000
0#
0(
#893640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#893690000000
0$
0)
#893700000000
1"
1'
b0 +
b0 1
#893750000000
0"
0'
#893760000000
1#
1(
b101111101100100 +
b101111101100100 1
#893810000000
0#
0(
#893820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#893870000000
0$
0)
#893880000000
1"
1'
b0 +
b0 1
#893930000000
0"
0'
#893940000000
1#
1(
b101111101100100 +
b101111101100100 1
#893990000000
0#
0(
#894000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#894050000000
0$
0)
#894060000000
1"
1'
b0 +
b0 1
#894110000000
0"
0'
#894120000000
1#
1(
b101111101100100 +
b101111101100100 1
#894170000000
0#
0(
#894180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#894230000000
0$
0)
#894240000000
1"
1'
b0 +
b0 1
#894290000000
0"
0'
#894300000000
1#
1(
b101111101100100 +
b101111101100100 1
#894350000000
0#
0(
#894360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#894410000000
0$
0)
#894420000000
1"
1'
b0 +
b0 1
#894470000000
0"
0'
#894480000000
1#
1(
b101111101100100 +
b101111101100100 1
#894530000000
0#
0(
#894540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#894590000000
0$
0)
#894600000000
1"
1'
b0 +
b0 1
#894650000000
0"
0'
#894660000000
1#
1(
b101111101100100 +
b101111101100100 1
#894710000000
0#
0(
#894720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#894770000000
0$
0)
#894780000000
1"
1'
b0 +
b0 1
#894830000000
0"
0'
#894840000000
1#
1(
b101111101100100 +
b101111101100100 1
#894890000000
0#
0(
#894900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#894950000000
0$
0)
#894960000000
1"
1'
b0 +
b0 1
#895010000000
0"
0'
#895020000000
1#
1(
b101111101100100 +
b101111101100100 1
#895070000000
0#
0(
#895080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#895130000000
0$
0)
#895140000000
1"
1'
b0 +
b0 1
#895190000000
0"
0'
#895200000000
1#
1(
b101111101100100 +
b101111101100100 1
#895250000000
0#
0(
#895260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#895310000000
0$
0)
#895320000000
1"
1'
b0 +
b0 1
#895370000000
0"
0'
#895380000000
1#
1(
b101111101100100 +
b101111101100100 1
#895430000000
0#
0(
#895440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#895490000000
0$
0)
#895500000000
1"
1'
b0 +
b0 1
#895550000000
0"
0'
#895560000000
1#
1(
b101111101100100 +
b101111101100100 1
#895610000000
0#
0(
#895620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#895670000000
0$
0)
#895680000000
1"
1'
b0 +
b0 1
#895730000000
0"
0'
#895740000000
1#
1(
b101111101100100 +
b101111101100100 1
#895790000000
0#
0(
#895800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#895850000000
0$
0)
#895860000000
1"
1'
b0 +
b0 1
#895910000000
0"
0'
#895920000000
1#
1(
b101111101100100 +
b101111101100100 1
#895970000000
0#
0(
#895980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#896030000000
0$
0)
#896040000000
1"
1'
b0 +
b0 1
#896090000000
0"
0'
#896100000000
1#
1(
b101111101100100 +
b101111101100100 1
#896150000000
0#
0(
#896160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#896210000000
0$
0)
#896220000000
1"
1'
b0 +
b0 1
#896270000000
0"
0'
#896280000000
1#
1(
b101111101100100 +
b101111101100100 1
#896330000000
0#
0(
#896340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#896390000000
0$
0)
#896400000000
1"
1'
b0 +
b0 1
#896450000000
0"
0'
#896460000000
1#
1(
b101111101100100 +
b101111101100100 1
#896510000000
0#
0(
#896520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#896570000000
0$
0)
#896580000000
1"
1'
b0 +
b0 1
#896630000000
0"
0'
#896640000000
1#
1(
b101111101100100 +
b101111101100100 1
#896690000000
0#
0(
#896700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#896750000000
0$
0)
#896760000000
1"
1'
b0 +
b0 1
#896810000000
0"
0'
#896820000000
1#
1(
b101111101100100 +
b101111101100100 1
#896870000000
0#
0(
#896880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#896930000000
0$
0)
#896940000000
1"
1'
b0 +
b0 1
#896990000000
0"
0'
#897000000000
1#
1(
b101111101100100 +
b101111101100100 1
#897050000000
0#
0(
#897060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#897110000000
0$
0)
#897120000000
1"
1'
b0 +
b0 1
#897170000000
0"
0'
#897180000000
1#
1(
b101111101100100 +
b101111101100100 1
#897230000000
0#
0(
#897240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#897290000000
0$
0)
#897300000000
1"
1'
b0 +
b0 1
#897350000000
0"
0'
#897360000000
1#
1(
b101111101100100 +
b101111101100100 1
#897410000000
0#
0(
#897420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#897470000000
0$
0)
#897480000000
1"
1'
b0 +
b0 1
#897530000000
0"
0'
#897540000000
1#
1(
b101111101100100 +
b101111101100100 1
#897590000000
0#
0(
#897600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#897650000000
0$
0)
#897660000000
1"
1'
b0 +
b0 1
#897710000000
0"
0'
#897720000000
1#
1(
b101111101100100 +
b101111101100100 1
#897770000000
0#
0(
#897780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#897830000000
0$
0)
#897840000000
1"
1'
b0 +
b0 1
#897890000000
0"
0'
#897900000000
1#
1(
b101111101100100 +
b101111101100100 1
#897950000000
0#
0(
#897960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#898010000000
0$
0)
#898020000000
1"
1'
b0 +
b0 1
#898070000000
0"
0'
#898080000000
1#
1(
b101111101100100 +
b101111101100100 1
#898130000000
0#
0(
#898140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#898190000000
0$
0)
#898200000000
1"
1'
b0 +
b0 1
#898250000000
0"
0'
#898260000000
1#
1(
b101111101100100 +
b101111101100100 1
#898310000000
0#
0(
#898320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#898370000000
0$
0)
#898380000000
1"
1'
b0 +
b0 1
#898430000000
0"
0'
#898440000000
1#
1(
b101111101100100 +
b101111101100100 1
#898490000000
0#
0(
#898500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#898550000000
0$
0)
#898560000000
1"
1'
b0 +
b0 1
#898610000000
0"
0'
#898620000000
1#
1(
b101111101100100 +
b101111101100100 1
#898670000000
0#
0(
#898680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#898730000000
0$
0)
#898740000000
1"
1'
b0 +
b0 1
#898790000000
0"
0'
#898800000000
1#
1(
b101111101100100 +
b101111101100100 1
#898850000000
0#
0(
#898860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#898910000000
0$
0)
#898920000000
1"
1'
b0 +
b0 1
#898970000000
0"
0'
#898980000000
1#
1(
b101111101100100 +
b101111101100100 1
#899030000000
0#
0(
#899040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#899090000000
0$
0)
#899100000000
1"
1'
b0 +
b0 1
#899150000000
0"
0'
#899160000000
1#
1(
b101111101100100 +
b101111101100100 1
#899210000000
0#
0(
#899220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#899270000000
0$
0)
#899280000000
1"
1'
b0 +
b0 1
#899330000000
0"
0'
#899340000000
1#
1(
b101111101100100 +
b101111101100100 1
#899390000000
0#
0(
#899400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#899450000000
0$
0)
#899460000000
1"
1'
b0 +
b0 1
#899510000000
0"
0'
#899520000000
1#
1(
b101111101100100 +
b101111101100100 1
#899570000000
0#
0(
#899580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#899630000000
0$
0)
#899640000000
1"
1'
b0 +
b0 1
#899690000000
0"
0'
#899700000000
1#
1(
b101111101100100 +
b101111101100100 1
#899750000000
0#
0(
#899760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#899810000000
0$
0)
#899820000000
1"
1'
b0 +
b0 1
#899870000000
0"
0'
#899880000000
1#
1(
b101111101100100 +
b101111101100100 1
#899930000000
0#
0(
#899940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#899990000000
0$
0)
#900000000000
1"
1'
b0 +
b0 1
#900050000000
0"
0'
#900060000000
1#
1(
b101111101100100 +
b101111101100100 1
#900110000000
0#
0(
#900120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#900170000000
0$
0)
#900180000000
1"
1'
b0 +
b0 1
#900230000000
0"
0'
#900240000000
1#
1(
b101111101100100 +
b101111101100100 1
#900290000000
0#
0(
#900300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#900350000000
0$
0)
#900360000000
1"
1'
b0 +
b0 1
#900410000000
0"
0'
#900420000000
1#
1(
b101111101100100 +
b101111101100100 1
#900470000000
0#
0(
#900480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#900530000000
0$
0)
#900540000000
1"
1'
b0 +
b0 1
#900590000000
0"
0'
#900600000000
1#
1(
b101111101100100 +
b101111101100100 1
#900650000000
0#
0(
#900660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#900710000000
0$
0)
#900720000000
1"
1'
b0 +
b0 1
#900770000000
0"
0'
#900780000000
1#
1(
b101111101100100 +
b101111101100100 1
#900830000000
0#
0(
#900840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#900890000000
0$
0)
#900900000000
1"
1'
b0 +
b0 1
#900950000000
0"
0'
#900960000000
1#
1(
b101111101100100 +
b101111101100100 1
#901010000000
0#
0(
#901020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#901070000000
0$
0)
#901080000000
1"
1'
b0 +
b0 1
#901130000000
0"
0'
#901140000000
1#
1(
b101111101100100 +
b101111101100100 1
#901190000000
0#
0(
#901200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#901250000000
0$
0)
#901260000000
1"
1'
b0 +
b0 1
#901310000000
0"
0'
#901320000000
1#
1(
b101111101100100 +
b101111101100100 1
#901370000000
0#
0(
#901380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#901430000000
0$
0)
#901440000000
1"
1'
b0 +
b0 1
#901490000000
0"
0'
#901500000000
1#
1(
b101111101100100 +
b101111101100100 1
#901550000000
0#
0(
#901560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#901610000000
0$
0)
#901620000000
1"
1'
b0 +
b0 1
#901670000000
0"
0'
#901680000000
1#
1(
b101111101100100 +
b101111101100100 1
#901730000000
0#
0(
#901740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#901790000000
0$
0)
#901800000000
1"
1'
b0 +
b0 1
#901850000000
0"
0'
#901860000000
1#
1(
b101111101100100 +
b101111101100100 1
#901910000000
0#
0(
#901920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#901970000000
0$
0)
#901980000000
1"
1'
b0 +
b0 1
#902030000000
0"
0'
#902040000000
1#
1(
b101111101100100 +
b101111101100100 1
#902090000000
0#
0(
#902100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#902150000000
0$
0)
#902160000000
1"
1'
b0 +
b0 1
#902210000000
0"
0'
#902220000000
1#
1(
b101111101100100 +
b101111101100100 1
#902270000000
0#
0(
#902280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#902330000000
0$
0)
#902340000000
1"
1'
b0 +
b0 1
#902390000000
0"
0'
#902400000000
1#
1(
b101111101100100 +
b101111101100100 1
#902450000000
0#
0(
#902460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#902510000000
0$
0)
#902520000000
1"
1'
b0 +
b0 1
#902570000000
0"
0'
#902580000000
1#
1(
b101111101100100 +
b101111101100100 1
#902630000000
0#
0(
#902640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#902690000000
0$
0)
#902700000000
1"
1'
b0 +
b0 1
#902750000000
0"
0'
#902760000000
1#
1(
b101111101100100 +
b101111101100100 1
#902810000000
0#
0(
#902820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#902870000000
0$
0)
#902880000000
1"
1'
b0 +
b0 1
#902930000000
0"
0'
#902940000000
1#
1(
b101111101100100 +
b101111101100100 1
#902990000000
0#
0(
#903000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#903050000000
0$
0)
#903060000000
1"
1'
b0 +
b0 1
#903110000000
0"
0'
#903120000000
1#
1(
b101111101100100 +
b101111101100100 1
#903170000000
0#
0(
#903180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#903230000000
0$
0)
#903240000000
1"
1'
b0 +
b0 1
#903290000000
0"
0'
#903300000000
1#
1(
b101111101100100 +
b101111101100100 1
#903350000000
0#
0(
#903360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#903410000000
0$
0)
#903420000000
1"
1'
b0 +
b0 1
#903470000000
0"
0'
#903480000000
1#
1(
b101111101100100 +
b101111101100100 1
#903530000000
0#
0(
#903540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#903590000000
0$
0)
#903600000000
1"
1'
b0 +
b0 1
#903650000000
0"
0'
#903660000000
1#
1(
b101111101100100 +
b101111101100100 1
#903710000000
0#
0(
#903720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#903770000000
0$
0)
#903780000000
1"
1'
b0 +
b0 1
#903830000000
0"
0'
#903840000000
1#
1(
b101111101100100 +
b101111101100100 1
#903890000000
0#
0(
#903900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#903950000000
0$
0)
#903960000000
1"
1'
b0 +
b0 1
#904010000000
0"
0'
#904020000000
1#
1(
b101111101100100 +
b101111101100100 1
#904070000000
0#
0(
#904080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#904130000000
0$
0)
#904140000000
1"
1'
b0 +
b0 1
#904190000000
0"
0'
#904200000000
1#
1(
b101111101100100 +
b101111101100100 1
#904250000000
0#
0(
#904260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#904310000000
0$
0)
#904320000000
1"
1'
b0 +
b0 1
#904370000000
0"
0'
#904380000000
1#
1(
b101111101100100 +
b101111101100100 1
#904430000000
0#
0(
#904440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#904490000000
0$
0)
#904500000000
1"
1'
b0 +
b0 1
#904550000000
0"
0'
#904560000000
1#
1(
b101111101100100 +
b101111101100100 1
#904610000000
0#
0(
#904620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#904670000000
0$
0)
#904680000000
1"
1'
b0 +
b0 1
#904730000000
0"
0'
#904740000000
1#
1(
b101111101100100 +
b101111101100100 1
#904790000000
0#
0(
#904800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#904850000000
0$
0)
#904860000000
1"
1'
b0 +
b0 1
#904910000000
0"
0'
#904920000000
1#
1(
b101111101100100 +
b101111101100100 1
#904970000000
0#
0(
#904980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#905030000000
0$
0)
#905040000000
1"
1'
b0 +
b0 1
#905090000000
0"
0'
#905100000000
1#
1(
b101111101100100 +
b101111101100100 1
#905150000000
0#
0(
#905160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#905210000000
0$
0)
#905220000000
1"
1'
b0 +
b0 1
#905270000000
0"
0'
#905280000000
1#
1(
b101111101100100 +
b101111101100100 1
#905330000000
0#
0(
#905340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#905390000000
0$
0)
#905400000000
1"
1'
b0 +
b0 1
#905450000000
0"
0'
#905460000000
1#
1(
b101111101100100 +
b101111101100100 1
#905510000000
0#
0(
#905520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#905570000000
0$
0)
#905580000000
1"
1'
b0 +
b0 1
#905630000000
0"
0'
#905640000000
1#
1(
b101111101100100 +
b101111101100100 1
#905690000000
0#
0(
#905700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#905750000000
0$
0)
#905760000000
1"
1'
b0 +
b0 1
#905810000000
0"
0'
#905820000000
1#
1(
b101111101100100 +
b101111101100100 1
#905870000000
0#
0(
#905880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#905930000000
0$
0)
#905940000000
1"
1'
b0 +
b0 1
#905990000000
0"
0'
#906000000000
1#
1(
b101111101100100 +
b101111101100100 1
#906050000000
0#
0(
#906060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#906110000000
0$
0)
#906120000000
1"
1'
b0 +
b0 1
#906170000000
0"
0'
#906180000000
1#
1(
b101111101100100 +
b101111101100100 1
#906230000000
0#
0(
#906240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#906290000000
0$
0)
#906300000000
1"
1'
b0 +
b0 1
#906350000000
0"
0'
#906360000000
1#
1(
b101111101100100 +
b101111101100100 1
#906410000000
0#
0(
#906420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#906470000000
0$
0)
#906480000000
1"
1'
b0 +
b0 1
#906530000000
0"
0'
#906540000000
1#
1(
b101111101100100 +
b101111101100100 1
#906590000000
0#
0(
#906600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#906650000000
0$
0)
#906660000000
1"
1'
b0 +
b0 1
#906710000000
0"
0'
#906720000000
1#
1(
b101111101100100 +
b101111101100100 1
#906770000000
0#
0(
#906780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#906830000000
0$
0)
#906840000000
1"
1'
b0 +
b0 1
#906890000000
0"
0'
#906900000000
1#
1(
b101111101100100 +
b101111101100100 1
#906950000000
0#
0(
#906960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#907010000000
0$
0)
#907020000000
1"
1'
b0 +
b0 1
#907070000000
0"
0'
#907080000000
1#
1(
b101111101100100 +
b101111101100100 1
#907130000000
0#
0(
#907140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#907190000000
0$
0)
#907200000000
1"
1'
b0 +
b0 1
#907250000000
0"
0'
#907260000000
1#
1(
b101111101100100 +
b101111101100100 1
#907310000000
0#
0(
#907320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#907370000000
0$
0)
#907380000000
1"
1'
b0 +
b0 1
#907430000000
0"
0'
#907440000000
1#
1(
b101111101100100 +
b101111101100100 1
#907490000000
0#
0(
#907500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#907550000000
0$
0)
#907560000000
1"
1'
b0 +
b0 1
#907610000000
0"
0'
#907620000000
1#
1(
b101111101100100 +
b101111101100100 1
#907670000000
0#
0(
#907680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#907730000000
0$
0)
#907740000000
1"
1'
b0 +
b0 1
#907790000000
0"
0'
#907800000000
1#
1(
b101111101100100 +
b101111101100100 1
#907850000000
0#
0(
#907860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#907910000000
0$
0)
#907920000000
1"
1'
b0 +
b0 1
#907970000000
0"
0'
#907980000000
1#
1(
b101111101100100 +
b101111101100100 1
#908030000000
0#
0(
#908040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#908090000000
0$
0)
#908100000000
1"
1'
b0 +
b0 1
#908150000000
0"
0'
#908160000000
1#
1(
b101111101100100 +
b101111101100100 1
#908210000000
0#
0(
#908220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#908270000000
0$
0)
#908280000000
1"
1'
b0 +
b0 1
#908330000000
0"
0'
#908340000000
1#
1(
b101111101100100 +
b101111101100100 1
#908390000000
0#
0(
#908400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#908450000000
0$
0)
#908460000000
1"
1'
b0 +
b0 1
#908510000000
0"
0'
#908520000000
1#
1(
b101111101100100 +
b101111101100100 1
#908570000000
0#
0(
#908580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#908630000000
0$
0)
#908640000000
1"
1'
b0 +
b0 1
#908690000000
0"
0'
#908700000000
1#
1(
b101111101100100 +
b101111101100100 1
#908750000000
0#
0(
#908760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#908810000000
0$
0)
#908820000000
1"
1'
b0 +
b0 1
#908870000000
0"
0'
#908880000000
1#
1(
b101111101100100 +
b101111101100100 1
#908930000000
0#
0(
#908940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#908990000000
0$
0)
#909000000000
1"
1'
b0 +
b0 1
#909050000000
0"
0'
#909060000000
1#
1(
b101111101100100 +
b101111101100100 1
#909110000000
0#
0(
#909120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#909170000000
0$
0)
#909180000000
1"
1'
b0 +
b0 1
#909230000000
0"
0'
#909240000000
1#
1(
b101111101100100 +
b101111101100100 1
#909290000000
0#
0(
#909300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#909350000000
0$
0)
#909360000000
1"
1'
b0 +
b0 1
#909410000000
0"
0'
#909420000000
1#
1(
b101111101100100 +
b101111101100100 1
#909470000000
0#
0(
#909480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#909530000000
0$
0)
#909540000000
1"
1'
b0 +
b0 1
#909590000000
0"
0'
#909600000000
1#
1(
b101111101100100 +
b101111101100100 1
#909650000000
0#
0(
#909660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#909710000000
0$
0)
#909720000000
1"
1'
b0 +
b0 1
#909770000000
0"
0'
#909780000000
1#
1(
b101111101100100 +
b101111101100100 1
#909830000000
0#
0(
#909840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#909890000000
0$
0)
#909900000000
1"
1'
b0 +
b0 1
#909950000000
0"
0'
#909960000000
1#
1(
b101111101100100 +
b101111101100100 1
#910010000000
0#
0(
#910020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#910070000000
0$
0)
#910080000000
1"
1'
b0 +
b0 1
#910130000000
0"
0'
#910140000000
1#
1(
b101111101100100 +
b101111101100100 1
#910190000000
0#
0(
#910200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#910250000000
0$
0)
#910260000000
1"
1'
b0 +
b0 1
#910310000000
0"
0'
#910320000000
1#
1(
b101111101100100 +
b101111101100100 1
#910370000000
0#
0(
#910380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#910430000000
0$
0)
#910440000000
1"
1'
b0 +
b0 1
#910490000000
0"
0'
#910500000000
1#
1(
b101111101100100 +
b101111101100100 1
#910550000000
0#
0(
#910560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#910610000000
0$
0)
#910620000000
1"
1'
b0 +
b0 1
#910670000000
0"
0'
#910680000000
1#
1(
b101111101100100 +
b101111101100100 1
#910730000000
0#
0(
#910740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#910790000000
0$
0)
#910800000000
1"
1'
b0 +
b0 1
#910850000000
0"
0'
#910860000000
1#
1(
b101111101100100 +
b101111101100100 1
#910910000000
0#
0(
#910920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#910970000000
0$
0)
#910980000000
1"
1'
b0 +
b0 1
#911030000000
0"
0'
#911040000000
1#
1(
b101111101100100 +
b101111101100100 1
#911090000000
0#
0(
#911100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#911150000000
0$
0)
#911160000000
1"
1'
b0 +
b0 1
#911210000000
0"
0'
#911220000000
1#
1(
b101111101100100 +
b101111101100100 1
#911270000000
0#
0(
#911280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#911330000000
0$
0)
#911340000000
1"
1'
b0 +
b0 1
#911390000000
0"
0'
#911400000000
1#
1(
b101111101100100 +
b101111101100100 1
#911450000000
0#
0(
#911460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#911510000000
0$
0)
#911520000000
1"
1'
b0 +
b0 1
#911570000000
0"
0'
#911580000000
1#
1(
b101111101100100 +
b101111101100100 1
#911630000000
0#
0(
#911640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#911690000000
0$
0)
#911700000000
1"
1'
b0 +
b0 1
#911750000000
0"
0'
#911760000000
1#
1(
b101111101100100 +
b101111101100100 1
#911810000000
0#
0(
#911820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#911870000000
0$
0)
#911880000000
1"
1'
b0 +
b0 1
#911930000000
0"
0'
#911940000000
1#
1(
b101111101100100 +
b101111101100100 1
#911990000000
0#
0(
#912000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#912050000000
0$
0)
#912060000000
1"
1'
b0 +
b0 1
#912110000000
0"
0'
#912120000000
1#
1(
b101111101100100 +
b101111101100100 1
#912170000000
0#
0(
#912180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#912230000000
0$
0)
#912240000000
1"
1'
b0 +
b0 1
#912290000000
0"
0'
#912300000000
1#
1(
b101111101100100 +
b101111101100100 1
#912350000000
0#
0(
#912360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#912410000000
0$
0)
#912420000000
1"
1'
b0 +
b0 1
#912470000000
0"
0'
#912480000000
1#
1(
b101111101100100 +
b101111101100100 1
#912530000000
0#
0(
#912540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#912590000000
0$
0)
#912600000000
1"
1'
b0 +
b0 1
#912650000000
0"
0'
#912660000000
1#
1(
b101111101100100 +
b101111101100100 1
#912710000000
0#
0(
#912720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#912770000000
0$
0)
#912780000000
1"
1'
b0 +
b0 1
#912830000000
0"
0'
#912840000000
1#
1(
b101111101100100 +
b101111101100100 1
#912890000000
0#
0(
#912900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#912950000000
0$
0)
#912960000000
1"
1'
b0 +
b0 1
#913010000000
0"
0'
#913020000000
1#
1(
b101111101100100 +
b101111101100100 1
#913070000000
0#
0(
#913080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#913130000000
0$
0)
#913140000000
1"
1'
b0 +
b0 1
#913190000000
0"
0'
#913200000000
1#
1(
b101111101100100 +
b101111101100100 1
#913250000000
0#
0(
#913260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#913310000000
0$
0)
#913320000000
1"
1'
b0 +
b0 1
#913370000000
0"
0'
#913380000000
1#
1(
b101111101100100 +
b101111101100100 1
#913430000000
0#
0(
#913440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#913490000000
0$
0)
#913500000000
1"
1'
b0 +
b0 1
#913550000000
0"
0'
#913560000000
1#
1(
b101111101100100 +
b101111101100100 1
#913610000000
0#
0(
#913620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#913670000000
0$
0)
#913680000000
1"
1'
b0 +
b0 1
#913730000000
0"
0'
#913740000000
1#
1(
b101111101100100 +
b101111101100100 1
#913790000000
0#
0(
#913800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#913850000000
0$
0)
#913860000000
1"
1'
b0 +
b0 1
#913910000000
0"
0'
#913920000000
1#
1(
b101111101100100 +
b101111101100100 1
#913970000000
0#
0(
#913980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#914030000000
0$
0)
#914040000000
1"
1'
b0 +
b0 1
#914090000000
0"
0'
#914100000000
1#
1(
b101111101100100 +
b101111101100100 1
#914150000000
0#
0(
#914160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#914210000000
0$
0)
#914220000000
1"
1'
b0 +
b0 1
#914270000000
0"
0'
#914280000000
1#
1(
b101111101100100 +
b101111101100100 1
#914330000000
0#
0(
#914340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#914390000000
0$
0)
#914400000000
1"
1'
b0 +
b0 1
#914450000000
0"
0'
#914460000000
1#
1(
b101111101100100 +
b101111101100100 1
#914510000000
0#
0(
#914520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#914570000000
0$
0)
#914580000000
1"
1'
b0 +
b0 1
#914630000000
0"
0'
#914640000000
1#
1(
b101111101100100 +
b101111101100100 1
#914690000000
0#
0(
#914700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#914750000000
0$
0)
#914760000000
1"
1'
b0 +
b0 1
#914810000000
0"
0'
#914820000000
1#
1(
b101111101100100 +
b101111101100100 1
#914870000000
0#
0(
#914880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#914930000000
0$
0)
#914940000000
1"
1'
b0 +
b0 1
#914990000000
0"
0'
#915000000000
1#
1(
b101111101100100 +
b101111101100100 1
#915050000000
0#
0(
#915060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#915110000000
0$
0)
#915120000000
1"
1'
b0 +
b0 1
#915170000000
0"
0'
#915180000000
1#
1(
b101111101100100 +
b101111101100100 1
#915230000000
0#
0(
#915240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#915290000000
0$
0)
#915300000000
1"
1'
b0 +
b0 1
#915350000000
0"
0'
#915360000000
1#
1(
b101111101100100 +
b101111101100100 1
#915410000000
0#
0(
#915420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#915470000000
0$
0)
#915480000000
1"
1'
b0 +
b0 1
#915530000000
0"
0'
#915540000000
1#
1(
b101111101100100 +
b101111101100100 1
#915590000000
0#
0(
#915600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#915650000000
0$
0)
#915660000000
1"
1'
b0 +
b0 1
#915710000000
0"
0'
#915720000000
1#
1(
b101111101100100 +
b101111101100100 1
#915770000000
0#
0(
#915780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#915830000000
0$
0)
#915840000000
1"
1'
b0 +
b0 1
#915890000000
0"
0'
#915900000000
1#
1(
b101111101100100 +
b101111101100100 1
#915950000000
0#
0(
#915960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#916010000000
0$
0)
#916020000000
1"
1'
b0 +
b0 1
#916070000000
0"
0'
#916080000000
1#
1(
b101111101100100 +
b101111101100100 1
#916130000000
0#
0(
#916140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#916190000000
0$
0)
#916200000000
1"
1'
b0 +
b0 1
#916250000000
0"
0'
#916260000000
1#
1(
b101111101100100 +
b101111101100100 1
#916310000000
0#
0(
#916320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#916370000000
0$
0)
#916380000000
1"
1'
b0 +
b0 1
#916430000000
0"
0'
#916440000000
1#
1(
b101111101100100 +
b101111101100100 1
#916490000000
0#
0(
#916500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#916550000000
0$
0)
#916560000000
1"
1'
b0 +
b0 1
#916610000000
0"
0'
#916620000000
1#
1(
b101111101100100 +
b101111101100100 1
#916670000000
0#
0(
#916680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#916730000000
0$
0)
#916740000000
1"
1'
b0 +
b0 1
#916790000000
0"
0'
#916800000000
1#
1(
b101111101100100 +
b101111101100100 1
#916850000000
0#
0(
#916860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#916910000000
0$
0)
#916920000000
1"
1'
b0 +
b0 1
#916970000000
0"
0'
#916980000000
1#
1(
b101111101100100 +
b101111101100100 1
#917030000000
0#
0(
#917040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#917090000000
0$
0)
#917100000000
1"
1'
b0 +
b0 1
#917150000000
0"
0'
#917160000000
1#
1(
b101111101100100 +
b101111101100100 1
#917210000000
0#
0(
#917220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#917270000000
0$
0)
#917280000000
1"
1'
b0 +
b0 1
#917330000000
0"
0'
#917340000000
1#
1(
b101111101100100 +
b101111101100100 1
#917390000000
0#
0(
#917400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#917450000000
0$
0)
#917460000000
1"
1'
b0 +
b0 1
#917510000000
0"
0'
#917520000000
1#
1(
b101111101100100 +
b101111101100100 1
#917570000000
0#
0(
#917580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#917630000000
0$
0)
#917640000000
1"
1'
b0 +
b0 1
#917690000000
0"
0'
#917700000000
1#
1(
b101111101100100 +
b101111101100100 1
#917750000000
0#
0(
#917760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#917810000000
0$
0)
#917820000000
1"
1'
b0 +
b0 1
#917870000000
0"
0'
#917880000000
1#
1(
b101111101100100 +
b101111101100100 1
#917930000000
0#
0(
#917940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#917990000000
0$
0)
#918000000000
1"
1'
b0 +
b0 1
#918050000000
0"
0'
#918060000000
1#
1(
b101111101100100 +
b101111101100100 1
#918110000000
0#
0(
#918120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#918170000000
0$
0)
#918180000000
1"
1'
b0 +
b0 1
#918230000000
0"
0'
#918240000000
1#
1(
b101111101100100 +
b101111101100100 1
#918290000000
0#
0(
#918300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#918350000000
0$
0)
#918360000000
1"
1'
b0 +
b0 1
#918410000000
0"
0'
#918420000000
1#
1(
b101111101100100 +
b101111101100100 1
#918470000000
0#
0(
#918480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#918530000000
0$
0)
#918540000000
1"
1'
b0 +
b0 1
#918590000000
0"
0'
#918600000000
1#
1(
b101111101100100 +
b101111101100100 1
#918650000000
0#
0(
#918660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#918710000000
0$
0)
#918720000000
1"
1'
b0 +
b0 1
#918770000000
0"
0'
#918780000000
1#
1(
b101111101100100 +
b101111101100100 1
#918830000000
0#
0(
#918840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#918890000000
0$
0)
#918900000000
1"
1'
b0 +
b0 1
#918950000000
0"
0'
#918960000000
1#
1(
b101111101100100 +
b101111101100100 1
#919010000000
0#
0(
#919020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#919070000000
0$
0)
#919080000000
1"
1'
b0 +
b0 1
#919130000000
0"
0'
#919140000000
1#
1(
b101111101100100 +
b101111101100100 1
#919190000000
0#
0(
#919200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#919250000000
0$
0)
#919260000000
1"
1'
b0 +
b0 1
#919310000000
0"
0'
#919320000000
1#
1(
b101111101100100 +
b101111101100100 1
#919370000000
0#
0(
#919380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#919430000000
0$
0)
#919440000000
1"
1'
b0 +
b0 1
#919490000000
0"
0'
#919500000000
1#
1(
b101111101100100 +
b101111101100100 1
#919550000000
0#
0(
#919560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#919610000000
0$
0)
#919620000000
1"
1'
b0 +
b0 1
#919670000000
0"
0'
#919680000000
1#
1(
b101111101100100 +
b101111101100100 1
#919730000000
0#
0(
#919740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#919790000000
0$
0)
#919800000000
1"
1'
b0 +
b0 1
#919850000000
0"
0'
#919860000000
1#
1(
b101111101100100 +
b101111101100100 1
#919910000000
0#
0(
#919920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#919970000000
0$
0)
#919980000000
1"
1'
b0 +
b0 1
#920030000000
0"
0'
#920040000000
1#
1(
b101111101100100 +
b101111101100100 1
#920090000000
0#
0(
#920100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#920150000000
0$
0)
#920160000000
1"
1'
b0 +
b0 1
#920210000000
0"
0'
#920220000000
1#
1(
b101111101100100 +
b101111101100100 1
#920270000000
0#
0(
#920280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#920330000000
0$
0)
#920340000000
1"
1'
b0 +
b0 1
#920390000000
0"
0'
#920400000000
1#
1(
b101111101100100 +
b101111101100100 1
#920450000000
0#
0(
#920460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#920510000000
0$
0)
#920520000000
1"
1'
b0 +
b0 1
#920570000000
0"
0'
#920580000000
1#
1(
b101111101100100 +
b101111101100100 1
#920630000000
0#
0(
#920640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#920690000000
0$
0)
#920700000000
1"
1'
b0 +
b0 1
#920750000000
0"
0'
#920760000000
1#
1(
b101111101100100 +
b101111101100100 1
#920810000000
0#
0(
#920820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#920870000000
0$
0)
#920880000000
1"
1'
b0 +
b0 1
#920930000000
0"
0'
#920940000000
1#
1(
b101111101100100 +
b101111101100100 1
#920990000000
0#
0(
#921000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#921050000000
0$
0)
#921060000000
1"
1'
b0 +
b0 1
#921110000000
0"
0'
#921120000000
1#
1(
b101111101100100 +
b101111101100100 1
#921170000000
0#
0(
#921180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#921230000000
0$
0)
#921240000000
1"
1'
b0 +
b0 1
#921290000000
0"
0'
#921300000000
1#
1(
b101111101100100 +
b101111101100100 1
#921350000000
0#
0(
#921360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#921410000000
0$
0)
#921420000000
1"
1'
b0 +
b0 1
#921470000000
0"
0'
#921480000000
1#
1(
b101111101100100 +
b101111101100100 1
#921530000000
0#
0(
#921540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#921590000000
0$
0)
#921600000000
1"
1'
b0 +
b0 1
#921650000000
0"
0'
#921660000000
1#
1(
b101111101100100 +
b101111101100100 1
#921710000000
0#
0(
#921720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#921770000000
0$
0)
#921780000000
1"
1'
b0 +
b0 1
#921830000000
0"
0'
#921840000000
1#
1(
b101111101100100 +
b101111101100100 1
#921890000000
0#
0(
#921900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#921950000000
0$
0)
#921960000000
1"
1'
b0 +
b0 1
#922010000000
0"
0'
#922020000000
1#
1(
b101111101100100 +
b101111101100100 1
#922070000000
0#
0(
#922080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#922130000000
0$
0)
#922140000000
1"
1'
b0 +
b0 1
#922190000000
0"
0'
#922200000000
1#
1(
b101111101100100 +
b101111101100100 1
#922250000000
0#
0(
#922260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#922310000000
0$
0)
#922320000000
1"
1'
b0 +
b0 1
#922370000000
0"
0'
#922380000000
1#
1(
b101111101100100 +
b101111101100100 1
#922430000000
0#
0(
#922440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#922490000000
0$
0)
#922500000000
1"
1'
b0 +
b0 1
#922550000000
0"
0'
#922560000000
1#
1(
b101111101100100 +
b101111101100100 1
#922610000000
0#
0(
#922620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#922670000000
0$
0)
#922680000000
1"
1'
b0 +
b0 1
#922730000000
0"
0'
#922740000000
1#
1(
b101111101100100 +
b101111101100100 1
#922790000000
0#
0(
#922800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#922850000000
0$
0)
#922860000000
1"
1'
b0 +
b0 1
#922910000000
0"
0'
#922920000000
1#
1(
b101111101100100 +
b101111101100100 1
#922970000000
0#
0(
#922980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#923030000000
0$
0)
#923040000000
1"
1'
b0 +
b0 1
#923090000000
0"
0'
#923100000000
1#
1(
b101111101100100 +
b101111101100100 1
#923150000000
0#
0(
#923160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#923210000000
0$
0)
#923220000000
1"
1'
b0 +
b0 1
#923270000000
0"
0'
#923280000000
1#
1(
b101111101100100 +
b101111101100100 1
#923330000000
0#
0(
#923340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#923390000000
0$
0)
#923400000000
1"
1'
b0 +
b0 1
#923450000000
0"
0'
#923460000000
1#
1(
b101111101100100 +
b101111101100100 1
#923510000000
0#
0(
#923520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#923570000000
0$
0)
#923580000000
1"
1'
b0 +
b0 1
#923630000000
0"
0'
#923640000000
1#
1(
b101111101100100 +
b101111101100100 1
#923690000000
0#
0(
#923700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#923750000000
0$
0)
#923760000000
1"
1'
b0 +
b0 1
#923810000000
0"
0'
#923820000000
1#
1(
b101111101100100 +
b101111101100100 1
#923870000000
0#
0(
#923880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#923930000000
0$
0)
#923940000000
1"
1'
b0 +
b0 1
#923990000000
0"
0'
#924000000000
1#
1(
b101111101100100 +
b101111101100100 1
#924050000000
0#
0(
#924060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#924110000000
0$
0)
#924120000000
1"
1'
b0 +
b0 1
#924170000000
0"
0'
#924180000000
1#
1(
b101111101100100 +
b101111101100100 1
#924230000000
0#
0(
#924240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#924290000000
0$
0)
#924300000000
1"
1'
b0 +
b0 1
#924350000000
0"
0'
#924360000000
1#
1(
b101111101100100 +
b101111101100100 1
#924410000000
0#
0(
#924420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#924470000000
0$
0)
#924480000000
1"
1'
b0 +
b0 1
#924530000000
0"
0'
#924540000000
1#
1(
b101111101100100 +
b101111101100100 1
#924590000000
0#
0(
#924600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#924650000000
0$
0)
#924660000000
1"
1'
b0 +
b0 1
#924710000000
0"
0'
#924720000000
1#
1(
b101111101100100 +
b101111101100100 1
#924770000000
0#
0(
#924780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#924830000000
0$
0)
#924840000000
1"
1'
b0 +
b0 1
#924890000000
0"
0'
#924900000000
1#
1(
b101111101100100 +
b101111101100100 1
#924950000000
0#
0(
#924960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#925010000000
0$
0)
#925020000000
1"
1'
b0 +
b0 1
#925070000000
0"
0'
#925080000000
1#
1(
b101111101100100 +
b101111101100100 1
#925130000000
0#
0(
#925140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#925190000000
0$
0)
#925200000000
1"
1'
b0 +
b0 1
#925250000000
0"
0'
#925260000000
1#
1(
b101111101100100 +
b101111101100100 1
#925310000000
0#
0(
#925320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#925370000000
0$
0)
#925380000000
1"
1'
b0 +
b0 1
#925430000000
0"
0'
#925440000000
1#
1(
b101111101100100 +
b101111101100100 1
#925490000000
0#
0(
#925500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#925550000000
0$
0)
#925560000000
1"
1'
b0 +
b0 1
#925610000000
0"
0'
#925620000000
1#
1(
b101111101100100 +
b101111101100100 1
#925670000000
0#
0(
#925680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#925730000000
0$
0)
#925740000000
1"
1'
b0 +
b0 1
#925790000000
0"
0'
#925800000000
1#
1(
b101111101100100 +
b101111101100100 1
#925850000000
0#
0(
#925860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#925910000000
0$
0)
#925920000000
1"
1'
b0 +
b0 1
#925970000000
0"
0'
#925980000000
1#
1(
b101111101100100 +
b101111101100100 1
#926030000000
0#
0(
#926040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#926090000000
0$
0)
#926100000000
1"
1'
b0 +
b0 1
#926150000000
0"
0'
#926160000000
1#
1(
b101111101100100 +
b101111101100100 1
#926210000000
0#
0(
#926220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#926270000000
0$
0)
#926280000000
1"
1'
b0 +
b0 1
#926330000000
0"
0'
#926340000000
1#
1(
b101111101100100 +
b101111101100100 1
#926390000000
0#
0(
#926400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#926450000000
0$
0)
#926460000000
1"
1'
b0 +
b0 1
#926510000000
0"
0'
#926520000000
1#
1(
b101111101100100 +
b101111101100100 1
#926570000000
0#
0(
#926580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#926630000000
0$
0)
#926640000000
1"
1'
b0 +
b0 1
#926690000000
0"
0'
#926700000000
1#
1(
b101111101100100 +
b101111101100100 1
#926750000000
0#
0(
#926760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#926810000000
0$
0)
#926820000000
1"
1'
b0 +
b0 1
#926870000000
0"
0'
#926880000000
1#
1(
b101111101100100 +
b101111101100100 1
#926930000000
0#
0(
#926940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#926990000000
0$
0)
#927000000000
1"
1'
b0 +
b0 1
#927050000000
0"
0'
#927060000000
1#
1(
b101111101100100 +
b101111101100100 1
#927110000000
0#
0(
#927120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#927170000000
0$
0)
#927180000000
1"
1'
b0 +
b0 1
#927230000000
0"
0'
#927240000000
1#
1(
b101111101100100 +
b101111101100100 1
#927290000000
0#
0(
#927300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#927350000000
0$
0)
#927360000000
1"
1'
b0 +
b0 1
#927410000000
0"
0'
#927420000000
1#
1(
b101111101100100 +
b101111101100100 1
#927470000000
0#
0(
#927480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#927530000000
0$
0)
#927540000000
1"
1'
b0 +
b0 1
#927590000000
0"
0'
#927600000000
1#
1(
b101111101100100 +
b101111101100100 1
#927650000000
0#
0(
#927660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#927710000000
0$
0)
#927720000000
1"
1'
b0 +
b0 1
#927770000000
0"
0'
#927780000000
1#
1(
b101111101100100 +
b101111101100100 1
#927830000000
0#
0(
#927840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#927890000000
0$
0)
#927900000000
1"
1'
b0 +
b0 1
#927950000000
0"
0'
#927960000000
1#
1(
b101111101100100 +
b101111101100100 1
#928010000000
0#
0(
#928020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#928070000000
0$
0)
#928080000000
1"
1'
b0 +
b0 1
#928130000000
0"
0'
#928140000000
1#
1(
b101111101100100 +
b101111101100100 1
#928190000000
0#
0(
#928200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#928250000000
0$
0)
#928260000000
1"
1'
b0 +
b0 1
#928310000000
0"
0'
#928320000000
1#
1(
b101111101100100 +
b101111101100100 1
#928370000000
0#
0(
#928380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#928430000000
0$
0)
#928440000000
1"
1'
b0 +
b0 1
#928490000000
0"
0'
#928500000000
1#
1(
b101111101100100 +
b101111101100100 1
#928550000000
0#
0(
#928560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#928610000000
0$
0)
#928620000000
1"
1'
b0 +
b0 1
#928670000000
0"
0'
#928680000000
1#
1(
b101111101100100 +
b101111101100100 1
#928730000000
0#
0(
#928740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#928790000000
0$
0)
#928800000000
1"
1'
b0 +
b0 1
#928850000000
0"
0'
#928860000000
1#
1(
b101111101100100 +
b101111101100100 1
#928910000000
0#
0(
#928920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#928970000000
0$
0)
#928980000000
1"
1'
b0 +
b0 1
#929030000000
0"
0'
#929040000000
1#
1(
b101111101100100 +
b101111101100100 1
#929090000000
0#
0(
#929100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#929150000000
0$
0)
#929160000000
1"
1'
b0 +
b0 1
#929210000000
0"
0'
#929220000000
1#
1(
b101111101100100 +
b101111101100100 1
#929270000000
0#
0(
#929280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#929330000000
0$
0)
#929340000000
1"
1'
b0 +
b0 1
#929390000000
0"
0'
#929400000000
1#
1(
b101111101100100 +
b101111101100100 1
#929450000000
0#
0(
#929460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#929510000000
0$
0)
#929520000000
1"
1'
b0 +
b0 1
#929570000000
0"
0'
#929580000000
1#
1(
b101111101100100 +
b101111101100100 1
#929630000000
0#
0(
#929640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#929690000000
0$
0)
#929700000000
1"
1'
b0 +
b0 1
#929750000000
0"
0'
#929760000000
1#
1(
b101111101100100 +
b101111101100100 1
#929810000000
0#
0(
#929820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#929870000000
0$
0)
#929880000000
1"
1'
b0 +
b0 1
#929930000000
0"
0'
#929940000000
1#
1(
b101111101100100 +
b101111101100100 1
#929990000000
0#
0(
#930000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#930050000000
0$
0)
#930060000000
1"
1'
b0 +
b0 1
#930110000000
0"
0'
#930120000000
1#
1(
b101111101100100 +
b101111101100100 1
#930170000000
0#
0(
#930180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#930230000000
0$
0)
#930240000000
1"
1'
b0 +
b0 1
#930290000000
0"
0'
#930300000000
1#
1(
b101111101100100 +
b101111101100100 1
#930350000000
0#
0(
#930360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#930410000000
0$
0)
#930420000000
1"
1'
b0 +
b0 1
#930470000000
0"
0'
#930480000000
1#
1(
b101111101100100 +
b101111101100100 1
#930530000000
0#
0(
#930540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#930590000000
0$
0)
#930600000000
1"
1'
b0 +
b0 1
#930650000000
0"
0'
#930660000000
1#
1(
b101111101100100 +
b101111101100100 1
#930710000000
0#
0(
#930720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#930770000000
0$
0)
#930780000000
1"
1'
b0 +
b0 1
#930830000000
0"
0'
#930840000000
1#
1(
b101111101100100 +
b101111101100100 1
#930890000000
0#
0(
#930900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#930950000000
0$
0)
#930960000000
1"
1'
b0 +
b0 1
#931010000000
0"
0'
#931020000000
1#
1(
b101111101100100 +
b101111101100100 1
#931070000000
0#
0(
#931080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#931130000000
0$
0)
#931140000000
1"
1'
b0 +
b0 1
#931190000000
0"
0'
#931200000000
1#
1(
b101111101100100 +
b101111101100100 1
#931250000000
0#
0(
#931260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#931310000000
0$
0)
#931320000000
1"
1'
b0 +
b0 1
#931370000000
0"
0'
#931380000000
1#
1(
b101111101100100 +
b101111101100100 1
#931430000000
0#
0(
#931440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#931490000000
0$
0)
#931500000000
1"
1'
b0 +
b0 1
#931550000000
0"
0'
#931560000000
1#
1(
b101111101100100 +
b101111101100100 1
#931610000000
0#
0(
#931620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#931670000000
0$
0)
#931680000000
1"
1'
b0 +
b0 1
#931730000000
0"
0'
#931740000000
1#
1(
b101111101100100 +
b101111101100100 1
#931790000000
0#
0(
#931800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#931850000000
0$
0)
#931860000000
1"
1'
b0 +
b0 1
#931910000000
0"
0'
#931920000000
1#
1(
b101111101100100 +
b101111101100100 1
#931970000000
0#
0(
#931980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#932030000000
0$
0)
#932040000000
1"
1'
b0 +
b0 1
#932090000000
0"
0'
#932100000000
1#
1(
b101111101100100 +
b101111101100100 1
#932150000000
0#
0(
#932160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#932210000000
0$
0)
#932220000000
1"
1'
b0 +
b0 1
#932270000000
0"
0'
#932280000000
1#
1(
b101111101100100 +
b101111101100100 1
#932330000000
0#
0(
#932340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#932390000000
0$
0)
#932400000000
1"
1'
b0 +
b0 1
#932450000000
0"
0'
#932460000000
1#
1(
b101111101100100 +
b101111101100100 1
#932510000000
0#
0(
#932520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#932570000000
0$
0)
#932580000000
1"
1'
b0 +
b0 1
#932630000000
0"
0'
#932640000000
1#
1(
b101111101100100 +
b101111101100100 1
#932690000000
0#
0(
#932700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#932750000000
0$
0)
#932760000000
1"
1'
b0 +
b0 1
#932810000000
0"
0'
#932820000000
1#
1(
b101111101100100 +
b101111101100100 1
#932870000000
0#
0(
#932880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#932930000000
0$
0)
#932940000000
1"
1'
b0 +
b0 1
#932990000000
0"
0'
#933000000000
1#
1(
b101111101100100 +
b101111101100100 1
#933050000000
0#
0(
#933060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#933110000000
0$
0)
#933120000000
1"
1'
b0 +
b0 1
#933170000000
0"
0'
#933180000000
1#
1(
b101111101100100 +
b101111101100100 1
#933230000000
0#
0(
#933240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#933290000000
0$
0)
#933300000000
1"
1'
b0 +
b0 1
#933350000000
0"
0'
#933360000000
1#
1(
b101111101100100 +
b101111101100100 1
#933410000000
0#
0(
#933420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#933470000000
0$
0)
#933480000000
1"
1'
b0 +
b0 1
#933530000000
0"
0'
#933540000000
1#
1(
b101111101100100 +
b101111101100100 1
#933590000000
0#
0(
#933600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#933650000000
0$
0)
#933660000000
1"
1'
b0 +
b0 1
#933710000000
0"
0'
#933720000000
1#
1(
b101111101100100 +
b101111101100100 1
#933770000000
0#
0(
#933780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#933830000000
0$
0)
#933840000000
1"
1'
b0 +
b0 1
#933890000000
0"
0'
#933900000000
1#
1(
b101111101100100 +
b101111101100100 1
#933950000000
0#
0(
#933960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#934010000000
0$
0)
#934020000000
1"
1'
b0 +
b0 1
#934070000000
0"
0'
#934080000000
1#
1(
b101111101100100 +
b101111101100100 1
#934130000000
0#
0(
#934140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#934190000000
0$
0)
#934200000000
1"
1'
b0 +
b0 1
#934250000000
0"
0'
#934260000000
1#
1(
b101111101100100 +
b101111101100100 1
#934310000000
0#
0(
#934320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#934370000000
0$
0)
#934380000000
1"
1'
b0 +
b0 1
#934430000000
0"
0'
#934440000000
1#
1(
b101111101100100 +
b101111101100100 1
#934490000000
0#
0(
#934500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#934550000000
0$
0)
#934560000000
1"
1'
b0 +
b0 1
#934610000000
0"
0'
#934620000000
1#
1(
b101111101100100 +
b101111101100100 1
#934670000000
0#
0(
#934680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#934730000000
0$
0)
#934740000000
1"
1'
b0 +
b0 1
#934790000000
0"
0'
#934800000000
1#
1(
b101111101100100 +
b101111101100100 1
#934850000000
0#
0(
#934860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#934910000000
0$
0)
#934920000000
1"
1'
b0 +
b0 1
#934970000000
0"
0'
#934980000000
1#
1(
b101111101100100 +
b101111101100100 1
#935030000000
0#
0(
#935040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#935090000000
0$
0)
#935100000000
1"
1'
b0 +
b0 1
#935150000000
0"
0'
#935160000000
1#
1(
b101111101100100 +
b101111101100100 1
#935210000000
0#
0(
#935220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#935270000000
0$
0)
#935280000000
1"
1'
b0 +
b0 1
#935330000000
0"
0'
#935340000000
1#
1(
b101111101100100 +
b101111101100100 1
#935390000000
0#
0(
#935400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#935450000000
0$
0)
#935460000000
1"
1'
b0 +
b0 1
#935510000000
0"
0'
#935520000000
1#
1(
b101111101100100 +
b101111101100100 1
#935570000000
0#
0(
#935580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#935630000000
0$
0)
#935640000000
1"
1'
b0 +
b0 1
#935690000000
0"
0'
#935700000000
1#
1(
b101111101100100 +
b101111101100100 1
#935750000000
0#
0(
#935760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#935810000000
0$
0)
#935820000000
1"
1'
b0 +
b0 1
#935870000000
0"
0'
#935880000000
1#
1(
b101111101100100 +
b101111101100100 1
#935930000000
0#
0(
#935940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#935990000000
0$
0)
#936000000000
1"
1'
b0 +
b0 1
#936050000000
0"
0'
#936060000000
1#
1(
b101111101100100 +
b101111101100100 1
#936110000000
0#
0(
#936120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#936170000000
0$
0)
#936180000000
1"
1'
b0 +
b0 1
#936230000000
0"
0'
#936240000000
1#
1(
b101111101100100 +
b101111101100100 1
#936290000000
0#
0(
#936300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#936350000000
0$
0)
#936360000000
1"
1'
b0 +
b0 1
#936410000000
0"
0'
#936420000000
1#
1(
b101111101100100 +
b101111101100100 1
#936470000000
0#
0(
#936480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#936530000000
0$
0)
#936540000000
1"
1'
b0 +
b0 1
#936590000000
0"
0'
#936600000000
1#
1(
b101111101100100 +
b101111101100100 1
#936650000000
0#
0(
#936660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#936710000000
0$
0)
#936720000000
1"
1'
b0 +
b0 1
#936770000000
0"
0'
#936780000000
1#
1(
b101111101100100 +
b101111101100100 1
#936830000000
0#
0(
#936840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#936890000000
0$
0)
#936900000000
1"
1'
b0 +
b0 1
#936950000000
0"
0'
#936960000000
1#
1(
b101111101100100 +
b101111101100100 1
#937010000000
0#
0(
#937020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#937070000000
0$
0)
#937080000000
1"
1'
b0 +
b0 1
#937130000000
0"
0'
#937140000000
1#
1(
b101111101100100 +
b101111101100100 1
#937190000000
0#
0(
#937200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#937250000000
0$
0)
#937260000000
1"
1'
b0 +
b0 1
#937310000000
0"
0'
#937320000000
1#
1(
b101111101100100 +
b101111101100100 1
#937370000000
0#
0(
#937380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#937430000000
0$
0)
#937440000000
1"
1'
b0 +
b0 1
#937490000000
0"
0'
#937500000000
1#
1(
b101111101100100 +
b101111101100100 1
#937550000000
0#
0(
#937560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#937610000000
0$
0)
#937620000000
1"
1'
b0 +
b0 1
#937670000000
0"
0'
#937680000000
1#
1(
b101111101100100 +
b101111101100100 1
#937730000000
0#
0(
#937740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#937790000000
0$
0)
#937800000000
1"
1'
b0 +
b0 1
#937850000000
0"
0'
#937860000000
1#
1(
b101111101100100 +
b101111101100100 1
#937910000000
0#
0(
#937920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#937970000000
0$
0)
#937980000000
1"
1'
b0 +
b0 1
#938030000000
0"
0'
#938040000000
1#
1(
b101111101100100 +
b101111101100100 1
#938090000000
0#
0(
#938100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#938150000000
0$
0)
#938160000000
1"
1'
b0 +
b0 1
#938210000000
0"
0'
#938220000000
1#
1(
b101111101100100 +
b101111101100100 1
#938270000000
0#
0(
#938280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#938330000000
0$
0)
#938340000000
1"
1'
b0 +
b0 1
#938390000000
0"
0'
#938400000000
1#
1(
b101111101100100 +
b101111101100100 1
#938450000000
0#
0(
#938460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#938510000000
0$
0)
#938520000000
1"
1'
b0 +
b0 1
#938570000000
0"
0'
#938580000000
1#
1(
b101111101100100 +
b101111101100100 1
#938630000000
0#
0(
#938640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#938690000000
0$
0)
#938700000000
1"
1'
b0 +
b0 1
#938750000000
0"
0'
#938760000000
1#
1(
b101111101100100 +
b101111101100100 1
#938810000000
0#
0(
#938820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#938870000000
0$
0)
#938880000000
1"
1'
b0 +
b0 1
#938930000000
0"
0'
#938940000000
1#
1(
b101111101100100 +
b101111101100100 1
#938990000000
0#
0(
#939000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#939050000000
0$
0)
#939060000000
1"
1'
b0 +
b0 1
#939110000000
0"
0'
#939120000000
1#
1(
b101111101100100 +
b101111101100100 1
#939170000000
0#
0(
#939180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#939230000000
0$
0)
#939240000000
1"
1'
b0 +
b0 1
#939290000000
0"
0'
#939300000000
1#
1(
b101111101100100 +
b101111101100100 1
#939350000000
0#
0(
#939360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#939410000000
0$
0)
#939420000000
1"
1'
b0 +
b0 1
#939470000000
0"
0'
#939480000000
1#
1(
b101111101100100 +
b101111101100100 1
#939530000000
0#
0(
#939540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#939590000000
0$
0)
#939600000000
1"
1'
b0 +
b0 1
#939650000000
0"
0'
#939660000000
1#
1(
b101111101100100 +
b101111101100100 1
#939710000000
0#
0(
#939720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#939770000000
0$
0)
#939780000000
1"
1'
b0 +
b0 1
#939830000000
0"
0'
#939840000000
1#
1(
b101111101100100 +
b101111101100100 1
#939890000000
0#
0(
#939900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#939950000000
0$
0)
#939960000000
1"
1'
b0 +
b0 1
#940010000000
0"
0'
#940020000000
1#
1(
b101111101100100 +
b101111101100100 1
#940070000000
0#
0(
#940080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#940130000000
0$
0)
#940140000000
1"
1'
b0 +
b0 1
#940190000000
0"
0'
#940200000000
1#
1(
b101111101100100 +
b101111101100100 1
#940250000000
0#
0(
#940260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#940310000000
0$
0)
#940320000000
1"
1'
b0 +
b0 1
#940370000000
0"
0'
#940380000000
1#
1(
b101111101100100 +
b101111101100100 1
#940430000000
0#
0(
#940440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#940490000000
0$
0)
#940500000000
1"
1'
b0 +
b0 1
#940550000000
0"
0'
#940560000000
1#
1(
b101111101100100 +
b101111101100100 1
#940610000000
0#
0(
#940620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#940670000000
0$
0)
#940680000000
1"
1'
b0 +
b0 1
#940730000000
0"
0'
#940740000000
1#
1(
b101111101100100 +
b101111101100100 1
#940790000000
0#
0(
#940800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#940850000000
0$
0)
#940860000000
1"
1'
b0 +
b0 1
#940910000000
0"
0'
#940920000000
1#
1(
b101111101100100 +
b101111101100100 1
#940970000000
0#
0(
#940980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#941030000000
0$
0)
#941040000000
1"
1'
b0 +
b0 1
#941090000000
0"
0'
#941100000000
1#
1(
b101111101100100 +
b101111101100100 1
#941150000000
0#
0(
#941160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#941210000000
0$
0)
#941220000000
1"
1'
b0 +
b0 1
#941270000000
0"
0'
#941280000000
1#
1(
b101111101100100 +
b101111101100100 1
#941330000000
0#
0(
#941340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#941390000000
0$
0)
#941400000000
1"
1'
b0 +
b0 1
#941450000000
0"
0'
#941460000000
1#
1(
b101111101100100 +
b101111101100100 1
#941510000000
0#
0(
#941520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#941570000000
0$
0)
#941580000000
1"
1'
b0 +
b0 1
#941630000000
0"
0'
#941640000000
1#
1(
b101111101100100 +
b101111101100100 1
#941690000000
0#
0(
#941700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#941750000000
0$
0)
#941760000000
1"
1'
b0 +
b0 1
#941810000000
0"
0'
#941820000000
1#
1(
b101111101100100 +
b101111101100100 1
#941870000000
0#
0(
#941880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#941930000000
0$
0)
#941940000000
1"
1'
b0 +
b0 1
#941990000000
0"
0'
#942000000000
1#
1(
b101111101100100 +
b101111101100100 1
#942050000000
0#
0(
#942060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#942110000000
0$
0)
#942120000000
1"
1'
b0 +
b0 1
#942170000000
0"
0'
#942180000000
1#
1(
b101111101100100 +
b101111101100100 1
#942230000000
0#
0(
#942240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#942290000000
0$
0)
#942300000000
1"
1'
b0 +
b0 1
#942350000000
0"
0'
#942360000000
1#
1(
b101111101100100 +
b101111101100100 1
#942410000000
0#
0(
#942420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#942470000000
0$
0)
#942480000000
1"
1'
b0 +
b0 1
#942530000000
0"
0'
#942540000000
1#
1(
b101111101100100 +
b101111101100100 1
#942590000000
0#
0(
#942600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#942650000000
0$
0)
#942660000000
1"
1'
b0 +
b0 1
#942710000000
0"
0'
#942720000000
1#
1(
b101111101100100 +
b101111101100100 1
#942770000000
0#
0(
#942780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#942830000000
0$
0)
#942840000000
1"
1'
b0 +
b0 1
#942890000000
0"
0'
#942900000000
1#
1(
b101111101100100 +
b101111101100100 1
#942950000000
0#
0(
#942960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#943010000000
0$
0)
#943020000000
1"
1'
b0 +
b0 1
#943070000000
0"
0'
#943080000000
1#
1(
b101111101100100 +
b101111101100100 1
#943130000000
0#
0(
#943140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#943190000000
0$
0)
#943200000000
1"
1'
b0 +
b0 1
#943250000000
0"
0'
#943260000000
1#
1(
b101111101100100 +
b101111101100100 1
#943310000000
0#
0(
#943320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#943370000000
0$
0)
#943380000000
1"
1'
b0 +
b0 1
#943430000000
0"
0'
#943440000000
1#
1(
b101111101100100 +
b101111101100100 1
#943490000000
0#
0(
#943500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#943550000000
0$
0)
#943560000000
1"
1'
b0 +
b0 1
#943610000000
0"
0'
#943620000000
1#
1(
b101111101100100 +
b101111101100100 1
#943670000000
0#
0(
#943680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#943730000000
0$
0)
#943740000000
1"
1'
b0 +
b0 1
#943790000000
0"
0'
#943800000000
1#
1(
b101111101100100 +
b101111101100100 1
#943850000000
0#
0(
#943860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#943910000000
0$
0)
#943920000000
1"
1'
b0 +
b0 1
#943970000000
0"
0'
#943980000000
1#
1(
b101111101100100 +
b101111101100100 1
#944030000000
0#
0(
#944040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#944090000000
0$
0)
#944100000000
1"
1'
b0 +
b0 1
#944150000000
0"
0'
#944160000000
1#
1(
b101111101100100 +
b101111101100100 1
#944210000000
0#
0(
#944220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#944270000000
0$
0)
#944280000000
1"
1'
b0 +
b0 1
#944330000000
0"
0'
#944340000000
1#
1(
b101111101100100 +
b101111101100100 1
#944390000000
0#
0(
#944400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#944450000000
0$
0)
#944460000000
1"
1'
b0 +
b0 1
#944510000000
0"
0'
#944520000000
1#
1(
b101111101100100 +
b101111101100100 1
#944570000000
0#
0(
#944580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#944630000000
0$
0)
#944640000000
1"
1'
b0 +
b0 1
#944690000000
0"
0'
#944700000000
1#
1(
b101111101100100 +
b101111101100100 1
#944750000000
0#
0(
#944760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#944810000000
0$
0)
#944820000000
1"
1'
b0 +
b0 1
#944870000000
0"
0'
#944880000000
1#
1(
b101111101100100 +
b101111101100100 1
#944930000000
0#
0(
#944940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#944990000000
0$
0)
#945000000000
1"
1'
b0 +
b0 1
#945050000000
0"
0'
#945060000000
1#
1(
b101111101100100 +
b101111101100100 1
#945110000000
0#
0(
#945120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#945170000000
0$
0)
#945180000000
1"
1'
b0 +
b0 1
#945230000000
0"
0'
#945240000000
1#
1(
b101111101100100 +
b101111101100100 1
#945290000000
0#
0(
#945300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#945350000000
0$
0)
#945360000000
1"
1'
b0 +
b0 1
#945410000000
0"
0'
#945420000000
1#
1(
b101111101100100 +
b101111101100100 1
#945470000000
0#
0(
#945480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#945530000000
0$
0)
#945540000000
1"
1'
b0 +
b0 1
#945590000000
0"
0'
#945600000000
1#
1(
b101111101100100 +
b101111101100100 1
#945650000000
0#
0(
#945660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#945710000000
0$
0)
#945720000000
1"
1'
b0 +
b0 1
#945770000000
0"
0'
#945780000000
1#
1(
b101111101100100 +
b101111101100100 1
#945830000000
0#
0(
#945840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#945890000000
0$
0)
#945900000000
1"
1'
b0 +
b0 1
#945950000000
0"
0'
#945960000000
1#
1(
b101111101100100 +
b101111101100100 1
#946010000000
0#
0(
#946020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#946070000000
0$
0)
#946080000000
1"
1'
b0 +
b0 1
#946130000000
0"
0'
#946140000000
1#
1(
b101111101100100 +
b101111101100100 1
#946190000000
0#
0(
#946200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#946250000000
0$
0)
#946260000000
1"
1'
b0 +
b0 1
#946310000000
0"
0'
#946320000000
1#
1(
b101111101100100 +
b101111101100100 1
#946370000000
0#
0(
#946380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#946430000000
0$
0)
#946440000000
1"
1'
b0 +
b0 1
#946490000000
0"
0'
#946500000000
1#
1(
b101111101100100 +
b101111101100100 1
#946550000000
0#
0(
#946560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#946610000000
0$
0)
#946620000000
1"
1'
b0 +
b0 1
#946670000000
0"
0'
#946680000000
1#
1(
b101111101100100 +
b101111101100100 1
#946730000000
0#
0(
#946740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#946790000000
0$
0)
#946800000000
1"
1'
b0 +
b0 1
#946850000000
0"
0'
#946860000000
1#
1(
b101111101100100 +
b101111101100100 1
#946910000000
0#
0(
#946920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#946970000000
0$
0)
#946980000000
1"
1'
b0 +
b0 1
#947030000000
0"
0'
#947040000000
1#
1(
b101111101100100 +
b101111101100100 1
#947090000000
0#
0(
#947100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#947150000000
0$
0)
#947160000000
1"
1'
b0 +
b0 1
#947210000000
0"
0'
#947220000000
1#
1(
b101111101100100 +
b101111101100100 1
#947270000000
0#
0(
#947280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#947330000000
0$
0)
#947340000000
1"
1'
b0 +
b0 1
#947390000000
0"
0'
#947400000000
1#
1(
b101111101100100 +
b101111101100100 1
#947450000000
0#
0(
#947460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#947510000000
0$
0)
#947520000000
1"
1'
b0 +
b0 1
#947570000000
0"
0'
#947580000000
1#
1(
b101111101100100 +
b101111101100100 1
#947630000000
0#
0(
#947640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#947690000000
0$
0)
#947700000000
1"
1'
b0 +
b0 1
#947750000000
0"
0'
#947760000000
1#
1(
b101111101100100 +
b101111101100100 1
#947810000000
0#
0(
#947820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#947870000000
0$
0)
#947880000000
1"
1'
b0 +
b0 1
#947930000000
0"
0'
#947940000000
1#
1(
b101111101100100 +
b101111101100100 1
#947990000000
0#
0(
#948000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#948050000000
0$
0)
#948060000000
1"
1'
b0 +
b0 1
#948110000000
0"
0'
#948120000000
1#
1(
b101111101100100 +
b101111101100100 1
#948170000000
0#
0(
#948180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#948230000000
0$
0)
#948240000000
1"
1'
b0 +
b0 1
#948290000000
0"
0'
#948300000000
1#
1(
b101111101100100 +
b101111101100100 1
#948350000000
0#
0(
#948360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#948410000000
0$
0)
#948420000000
1"
1'
b0 +
b0 1
#948470000000
0"
0'
#948480000000
1#
1(
b101111101100100 +
b101111101100100 1
#948530000000
0#
0(
#948540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#948590000000
0$
0)
#948600000000
1"
1'
b0 +
b0 1
#948650000000
0"
0'
#948660000000
1#
1(
b101111101100100 +
b101111101100100 1
#948710000000
0#
0(
#948720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#948770000000
0$
0)
#948780000000
1"
1'
b0 +
b0 1
#948830000000
0"
0'
#948840000000
1#
1(
b101111101100100 +
b101111101100100 1
#948890000000
0#
0(
#948900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#948950000000
0$
0)
#948960000000
1"
1'
b0 +
b0 1
#949010000000
0"
0'
#949020000000
1#
1(
b101111101100100 +
b101111101100100 1
#949070000000
0#
0(
#949080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#949130000000
0$
0)
#949140000000
1"
1'
b0 +
b0 1
#949190000000
0"
0'
#949200000000
1#
1(
b101111101100100 +
b101111101100100 1
#949250000000
0#
0(
#949260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#949310000000
0$
0)
#949320000000
1"
1'
b0 +
b0 1
#949370000000
0"
0'
#949380000000
1#
1(
b101111101100100 +
b101111101100100 1
#949430000000
0#
0(
#949440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#949490000000
0$
0)
#949500000000
1"
1'
b0 +
b0 1
#949550000000
0"
0'
#949560000000
1#
1(
b101111101100100 +
b101111101100100 1
#949610000000
0#
0(
#949620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#949670000000
0$
0)
#949680000000
1"
1'
b0 +
b0 1
#949730000000
0"
0'
#949740000000
1#
1(
b101111101100100 +
b101111101100100 1
#949790000000
0#
0(
#949800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#949850000000
0$
0)
#949860000000
1"
1'
b0 +
b0 1
#949910000000
0"
0'
#949920000000
1#
1(
b101111101100100 +
b101111101100100 1
#949970000000
0#
0(
#949980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#950030000000
0$
0)
#950040000000
1"
1'
b0 +
b0 1
#950090000000
0"
0'
#950100000000
1#
1(
b101111101100100 +
b101111101100100 1
#950150000000
0#
0(
#950160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#950210000000
0$
0)
#950220000000
1"
1'
b0 +
b0 1
#950270000000
0"
0'
#950280000000
1#
1(
b101111101100100 +
b101111101100100 1
#950330000000
0#
0(
#950340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#950390000000
0$
0)
#950400000000
1"
1'
b0 +
b0 1
#950450000000
0"
0'
#950460000000
1#
1(
b101111101100100 +
b101111101100100 1
#950510000000
0#
0(
#950520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#950570000000
0$
0)
#950580000000
1"
1'
b0 +
b0 1
#950630000000
0"
0'
#950640000000
1#
1(
b101111101100100 +
b101111101100100 1
#950690000000
0#
0(
#950700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#950750000000
0$
0)
#950760000000
1"
1'
b0 +
b0 1
#950810000000
0"
0'
#950820000000
1#
1(
b101111101100100 +
b101111101100100 1
#950870000000
0#
0(
#950880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#950930000000
0$
0)
#950940000000
1"
1'
b0 +
b0 1
#950990000000
0"
0'
#951000000000
1#
1(
b101111101100100 +
b101111101100100 1
#951050000000
0#
0(
#951060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#951110000000
0$
0)
#951120000000
1"
1'
b0 +
b0 1
#951170000000
0"
0'
#951180000000
1#
1(
b101111101100100 +
b101111101100100 1
#951230000000
0#
0(
#951240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#951290000000
0$
0)
#951300000000
1"
1'
b0 +
b0 1
#951350000000
0"
0'
#951360000000
1#
1(
b101111101100100 +
b101111101100100 1
#951410000000
0#
0(
#951420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#951470000000
0$
0)
#951480000000
1"
1'
b0 +
b0 1
#951530000000
0"
0'
#951540000000
1#
1(
b101111101100100 +
b101111101100100 1
#951590000000
0#
0(
#951600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#951650000000
0$
0)
#951660000000
1"
1'
b0 +
b0 1
#951710000000
0"
0'
#951720000000
1#
1(
b101111101100100 +
b101111101100100 1
#951770000000
0#
0(
#951780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#951830000000
0$
0)
#951840000000
1"
1'
b0 +
b0 1
#951890000000
0"
0'
#951900000000
1#
1(
b101111101100100 +
b101111101100100 1
#951950000000
0#
0(
#951960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#952010000000
0$
0)
#952020000000
1"
1'
b0 +
b0 1
#952070000000
0"
0'
#952080000000
1#
1(
b101111101100100 +
b101111101100100 1
#952130000000
0#
0(
#952140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#952190000000
0$
0)
#952200000000
1"
1'
b0 +
b0 1
#952250000000
0"
0'
#952260000000
1#
1(
b101111101100100 +
b101111101100100 1
#952310000000
0#
0(
#952320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#952370000000
0$
0)
#952380000000
1"
1'
b0 +
b0 1
#952430000000
0"
0'
#952440000000
1#
1(
b101111101100100 +
b101111101100100 1
#952490000000
0#
0(
#952500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#952550000000
0$
0)
#952560000000
1"
1'
b0 +
b0 1
#952610000000
0"
0'
#952620000000
1#
1(
b101111101100100 +
b101111101100100 1
#952670000000
0#
0(
#952680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#952730000000
0$
0)
#952740000000
1"
1'
b0 +
b0 1
#952790000000
0"
0'
#952800000000
1#
1(
b101111101100100 +
b101111101100100 1
#952850000000
0#
0(
#952860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#952910000000
0$
0)
#952920000000
1"
1'
b0 +
b0 1
#952970000000
0"
0'
#952980000000
1#
1(
b101111101100100 +
b101111101100100 1
#953030000000
0#
0(
#953040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#953090000000
0$
0)
#953100000000
1"
1'
b0 +
b0 1
#953150000000
0"
0'
#953160000000
1#
1(
b101111101100100 +
b101111101100100 1
#953210000000
0#
0(
#953220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#953270000000
0$
0)
#953280000000
1"
1'
b0 +
b0 1
#953330000000
0"
0'
#953340000000
1#
1(
b101111101100100 +
b101111101100100 1
#953390000000
0#
0(
#953400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#953450000000
0$
0)
#953460000000
1"
1'
b0 +
b0 1
#953510000000
0"
0'
#953520000000
1#
1(
b101111101100100 +
b101111101100100 1
#953570000000
0#
0(
#953580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#953630000000
0$
0)
#953640000000
1"
1'
b0 +
b0 1
#953690000000
0"
0'
#953700000000
1#
1(
b101111101100100 +
b101111101100100 1
#953750000000
0#
0(
#953760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#953810000000
0$
0)
#953820000000
1"
1'
b0 +
b0 1
#953870000000
0"
0'
#953880000000
1#
1(
b101111101100100 +
b101111101100100 1
#953930000000
0#
0(
#953940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#953990000000
0$
0)
#954000000000
1"
1'
b0 +
b0 1
#954050000000
0"
0'
#954060000000
1#
1(
b101111101100100 +
b101111101100100 1
#954110000000
0#
0(
#954120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#954170000000
0$
0)
#954180000000
1"
1'
b0 +
b0 1
#954230000000
0"
0'
#954240000000
1#
1(
b101111101100100 +
b101111101100100 1
#954290000000
0#
0(
#954300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#954350000000
0$
0)
#954360000000
1"
1'
b0 +
b0 1
#954410000000
0"
0'
#954420000000
1#
1(
b101111101100100 +
b101111101100100 1
#954470000000
0#
0(
#954480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#954530000000
0$
0)
#954540000000
1"
1'
b0 +
b0 1
#954590000000
0"
0'
#954600000000
1#
1(
b101111101100100 +
b101111101100100 1
#954650000000
0#
0(
#954660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#954710000000
0$
0)
#954720000000
1"
1'
b0 +
b0 1
#954770000000
0"
0'
#954780000000
1#
1(
b101111101100100 +
b101111101100100 1
#954830000000
0#
0(
#954840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#954890000000
0$
0)
#954900000000
1"
1'
b0 +
b0 1
#954950000000
0"
0'
#954960000000
1#
1(
b101111101100100 +
b101111101100100 1
#955010000000
0#
0(
#955020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#955070000000
0$
0)
#955080000000
1"
1'
b0 +
b0 1
#955130000000
0"
0'
#955140000000
1#
1(
b101111101100100 +
b101111101100100 1
#955190000000
0#
0(
#955200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#955250000000
0$
0)
#955260000000
1"
1'
b0 +
b0 1
#955310000000
0"
0'
#955320000000
1#
1(
b101111101100100 +
b101111101100100 1
#955370000000
0#
0(
#955380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#955430000000
0$
0)
#955440000000
1"
1'
b0 +
b0 1
#955490000000
0"
0'
#955500000000
1#
1(
b101111101100100 +
b101111101100100 1
#955550000000
0#
0(
#955560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#955610000000
0$
0)
#955620000000
1"
1'
b0 +
b0 1
#955670000000
0"
0'
#955680000000
1#
1(
b101111101100100 +
b101111101100100 1
#955730000000
0#
0(
#955740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#955790000000
0$
0)
#955800000000
1"
1'
b0 +
b0 1
#955850000000
0"
0'
#955860000000
1#
1(
b101111101100100 +
b101111101100100 1
#955910000000
0#
0(
#955920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#955970000000
0$
0)
#955980000000
1"
1'
b0 +
b0 1
#956030000000
0"
0'
#956040000000
1#
1(
b101111101100100 +
b101111101100100 1
#956090000000
0#
0(
#956100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#956150000000
0$
0)
#956160000000
1"
1'
b0 +
b0 1
#956210000000
0"
0'
#956220000000
1#
1(
b101111101100100 +
b101111101100100 1
#956270000000
0#
0(
#956280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#956330000000
0$
0)
#956340000000
1"
1'
b0 +
b0 1
#956390000000
0"
0'
#956400000000
1#
1(
b101111101100100 +
b101111101100100 1
#956450000000
0#
0(
#956460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#956510000000
0$
0)
#956520000000
1"
1'
b0 +
b0 1
#956570000000
0"
0'
#956580000000
1#
1(
b101111101100100 +
b101111101100100 1
#956630000000
0#
0(
#956640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#956690000000
0$
0)
#956700000000
1"
1'
b0 +
b0 1
#956750000000
0"
0'
#956760000000
1#
1(
b101111101100100 +
b101111101100100 1
#956810000000
0#
0(
#956820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#956870000000
0$
0)
#956880000000
1"
1'
b0 +
b0 1
#956930000000
0"
0'
#956940000000
1#
1(
b101111101100100 +
b101111101100100 1
#956990000000
0#
0(
#957000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#957050000000
0$
0)
#957060000000
1"
1'
b0 +
b0 1
#957110000000
0"
0'
#957120000000
1#
1(
b101111101100100 +
b101111101100100 1
#957170000000
0#
0(
#957180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#957230000000
0$
0)
#957240000000
1"
1'
b0 +
b0 1
#957290000000
0"
0'
#957300000000
1#
1(
b101111101100100 +
b101111101100100 1
#957350000000
0#
0(
#957360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#957410000000
0$
0)
#957420000000
1"
1'
b0 +
b0 1
#957470000000
0"
0'
#957480000000
1#
1(
b101111101100100 +
b101111101100100 1
#957530000000
0#
0(
#957540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#957590000000
0$
0)
#957600000000
1"
1'
b0 +
b0 1
#957650000000
0"
0'
#957660000000
1#
1(
b101111101100100 +
b101111101100100 1
#957710000000
0#
0(
#957720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#957770000000
0$
0)
#957780000000
1"
1'
b0 +
b0 1
#957830000000
0"
0'
#957840000000
1#
1(
b101111101100100 +
b101111101100100 1
#957890000000
0#
0(
#957900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#957950000000
0$
0)
#957960000000
1"
1'
b0 +
b0 1
#958010000000
0"
0'
#958020000000
1#
1(
b101111101100100 +
b101111101100100 1
#958070000000
0#
0(
#958080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#958130000000
0$
0)
#958140000000
1"
1'
b0 +
b0 1
#958190000000
0"
0'
#958200000000
1#
1(
b101111101100100 +
b101111101100100 1
#958250000000
0#
0(
#958260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#958310000000
0$
0)
#958320000000
1"
1'
b0 +
b0 1
#958370000000
0"
0'
#958380000000
1#
1(
b101111101100100 +
b101111101100100 1
#958430000000
0#
0(
#958440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#958490000000
0$
0)
#958500000000
1"
1'
b0 +
b0 1
#958550000000
0"
0'
#958560000000
1#
1(
b101111101100100 +
b101111101100100 1
#958610000000
0#
0(
#958620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#958670000000
0$
0)
#958680000000
1"
1'
b0 +
b0 1
#958730000000
0"
0'
#958740000000
1#
1(
b101111101100100 +
b101111101100100 1
#958790000000
0#
0(
#958800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#958850000000
0$
0)
#958860000000
1"
1'
b0 +
b0 1
#958910000000
0"
0'
#958920000000
1#
1(
b101111101100100 +
b101111101100100 1
#958970000000
0#
0(
#958980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#959030000000
0$
0)
#959040000000
1"
1'
b0 +
b0 1
#959090000000
0"
0'
#959100000000
1#
1(
b101111101100100 +
b101111101100100 1
#959150000000
0#
0(
#959160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#959210000000
0$
0)
#959220000000
1"
1'
b0 +
b0 1
#959270000000
0"
0'
#959280000000
1#
1(
b101111101100100 +
b101111101100100 1
#959330000000
0#
0(
#959340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#959390000000
0$
0)
#959400000000
1"
1'
b0 +
b0 1
#959450000000
0"
0'
#959460000000
1#
1(
b101111101100100 +
b101111101100100 1
#959510000000
0#
0(
#959520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#959570000000
0$
0)
#959580000000
1"
1'
b0 +
b0 1
#959630000000
0"
0'
#959640000000
1#
1(
b101111101100100 +
b101111101100100 1
#959690000000
0#
0(
#959700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#959750000000
0$
0)
#959760000000
1"
1'
b0 +
b0 1
#959810000000
0"
0'
#959820000000
1#
1(
b101111101100100 +
b101111101100100 1
#959870000000
0#
0(
#959880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#959930000000
0$
0)
#959940000000
1"
1'
b0 +
b0 1
#959990000000
0"
0'
#960000000000
1#
1(
b101111101100100 +
b101111101100100 1
#960050000000
0#
0(
#960060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#960110000000
0$
0)
#960120000000
1"
1'
b0 +
b0 1
#960170000000
0"
0'
#960180000000
1#
1(
b101111101100100 +
b101111101100100 1
#960230000000
0#
0(
#960240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#960290000000
0$
0)
#960300000000
1"
1'
b0 +
b0 1
#960350000000
0"
0'
#960360000000
1#
1(
b101111101100100 +
b101111101100100 1
#960410000000
0#
0(
#960420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#960470000000
0$
0)
#960480000000
1"
1'
b0 +
b0 1
#960530000000
0"
0'
#960540000000
1#
1(
b101111101100100 +
b101111101100100 1
#960590000000
0#
0(
#960600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#960650000000
0$
0)
#960660000000
1"
1'
b0 +
b0 1
#960710000000
0"
0'
#960720000000
1#
1(
b101111101100100 +
b101111101100100 1
#960770000000
0#
0(
#960780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#960830000000
0$
0)
#960840000000
1"
1'
b0 +
b0 1
#960890000000
0"
0'
#960900000000
1#
1(
b101111101100100 +
b101111101100100 1
#960950000000
0#
0(
#960960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#961010000000
0$
0)
#961020000000
1"
1'
b0 +
b0 1
#961070000000
0"
0'
#961080000000
1#
1(
b101111101100100 +
b101111101100100 1
#961130000000
0#
0(
#961140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#961190000000
0$
0)
#961200000000
1"
1'
b0 +
b0 1
#961250000000
0"
0'
#961260000000
1#
1(
b101111101100100 +
b101111101100100 1
#961310000000
0#
0(
#961320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#961370000000
0$
0)
#961380000000
1"
1'
b0 +
b0 1
#961430000000
0"
0'
#961440000000
1#
1(
b101111101100100 +
b101111101100100 1
#961490000000
0#
0(
#961500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#961550000000
0$
0)
#961560000000
1"
1'
b0 +
b0 1
#961610000000
0"
0'
#961620000000
1#
1(
b101111101100100 +
b101111101100100 1
#961670000000
0#
0(
#961680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#961730000000
0$
0)
#961740000000
1"
1'
b0 +
b0 1
#961790000000
0"
0'
#961800000000
1#
1(
b101111101100100 +
b101111101100100 1
#961850000000
0#
0(
#961860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#961910000000
0$
0)
#961920000000
1"
1'
b0 +
b0 1
#961970000000
0"
0'
#961980000000
1#
1(
b101111101100100 +
b101111101100100 1
#962030000000
0#
0(
#962040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#962090000000
0$
0)
#962100000000
1"
1'
b0 +
b0 1
#962150000000
0"
0'
#962160000000
1#
1(
b101111101100100 +
b101111101100100 1
#962210000000
0#
0(
#962220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#962270000000
0$
0)
#962280000000
1"
1'
b0 +
b0 1
#962330000000
0"
0'
#962340000000
1#
1(
b101111101100100 +
b101111101100100 1
#962390000000
0#
0(
#962400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#962450000000
0$
0)
#962460000000
1"
1'
b0 +
b0 1
#962510000000
0"
0'
#962520000000
1#
1(
b101111101100100 +
b101111101100100 1
#962570000000
0#
0(
#962580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#962630000000
0$
0)
#962640000000
1"
1'
b0 +
b0 1
#962690000000
0"
0'
#962700000000
1#
1(
b101111101100100 +
b101111101100100 1
#962750000000
0#
0(
#962760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#962810000000
0$
0)
#962820000000
1"
1'
b0 +
b0 1
#962870000000
0"
0'
#962880000000
1#
1(
b101111101100100 +
b101111101100100 1
#962930000000
0#
0(
#962940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#962990000000
0$
0)
#963000000000
1"
1'
b0 +
b0 1
#963050000000
0"
0'
#963060000000
1#
1(
b101111101100100 +
b101111101100100 1
#963110000000
0#
0(
#963120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#963170000000
0$
0)
#963180000000
1"
1'
b0 +
b0 1
#963230000000
0"
0'
#963240000000
1#
1(
b101111101100100 +
b101111101100100 1
#963290000000
0#
0(
#963300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#963350000000
0$
0)
#963360000000
1"
1'
b0 +
b0 1
#963410000000
0"
0'
#963420000000
1#
1(
b101111101100100 +
b101111101100100 1
#963470000000
0#
0(
#963480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#963530000000
0$
0)
#963540000000
1"
1'
b0 +
b0 1
#963590000000
0"
0'
#963600000000
1#
1(
b101111101100100 +
b101111101100100 1
#963650000000
0#
0(
#963660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#963710000000
0$
0)
#963720000000
1"
1'
b0 +
b0 1
#963770000000
0"
0'
#963780000000
1#
1(
b101111101100100 +
b101111101100100 1
#963830000000
0#
0(
#963840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#963890000000
0$
0)
#963900000000
1"
1'
b0 +
b0 1
#963950000000
0"
0'
#963960000000
1#
1(
b101111101100100 +
b101111101100100 1
#964010000000
0#
0(
#964020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#964070000000
0$
0)
#964080000000
1"
1'
b0 +
b0 1
#964130000000
0"
0'
#964140000000
1#
1(
b101111101100100 +
b101111101100100 1
#964190000000
0#
0(
#964200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#964250000000
0$
0)
#964260000000
1"
1'
b0 +
b0 1
#964310000000
0"
0'
#964320000000
1#
1(
b101111101100100 +
b101111101100100 1
#964370000000
0#
0(
#964380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#964430000000
0$
0)
#964440000000
1"
1'
b0 +
b0 1
#964490000000
0"
0'
#964500000000
1#
1(
b101111101100100 +
b101111101100100 1
#964550000000
0#
0(
#964560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#964610000000
0$
0)
#964620000000
1"
1'
b0 +
b0 1
#964670000000
0"
0'
#964680000000
1#
1(
b101111101100100 +
b101111101100100 1
#964730000000
0#
0(
#964740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#964790000000
0$
0)
#964800000000
1"
1'
b0 +
b0 1
#964850000000
0"
0'
#964860000000
1#
1(
b101111101100100 +
b101111101100100 1
#964910000000
0#
0(
#964920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#964970000000
0$
0)
#964980000000
1"
1'
b0 +
b0 1
#965030000000
0"
0'
#965040000000
1#
1(
b101111101100100 +
b101111101100100 1
#965090000000
0#
0(
#965100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#965150000000
0$
0)
#965160000000
1"
1'
b0 +
b0 1
#965210000000
0"
0'
#965220000000
1#
1(
b101111101100100 +
b101111101100100 1
#965270000000
0#
0(
#965280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#965330000000
0$
0)
#965340000000
1"
1'
b0 +
b0 1
#965390000000
0"
0'
#965400000000
1#
1(
b101111101100100 +
b101111101100100 1
#965450000000
0#
0(
#965460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#965510000000
0$
0)
#965520000000
1"
1'
b0 +
b0 1
#965570000000
0"
0'
#965580000000
1#
1(
b101111101100100 +
b101111101100100 1
#965630000000
0#
0(
#965640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#965690000000
0$
0)
#965700000000
1"
1'
b0 +
b0 1
#965750000000
0"
0'
#965760000000
1#
1(
b101111101100100 +
b101111101100100 1
#965810000000
0#
0(
#965820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#965870000000
0$
0)
#965880000000
1"
1'
b0 +
b0 1
#965930000000
0"
0'
#965940000000
1#
1(
b101111101100100 +
b101111101100100 1
#965990000000
0#
0(
#966000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#966050000000
0$
0)
#966060000000
1"
1'
b0 +
b0 1
#966110000000
0"
0'
#966120000000
1#
1(
b101111101100100 +
b101111101100100 1
#966170000000
0#
0(
#966180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#966230000000
0$
0)
#966240000000
1"
1'
b0 +
b0 1
#966290000000
0"
0'
#966300000000
1#
1(
b101111101100100 +
b101111101100100 1
#966350000000
0#
0(
#966360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#966410000000
0$
0)
#966420000000
1"
1'
b0 +
b0 1
#966470000000
0"
0'
#966480000000
1#
1(
b101111101100100 +
b101111101100100 1
#966530000000
0#
0(
#966540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#966590000000
0$
0)
#966600000000
1"
1'
b0 +
b0 1
#966650000000
0"
0'
#966660000000
1#
1(
b101111101100100 +
b101111101100100 1
#966710000000
0#
0(
#966720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#966770000000
0$
0)
#966780000000
1"
1'
b0 +
b0 1
#966830000000
0"
0'
#966840000000
1#
1(
b101111101100100 +
b101111101100100 1
#966890000000
0#
0(
#966900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#966950000000
0$
0)
#966960000000
1"
1'
b0 +
b0 1
#967010000000
0"
0'
#967020000000
1#
1(
b101111101100100 +
b101111101100100 1
#967070000000
0#
0(
#967080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#967130000000
0$
0)
#967140000000
1"
1'
b0 +
b0 1
#967190000000
0"
0'
#967200000000
1#
1(
b101111101100100 +
b101111101100100 1
#967250000000
0#
0(
#967260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#967310000000
0$
0)
#967320000000
1"
1'
b0 +
b0 1
#967370000000
0"
0'
#967380000000
1#
1(
b101111101100100 +
b101111101100100 1
#967430000000
0#
0(
#967440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#967490000000
0$
0)
#967500000000
1"
1'
b0 +
b0 1
#967550000000
0"
0'
#967560000000
1#
1(
b101111101100100 +
b101111101100100 1
#967610000000
0#
0(
#967620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#967670000000
0$
0)
#967680000000
1"
1'
b0 +
b0 1
#967730000000
0"
0'
#967740000000
1#
1(
b101111101100100 +
b101111101100100 1
#967790000000
0#
0(
#967800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#967850000000
0$
0)
#967860000000
1"
1'
b0 +
b0 1
#967910000000
0"
0'
#967920000000
1#
1(
b101111101100100 +
b101111101100100 1
#967970000000
0#
0(
#967980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#968030000000
0$
0)
#968040000000
1"
1'
b0 +
b0 1
#968090000000
0"
0'
#968100000000
1#
1(
b101111101100100 +
b101111101100100 1
#968150000000
0#
0(
#968160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#968210000000
0$
0)
#968220000000
1"
1'
b0 +
b0 1
#968270000000
0"
0'
#968280000000
1#
1(
b101111101100100 +
b101111101100100 1
#968330000000
0#
0(
#968340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#968390000000
0$
0)
#968400000000
1"
1'
b0 +
b0 1
#968450000000
0"
0'
#968460000000
1#
1(
b101111101100100 +
b101111101100100 1
#968510000000
0#
0(
#968520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#968570000000
0$
0)
#968580000000
1"
1'
b0 +
b0 1
#968630000000
0"
0'
#968640000000
1#
1(
b101111101100100 +
b101111101100100 1
#968690000000
0#
0(
#968700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#968750000000
0$
0)
#968760000000
1"
1'
b0 +
b0 1
#968810000000
0"
0'
#968820000000
1#
1(
b101111101100100 +
b101111101100100 1
#968870000000
0#
0(
#968880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#968930000000
0$
0)
#968940000000
1"
1'
b0 +
b0 1
#968990000000
0"
0'
#969000000000
1#
1(
b101111101100100 +
b101111101100100 1
#969050000000
0#
0(
#969060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#969110000000
0$
0)
#969120000000
1"
1'
b0 +
b0 1
#969170000000
0"
0'
#969180000000
1#
1(
b101111101100100 +
b101111101100100 1
#969230000000
0#
0(
#969240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#969290000000
0$
0)
#969300000000
1"
1'
b0 +
b0 1
#969350000000
0"
0'
#969360000000
1#
1(
b101111101100100 +
b101111101100100 1
#969410000000
0#
0(
#969420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#969470000000
0$
0)
#969480000000
1"
1'
b0 +
b0 1
#969530000000
0"
0'
#969540000000
1#
1(
b101111101100100 +
b101111101100100 1
#969590000000
0#
0(
#969600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#969650000000
0$
0)
#969660000000
1"
1'
b0 +
b0 1
#969710000000
0"
0'
#969720000000
1#
1(
b101111101100100 +
b101111101100100 1
#969770000000
0#
0(
#969780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#969830000000
0$
0)
#969840000000
1"
1'
b0 +
b0 1
#969890000000
0"
0'
#969900000000
1#
1(
b101111101100100 +
b101111101100100 1
#969950000000
0#
0(
#969960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#970010000000
0$
0)
#970020000000
1"
1'
b0 +
b0 1
#970070000000
0"
0'
#970080000000
1#
1(
b101111101100100 +
b101111101100100 1
#970130000000
0#
0(
#970140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#970190000000
0$
0)
#970200000000
1"
1'
b0 +
b0 1
#970250000000
0"
0'
#970260000000
1#
1(
b101111101100100 +
b101111101100100 1
#970310000000
0#
0(
#970320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#970370000000
0$
0)
#970380000000
1"
1'
b0 +
b0 1
#970430000000
0"
0'
#970440000000
1#
1(
b101111101100100 +
b101111101100100 1
#970490000000
0#
0(
#970500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#970550000000
0$
0)
#970560000000
1"
1'
b0 +
b0 1
#970610000000
0"
0'
#970620000000
1#
1(
b101111101100100 +
b101111101100100 1
#970670000000
0#
0(
#970680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#970730000000
0$
0)
#970740000000
1"
1'
b0 +
b0 1
#970790000000
0"
0'
#970800000000
1#
1(
b101111101100100 +
b101111101100100 1
#970850000000
0#
0(
#970860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#970910000000
0$
0)
#970920000000
1"
1'
b0 +
b0 1
#970970000000
0"
0'
#970980000000
1#
1(
b101111101100100 +
b101111101100100 1
#971030000000
0#
0(
#971040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#971090000000
0$
0)
#971100000000
1"
1'
b0 +
b0 1
#971150000000
0"
0'
#971160000000
1#
1(
b101111101100100 +
b101111101100100 1
#971210000000
0#
0(
#971220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#971270000000
0$
0)
#971280000000
1"
1'
b0 +
b0 1
#971330000000
0"
0'
#971340000000
1#
1(
b101111101100100 +
b101111101100100 1
#971390000000
0#
0(
#971400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#971450000000
0$
0)
#971460000000
1"
1'
b0 +
b0 1
#971510000000
0"
0'
#971520000000
1#
1(
b101111101100100 +
b101111101100100 1
#971570000000
0#
0(
#971580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#971630000000
0$
0)
#971640000000
1"
1'
b0 +
b0 1
#971690000000
0"
0'
#971700000000
1#
1(
b101111101100100 +
b101111101100100 1
#971750000000
0#
0(
#971760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#971810000000
0$
0)
#971820000000
1"
1'
b0 +
b0 1
#971870000000
0"
0'
#971880000000
1#
1(
b101111101100100 +
b101111101100100 1
#971930000000
0#
0(
#971940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#971990000000
0$
0)
#972000000000
1"
1'
b0 +
b0 1
#972050000000
0"
0'
#972060000000
1#
1(
b101111101100100 +
b101111101100100 1
#972110000000
0#
0(
#972120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#972170000000
0$
0)
#972180000000
1"
1'
b0 +
b0 1
#972230000000
0"
0'
#972240000000
1#
1(
b101111101100100 +
b101111101100100 1
#972290000000
0#
0(
#972300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#972350000000
0$
0)
#972360000000
1"
1'
b0 +
b0 1
#972410000000
0"
0'
#972420000000
1#
1(
b101111101100100 +
b101111101100100 1
#972470000000
0#
0(
#972480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#972530000000
0$
0)
#972540000000
1"
1'
b0 +
b0 1
#972590000000
0"
0'
#972600000000
1#
1(
b101111101100100 +
b101111101100100 1
#972650000000
0#
0(
#972660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#972710000000
0$
0)
#972720000000
1"
1'
b0 +
b0 1
#972770000000
0"
0'
#972780000000
1#
1(
b101111101100100 +
b101111101100100 1
#972830000000
0#
0(
#972840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#972890000000
0$
0)
#972900000000
1"
1'
b0 +
b0 1
#972950000000
0"
0'
#972960000000
1#
1(
b101111101100100 +
b101111101100100 1
#973010000000
0#
0(
#973020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#973070000000
0$
0)
#973080000000
1"
1'
b0 +
b0 1
#973130000000
0"
0'
#973140000000
1#
1(
b101111101100100 +
b101111101100100 1
#973190000000
0#
0(
#973200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#973250000000
0$
0)
#973260000000
1"
1'
b0 +
b0 1
#973310000000
0"
0'
#973320000000
1#
1(
b101111101100100 +
b101111101100100 1
#973370000000
0#
0(
#973380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#973430000000
0$
0)
#973440000000
1"
1'
b0 +
b0 1
#973490000000
0"
0'
#973500000000
1#
1(
b101111101100100 +
b101111101100100 1
#973550000000
0#
0(
#973560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#973610000000
0$
0)
#973620000000
1"
1'
b0 +
b0 1
#973670000000
0"
0'
#973680000000
1#
1(
b101111101100100 +
b101111101100100 1
#973730000000
0#
0(
#973740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#973790000000
0$
0)
#973800000000
1"
1'
b0 +
b0 1
#973850000000
0"
0'
#973860000000
1#
1(
b101111101100100 +
b101111101100100 1
#973910000000
0#
0(
#973920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#973970000000
0$
0)
#973980000000
1"
1'
b0 +
b0 1
#974030000000
0"
0'
#974040000000
1#
1(
b101111101100100 +
b101111101100100 1
#974090000000
0#
0(
#974100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#974150000000
0$
0)
#974160000000
1"
1'
b0 +
b0 1
#974210000000
0"
0'
#974220000000
1#
1(
b101111101100100 +
b101111101100100 1
#974270000000
0#
0(
#974280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#974330000000
0$
0)
#974340000000
1"
1'
b0 +
b0 1
#974390000000
0"
0'
#974400000000
1#
1(
b101111101100100 +
b101111101100100 1
#974450000000
0#
0(
#974460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#974510000000
0$
0)
#974520000000
1"
1'
b0 +
b0 1
#974570000000
0"
0'
#974580000000
1#
1(
b101111101100100 +
b101111101100100 1
#974630000000
0#
0(
#974640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#974690000000
0$
0)
#974700000000
1"
1'
b0 +
b0 1
#974750000000
0"
0'
#974760000000
1#
1(
b101111101100100 +
b101111101100100 1
#974810000000
0#
0(
#974820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#974870000000
0$
0)
#974880000000
1"
1'
b0 +
b0 1
#974930000000
0"
0'
#974940000000
1#
1(
b101111101100100 +
b101111101100100 1
#974990000000
0#
0(
#975000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#975050000000
0$
0)
#975060000000
1"
1'
b0 +
b0 1
#975110000000
0"
0'
#975120000000
1#
1(
b101111101100100 +
b101111101100100 1
#975170000000
0#
0(
#975180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#975230000000
0$
0)
#975240000000
1"
1'
b0 +
b0 1
#975290000000
0"
0'
#975300000000
1#
1(
b101111101100100 +
b101111101100100 1
#975350000000
0#
0(
#975360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#975410000000
0$
0)
#975420000000
1"
1'
b0 +
b0 1
#975470000000
0"
0'
#975480000000
1#
1(
b101111101100100 +
b101111101100100 1
#975530000000
0#
0(
#975540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#975590000000
0$
0)
#975600000000
1"
1'
b0 +
b0 1
#975650000000
0"
0'
#975660000000
1#
1(
b101111101100100 +
b101111101100100 1
#975710000000
0#
0(
#975720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#975770000000
0$
0)
#975780000000
1"
1'
b0 +
b0 1
#975830000000
0"
0'
#975840000000
1#
1(
b101111101100100 +
b101111101100100 1
#975890000000
0#
0(
#975900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#975950000000
0$
0)
#975960000000
1"
1'
b0 +
b0 1
#976010000000
0"
0'
#976020000000
1#
1(
b101111101100100 +
b101111101100100 1
#976070000000
0#
0(
#976080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#976130000000
0$
0)
#976140000000
1"
1'
b0 +
b0 1
#976190000000
0"
0'
#976200000000
1#
1(
b101111101100100 +
b101111101100100 1
#976250000000
0#
0(
#976260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#976310000000
0$
0)
#976320000000
1"
1'
b0 +
b0 1
#976370000000
0"
0'
#976380000000
1#
1(
b101111101100100 +
b101111101100100 1
#976430000000
0#
0(
#976440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#976490000000
0$
0)
#976500000000
1"
1'
b0 +
b0 1
#976550000000
0"
0'
#976560000000
1#
1(
b101111101100100 +
b101111101100100 1
#976610000000
0#
0(
#976620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#976670000000
0$
0)
#976680000000
1"
1'
b0 +
b0 1
#976730000000
0"
0'
#976740000000
1#
1(
b101111101100100 +
b101111101100100 1
#976790000000
0#
0(
#976800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#976850000000
0$
0)
#976860000000
1"
1'
b0 +
b0 1
#976910000000
0"
0'
#976920000000
1#
1(
b101111101100100 +
b101111101100100 1
#976970000000
0#
0(
#976980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#977030000000
0$
0)
#977040000000
1"
1'
b0 +
b0 1
#977090000000
0"
0'
#977100000000
1#
1(
b101111101100100 +
b101111101100100 1
#977150000000
0#
0(
#977160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#977210000000
0$
0)
#977220000000
1"
1'
b0 +
b0 1
#977270000000
0"
0'
#977280000000
1#
1(
b101111101100100 +
b101111101100100 1
#977330000000
0#
0(
#977340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#977390000000
0$
0)
#977400000000
1"
1'
b0 +
b0 1
#977450000000
0"
0'
#977460000000
1#
1(
b101111101100100 +
b101111101100100 1
#977510000000
0#
0(
#977520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#977570000000
0$
0)
#977580000000
1"
1'
b0 +
b0 1
#977630000000
0"
0'
#977640000000
1#
1(
b101111101100100 +
b101111101100100 1
#977690000000
0#
0(
#977700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#977750000000
0$
0)
#977760000000
1"
1'
b0 +
b0 1
#977810000000
0"
0'
#977820000000
1#
1(
b101111101100100 +
b101111101100100 1
#977870000000
0#
0(
#977880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#977930000000
0$
0)
#977940000000
1"
1'
b0 +
b0 1
#977990000000
0"
0'
#978000000000
1#
1(
b101111101100100 +
b101111101100100 1
#978050000000
0#
0(
#978060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#978110000000
0$
0)
#978120000000
1"
1'
b0 +
b0 1
#978170000000
0"
0'
#978180000000
1#
1(
b101111101100100 +
b101111101100100 1
#978230000000
0#
0(
#978240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#978290000000
0$
0)
#978300000000
1"
1'
b0 +
b0 1
#978350000000
0"
0'
#978360000000
1#
1(
b101111101100100 +
b101111101100100 1
#978410000000
0#
0(
#978420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#978470000000
0$
0)
#978480000000
1"
1'
b0 +
b0 1
#978530000000
0"
0'
#978540000000
1#
1(
b101111101100100 +
b101111101100100 1
#978590000000
0#
0(
#978600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#978650000000
0$
0)
#978660000000
1"
1'
b0 +
b0 1
#978710000000
0"
0'
#978720000000
1#
1(
b101111101100100 +
b101111101100100 1
#978770000000
0#
0(
#978780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#978830000000
0$
0)
#978840000000
1"
1'
b0 +
b0 1
#978890000000
0"
0'
#978900000000
1#
1(
b101111101100100 +
b101111101100100 1
#978950000000
0#
0(
#978960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#979010000000
0$
0)
#979020000000
1"
1'
b0 +
b0 1
#979070000000
0"
0'
#979080000000
1#
1(
b101111101100100 +
b101111101100100 1
#979130000000
0#
0(
#979140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#979190000000
0$
0)
#979200000000
1"
1'
b0 +
b0 1
#979250000000
0"
0'
#979260000000
1#
1(
b101111101100100 +
b101111101100100 1
#979310000000
0#
0(
#979320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#979370000000
0$
0)
#979380000000
1"
1'
b0 +
b0 1
#979430000000
0"
0'
#979440000000
1#
1(
b101111101100100 +
b101111101100100 1
#979490000000
0#
0(
#979500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#979550000000
0$
0)
#979560000000
1"
1'
b0 +
b0 1
#979610000000
0"
0'
#979620000000
1#
1(
b101111101100100 +
b101111101100100 1
#979670000000
0#
0(
#979680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#979730000000
0$
0)
#979740000000
1"
1'
b0 +
b0 1
#979790000000
0"
0'
#979800000000
1#
1(
b101111101100100 +
b101111101100100 1
#979850000000
0#
0(
#979860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#979910000000
0$
0)
#979920000000
1"
1'
b0 +
b0 1
#979970000000
0"
0'
#979980000000
1#
1(
b101111101100100 +
b101111101100100 1
#980030000000
0#
0(
#980040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#980090000000
0$
0)
#980100000000
1"
1'
b0 +
b0 1
#980150000000
0"
0'
#980160000000
1#
1(
b101111101100100 +
b101111101100100 1
#980210000000
0#
0(
#980220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#980270000000
0$
0)
#980280000000
1"
1'
b0 +
b0 1
#980330000000
0"
0'
#980340000000
1#
1(
b101111101100100 +
b101111101100100 1
#980390000000
0#
0(
#980400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#980450000000
0$
0)
#980460000000
1"
1'
b0 +
b0 1
#980510000000
0"
0'
#980520000000
1#
1(
b101111101100100 +
b101111101100100 1
#980570000000
0#
0(
#980580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#980630000000
0$
0)
#980640000000
1"
1'
b0 +
b0 1
#980690000000
0"
0'
#980700000000
1#
1(
b101111101100100 +
b101111101100100 1
#980750000000
0#
0(
#980760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#980810000000
0$
0)
#980820000000
1"
1'
b0 +
b0 1
#980870000000
0"
0'
#980880000000
1#
1(
b101111101100100 +
b101111101100100 1
#980930000000
0#
0(
#980940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#980990000000
0$
0)
#981000000000
1"
1'
b0 +
b0 1
#981050000000
0"
0'
#981060000000
1#
1(
b101111101100100 +
b101111101100100 1
#981110000000
0#
0(
#981120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#981170000000
0$
0)
#981180000000
1"
1'
b0 +
b0 1
#981230000000
0"
0'
#981240000000
1#
1(
b101111101100100 +
b101111101100100 1
#981290000000
0#
0(
#981300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#981350000000
0$
0)
#981360000000
1"
1'
b0 +
b0 1
#981410000000
0"
0'
#981420000000
1#
1(
b101111101100100 +
b101111101100100 1
#981470000000
0#
0(
#981480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#981530000000
0$
0)
#981540000000
1"
1'
b0 +
b0 1
#981590000000
0"
0'
#981600000000
1#
1(
b101111101100100 +
b101111101100100 1
#981650000000
0#
0(
#981660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#981710000000
0$
0)
#981720000000
1"
1'
b0 +
b0 1
#981770000000
0"
0'
#981780000000
1#
1(
b101111101100100 +
b101111101100100 1
#981830000000
0#
0(
#981840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#981890000000
0$
0)
#981900000000
1"
1'
b0 +
b0 1
#981950000000
0"
0'
#981960000000
1#
1(
b101111101100100 +
b101111101100100 1
#982010000000
0#
0(
#982020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#982070000000
0$
0)
#982080000000
1"
1'
b0 +
b0 1
#982130000000
0"
0'
#982140000000
1#
1(
b101111101100100 +
b101111101100100 1
#982190000000
0#
0(
#982200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#982250000000
0$
0)
#982260000000
1"
1'
b0 +
b0 1
#982310000000
0"
0'
#982320000000
1#
1(
b101111101100100 +
b101111101100100 1
#982370000000
0#
0(
#982380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#982430000000
0$
0)
#982440000000
1"
1'
b0 +
b0 1
#982490000000
0"
0'
#982500000000
1#
1(
b101111101100100 +
b101111101100100 1
#982550000000
0#
0(
#982560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#982610000000
0$
0)
#982620000000
1"
1'
b0 +
b0 1
#982670000000
0"
0'
#982680000000
1#
1(
b101111101100100 +
b101111101100100 1
#982730000000
0#
0(
#982740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#982790000000
0$
0)
#982800000000
1"
1'
b0 +
b0 1
#982850000000
0"
0'
#982860000000
1#
1(
b101111101100100 +
b101111101100100 1
#982910000000
0#
0(
#982920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#982970000000
0$
0)
#982980000000
1"
1'
b0 +
b0 1
#983030000000
0"
0'
#983040000000
1#
1(
b101111101100100 +
b101111101100100 1
#983090000000
0#
0(
#983100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#983150000000
0$
0)
#983160000000
1"
1'
b0 +
b0 1
#983210000000
0"
0'
#983220000000
1#
1(
b101111101100100 +
b101111101100100 1
#983270000000
0#
0(
#983280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#983330000000
0$
0)
#983340000000
1"
1'
b0 +
b0 1
#983390000000
0"
0'
#983400000000
1#
1(
b101111101100100 +
b101111101100100 1
#983450000000
0#
0(
#983460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#983510000000
0$
0)
#983520000000
1"
1'
b0 +
b0 1
#983570000000
0"
0'
#983580000000
1#
1(
b101111101100100 +
b101111101100100 1
#983630000000
0#
0(
#983640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#983690000000
0$
0)
#983700000000
1"
1'
b0 +
b0 1
#983750000000
0"
0'
#983760000000
1#
1(
b101111101100100 +
b101111101100100 1
#983810000000
0#
0(
#983820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#983870000000
0$
0)
#983880000000
1"
1'
b0 +
b0 1
#983930000000
0"
0'
#983940000000
1#
1(
b101111101100100 +
b101111101100100 1
#983990000000
0#
0(
#984000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#984050000000
0$
0)
#984060000000
1"
1'
b0 +
b0 1
#984110000000
0"
0'
#984120000000
1#
1(
b101111101100100 +
b101111101100100 1
#984170000000
0#
0(
#984180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#984230000000
0$
0)
#984240000000
1"
1'
b0 +
b0 1
#984290000000
0"
0'
#984300000000
1#
1(
b101111101100100 +
b101111101100100 1
#984350000000
0#
0(
#984360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#984410000000
0$
0)
#984420000000
1"
1'
b0 +
b0 1
#984470000000
0"
0'
#984480000000
1#
1(
b101111101100100 +
b101111101100100 1
#984530000000
0#
0(
#984540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#984590000000
0$
0)
#984600000000
1"
1'
b0 +
b0 1
#984650000000
0"
0'
#984660000000
1#
1(
b101111101100100 +
b101111101100100 1
#984710000000
0#
0(
#984720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#984770000000
0$
0)
#984780000000
1"
1'
b0 +
b0 1
#984830000000
0"
0'
#984840000000
1#
1(
b101111101100100 +
b101111101100100 1
#984890000000
0#
0(
#984900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#984950000000
0$
0)
#984960000000
1"
1'
b0 +
b0 1
#985010000000
0"
0'
#985020000000
1#
1(
b101111101100100 +
b101111101100100 1
#985070000000
0#
0(
#985080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#985130000000
0$
0)
#985140000000
1"
1'
b0 +
b0 1
#985190000000
0"
0'
#985200000000
1#
1(
b101111101100100 +
b101111101100100 1
#985250000000
0#
0(
#985260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#985310000000
0$
0)
#985320000000
1"
1'
b0 +
b0 1
#985370000000
0"
0'
#985380000000
1#
1(
b101111101100100 +
b101111101100100 1
#985430000000
0#
0(
#985440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#985490000000
0$
0)
#985500000000
1"
1'
b0 +
b0 1
#985550000000
0"
0'
#985560000000
1#
1(
b101111101100100 +
b101111101100100 1
#985610000000
0#
0(
#985620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#985670000000
0$
0)
#985680000000
1"
1'
b0 +
b0 1
#985730000000
0"
0'
#985740000000
1#
1(
b101111101100100 +
b101111101100100 1
#985790000000
0#
0(
#985800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#985850000000
0$
0)
#985860000000
1"
1'
b0 +
b0 1
#985910000000
0"
0'
#985920000000
1#
1(
b101111101100100 +
b101111101100100 1
#985970000000
0#
0(
#985980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#986030000000
0$
0)
#986040000000
1"
1'
b0 +
b0 1
#986090000000
0"
0'
#986100000000
1#
1(
b101111101100100 +
b101111101100100 1
#986150000000
0#
0(
#986160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#986210000000
0$
0)
#986220000000
1"
1'
b0 +
b0 1
#986270000000
0"
0'
#986280000000
1#
1(
b101111101100100 +
b101111101100100 1
#986330000000
0#
0(
#986340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#986390000000
0$
0)
#986400000000
1"
1'
b0 +
b0 1
#986450000000
0"
0'
#986460000000
1#
1(
b101111101100100 +
b101111101100100 1
#986510000000
0#
0(
#986520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#986570000000
0$
0)
#986580000000
1"
1'
b0 +
b0 1
#986630000000
0"
0'
#986640000000
1#
1(
b101111101100100 +
b101111101100100 1
#986690000000
0#
0(
#986700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#986750000000
0$
0)
#986760000000
1"
1'
b0 +
b0 1
#986810000000
0"
0'
#986820000000
1#
1(
b101111101100100 +
b101111101100100 1
#986870000000
0#
0(
#986880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#986930000000
0$
0)
#986940000000
1"
1'
b0 +
b0 1
#986990000000
0"
0'
#987000000000
1#
1(
b101111101100100 +
b101111101100100 1
#987050000000
0#
0(
#987060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#987110000000
0$
0)
#987120000000
1"
1'
b0 +
b0 1
#987170000000
0"
0'
#987180000000
1#
1(
b101111101100100 +
b101111101100100 1
#987230000000
0#
0(
#987240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#987290000000
0$
0)
#987300000000
1"
1'
b0 +
b0 1
#987350000000
0"
0'
#987360000000
1#
1(
b101111101100100 +
b101111101100100 1
#987410000000
0#
0(
#987420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#987470000000
0$
0)
#987480000000
1"
1'
b0 +
b0 1
#987530000000
0"
0'
#987540000000
1#
1(
b101111101100100 +
b101111101100100 1
#987590000000
0#
0(
#987600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#987650000000
0$
0)
#987660000000
1"
1'
b0 +
b0 1
#987710000000
0"
0'
#987720000000
1#
1(
b101111101100100 +
b101111101100100 1
#987770000000
0#
0(
#987780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#987830000000
0$
0)
#987840000000
1"
1'
b0 +
b0 1
#987890000000
0"
0'
#987900000000
1#
1(
b101111101100100 +
b101111101100100 1
#987950000000
0#
0(
#987960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#988010000000
0$
0)
#988020000000
1"
1'
b0 +
b0 1
#988070000000
0"
0'
#988080000000
1#
1(
b101111101100100 +
b101111101100100 1
#988130000000
0#
0(
#988140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#988190000000
0$
0)
#988200000000
1"
1'
b0 +
b0 1
#988250000000
0"
0'
#988260000000
1#
1(
b101111101100100 +
b101111101100100 1
#988310000000
0#
0(
#988320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#988370000000
0$
0)
#988380000000
1"
1'
b0 +
b0 1
#988430000000
0"
0'
#988440000000
1#
1(
b101111101100100 +
b101111101100100 1
#988490000000
0#
0(
#988500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#988550000000
0$
0)
#988560000000
1"
1'
b0 +
b0 1
#988610000000
0"
0'
#988620000000
1#
1(
b101111101100100 +
b101111101100100 1
#988670000000
0#
0(
#988680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#988730000000
0$
0)
#988740000000
1"
1'
b0 +
b0 1
#988790000000
0"
0'
#988800000000
1#
1(
b101111101100100 +
b101111101100100 1
#988850000000
0#
0(
#988860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#988910000000
0$
0)
#988920000000
1"
1'
b0 +
b0 1
#988970000000
0"
0'
#988980000000
1#
1(
b101111101100100 +
b101111101100100 1
#989030000000
0#
0(
#989040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#989090000000
0$
0)
#989100000000
1"
1'
b0 +
b0 1
#989150000000
0"
0'
#989160000000
1#
1(
b101111101100100 +
b101111101100100 1
#989210000000
0#
0(
#989220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#989270000000
0$
0)
#989280000000
1"
1'
b0 +
b0 1
#989330000000
0"
0'
#989340000000
1#
1(
b101111101100100 +
b101111101100100 1
#989390000000
0#
0(
#989400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#989450000000
0$
0)
#989460000000
1"
1'
b0 +
b0 1
#989510000000
0"
0'
#989520000000
1#
1(
b101111101100100 +
b101111101100100 1
#989570000000
0#
0(
#989580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#989630000000
0$
0)
#989640000000
1"
1'
b0 +
b0 1
#989690000000
0"
0'
#989700000000
1#
1(
b101111101100100 +
b101111101100100 1
#989750000000
0#
0(
#989760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#989810000000
0$
0)
#989820000000
1"
1'
b0 +
b0 1
#989870000000
0"
0'
#989880000000
1#
1(
b101111101100100 +
b101111101100100 1
#989930000000
0#
0(
#989940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#989990000000
0$
0)
#990000000000
1"
1'
b0 +
b0 1
#990050000000
0"
0'
#990060000000
1#
1(
b101111101100100 +
b101111101100100 1
#990110000000
0#
0(
#990120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#990170000000
0$
0)
#990180000000
1"
1'
b0 +
b0 1
#990230000000
0"
0'
#990240000000
1#
1(
b101111101100100 +
b101111101100100 1
#990290000000
0#
0(
#990300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#990350000000
0$
0)
#990360000000
1"
1'
b0 +
b0 1
#990410000000
0"
0'
#990420000000
1#
1(
b101111101100100 +
b101111101100100 1
#990470000000
0#
0(
#990480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#990530000000
0$
0)
#990540000000
1"
1'
b0 +
b0 1
#990590000000
0"
0'
#990600000000
1#
1(
b101111101100100 +
b101111101100100 1
#990650000000
0#
0(
#990660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#990710000000
0$
0)
#990720000000
1"
1'
b0 +
b0 1
#990770000000
0"
0'
#990780000000
1#
1(
b101111101100100 +
b101111101100100 1
#990830000000
0#
0(
#990840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#990890000000
0$
0)
#990900000000
1"
1'
b0 +
b0 1
#990950000000
0"
0'
#990960000000
1#
1(
b101111101100100 +
b101111101100100 1
#991010000000
0#
0(
#991020000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#991070000000
0$
0)
#991080000000
1"
1'
b0 +
b0 1
#991130000000
0"
0'
#991140000000
1#
1(
b101111101100100 +
b101111101100100 1
#991190000000
0#
0(
#991200000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#991250000000
0$
0)
#991260000000
1"
1'
b0 +
b0 1
#991310000000
0"
0'
#991320000000
1#
1(
b101111101100100 +
b101111101100100 1
#991370000000
0#
0(
#991380000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#991430000000
0$
0)
#991440000000
1"
1'
b0 +
b0 1
#991490000000
0"
0'
#991500000000
1#
1(
b101111101100100 +
b101111101100100 1
#991550000000
0#
0(
#991560000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#991610000000
0$
0)
#991620000000
1"
1'
b0 +
b0 1
#991670000000
0"
0'
#991680000000
1#
1(
b101111101100100 +
b101111101100100 1
#991730000000
0#
0(
#991740000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#991790000000
0$
0)
#991800000000
1"
1'
b0 +
b0 1
#991850000000
0"
0'
#991860000000
1#
1(
b101111101100100 +
b101111101100100 1
#991910000000
0#
0(
#991920000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#991970000000
0$
0)
#991980000000
1"
1'
b0 +
b0 1
#992030000000
0"
0'
#992040000000
1#
1(
b101111101100100 +
b101111101100100 1
#992090000000
0#
0(
#992100000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#992150000000
0$
0)
#992160000000
1"
1'
b0 +
b0 1
#992210000000
0"
0'
#992220000000
1#
1(
b101111101100100 +
b101111101100100 1
#992270000000
0#
0(
#992280000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#992330000000
0$
0)
#992340000000
1"
1'
b0 +
b0 1
#992390000000
0"
0'
#992400000000
1#
1(
b101111101100100 +
b101111101100100 1
#992450000000
0#
0(
#992460000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#992510000000
0$
0)
#992520000000
1"
1'
b0 +
b0 1
#992570000000
0"
0'
#992580000000
1#
1(
b101111101100100 +
b101111101100100 1
#992630000000
0#
0(
#992640000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#992690000000
0$
0)
#992700000000
1"
1'
b0 +
b0 1
#992750000000
0"
0'
#992760000000
1#
1(
b101111101100100 +
b101111101100100 1
#992810000000
0#
0(
#992820000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#992870000000
0$
0)
#992880000000
1"
1'
b0 +
b0 1
#992930000000
0"
0'
#992940000000
1#
1(
b101111101100100 +
b101111101100100 1
#992990000000
0#
0(
#993000000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#993050000000
0$
0)
#993060000000
1"
1'
b0 +
b0 1
#993110000000
0"
0'
#993120000000
1#
1(
b101111101100100 +
b101111101100100 1
#993170000000
0#
0(
#993180000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#993230000000
0$
0)
#993240000000
1"
1'
b0 +
b0 1
#993290000000
0"
0'
#993300000000
1#
1(
b101111101100100 +
b101111101100100 1
#993350000000
0#
0(
#993360000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#993410000000
0$
0)
#993420000000
1"
1'
b0 +
b0 1
#993470000000
0"
0'
#993480000000
1#
1(
b101111101100100 +
b101111101100100 1
#993530000000
0#
0(
#993540000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#993590000000
0$
0)
#993600000000
1"
1'
b0 +
b0 1
#993650000000
0"
0'
#993660000000
1#
1(
b101111101100100 +
b101111101100100 1
#993710000000
0#
0(
#993720000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#993770000000
0$
0)
#993780000000
1"
1'
b0 +
b0 1
#993830000000
0"
0'
#993840000000
1#
1(
b101111101100100 +
b101111101100100 1
#993890000000
0#
0(
#993900000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#993950000000
0$
0)
#993960000000
1"
1'
b0 +
b0 1
#994010000000
0"
0'
#994020000000
1#
1(
b101111101100100 +
b101111101100100 1
#994070000000
0#
0(
#994080000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#994130000000
0$
0)
#994140000000
1"
1'
b0 +
b0 1
#994190000000
0"
0'
#994200000000
1#
1(
b101111101100100 +
b101111101100100 1
#994250000000
0#
0(
#994260000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#994310000000
0$
0)
#994320000000
1"
1'
b0 +
b0 1
#994370000000
0"
0'
#994380000000
1#
1(
b101111101100100 +
b101111101100100 1
#994430000000
0#
0(
#994440000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#994490000000
0$
0)
#994500000000
1"
1'
b0 +
b0 1
#994550000000
0"
0'
#994560000000
1#
1(
b101111101100100 +
b101111101100100 1
#994610000000
0#
0(
#994620000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#994670000000
0$
0)
#994680000000
1"
1'
b0 +
b0 1
#994730000000
0"
0'
#994740000000
1#
1(
b101111101100100 +
b101111101100100 1
#994790000000
0#
0(
#994800000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#994850000000
0$
0)
#994860000000
1"
1'
b0 +
b0 1
#994910000000
0"
0'
#994920000000
1#
1(
b101111101100100 +
b101111101100100 1
#994970000000
0#
0(
#994980000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#995030000000
0$
0)
#995040000000
1"
1'
b0 +
b0 1
#995090000000
0"
0'
#995100000000
1#
1(
b101111101100100 +
b101111101100100 1
#995150000000
0#
0(
#995160000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#995210000000
0$
0)
#995220000000
1"
1'
b0 +
b0 1
#995270000000
0"
0'
#995280000000
1#
1(
b101111101100100 +
b101111101100100 1
#995330000000
0#
0(
#995340000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#995390000000
0$
0)
#995400000000
1"
1'
b0 +
b0 1
#995450000000
0"
0'
#995460000000
1#
1(
b101111101100100 +
b101111101100100 1
#995510000000
0#
0(
#995520000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#995570000000
0$
0)
#995580000000
1"
1'
b0 +
b0 1
#995630000000
0"
0'
#995640000000
1#
1(
b101111101100100 +
b101111101100100 1
#995690000000
0#
0(
#995700000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#995750000000
0$
0)
#995760000000
1"
1'
b0 +
b0 1
#995810000000
0"
0'
#995820000000
1#
1(
b101111101100100 +
b101111101100100 1
#995870000000
0#
0(
#995880000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#995930000000
0$
0)
#995940000000
1"
1'
b0 +
b0 1
#995990000000
0"
0'
#996000000000
1#
1(
b101111101100100 +
b101111101100100 1
#996050000000
0#
0(
#996060000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#996110000000
0$
0)
#996120000000
1"
1'
b0 +
b0 1
#996170000000
0"
0'
#996180000000
1#
1(
b101111101100100 +
b101111101100100 1
#996230000000
0#
0(
#996240000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#996290000000
0$
0)
#996300000000
1"
1'
b0 +
b0 1
#996350000000
0"
0'
#996360000000
1#
1(
b101111101100100 +
b101111101100100 1
#996410000000
0#
0(
#996420000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#996470000000
0$
0)
#996480000000
1"
1'
b0 +
b0 1
#996530000000
0"
0'
#996540000000
1#
1(
b101111101100100 +
b101111101100100 1
#996590000000
0#
0(
#996600000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#996650000000
0$
0)
#996660000000
1"
1'
b0 +
b0 1
#996710000000
0"
0'
#996720000000
1#
1(
b101111101100100 +
b101111101100100 1
#996770000000
0#
0(
#996780000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#996830000000
0$
0)
#996840000000
1"
1'
b0 +
b0 1
#996890000000
0"
0'
#996900000000
1#
1(
b101111101100100 +
b101111101100100 1
#996950000000
0#
0(
#996960000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#997010000000
0$
0)
#997020000000
1"
1'
b0 +
b0 1
#997070000000
0"
0'
#997080000000
1#
1(
b101111101100100 +
b101111101100100 1
#997130000000
0#
0(
#997140000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#997190000000
0$
0)
#997200000000
1"
1'
b0 +
b0 1
#997250000000
0"
0'
#997260000000
1#
1(
b101111101100100 +
b101111101100100 1
#997310000000
0#
0(
#997320000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#997370000000
0$
0)
#997380000000
1"
1'
b0 +
b0 1
#997430000000
0"
0'
#997440000000
1#
1(
b101111101100100 +
b101111101100100 1
#997490000000
0#
0(
#997500000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#997550000000
0$
0)
#997560000000
1"
1'
b0 +
b0 1
#997610000000
0"
0'
#997620000000
1#
1(
b101111101100100 +
b101111101100100 1
#997670000000
0#
0(
#997680000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#997730000000
0$
0)
#997740000000
1"
1'
b0 +
b0 1
#997790000000
0"
0'
#997800000000
1#
1(
b101111101100100 +
b101111101100100 1
#997850000000
0#
0(
#997860000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#997910000000
0$
0)
#997920000000
1"
1'
b0 +
b0 1
#997970000000
0"
0'
#997980000000
1#
1(
b101111101100100 +
b101111101100100 1
#998030000000
0#
0(
#998040000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#998090000000
0$
0)
#998100000000
1"
1'
b0 +
b0 1
#998150000000
0"
0'
#998160000000
1#
1(
b101111101100100 +
b101111101100100 1
#998210000000
0#
0(
#998220000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#998270000000
0$
0)
#998280000000
1"
1'
b0 +
b0 1
#998330000000
0"
0'
#998340000000
1#
1(
b101111101100100 +
b101111101100100 1
#998390000000
0#
0(
#998400000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#998450000000
0$
0)
#998460000000
1"
1'
b0 +
b0 1
#998510000000
0"
0'
#998520000000
1#
1(
b101111101100100 +
b101111101100100 1
#998570000000
0#
0(
#998580000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#998630000000
0$
0)
#998640000000
1"
1'
b0 +
b0 1
#998690000000
0"
0'
#998700000000
1#
1(
b101111101100100 +
b101111101100100 1
#998750000000
0#
0(
#998760000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#998810000000
0$
0)
#998820000000
1"
1'
b0 +
b0 1
#998870000000
0"
0'
#998880000000
1#
1(
b101111101100100 +
b101111101100100 1
#998930000000
0#
0(
#998940000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#998990000000
0$
0)
#999000000000
1"
1'
b0 +
b0 1
#999050000000
0"
0'
#999060000000
1#
1(
b101111101100100 +
b101111101100100 1
#999110000000
0#
0(
#999120000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#999170000000
0$
0)
#999180000000
1"
1'
b0 +
b0 1
#999230000000
0"
0'
#999240000000
1#
1(
b101111101100100 +
b101111101100100 1
#999290000000
0#
0(
#999300000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#999350000000
0$
0)
#999360000000
1"
1'
b0 +
b0 1
#999410000000
0"
0'
#999420000000
1#
1(
b101111101100100 +
b101111101100100 1
#999470000000
0#
0(
#999480000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#999530000000
0$
0)
#999540000000
1"
1'
b0 +
b0 1
#999590000000
0"
0'
#999600000000
1#
1(
b101111101100100 +
b101111101100100 1
#999650000000
0#
0(
#999660000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#999710000000
0$
0)
#999720000000
1"
1'
b0 +
b0 1
#999770000000
0"
0'
#999780000000
1#
1(
b101111101100100 +
b101111101100100 1
#999830000000
0#
0(
#999840000000
1$
1)
b1100001101000011 +
b1100001101000011 1
#999890000000
0$
0)
#999900000000
1"
1'
b0 +
b0 1
#999950000000
0"
0'
#999960000000
1#
1(
b101111101100100 +
b101111101100100 1
