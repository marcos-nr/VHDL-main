$date
  Tue May 07 00:24:10 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp2_3 $end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 4 # enable_disp[3:0] $end
$var reg 7 $ segmentos[6:0] $end
$scope module uut $end
$var reg 1 % clk $end
$var reg 1 & reset $end
$var reg 4 ' enable_disp[3:0] $end
$var reg 7 ( segmentos[6:0] $end
$comment state is not handled $end
$var reg 4 ) bcd[3:0] $end
$var integer 32 * cuenta $end
$var reg 1 + debounced_reset $end
$var reg 1 , clk_reset $end
$var reg 1 - enable_conta $end
$scope module a $end
$var reg 1 . clk $end
$var reg 1 / key $end
$var reg 1 0 debounced_key $end
$var reg 1 1 key_stable $end
$var reg 1 2 last_key $end
$upscope $end
$scope module b $end
$var reg 1 3 clk $end
$var reg 1 4 reset $end
$var reg 1 5 enable $end
$var reg 1 6 cout $end
$var integer 32 7 q $end
$upscope $end
$scope module d $end
$var reg 7 8 segmentos[6:0] $end
$var reg 4 9 bcd[3:0] $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
1"
b1000 #
b0110000 $
0%
1&
b1000 '
b0110000 (
b0001 )
b0 *
U+
0,
1-
0.
1/
U0
U1
U2
03
04
15
U6
b0 7
b0110000 8
b0001 9
#10000000
1!
1%
1+
1.
10
11
12
13
06
#20000000
0!
0%
b1 *
0.
03
b1 7
#30000000
1!
1%
1.
13
#40000000
0!
0%
b10 *
0.
03
b10 7
#50000000
1!
1%
1.
13
#60000000
0!
0%
b11 *
0.
03
b11 7
#70000000
1!
1%
1.
13
16
#80000000
0!
0%
b100 *
0.
03
b100 7
#90000000
1!
1%
1.
13
#100000000
0!
0%
b101 *
0.
03
b101 7
#110000000
1!
1%
1.
13
#120000000
0!
0%
b110 *
0.
03
b110 7
#130000000
1!
1%
1.
13
#140000000
0!
0%
b111 *
0.
03
b111 7
#150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#160000000
0!
0"
0%
0&
b0 *
0.
0/
03
b0 7
#170000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#180000000
0!
0%
b1 *
0.
03
b1 7
#190000000
1!
1%
1.
13
#200000000
0!
0%
b10 *
0.
03
b10 7
#210000000
1!
1%
1.
13
#220000000
0!
0%
b11 *
0.
03
b11 7
#230000000
1!
1%
1.
13
16
#240000000
0!
0%
b100 *
0.
03
b100 7
#250000000
1!
1%
1.
13
#260000000
0!
0%
b101 *
0.
03
b101 7
#270000000
1!
1%
1.
13
#280000000
0!
0%
b110 *
0.
03
b110 7
#290000000
1!
1%
1.
13
#300000000
0!
0%
b111 *
0.
03
b111 7
#310000000
1!
1%
1.
13
06
#320000000
0!
0%
b0 *
0.
03
b0 7
#330000000
1!
1%
1.
13
#340000000
0!
0%
b1 *
0.
03
b1 7
#350000000
1!
1%
1.
13
#360000000
0!
0%
b10 *
0.
03
b10 7
#370000000
1!
1%
1.
13
#380000000
0!
0%
b11 *
0.
03
b11 7
#390000000
1!
1%
1.
13
16
#400000000
0!
0%
b100 *
0.
03
b100 7
#410000000
1!
1%
1.
13
#420000000
0!
0%
b101 *
0.
03
b101 7
#430000000
1!
1%
1.
13
#440000000
0!
0%
b110 *
0.
03
b110 7
#450000000
1!
1%
1.
13
#460000000
0!
0%
b111 *
0.
03
b111 7
#470000000
1!
1%
1.
13
06
#480000000
0!
0%
b0 *
0.
03
b0 7
#490000000
1!
1%
1.
13
#500000000
0!
0%
b1 *
0.
03
b1 7
#510000000
1!
1%
1.
13
#520000000
0!
0%
b10 *
0.
03
b10 7
#530000000
1!
1%
1.
13
#540000000
0!
0%
b11 *
0.
03
b11 7
#550000000
1!
1%
1.
13
16
#560000000
0!
0%
b100 *
0.
03
b100 7
#570000000
1!
1%
1.
13
#580000000
0!
0%
b101 *
0.
03
b101 7
#590000000
1!
1%
1.
13
#600000000
0!
0%
b110 *
0.
03
b110 7
#610000000
1!
1%
1.
13
#620000000
0!
0%
b111 *
0.
03
b111 7
#630000000
1!
1%
1.
13
06
#640000000
0!
0%
b0 *
0.
03
b0 7
#650000000
1!
1%
1.
13
#660000000
0!
0%
b1 *
0.
03
b1 7
#670000000
1!
1%
1.
13
#680000000
0!
1"
0%
1&
b10 *
0.
1/
03
b10 7
#690000000
1!
1%
1+
1.
10
11
12
13
#700000000
0!
0%
b11 *
0.
03
b11 7
#710000000
1!
1%
1.
13
16
#720000000
0!
0%
b100 *
0.
03
b100 7
#730000000
1!
1%
1.
13
#740000000
0!
0%
b101 *
0.
03
b101 7
#750000000
1!
1%
1.
13
#760000000
0!
0%
b110 *
0.
03
b110 7
#770000000
1!
1%
1.
13
#780000000
0!
0%
b111 *
0.
03
b111 7
#790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#800000000
0!
0%
b0 *
0.
03
b0 7
#810000000
1!
1%
1.
13
#820000000
0!
0%
b1 *
0.
03
b1 7
#830000000
1!
1%
1.
13
#840000000
0!
0"
0%
0&
b10 *
0.
0/
03
b10 7
#850000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#860000000
0!
0%
b11 *
0.
03
b11 7
#870000000
1!
1%
1.
13
16
#880000000
0!
0%
b100 *
0.
03
b100 7
#890000000
1!
1%
1.
13
#900000000
0!
0%
b101 *
0.
03
b101 7
#910000000
1!
1%
1.
13
#920000000
0!
0%
b110 *
0.
03
b110 7
#930000000
1!
1%
1.
13
#940000000
0!
0%
b111 *
0.
03
b111 7
#950000000
1!
1%
1.
13
06
#960000000
0!
0%
b0 *
0.
03
b0 7
#970000000
1!
1%
1.
13
#980000000
0!
0%
b1 *
0.
03
b1 7
#990000000
1!
1%
1.
13
#1000000000
0!
0%
b10 *
0.
03
b10 7
#1010000000
1!
1%
1.
13
#1020000000
0!
0%
b11 *
0.
03
b11 7
#1030000000
1!
1%
1.
13
16
#1040000000
0!
0%
b100 *
0.
03
b100 7
#1050000000
1!
1%
1.
13
#1060000000
0!
0%
b101 *
0.
03
b101 7
#1070000000
1!
1%
1.
13
#1080000000
0!
0%
b110 *
0.
03
b110 7
#1090000000
1!
1%
1.
13
#1100000000
0!
0%
b111 *
0.
03
b111 7
#1110000000
1!
1%
1.
13
06
#1120000000
0!
0%
b0 *
0.
03
b0 7
#1130000000
1!
1%
1.
13
#1140000000
0!
0%
b1 *
0.
03
b1 7
#1150000000
1!
1%
1.
13
#1160000000
0!
0%
b10 *
0.
03
b10 7
#1170000000
1!
1%
1.
13
#1180000000
0!
0%
b11 *
0.
03
b11 7
#1190000000
1!
1%
1.
13
16
#1200000000
0!
0%
b100 *
0.
03
b100 7
#1210000000
1!
1%
1.
13
#1220000000
0!
0%
b101 *
0.
03
b101 7
#1230000000
1!
1%
1.
13
#1240000000
0!
0%
b110 *
0.
03
b110 7
#1250000000
1!
1%
1.
13
#1260000000
0!
0%
b111 *
0.
03
b111 7
#1270000000
1!
1%
1.
13
06
#1280000000
0!
0%
b0 *
0.
03
b0 7
#1290000000
1!
1%
1.
13
#1300000000
0!
0%
b1 *
0.
03
b1 7
#1310000000
1!
1%
1.
13
#1320000000
0!
0%
b10 *
0.
03
b10 7
#1330000000
1!
1%
1.
13
#1340000000
0!
0%
b11 *
0.
03
b11 7
#1350000000
1!
1%
1.
13
16
#1360000000
0!
1"
0%
1&
b100 *
0.
1/
03
b100 7
#1370000000
1!
1%
1+
1.
10
11
12
13
#1380000000
0!
0%
b101 *
0.
03
b101 7
#1390000000
1!
1%
1.
13
#1400000000
0!
0%
b110 *
0.
03
b110 7
#1410000000
1!
1%
1.
13
#1420000000
0!
0%
b111 *
0.
03
b111 7
#1430000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#1440000000
0!
0%
b0 *
0.
03
b0 7
#1450000000
1!
1%
1.
13
#1460000000
0!
0%
b1 *
0.
03
b1 7
#1470000000
1!
1%
1.
13
#1480000000
0!
0%
b10 *
0.
03
b10 7
#1490000000
1!
1%
1.
13
#1500000000
0!
0%
b11 *
0.
03
b11 7
#1510000000
1!
1%
1.
13
16
#1520000000
0!
0"
0%
0&
b100 *
0.
0/
03
b100 7
#1530000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#1540000000
0!
0%
b101 *
0.
03
b101 7
#1550000000
1!
1%
1.
13
#1560000000
0!
0%
b110 *
0.
03
b110 7
#1570000000
1!
1%
1.
13
#1580000000
0!
0%
b111 *
0.
03
b111 7
#1590000000
1!
1%
1.
13
06
#1600000000
0!
0%
b0 *
0.
03
b0 7
#1610000000
1!
1%
1.
13
#1620000000
0!
0%
b1 *
0.
03
b1 7
#1630000000
1!
1%
1.
13
#1640000000
0!
0%
b10 *
0.
03
b10 7
#1650000000
1!
1%
1.
13
#1660000000
0!
0%
b11 *
0.
03
b11 7
#1670000000
1!
1%
1.
13
16
#1680000000
0!
0%
b100 *
0.
03
b100 7
#1690000000
1!
1%
1.
13
#1700000000
0!
0%
b101 *
0.
03
b101 7
#1710000000
1!
1%
1.
13
#1720000000
0!
0%
b110 *
0.
03
b110 7
#1730000000
1!
1%
1.
13
#1740000000
0!
0%
b111 *
0.
03
b111 7
#1750000000
1!
1%
1.
13
06
#1760000000
0!
0%
b0 *
0.
03
b0 7
#1770000000
1!
1%
1.
13
#1780000000
0!
0%
b1 *
0.
03
b1 7
#1790000000
1!
1%
1.
13
#1800000000
0!
0%
b10 *
0.
03
b10 7
#1810000000
1!
1%
1.
13
#1820000000
0!
0%
b11 *
0.
03
b11 7
#1830000000
1!
1%
1.
13
16
#1840000000
0!
0%
b100 *
0.
03
b100 7
#1850000000
1!
1%
1.
13
#1860000000
0!
0%
b101 *
0.
03
b101 7
#1870000000
1!
1%
1.
13
#1880000000
0!
0%
b110 *
0.
03
b110 7
#1890000000
1!
1%
1.
13
#1900000000
0!
0%
b111 *
0.
03
b111 7
#1910000000
1!
1%
1.
13
06
#1920000000
0!
0%
b0 *
0.
03
b0 7
#1930000000
1!
1%
1.
13
#1940000000
0!
0%
b1 *
0.
03
b1 7
#1950000000
1!
1%
1.
13
#1960000000
0!
0%
b10 *
0.
03
b10 7
#1970000000
1!
1%
1.
13
#1980000000
0!
0%
b11 *
0.
03
b11 7
#1990000000
1!
1%
1.
13
16
#2000000000
0!
0%
b100 *
0.
03
b100 7
#2010000000
1!
1%
1.
13
#2020000000
0!
0%
b101 *
0.
03
b101 7
#2030000000
1!
1%
1.
13
#2040000000
0!
1"
0%
1&
b110 *
0.
1/
03
b110 7
#2050000000
1!
1%
1+
1.
10
11
12
13
#2060000000
0!
0%
b111 *
0.
03
b111 7
#2070000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#2080000000
0!
0%
b0 *
0.
03
b0 7
#2090000000
1!
1%
1.
13
#2100000000
0!
0%
b1 *
0.
03
b1 7
#2110000000
1!
1%
1.
13
#2120000000
0!
0%
b10 *
0.
03
b10 7
#2130000000
1!
1%
1.
13
#2140000000
0!
0%
b11 *
0.
03
b11 7
#2150000000
1!
1%
1.
13
16
#2160000000
0!
0%
b100 *
0.
03
b100 7
#2170000000
1!
1%
1.
13
#2180000000
0!
0%
b101 *
0.
03
b101 7
#2190000000
1!
1%
1.
13
#2200000000
0!
0"
0%
0&
b110 *
0.
0/
03
b110 7
#2210000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#2220000000
0!
0%
b111 *
0.
03
b111 7
#2230000000
1!
1%
1.
13
06
#2240000000
0!
0%
b0 *
0.
03
b0 7
#2250000000
1!
1%
1.
13
#2260000000
0!
0%
b1 *
0.
03
b1 7
#2270000000
1!
1%
1.
13
#2280000000
0!
0%
b10 *
0.
03
b10 7
#2290000000
1!
1%
1.
13
#2300000000
0!
0%
b11 *
0.
03
b11 7
#2310000000
1!
1%
1.
13
16
#2320000000
0!
0%
b100 *
0.
03
b100 7
#2330000000
1!
1%
1.
13
#2340000000
0!
0%
b101 *
0.
03
b101 7
#2350000000
1!
1%
1.
13
#2360000000
0!
0%
b110 *
0.
03
b110 7
#2370000000
1!
1%
1.
13
#2380000000
0!
0%
b111 *
0.
03
b111 7
#2390000000
1!
1%
1.
13
06
#2400000000
0!
0%
b0 *
0.
03
b0 7
#2410000000
1!
1%
1.
13
#2420000000
0!
0%
b1 *
0.
03
b1 7
#2430000000
1!
1%
1.
13
#2440000000
0!
0%
b10 *
0.
03
b10 7
#2450000000
1!
1%
1.
13
#2460000000
0!
0%
b11 *
0.
03
b11 7
#2470000000
1!
1%
1.
13
16
#2480000000
0!
0%
b100 *
0.
03
b100 7
#2490000000
1!
1%
1.
13
#2500000000
0!
0%
b101 *
0.
03
b101 7
#2510000000
1!
1%
1.
13
#2520000000
0!
0%
b110 *
0.
03
b110 7
#2530000000
1!
1%
1.
13
#2540000000
0!
0%
b111 *
0.
03
b111 7
#2550000000
1!
1%
1.
13
06
#2560000000
0!
0%
b0 *
0.
03
b0 7
#2570000000
1!
1%
1.
13
#2580000000
0!
0%
b1 *
0.
03
b1 7
#2590000000
1!
1%
1.
13
#2600000000
0!
0%
b10 *
0.
03
b10 7
#2610000000
1!
1%
1.
13
#2620000000
0!
0%
b11 *
0.
03
b11 7
#2630000000
1!
1%
1.
13
16
#2640000000
0!
0%
b100 *
0.
03
b100 7
#2650000000
1!
1%
1.
13
#2660000000
0!
0%
b101 *
0.
03
b101 7
#2670000000
1!
1%
1.
13
#2680000000
0!
0%
b110 *
0.
03
b110 7
#2690000000
1!
1%
1.
13
#2700000000
0!
0%
b111 *
0.
03
b111 7
#2710000000
1!
1%
1.
13
06
#2720000000
0!
1"
0%
1&
b0 *
0.
1/
03
b0 7
#2730000000
1!
1%
1+
1.
10
11
12
13
#2740000000
0!
0%
b1 *
0.
03
b1 7
#2750000000
1!
1%
1.
13
#2760000000
0!
0%
b10 *
0.
03
b10 7
#2770000000
1!
1%
1.
13
#2780000000
0!
0%
b11 *
0.
03
b11 7
#2790000000
1!
1%
1.
13
16
#2800000000
0!
0%
b100 *
0.
03
b100 7
#2810000000
1!
1%
1.
13
#2820000000
0!
0%
b101 *
0.
03
b101 7
#2830000000
1!
1%
1.
13
#2840000000
0!
0%
b110 *
0.
03
b110 7
#2850000000
1!
1%
1.
13
#2860000000
0!
0%
b111 *
0.
03
b111 7
#2870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#2880000000
0!
0"
0%
0&
b0 *
0.
0/
03
b0 7
#2890000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#2900000000
0!
0%
b1 *
0.
03
b1 7
#2910000000
1!
1%
1.
13
#2920000000
0!
0%
b10 *
0.
03
b10 7
#2930000000
1!
1%
1.
13
#2940000000
0!
0%
b11 *
0.
03
b11 7
#2950000000
1!
1%
1.
13
16
#2960000000
0!
0%
b100 *
0.
03
b100 7
#2970000000
1!
1%
1.
13
#2980000000
0!
0%
b101 *
0.
03
b101 7
#2990000000
1!
1%
1.
13
#3000000000
0!
0%
b110 *
0.
03
b110 7
#3010000000
1!
1%
1.
13
#3020000000
0!
0%
b111 *
0.
03
b111 7
#3030000000
1!
1%
1.
13
06
#3040000000
0!
0%
b0 *
0.
03
b0 7
#3050000000
1!
1%
1.
13
#3060000000
0!
0%
b1 *
0.
03
b1 7
#3070000000
1!
1%
1.
13
#3080000000
0!
0%
b10 *
0.
03
b10 7
#3090000000
1!
1%
1.
13
#3100000000
0!
0%
b11 *
0.
03
b11 7
#3110000000
1!
1%
1.
13
16
#3120000000
0!
0%
b100 *
0.
03
b100 7
#3130000000
1!
1%
1.
13
#3140000000
0!
0%
b101 *
0.
03
b101 7
#3150000000
1!
1%
1.
13
#3160000000
0!
0%
b110 *
0.
03
b110 7
#3170000000
1!
1%
1.
13
#3180000000
0!
0%
b111 *
0.
03
b111 7
#3190000000
1!
1%
1.
13
06
#3200000000
0!
0%
b0 *
0.
03
b0 7
#3210000000
1!
1%
1.
13
#3220000000
0!
0%
b1 *
0.
03
b1 7
#3230000000
1!
1%
1.
13
#3240000000
0!
0%
b10 *
0.
03
b10 7
#3250000000
1!
1%
1.
13
#3260000000
0!
0%
b11 *
0.
03
b11 7
#3270000000
1!
1%
1.
13
16
#3280000000
0!
0%
b100 *
0.
03
b100 7
#3290000000
1!
1%
1.
13
#3300000000
0!
0%
b101 *
0.
03
b101 7
#3310000000
1!
1%
1.
13
#3320000000
0!
0%
b110 *
0.
03
b110 7
#3330000000
1!
1%
1.
13
#3340000000
0!
0%
b111 *
0.
03
b111 7
#3350000000
1!
1%
1.
13
06
#3360000000
0!
0%
b0 *
0.
03
b0 7
#3370000000
1!
1%
1.
13
#3380000000
0!
0%
b1 *
0.
03
b1 7
#3390000000
1!
1%
1.
13
#3400000000
0!
1"
0%
1&
b10 *
0.
1/
03
b10 7
#3410000000
1!
1%
1+
1.
10
11
12
13
#3420000000
0!
0%
b11 *
0.
03
b11 7
#3430000000
1!
1%
1.
13
16
#3440000000
0!
0%
b100 *
0.
03
b100 7
#3450000000
1!
1%
1.
13
#3460000000
0!
0%
b101 *
0.
03
b101 7
#3470000000
1!
1%
1.
13
#3480000000
0!
0%
b110 *
0.
03
b110 7
#3490000000
1!
1%
1.
13
#3500000000
0!
0%
b111 *
0.
03
b111 7
#3510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#3520000000
0!
0%
b0 *
0.
03
b0 7
#3530000000
1!
1%
1.
13
#3540000000
0!
0%
b1 *
0.
03
b1 7
#3550000000
1!
1%
1.
13
#3560000000
0!
0"
0%
0&
b10 *
0.
0/
03
b10 7
#3570000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#3580000000
0!
0%
b11 *
0.
03
b11 7
#3590000000
1!
1%
1.
13
16
#3600000000
0!
0%
b100 *
0.
03
b100 7
#3610000000
1!
1%
1.
13
#3620000000
0!
0%
b101 *
0.
03
b101 7
#3630000000
1!
1%
1.
13
#3640000000
0!
0%
b110 *
0.
03
b110 7
#3650000000
1!
1%
1.
13
#3660000000
0!
0%
b111 *
0.
03
b111 7
#3670000000
1!
1%
1.
13
06
#3680000000
0!
0%
b0 *
0.
03
b0 7
#3690000000
1!
1%
1.
13
#3700000000
0!
0%
b1 *
0.
03
b1 7
#3710000000
1!
1%
1.
13
#3720000000
0!
0%
b10 *
0.
03
b10 7
#3730000000
1!
1%
1.
13
#3740000000
0!
0%
b11 *
0.
03
b11 7
#3750000000
1!
1%
1.
13
16
#3760000000
0!
0%
b100 *
0.
03
b100 7
#3770000000
1!
1%
1.
13
#3780000000
0!
0%
b101 *
0.
03
b101 7
#3790000000
1!
1%
1.
13
#3800000000
0!
0%
b110 *
0.
03
b110 7
#3810000000
1!
1%
1.
13
#3820000000
0!
0%
b111 *
0.
03
b111 7
#3830000000
1!
1%
1.
13
06
#3840000000
0!
0%
b0 *
0.
03
b0 7
#3850000000
1!
1%
1.
13
#3860000000
0!
0%
b1 *
0.
03
b1 7
#3870000000
1!
1%
1.
13
#3880000000
0!
0%
b10 *
0.
03
b10 7
#3890000000
1!
1%
1.
13
#3900000000
0!
0%
b11 *
0.
03
b11 7
#3910000000
1!
1%
1.
13
16
#3920000000
0!
0%
b100 *
0.
03
b100 7
#3930000000
1!
1%
1.
13
#3940000000
0!
0%
b101 *
0.
03
b101 7
#3950000000
1!
1%
1.
13
#3960000000
0!
0%
b110 *
0.
03
b110 7
#3970000000
1!
1%
1.
13
#3980000000
0!
0%
b111 *
0.
03
b111 7
#3990000000
1!
1%
1.
13
06
#4000000000
0!
0%
b0 *
0.
03
b0 7
#4010000000
1!
1%
1.
13
#4020000000
0!
0%
b1 *
0.
03
b1 7
#4030000000
1!
1%
1.
13
#4040000000
0!
0%
b10 *
0.
03
b10 7
#4050000000
1!
1%
1.
13
#4060000000
0!
0%
b11 *
0.
03
b11 7
#4070000000
1!
1%
1.
13
16
#4080000000
0!
1"
0%
1&
b100 *
0.
1/
03
b100 7
#4090000000
1!
1%
1+
1.
10
11
12
13
#4100000000
0!
0%
b101 *
0.
03
b101 7
#4110000000
1!
1%
1.
13
#4120000000
0!
0%
b110 *
0.
03
b110 7
#4130000000
1!
1%
1.
13
#4140000000
0!
0%
b111 *
0.
03
b111 7
#4150000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#4160000000
0!
0%
b0 *
0.
03
b0 7
#4170000000
1!
1%
1.
13
#4180000000
0!
0%
b1 *
0.
03
b1 7
#4190000000
1!
1%
1.
13
#4200000000
0!
0%
b10 *
0.
03
b10 7
#4210000000
1!
1%
1.
13
#4220000000
0!
0%
b11 *
0.
03
b11 7
#4230000000
1!
1%
1.
13
16
#4240000000
0!
0"
0%
0&
b100 *
0.
0/
03
b100 7
#4250000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#4260000000
0!
0%
b101 *
0.
03
b101 7
#4270000000
1!
1%
1.
13
#4280000000
0!
0%
b110 *
0.
03
b110 7
#4290000000
1!
1%
1.
13
#4300000000
0!
0%
b111 *
0.
03
b111 7
#4310000000
1!
1%
1.
13
06
#4320000000
0!
0%
b0 *
0.
03
b0 7
#4330000000
1!
1%
1.
13
#4340000000
0!
0%
b1 *
0.
03
b1 7
#4350000000
1!
1%
1.
13
#4360000000
0!
0%
b10 *
0.
03
b10 7
#4370000000
1!
1%
1.
13
#4380000000
0!
0%
b11 *
0.
03
b11 7
#4390000000
1!
1%
1.
13
16
#4400000000
0!
0%
b100 *
0.
03
b100 7
#4410000000
1!
1%
1.
13
#4420000000
0!
0%
b101 *
0.
03
b101 7
#4430000000
1!
1%
1.
13
#4440000000
0!
0%
b110 *
0.
03
b110 7
#4450000000
1!
1%
1.
13
#4460000000
0!
0%
b111 *
0.
03
b111 7
#4470000000
1!
1%
1.
13
06
#4480000000
0!
0%
b0 *
0.
03
b0 7
#4490000000
1!
1%
1.
13
#4500000000
0!
0%
b1 *
0.
03
b1 7
#4510000000
1!
1%
1.
13
#4520000000
0!
0%
b10 *
0.
03
b10 7
#4530000000
1!
1%
1.
13
#4540000000
0!
0%
b11 *
0.
03
b11 7
#4550000000
1!
1%
1.
13
16
#4560000000
0!
0%
b100 *
0.
03
b100 7
#4570000000
1!
1%
1.
13
#4580000000
0!
0%
b101 *
0.
03
b101 7
#4590000000
1!
1%
1.
13
#4600000000
0!
0%
b110 *
0.
03
b110 7
#4610000000
1!
1%
1.
13
#4620000000
0!
0%
b111 *
0.
03
b111 7
#4630000000
1!
1%
1.
13
06
#4640000000
0!
0%
b0 *
0.
03
b0 7
#4650000000
1!
1%
1.
13
#4660000000
0!
0%
b1 *
0.
03
b1 7
#4670000000
1!
1%
1.
13
#4680000000
0!
0%
b10 *
0.
03
b10 7
#4690000000
1!
1%
1.
13
#4700000000
0!
0%
b11 *
0.
03
b11 7
#4710000000
1!
1%
1.
13
16
#4720000000
0!
0%
b100 *
0.
03
b100 7
#4730000000
1!
1%
1.
13
#4740000000
0!
0%
b101 *
0.
03
b101 7
#4750000000
1!
1%
1.
13
#4760000000
0!
1"
0%
1&
b110 *
0.
1/
03
b110 7
#4770000000
1!
1%
1+
1.
10
11
12
13
#4780000000
0!
0%
b111 *
0.
03
b111 7
#4790000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#4800000000
0!
0%
b0 *
0.
03
b0 7
#4810000000
1!
1%
1.
13
#4820000000
0!
0%
b1 *
0.
03
b1 7
#4830000000
1!
1%
1.
13
#4840000000
0!
0%
b10 *
0.
03
b10 7
#4850000000
1!
1%
1.
13
#4860000000
0!
0%
b11 *
0.
03
b11 7
#4870000000
1!
1%
1.
13
16
#4880000000
0!
0%
b100 *
0.
03
b100 7
#4890000000
1!
1%
1.
13
#4900000000
0!
0%
b101 *
0.
03
b101 7
#4910000000
1!
1%
1.
13
#4920000000
0!
0"
0%
0&
b110 *
0.
0/
03
b110 7
#4930000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#4940000000
0!
0%
b111 *
0.
03
b111 7
#4950000000
1!
1%
1.
13
06
#4960000000
0!
0%
b0 *
0.
03
b0 7
#4970000000
1!
1%
1.
13
#4980000000
0!
0%
b1 *
0.
03
b1 7
#4990000000
1!
1%
1.
13
#5000000000
0!
0%
b10 *
0.
03
b10 7
#5010000000
1!
1%
1.
13
#5020000000
0!
0%
b11 *
0.
03
b11 7
#5030000000
1!
1%
1.
13
16
#5040000000
0!
0%
b100 *
0.
03
b100 7
#5050000000
1!
1%
1.
13
#5060000000
0!
0%
b101 *
0.
03
b101 7
#5070000000
1!
1%
1.
13
#5080000000
0!
0%
b110 *
0.
03
b110 7
#5090000000
1!
1%
1.
13
#5100000000
0!
0%
b111 *
0.
03
b111 7
#5110000000
1!
1%
1.
13
06
#5120000000
0!
0%
b0 *
0.
03
b0 7
#5130000000
1!
1%
1.
13
#5140000000
0!
0%
b1 *
0.
03
b1 7
#5150000000
1!
1%
1.
13
#5160000000
0!
0%
b10 *
0.
03
b10 7
#5170000000
1!
1%
1.
13
#5180000000
0!
0%
b11 *
0.
03
b11 7
#5190000000
1!
1%
1.
13
16
#5200000000
0!
0%
b100 *
0.
03
b100 7
#5210000000
1!
1%
1.
13
#5220000000
0!
0%
b101 *
0.
03
b101 7
#5230000000
1!
1%
1.
13
#5240000000
0!
0%
b110 *
0.
03
b110 7
#5250000000
1!
1%
1.
13
#5260000000
0!
0%
b111 *
0.
03
b111 7
#5270000000
1!
1%
1.
13
06
#5280000000
0!
0%
b0 *
0.
03
b0 7
#5290000000
1!
1%
1.
13
#5300000000
0!
0%
b1 *
0.
03
b1 7
#5310000000
1!
1%
1.
13
#5320000000
0!
0%
b10 *
0.
03
b10 7
#5330000000
1!
1%
1.
13
#5340000000
0!
0%
b11 *
0.
03
b11 7
#5350000000
1!
1%
1.
13
16
#5360000000
0!
0%
b100 *
0.
03
b100 7
#5370000000
1!
1%
1.
13
#5380000000
0!
0%
b101 *
0.
03
b101 7
#5390000000
1!
1%
1.
13
#5400000000
0!
0%
b110 *
0.
03
b110 7
#5410000000
1!
1%
1.
13
#5420000000
0!
0%
b111 *
0.
03
b111 7
#5430000000
1!
1%
1.
13
06
#5440000000
0!
1"
0%
1&
b0 *
0.
1/
03
b0 7
#5450000000
1!
1%
1+
1.
10
11
12
13
#5460000000
0!
0%
b1 *
0.
03
b1 7
#5470000000
1!
1%
1.
13
#5480000000
0!
0%
b10 *
0.
03
b10 7
#5490000000
1!
1%
1.
13
#5500000000
0!
0%
b11 *
0.
03
b11 7
#5510000000
1!
1%
1.
13
16
#5520000000
0!
0%
b100 *
0.
03
b100 7
#5530000000
1!
1%
1.
13
#5540000000
0!
0%
b101 *
0.
03
b101 7
#5550000000
1!
1%
1.
13
#5560000000
0!
0%
b110 *
0.
03
b110 7
#5570000000
1!
1%
1.
13
#5580000000
0!
0%
b111 *
0.
03
b111 7
#5590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#5600000000
0!
0"
0%
0&
b0 *
0.
0/
03
b0 7
#5610000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#5620000000
0!
0%
b1 *
0.
03
b1 7
#5630000000
1!
1%
1.
13
#5640000000
0!
0%
b10 *
0.
03
b10 7
#5650000000
1!
1%
1.
13
#5660000000
0!
0%
b11 *
0.
03
b11 7
#5670000000
1!
1%
1.
13
16
#5680000000
0!
0%
b100 *
0.
03
b100 7
#5690000000
1!
1%
1.
13
#5700000000
0!
0%
b101 *
0.
03
b101 7
#5710000000
1!
1%
1.
13
#5720000000
0!
0%
b110 *
0.
03
b110 7
#5730000000
1!
1%
1.
13
#5740000000
0!
0%
b111 *
0.
03
b111 7
#5750000000
1!
1%
1.
13
06
#5760000000
0!
0%
b0 *
0.
03
b0 7
#5770000000
1!
1%
1.
13
#5780000000
0!
0%
b1 *
0.
03
b1 7
#5790000000
1!
1%
1.
13
#5800000000
0!
0%
b10 *
0.
03
b10 7
#5810000000
1!
1%
1.
13
#5820000000
0!
0%
b11 *
0.
03
b11 7
#5830000000
1!
1%
1.
13
16
#5840000000
0!
0%
b100 *
0.
03
b100 7
#5850000000
1!
1%
1.
13
#5860000000
0!
0%
b101 *
0.
03
b101 7
#5870000000
1!
1%
1.
13
#5880000000
0!
0%
b110 *
0.
03
b110 7
#5890000000
1!
1%
1.
13
#5900000000
0!
0%
b111 *
0.
03
b111 7
#5910000000
1!
1%
1.
13
06
#5920000000
0!
0%
b0 *
0.
03
b0 7
#5930000000
1!
1%
1.
13
#5940000000
0!
0%
b1 *
0.
03
b1 7
#5950000000
1!
1%
1.
13
#5960000000
0!
0%
b10 *
0.
03
b10 7
#5970000000
1!
1%
1.
13
#5980000000
0!
0%
b11 *
0.
03
b11 7
#5990000000
1!
1%
1.
13
16
#6000000000
0!
0%
b100 *
0.
03
b100 7
#6010000000
1!
1%
1.
13
#6020000000
0!
0%
b101 *
0.
03
b101 7
#6030000000
1!
1%
1.
13
#6040000000
0!
0%
b110 *
0.
03
b110 7
#6050000000
1!
1%
1.
13
#6060000000
0!
0%
b111 *
0.
03
b111 7
#6070000000
1!
1%
1.
13
06
#6080000000
0!
0%
b0 *
0.
03
b0 7
#6090000000
1!
1%
1.
13
#6100000000
0!
0%
b1 *
0.
03
b1 7
#6110000000
1!
1%
1.
13
#6120000000
0!
1"
0%
1&
b10 *
0.
1/
03
b10 7
#6130000000
1!
1%
1+
1.
10
11
12
13
#6140000000
0!
0%
b11 *
0.
03
b11 7
#6150000000
1!
1%
1.
13
16
#6160000000
0!
0%
b100 *
0.
03
b100 7
#6170000000
1!
1%
1.
13
#6180000000
0!
0%
b101 *
0.
03
b101 7
#6190000000
1!
1%
1.
13
#6200000000
0!
0%
b110 *
0.
03
b110 7
#6210000000
1!
1%
1.
13
#6220000000
0!
0%
b111 *
0.
03
b111 7
#6230000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#6240000000
0!
0%
b0 *
0.
03
b0 7
#6250000000
1!
1%
1.
13
#6260000000
0!
0%
b1 *
0.
03
b1 7
#6270000000
1!
1%
1.
13
#6280000000
0!
0"
0%
0&
b10 *
0.
0/
03
b10 7
#6290000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#6300000000
0!
0%
b11 *
0.
03
b11 7
#6310000000
1!
1%
1.
13
16
#6320000000
0!
0%
b100 *
0.
03
b100 7
#6330000000
1!
1%
1.
13
#6340000000
0!
0%
b101 *
0.
03
b101 7
#6350000000
1!
1%
1.
13
#6360000000
0!
0%
b110 *
0.
03
b110 7
#6370000000
1!
1%
1.
13
#6380000000
0!
0%
b111 *
0.
03
b111 7
#6390000000
1!
1%
1.
13
06
#6400000000
0!
0%
b0 *
0.
03
b0 7
#6410000000
1!
1%
1.
13
#6420000000
0!
0%
b1 *
0.
03
b1 7
#6430000000
1!
1%
1.
13
#6440000000
0!
0%
b10 *
0.
03
b10 7
#6450000000
1!
1%
1.
13
#6460000000
0!
0%
b11 *
0.
03
b11 7
#6470000000
1!
1%
1.
13
16
#6480000000
0!
0%
b100 *
0.
03
b100 7
#6490000000
1!
1%
1.
13
#6500000000
0!
0%
b101 *
0.
03
b101 7
#6510000000
1!
1%
1.
13
#6520000000
0!
0%
b110 *
0.
03
b110 7
#6530000000
1!
1%
1.
13
#6540000000
0!
0%
b111 *
0.
03
b111 7
#6550000000
1!
1%
1.
13
06
#6560000000
0!
0%
b0 *
0.
03
b0 7
#6570000000
1!
1%
1.
13
#6580000000
0!
0%
b1 *
0.
03
b1 7
#6590000000
1!
1%
1.
13
#6600000000
0!
0%
b10 *
0.
03
b10 7
#6610000000
1!
1%
1.
13
#6620000000
0!
0%
b11 *
0.
03
b11 7
#6630000000
1!
1%
1.
13
16
#6640000000
0!
0%
b100 *
0.
03
b100 7
#6650000000
1!
1%
1.
13
#6660000000
0!
0%
b101 *
0.
03
b101 7
#6670000000
1!
1%
1.
13
#6680000000
0!
0%
b110 *
0.
03
b110 7
#6690000000
1!
1%
1.
13
#6700000000
0!
0%
b111 *
0.
03
b111 7
#6710000000
1!
1%
1.
13
06
#6720000000
0!
0%
b0 *
0.
03
b0 7
#6730000000
1!
1%
1.
13
#6740000000
0!
0%
b1 *
0.
03
b1 7
#6750000000
1!
1%
1.
13
#6760000000
0!
0%
b10 *
0.
03
b10 7
#6770000000
1!
1%
1.
13
#6780000000
0!
0%
b11 *
0.
03
b11 7
#6790000000
1!
1%
1.
13
16
#6800000000
0!
1"
0%
1&
b100 *
0.
1/
03
b100 7
#6810000000
1!
1%
1+
1.
10
11
12
13
#6820000000
0!
0%
b101 *
0.
03
b101 7
#6830000000
1!
1%
1.
13
#6840000000
0!
0%
b110 *
0.
03
b110 7
#6850000000
1!
1%
1.
13
#6860000000
0!
0%
b111 *
0.
03
b111 7
#6870000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#6880000000
0!
0%
b0 *
0.
03
b0 7
#6890000000
1!
1%
1.
13
#6900000000
0!
0%
b1 *
0.
03
b1 7
#6910000000
1!
1%
1.
13
#6920000000
0!
0%
b10 *
0.
03
b10 7
#6930000000
1!
1%
1.
13
#6940000000
0!
0%
b11 *
0.
03
b11 7
#6950000000
1!
1%
1.
13
16
#6960000000
0!
0"
0%
0&
b100 *
0.
0/
03
b100 7
#6970000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#6980000000
0!
0%
b101 *
0.
03
b101 7
#6990000000
1!
1%
1.
13
#7000000000
0!
0%
b110 *
0.
03
b110 7
#7010000000
1!
1%
1.
13
#7020000000
0!
0%
b111 *
0.
03
b111 7
#7030000000
1!
1%
1.
13
06
#7040000000
0!
0%
b0 *
0.
03
b0 7
#7050000000
1!
1%
1.
13
#7060000000
0!
0%
b1 *
0.
03
b1 7
#7070000000
1!
1%
1.
13
#7080000000
0!
0%
b10 *
0.
03
b10 7
#7090000000
1!
1%
1.
13
#7100000000
0!
0%
b11 *
0.
03
b11 7
#7110000000
1!
1%
1.
13
16
#7120000000
0!
0%
b100 *
0.
03
b100 7
#7130000000
1!
1%
1.
13
#7140000000
0!
0%
b101 *
0.
03
b101 7
#7150000000
1!
1%
1.
13
#7160000000
0!
0%
b110 *
0.
03
b110 7
#7170000000
1!
1%
1.
13
#7180000000
0!
0%
b111 *
0.
03
b111 7
#7190000000
1!
1%
1.
13
06
#7200000000
0!
0%
b0 *
0.
03
b0 7
#7210000000
1!
1%
1.
13
#7220000000
0!
0%
b1 *
0.
03
b1 7
#7230000000
1!
1%
1.
13
#7240000000
0!
0%
b10 *
0.
03
b10 7
#7250000000
1!
1%
1.
13
#7260000000
0!
0%
b11 *
0.
03
b11 7
#7270000000
1!
1%
1.
13
16
#7280000000
0!
0%
b100 *
0.
03
b100 7
#7290000000
1!
1%
1.
13
#7300000000
0!
0%
b101 *
0.
03
b101 7
#7310000000
1!
1%
1.
13
#7320000000
0!
0%
b110 *
0.
03
b110 7
#7330000000
1!
1%
1.
13
#7340000000
0!
0%
b111 *
0.
03
b111 7
#7350000000
1!
1%
1.
13
06
#7360000000
0!
0%
b0 *
0.
03
b0 7
#7370000000
1!
1%
1.
13
#7380000000
0!
0%
b1 *
0.
03
b1 7
#7390000000
1!
1%
1.
13
#7400000000
0!
0%
b10 *
0.
03
b10 7
#7410000000
1!
1%
1.
13
#7420000000
0!
0%
b11 *
0.
03
b11 7
#7430000000
1!
1%
1.
13
16
#7440000000
0!
0%
b100 *
0.
03
b100 7
#7450000000
1!
1%
1.
13
#7460000000
0!
0%
b101 *
0.
03
b101 7
#7470000000
1!
1%
1.
13
#7480000000
0!
1"
0%
1&
b110 *
0.
1/
03
b110 7
#7490000000
1!
1%
1+
1.
10
11
12
13
#7500000000
0!
0%
b111 *
0.
03
b111 7
#7510000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#7520000000
0!
0%
b0 *
0.
03
b0 7
#7530000000
1!
1%
1.
13
#7540000000
0!
0%
b1 *
0.
03
b1 7
#7550000000
1!
1%
1.
13
#7560000000
0!
0%
b10 *
0.
03
b10 7
#7570000000
1!
1%
1.
13
#7580000000
0!
0%
b11 *
0.
03
b11 7
#7590000000
1!
1%
1.
13
16
#7600000000
0!
0%
b100 *
0.
03
b100 7
#7610000000
1!
1%
1.
13
#7620000000
0!
0%
b101 *
0.
03
b101 7
#7630000000
1!
1%
1.
13
#7640000000
0!
0"
0%
0&
b110 *
0.
0/
03
b110 7
#7650000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#7660000000
0!
0%
b111 *
0.
03
b111 7
#7670000000
1!
1%
1.
13
06
#7680000000
0!
0%
b0 *
0.
03
b0 7
#7690000000
1!
1%
1.
13
#7700000000
0!
0%
b1 *
0.
03
b1 7
#7710000000
1!
1%
1.
13
#7720000000
0!
0%
b10 *
0.
03
b10 7
#7730000000
1!
1%
1.
13
#7740000000
0!
0%
b11 *
0.
03
b11 7
#7750000000
1!
1%
1.
13
16
#7760000000
0!
0%
b100 *
0.
03
b100 7
#7770000000
1!
1%
1.
13
#7780000000
0!
0%
b101 *
0.
03
b101 7
#7790000000
1!
1%
1.
13
#7800000000
0!
0%
b110 *
0.
03
b110 7
#7810000000
1!
1%
1.
13
#7820000000
0!
0%
b111 *
0.
03
b111 7
#7830000000
1!
1%
1.
13
06
#7840000000
0!
0%
b0 *
0.
03
b0 7
#7850000000
1!
1%
1.
13
#7860000000
0!
0%
b1 *
0.
03
b1 7
#7870000000
1!
1%
1.
13
#7880000000
0!
0%
b10 *
0.
03
b10 7
#7890000000
1!
1%
1.
13
#7900000000
0!
0%
b11 *
0.
03
b11 7
#7910000000
1!
1%
1.
13
16
#7920000000
0!
0%
b100 *
0.
03
b100 7
#7930000000
1!
1%
1.
13
#7940000000
0!
0%
b101 *
0.
03
b101 7
#7950000000
1!
1%
1.
13
#7960000000
0!
0%
b110 *
0.
03
b110 7
#7970000000
1!
1%
1.
13
#7980000000
0!
0%
b111 *
0.
03
b111 7
#7990000000
1!
1%
1.
13
06
#8000000000
0!
0%
b0 *
0.
03
b0 7
#8010000000
1!
1%
1.
13
#8020000000
0!
0%
b1 *
0.
03
b1 7
#8030000000
1!
1%
1.
13
#8040000000
0!
0%
b10 *
0.
03
b10 7
#8050000000
1!
1%
1.
13
#8060000000
0!
0%
b11 *
0.
03
b11 7
#8070000000
1!
1%
1.
13
16
#8080000000
0!
0%
b100 *
0.
03
b100 7
#8090000000
1!
1%
1.
13
#8100000000
0!
0%
b101 *
0.
03
b101 7
#8110000000
1!
1%
1.
13
#8120000000
0!
0%
b110 *
0.
03
b110 7
#8130000000
1!
1%
1.
13
#8140000000
0!
0%
b111 *
0.
03
b111 7
#8150000000
1!
1%
1.
13
06
#8160000000
0!
1"
0%
1&
b0 *
0.
1/
03
b0 7
#8170000000
1!
1%
1+
1.
10
11
12
13
#8180000000
0!
0%
b1 *
0.
03
b1 7
#8190000000
1!
1%
1.
13
#8200000000
0!
0%
b10 *
0.
03
b10 7
#8210000000
1!
1%
1.
13
#8220000000
0!
0%
b11 *
0.
03
b11 7
#8230000000
1!
1%
1.
13
16
#8240000000
0!
0%
b100 *
0.
03
b100 7
#8250000000
1!
1%
1.
13
#8260000000
0!
0%
b101 *
0.
03
b101 7
#8270000000
1!
1%
1.
13
#8280000000
0!
0%
b110 *
0.
03
b110 7
#8290000000
1!
1%
1.
13
#8300000000
0!
0%
b111 *
0.
03
b111 7
#8310000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#8320000000
0!
0"
0%
0&
b0 *
0.
0/
03
b0 7
#8330000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#8340000000
0!
0%
b1 *
0.
03
b1 7
#8350000000
1!
1%
1.
13
#8360000000
0!
0%
b10 *
0.
03
b10 7
#8370000000
1!
1%
1.
13
#8380000000
0!
0%
b11 *
0.
03
b11 7
#8390000000
1!
1%
1.
13
16
#8400000000
0!
0%
b100 *
0.
03
b100 7
#8410000000
1!
1%
1.
13
#8420000000
0!
0%
b101 *
0.
03
b101 7
#8430000000
1!
1%
1.
13
#8440000000
0!
0%
b110 *
0.
03
b110 7
#8450000000
1!
1%
1.
13
#8460000000
0!
0%
b111 *
0.
03
b111 7
#8470000000
1!
1%
1.
13
06
#8480000000
0!
0%
b0 *
0.
03
b0 7
#8490000000
1!
1%
1.
13
#8500000000
0!
0%
b1 *
0.
03
b1 7
#8510000000
1!
1%
1.
13
#8520000000
0!
0%
b10 *
0.
03
b10 7
#8530000000
1!
1%
1.
13
#8540000000
0!
0%
b11 *
0.
03
b11 7
#8550000000
1!
1%
1.
13
16
#8560000000
0!
0%
b100 *
0.
03
b100 7
#8570000000
1!
1%
1.
13
#8580000000
0!
0%
b101 *
0.
03
b101 7
#8590000000
1!
1%
1.
13
#8600000000
0!
0%
b110 *
0.
03
b110 7
#8610000000
1!
1%
1.
13
#8620000000
0!
0%
b111 *
0.
03
b111 7
#8630000000
1!
1%
1.
13
06
#8640000000
0!
0%
b0 *
0.
03
b0 7
#8650000000
1!
1%
1.
13
#8660000000
0!
0%
b1 *
0.
03
b1 7
#8670000000
1!
1%
1.
13
#8680000000
0!
0%
b10 *
0.
03
b10 7
#8690000000
1!
1%
1.
13
#8700000000
0!
0%
b11 *
0.
03
b11 7
#8710000000
1!
1%
1.
13
16
#8720000000
0!
0%
b100 *
0.
03
b100 7
#8730000000
1!
1%
1.
13
#8740000000
0!
0%
b101 *
0.
03
b101 7
#8750000000
1!
1%
1.
13
#8760000000
0!
0%
b110 *
0.
03
b110 7
#8770000000
1!
1%
1.
13
#8780000000
0!
0%
b111 *
0.
03
b111 7
#8790000000
1!
1%
1.
13
06
#8800000000
0!
0%
b0 *
0.
03
b0 7
#8810000000
1!
1%
1.
13
#8820000000
0!
0%
b1 *
0.
03
b1 7
#8830000000
1!
1%
1.
13
#8840000000
0!
1"
0%
1&
b10 *
0.
1/
03
b10 7
#8850000000
1!
1%
1+
1.
10
11
12
13
#8860000000
0!
0%
b11 *
0.
03
b11 7
#8870000000
1!
1%
1.
13
16
#8880000000
0!
0%
b100 *
0.
03
b100 7
#8890000000
1!
1%
1.
13
#8900000000
0!
0%
b101 *
0.
03
b101 7
#8910000000
1!
1%
1.
13
#8920000000
0!
0%
b110 *
0.
03
b110 7
#8930000000
1!
1%
1.
13
#8940000000
0!
0%
b111 *
0.
03
b111 7
#8950000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#8960000000
0!
0%
b0 *
0.
03
b0 7
#8970000000
1!
1%
1.
13
#8980000000
0!
0%
b1 *
0.
03
b1 7
#8990000000
1!
1%
1.
13
#9000000000
0!
0"
0%
0&
b10 *
0.
0/
03
b10 7
#9010000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#9020000000
0!
0%
b11 *
0.
03
b11 7
#9030000000
1!
1%
1.
13
16
#9040000000
0!
0%
b100 *
0.
03
b100 7
#9050000000
1!
1%
1.
13
#9060000000
0!
0%
b101 *
0.
03
b101 7
#9070000000
1!
1%
1.
13
#9080000000
0!
0%
b110 *
0.
03
b110 7
#9090000000
1!
1%
1.
13
#9100000000
0!
0%
b111 *
0.
03
b111 7
#9110000000
1!
1%
1.
13
06
#9120000000
0!
0%
b0 *
0.
03
b0 7
#9130000000
1!
1%
1.
13
#9140000000
0!
0%
b1 *
0.
03
b1 7
#9150000000
1!
1%
1.
13
#9160000000
0!
0%
b10 *
0.
03
b10 7
#9170000000
1!
1%
1.
13
#9180000000
0!
0%
b11 *
0.
03
b11 7
#9190000000
1!
1%
1.
13
16
#9200000000
0!
0%
b100 *
0.
03
b100 7
#9210000000
1!
1%
1.
13
#9220000000
0!
0%
b101 *
0.
03
b101 7
#9230000000
1!
1%
1.
13
#9240000000
0!
0%
b110 *
0.
03
b110 7
#9250000000
1!
1%
1.
13
#9260000000
0!
0%
b111 *
0.
03
b111 7
#9270000000
1!
1%
1.
13
06
#9280000000
0!
0%
b0 *
0.
03
b0 7
#9290000000
1!
1%
1.
13
#9300000000
0!
0%
b1 *
0.
03
b1 7
#9310000000
1!
1%
1.
13
#9320000000
0!
0%
b10 *
0.
03
b10 7
#9330000000
1!
1%
1.
13
#9340000000
0!
0%
b11 *
0.
03
b11 7
#9350000000
1!
1%
1.
13
16
#9360000000
0!
0%
b100 *
0.
03
b100 7
#9370000000
1!
1%
1.
13
#9380000000
0!
0%
b101 *
0.
03
b101 7
#9390000000
1!
1%
1.
13
#9400000000
0!
0%
b110 *
0.
03
b110 7
#9410000000
1!
1%
1.
13
#9420000000
0!
0%
b111 *
0.
03
b111 7
#9430000000
1!
1%
1.
13
06
#9440000000
0!
0%
b0 *
0.
03
b0 7
#9450000000
1!
1%
1.
13
#9460000000
0!
0%
b1 *
0.
03
b1 7
#9470000000
1!
1%
1.
13
#9480000000
0!
0%
b10 *
0.
03
b10 7
#9490000000
1!
1%
1.
13
#9500000000
0!
0%
b11 *
0.
03
b11 7
#9510000000
1!
1%
1.
13
16
#9520000000
0!
1"
0%
1&
b100 *
0.
1/
03
b100 7
#9530000000
1!
1%
1+
1.
10
11
12
13
#9540000000
0!
0%
b101 *
0.
03
b101 7
#9550000000
1!
1%
1.
13
#9560000000
0!
0%
b110 *
0.
03
b110 7
#9570000000
1!
1%
1.
13
#9580000000
0!
0%
b111 *
0.
03
b111 7
#9590000000
1!
b0100 #
b1101101 $
1%
b0100 '
b1101101 (
b0010 )
1.
13
06
b1101101 8
b0010 9
#9600000000
0!
0%
b0 *
0.
03
b0 7
#9610000000
1!
1%
1.
13
#9620000000
0!
0%
b1 *
0.
03
b1 7
#9630000000
1!
1%
1.
13
#9640000000
0!
0%
b10 *
0.
03
b10 7
#9650000000
1!
1%
1.
13
#9660000000
0!
0%
b11 *
0.
03
b11 7
#9670000000
1!
1%
1.
13
16
#9680000000
0!
0"
0%
0&
b100 *
0.
0/
03
b100 7
#9690000000
1!
b1000 #
b0110000 $
1%
b1000 '
b0110000 (
b0001 )
0+
1.
00
01
02
13
b0110000 8
b0001 9
#9700000000
0!
0%
b101 *
0.
03
b101 7
#9710000000
1!
1%
1.
13
#9720000000
0!
0%
b110 *
0.
03
b110 7
#9730000000
1!
1%
1.
13
#9740000000
0!
0%
b111 *
0.
03
b111 7
#9750000000
1!
1%
1.
13
06
#9760000000
0!
0%
b0 *
0.
03
b0 7
#9770000000
1!
1%
1.
13
#9780000000
0!
0%
b1 *
0.
03
b1 7
#9790000000
1!
1%
1.
13
#9800000000
0!
0%
b10 *
0.
03
b10 7
#9810000000
1!
1%
1.
13
#9820000000
0!
0%
b11 *
0.
03
b11 7
#9830000000
1!
1%
1.
13
16
#9840000000
0!
0%
b100 *
0.
03
b100 7
#9850000000
1!
1%
1.
13
#9860000000
0!
0%
b101 *
0.
03
b101 7
#9870000000
1!
1%
1.
13
#9880000000
0!
0%
b110 *
0.
03
b110 7
#9890000000
1!
1%
1.
13
#9900000000
0!
0%
b111 *
0.
03
b111 7
#9910000000
1!
1%
1.
13
06
#9920000000
0!
0%
b0 *
0.
03
b0 7
#9930000000
1!
1%
1.
13
#9940000000
0!
0%
b1 *
0.
03
b1 7
#9950000000
1!
1%
1.
13
#9960000000
0!
0%
b10 *
0.
03
b10 7
#9970000000
1!
1%
1.
13
#9980000000
0!
0%
b11 *
0.
03
b11 7
#9990000000
1!
1%
1.
13
16
#10000000000
0!
0%
b100 *
0.
03
b100 7
