$date
  Tue May 14 11:25:49 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_motor $end
$var reg 1 ! clk $end
$var reg 1 " key_asc $end
$var reg 1 # key_desc $end
$var reg 1 $ key_frec $end
$var reg 1 % enable_disp $end
$var reg 7 & segmentos[6:0] $end
$var reg 4 ' salida[3:0] $end
$scope module uut $end
$var reg 1 ( clk $end
$var reg 1 ) key_asc $end
$var reg 1 * key_desc $end
$var reg 1 + key_frec $end
$var reg 1 , enable_disp $end
$var reg 7 - segmentos[6:0] $end
$var reg 4 . salida[3:0] $end
$comment state is not handled $end
$var integer 32 / cuenta $end
$var integer 32 0 cuenta_maxima $end
$var integer 32 1 aux $end
$var integer 32 2 cuenta2 $end
$var reg 4 3 bcd_disp[3:0] $end
$scope module a $end
$var reg 1 4 clk $end
$var reg 1 5 reset $end
$var reg 1 6 enable $end
$var reg 1 7 cout $end
$var integer 32 8 q $end
$upscope $end
$scope module a2 $end
$var reg 1 9 clk $end
$var reg 1 : reset $end
$var reg 1 ; enable $end
$var reg 1 < cout $end
$var integer 32 = q $end
$upscope $end
$scope module b $end
$var reg 7 > segmentos[6:0] $end
$var reg 4 ? bcd[3:0] $end
$var reg 1 @ enable $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
0#
U$
0%
b0000001 &
b1000 '
0(
0)
0*
U+
0,
b0000001 -
b1000 .
b0 /
b1010 0
b0 1
b0 2
b0000 3
04
05
16
U7
b0 8
09
0:
1;
U<
b0 =
b0000001 >
b0000 ?
0@
#10000000
1!
1(
14
07
19
1<
#20000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#30000000
1!
1(
b1 1
14
19
0<
#40000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#50000000
1!
1(
b10 1
14
19
1<
#60000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#70000000
1!
1(
b11 1
14
19
0<
#80000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#90000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b100 1
b0001 3
14
17
19
1<
b1001111 >
b0001 ?
#100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#110000000
1!
1(
b101 1
14
19
0<
#120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#130000000
1!
1(
b110 1
14
19
1<
#140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#150000000
1!
1(
b111 1
14
19
0<
#160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#170000000
1!
1(
b1000 1
14
19
1<
#180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#190000000
1!
1(
b1001 1
14
07
19
0<
#200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#210000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
1<
#220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#230000000
1!
1(
b1 1
14
19
0<
#240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#250000000
1!
1(
b10 1
14
19
1<
#260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#270000000
1!
1(
b11 1
14
19
0<
#280000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#290000000
1!
1(
b100 1
14
17
19
1<
#300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#310000000
1!
1(
b101 1
14
19
0<
#320000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#330000000
1!
1(
b110 1
14
19
1<
#340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#350000000
1!
1(
b111 1
14
19
0<
#360000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#370000000
1!
1(
b1000 1
14
19
1<
#380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#390000000
1!
1(
b1001 1
14
07
19
0<
#400000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#410000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
1<
#420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#430000000
1!
1(
b1 1
14
19
0<
#440000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#450000000
1!
1(
b10 1
14
19
1<
#460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#470000000
1!
1(
b11 1
14
19
0<
#480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#490000000
1!
1(
b100 1
14
17
19
1<
#500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#510000000
1!
1(
b101 1
14
19
0<
#520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#530000000
1!
1(
b110 1
14
19
1<
#540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#550000000
1!
1(
b111 1
14
19
0<
#560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#570000000
1!
1(
b1000 1
14
19
1<
#580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#590000000
1!
1(
b1001 1
14
07
19
0<
#600000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b0 /
b0 2
b0000 3
04
b0 8
09
b0 =
b0000001 >
b0000 ?
#610000000
1!
1(
b0 1
14
19
1<
#620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#630000000
1!
1(
b1 1
14
19
0<
#640000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#650000000
1!
1(
b10 1
14
19
1<
#660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#670000000
1!
1(
b11 1
14
19
0<
#680000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#690000000
1!
1(
b100 1
14
17
19
1<
#700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#710000000
1!
1(
b101 1
14
19
0<
#720000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#730000000
1!
1(
b110 1
14
19
1<
#740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#750000000
1!
1(
b111 1
14
19
0<
#760000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#770000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b1000 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#790000000
1!
1(
b1001 1
14
07
19
0<
#800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#810000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
1<
#820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#830000000
1!
1(
b1 1
14
19
0<
#840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#850000000
1!
1(
b10 1
14
19
1<
#860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#870000000
1!
1(
b11 1
14
19
0<
#880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#890000000
1!
1(
b100 1
14
17
19
1<
#900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#910000000
1!
1(
b101 1
14
19
0<
#920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#930000000
1!
1(
b110 1
14
19
1<
#940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#950000000
1!
1(
b111 1
14
19
0<
#960000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#970000000
1!
1(
b1000 1
14
19
1<
#980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#990000000
1!
1(
b1001 1
14
07
19
0<
#1000000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#1010000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
1<
#1020000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#1030000000
1!
1(
b1 1
14
19
0<
#1040000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#1050000000
1!
1(
b10 1
14
19
1<
#1060000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#1070000000
1!
1(
b11 1
14
19
0<
#1080000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#1090000000
1!
1(
b100 1
14
17
19
1<
#1100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#1110000000
1!
1(
b101 1
14
19
0<
#1120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#1130000000
1!
1(
b110 1
14
19
1<
#1140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#1150000000
1!
1(
b111 1
14
19
0<
#1160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#1170000000
1!
1(
b1000 1
14
19
1<
#1180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#1190000000
1!
1(
b1001 1
14
07
19
0<
#1200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#1210000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
1<
#1220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#1230000000
1!
1(
b1 1
14
19
0<
#1240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#1250000000
1!
1(
b10 1
14
19
1<
#1260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#1270000000
1!
1(
b11 1
14
19
0<
#1280000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b100 /
b0 2
b0000 3
04
b100 8
09
b0 =
b0000001 >
b0000 ?
#1290000000
1!
1(
b100 1
14
17
19
1<
#1300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#1310000000
1!
1(
b101 1
14
19
0<
#1320000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#1330000000
1!
1(
b110 1
14
19
1<
#1340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#1350000000
1!
1(
b111 1
14
19
0<
#1360000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#1370000000
1!
1(
b1000 1
14
19
1<
#1380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#1390000000
1!
1(
b1001 1
14
07
19
0<
#1400000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#1410000000
1!
1(
b0 1
14
19
1<
#1420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#1430000000
1!
1(
b1 1
14
19
0<
#1440000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#1450000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b10 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#1460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#1470000000
1!
1(
b11 1
14
19
0<
#1480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#1490000000
1!
1(
b100 1
14
17
19
1<
#1500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#1510000000
1!
1(
b101 1
14
19
0<
#1520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#1530000000
1!
1(
b110 1
14
19
1<
#1540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#1550000000
1!
1(
b111 1
14
19
0<
#1560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#1570000000
1!
1(
b1000 1
14
19
1<
#1580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#1590000000
1!
1(
b1001 1
14
07
19
0<
#1600000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#1610000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
1<
#1620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#1630000000
1!
1(
b1 1
14
19
0<
#1640000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#1650000000
1!
1(
b10 1
14
19
1<
#1660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#1670000000
1!
1(
b11 1
14
19
0<
#1680000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#1690000000
1!
1(
b100 1
14
17
19
1<
#1700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#1710000000
1!
1(
b101 1
14
19
0<
#1720000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#1730000000
1!
1(
b110 1
14
19
1<
#1740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#1750000000
1!
1(
b111 1
14
19
0<
#1760000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#1770000000
1!
1(
b1000 1
14
19
1<
#1780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#1790000000
1!
1(
b1001 1
14
07
19
0<
#1800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#1810000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
1<
#1820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#1830000000
1!
1(
b1 1
14
19
0<
#1840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#1850000000
1!
1(
b10 1
14
19
1<
#1860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#1870000000
1!
1(
b11 1
14
19
0<
#1880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#1890000000
1!
1(
b100 1
14
17
19
1<
#1900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#1910000000
1!
1(
b101 1
14
19
0<
#1920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#1930000000
1!
1(
b110 1
14
19
1<
#1940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#1950000000
1!
1(
b111 1
14
19
0<
#1960000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b1000 /
b0 2
b0000 3
04
b1000 8
09
b0 =
b0000001 >
b0000 ?
#1970000000
1!
1(
b1000 1
14
19
1<
#1980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#1990000000
1!
1(
b1001 1
14
07
19
0<
#2000000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#2010000000
1!
1(
b0 1
14
19
1<
#2020000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#2030000000
1!
1(
b1 1
14
19
0<
#2040000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#2050000000
1!
1(
b10 1
14
19
1<
#2060000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#2070000000
1!
1(
b11 1
14
19
0<
#2080000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#2090000000
1!
1(
b100 1
14
17
19
1<
#2100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#2110000000
1!
1(
b101 1
14
19
0<
#2120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#2130000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b110 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#2140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#2150000000
1!
1(
b111 1
14
19
0<
#2160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#2170000000
1!
1(
b1000 1
14
19
1<
#2180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#2190000000
1!
1(
b1001 1
14
07
19
0<
#2200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#2210000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
1<
#2220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#2230000000
1!
1(
b1 1
14
19
0<
#2240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#2250000000
1!
1(
b10 1
14
19
1<
#2260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#2270000000
1!
1(
b11 1
14
19
0<
#2280000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#2290000000
1!
1(
b100 1
14
17
19
1<
#2300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#2310000000
1!
1(
b101 1
14
19
0<
#2320000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#2330000000
1!
1(
b110 1
14
19
1<
#2340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#2350000000
1!
1(
b111 1
14
19
0<
#2360000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#2370000000
1!
1(
b1000 1
14
19
1<
#2380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#2390000000
1!
1(
b1001 1
14
07
19
0<
#2400000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#2410000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
1<
#2420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#2430000000
1!
1(
b1 1
14
19
0<
#2440000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#2450000000
1!
1(
b10 1
14
19
1<
#2460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#2470000000
1!
1(
b11 1
14
19
0<
#2480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#2490000000
1!
1(
b100 1
14
17
19
1<
#2500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#2510000000
1!
1(
b101 1
14
19
0<
#2520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#2530000000
1!
1(
b110 1
14
19
1<
#2540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#2550000000
1!
1(
b111 1
14
19
0<
#2560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#2570000000
1!
1(
b1000 1
14
19
1<
#2580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#2590000000
1!
1(
b1001 1
14
07
19
0<
#2600000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#2610000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
1<
#2620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#2630000000
1!
1(
b1 1
14
19
0<
#2640000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b10 /
b0 2
b0000 3
04
b10 8
09
b0 =
b0000001 >
b0000 ?
#2650000000
1!
1(
b10 1
14
19
1<
#2660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#2670000000
1!
1(
b11 1
14
19
0<
#2680000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#2690000000
1!
1(
b100 1
14
17
19
1<
#2700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#2710000000
1!
1(
b101 1
14
19
0<
#2720000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#2730000000
1!
1(
b110 1
14
19
1<
#2740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#2750000000
1!
1(
b111 1
14
19
0<
#2760000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#2770000000
1!
1(
b1000 1
14
19
1<
#2780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#2790000000
1!
1(
b1001 1
14
07
19
0<
#2800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#2810000000
1!
1"
b1001111 &
b0110 '
1(
1)
b1001111 -
b0110 .
b0 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#2820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#2830000000
1!
1(
b1 1
14
19
0<
#2840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#2850000000
1!
1(
b10 1
14
19
1<
#2860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#2870000000
1!
1(
b11 1
14
19
0<
#2880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#2890000000
1!
1(
b100 1
14
17
19
1<
#2900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#2910000000
1!
1(
b101 1
14
19
0<
#2920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#2930000000
1!
1(
b110 1
14
19
1<
#2940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#2950000000
1!
1(
b111 1
14
19
0<
#2960000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#2970000000
1!
1(
b1000 1
14
19
1<
#2980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#2990000000
1!
1(
b1001 1
14
07
19
0<
#3000000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#3010000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
1<
#3020000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#3030000000
1!
1(
b1 1
14
19
0<
#3040000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#3050000000
1!
1(
b10 1
14
19
1<
#3060000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#3070000000
1!
1(
b11 1
14
19
0<
#3080000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#3090000000
1!
1(
b100 1
14
17
19
1<
#3100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#3110000000
1!
1(
b101 1
14
19
0<
#3120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#3130000000
1!
1(
b110 1
14
19
1<
#3140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#3150000000
1!
1(
b111 1
14
19
0<
#3160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#3170000000
1!
1(
b1000 1
14
19
1<
#3180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#3190000000
1!
1(
b1001 1
14
07
19
0<
#3200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#3210000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
1<
#3220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#3230000000
1!
1(
b1 1
14
19
0<
#3240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#3250000000
1!
1(
b10 1
14
19
1<
#3260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#3270000000
1!
1(
b11 1
14
19
0<
#3280000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#3290000000
1!
1(
b100 1
14
17
19
1<
#3300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#3310000000
1!
1(
b101 1
14
19
0<
#3320000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b110 /
b0 2
b0000 3
04
b110 8
09
b0 =
b0000001 >
b0000 ?
#3330000000
1!
1(
b110 1
14
19
1<
#3340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#3350000000
1!
1(
b111 1
14
19
0<
#3360000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#3370000000
1!
1(
b1000 1
14
19
1<
#3380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#3390000000
1!
1(
b1001 1
14
07
19
0<
#3400000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#3410000000
1!
1(
b0 1
14
19
1<
#3420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#3430000000
1!
1(
b1 1
14
19
0<
#3440000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#3450000000
1!
1(
b10 1
14
19
1<
#3460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#3470000000
1!
1(
b11 1
14
19
0<
#3480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#3490000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b100 1
b0001 3
14
17
19
1<
b1001111 >
b0001 ?
#3500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#3510000000
1!
1(
b101 1
14
19
0<
#3520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#3530000000
1!
1(
b110 1
14
19
1<
#3540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#3550000000
1!
1(
b111 1
14
19
0<
#3560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#3570000000
1!
1(
b1000 1
14
19
1<
#3580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#3590000000
1!
1(
b1001 1
14
07
19
0<
#3600000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#3610000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
1<
#3620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#3630000000
1!
1(
b1 1
14
19
0<
#3640000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#3650000000
1!
1(
b10 1
14
19
1<
#3660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#3670000000
1!
1(
b11 1
14
19
0<
#3680000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#3690000000
1!
1(
b100 1
14
17
19
1<
#3700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#3710000000
1!
1(
b101 1
14
19
0<
#3720000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#3730000000
1!
1(
b110 1
14
19
1<
#3740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#3750000000
1!
1(
b111 1
14
19
0<
#3760000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#3770000000
1!
1(
b1000 1
14
19
1<
#3780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#3790000000
1!
1(
b1001 1
14
07
19
0<
#3800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#3810000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
1<
#3820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#3830000000
1!
1(
b1 1
14
19
0<
#3840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#3850000000
1!
1(
b10 1
14
19
1<
#3860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#3870000000
1!
1(
b11 1
14
19
0<
#3880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#3890000000
1!
1(
b100 1
14
17
19
1<
#3900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#3910000000
1!
1(
b101 1
14
19
0<
#3920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#3930000000
1!
1(
b110 1
14
19
1<
#3940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#3950000000
1!
1(
b111 1
14
19
0<
#3960000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#3970000000
1!
1(
b1000 1
14
19
1<
#3980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#3990000000
1!
1(
b1001 1
14
07
19
0<
#4000000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b0 /
b0 2
b0000 3
04
b0 8
09
b0 =
b0000001 >
b0000 ?
#4010000000
1!
1(
b0 1
14
19
1<
#4020000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#4030000000
1!
1(
b1 1
14
19
0<
#4040000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#4050000000
1!
1(
b10 1
14
19
1<
#4060000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#4070000000
1!
1(
b11 1
14
19
0<
#4080000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#4090000000
1!
1(
b100 1
14
17
19
1<
#4100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#4110000000
1!
1(
b101 1
14
19
0<
#4120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#4130000000
1!
1(
b110 1
14
19
1<
#4140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#4150000000
1!
1(
b111 1
14
19
0<
#4160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#4170000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b1000 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#4180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#4190000000
1!
1(
b1001 1
14
07
19
0<
#4200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#4210000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
1<
#4220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#4230000000
1!
1(
b1 1
14
19
0<
#4240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#4250000000
1!
1(
b10 1
14
19
1<
#4260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#4270000000
1!
1(
b11 1
14
19
0<
#4280000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#4290000000
1!
1(
b100 1
14
17
19
1<
#4300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#4310000000
1!
1(
b101 1
14
19
0<
#4320000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#4330000000
1!
1(
b110 1
14
19
1<
#4340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#4350000000
1!
1(
b111 1
14
19
0<
#4360000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#4370000000
1!
1(
b1000 1
14
19
1<
#4380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#4390000000
1!
1(
b1001 1
14
07
19
0<
#4400000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#4410000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
1<
#4420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#4430000000
1!
1(
b1 1
14
19
0<
#4440000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#4450000000
1!
1(
b10 1
14
19
1<
#4460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#4470000000
1!
1(
b11 1
14
19
0<
#4480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#4490000000
1!
1(
b100 1
14
17
19
1<
#4500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#4510000000
1!
1(
b101 1
14
19
0<
#4520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#4530000000
1!
1(
b110 1
14
19
1<
#4540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#4550000000
1!
1(
b111 1
14
19
0<
#4560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#4570000000
1!
1(
b1000 1
14
19
1<
#4580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#4590000000
1!
1(
b1001 1
14
07
19
0<
#4600000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#4610000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
1<
#4620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#4630000000
1!
1(
b1 1
14
19
0<
#4640000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#4650000000
1!
1(
b10 1
14
19
1<
#4660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#4670000000
1!
1(
b11 1
14
19
0<
#4680000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b100 /
b0 2
b0000 3
04
b100 8
09
b0 =
b0000001 >
b0000 ?
#4690000000
1!
1(
b100 1
14
17
19
1<
#4700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#4710000000
1!
1(
b101 1
14
19
0<
#4720000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#4730000000
1!
1(
b110 1
14
19
1<
#4740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#4750000000
1!
1(
b111 1
14
19
0<
#4760000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#4770000000
1!
1(
b1000 1
14
19
1<
#4780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#4790000000
1!
1(
b1001 1
14
07
19
0<
#4800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#4810000000
1!
1(
b0 1
14
19
1<
#4820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#4830000000
1!
1(
b1 1
14
19
0<
#4840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#4850000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b10 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#4860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#4870000000
1!
1(
b11 1
14
19
0<
#4880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#4890000000
1!
1(
b100 1
14
17
19
1<
#4900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#4910000000
1!
1(
b101 1
14
19
0<
#4920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#4930000000
1!
1(
b110 1
14
19
1<
#4940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#4950000000
1!
1(
b111 1
14
19
0<
#4960000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#4970000000
1!
1(
b1000 1
14
19
1<
#4980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#4990000000
1!
1(
b1001 1
14
07
19
0<
#5000000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#5010000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
1<
#5020000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#5030000000
1!
1(
b1 1
14
19
0<
#5040000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#5050000000
1!
1(
b10 1
14
19
1<
#5060000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#5070000000
1!
1(
b11 1
14
19
0<
#5080000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#5090000000
1!
1(
b100 1
14
17
19
1<
#5100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#5110000000
1!
1(
b101 1
14
19
0<
#5120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#5130000000
1!
1(
b110 1
14
19
1<
#5140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#5150000000
1!
1(
b111 1
14
19
0<
#5160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#5170000000
1!
1(
b1000 1
14
19
1<
#5180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#5190000000
1!
1(
b1001 1
14
07
19
0<
#5200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#5210000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
1<
#5220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#5230000000
1!
1(
b1 1
14
19
0<
#5240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#5250000000
1!
1(
b10 1
14
19
1<
#5260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#5270000000
1!
1(
b11 1
14
19
0<
#5280000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#5290000000
1!
1(
b100 1
14
17
19
1<
#5300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#5310000000
1!
1(
b101 1
14
19
0<
#5320000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#5330000000
1!
1(
b110 1
14
19
1<
#5340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#5350000000
1!
1(
b111 1
14
19
0<
#5360000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b1000 /
b0 2
b0000 3
04
b1000 8
09
b0 =
b0000001 >
b0000 ?
#5370000000
1!
1(
b1000 1
14
19
1<
#5380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#5390000000
1!
1(
b1001 1
14
07
19
0<
#5400000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#5410000000
1!
1(
b0 1
14
19
1<
#5420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#5430000000
1!
1(
b1 1
14
19
0<
#5440000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#5450000000
1!
1(
b10 1
14
19
1<
#5460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#5470000000
1!
1(
b11 1
14
19
0<
#5480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#5490000000
1!
1(
b100 1
14
17
19
1<
#5500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#5510000000
1!
1(
b101 1
14
19
0<
#5520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#5530000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b110 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#5540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#5550000000
1!
1(
b111 1
14
19
0<
#5560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#5570000000
1!
1(
b1000 1
14
19
1<
#5580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#5590000000
1!
1(
b1001 1
14
07
19
0<
#5600000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#5610000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
1<
#5620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#5630000000
1!
1(
b1 1
14
19
0<
#5640000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#5650000000
1!
1(
b10 1
14
19
1<
#5660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#5670000000
1!
1(
b11 1
14
19
0<
#5680000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#5690000000
1!
1(
b100 1
14
17
19
1<
#5700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#5710000000
1!
1(
b101 1
14
19
0<
#5720000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#5730000000
1!
1(
b110 1
14
19
1<
#5740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#5750000000
1!
1(
b111 1
14
19
0<
#5760000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#5770000000
1!
1(
b1000 1
14
19
1<
#5780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#5790000000
1!
1(
b1001 1
14
07
19
0<
#5800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#5810000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
1<
#5820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#5830000000
1!
1(
b1 1
14
19
0<
#5840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#5850000000
1!
1(
b10 1
14
19
1<
#5860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#5870000000
1!
1(
b11 1
14
19
0<
#5880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#5890000000
1!
1(
b100 1
14
17
19
1<
#5900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#5910000000
1!
1(
b101 1
14
19
0<
#5920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#5930000000
1!
1(
b110 1
14
19
1<
#5940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#5950000000
1!
1(
b111 1
14
19
0<
#5960000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#5970000000
1!
1(
b1000 1
14
19
1<
#5980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#5990000000
1!
1(
b1001 1
14
07
19
0<
#6000000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#6010000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
1<
#6020000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#6030000000
1!
1(
b1 1
14
19
0<
#6040000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b10 /
b0 2
b0000 3
04
b10 8
09
b0 =
b0000001 >
b0000 ?
#6050000000
1!
1(
b10 1
14
19
1<
#6060000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#6070000000
1!
1(
b11 1
14
19
0<
#6080000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#6090000000
1!
1(
b100 1
14
17
19
1<
#6100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#6110000000
1!
1(
b101 1
14
19
0<
#6120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#6130000000
1!
1(
b110 1
14
19
1<
#6140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#6150000000
1!
1(
b111 1
14
19
0<
#6160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#6170000000
1!
1(
b1000 1
14
19
1<
#6180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#6190000000
1!
1(
b1001 1
14
07
19
0<
#6200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#6210000000
1!
1"
b1001111 &
b1000 '
1(
1)
b1001111 -
b1000 .
b0 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#6220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#6230000000
1!
1(
b1 1
14
19
0<
#6240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#6250000000
1!
1(
b10 1
14
19
1<
#6260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#6270000000
1!
1(
b11 1
14
19
0<
#6280000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#6290000000
1!
1(
b100 1
14
17
19
1<
#6300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#6310000000
1!
1(
b101 1
14
19
0<
#6320000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#6330000000
1!
1(
b110 1
14
19
1<
#6340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#6350000000
1!
1(
b111 1
14
19
0<
#6360000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#6370000000
1!
1(
b1000 1
14
19
1<
#6380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#6390000000
1!
1(
b1001 1
14
07
19
0<
#6400000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#6410000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
1<
#6420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#6430000000
1!
1(
b1 1
14
19
0<
#6440000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#6450000000
1!
1(
b10 1
14
19
1<
#6460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#6470000000
1!
1(
b11 1
14
19
0<
#6480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#6490000000
1!
1(
b100 1
14
17
19
1<
#6500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#6510000000
1!
1(
b101 1
14
19
0<
#6520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#6530000000
1!
1(
b110 1
14
19
1<
#6540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#6550000000
1!
1(
b111 1
14
19
0<
#6560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#6570000000
1!
1(
b1000 1
14
19
1<
#6580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#6590000000
1!
1(
b1001 1
14
07
19
0<
#6600000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#6610000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
1<
#6620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#6630000000
1!
1(
b1 1
14
19
0<
#6640000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#6650000000
1!
1(
b10 1
14
19
1<
#6660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#6670000000
1!
1(
b11 1
14
19
0<
#6680000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#6690000000
1!
1(
b100 1
14
17
19
1<
#6700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#6710000000
1!
1(
b101 1
14
19
0<
#6720000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b110 /
b0 2
b0000 3
04
b110 8
09
b0 =
b0000001 >
b0000 ?
#6730000000
1!
1(
b110 1
14
19
1<
#6740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#6750000000
1!
1(
b111 1
14
19
0<
#6760000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#6770000000
1!
1(
b1000 1
14
19
1<
#6780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#6790000000
1!
1(
b1001 1
14
07
19
0<
#6800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#6810000000
1!
1(
b0 1
14
19
1<
#6820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#6830000000
1!
1(
b1 1
14
19
0<
#6840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#6850000000
1!
1(
b10 1
14
19
1<
#6860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#6870000000
1!
1(
b11 1
14
19
0<
#6880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#6890000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b100 1
b0001 3
14
17
19
1<
b1001111 >
b0001 ?
#6900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#6910000000
1!
1(
b101 1
14
19
0<
#6920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#6930000000
1!
1(
b110 1
14
19
1<
#6940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#6950000000
1!
1(
b111 1
14
19
0<
#6960000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#6970000000
1!
1(
b1000 1
14
19
1<
#6980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#6990000000
1!
1(
b1001 1
14
07
19
0<
#7000000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#7010000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
1<
#7020000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#7030000000
1!
1(
b1 1
14
19
0<
#7040000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#7050000000
1!
1(
b10 1
14
19
1<
#7060000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#7070000000
1!
1(
b11 1
14
19
0<
#7080000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#7090000000
1!
1(
b100 1
14
17
19
1<
#7100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#7110000000
1!
1(
b101 1
14
19
0<
#7120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#7130000000
1!
1(
b110 1
14
19
1<
#7140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#7150000000
1!
1(
b111 1
14
19
0<
#7160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#7170000000
1!
1(
b1000 1
14
19
1<
#7180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#7190000000
1!
1(
b1001 1
14
07
19
0<
#7200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#7210000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
1<
#7220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#7230000000
1!
1(
b1 1
14
19
0<
#7240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#7250000000
1!
1(
b10 1
14
19
1<
#7260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#7270000000
1!
1(
b11 1
14
19
0<
#7280000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#7290000000
1!
1(
b100 1
14
17
19
1<
#7300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#7310000000
1!
1(
b101 1
14
19
0<
#7320000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#7330000000
1!
1(
b110 1
14
19
1<
#7340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#7350000000
1!
1(
b111 1
14
19
0<
#7360000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#7370000000
1!
1(
b1000 1
14
19
1<
#7380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#7390000000
1!
1(
b1001 1
14
07
19
0<
#7400000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b0 /
b0 2
b0000 3
04
b0 8
09
b0 =
b0000001 >
b0000 ?
#7410000000
1!
1(
b0 1
14
19
1<
#7420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#7430000000
1!
1(
b1 1
14
19
0<
#7440000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#7450000000
1!
1(
b10 1
14
19
1<
#7460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#7470000000
1!
1(
b11 1
14
19
0<
#7480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#7490000000
1!
1(
b100 1
14
17
19
1<
#7500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#7510000000
1!
1(
b101 1
14
19
0<
#7520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#7530000000
1!
1(
b110 1
14
19
1<
#7540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#7550000000
1!
1(
b111 1
14
19
0<
#7560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#7570000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b1000 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#7580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#7590000000
1!
1(
b1001 1
14
07
19
0<
#7600000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#7610000000
1!
b0011 '
1(
b0011 .
b0 1
14
19
1<
#7620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#7630000000
1!
1(
b1 1
14
19
0<
#7640000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#7650000000
1!
1(
b10 1
14
19
1<
#7660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#7670000000
1!
1(
b11 1
14
19
0<
#7680000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#7690000000
1!
1(
b100 1
14
17
19
1<
#7700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#7710000000
1!
1(
b101 1
14
19
0<
#7720000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#7730000000
1!
1(
b110 1
14
19
1<
#7740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#7750000000
1!
1(
b111 1
14
19
0<
#7760000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#7770000000
1!
1(
b1000 1
14
19
1<
#7780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#7790000000
1!
1(
b1001 1
14
07
19
0<
#7800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#7810000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
1<
#7820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#7830000000
1!
1(
b1 1
14
19
0<
#7840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#7850000000
1!
1(
b10 1
14
19
1<
#7860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#7870000000
1!
1(
b11 1
14
19
0<
#7880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#7890000000
1!
1(
b100 1
14
17
19
1<
#7900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#7910000000
1!
1(
b101 1
14
19
0<
#7920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#7930000000
1!
1(
b110 1
14
19
1<
#7940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#7950000000
1!
1(
b111 1
14
19
0<
#7960000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#7970000000
1!
1(
b1000 1
14
19
1<
#7980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#7990000000
1!
1(
b1001 1
14
07
19
0<
#8000000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#8010000000
1!
b1001 '
1(
b1001 .
b0 1
14
19
1<
#8020000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#8030000000
1!
1(
b1 1
14
19
0<
#8040000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#8050000000
1!
1(
b10 1
14
19
1<
#8060000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#8070000000
1!
1(
b11 1
14
19
0<
#8080000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b100 /
b0 2
b0000 3
04
b100 8
09
b0 =
b0000001 >
b0000 ?
#8090000000
1!
1(
b100 1
14
17
19
1<
#8100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#8110000000
1!
1(
b101 1
14
19
0<
#8120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#8130000000
1!
1(
b110 1
14
19
1<
#8140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#8150000000
1!
1(
b111 1
14
19
0<
#8160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#8170000000
1!
1(
b1000 1
14
19
1<
#8180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#8190000000
1!
1(
b1001 1
14
07
19
0<
#8200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#8210000000
1!
1(
b0 1
14
19
1<
#8220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#8230000000
1!
1(
b1 1
14
19
0<
#8240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#8250000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b10 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#8260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#8270000000
1!
1(
b11 1
14
19
0<
#8280000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#8290000000
1!
1(
b100 1
14
17
19
1<
#8300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#8310000000
1!
1(
b101 1
14
19
0<
#8320000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#8330000000
1!
1(
b110 1
14
19
1<
#8340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#8350000000
1!
1(
b111 1
14
19
0<
#8360000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#8370000000
1!
1(
b1000 1
14
19
1<
#8380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#8390000000
1!
1(
b1001 1
14
07
19
0<
#8400000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#8410000000
1!
b1000 '
1(
b1000 .
b0 1
14
19
1<
#8420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#8430000000
1!
1(
b1 1
14
19
0<
#8440000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#8450000000
1!
1(
b10 1
14
19
1<
#8460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#8470000000
1!
1(
b11 1
14
19
0<
#8480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#8490000000
1!
1(
b100 1
14
17
19
1<
#8500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#8510000000
1!
1(
b101 1
14
19
0<
#8520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#8530000000
1!
1(
b110 1
14
19
1<
#8540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#8550000000
1!
1(
b111 1
14
19
0<
#8560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#8570000000
1!
1(
b1000 1
14
19
1<
#8580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#8590000000
1!
1(
b1001 1
14
07
19
0<
#8600000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#8610000000
1!
b1100 '
1(
b1100 .
b0 1
14
19
1<
#8620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#8630000000
1!
1(
b1 1
14
19
0<
#8640000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#8650000000
1!
1(
b10 1
14
19
1<
#8660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#8670000000
1!
1(
b11 1
14
19
0<
#8680000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#8690000000
1!
1(
b100 1
14
17
19
1<
#8700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#8710000000
1!
1(
b101 1
14
19
0<
#8720000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#8730000000
1!
1(
b110 1
14
19
1<
#8740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#8750000000
1!
1(
b111 1
14
19
0<
#8760000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b1000 /
b0 2
b0000 3
04
b1000 8
09
b0 =
b0000001 >
b0000 ?
#8770000000
1!
1(
b1000 1
14
19
1<
#8780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#8790000000
1!
1(
b1001 1
14
07
19
0<
#8800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#8810000000
1!
1(
b0 1
14
19
1<
#8820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#8830000000
1!
1(
b1 1
14
19
0<
#8840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#8850000000
1!
1(
b10 1
14
19
1<
#8860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#8870000000
1!
1(
b11 1
14
19
0<
#8880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#8890000000
1!
1(
b100 1
14
17
19
1<
#8900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#8910000000
1!
1(
b101 1
14
19
0<
#8920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#8930000000
1!
1"
b1001111 &
1(
1)
b1001111 -
b110 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#8940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#8950000000
1!
1(
b111 1
14
19
0<
#8960000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#8970000000
1!
1(
b1000 1
14
19
1<
#8980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#8990000000
1!
1(
b1001 1
14
07
19
0<
#9000000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#9010000000
1!
b0100 '
1(
b0100 .
b0 1
14
19
1<
#9020000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#9030000000
1!
1(
b1 1
14
19
0<
#9040000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#9050000000
1!
1(
b10 1
14
19
1<
#9060000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#9070000000
1!
1(
b11 1
14
19
0<
#9080000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#9090000000
1!
1(
b100 1
14
17
19
1<
#9100000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#9110000000
1!
1(
b101 1
14
19
0<
#9120000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#9130000000
1!
1(
b110 1
14
19
1<
#9140000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#9150000000
1!
1(
b111 1
14
19
0<
#9160000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#9170000000
1!
1(
b1000 1
14
19
1<
#9180000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#9190000000
1!
1(
b1001 1
14
07
19
0<
#9200000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#9210000000
1!
b0110 '
1(
b0110 .
b0 1
14
19
1<
#9220000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#9230000000
1!
1(
b1 1
14
19
0<
#9240000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#9250000000
1!
1(
b10 1
14
19
1<
#9260000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#9270000000
1!
1(
b11 1
14
19
0<
#9280000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#9290000000
1!
1(
b100 1
14
17
19
1<
#9300000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#9310000000
1!
1(
b101 1
14
19
0<
#9320000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#9330000000
1!
1(
b110 1
14
19
1<
#9340000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#9350000000
1!
1(
b111 1
14
19
0<
#9360000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#9370000000
1!
1(
b1000 1
14
19
1<
#9380000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#9390000000
1!
1(
b1001 1
14
07
19
0<
#9400000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#9410000000
1!
b0010 '
1(
b0010 .
b0 1
14
19
1<
#9420000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#9430000000
1!
1(
b1 1
14
19
0<
#9440000000
0!
0"
b0000001 &
0(
0)
b0000001 -
b10 /
b0 2
b0000 3
04
b10 8
09
b0 =
b0000001 >
b0000 ?
#9450000000
1!
1(
b10 1
14
19
1<
#9460000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#9470000000
1!
1(
b11 1
14
19
0<
#9480000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#9490000000
1!
1(
b100 1
14
17
19
1<
#9500000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#9510000000
1!
1(
b101 1
14
19
0<
#9520000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#9530000000
1!
1(
b110 1
14
19
1<
#9540000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#9550000000
1!
1(
b111 1
14
19
0<
#9560000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#9570000000
1!
1(
b1000 1
14
19
1<
#9580000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#9590000000
1!
1(
b1001 1
14
07
19
0<
#9600000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#9610000000
1!
1"
b1001111 &
b0011 '
1(
1)
b1001111 -
b0011 .
b0 1
b0001 3
14
19
1<
b1001111 >
b0001 ?
#9620000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#9630000000
1!
1(
b1 1
14
19
0<
#9640000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#9650000000
1!
1(
b10 1
14
19
1<
#9660000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#9670000000
1!
1(
b11 1
14
19
0<
#9680000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#9690000000
1!
1(
b100 1
14
17
19
1<
#9700000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#9710000000
1!
1(
b101 1
14
19
0<
#9720000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#9730000000
1!
1(
b110 1
14
19
1<
#9740000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#9750000000
1!
1(
b111 1
14
19
0<
#9760000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#9770000000
1!
1(
b1000 1
14
19
1<
#9780000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#9790000000
1!
1(
b1001 1
14
07
19
0<
#9800000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
#9810000000
1!
b0001 '
1(
b0001 .
b0 1
14
19
1<
#9820000000
0!
0(
b1 /
b1 2
04
b1 8
09
b1 =
#9830000000
1!
1(
b1 1
14
19
0<
#9840000000
0!
0(
b10 /
b0 2
04
b10 8
09
b0 =
#9850000000
1!
1(
b10 1
14
19
1<
#9860000000
0!
0(
b11 /
b1 2
04
b11 8
09
b1 =
#9870000000
1!
1(
b11 1
14
19
0<
#9880000000
0!
0(
b100 /
b0 2
04
b100 8
09
b0 =
#9890000000
1!
1(
b100 1
14
17
19
1<
#9900000000
0!
0(
b101 /
b1 2
04
b101 8
09
b1 =
#9910000000
1!
1(
b101 1
14
19
0<
#9920000000
0!
0(
b110 /
b0 2
04
b110 8
09
b0 =
#9930000000
1!
1(
b110 1
14
19
1<
#9940000000
0!
0(
b111 /
b1 2
04
b111 8
09
b1 =
#9950000000
1!
1(
b111 1
14
19
0<
#9960000000
0!
0(
b1000 /
b0 2
04
b1000 8
09
b0 =
#9970000000
1!
1(
b1000 1
14
19
1<
#9980000000
0!
0(
b1001 /
b1 2
04
b1001 8
09
b1 =
#9990000000
1!
1(
b1001 1
14
07
19
0<
#10000000000
0!
0(
b0 /
b0 2
04
b0 8
09
b0 =
