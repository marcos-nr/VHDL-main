$date
  Fri Apr 26 22:35:24 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_tp2_2 $end
$var reg 1 ! clk $end
$var reg 1 " start $end
$var reg 1 # reset $end
$var reg 1 $ led_uv $end
$var reg 1 % led_rojo $end
$var reg 1 & led_conta $end
$var reg 7 ' segmentos[6:0] $end
$var integer 32 ( min_count $end
$var integer 32 ) max_count $end
$scope module uut $end
$var reg 1 * clk $end
$var reg 1 + start $end
$var reg 1 , reset $end
$var reg 1 - led_uv $end
$var reg 1 . led_rojo $end
$var reg 1 / led_conta $end
$var reg 7 0 segmentos[6:0] $end
$var reg 1 1 debounced_start $end
$var reg 1 2 debounced_recet $end
$var reg 1 3 enable_conta $end
$var reg 1 4 reset_conta $end
$var reg 4 5 bcd[3:0] $end
$var integer 32 6 cuenta $end
$var reg 1 7 enable_display $end
$var integer 32 8 segundos $end
$scope module a $end
$var reg 1 9 clk $end
$var reg 1 : key $end
$var reg 1 ; debounced_key $end
$var reg 1 < key_stable $end
$var reg 1 = last_key $end
$upscope $end
$scope module b $end
$var reg 1 > clk $end
$var reg 1 ? key $end
$var reg 1 @ debounced_key $end
$var reg 1 A key_stable $end
$var reg 1 B last_key $end
$upscope $end
$scope module c $end
$var reg 1 C clk $end
$var reg 1 D reset $end
$var reg 1 E enable $end
$var reg 1 F cout $end
$var integer 32 G q $end
$upscope $end
$scope module d $end
$var reg 7 H segmentos[6:0] $end
$var reg 4 I bcd[3:0] $end
$var reg 1 J enable $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
0#
U$
U%
U&
b1111110 '
b0 (
b0 )
0*
0+
0,
U-
U.
U/
b1111110 0
U1
U2
U3
U4
b0000 5
b0 6
17
b0 8
09
0:
U;
U<
U=
0>
0?
U@
UA
UB
0C
UD
UE
UF
b0 G
b1111110 H
b0000 I
1J
#10000000
1!
0&
1*
0/
01
02
19
0;
0<
0=
1>
0@
0A
0B
1C
0F
#20000000
0!
0*
09
0>
0C
#30000000
1!
1*
19
1>
1C
#40000000
0!
1"
0*
1+
09
1:
0>
0C
#50000000
1!
1*
11
19
1;
1<
1=
1>
1C
#60000000
0!
0*
09
0>
0C
#70000000
1!
1*
19
1>
1C
#80000000
0!
0*
09
0>
0C
#90000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#100000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#110000000
1!
1#
1*
1,
12
b1 6
19
1>
1?
1@
1A
1B
1C
b1 G
#120000000
0!
0*
09
0>
0C
#130000000
1!
1*
b10 6
19
1>
1C
b10 G
#140000000
0!
0*
09
0>
0C
#150000000
1!
1*
b11 6
19
1>
1C
b11 G
#160000000
0!
0#
0*
0,
09
0>
0?
0C
#170000000
1!
1&
1*
1/
02
03
14
b100 6
19
1>
0@
0A
0B
1C
1D
0E
1F
b100 G
#180000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#190000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#200000000
0!
0*
09
0>
0C
#210000000
1!
1*
19
1>
1C
#220000000
0!
0*
09
0>
0C
#230000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#240000000
0!
0*
09
0>
0C
#250000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#260000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#270000000
1!
1*
b1 6
19
1>
1C
b1 G
#280000000
0!
0*
09
0>
0C
#290000000
1!
1*
b10 6
19
1>
1C
b10 G
#300000000
0!
0*
09
0>
0C
#310000000
1!
1*
b11 6
19
1>
1C
b11 G
#320000000
0!
0*
09
0>
0C
#330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#340000000
0!
0*
09
0>
0C
#350000000
1!
1*
b101 6
19
1>
1C
b101 G
#360000000
0!
0*
09
0>
0C
#370000000
1!
1*
b110 6
19
1>
1C
b110 G
#380000000
0!
0*
09
0>
0C
#390000000
1!
1*
b111 6
19
1>
1C
b111 G
#400000000
0!
0*
09
0>
0C
#410000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#420000000
0!
0*
09
0>
0C
#430000000
1!
1*
b1 6
19
1>
1C
b1 G
#440000000
0!
0*
09
0>
0C
#450000000
1!
1*
b10 6
19
1>
1C
b10 G
#460000000
0!
0*
09
0>
0C
#470000000
1!
1*
b11 6
19
1>
1C
b11 G
#480000000
0!
0*
09
0>
0C
#490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#500000000
0!
0*
09
0>
0C
#510000000
1!
1*
b101 6
19
1>
1C
b101 G
#520000000
0!
0*
09
0>
0C
#530000000
1!
1*
b110 6
19
1>
1C
b110 G
#540000000
0!
0*
09
0>
0C
#550000000
1!
1*
b111 6
19
1>
1C
b111 G
#560000000
0!
0*
09
0>
0C
#570000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#580000000
0!
0*
09
0>
0C
#590000000
1!
1*
b1 6
19
1>
1C
b1 G
#600000000
0!
0*
09
0>
0C
#610000000
1!
1*
b10 6
19
1>
1C
b10 G
#620000000
0!
0*
09
0>
0C
#630000000
1!
1*
b11 6
19
1>
1C
b11 G
#640000000
0!
0*
09
0>
0C
#650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#660000000
0!
0*
09
0>
0C
#670000000
1!
1*
b101 6
19
1>
1C
b101 G
#680000000
0!
0*
09
0>
0C
#690000000
1!
1*
b110 6
19
1>
1C
b110 G
#700000000
0!
0*
09
0>
0C
#710000000
1!
1*
b111 6
19
1>
1C
b111 G
#720000000
0!
1"
0*
1+
09
1:
0>
0C
#730000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#740000000
0!
0*
09
0>
0C
#750000000
1!
1*
b1 6
19
1>
1C
b1 G
#760000000
0!
0*
09
0>
0C
#770000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#780000000
0!
0*
09
0>
0C
#790000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#800000000
0!
0*
09
0>
0C
#810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#820000000
0!
0*
09
0>
0C
#830000000
1!
1*
b101 6
19
1>
1C
b101 G
#840000000
0!
0#
0*
0,
09
0>
0?
0C
#850000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#860000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#870000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#880000000
0!
0*
09
0>
0C
#890000000
1!
1*
19
1>
1C
#900000000
0!
0*
09
0>
0C
#910000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#920000000
0!
0*
09
0>
0C
#930000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#940000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#950000000
1!
1*
b1 6
19
1>
1C
b1 G
#960000000
0!
0*
09
0>
0C
#970000000
1!
1*
b10 6
19
1>
1C
b10 G
#980000000
0!
0*
09
0>
0C
#990000000
1!
1*
b11 6
19
1>
1C
b11 G
#1000000000
0!
0*
09
0>
0C
#1010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1020000000
0!
0*
09
0>
0C
#1030000000
1!
1*
b101 6
19
1>
1C
b101 G
#1040000000
0!
0*
09
0>
0C
#1050000000
1!
1*
b110 6
19
1>
1C
b110 G
#1060000000
0!
0*
09
0>
0C
#1070000000
1!
1*
b111 6
19
1>
1C
b111 G
#1080000000
0!
0*
09
0>
0C
#1090000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#1100000000
0!
0*
09
0>
0C
#1110000000
1!
1*
b1 6
19
1>
1C
b1 G
#1120000000
0!
0*
09
0>
0C
#1130000000
1!
1*
b10 6
19
1>
1C
b10 G
#1140000000
0!
0*
09
0>
0C
#1150000000
1!
1*
b11 6
19
1>
1C
b11 G
#1160000000
0!
0*
09
0>
0C
#1170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1180000000
0!
0*
09
0>
0C
#1190000000
1!
1*
b101 6
19
1>
1C
b101 G
#1200000000
0!
0*
09
0>
0C
#1210000000
1!
1*
b110 6
19
1>
1C
b110 G
#1220000000
0!
0*
09
0>
0C
#1230000000
1!
1*
b111 6
19
1>
1C
b111 G
#1240000000
0!
0*
09
0>
0C
#1250000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#1260000000
0!
0*
09
0>
0C
#1270000000
1!
1*
b1 6
19
1>
1C
b1 G
#1280000000
0!
0*
09
0>
0C
#1290000000
1!
1*
b10 6
19
1>
1C
b10 G
#1300000000
0!
0*
09
0>
0C
#1310000000
1!
1*
b11 6
19
1>
1C
b11 G
#1320000000
0!
0*
09
0>
0C
#1330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1340000000
0!
0*
09
0>
0C
#1350000000
1!
1*
b101 6
19
1>
1C
b101 G
#1360000000
0!
0*
09
0>
0C
#1370000000
1!
1*
b110 6
19
1>
1C
b110 G
#1380000000
0!
0*
09
0>
0C
#1390000000
1!
1*
b111 6
19
1>
1C
b111 G
#1400000000
0!
1"
0*
1+
09
1:
0>
0C
#1410000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#1420000000
0!
0*
09
0>
0C
#1430000000
1!
1*
b1 6
19
1>
1C
b1 G
#1440000000
0!
0*
09
0>
0C
#1450000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#1460000000
0!
0*
09
0>
0C
#1470000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#1480000000
0!
0*
09
0>
0C
#1490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1500000000
0!
0*
09
0>
0C
#1510000000
1!
1*
b101 6
19
1>
1C
b101 G
#1520000000
0!
0#
0*
0,
09
0>
0?
0C
#1530000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#1540000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#1550000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#1560000000
0!
0*
09
0>
0C
#1570000000
1!
1*
19
1>
1C
#1580000000
0!
0*
09
0>
0C
#1590000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#1600000000
0!
0*
09
0>
0C
#1610000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#1620000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#1630000000
1!
1*
b1 6
19
1>
1C
b1 G
#1640000000
0!
0*
09
0>
0C
#1650000000
1!
1*
b10 6
19
1>
1C
b10 G
#1660000000
0!
0*
09
0>
0C
#1670000000
1!
1*
b11 6
19
1>
1C
b11 G
#1680000000
0!
0*
09
0>
0C
#1690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1700000000
0!
0*
09
0>
0C
#1710000000
1!
1*
b101 6
19
1>
1C
b101 G
#1720000000
0!
0*
09
0>
0C
#1730000000
1!
1*
b110 6
19
1>
1C
b110 G
#1740000000
0!
0*
09
0>
0C
#1750000000
1!
1*
b111 6
19
1>
1C
b111 G
#1760000000
0!
0*
09
0>
0C
#1770000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#1780000000
0!
0*
09
0>
0C
#1790000000
1!
1*
b1 6
19
1>
1C
b1 G
#1800000000
0!
0*
09
0>
0C
#1810000000
1!
1*
b10 6
19
1>
1C
b10 G
#1820000000
0!
0*
09
0>
0C
#1830000000
1!
1*
b11 6
19
1>
1C
b11 G
#1840000000
0!
0*
09
0>
0C
#1850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#1860000000
0!
0*
09
0>
0C
#1870000000
1!
1*
b101 6
19
1>
1C
b101 G
#1880000000
0!
0*
09
0>
0C
#1890000000
1!
1*
b110 6
19
1>
1C
b110 G
#1900000000
0!
0*
09
0>
0C
#1910000000
1!
1*
b111 6
19
1>
1C
b111 G
#1920000000
0!
0*
09
0>
0C
#1930000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#1940000000
0!
0*
09
0>
0C
#1950000000
1!
1*
b1 6
19
1>
1C
b1 G
#1960000000
0!
0*
09
0>
0C
#1970000000
1!
1*
b10 6
19
1>
1C
b10 G
#1980000000
0!
0*
09
0>
0C
#1990000000
1!
1*
b11 6
19
1>
1C
b11 G
#2000000000
0!
0*
09
0>
0C
#2010000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2020000000
0!
0*
09
0>
0C
#2030000000
1!
1*
b101 6
19
1>
1C
b101 G
#2040000000
0!
0*
09
0>
0C
#2050000000
1!
1*
b110 6
19
1>
1C
b110 G
#2060000000
0!
0*
09
0>
0C
#2070000000
1!
1*
b111 6
19
1>
1C
b111 G
#2080000000
0!
1"
0*
1+
09
1:
0>
0C
#2090000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#2100000000
0!
0*
09
0>
0C
#2110000000
1!
1*
b1 6
19
1>
1C
b1 G
#2120000000
0!
0*
09
0>
0C
#2130000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#2140000000
0!
0*
09
0>
0C
#2150000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#2160000000
0!
0*
09
0>
0C
#2170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2180000000
0!
0*
09
0>
0C
#2190000000
1!
1*
b101 6
19
1>
1C
b101 G
#2200000000
0!
0#
0*
0,
09
0>
0?
0C
#2210000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#2220000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#2230000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#2240000000
0!
0*
09
0>
0C
#2250000000
1!
1*
19
1>
1C
#2260000000
0!
0*
09
0>
0C
#2270000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#2280000000
0!
0*
09
0>
0C
#2290000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#2300000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#2310000000
1!
1*
b1 6
19
1>
1C
b1 G
#2320000000
0!
0*
09
0>
0C
#2330000000
1!
1*
b10 6
19
1>
1C
b10 G
#2340000000
0!
0*
09
0>
0C
#2350000000
1!
1*
b11 6
19
1>
1C
b11 G
#2360000000
0!
0*
09
0>
0C
#2370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2380000000
0!
0*
09
0>
0C
#2390000000
1!
1*
b101 6
19
1>
1C
b101 G
#2400000000
0!
0*
09
0>
0C
#2410000000
1!
1*
b110 6
19
1>
1C
b110 G
#2420000000
0!
0*
09
0>
0C
#2430000000
1!
1*
b111 6
19
1>
1C
b111 G
#2440000000
0!
0*
09
0>
0C
#2450000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#2460000000
0!
0*
09
0>
0C
#2470000000
1!
1*
b1 6
19
1>
1C
b1 G
#2480000000
0!
0*
09
0>
0C
#2490000000
1!
1*
b10 6
19
1>
1C
b10 G
#2500000000
0!
0*
09
0>
0C
#2510000000
1!
1*
b11 6
19
1>
1C
b11 G
#2520000000
0!
0*
09
0>
0C
#2530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2540000000
0!
0*
09
0>
0C
#2550000000
1!
1*
b101 6
19
1>
1C
b101 G
#2560000000
0!
0*
09
0>
0C
#2570000000
1!
1*
b110 6
19
1>
1C
b110 G
#2580000000
0!
0*
09
0>
0C
#2590000000
1!
1*
b111 6
19
1>
1C
b111 G
#2600000000
0!
0*
09
0>
0C
#2610000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#2620000000
0!
0*
09
0>
0C
#2630000000
1!
1*
b1 6
19
1>
1C
b1 G
#2640000000
0!
0*
09
0>
0C
#2650000000
1!
1*
b10 6
19
1>
1C
b10 G
#2660000000
0!
0*
09
0>
0C
#2670000000
1!
1*
b11 6
19
1>
1C
b11 G
#2680000000
0!
0*
09
0>
0C
#2690000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2700000000
0!
0*
09
0>
0C
#2710000000
1!
1*
b101 6
19
1>
1C
b101 G
#2720000000
0!
0*
09
0>
0C
#2730000000
1!
1*
b110 6
19
1>
1C
b110 G
#2740000000
0!
0*
09
0>
0C
#2750000000
1!
1*
b111 6
19
1>
1C
b111 G
#2760000000
0!
1"
0*
1+
09
1:
0>
0C
#2770000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#2780000000
0!
0*
09
0>
0C
#2790000000
1!
1*
b1 6
19
1>
1C
b1 G
#2800000000
0!
0*
09
0>
0C
#2810000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#2820000000
0!
0*
09
0>
0C
#2830000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#2840000000
0!
0*
09
0>
0C
#2850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#2860000000
0!
0*
09
0>
0C
#2870000000
1!
1*
b101 6
19
1>
1C
b101 G
#2880000000
0!
0#
0*
0,
09
0>
0?
0C
#2890000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#2900000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#2910000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#2920000000
0!
0*
09
0>
0C
#2930000000
1!
1*
19
1>
1C
#2940000000
0!
0*
09
0>
0C
#2950000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#2960000000
0!
0*
09
0>
0C
#2970000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#2980000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#2990000000
1!
1*
b1 6
19
1>
1C
b1 G
#3000000000
0!
0*
09
0>
0C
#3010000000
1!
1*
b10 6
19
1>
1C
b10 G
#3020000000
0!
0*
09
0>
0C
#3030000000
1!
1*
b11 6
19
1>
1C
b11 G
#3040000000
0!
0*
09
0>
0C
#3050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3060000000
0!
0*
09
0>
0C
#3070000000
1!
1*
b101 6
19
1>
1C
b101 G
#3080000000
0!
0*
09
0>
0C
#3090000000
1!
1*
b110 6
19
1>
1C
b110 G
#3100000000
0!
0*
09
0>
0C
#3110000000
1!
1*
b111 6
19
1>
1C
b111 G
#3120000000
0!
0*
09
0>
0C
#3130000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#3140000000
0!
0*
09
0>
0C
#3150000000
1!
1*
b1 6
19
1>
1C
b1 G
#3160000000
0!
0*
09
0>
0C
#3170000000
1!
1*
b10 6
19
1>
1C
b10 G
#3180000000
0!
0*
09
0>
0C
#3190000000
1!
1*
b11 6
19
1>
1C
b11 G
#3200000000
0!
0*
09
0>
0C
#3210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3220000000
0!
0*
09
0>
0C
#3230000000
1!
1*
b101 6
19
1>
1C
b101 G
#3240000000
0!
0*
09
0>
0C
#3250000000
1!
1*
b110 6
19
1>
1C
b110 G
#3260000000
0!
0*
09
0>
0C
#3270000000
1!
1*
b111 6
19
1>
1C
b111 G
#3280000000
0!
0*
09
0>
0C
#3290000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#3300000000
0!
0*
09
0>
0C
#3310000000
1!
1*
b1 6
19
1>
1C
b1 G
#3320000000
0!
0*
09
0>
0C
#3330000000
1!
1*
b10 6
19
1>
1C
b10 G
#3340000000
0!
0*
09
0>
0C
#3350000000
1!
1*
b11 6
19
1>
1C
b11 G
#3360000000
0!
0*
09
0>
0C
#3370000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3380000000
0!
0*
09
0>
0C
#3390000000
1!
1*
b101 6
19
1>
1C
b101 G
#3400000000
0!
0*
09
0>
0C
#3410000000
1!
1*
b110 6
19
1>
1C
b110 G
#3420000000
0!
0*
09
0>
0C
#3430000000
1!
1*
b111 6
19
1>
1C
b111 G
#3440000000
0!
1"
0*
1+
09
1:
0>
0C
#3450000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#3460000000
0!
0*
09
0>
0C
#3470000000
1!
1*
b1 6
19
1>
1C
b1 G
#3480000000
0!
0*
09
0>
0C
#3490000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#3500000000
0!
0*
09
0>
0C
#3510000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#3520000000
0!
0*
09
0>
0C
#3530000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3540000000
0!
0*
09
0>
0C
#3550000000
1!
1*
b101 6
19
1>
1C
b101 G
#3560000000
0!
0#
0*
0,
09
0>
0?
0C
#3570000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#3580000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#3590000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#3600000000
0!
0*
09
0>
0C
#3610000000
1!
1*
19
1>
1C
#3620000000
0!
0*
09
0>
0C
#3630000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#3640000000
0!
0*
09
0>
0C
#3650000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#3660000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#3670000000
1!
1*
b1 6
19
1>
1C
b1 G
#3680000000
0!
0*
09
0>
0C
#3690000000
1!
1*
b10 6
19
1>
1C
b10 G
#3700000000
0!
0*
09
0>
0C
#3710000000
1!
1*
b11 6
19
1>
1C
b11 G
#3720000000
0!
0*
09
0>
0C
#3730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3740000000
0!
0*
09
0>
0C
#3750000000
1!
1*
b101 6
19
1>
1C
b101 G
#3760000000
0!
0*
09
0>
0C
#3770000000
1!
1*
b110 6
19
1>
1C
b110 G
#3780000000
0!
0*
09
0>
0C
#3790000000
1!
1*
b111 6
19
1>
1C
b111 G
#3800000000
0!
0*
09
0>
0C
#3810000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#3820000000
0!
0*
09
0>
0C
#3830000000
1!
1*
b1 6
19
1>
1C
b1 G
#3840000000
0!
0*
09
0>
0C
#3850000000
1!
1*
b10 6
19
1>
1C
b10 G
#3860000000
0!
0*
09
0>
0C
#3870000000
1!
1*
b11 6
19
1>
1C
b11 G
#3880000000
0!
0*
09
0>
0C
#3890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#3900000000
0!
0*
09
0>
0C
#3910000000
1!
1*
b101 6
19
1>
1C
b101 G
#3920000000
0!
0*
09
0>
0C
#3930000000
1!
1*
b110 6
19
1>
1C
b110 G
#3940000000
0!
0*
09
0>
0C
#3950000000
1!
1*
b111 6
19
1>
1C
b111 G
#3960000000
0!
0*
09
0>
0C
#3970000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#3980000000
0!
0*
09
0>
0C
#3990000000
1!
1*
b1 6
19
1>
1C
b1 G
#4000000000
0!
0*
09
0>
0C
#4010000000
1!
1*
b10 6
19
1>
1C
b10 G
#4020000000
0!
0*
09
0>
0C
#4030000000
1!
1*
b11 6
19
1>
1C
b11 G
#4040000000
0!
0*
09
0>
0C
#4050000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4060000000
0!
0*
09
0>
0C
#4070000000
1!
1*
b101 6
19
1>
1C
b101 G
#4080000000
0!
0*
09
0>
0C
#4090000000
1!
1*
b110 6
19
1>
1C
b110 G
#4100000000
0!
0*
09
0>
0C
#4110000000
1!
1*
b111 6
19
1>
1C
b111 G
#4120000000
0!
1"
0*
1+
09
1:
0>
0C
#4130000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#4140000000
0!
0*
09
0>
0C
#4150000000
1!
1*
b1 6
19
1>
1C
b1 G
#4160000000
0!
0*
09
0>
0C
#4170000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#4180000000
0!
0*
09
0>
0C
#4190000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#4200000000
0!
0*
09
0>
0C
#4210000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4220000000
0!
0*
09
0>
0C
#4230000000
1!
1*
b101 6
19
1>
1C
b101 G
#4240000000
0!
0#
0*
0,
09
0>
0?
0C
#4250000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#4260000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#4270000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#4280000000
0!
0*
09
0>
0C
#4290000000
1!
1*
19
1>
1C
#4300000000
0!
0*
09
0>
0C
#4310000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#4320000000
0!
0*
09
0>
0C
#4330000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#4340000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#4350000000
1!
1*
b1 6
19
1>
1C
b1 G
#4360000000
0!
0*
09
0>
0C
#4370000000
1!
1*
b10 6
19
1>
1C
b10 G
#4380000000
0!
0*
09
0>
0C
#4390000000
1!
1*
b11 6
19
1>
1C
b11 G
#4400000000
0!
0*
09
0>
0C
#4410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4420000000
0!
0*
09
0>
0C
#4430000000
1!
1*
b101 6
19
1>
1C
b101 G
#4440000000
0!
0*
09
0>
0C
#4450000000
1!
1*
b110 6
19
1>
1C
b110 G
#4460000000
0!
0*
09
0>
0C
#4470000000
1!
1*
b111 6
19
1>
1C
b111 G
#4480000000
0!
0*
09
0>
0C
#4490000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#4500000000
0!
0*
09
0>
0C
#4510000000
1!
1*
b1 6
19
1>
1C
b1 G
#4520000000
0!
0*
09
0>
0C
#4530000000
1!
1*
b10 6
19
1>
1C
b10 G
#4540000000
0!
0*
09
0>
0C
#4550000000
1!
1*
b11 6
19
1>
1C
b11 G
#4560000000
0!
0*
09
0>
0C
#4570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4580000000
0!
0*
09
0>
0C
#4590000000
1!
1*
b101 6
19
1>
1C
b101 G
#4600000000
0!
0*
09
0>
0C
#4610000000
1!
1*
b110 6
19
1>
1C
b110 G
#4620000000
0!
0*
09
0>
0C
#4630000000
1!
1*
b111 6
19
1>
1C
b111 G
#4640000000
0!
0*
09
0>
0C
#4650000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#4660000000
0!
0*
09
0>
0C
#4670000000
1!
1*
b1 6
19
1>
1C
b1 G
#4680000000
0!
0*
09
0>
0C
#4690000000
1!
1*
b10 6
19
1>
1C
b10 G
#4700000000
0!
0*
09
0>
0C
#4710000000
1!
1*
b11 6
19
1>
1C
b11 G
#4720000000
0!
0*
09
0>
0C
#4730000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4740000000
0!
0*
09
0>
0C
#4750000000
1!
1*
b101 6
19
1>
1C
b101 G
#4760000000
0!
0*
09
0>
0C
#4770000000
1!
1*
b110 6
19
1>
1C
b110 G
#4780000000
0!
0*
09
0>
0C
#4790000000
1!
1*
b111 6
19
1>
1C
b111 G
#4800000000
0!
1"
0*
1+
09
1:
0>
0C
#4810000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#4820000000
0!
0*
09
0>
0C
#4830000000
1!
1*
b1 6
19
1>
1C
b1 G
#4840000000
0!
0*
09
0>
0C
#4850000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#4860000000
0!
0*
09
0>
0C
#4870000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#4880000000
0!
0*
09
0>
0C
#4890000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#4900000000
0!
0*
09
0>
0C
#4910000000
1!
1*
b101 6
19
1>
1C
b101 G
#4920000000
0!
0#
0*
0,
09
0>
0?
0C
#4930000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#4940000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#4950000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#4960000000
0!
0*
09
0>
0C
#4970000000
1!
1*
19
1>
1C
#4980000000
0!
0*
09
0>
0C
#4990000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#5000000000
0!
0*
09
0>
0C
#5010000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#5020000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#5030000000
1!
1*
b1 6
19
1>
1C
b1 G
#5040000000
0!
0*
09
0>
0C
#5050000000
1!
1*
b10 6
19
1>
1C
b10 G
#5060000000
0!
0*
09
0>
0C
#5070000000
1!
1*
b11 6
19
1>
1C
b11 G
#5080000000
0!
0*
09
0>
0C
#5090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5100000000
0!
0*
09
0>
0C
#5110000000
1!
1*
b101 6
19
1>
1C
b101 G
#5120000000
0!
0*
09
0>
0C
#5130000000
1!
1*
b110 6
19
1>
1C
b110 G
#5140000000
0!
0*
09
0>
0C
#5150000000
1!
1*
b111 6
19
1>
1C
b111 G
#5160000000
0!
0*
09
0>
0C
#5170000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#5180000000
0!
0*
09
0>
0C
#5190000000
1!
1*
b1 6
19
1>
1C
b1 G
#5200000000
0!
0*
09
0>
0C
#5210000000
1!
1*
b10 6
19
1>
1C
b10 G
#5220000000
0!
0*
09
0>
0C
#5230000000
1!
1*
b11 6
19
1>
1C
b11 G
#5240000000
0!
0*
09
0>
0C
#5250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5260000000
0!
0*
09
0>
0C
#5270000000
1!
1*
b101 6
19
1>
1C
b101 G
#5280000000
0!
0*
09
0>
0C
#5290000000
1!
1*
b110 6
19
1>
1C
b110 G
#5300000000
0!
0*
09
0>
0C
#5310000000
1!
1*
b111 6
19
1>
1C
b111 G
#5320000000
0!
0*
09
0>
0C
#5330000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#5340000000
0!
0*
09
0>
0C
#5350000000
1!
1*
b1 6
19
1>
1C
b1 G
#5360000000
0!
0*
09
0>
0C
#5370000000
1!
1*
b10 6
19
1>
1C
b10 G
#5380000000
0!
0*
09
0>
0C
#5390000000
1!
1*
b11 6
19
1>
1C
b11 G
#5400000000
0!
0*
09
0>
0C
#5410000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5420000000
0!
0*
09
0>
0C
#5430000000
1!
1*
b101 6
19
1>
1C
b101 G
#5440000000
0!
0*
09
0>
0C
#5450000000
1!
1*
b110 6
19
1>
1C
b110 G
#5460000000
0!
0*
09
0>
0C
#5470000000
1!
1*
b111 6
19
1>
1C
b111 G
#5480000000
0!
1"
0*
1+
09
1:
0>
0C
#5490000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#5500000000
0!
0*
09
0>
0C
#5510000000
1!
1*
b1 6
19
1>
1C
b1 G
#5520000000
0!
0*
09
0>
0C
#5530000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#5540000000
0!
0*
09
0>
0C
#5550000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#5560000000
0!
0*
09
0>
0C
#5570000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5580000000
0!
0*
09
0>
0C
#5590000000
1!
1*
b101 6
19
1>
1C
b101 G
#5600000000
0!
0#
0*
0,
09
0>
0?
0C
#5610000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#5620000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#5630000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#5640000000
0!
0*
09
0>
0C
#5650000000
1!
1*
19
1>
1C
#5660000000
0!
0*
09
0>
0C
#5670000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#5680000000
0!
0*
09
0>
0C
#5690000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#5700000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#5710000000
1!
1*
b1 6
19
1>
1C
b1 G
#5720000000
0!
0*
09
0>
0C
#5730000000
1!
1*
b10 6
19
1>
1C
b10 G
#5740000000
0!
0*
09
0>
0C
#5750000000
1!
1*
b11 6
19
1>
1C
b11 G
#5760000000
0!
0*
09
0>
0C
#5770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5780000000
0!
0*
09
0>
0C
#5790000000
1!
1*
b101 6
19
1>
1C
b101 G
#5800000000
0!
0*
09
0>
0C
#5810000000
1!
1*
b110 6
19
1>
1C
b110 G
#5820000000
0!
0*
09
0>
0C
#5830000000
1!
1*
b111 6
19
1>
1C
b111 G
#5840000000
0!
0*
09
0>
0C
#5850000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#5860000000
0!
0*
09
0>
0C
#5870000000
1!
1*
b1 6
19
1>
1C
b1 G
#5880000000
0!
0*
09
0>
0C
#5890000000
1!
1*
b10 6
19
1>
1C
b10 G
#5900000000
0!
0*
09
0>
0C
#5910000000
1!
1*
b11 6
19
1>
1C
b11 G
#5920000000
0!
0*
09
0>
0C
#5930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#5940000000
0!
0*
09
0>
0C
#5950000000
1!
1*
b101 6
19
1>
1C
b101 G
#5960000000
0!
0*
09
0>
0C
#5970000000
1!
1*
b110 6
19
1>
1C
b110 G
#5980000000
0!
0*
09
0>
0C
#5990000000
1!
1*
b111 6
19
1>
1C
b111 G
#6000000000
0!
0*
09
0>
0C
#6010000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#6020000000
0!
0*
09
0>
0C
#6030000000
1!
1*
b1 6
19
1>
1C
b1 G
#6040000000
0!
0*
09
0>
0C
#6050000000
1!
1*
b10 6
19
1>
1C
b10 G
#6060000000
0!
0*
09
0>
0C
#6070000000
1!
1*
b11 6
19
1>
1C
b11 G
#6080000000
0!
0*
09
0>
0C
#6090000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6100000000
0!
0*
09
0>
0C
#6110000000
1!
1*
b101 6
19
1>
1C
b101 G
#6120000000
0!
0*
09
0>
0C
#6130000000
1!
1*
b110 6
19
1>
1C
b110 G
#6140000000
0!
0*
09
0>
0C
#6150000000
1!
1*
b111 6
19
1>
1C
b111 G
#6160000000
0!
1"
0*
1+
09
1:
0>
0C
#6170000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#6180000000
0!
0*
09
0>
0C
#6190000000
1!
1*
b1 6
19
1>
1C
b1 G
#6200000000
0!
0*
09
0>
0C
#6210000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#6220000000
0!
0*
09
0>
0C
#6230000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#6240000000
0!
0*
09
0>
0C
#6250000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6260000000
0!
0*
09
0>
0C
#6270000000
1!
1*
b101 6
19
1>
1C
b101 G
#6280000000
0!
0#
0*
0,
09
0>
0?
0C
#6290000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#6300000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#6310000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#6320000000
0!
0*
09
0>
0C
#6330000000
1!
1*
19
1>
1C
#6340000000
0!
0*
09
0>
0C
#6350000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#6360000000
0!
0*
09
0>
0C
#6370000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#6380000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#6390000000
1!
1*
b1 6
19
1>
1C
b1 G
#6400000000
0!
0*
09
0>
0C
#6410000000
1!
1*
b10 6
19
1>
1C
b10 G
#6420000000
0!
0*
09
0>
0C
#6430000000
1!
1*
b11 6
19
1>
1C
b11 G
#6440000000
0!
0*
09
0>
0C
#6450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6460000000
0!
0*
09
0>
0C
#6470000000
1!
1*
b101 6
19
1>
1C
b101 G
#6480000000
0!
0*
09
0>
0C
#6490000000
1!
1*
b110 6
19
1>
1C
b110 G
#6500000000
0!
0*
09
0>
0C
#6510000000
1!
1*
b111 6
19
1>
1C
b111 G
#6520000000
0!
0*
09
0>
0C
#6530000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#6540000000
0!
0*
09
0>
0C
#6550000000
1!
1*
b1 6
19
1>
1C
b1 G
#6560000000
0!
0*
09
0>
0C
#6570000000
1!
1*
b10 6
19
1>
1C
b10 G
#6580000000
0!
0*
09
0>
0C
#6590000000
1!
1*
b11 6
19
1>
1C
b11 G
#6600000000
0!
0*
09
0>
0C
#6610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6620000000
0!
0*
09
0>
0C
#6630000000
1!
1*
b101 6
19
1>
1C
b101 G
#6640000000
0!
0*
09
0>
0C
#6650000000
1!
1*
b110 6
19
1>
1C
b110 G
#6660000000
0!
0*
09
0>
0C
#6670000000
1!
1*
b111 6
19
1>
1C
b111 G
#6680000000
0!
0*
09
0>
0C
#6690000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#6700000000
0!
0*
09
0>
0C
#6710000000
1!
1*
b1 6
19
1>
1C
b1 G
#6720000000
0!
0*
09
0>
0C
#6730000000
1!
1*
b10 6
19
1>
1C
b10 G
#6740000000
0!
0*
09
0>
0C
#6750000000
1!
1*
b11 6
19
1>
1C
b11 G
#6760000000
0!
0*
09
0>
0C
#6770000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6780000000
0!
0*
09
0>
0C
#6790000000
1!
1*
b101 6
19
1>
1C
b101 G
#6800000000
0!
0*
09
0>
0C
#6810000000
1!
1*
b110 6
19
1>
1C
b110 G
#6820000000
0!
0*
09
0>
0C
#6830000000
1!
1*
b111 6
19
1>
1C
b111 G
#6840000000
0!
1"
0*
1+
09
1:
0>
0C
#6850000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#6860000000
0!
0*
09
0>
0C
#6870000000
1!
1*
b1 6
19
1>
1C
b1 G
#6880000000
0!
0*
09
0>
0C
#6890000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#6900000000
0!
0*
09
0>
0C
#6910000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#6920000000
0!
0*
09
0>
0C
#6930000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#6940000000
0!
0*
09
0>
0C
#6950000000
1!
1*
b101 6
19
1>
1C
b101 G
#6960000000
0!
0#
0*
0,
09
0>
0?
0C
#6970000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#6980000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#6990000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#7000000000
0!
0*
09
0>
0C
#7010000000
1!
1*
19
1>
1C
#7020000000
0!
0*
09
0>
0C
#7030000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#7040000000
0!
0*
09
0>
0C
#7050000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#7060000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#7070000000
1!
1*
b1 6
19
1>
1C
b1 G
#7080000000
0!
0*
09
0>
0C
#7090000000
1!
1*
b10 6
19
1>
1C
b10 G
#7100000000
0!
0*
09
0>
0C
#7110000000
1!
1*
b11 6
19
1>
1C
b11 G
#7120000000
0!
0*
09
0>
0C
#7130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7140000000
0!
0*
09
0>
0C
#7150000000
1!
1*
b101 6
19
1>
1C
b101 G
#7160000000
0!
0*
09
0>
0C
#7170000000
1!
1*
b110 6
19
1>
1C
b110 G
#7180000000
0!
0*
09
0>
0C
#7190000000
1!
1*
b111 6
19
1>
1C
b111 G
#7200000000
0!
0*
09
0>
0C
#7210000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#7220000000
0!
0*
09
0>
0C
#7230000000
1!
1*
b1 6
19
1>
1C
b1 G
#7240000000
0!
0*
09
0>
0C
#7250000000
1!
1*
b10 6
19
1>
1C
b10 G
#7260000000
0!
0*
09
0>
0C
#7270000000
1!
1*
b11 6
19
1>
1C
b11 G
#7280000000
0!
0*
09
0>
0C
#7290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7300000000
0!
0*
09
0>
0C
#7310000000
1!
1*
b101 6
19
1>
1C
b101 G
#7320000000
0!
0*
09
0>
0C
#7330000000
1!
1*
b110 6
19
1>
1C
b110 G
#7340000000
0!
0*
09
0>
0C
#7350000000
1!
1*
b111 6
19
1>
1C
b111 G
#7360000000
0!
0*
09
0>
0C
#7370000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#7380000000
0!
0*
09
0>
0C
#7390000000
1!
1*
b1 6
19
1>
1C
b1 G
#7400000000
0!
0*
09
0>
0C
#7410000000
1!
1*
b10 6
19
1>
1C
b10 G
#7420000000
0!
0*
09
0>
0C
#7430000000
1!
1*
b11 6
19
1>
1C
b11 G
#7440000000
0!
0*
09
0>
0C
#7450000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7460000000
0!
0*
09
0>
0C
#7470000000
1!
1*
b101 6
19
1>
1C
b101 G
#7480000000
0!
0*
09
0>
0C
#7490000000
1!
1*
b110 6
19
1>
1C
b110 G
#7500000000
0!
0*
09
0>
0C
#7510000000
1!
1*
b111 6
19
1>
1C
b111 G
#7520000000
0!
1"
0*
1+
09
1:
0>
0C
#7530000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#7540000000
0!
0*
09
0>
0C
#7550000000
1!
1*
b1 6
19
1>
1C
b1 G
#7560000000
0!
0*
09
0>
0C
#7570000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#7580000000
0!
0*
09
0>
0C
#7590000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#7600000000
0!
0*
09
0>
0C
#7610000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7620000000
0!
0*
09
0>
0C
#7630000000
1!
1*
b101 6
19
1>
1C
b101 G
#7640000000
0!
0#
0*
0,
09
0>
0?
0C
#7650000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#7660000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#7670000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#7680000000
0!
0*
09
0>
0C
#7690000000
1!
1*
19
1>
1C
#7700000000
0!
0*
09
0>
0C
#7710000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#7720000000
0!
0*
09
0>
0C
#7730000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#7740000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#7750000000
1!
1*
b1 6
19
1>
1C
b1 G
#7760000000
0!
0*
09
0>
0C
#7770000000
1!
1*
b10 6
19
1>
1C
b10 G
#7780000000
0!
0*
09
0>
0C
#7790000000
1!
1*
b11 6
19
1>
1C
b11 G
#7800000000
0!
0*
09
0>
0C
#7810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7820000000
0!
0*
09
0>
0C
#7830000000
1!
1*
b101 6
19
1>
1C
b101 G
#7840000000
0!
0*
09
0>
0C
#7850000000
1!
1*
b110 6
19
1>
1C
b110 G
#7860000000
0!
0*
09
0>
0C
#7870000000
1!
1*
b111 6
19
1>
1C
b111 G
#7880000000
0!
0*
09
0>
0C
#7890000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#7900000000
0!
0*
09
0>
0C
#7910000000
1!
1*
b1 6
19
1>
1C
b1 G
#7920000000
0!
0*
09
0>
0C
#7930000000
1!
1*
b10 6
19
1>
1C
b10 G
#7940000000
0!
0*
09
0>
0C
#7950000000
1!
1*
b11 6
19
1>
1C
b11 G
#7960000000
0!
0*
09
0>
0C
#7970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#7980000000
0!
0*
09
0>
0C
#7990000000
1!
1*
b101 6
19
1>
1C
b101 G
#8000000000
0!
0*
09
0>
0C
#8010000000
1!
1*
b110 6
19
1>
1C
b110 G
#8020000000
0!
0*
09
0>
0C
#8030000000
1!
1*
b111 6
19
1>
1C
b111 G
#8040000000
0!
0*
09
0>
0C
#8050000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#8060000000
0!
0*
09
0>
0C
#8070000000
1!
1*
b1 6
19
1>
1C
b1 G
#8080000000
0!
0*
09
0>
0C
#8090000000
1!
1*
b10 6
19
1>
1C
b10 G
#8100000000
0!
0*
09
0>
0C
#8110000000
1!
1*
b11 6
19
1>
1C
b11 G
#8120000000
0!
0*
09
0>
0C
#8130000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8140000000
0!
0*
09
0>
0C
#8150000000
1!
1*
b101 6
19
1>
1C
b101 G
#8160000000
0!
0*
09
0>
0C
#8170000000
1!
1*
b110 6
19
1>
1C
b110 G
#8180000000
0!
0*
09
0>
0C
#8190000000
1!
1*
b111 6
19
1>
1C
b111 G
#8200000000
0!
1"
0*
1+
09
1:
0>
0C
#8210000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#8220000000
0!
0*
09
0>
0C
#8230000000
1!
1*
b1 6
19
1>
1C
b1 G
#8240000000
0!
0*
09
0>
0C
#8250000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#8260000000
0!
0*
09
0>
0C
#8270000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#8280000000
0!
0*
09
0>
0C
#8290000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8300000000
0!
0*
09
0>
0C
#8310000000
1!
1*
b101 6
19
1>
1C
b101 G
#8320000000
0!
0#
0*
0,
09
0>
0?
0C
#8330000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#8340000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#8350000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#8360000000
0!
0*
09
0>
0C
#8370000000
1!
1*
19
1>
1C
#8380000000
0!
0*
09
0>
0C
#8390000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#8400000000
0!
0*
09
0>
0C
#8410000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#8420000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#8430000000
1!
1*
b1 6
19
1>
1C
b1 G
#8440000000
0!
0*
09
0>
0C
#8450000000
1!
1*
b10 6
19
1>
1C
b10 G
#8460000000
0!
0*
09
0>
0C
#8470000000
1!
1*
b11 6
19
1>
1C
b11 G
#8480000000
0!
0*
09
0>
0C
#8490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8500000000
0!
0*
09
0>
0C
#8510000000
1!
1*
b101 6
19
1>
1C
b101 G
#8520000000
0!
0*
09
0>
0C
#8530000000
1!
1*
b110 6
19
1>
1C
b110 G
#8540000000
0!
0*
09
0>
0C
#8550000000
1!
1*
b111 6
19
1>
1C
b111 G
#8560000000
0!
0*
09
0>
0C
#8570000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#8580000000
0!
0*
09
0>
0C
#8590000000
1!
1*
b1 6
19
1>
1C
b1 G
#8600000000
0!
0*
09
0>
0C
#8610000000
1!
1*
b10 6
19
1>
1C
b10 G
#8620000000
0!
0*
09
0>
0C
#8630000000
1!
1*
b11 6
19
1>
1C
b11 G
#8640000000
0!
0*
09
0>
0C
#8650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8660000000
0!
0*
09
0>
0C
#8670000000
1!
1*
b101 6
19
1>
1C
b101 G
#8680000000
0!
0*
09
0>
0C
#8690000000
1!
1*
b110 6
19
1>
1C
b110 G
#8700000000
0!
0*
09
0>
0C
#8710000000
1!
1*
b111 6
19
1>
1C
b111 G
#8720000000
0!
0*
09
0>
0C
#8730000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#8740000000
0!
0*
09
0>
0C
#8750000000
1!
1*
b1 6
19
1>
1C
b1 G
#8760000000
0!
0*
09
0>
0C
#8770000000
1!
1*
b10 6
19
1>
1C
b10 G
#8780000000
0!
0*
09
0>
0C
#8790000000
1!
1*
b11 6
19
1>
1C
b11 G
#8800000000
0!
0*
09
0>
0C
#8810000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8820000000
0!
0*
09
0>
0C
#8830000000
1!
1*
b101 6
19
1>
1C
b101 G
#8840000000
0!
0*
09
0>
0C
#8850000000
1!
1*
b110 6
19
1>
1C
b110 G
#8860000000
0!
0*
09
0>
0C
#8870000000
1!
1*
b111 6
19
1>
1C
b111 G
#8880000000
0!
1"
0*
1+
09
1:
0>
0C
#8890000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#8900000000
0!
0*
09
0>
0C
#8910000000
1!
1*
b1 6
19
1>
1C
b1 G
#8920000000
0!
0*
09
0>
0C
#8930000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#8940000000
0!
0*
09
0>
0C
#8950000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#8960000000
0!
0*
09
0>
0C
#8970000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#8980000000
0!
0*
09
0>
0C
#8990000000
1!
1*
b101 6
19
1>
1C
b101 G
#9000000000
0!
0#
0*
0,
09
0>
0?
0C
#9010000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#9020000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#9030000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#9040000000
0!
0*
09
0>
0C
#9050000000
1!
1*
19
1>
1C
#9060000000
0!
0*
09
0>
0C
#9070000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#9080000000
0!
0*
09
0>
0C
#9090000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#9100000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#9110000000
1!
1*
b1 6
19
1>
1C
b1 G
#9120000000
0!
0*
09
0>
0C
#9130000000
1!
1*
b10 6
19
1>
1C
b10 G
#9140000000
0!
0*
09
0>
0C
#9150000000
1!
1*
b11 6
19
1>
1C
b11 G
#9160000000
0!
0*
09
0>
0C
#9170000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#9180000000
0!
0*
09
0>
0C
#9190000000
1!
1*
b101 6
19
1>
1C
b101 G
#9200000000
0!
0*
09
0>
0C
#9210000000
1!
1*
b110 6
19
1>
1C
b110 G
#9220000000
0!
0*
09
0>
0C
#9230000000
1!
1*
b111 6
19
1>
1C
b111 G
#9240000000
0!
0*
09
0>
0C
#9250000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#9260000000
0!
0*
09
0>
0C
#9270000000
1!
1*
b1 6
19
1>
1C
b1 G
#9280000000
0!
0*
09
0>
0C
#9290000000
1!
1*
b10 6
19
1>
1C
b10 G
#9300000000
0!
0*
09
0>
0C
#9310000000
1!
1*
b11 6
19
1>
1C
b11 G
#9320000000
0!
0*
09
0>
0C
#9330000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#9340000000
0!
0*
09
0>
0C
#9350000000
1!
1*
b101 6
19
1>
1C
b101 G
#9360000000
0!
0*
09
0>
0C
#9370000000
1!
1*
b110 6
19
1>
1C
b110 G
#9380000000
0!
0*
09
0>
0C
#9390000000
1!
1*
b111 6
19
1>
1C
b111 G
#9400000000
0!
0*
09
0>
0C
#9410000000
1!
0&
b1101101 '
1*
0/
b1101101 0
b0010 5
b0 6
b10 8
19
1>
1C
0F
b0 G
b1101101 H
b0010 I
#9420000000
0!
0*
09
0>
0C
#9430000000
1!
1*
b1 6
19
1>
1C
b1 G
#9440000000
0!
0*
09
0>
0C
#9450000000
1!
1*
b10 6
19
1>
1C
b10 G
#9460000000
0!
0*
09
0>
0C
#9470000000
1!
1*
b11 6
19
1>
1C
b11 G
#9480000000
0!
0*
09
0>
0C
#9490000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#9500000000
0!
0*
09
0>
0C
#9510000000
1!
1*
b101 6
19
1>
1C
b101 G
#9520000000
0!
0*
09
0>
0C
#9530000000
1!
1*
b110 6
19
1>
1C
b110 G
#9540000000
0!
0*
09
0>
0C
#9550000000
1!
1*
b111 6
19
1>
1C
b111 G
#9560000000
0!
1"
0*
1+
09
1:
0>
0C
#9570000000
1!
0&
b1111001 '
1*
0/
b1111001 0
11
b0011 5
b0 6
b11 8
19
1;
1<
1=
1>
1C
0F
b0 G
b1111001 H
b0011 I
#9580000000
0!
0*
09
0>
0C
#9590000000
1!
1*
b1 6
19
1>
1C
b1 G
#9600000000
0!
0*
09
0>
0C
#9610000000
1!
0"
1*
0+
01
b10 6
19
0:
0;
0<
0=
1>
1C
b10 G
#9620000000
0!
0*
09
0>
0C
#9630000000
1!
1#
1*
1,
12
b11 6
19
1>
1?
1@
1A
1B
1C
b11 G
#9640000000
0!
0*
09
0>
0C
#9650000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#9660000000
0!
0*
09
0>
0C
#9670000000
1!
1*
b101 6
19
1>
1C
b101 G
#9680000000
0!
0#
0*
0,
09
0>
0?
0C
#9690000000
1!
b1111110 '
1*
b1111110 0
02
03
14
b0000 5
b110 6
b0 8
19
1>
0@
0A
0B
1C
1D
0E
b110 G
b1111110 H
b0000 I
#9700000000
0!
0$
1%
0*
0-
1.
09
0>
0C
#9710000000
1!
0&
1*
0/
b0 6
19
1>
1C
0F
b0 G
#9720000000
0!
0*
09
0>
0C
#9730000000
1!
1*
19
1>
1C
#9740000000
0!
0*
09
0>
0C
#9750000000
1!
1"
1*
1+
11
19
1:
1;
1<
1=
1>
1C
#9760000000
0!
0*
09
0>
0C
#9770000000
1!
0"
1*
0+
01
13
04
19
0:
0;
0<
0=
1>
1C
0D
1E
#9780000000
0!
1$
0%
0*
1-
0.
09
0>
0C
#9790000000
1!
1*
b1 6
19
1>
1C
b1 G
#9800000000
0!
0*
09
0>
0C
#9810000000
1!
1*
b10 6
19
1>
1C
b10 G
#9820000000
0!
0*
09
0>
0C
#9830000000
1!
1*
b11 6
19
1>
1C
b11 G
#9840000000
0!
0*
09
0>
0C
#9850000000
1!
1&
1*
1/
b100 6
19
1>
1C
1F
b100 G
#9860000000
0!
0*
09
0>
0C
#9870000000
1!
1*
b101 6
19
1>
1C
b101 G
#9880000000
0!
0*
09
0>
0C
#9890000000
1!
1*
b110 6
19
1>
1C
b110 G
#9900000000
0!
0*
09
0>
0C
#9910000000
1!
1*
b111 6
19
1>
1C
b111 G
#9920000000
0!
0*
09
0>
0C
#9930000000
1!
0&
b0110000 '
1*
0/
b0110000 0
b0001 5
b0 6
b1 8
19
1>
1C
0F
b0 G
b0110000 H
b0001 I
#9940000000
0!
0*
09
0>
0C
#9950000000
1!
1*
b1 6
19
1>
1C
b1 G
#9960000000
0!
0*
09
0>
0C
#9970000000
1!
1*
b10 6
19
1>
1C
b10 G
#9980000000
0!
0*
09
0>
0C
#9990000000
1!
1*
b11 6
19
1>
1C
b11 G
#10000000000
0!
0*
09
0>
0C
