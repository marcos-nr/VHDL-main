$date
  Fri Apr 19 21:55:13 2024
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb_display_cyclone4 $end
$var reg 7 ! seg[6:0] $end
$var reg 4 " bcd[3:0] $end
$var reg 1 # en $end
$scope module uut $end
$var reg 7 $ segmentos[6:0] $end
$var reg 4 % bcd[3:0] $end
$var reg 1 & enable $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
b0000001 !
b0000 "
1#
b0000001 $
b0000 %
1&
#10000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#20000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#30000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#40000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#50000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#60000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#70000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#80000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#90000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#100000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#110000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#120000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#130000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#140000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#150000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#160000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#170000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#180000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#190000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#200000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#210000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#220000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#230000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#240000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#250000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#260000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#270000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#280000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#290000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#300000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#310000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#320000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#330000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#340000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#350000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#360000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#370000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#380000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#390000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#400000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#410000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#420000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#430000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#440000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#450000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#460000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#470000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#480000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#490000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#500000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#510000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#520000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#530000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#540000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#550000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#560000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#570000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#580000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#590000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#600000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#610000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#620000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#630000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#640000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#650000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#660000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#670000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#680000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#690000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#700000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#710000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#720000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#730000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#740000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#750000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#760000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#770000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#780000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#790000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#800000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#810000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#820000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#830000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#840000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#850000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#860000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#870000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#880000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#890000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#900000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#910000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#920000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#930000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#940000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#950000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#960000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#970000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#980000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#990000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#1000000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#1010000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#1020000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#1030000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#1040000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#1050000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#1060000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#1070000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#1080000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#1090000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#1100000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#1110000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#1120000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#1130000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#1140000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#1150000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#1160000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#1170000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#1180000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#1190000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#1200000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#1210000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#1220000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#1230000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#1240000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#1250000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#1260000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#1270000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#1280000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#1290000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#1300000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#1310000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#1320000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#1330000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#1340000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#1350000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#1360000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#1370000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#1380000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#1390000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#1400000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#1410000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#1420000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#1430000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#1440000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#1450000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#1460000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#1470000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#1480000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#1490000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#1500000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#1510000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#1520000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#1530000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#1540000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#1550000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#1560000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#1570000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#1580000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#1590000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#1600000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#1610000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#1620000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#1630000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#1640000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#1650000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#1660000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#1670000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#1680000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#1690000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#1700000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#1710000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#1720000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#1730000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#1740000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#1750000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#1760000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#1770000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#1780000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#1790000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#1800000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#1810000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#1820000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#1830000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#1840000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#1850000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#1860000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#1870000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#1880000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#1890000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#1900000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#1910000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#1920000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#1930000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#1940000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#1950000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#1960000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#1970000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#1980000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#1990000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#2000000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#2010000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#2020000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#2030000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#2040000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#2050000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#2060000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#2070000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#2080000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#2090000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#2100000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#2110000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#2120000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#2130000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#2140000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#2150000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#2160000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#2170000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#2180000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#2190000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#2200000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#2210000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#2220000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#2230000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#2240000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#2250000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#2260000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#2270000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#2280000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#2290000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#2300000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#2310000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#2320000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#2330000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#2340000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#2350000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#2360000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#2370000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#2380000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#2390000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#2400000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#2410000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#2420000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#2430000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#2440000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#2450000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#2460000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#2470000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#2480000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#2490000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#2500000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#2510000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#2520000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#2530000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#2540000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#2550000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#2560000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#2570000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#2580000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#2590000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#2600000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#2610000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#2620000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#2630000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#2640000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#2650000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#2660000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#2670000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#2680000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#2690000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#2700000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#2710000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#2720000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#2730000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#2740000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#2750000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#2760000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#2770000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#2780000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#2790000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#2800000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#2810000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#2820000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#2830000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#2840000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#2850000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#2860000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#2870000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#2880000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#2890000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#2900000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#2910000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#2920000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#2930000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#2940000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#2950000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#2960000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#2970000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#2980000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#2990000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#3000000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#3010000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#3020000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#3030000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#3040000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#3050000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#3060000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#3070000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#3080000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#3090000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#3100000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#3110000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#3120000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#3130000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#3140000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#3150000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#3160000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#3170000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#3180000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#3190000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#3200000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#3210000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#3220000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#3230000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#3240000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#3250000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#3260000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#3270000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#3280000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#3290000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#3300000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#3310000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#3320000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#3330000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#3340000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#3350000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#3360000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#3370000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#3380000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#3390000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#3400000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#3410000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#3420000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#3430000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#3440000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#3450000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#3460000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#3470000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#3480000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#3490000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#3500000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#3510000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#3520000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#3530000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#3540000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#3550000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#3560000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#3570000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#3580000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#3590000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#3600000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#3610000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#3620000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#3630000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#3640000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#3650000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#3660000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#3670000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#3680000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#3690000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#3700000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#3710000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#3720000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#3730000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#3740000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#3750000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#3760000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#3770000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#3780000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#3790000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#3800000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#3810000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#3820000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#3830000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#3840000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#3850000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#3860000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#3870000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#3880000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#3890000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#3900000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#3910000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#3920000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#3930000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#3940000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#3950000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#3960000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#3970000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#3980000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#3990000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#4000000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#4010000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#4020000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#4030000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#4040000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#4050000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#4060000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#4070000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#4080000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#4090000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#4100000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#4110000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#4120000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#4130000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#4140000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#4150000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#4160000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#4170000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#4180000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#4190000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#4200000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#4210000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#4220000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#4230000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#4240000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#4250000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#4260000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#4270000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#4280000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#4290000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#4300000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#4310000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#4320000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#4330000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#4340000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#4350000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#4360000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#4370000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#4380000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#4390000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#4400000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#4410000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#4420000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#4430000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#4440000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#4450000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#4460000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#4470000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#4480000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#4490000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#4500000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#4510000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#4520000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#4530000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#4540000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#4550000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#4560000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#4570000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#4580000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#4590000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#4600000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#4610000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#4620000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#4630000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#4640000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#4650000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#4660000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#4670000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#4680000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#4690000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#4700000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#4710000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#4720000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#4730000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#4740000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#4750000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#4760000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#4770000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#4780000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#4790000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#4800000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#4810000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#4820000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#4830000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#4840000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#4850000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#4860000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#4870000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#4880000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#4890000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#4900000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#4910000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#4920000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#4930000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#4940000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#4950000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#4960000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#4970000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#4980000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#4990000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#5000000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#5010000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#5020000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#5030000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#5040000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#5050000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#5060000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#5070000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#5080000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#5090000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#5100000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#5110000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#5120000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#5130000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#5140000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#5150000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#5160000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#5170000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#5180000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#5190000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#5200000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#5210000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#5220000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#5230000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#5240000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#5250000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#5260000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#5270000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#5280000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#5290000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#5300000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#5310000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#5320000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#5330000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#5340000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#5350000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#5360000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#5370000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#5380000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#5390000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#5400000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#5410000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#5420000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#5430000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#5440000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#5450000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#5460000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#5470000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#5480000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#5490000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#5500000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#5510000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#5520000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#5530000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#5540000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#5550000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#5560000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#5570000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#5580000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#5590000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#5600000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#5610000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#5620000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#5630000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#5640000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#5650000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#5660000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#5670000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#5680000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#5690000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#5700000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#5710000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#5720000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#5730000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#5740000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#5750000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#5760000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#5770000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#5780000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#5790000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#5800000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#5810000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#5820000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#5830000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#5840000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#5850000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#5860000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#5870000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#5880000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#5890000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#5900000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#5910000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#5920000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#5930000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#5940000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#5950000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#5960000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#5970000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#5980000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#5990000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#6000000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#6010000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#6020000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#6030000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#6040000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#6050000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#6060000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#6070000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#6080000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#6090000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#6100000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#6110000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#6120000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#6130000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#6140000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#6150000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#6160000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#6170000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#6180000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#6190000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#6200000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#6210000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#6220000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#6230000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#6240000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#6250000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#6260000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#6270000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#6280000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#6290000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#6300000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#6310000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#6320000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#6330000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#6340000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#6350000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#6360000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#6370000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#6380000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#6390000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#6400000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#6410000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#6420000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#6430000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#6440000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#6450000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#6460000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#6470000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#6480000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#6490000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#6500000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#6510000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#6520000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#6530000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#6540000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#6550000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#6560000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#6570000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#6580000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#6590000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#6600000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#6610000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#6620000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#6630000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#6640000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#6650000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#6660000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#6670000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#6680000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#6690000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#6700000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#6710000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#6720000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#6730000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#6740000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#6750000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#6760000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#6770000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#6780000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#6790000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#6800000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#6810000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#6820000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#6830000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#6840000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#6850000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#6860000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#6870000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#6880000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#6890000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#6900000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#6910000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#6920000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#6930000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#6940000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#6950000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#6960000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#6970000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#6980000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#6990000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#7000000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#7010000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#7020000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#7030000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#7040000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#7050000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#7060000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#7070000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#7080000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#7090000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#7100000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#7110000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#7120000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#7130000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#7140000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#7150000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#7160000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#7170000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#7180000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#7190000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#7200000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#7210000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#7220000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#7230000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#7240000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#7250000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#7260000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#7270000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#7280000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#7290000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#7300000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#7310000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#7320000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#7330000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#7340000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#7350000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#7360000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#7370000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#7380000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#7390000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#7400000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#7410000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#7420000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#7430000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#7440000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#7450000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#7460000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#7470000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#7480000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#7490000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#7500000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#7510000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#7520000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#7530000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#7540000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#7550000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#7560000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#7570000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#7580000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#7590000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#7600000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#7610000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#7620000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#7630000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#7640000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#7650000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#7660000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#7670000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#7680000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#7690000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#7700000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#7710000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#7720000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#7730000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#7740000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#7750000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#7760000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#7770000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#7780000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#7790000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#7800000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#7810000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#7820000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#7830000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#7840000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#7850000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#7860000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#7870000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#7880000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#7890000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#7900000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#7910000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#7920000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#7930000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#7940000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#7950000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#7960000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#7970000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#7980000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#7990000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#8000000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#8010000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#8020000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#8030000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#8040000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#8050000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#8060000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#8070000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#8080000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#8090000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#8100000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#8110000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#8120000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#8130000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#8140000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#8150000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#8160000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#8170000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#8180000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#8190000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#8200000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#8210000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#8220000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#8230000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#8240000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#8250000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#8260000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#8270000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#8280000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#8290000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#8300000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#8310000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#8320000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#8330000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#8340000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#8350000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#8360000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#8370000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#8380000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#8390000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#8400000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#8410000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#8420000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#8430000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#8440000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#8450000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#8460000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#8470000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#8480000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#8490000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#8500000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#8510000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#8520000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#8530000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#8540000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#8550000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#8560000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#8570000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#8580000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#8590000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#8600000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#8610000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#8620000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#8630000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#8640000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#8650000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#8660000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#8670000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#8680000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#8690000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#8700000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#8710000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#8720000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#8730000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#8740000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#8750000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#8760000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#8770000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#8780000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#8790000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#8800000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#8810000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#8820000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#8830000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#8840000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#8850000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#8860000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#8870000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#8880000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#8890000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#8900000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#8910000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#8920000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#8930000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#8940000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#8950000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#8960000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#8970000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#8980000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#8990000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#9000000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#9010000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#9020000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#9030000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#9040000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#9050000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#9060000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#9070000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#9080000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#9090000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#9100000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#9110000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#9120000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#9130000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#9140000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#9150000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#9160000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#9170000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#9180000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#9190000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#9200000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#9210000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#9220000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#9230000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#9240000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#9250000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#9260000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#9270000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#9280000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#9290000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#9300000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#9310000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#9320000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#9330000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#9340000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#9350000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#9360000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#9370000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#9380000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#9390000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#9400000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#9410000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#9420000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#9430000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#9440000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#9450000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#9460000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#9470000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#9480000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#9490000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#9500000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#9510000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#9520000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#9530000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#9540000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#9550000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#9560000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#9570000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#9580000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#9590000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#9600000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#9610000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#9620000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#9630000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#9640000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#9650000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#9660000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#9670000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#9680000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#9690000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#9700000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#9710000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#9720000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#9730000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#9740000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#9750000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#9760000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#9770000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#9780000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#9790000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#9800000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#9810000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#9820000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#9830000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#9840000000
b0000000 !
b1000 "
b0000000 $
b1000 %
#9850000000
b0000100 !
b1001 "
b0000100 $
b1001 %
#9860000000
b0001000 !
b1010 "
b0001000 $
b1010 %
#9870000000
b1100000 !
b1011 "
b1100000 $
b1011 %
#9880000000
b0110001 !
b1100 "
b0110001 $
b1100 %
#9890000000
b1000010 !
b1101 "
b1000010 $
b1101 %
#9900000000
b0110000 !
b1110 "
b0110000 $
b1110 %
#9910000000
b0111000 !
b1111 "
b0111000 $
b1111 %
#9920000000
b0000001 !
b0000 "
b0000001 $
b0000 %
#9930000000
b1001111 !
b0001 "
b1001111 $
b0001 %
#9940000000
b0010010 !
b0010 "
b0010010 $
b0010 %
#9950000000
b0000110 !
b0011 "
b0000110 $
b0011 %
#9960000000
b1001100 !
b0100 "
b1001100 $
b0100 %
#9970000000
b0100100 !
b0101 "
b0100100 $
b0101 %
#9980000000
b0100000 !
b0110 "
b0100000 $
b0110 %
#9990000000
b0001111 !
b0111 "
b0001111 $
b0111 %
#10000000000
b0000000 !
b1000 "
b0000000 $
b1000 %
